

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
         n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
         n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
         n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
         n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
         n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
         n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
         n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
         n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
         n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
         n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
         n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
         n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
         n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
         n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
         n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
         n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487,
         n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
         n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
         n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
         n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
         n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527,
         n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
         n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
         n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
         n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559,
         n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
         n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
         n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583,
         n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
         n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599,
         n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
         n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
         n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
         n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
         n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
         n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
         n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655,
         n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
         n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671,
         n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
         n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
         n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
         n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703,
         n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
         n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
         n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743,
         n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
         n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
         n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
         n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
         n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111,
         n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119,
         n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
         n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135,
         n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
         n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
         n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159,
         n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167,
         n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
         n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183,
         n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191,
         n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199,
         n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207,
         n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215,
         n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223,
         n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231,
         n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
         n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247,
         n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255,
         n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263,
         n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
         n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279,
         n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287,
         n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295,
         n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303,
         n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311,
         n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319,
         n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327,
         n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335,
         n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343,
         n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351,
         n21352, n21353, n21354, n21355;

  OR2_X1 U11032 ( .A1(n19988), .A2(n20030), .ZN(n20152) );
  NAND2_X1 U11033 ( .A1(n13505), .A2(n13504), .ZN(n20102) );
  INV_X2 U11034 ( .A(n18228), .ZN(n10304) );
  INV_X1 U11035 ( .A(n21355), .ZN(n9613) );
  CLKBUF_X2 U11037 ( .A(n11741), .Z(n10064) );
  AND2_X1 U11038 ( .A1(n13517), .A2(n20104), .ZN(n12045) );
  CLKBUF_X2 U11039 ( .A(n12833), .Z(n9590) );
  CLKBUF_X2 U11040 ( .A(n12787), .Z(n14270) );
  OAI211_X2 U11041 ( .C1(n12371), .C2(n12543), .A(n9908), .B(n12392), .ZN(
        n12395) );
  CLKBUF_X2 U11042 ( .A(n12369), .Z(n12543) );
  NAND2_X1 U11043 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18339) );
  AND2_X1 U11044 ( .A1(n11763), .A2(n10422), .ZN(n13913) );
  AND2_X1 U11045 ( .A1(n11448), .A2(n10811), .ZN(n10851) );
  NAND4_X1 U11046 ( .A1(n10826), .A2(n11442), .A3(n10816), .A4(n14008), .ZN(
        n13454) );
  OR2_X1 U11047 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12619) );
  AND2_X2 U11048 ( .A1(n9605), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11662) );
  BUF_X1 U11049 ( .A(n11777), .Z(n12008) );
  AND2_X1 U11050 ( .A1(n11579), .A2(n14443), .ZN(n14470) );
  AND2_X2 U11051 ( .A1(n14454), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11612) );
  AND2_X1 U11052 ( .A1(n11581), .A2(n11582), .ZN(n14472) );
  INV_X1 U11053 ( .A(n14010), .ZN(n10837) );
  BUF_X1 U11054 ( .A(n10819), .Z(n13722) );
  CLKBUF_X1 U11055 ( .A(n10823), .Z(n20524) );
  AND4_X1 U11056 ( .A1(n10754), .A2(n10753), .A3(n10752), .A4(n10751), .ZN(
        n10766) );
  BUF_X2 U11057 ( .A(n11732), .Z(n14601) );
  CLKBUF_X2 U11058 ( .A(n10804), .Z(n13140) );
  CLKBUF_X2 U11060 ( .A(n10804), .Z(n11310) );
  BUF_X2 U11061 ( .A(n10705), .Z(n11286) );
  AND2_X1 U11062 ( .A1(n13485), .A2(n10606), .ZN(n10732) );
  AND2_X1 U11063 ( .A1(n10465), .A2(n13457), .ZN(n10683) );
  AND2_X1 U11064 ( .A1(n10465), .A2(n10607), .ZN(n10625) );
  AND4_X1 U11065 ( .A1(n10225), .A2(n9816), .A3(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A4(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9619) );
  AND2_X1 U11067 ( .A1(n10225), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10606) );
  INV_X1 U11068 ( .A(n19545), .ZN(n11803) );
  INV_X1 U11069 ( .A(n16778), .ZN(n11773) );
  NAND2_X1 U11070 ( .A1(n19325), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12618) );
  INV_X1 U11071 ( .A(n12786), .ZN(n17489) );
  INV_X1 U11072 ( .A(n17732), .ZN(n12627) );
  NAND2_X1 U11073 ( .A1(n11434), .A2(n13722), .ZN(n10820) );
  NOR2_X1 U11074 ( .A1(n9614), .A2(n14671), .ZN(n11548) );
  INV_X1 U11075 ( .A(n21355), .ZN(n9614) );
  INV_X2 U11077 ( .A(n12193), .ZN(n12559) );
  NOR2_X1 U11078 ( .A1(n13084), .A2(n15815), .ZN(n13086) );
  INV_X1 U11079 ( .A(n17736), .ZN(n17684) );
  OR2_X1 U11080 ( .A1(n18342), .A2(n9807), .ZN(n9982) );
  CLKBUF_X2 U11081 ( .A(n12833), .Z(n9591) );
  BUF_X1 U11082 ( .A(n12833), .Z(n9592) );
  AND2_X1 U11083 ( .A1(n14718), .A2(n10498), .ZN(n13293) );
  NAND2_X1 U11084 ( .A1(n10823), .A2(n10819), .ZN(n11390) );
  NOR2_X1 U11085 ( .A1(n13075), .A2(n21303), .ZN(n13074) );
  AND2_X1 U11086 ( .A1(n11863), .A2(n11871), .ZN(n16774) );
  NOR2_X1 U11087 ( .A1(n18044), .A2(n17146), .ZN(n17145) );
  INV_X1 U11088 ( .A(n17470), .ZN(n17481) );
  INV_X2 U11089 ( .A(n17434), .ZN(n10321) );
  NAND2_X1 U11090 ( .A1(n13524), .A2(n11777), .ZN(n11794) );
  INV_X1 U11091 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20104) );
  NOR2_X1 U11092 ( .A1(n12727), .A2(n12731), .ZN(n17462) );
  INV_X1 U11093 ( .A(n18248), .ZN(n18293) );
  NAND2_X1 U11094 ( .A1(n16805), .A2(n18381), .ZN(n18374) );
  NOR2_X1 U11095 ( .A1(n17972), .A2(n17104), .ZN(n18371) );
  INV_X2 U11096 ( .A(n20375), .ZN(n20358) );
  OR2_X1 U11097 ( .A1(n13725), .A2(n13724), .ZN(n20481) );
  AOI211_X1 U11098 ( .C1(n19414), .C2(n15607), .A(n15606), .B(n15605), .ZN(
        n15608) );
  INV_X2 U11099 ( .A(n20284), .ZN(n20287) );
  NAND2_X1 U11100 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17485), .ZN(n17471) );
  NOR2_X1 U11101 ( .A1(n12782), .A2(n12781), .ZN(n17916) );
  AOI21_X1 U11102 ( .B1(n18371), .B2(n18544), .A(n10294), .ZN(n18283) );
  NOR2_X1 U11103 ( .A1(n10181), .A2(n13275), .ZN(n16826) );
  OR2_X1 U11104 ( .A1(n14229), .A2(n17466), .ZN(n9588) );
  INV_X1 U11105 ( .A(n12812), .ZN(n17736) );
  OR2_X1 U11106 ( .A1(n11838), .A2(n13702), .ZN(n9589) );
  INV_X4 U11107 ( .A(n17489), .ZN(n17643) );
  NAND3_X2 U11109 ( .A1(n18071), .A2(n18061), .A3(n10305), .ZN(n18045) );
  OAI211_X2 U11110 ( .C1(n18413), .C2(n10281), .A(n10169), .B(n10171), .ZN(
        n18061) );
  NAND2_X2 U11111 ( .A1(n12710), .A2(n12709), .ZN(n17466) );
  NAND2_X4 U11112 ( .A1(n9948), .A2(n9947), .ZN(n16267) );
  AND4_X2 U11113 ( .A1(n10693), .A2(n10692), .A3(n10691), .A4(n10690), .ZN(
        n10581) );
  NAND2_X2 U11114 ( .A1(n13968), .A2(n11929), .ZN(n11931) );
  NAND2_X4 U11115 ( .A1(n10581), .A2(n10698), .ZN(n10818) );
  NAND2_X2 U11116 ( .A1(n10049), .A2(n10047), .ZN(n11810) );
  NOR2_X1 U11117 ( .A1(n17466), .A2(n12618), .ZN(n12833) );
  CLKBUF_X1 U11118 ( .A(n10624), .Z(n9593) );
  AND2_X1 U11119 ( .A1(n10465), .A2(n13485), .ZN(n10624) );
  CLKBUF_X1 U11120 ( .A(n10624), .Z(n13139) );
  AND2_X4 U11121 ( .A1(n13166), .A2(n13165), .ZN(n10583) );
  NOR2_X1 U11122 ( .A1(n10167), .A2(n12619), .ZN(n9594) );
  NOR2_X2 U11123 ( .A1(n10167), .A2(n12619), .ZN(n17676) );
  INV_X1 U11124 ( .A(n17676), .ZN(n12835) );
  AOI21_X2 U11125 ( .B1(n11840), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11834), .ZN(n12202) );
  INV_X4 U11126 ( .A(n12627), .ZN(n17719) );
  XNOR2_X2 U11127 ( .A(n11827), .B(n11829), .ZN(n11853) );
  NAND2_X2 U11128 ( .A1(n11704), .A2(n11703), .ZN(n19545) );
  XNOR2_X2 U11129 ( .A(n11999), .B(n12048), .ZN(n16417) );
  BUF_X1 U11130 ( .A(n12803), .Z(n9595) );
  MUX2_X1 U11131 ( .A(n14342), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n9596) );
  NOR2_X2 U11132 ( .A1(n12619), .A2(n12617), .ZN(n12752) );
  XNOR2_X1 U11133 ( .A(n9888), .B(n16205), .ZN(n16464) );
  NAND2_X1 U11134 ( .A1(n9970), .A2(n9685), .ZN(n16574) );
  XNOR2_X1 U11135 ( .A(n16194), .B(n16192), .ZN(n16191) );
  NOR2_X1 U11136 ( .A1(n16342), .A2(n16591), .ZN(n16343) );
  AOI21_X1 U11137 ( .B1(n10203), .B2(n10202), .A(n10201), .ZN(n12990) );
  OAI21_X1 U11138 ( .B1(n16229), .B2(n10547), .A(n10217), .ZN(n10220) );
  AND2_X1 U11139 ( .A1(n9904), .A2(n9903), .ZN(n16229) );
  OAI21_X1 U11140 ( .B1(n13276), .B2(n9780), .A(n12930), .ZN(n16888) );
  NAND2_X1 U11141 ( .A1(n9716), .A2(n10157), .ZN(n9866) );
  OR2_X1 U11142 ( .A1(n9720), .A2(n9910), .ZN(n10199) );
  OR2_X1 U11143 ( .A1(n10596), .A2(n10595), .ZN(n14003) );
  OAI21_X1 U11144 ( .B1(n10228), .B2(n13645), .A(n13210), .ZN(n13211) );
  NAND3_X1 U11145 ( .A1(n10541), .A2(n11920), .A3(n13967), .ZN(n13968) );
  CLKBUF_X1 U11146 ( .A(n14975), .Z(n15020) );
  OR2_X1 U11147 ( .A1(n16455), .A2(n12361), .ZN(n13000) );
  INV_X4 U11148 ( .A(n10583), .ZN(n15236) );
  NAND2_X1 U11149 ( .A1(n10060), .A2(n11020), .ZN(n15560) );
  INV_X2 U11150 ( .A(n16929), .ZN(n15241) );
  OR2_X1 U11151 ( .A1(n12463), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12452) );
  NAND2_X1 U11152 ( .A1(n20293), .A2(n13256), .ZN(n16937) );
  INV_X2 U11153 ( .A(n18140), .ZN(n18239) );
  AND2_X1 U11154 ( .A1(n12465), .A2(n9762), .ZN(n12460) );
  INV_X1 U11155 ( .A(n11906), .ZN(n19530) );
  NAND2_X1 U11156 ( .A1(n12465), .A2(n12464), .ZN(n12463) );
  NAND2_X4 U11157 ( .A1(n9798), .A2(n11871), .ZN(n11904) );
  NAND2_X1 U11158 ( .A1(n12478), .A2(n12522), .ZN(n12465) );
  NAND2_X1 U11159 ( .A1(n11876), .A2(n11871), .ZN(n11906) );
  AND2_X1 U11160 ( .A1(n14937), .A2(n14936), .ZN(n14939) );
  OAI21_X2 U11161 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19352), .A(n17104), 
        .ZN(n18381) );
  NAND2_X4 U11162 ( .A1(n12443), .A2(n12522), .ZN(n12482) );
  INV_X1 U11163 ( .A(n13518), .ZN(n9836) );
  NAND2_X1 U11164 ( .A1(n10124), .A2(n11854), .ZN(n11852) );
  INV_X2 U11165 ( .A(n18703), .ZN(n19184) );
  NAND2_X1 U11166 ( .A1(n12385), .A2(n12386), .ZN(n12384) );
  NOR2_X2 U11167 ( .A1(n12390), .A2(n12395), .ZN(n12385) );
  INV_X2 U11168 ( .A(n12189), .ZN(n12003) );
  NOR2_X2 U11169 ( .A1(n17916), .A2(n12852), .ZN(n12854) );
  NAND2_X1 U11170 ( .A1(n11794), .A2(n19553), .ZN(n11782) );
  NAND2_X1 U11171 ( .A1(n20520), .A2(n20532), .ZN(n9821) );
  NAND2_X1 U11172 ( .A1(n11787), .A2(n13517), .ZN(n11793) );
  INV_X2 U11173 ( .A(n11800), .ZN(n11780) );
  NAND2_X1 U11174 ( .A1(n9667), .A2(n12810), .ZN(n17922) );
  NOR2_X1 U11175 ( .A1(n14561), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12009) );
  CLKBUF_X1 U11176 ( .A(n11810), .Z(n19566) );
  NAND2_X1 U11177 ( .A1(n20532), .A2(n10818), .ZN(n13318) );
  NAND2_X2 U11178 ( .A1(n14561), .A2(n16778), .ZN(n11800) );
  NAND2_X2 U11179 ( .A1(n10093), .A2(n10091), .ZN(n14561) );
  OR2_X2 U11180 ( .A1(n10742), .A2(n10741), .ZN(n20532) );
  CLKBUF_X2 U11181 ( .A(n11890), .Z(n12122) );
  BUF_X2 U11183 ( .A(n10759), .Z(n13138) );
  BUF_X2 U11184 ( .A(n10700), .Z(n11246) );
  BUF_X2 U11185 ( .A(n10625), .Z(n13146) );
  BUF_X2 U11186 ( .A(n10705), .Z(n13149) );
  AND2_X1 U11187 ( .A1(n10607), .A2(n15518), .ZN(n10672) );
  CLKBUF_X3 U11188 ( .A(n11732), .Z(n14607) );
  AND2_X2 U11189 ( .A1(n14447), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11676) );
  CLKBUF_X1 U11190 ( .A(n14610), .Z(n14598) );
  CLKBUF_X2 U11191 ( .A(n9619), .Z(n10646) );
  BUF_X4 U11192 ( .A(n12639), .Z(n9597) );
  BUF_X2 U11193 ( .A(n10883), .Z(n13147) );
  AND3_X1 U11194 ( .A1(n15524), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n16848), .ZN(n10773) );
  CLKBUF_X1 U11195 ( .A(n11580), .Z(n13887) );
  NOR2_X4 U11196 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13485) );
  INV_X2 U11197 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11564) );
  OAI21_X1 U11198 ( .B1(n10044), .B2(n15236), .A(n9825), .ZN(n15050) );
  OR2_X1 U11199 ( .A1(n12989), .A2(n12988), .ZN(n16190) );
  AOI21_X1 U11200 ( .B1(n9834), .B2(n16383), .A(n9711), .ZN(n16260) );
  AND2_X1 U11201 ( .A1(n10080), .A2(n10078), .ZN(n10077) );
  AOI21_X1 U11202 ( .B1(n16574), .B2(n16576), .A(n9882), .ZN(n16575) );
  AOI21_X1 U11203 ( .B1(n10214), .B2(n16426), .A(n10212), .ZN(n16201) );
  AOI21_X1 U11204 ( .B1(n10214), .B2(n16689), .A(n16451), .ZN(n16452) );
  AND2_X1 U11205 ( .A1(n9803), .A2(n9802), .ZN(n9834) );
  AND2_X1 U11206 ( .A1(n10538), .A2(n10540), .ZN(n16285) );
  AND2_X1 U11207 ( .A1(n9952), .A2(n9950), .ZN(n12988) );
  NAND2_X1 U11208 ( .A1(n15086), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13251) );
  AND2_X1 U11209 ( .A1(n15080), .A2(n15303), .ZN(n10044) );
  XNOR2_X1 U11210 ( .A(n13296), .B(n13295), .ZN(n14650) );
  INV_X1 U11211 ( .A(n10254), .ZN(n9952) );
  AND3_X1 U11212 ( .A1(n9789), .A2(n13250), .A3(n15107), .ZN(n15080) );
  XNOR2_X1 U11213 ( .A(n13293), .B(n10136), .ZN(n10397) );
  NAND2_X1 U11214 ( .A1(n16343), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16316) );
  AND2_X1 U11215 ( .A1(n10165), .A2(n9793), .ZN(n16310) );
  NAND2_X1 U11216 ( .A1(n13250), .A2(n15107), .ZN(n15099) );
  NOR2_X1 U11217 ( .A1(n12990), .A2(n12992), .ZN(n12582) );
  NAND2_X1 U11218 ( .A1(n15106), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13250) );
  AND2_X1 U11219 ( .A1(n14328), .A2(n14327), .ZN(n16354) );
  CLKBUF_X1 U11220 ( .A(n16400), .Z(n16401) );
  NAND2_X1 U11221 ( .A1(n10336), .A2(n16361), .ZN(n14327) );
  NAND2_X1 U11222 ( .A1(n10334), .A2(n16362), .ZN(n14328) );
  NAND2_X1 U11223 ( .A1(n12515), .A2(n12514), .ZN(n16222) );
  NAND2_X1 U11224 ( .A1(n16364), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10334) );
  NAND2_X1 U11225 ( .A1(n9958), .A2(n9955), .ZN(n16451) );
  NAND2_X1 U11226 ( .A1(n9928), .A2(n13236), .ZN(n9935) );
  NAND2_X1 U11227 ( .A1(n9866), .A2(n10385), .ZN(n16364) );
  AOI21_X1 U11228 ( .B1(n15287), .B2(n9876), .A(n9874), .ZN(n15291) );
  AND2_X1 U11229 ( .A1(n13041), .A2(n13040), .ZN(n13042) );
  OR2_X2 U11230 ( .A1(n14353), .A2(n14016), .ZN(n16908) );
  NOR2_X1 U11231 ( .A1(n9957), .A2(n9956), .ZN(n9955) );
  OR2_X1 U11232 ( .A1(n14110), .A2(n14902), .ZN(n14905) );
  NAND2_X1 U11233 ( .A1(n9875), .A2(n15289), .ZN(n9874) );
  AND2_X1 U11234 ( .A1(n9907), .A2(n10567), .ZN(n10385) );
  NOR2_X1 U11235 ( .A1(n18045), .A2(n18228), .ZN(n13027) );
  AND2_X1 U11236 ( .A1(n9949), .A2(n16403), .ZN(n9676) );
  AND2_X1 U11237 ( .A1(n11932), .A2(n10252), .ZN(n9848) );
  AND2_X1 U11238 ( .A1(n16417), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11998) );
  OR2_X1 U11239 ( .A1(n10281), .A2(n9979), .ZN(n9972) );
  CLKBUF_X1 U11240 ( .A(n13963), .Z(n14149) );
  NAND2_X1 U11241 ( .A1(n10281), .A2(n10284), .ZN(n12870) );
  NAND2_X1 U11242 ( .A1(n9799), .A2(n10028), .ZN(n9850) );
  OR2_X1 U11243 ( .A1(n12534), .A2(n12533), .ZN(n12547) );
  XNOR2_X1 U11244 ( .A(n13211), .B(n16979), .ZN(n16932) );
  NAND3_X1 U11245 ( .A1(n9902), .A2(n9901), .A3(n10256), .ZN(n12411) );
  NAND2_X1 U11246 ( .A1(n10282), .A2(n9809), .ZN(n10281) );
  NOR2_X1 U11247 ( .A1(n10216), .A2(n10215), .ZN(n16250) );
  AOI21_X1 U11248 ( .B1(n10258), .B2(n10028), .A(n19407), .ZN(n9901) );
  AOI221_X1 U11249 ( .B1(n18178), .B2(n18105), .C1(n18453), .C2(n18105), .A(
        n18133), .ZN(n18106) );
  NAND2_X1 U11250 ( .A1(n12383), .A2(n10258), .ZN(n10256) );
  NAND2_X1 U11251 ( .A1(n11006), .A2(n11005), .ZN(n13784) );
  AND3_X2 U11252 ( .A1(n11973), .A2(n12367), .A3(n11979), .ZN(n11999) );
  NOR2_X1 U11253 ( .A1(n9637), .A2(n10033), .ZN(n10240) );
  NOR2_X1 U11254 ( .A1(n12368), .A2(n12412), .ZN(n10258) );
  INV_X1 U11255 ( .A(n10028), .ZN(n11973) );
  NAND2_X1 U11256 ( .A1(n10089), .A2(n9809), .ZN(n10170) );
  NAND2_X1 U11257 ( .A1(n18544), .A2(n10179), .ZN(n18523) );
  AND2_X1 U11258 ( .A1(n19213), .A2(n10272), .ZN(n19207) );
  NAND2_X1 U11259 ( .A1(n15216), .A2(n13232), .ZN(n15247) );
  NAND2_X1 U11260 ( .A1(n10384), .A2(n11972), .ZN(n12368) );
  NAND2_X1 U11261 ( .A1(n9801), .A2(n9847), .ZN(n10028) );
  OR2_X1 U11262 ( .A1(n15236), .A2(n15429), .ZN(n15179) );
  OAI211_X1 U11263 ( .C1(n13213), .C2(n11189), .A(n11047), .B(n11046), .ZN(
        n14125) );
  AND2_X1 U11264 ( .A1(n10276), .A2(n10273), .ZN(n19213) );
  NAND2_X1 U11265 ( .A1(n18189), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18514) );
  NOR2_X1 U11266 ( .A1(n18168), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18167) );
  AND2_X1 U11267 ( .A1(n10178), .A2(n12866), .ZN(n18178) );
  NAND2_X1 U11268 ( .A1(n9846), .A2(n11953), .ZN(n12383) );
  AND2_X1 U11269 ( .A1(n12453), .A2(n12452), .ZN(n15743) );
  NAND2_X1 U11270 ( .A1(n9858), .A2(n9857), .ZN(n13169) );
  CLKBUF_X1 U11271 ( .A(n15556), .Z(n15562) );
  NAND2_X1 U11272 ( .A1(n10000), .A2(n12911), .ZN(n18285) );
  OAI211_X1 U11273 ( .C1(n18292), .C2(n18512), .A(n10176), .B(n12866), .ZN(
        n18168) );
  XNOR2_X1 U11274 ( .A(n13166), .B(n11051), .ZN(n14126) );
  INV_X1 U11275 ( .A(n10177), .ZN(n10176) );
  AOI22_X1 U11276 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19828), .B1(
        n16774), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11912) );
  AOI22_X1 U11277 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19727), .B1(
        n11956), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11909) );
  NOR2_X1 U11278 ( .A1(n10295), .A2(n12890), .ZN(n10294) );
  INV_X1 U11279 ( .A(n19630), .ZN(n19627) );
  INV_X1 U11280 ( .A(n11913), .ZN(n19587) );
  NAND2_X1 U11281 ( .A1(n9822), .A2(n10948), .ZN(n10949) );
  NAND2_X1 U11282 ( .A1(n14939), .A2(n9702), .ZN(n14875) );
  NAND2_X1 U11283 ( .A1(n11876), .A2(n11879), .ZN(n19630) );
  NAND2_X1 U11284 ( .A1(n15517), .A2(n10144), .ZN(n9822) );
  INV_X1 U11285 ( .A(n10394), .ZN(n18301) );
  NAND2_X1 U11286 ( .A1(n10395), .A2(n10394), .ZN(n18261) );
  NAND2_X1 U11287 ( .A1(n11876), .A2(n11875), .ZN(n11913) );
  CLKBUF_X1 U11288 ( .A(n15517), .Z(n20774) );
  NAND2_X1 U11289 ( .A1(n11863), .A2(n11879), .ZN(n20043) );
  NAND2_X1 U11290 ( .A1(n18312), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18311) );
  AND2_X1 U11291 ( .A1(n10306), .A2(n10321), .ZN(n17199) );
  NAND2_X1 U11292 ( .A1(n9880), .A2(n11433), .ZN(n16883) );
  XNOR2_X1 U11293 ( .A(n15542), .B(n20644), .ZN(n15517) );
  NOR2_X1 U11294 ( .A1(n15506), .A2(n14112), .ZN(n14937) );
  NAND2_X1 U11295 ( .A1(n10035), .A2(n10864), .ZN(n15542) );
  XNOR2_X1 U11296 ( .A(n13193), .B(n13189), .ZN(n20570) );
  NOR2_X1 U11297 ( .A1(n13120), .A2(n10365), .ZN(n13062) );
  XNOR2_X1 U11298 ( .A(n12908), .B(n10339), .ZN(n18312) );
  NAND3_X1 U11299 ( .A1(n11861), .A2(n11860), .A3(n11859), .ZN(n13703) );
  NAND2_X1 U11300 ( .A1(n19353), .A2(n19202), .ZN(n17104) );
  AND2_X1 U11301 ( .A1(n9988), .A2(n9987), .ZN(n12864) );
  INV_X2 U11302 ( .A(n16058), .ZN(n9598) );
  OAI21_X1 U11303 ( .B1(n13518), .B2(n13630), .A(n13498), .ZN(n13525) );
  XNOR2_X1 U11304 ( .A(n9844), .B(n11852), .ZN(n16714) );
  NAND2_X1 U11305 ( .A1(n18326), .A2(n12906), .ZN(n12908) );
  NAND2_X1 U11306 ( .A1(n10982), .A2(n10981), .ZN(n13193) );
  NAND2_X1 U11307 ( .A1(n11852), .A2(n10125), .ZN(n13518) );
  CLKBUF_X1 U11308 ( .A(n10985), .Z(n20606) );
  NAND2_X1 U11309 ( .A1(n9624), .A2(n9811), .ZN(n9810) );
  NOR2_X1 U11310 ( .A1(n9923), .A2(n10864), .ZN(n10865) );
  AOI21_X2 U11311 ( .B1(n11770), .B2(n11769), .A(n19381), .ZN(n12554) );
  NAND3_X1 U11312 ( .A1(n9997), .A2(n18328), .A3(n9998), .ZN(n18326) );
  AND2_X1 U11313 ( .A1(n10863), .A2(n10144), .ZN(n10137) );
  INV_X2 U11314 ( .A(n17950), .ZN(n17963) );
  AND2_X1 U11315 ( .A1(n9936), .A2(n10894), .ZN(n10880) );
  OR2_X1 U11316 ( .A1(n11829), .A2(n11828), .ZN(n11830) );
  NOR2_X1 U11317 ( .A1(n11488), .A2(n10479), .ZN(n10478) );
  XNOR2_X1 U11318 ( .A(n9851), .B(n11843), .ZN(n11850) );
  NAND2_X1 U11319 ( .A1(n13787), .A2(n13786), .ZN(n16974) );
  NAND2_X1 U11320 ( .A1(n11826), .A2(n11825), .ZN(n11829) );
  AND2_X1 U11321 ( .A1(n13755), .A2(n13754), .ZN(n13787) );
  OAI211_X1 U11322 ( .C1(n12218), .C2(n13634), .A(n11833), .B(n11832), .ZN(
        n12204) );
  NOR2_X1 U11323 ( .A1(n16972), .A2(n16973), .ZN(n11481) );
  NAND2_X1 U11324 ( .A1(n12378), .A2(n12377), .ZN(n12407) );
  NAND3_X1 U11325 ( .A1(n11837), .A2(n11836), .A3(n9589), .ZN(n9851) );
  NOR2_X1 U11326 ( .A1(n14232), .A2(n10270), .ZN(n19167) );
  AND2_X1 U11327 ( .A1(n11480), .A2(n11479), .ZN(n16973) );
  NAND2_X1 U11328 ( .A1(n12876), .A2(n17973), .ZN(n14232) );
  NAND2_X2 U11329 ( .A1(n13029), .A2(n12862), .ZN(n18228) );
  INV_X1 U11330 ( .A(n11555), .ZN(n11556) );
  CLKBUF_X1 U11331 ( .A(n12209), .Z(n12302) );
  OAI21_X1 U11332 ( .B1(n12328), .B2(n11803), .A(n12330), .ZN(n11784) );
  MUX2_X1 U11333 ( .A(n12374), .B(n13702), .S(n12543), .Z(n12386) );
  AND2_X1 U11334 ( .A1(n11776), .A2(n11775), .ZN(n13884) );
  AND2_X2 U11335 ( .A1(n11823), .A2(n11801), .ZN(n12230) );
  NAND3_X1 U11336 ( .A1(n10062), .A2(n11782), .A3(n19577), .ZN(n12328) );
  NAND4_X1 U11337 ( .A1(n12886), .A2(n12697), .A3(n12702), .A4(n17424), .ZN(
        n17973) );
  OAI211_X1 U11338 ( .C1(n11416), .C2(n10922), .A(n10921), .B(n10920), .ZN(
        n13189) );
  AND2_X1 U11339 ( .A1(n12850), .A2(n9999), .ZN(n12898) );
  XNOR2_X1 U11340 ( .A(n12852), .B(n17916), .ZN(n18353) );
  INV_X1 U11341 ( .A(n11808), .ZN(n11823) );
  CLKBUF_X1 U11342 ( .A(n11812), .Z(n13911) );
  OAI21_X1 U11343 ( .B1(n11783), .B2(n13913), .A(n11808), .ZN(n10090) );
  NAND2_X1 U11344 ( .A1(n13318), .A2(n9821), .ZN(n10826) );
  OR2_X1 U11345 ( .A1(n11762), .A2(n19553), .ZN(n10062) );
  NAND2_X2 U11346 ( .A1(n13534), .A2(n12009), .ZN(n12189) );
  NAND3_X1 U11348 ( .A1(n11763), .A2(n13534), .A3(n13524), .ZN(n11808) );
  CLKBUF_X1 U11349 ( .A(n10843), .Z(n14647) );
  OR2_X1 U11350 ( .A1(n11587), .A2(n11588), .ZN(n10211) );
  NAND4_X2 U11351 ( .A1(n11995), .A2(n11994), .A3(n11993), .A4(n11992), .ZN(
        n12412) );
  AND3_X1 U11352 ( .A1(n11778), .A2(n12369), .A3(n11810), .ZN(n11787) );
  NAND3_X1 U11353 ( .A1(n12666), .A2(n12665), .A3(n12664), .ZN(n18732) );
  NAND3_X1 U11354 ( .A1(n12687), .A2(n12686), .A3(n12685), .ZN(n18745) );
  AND2_X1 U11355 ( .A1(n11741), .A2(n16778), .ZN(n13928) );
  INV_X1 U11356 ( .A(n17785), .ZN(n18749) );
  INV_X1 U11357 ( .A(n20512), .ZN(n11436) );
  INV_X2 U11358 ( .A(n17035), .ZN(n17063) );
  INV_X1 U11359 ( .A(n11810), .ZN(n13524) );
  BUF_X2 U11360 ( .A(n11438), .Z(n20516) );
  OR2_X1 U11361 ( .A1(n10905), .A2(n10904), .ZN(n13229) );
  INV_X1 U11362 ( .A(n14561), .ZN(n11741) );
  AND4_X1 U11363 ( .A1(n12801), .A2(n12800), .A3(n12799), .A4(n12798), .ZN(
        n12810) );
  AND4_X1 U11364 ( .A1(n10795), .A2(n10794), .A3(n10793), .A4(n10792), .ZN(
        n10796) );
  AND4_X1 U11365 ( .A1(n10790), .A2(n10789), .A3(n10788), .A4(n10787), .ZN(
        n10797) );
  AND4_X1 U11367 ( .A1(n10719), .A2(n10718), .A3(n10717), .A4(n10716), .ZN(
        n10730) );
  AND4_X1 U11368 ( .A1(n10723), .A2(n10722), .A3(n10721), .A4(n10720), .ZN(
        n10729) );
  AND4_X1 U11369 ( .A1(n10772), .A2(n10771), .A3(n10770), .A4(n10769), .ZN(
        n10778) );
  AND4_X1 U11370 ( .A1(n10697), .A2(n10696), .A3(n10695), .A4(n10694), .ZN(
        n10698) );
  AND4_X1 U11371 ( .A1(n10786), .A2(n10785), .A3(n10784), .A4(n10783), .ZN(
        n10798) );
  AND4_X1 U11372 ( .A1(n10763), .A2(n10762), .A3(n10761), .A4(n10760), .ZN(
        n10764) );
  INV_X1 U11373 ( .A(n9588), .ZN(n9610) );
  INV_X2 U11374 ( .A(n9588), .ZN(n9609) );
  NOR2_X2 U11375 ( .A1(n20492), .A2(n20491), .ZN(n20493) );
  INV_X2 U11376 ( .A(n12678), .ZN(n17733) );
  INV_X1 U11377 ( .A(n9588), .ZN(n9611) );
  BUF_X2 U11378 ( .A(n10672), .Z(n10799) );
  INV_X1 U11379 ( .A(n12822), .ZN(n17714) );
  AND2_X2 U11380 ( .A1(n14607), .A2(n11839), .ZN(n14463) );
  NOR2_X1 U11381 ( .A1(n17340), .A2(n17330), .ZN(n18252) );
  CLKBUF_X1 U11382 ( .A(n13140), .Z(n11227) );
  INV_X2 U11383 ( .A(n17090), .ZN(U215) );
  BUF_X2 U11384 ( .A(n9595), .Z(n17734) );
  CLKBUF_X3 U11385 ( .A(n12752), .Z(n17570) );
  BUF_X2 U11386 ( .A(n9595), .Z(n12836) );
  BUF_X2 U11387 ( .A(n10683), .Z(n11281) );
  AND2_X1 U11388 ( .A1(n11726), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11728) );
  AND2_X1 U11389 ( .A1(n11734), .A2(n11839), .ZN(n11735) );
  NOR2_X1 U11390 ( .A1(n10167), .A2(n12620), .ZN(n12787) );
  INV_X2 U11391 ( .A(n17092), .ZN(n17095) );
  AND2_X2 U11392 ( .A1(n10605), .A2(n15518), .ZN(n10699) );
  BUF_X2 U11393 ( .A(n10773), .Z(n9607) );
  BUF_X4 U11394 ( .A(n10773), .Z(n9608) );
  NOR2_X1 U11395 ( .A1(n10997), .A2(n10584), .ZN(n10998) );
  AND2_X2 U11396 ( .A1(n11581), .A2(n11630), .ZN(n14610) );
  NAND2_X1 U11397 ( .A1(n12710), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10167) );
  NAND2_X1 U11398 ( .A1(n12709), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12617) );
  NAND2_X1 U11399 ( .A1(n17437), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12620) );
  NOR2_X1 U11400 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10600), .ZN(
        n10605) );
  NAND3_X2 U11401 ( .A1(n19330), .A2(n19215), .A3(n18707), .ZN(n18701) );
  NOR2_X1 U11402 ( .A1(n13066), .A2(n13069), .ZN(n13068) );
  AND2_X1 U11403 ( .A1(n9922), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10465) );
  AND2_X1 U11404 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15524) );
  INV_X2 U11405 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16848) );
  INV_X2 U11406 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12710) );
  INV_X1 U11407 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n9601) );
  AND2_X1 U11408 ( .A1(n9602), .A2(n9968), .ZN(n16360) );
  NOR2_X1 U11409 ( .A1(n10363), .A2(n9601), .ZN(n9602) );
  NAND2_X1 U11410 ( .A1(n11880), .A2(n11879), .ZN(n19755) );
  NAND2_X1 U11411 ( .A1(n11606), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10359) );
  AND2_X1 U11412 ( .A1(n9798), .A2(n11879), .ZN(n9621) );
  NAND2_X1 U11413 ( .A1(n10358), .A2(n11800), .ZN(n12320) );
  NAND2_X1 U11414 ( .A1(n11810), .A2(n11777), .ZN(n11786) );
  NOR2_X2 U11415 ( .A1(n12619), .A2(n17466), .ZN(n12812) );
  AND2_X1 U11416 ( .A1(n10457), .A2(n11564), .ZN(n9603) );
  AND2_X2 U11417 ( .A1(n10457), .A2(n11564), .ZN(n9604) );
  AND2_X1 U11418 ( .A1(n11581), .A2(n11630), .ZN(n9605) );
  AND2_X1 U11419 ( .A1(n11581), .A2(n11630), .ZN(n9606) );
  AND3_X1 U11420 ( .A1(n11778), .A2(n19545), .A3(n12331), .ZN(n11763) );
  NAND2_X1 U11421 ( .A1(n14147), .A2(n14207), .ZN(n9945) );
  INV_X2 U11422 ( .A(n11904), .ZN(n19828) );
  NOR2_X2 U11423 ( .A1(n15750), .A2(n16297), .ZN(n15738) );
  OR2_X2 U11424 ( .A1(n15763), .A2(n15765), .ZN(n15750) );
  NOR2_X2 U11425 ( .A1(n14734), .A2(n14721), .ZN(n14702) );
  NOR2_X4 U11426 ( .A1(n14066), .A2(n11048), .ZN(n14107) );
  NOR2_X2 U11427 ( .A1(n19413), .A2(n16419), .ZN(n15874) );
  OR2_X2 U11428 ( .A1(n19408), .A2(n19411), .ZN(n19413) );
  AOI21_X2 U11429 ( .B1(n15610), .B2(n19409), .A(n15611), .ZN(n15602) );
  NAND2_X1 U11430 ( .A1(n10141), .A2(n10144), .ZN(n10140) );
  AND2_X1 U11431 ( .A1(n20520), .A2(n9878), .ZN(n11398) );
  NOR2_X1 U11432 ( .A1(n14010), .A2(n10144), .ZN(n9878) );
  NAND2_X1 U11433 ( .A1(n10199), .A2(n16239), .ZN(n10160) );
  INV_X1 U11434 ( .A(n16430), .ZN(n9863) );
  AND2_X1 U11435 ( .A1(n11902), .A2(n11930), .ZN(n9845) );
  NAND2_X1 U11436 ( .A1(n11192), .A2(n10497), .ZN(n10496) );
  INV_X1 U11437 ( .A(n14855), .ZN(n10497) );
  INV_X1 U11438 ( .A(n11398), .ZN(n11416) );
  INV_X1 U11439 ( .A(n10918), .ZN(n10981) );
  AND4_X1 U11441 ( .A1(n11987), .A2(n11986), .A3(n11985), .A4(n11984), .ZN(
        n11994) );
  AND4_X1 U11442 ( .A1(n11983), .A2(n11982), .A3(n11981), .A4(n11980), .ZN(
        n11995) );
  NAND2_X1 U11443 ( .A1(n14561), .A2(n20104), .ZN(n12193) );
  NAND2_X1 U11444 ( .A1(n11639), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11642) );
  NAND2_X1 U11445 ( .A1(n10013), .A2(n9700), .ZN(n16248) );
  NOR2_X1 U11446 ( .A1(n13014), .A2(n11768), .ZN(n11769) );
  NAND2_X1 U11447 ( .A1(n13014), .A2(n13045), .ZN(n19383) );
  AND2_X1 U11448 ( .A1(n10845), .A2(n13254), .ZN(n10821) );
  NAND2_X1 U11449 ( .A1(n11394), .A2(n11419), .ZN(n11395) );
  AND4_X1 U11450 ( .A1(n11991), .A2(n11990), .A3(n11989), .A4(n11988), .ZN(
        n11993) );
  AND2_X1 U11451 ( .A1(n12368), .A2(n12048), .ZN(n10257) );
  OR2_X1 U11452 ( .A1(n11952), .A2(n11951), .ZN(n12379) );
  NOR2_X1 U11453 ( .A1(n14232), .A2(n10185), .ZN(n10183) );
  NAND2_X1 U11454 ( .A1(n10187), .A2(n10186), .ZN(n10185) );
  INV_X1 U11455 ( .A(n10270), .ZN(n10187) );
  NOR2_X1 U11456 ( .A1(n10149), .A2(n10147), .ZN(n10146) );
  INV_X1 U11457 ( .A(n14795), .ZN(n10147) );
  INV_X1 U11458 ( .A(n11364), .ZN(n13158) );
  NOR2_X1 U11459 ( .A1(n11191), .A2(n14871), .ZN(n11192) );
  OR2_X1 U11460 ( .A1(n15037), .A2(n14131), .ZN(n11091) );
  INV_X1 U11461 ( .A(n15048), .ZN(n10355) );
  NAND2_X1 U11462 ( .A1(n10180), .A2(n9694), .ZN(n10248) );
  INV_X1 U11463 ( .A(n15164), .ZN(n10180) );
  NAND2_X1 U11464 ( .A1(n10232), .A2(n15218), .ZN(n10234) );
  NOR2_X1 U11465 ( .A1(n13247), .A2(n10233), .ZN(n10232) );
  INV_X1 U11466 ( .A(n13238), .ZN(n10233) );
  NOR2_X1 U11467 ( .A1(n11019), .A2(n10038), .ZN(n10037) );
  INV_X1 U11468 ( .A(n11039), .ZN(n10038) );
  NAND2_X1 U11469 ( .A1(n10057), .A2(n9706), .ZN(n9928) );
  AND2_X1 U11470 ( .A1(n10227), .A2(n10226), .ZN(n10058) );
  NAND2_X1 U11471 ( .A1(n16916), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10226) );
  NAND2_X1 U11472 ( .A1(n16925), .A2(n16923), .ZN(n10057) );
  AND2_X1 U11473 ( .A1(n21355), .A2(n14671), .ZN(n11555) );
  NAND2_X1 U11474 ( .A1(n13197), .A2(n13196), .ZN(n13199) );
  NAND2_X1 U11475 ( .A1(n10153), .A2(n10879), .ZN(n10152) );
  AND2_X1 U11476 ( .A1(n20541), .A2(n10144), .ZN(n10153) );
  AND3_X1 U11477 ( .A1(n10927), .A2(n10926), .A3(n10925), .ZN(n10928) );
  NAND2_X1 U11478 ( .A1(n9883), .A2(n9884), .ZN(n10930) );
  NAND2_X1 U11479 ( .A1(n9715), .A2(n13189), .ZN(n9884) );
  NOR2_X1 U11480 ( .A1(n10551), .A2(n10572), .ZN(n10836) );
  NOR2_X1 U11481 ( .A1(n14559), .A2(n10096), .ZN(n10095) );
  INV_X1 U11482 ( .A(n10105), .ZN(n10096) );
  NAND2_X1 U11483 ( .A1(n10121), .A2(n10119), .ZN(n14502) );
  AND2_X1 U11484 ( .A1(n14499), .A2(n10120), .ZN(n10119) );
  INV_X1 U11485 ( .A(n10122), .ZN(n10120) );
  AND2_X1 U11486 ( .A1(n13524), .A2(n13523), .ZN(n14556) );
  NOR2_X1 U11487 ( .A1(n10064), .A2(n14059), .ZN(n13523) );
  NAND2_X1 U11488 ( .A1(n12529), .A2(n12522), .ZN(n12584) );
  NOR2_X1 U11489 ( .A1(n12547), .A2(n12546), .ZN(n12583) );
  NAND2_X1 U11490 ( .A1(n10220), .A2(n10445), .ZN(n16194) );
  AND2_X1 U11491 ( .A1(n10544), .A2(n10218), .ZN(n10217) );
  NAND2_X1 U11492 ( .A1(n10219), .A2(n10546), .ZN(n10218) );
  AND2_X1 U11493 ( .A1(n12295), .A2(n15703), .ZN(n10421) );
  NAND2_X1 U11494 ( .A1(n10160), .A2(n16238), .ZN(n10159) );
  NAND2_X1 U11495 ( .A1(n9705), .A2(n12499), .ZN(n9910) );
  NOR2_X1 U11496 ( .A1(n9665), .A2(n9965), .ZN(n9964) );
  INV_X1 U11497 ( .A(n15762), .ZN(n9965) );
  OR2_X1 U11498 ( .A1(n15768), .A2(n12048), .ZN(n12488) );
  AND2_X1 U11499 ( .A1(n12066), .A2(n13529), .ZN(n10487) );
  INV_X1 U11500 ( .A(n13637), .ZN(n12066) );
  NAND2_X1 U11501 ( .A1(n11822), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10001) );
  OAI21_X1 U11502 ( .B1(n11809), .B2(n11808), .A(n11807), .ZN(n10003) );
  NAND2_X1 U11503 ( .A1(n10541), .A2(n12035), .ZN(n9799) );
  AND2_X1 U11504 ( .A1(n11804), .A2(n12320), .ZN(n11776) );
  MUX2_X1 U11505 ( .A(n11774), .B(n11805), .S(n11803), .Z(n11775) );
  NAND2_X1 U11506 ( .A1(n13697), .A2(n10580), .ZN(n13766) );
  AND3_X1 U11507 ( .A1(n12337), .A2(n11765), .A3(n11764), .ZN(n13865) );
  NAND2_X1 U11508 ( .A1(n10050), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10049) );
  INV_X1 U11509 ( .A(n11741), .ZN(n10074) );
  INV_X1 U11510 ( .A(n12842), .ZN(n17578) );
  NOR2_X1 U11511 ( .A1(n12617), .A2(n12618), .ZN(n12639) );
  OR2_X1 U11512 ( .A1(n12617), .A2(n12620), .ZN(n17563) );
  NOR2_X1 U11513 ( .A1(n17466), .A2(n12620), .ZN(n12803) );
  NOR2_X1 U11514 ( .A1(n10173), .A2(n10172), .ZN(n10171) );
  OAI21_X1 U11515 ( .B1(n10284), .B2(n18413), .A(n18407), .ZN(n10172) );
  INV_X1 U11516 ( .A(n10386), .ZN(n10173) );
  NAND2_X1 U11517 ( .A1(n10283), .A2(n18120), .ZN(n10282) );
  AND2_X1 U11518 ( .A1(n12860), .A2(n12892), .ZN(n12862) );
  NOR2_X1 U11519 ( .A1(n18303), .A2(n18306), .ZN(n12910) );
  AOI21_X1 U11520 ( .B1(n18736), .B2(n12706), .A(n12954), .ZN(n12877) );
  AND3_X1 U11521 ( .A1(n12886), .A2(n12951), .A3(n19163), .ZN(n14234) );
  NOR2_X1 U11522 ( .A1(n18736), .A2(n18732), .ZN(n19162) );
  NAND2_X1 U11523 ( .A1(n13730), .A2(n11453), .ZN(n13470) );
  NOR2_X1 U11524 ( .A1(n10486), .A2(n14777), .ZN(n10485) );
  INV_X1 U11525 ( .A(n14783), .ZN(n10486) );
  CLKBUF_X1 U11526 ( .A(n10986), .Z(n11374) );
  NOR3_X1 U11527 ( .A1(n10501), .A2(n11382), .A3(n10499), .ZN(n10498) );
  INV_X1 U11528 ( .A(n14720), .ZN(n10499) );
  OR2_X1 U11529 ( .A1(n16883), .A2(n20288), .ZN(n13556) );
  NAND2_X1 U11530 ( .A1(n9877), .A2(n15263), .ZN(n15372) );
  OR2_X1 U11531 ( .A1(n15397), .A2(n15373), .ZN(n9877) );
  NAND2_X1 U11532 ( .A1(n15151), .A2(n9934), .ZN(n9933) );
  NOR2_X1 U11533 ( .A1(n15198), .A2(n15195), .ZN(n9934) );
  AND2_X1 U11534 ( .A1(n13738), .A2(n13731), .ZN(n15382) );
  INV_X1 U11535 ( .A(n16942), .ZN(n15469) );
  NAND2_X1 U11536 ( .A1(n9670), .A2(n9817), .ZN(n16933) );
  NAND2_X1 U11537 ( .A1(n13738), .A2(n13733), .ZN(n16939) );
  NAND2_X1 U11538 ( .A1(n15469), .A2(n16939), .ZN(n16944) );
  OR2_X1 U11539 ( .A1(n13472), .A2(n11390), .ZN(n16864) );
  AND2_X1 U11540 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11582) );
  NAND2_X1 U11541 ( .A1(n10435), .A2(n10436), .ZN(n10113) );
  NAND2_X1 U11542 ( .A1(n15981), .A2(n14592), .ZN(n10436) );
  NAND2_X1 U11543 ( .A1(n13764), .A2(n13763), .ZN(n10118) );
  INV_X1 U11544 ( .A(n20264), .ZN(n16766) );
  NAND2_X1 U11545 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12307) );
  INV_X1 U11547 ( .A(n12991), .ZN(n12580) );
  INV_X1 U11548 ( .A(n12579), .ZN(n10443) );
  NAND2_X1 U11549 ( .A1(n12994), .A2(n10414), .ZN(n12568) );
  AND2_X1 U11550 ( .A1(n12995), .A2(n12312), .ZN(n10414) );
  NAND2_X1 U11551 ( .A1(n16276), .A2(n16274), .ZN(n10216) );
  NAND2_X1 U11552 ( .A1(n10538), .A2(n9696), .ZN(n16262) );
  NAND2_X1 U11553 ( .A1(n16248), .A2(n16247), .ZN(n10538) );
  INV_X1 U11554 ( .A(n10516), .ZN(n10515) );
  OAI21_X1 U11555 ( .B1(n10520), .B2(n10517), .A(n16323), .ZN(n10516) );
  INV_X1 U11556 ( .A(n16322), .ZN(n10517) );
  INV_X1 U11557 ( .A(n16364), .ZN(n10336) );
  AOI21_X1 U11558 ( .B1(n9676), .B2(n11998), .A(n9622), .ZN(n9947) );
  NAND2_X1 U11559 ( .A1(n16400), .A2(n9676), .ZN(n9948) );
  AND3_X1 U11560 ( .A1(n12033), .A2(n12032), .A3(n12031), .ZN(n13972) );
  AOI21_X1 U11561 ( .B1(n12030), .B2(n10211), .A(n10210), .ZN(n12033) );
  NAND2_X1 U11562 ( .A1(n11658), .A2(n11657), .ZN(n13905) );
  CLKBUF_X1 U11563 ( .A(n12314), .Z(n13892) );
  INV_X1 U11564 ( .A(n19820), .ZN(n19857) );
  NAND2_X1 U11565 ( .A1(n11611), .A2(n11839), .ZN(n10360) );
  NOR2_X1 U11566 ( .A1(n17145), .A2(n17434), .ZN(n17137) );
  AOI22_X1 U11567 ( .A1(n14234), .A2(n9744), .B1(n10328), .B2(n10327), .ZN(
        n16896) );
  NOR2_X1 U11568 ( .A1(n17826), .A2(n14224), .ZN(n10327) );
  INV_X1 U11569 ( .A(n14223), .ZN(n10328) );
  NOR2_X1 U11570 ( .A1(n10083), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10082) );
  INV_X1 U11571 ( .A(n13038), .ZN(n10083) );
  INV_X1 U11572 ( .A(n18353), .ZN(n10166) );
  NOR3_X1 U11573 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n19215), .A3(n18707), 
        .ZN(n19353) );
  NOR2_X1 U11574 ( .A1(n16177), .A2(n15955), .ZN(n13058) );
  AND2_X1 U11575 ( .A1(n14345), .A2(n14344), .ZN(n14346) );
  NAND2_X1 U11576 ( .A1(n19383), .A2(n13016), .ZN(n16436) );
  INV_X1 U11577 ( .A(n16433), .ZN(n16413) );
  OR2_X1 U11578 ( .A1(n14369), .A2(n16708), .ZN(n12578) );
  INV_X1 U11579 ( .A(n16573), .ZN(n9969) );
  AND2_X1 U11580 ( .A1(n9620), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10018) );
  NAND2_X1 U11581 ( .A1(n11436), .A2(n20516), .ZN(n11439) );
  AND2_X1 U11582 ( .A1(n14647), .A2(n11383), .ZN(n11407) );
  NAND2_X1 U11583 ( .A1(n12209), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n11819) );
  NAND2_X1 U11584 ( .A1(n11741), .A2(n11674), .ZN(n10069) );
  NAND2_X1 U11585 ( .A1(n10064), .A2(n10067), .ZN(n10066) );
  BUF_X1 U11586 ( .A(n10699), .Z(n10667) );
  NOR2_X1 U11587 ( .A1(n10582), .A2(n14013), .ZN(n10151) );
  INV_X1 U11588 ( .A(n10032), .ZN(n10031) );
  AOI22_X1 U11589 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9619), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10701) );
  INV_X1 U11590 ( .A(n11407), .ZN(n9868) );
  AND3_X1 U11591 ( .A1(n11960), .A2(n11958), .A3(n11959), .ZN(n10383) );
  NOR2_X1 U11592 ( .A1(n9895), .A2(n9891), .ZN(n10381) );
  NAND2_X1 U11593 ( .A1(n16774), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n9894) );
  INV_X1 U11594 ( .A(n11793), .ZN(n11779) );
  XNOR2_X1 U11595 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11628) );
  NAND2_X1 U11596 ( .A1(n18379), .A2(n17926), .ZN(n9999) );
  AOI21_X1 U11597 ( .B1(n19189), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12711), .ZN(n12717) );
  AND2_X1 U11598 ( .A1(n12873), .A2(n12871), .ZN(n12711) );
  INV_X1 U11599 ( .A(n18736), .ZN(n12699) );
  NOR2_X1 U11600 ( .A1(n14753), .A2(n10504), .ZN(n10503) );
  INV_X1 U11601 ( .A(n10505), .ZN(n10504) );
  NAND2_X1 U11602 ( .A1(n16846), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11364) );
  AND2_X1 U11603 ( .A1(n13169), .A2(n14127), .ZN(n10960) );
  INV_X1 U11604 ( .A(n10986), .ZN(n11368) );
  INV_X1 U11605 ( .A(n10818), .ZN(n10983) );
  NOR2_X1 U11606 ( .A1(n10474), .A2(n10472), .ZN(n10471) );
  INV_X1 U11607 ( .A(n11558), .ZN(n10474) );
  INV_X1 U11608 ( .A(n14754), .ZN(n10484) );
  NOR2_X1 U11609 ( .A1(n10391), .A2(n15362), .ZN(n10388) );
  AND2_X1 U11610 ( .A1(n10388), .A2(n13238), .ZN(n10245) );
  INV_X1 U11611 ( .A(n14891), .ZN(n10480) );
  OAI21_X1 U11612 ( .B1(n15560), .B2(n9916), .A(n9914), .ZN(n9919) );
  NAND2_X1 U11613 ( .A1(n13222), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9916) );
  INV_X1 U11614 ( .A(n9915), .ZN(n9914) );
  OAI21_X1 U11615 ( .B1(n13205), .B2(n13206), .A(n20461), .ZN(n9915) );
  INV_X1 U11616 ( .A(n16974), .ZN(n11482) );
  NAND2_X1 U11617 ( .A1(n9880), .A2(n9704), .ZN(n13713) );
  NAND2_X1 U11619 ( .A1(n9924), .A2(n9754), .ZN(n10863) );
  INV_X1 U11620 ( .A(n10858), .ZN(n9924) );
  OAI21_X1 U11621 ( .B1(n10032), .B2(n9922), .A(n9920), .ZN(n10864) );
  INV_X1 U11622 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9922) );
  NOR2_X1 U11623 ( .A1(n9752), .A2(n9921), .ZN(n9920) );
  NOR2_X1 U11624 ( .A1(n16880), .A2(n20836), .ZN(n9921) );
  OR2_X1 U11625 ( .A1(n10930), .A2(n10929), .ZN(n10168) );
  NAND2_X1 U11626 ( .A1(n10877), .A2(n10907), .ZN(n10142) );
  XNOR2_X1 U11627 ( .A(n10967), .B(n9886), .ZN(n15556) );
  INV_X1 U11628 ( .A(n10968), .ZN(n9886) );
  NAND2_X1 U11629 ( .A1(n10285), .A2(n11434), .ZN(n13254) );
  AND2_X1 U11630 ( .A1(n13476), .A2(n13475), .ZN(n13716) );
  INV_X1 U11631 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20901) );
  NAND2_X1 U11632 ( .A1(n11415), .A2(n11414), .ZN(n13298) );
  OR2_X1 U11633 ( .A1(n11423), .A2(n11422), .ZN(n11415) );
  NAND2_X1 U11634 ( .A1(n10209), .A2(n10208), .ZN(n12374) );
  NAND2_X1 U11635 ( .A1(n11800), .A2(n11746), .ZN(n10208) );
  NAND2_X1 U11636 ( .A1(n10211), .A2(n11780), .ZN(n10209) );
  OR2_X1 U11637 ( .A1(n11686), .A2(n11685), .ZN(n11901) );
  AND2_X1 U11638 ( .A1(n10558), .A2(n12464), .ZN(n10456) );
  OR2_X1 U11639 ( .A1(n12407), .A2(n10451), .ZN(n12434) );
  NAND2_X1 U11640 ( .A1(n9714), .A2(n10207), .ZN(n12423) );
  INV_X1 U11641 ( .A(n12407), .ZN(n10207) );
  CLKBUF_X1 U11642 ( .A(n11942), .Z(n12094) );
  NOR2_X2 U11643 ( .A1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14443) );
  AND2_X1 U11644 ( .A1(n14592), .A2(n10063), .ZN(n14593) );
  AND2_X1 U11645 ( .A1(n15988), .A2(n14592), .ZN(n10437) );
  AOI21_X1 U11646 ( .B1(n14601), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A(n9778), .ZN(n14485) );
  NAND2_X1 U11647 ( .A1(n10578), .A2(n10441), .ZN(n10440) );
  INV_X1 U11648 ( .A(n16049), .ZN(n10441) );
  AND2_X1 U11649 ( .A1(n9733), .A2(n13765), .ZN(n10117) );
  NAND2_X1 U11650 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12301) );
  OR2_X1 U11651 ( .A1(n15674), .A2(n16023), .ZN(n15656) );
  NAND2_X1 U11652 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12289) );
  NAND2_X1 U11653 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12260) );
  INV_X1 U11654 ( .A(n15767), .ZN(n10408) );
  NOR2_X1 U11655 ( .A1(n10379), .A2(n10378), .ZN(n10377) );
  NAND2_X1 U11656 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12225) );
  INV_X1 U11657 ( .A(n10160), .ZN(n10158) );
  NAND2_X1 U11658 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12254) );
  INV_X1 U11659 ( .A(n14194), .ZN(n12257) );
  INV_X1 U11660 ( .A(n16329), .ZN(n10522) );
  INV_X1 U11661 ( .A(n13957), .ZN(n10413) );
  INV_X1 U11662 ( .A(n14098), .ZN(n12228) );
  INV_X1 U11663 ( .A(n13835), .ZN(n12229) );
  NAND2_X1 U11664 ( .A1(n11997), .A2(n16681), .ZN(n9949) );
  INV_X1 U11665 ( .A(n16417), .ZN(n11997) );
  NOR2_X1 U11666 ( .A1(n11998), .A2(n9622), .ZN(n10361) );
  OAI21_X1 U11667 ( .B1(n9676), .B2(n9622), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10363) );
  NOR2_X1 U11668 ( .A1(n11971), .A2(n11970), .ZN(n12381) );
  INV_X1 U11669 ( .A(n13773), .ZN(n12213) );
  INV_X1 U11670 ( .A(n13803), .ZN(n10417) );
  XNOR2_X1 U11671 ( .A(n10028), .B(n12383), .ZN(n11954) );
  NAND2_X1 U11672 ( .A1(n11779), .A2(n11803), .ZN(n12330) );
  NAND2_X1 U11673 ( .A1(n12328), .A2(n10063), .ZN(n13885) );
  NAND2_X1 U11674 ( .A1(n11880), .A2(n11875), .ZN(n11907) );
  AND2_X1 U11675 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19754) );
  INV_X1 U11676 ( .A(n11905), .ZN(n19990) );
  INV_X1 U11677 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20032) );
  NAND2_X1 U11678 ( .A1(n10321), .A2(n18081), .ZN(n10318) );
  INV_X1 U11679 ( .A(n18095), .ZN(n10316) );
  NAND2_X1 U11681 ( .A1(n19162), .A2(n12884), .ZN(n14223) );
  NAND2_X1 U11682 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10087) );
  INV_X1 U11683 ( .A(n12816), .ZN(n10086) );
  NAND2_X1 U11684 ( .A1(n9805), .A2(n9804), .ZN(n12678) );
  INV_X1 U11685 ( .A(n12618), .ZN(n9804) );
  INV_X1 U11686 ( .A(n10167), .ZN(n9805) );
  NAND2_X1 U11687 ( .A1(n10182), .A2(n10184), .ZN(n16898) );
  NAND2_X1 U11688 ( .A1(n9713), .A2(n10186), .ZN(n10184) );
  NOR3_X1 U11689 ( .A1(n18732), .A2(n18749), .A3(n14224), .ZN(n12702) );
  INV_X1 U11690 ( .A(n18721), .ZN(n17424) );
  AND2_X1 U11691 ( .A1(n10324), .A2(n10568), .ZN(n10323) );
  NOR2_X1 U11692 ( .A1(n12596), .A2(n17477), .ZN(n10324) );
  NAND2_X1 U11693 ( .A1(n10574), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9979) );
  NAND2_X1 U11694 ( .A1(n10170), .A2(n9976), .ZN(n9975) );
  NOR2_X1 U11695 ( .A1(n10304), .A2(n9980), .ZN(n9976) );
  NAND2_X1 U11696 ( .A1(n9978), .A2(n10574), .ZN(n9977) );
  INV_X1 U11697 ( .A(n10171), .ZN(n9978) );
  NAND2_X1 U11698 ( .A1(n10089), .A2(n18433), .ZN(n10283) );
  NOR2_X1 U11699 ( .A1(n18178), .A2(n18489), .ZN(n18120) );
  NAND2_X1 U11700 ( .A1(n9994), .A2(n18228), .ZN(n12866) );
  OR2_X1 U11701 ( .A1(n18261), .A2(n9995), .ZN(n9994) );
  NAND2_X1 U11702 ( .A1(n17926), .A2(n17922), .ZN(n12852) );
  NAND2_X1 U11703 ( .A1(n10338), .A2(n10337), .ZN(n12902) );
  OAI21_X1 U11704 ( .B1(n16901), .B2(n9983), .A(n17922), .ZN(n10337) );
  INV_X1 U11705 ( .A(n18745), .ZN(n12697) );
  NOR2_X1 U11706 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12709), .ZN(
        n12871) );
  AOI22_X1 U11707 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19189), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n12710), .ZN(n12873) );
  AOI21_X1 U11708 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n19197), .A(
        n12720), .ZN(n12875) );
  NOR2_X1 U11709 ( .A1(n12619), .A2(n19179), .ZN(n12802) );
  NAND2_X1 U11710 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12837) );
  NAND2_X1 U11711 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14229) );
  INV_X1 U11712 ( .A(n12678), .ZN(n12843) );
  NAND2_X1 U11713 ( .A1(n10267), .A2(n10266), .ZN(n10265) );
  NAND2_X1 U11714 ( .A1(n19336), .A2(n19189), .ZN(n10266) );
  OAI21_X1 U11715 ( .B1(n19336), .B2(n10268), .A(n19331), .ZN(n10267) );
  NAND2_X1 U11716 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10268) );
  AND2_X1 U11717 ( .A1(n11532), .A2(n11531), .ZN(n14777) );
  AND2_X1 U11718 ( .A1(n14859), .A2(n9760), .ZN(n14796) );
  INV_X1 U11719 ( .A(n14812), .ZN(n10475) );
  NOR2_X1 U11720 ( .A1(n14706), .A2(n10501), .ZN(n10500) );
  NAND2_X1 U11721 ( .A1(n11358), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11372) );
  NAND2_X1 U11722 ( .A1(n11340), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11350) );
  NAND2_X1 U11723 ( .A1(n11322), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11333) );
  OR2_X1 U11724 ( .A1(n15119), .A2(n11371), .ZN(n11298) );
  NOR2_X2 U11725 ( .A1(n11226), .A2(n15143), .ZN(n11243) );
  NOR2_X1 U11726 ( .A1(n10496), .A2(n10495), .ZN(n10494) );
  INV_X1 U11727 ( .A(n14841), .ZN(n10495) );
  NAND2_X1 U11728 ( .A1(n10587), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11157) );
  AND3_X1 U11729 ( .A1(n11079), .A2(n11078), .A3(n11077), .ZN(n15037) );
  OR2_X1 U11730 ( .A1(n14702), .A2(n14671), .ZN(n10467) );
  OR2_X1 U11731 ( .A1(n10471), .A2(n14671), .ZN(n10468) );
  AND2_X1 U11732 ( .A1(n15080), .A2(n9725), .ZN(n10040) );
  AND2_X1 U11733 ( .A1(n10402), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10401) );
  NOR2_X1 U11734 ( .A1(n15265), .A2(n10403), .ZN(n10402) );
  NAND2_X1 U11735 ( .A1(n13253), .A2(n10043), .ZN(n10041) );
  AND2_X1 U11736 ( .A1(n13252), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10043) );
  INV_X1 U11737 ( .A(n14352), .ZN(n13253) );
  INV_X1 U11738 ( .A(n10472), .ZN(n10470) );
  NAND2_X1 U11739 ( .A1(n15086), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10244) );
  INV_X1 U11740 ( .A(n15099), .ZN(n10243) );
  INV_X1 U11741 ( .A(n10244), .ZN(n15095) );
  NAND2_X1 U11742 ( .A1(n10352), .A2(n10583), .ZN(n15107) );
  AND2_X1 U11743 ( .A1(n13246), .A2(n10353), .ZN(n10231) );
  AND2_X1 U11744 ( .A1(n10555), .A2(n9790), .ZN(n10353) );
  INV_X1 U11745 ( .A(n10248), .ZN(n13246) );
  INV_X1 U11746 ( .A(n15154), .ZN(n9932) );
  NOR2_X1 U11747 ( .A1(n15236), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9930) );
  NAND2_X1 U11748 ( .A1(n15179), .A2(n15176), .ZN(n15164) );
  AND2_X1 U11749 ( .A1(n13751), .A2(n13750), .ZN(n15467) );
  NAND2_X1 U11750 ( .A1(n9926), .A2(n9693), .ZN(n15151) );
  OR2_X1 U11751 ( .A1(n9928), .A2(n9927), .ZN(n9926) );
  OR2_X1 U11752 ( .A1(n13236), .A2(n9927), .ZN(n9925) );
  OR2_X1 U11753 ( .A1(n20477), .A2(n15382), .ZN(n16942) );
  NAND2_X1 U11754 ( .A1(n9820), .A2(n13200), .ZN(n13944) );
  INV_X1 U11755 ( .A(n16939), .ZN(n20460) );
  OAI211_X1 U11756 ( .C1(n13193), .C2(n13192), .A(n13191), .B(n9937), .ZN(
        n13649) );
  NAND2_X1 U11757 ( .A1(n13193), .A2(n9938), .ZN(n9937) );
  NAND2_X1 U11758 ( .A1(n14651), .A2(n11466), .ZN(n14652) );
  XNOR2_X1 U11759 ( .A(n10930), .B(n10928), .ZN(n10974) );
  NAND2_X1 U11760 ( .A1(n15560), .A2(n20494), .ZN(n20610) );
  INV_X1 U11761 ( .A(n20648), .ZN(n20742) );
  AND2_X1 U11762 ( .A1(n20976), .A2(n20497), .ZN(n20842) );
  INV_X1 U11763 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20873) );
  AND2_X1 U11764 ( .A1(n15553), .A2(n20495), .ZN(n20871) );
  INV_X1 U11765 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20933) );
  NAND2_X1 U11766 ( .A1(n10882), .A2(n10881), .ZN(n20541) );
  INV_X1 U11767 ( .A(n10880), .ZN(n10881) );
  INV_X1 U11768 ( .A(n13484), .ZN(n20981) );
  NOR2_X1 U11769 ( .A1(n20834), .A2(n20649), .ZN(n20985) );
  INV_X1 U11770 ( .A(n20809), .ZN(n20932) );
  AND2_X1 U11771 ( .A1(n15562), .A2(n10949), .ZN(n20978) );
  AOI21_X1 U11772 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20933), .A(n20649), 
        .ZN(n21018) );
  NOR2_X1 U11773 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13926) );
  NOR2_X1 U11774 ( .A1(n11786), .A2(n13517), .ZN(n10422) );
  XNOR2_X1 U11775 ( .A(n12549), .B(n12548), .ZN(n12550) );
  AND2_X1 U11776 ( .A1(n10454), .A2(n15999), .ZN(n10453) );
  NAND2_X1 U11777 ( .A1(n12465), .A2(n10456), .ZN(n12456) );
  NAND2_X1 U11778 ( .A1(n12463), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10223) );
  NAND2_X1 U11779 ( .A1(n12482), .A2(n9701), .ZN(n12478) );
  AND2_X1 U11780 ( .A1(n9633), .A2(n12466), .ZN(n10224) );
  OR2_X1 U11781 ( .A1(n16750), .A2(n15940), .ZN(n15950) );
  NAND2_X1 U11782 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12305) );
  NAND2_X1 U11783 ( .A1(n10118), .A2(n10117), .ZN(n13821) );
  INV_X1 U11784 ( .A(n13525), .ZN(n13624) );
  NAND2_X1 U11785 ( .A1(n10425), .A2(n9695), .ZN(n10102) );
  NOR2_X1 U11786 ( .A1(n14559), .A2(n10098), .ZN(n10097) );
  NOR2_X1 U11787 ( .A1(n15981), .A2(n10099), .ZN(n15989) );
  AND2_X1 U11788 ( .A1(n10104), .A2(n10100), .ZN(n10099) );
  NAND2_X1 U11789 ( .A1(n10425), .A2(n9666), .ZN(n10104) );
  AOI21_X1 U11790 ( .B1(n15993), .B2(n15996), .A(n10103), .ZN(n10100) );
  AOI21_X1 U11791 ( .B1(n14502), .B2(n14501), .A(n14537), .ZN(n15993) );
  AND3_X1 U11792 ( .A1(n12093), .A2(n12092), .A3(n12091), .ZN(n13681) );
  NAND2_X1 U11793 ( .A1(n13793), .A2(n13792), .ZN(n13794) );
  OR2_X1 U11794 ( .A1(n19431), .A2(n13536), .ZN(n14366) );
  NAND2_X1 U11795 ( .A1(n13905), .A2(n10063), .ZN(n13868) );
  AND2_X1 U11796 ( .A1(n13348), .A2(n13057), .ZN(n19489) );
  NOR2_X1 U11797 ( .A1(n10064), .A2(n20166), .ZN(n13057) );
  AND2_X1 U11798 ( .A1(n10579), .A2(n10418), .ZN(n15597) );
  AND2_X1 U11799 ( .A1(n9675), .A2(n10419), .ZN(n10418) );
  INV_X1 U11800 ( .A(n12743), .ZN(n10419) );
  INV_X1 U11801 ( .A(n10380), .ZN(n13109) );
  AND2_X1 U11802 ( .A1(n12273), .A2(n12272), .ZN(n15718) );
  NAND2_X1 U11803 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12219) );
  XNOR2_X1 U11804 ( .A(n12204), .B(n11847), .ZN(n11835) );
  OR2_X1 U11805 ( .A1(n12198), .A2(n12562), .ZN(n14623) );
  AND2_X1 U11806 ( .A1(n13009), .A2(n13008), .ZN(n15580) );
  AND2_X1 U11807 ( .A1(n10543), .A2(n12542), .ZN(n10202) );
  NAND2_X1 U11808 ( .A1(n10446), .A2(n10445), .ZN(n10201) );
  NAND2_X1 U11809 ( .A1(n12515), .A2(n10546), .ZN(n10203) );
  AND2_X1 U11810 ( .A1(n10053), .A2(n12351), .ZN(n9950) );
  NOR2_X1 U11811 ( .A1(n9794), .A2(n12738), .ZN(n10511) );
  AND2_X1 U11812 ( .A1(n12518), .A2(n12412), .ZN(n10448) );
  NAND2_X1 U11813 ( .A1(n9961), .A2(n9775), .ZN(n15632) );
  INV_X1 U11814 ( .A(n15636), .ZN(n9960) );
  NAND2_X1 U11815 ( .A1(n10579), .A2(n9675), .ZN(n15624) );
  AND2_X1 U11816 ( .A1(n10510), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10255) );
  NAND2_X1 U11817 ( .A1(n9669), .A2(n10564), .ZN(n9907) );
  INV_X1 U11818 ( .A(n9910), .ZN(n12500) );
  NAND2_X1 U11819 ( .A1(n16362), .A2(n16361), .ZN(n10335) );
  NAND2_X1 U11820 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12292) );
  AND2_X1 U11821 ( .A1(n15717), .A2(n12274), .ZN(n10579) );
  INV_X1 U11822 ( .A(n15718), .ZN(n12274) );
  NAND2_X1 U11823 ( .A1(n9623), .A2(n15701), .ZN(n9962) );
  NAND2_X1 U11824 ( .A1(n16267), .A2(n16536), .ZN(n16290) );
  OR2_X1 U11825 ( .A1(n10528), .A2(n10522), .ZN(n10521) );
  OR3_X1 U11826 ( .A1(n12490), .A2(n12048), .A3(n21336), .ZN(n16322) );
  OR2_X1 U11827 ( .A1(n10524), .A2(n10522), .ZN(n10520) );
  AOI21_X1 U11828 ( .B1(n10527), .B2(n10526), .A(n10525), .ZN(n10524) );
  INV_X1 U11829 ( .A(n16330), .ZN(n10525) );
  INV_X1 U11830 ( .A(n10529), .ZN(n10526) );
  NOR2_X1 U11831 ( .A1(n14085), .A2(n10411), .ZN(n10409) );
  INV_X1 U11832 ( .A(n13933), .ZN(n10410) );
  NAND2_X1 U11833 ( .A1(n10412), .A2(n14161), .ZN(n10411) );
  AND2_X1 U11834 ( .A1(n16340), .A2(n16352), .ZN(n10529) );
  AND3_X1 U11835 ( .A1(n12149), .A2(n12148), .A3(n12147), .ZN(n13997) );
  NOR2_X1 U11836 ( .A1(n13675), .A2(n13745), .ZN(n13779) );
  AND3_X1 U11837 ( .A1(n12065), .A2(n12064), .A3(n12063), .ZN(n13637) );
  AND2_X1 U11838 ( .A1(n16695), .A2(n16693), .ZN(n12357) );
  NAND2_X1 U11839 ( .A1(n10405), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12222) );
  NAND2_X1 U11840 ( .A1(n9849), .A2(n9850), .ZN(n11932) );
  INV_X1 U11841 ( .A(n13972), .ZN(n12034) );
  INV_X1 U11842 ( .A(n11856), .ZN(n9844) );
  NAND4_X1 U11843 ( .A1(n10571), .A2(n11673), .A3(n11672), .A4(n11671), .ZN(
        n13428) );
  NAND2_X1 U11844 ( .A1(n13659), .A2(n13658), .ZN(n13661) );
  NAND2_X1 U11845 ( .A1(n13497), .A2(n20104), .ZN(n13693) );
  XNOR2_X1 U11846 ( .A(n13525), .B(n13623), .ZN(n13526) );
  AND2_X1 U11847 ( .A1(n13701), .A2(n13767), .ZN(n13763) );
  INV_X1 U11848 ( .A(n19696), .ZN(n19693) );
  INV_X1 U11849 ( .A(n11907), .ZN(n19727) );
  AND2_X1 U11850 ( .A1(n19598), .A2(n19522), .ZN(n19753) );
  NOR2_X1 U11851 ( .A1(n19897), .A2(n19896), .ZN(n10026) );
  NAND2_X1 U11852 ( .A1(n16766), .A2(n19523), .ZN(n19993) );
  OR2_X1 U11853 ( .A1(n19598), .A2(n19522), .ZN(n19988) );
  NAND2_X1 U11854 ( .A1(n16752), .A2(n14059), .ZN(n13505) );
  NAND2_X1 U11855 ( .A1(n10027), .A2(n19522), .ZN(n20031) );
  AND2_X1 U11856 ( .A1(n11744), .A2(n11743), .ZN(n13910) );
  NOR2_X1 U11857 ( .A1(n14230), .A2(n14232), .ZN(n19152) );
  INV_X1 U11858 ( .A(n12950), .ZN(n19153) );
  NAND2_X1 U11859 ( .A1(n10301), .A2(n10299), .ZN(n19202) );
  NAND2_X1 U11860 ( .A1(n10300), .A2(n19154), .ZN(n10299) );
  INV_X1 U11861 ( .A(n19155), .ZN(n10300) );
  OAI22_X1 U11862 ( .A1(n17137), .A2(n10325), .B1(n10321), .B2(n17118), .ZN(
        n17120) );
  OR2_X1 U11863 ( .A1(n17118), .A2(n17138), .ZN(n10325) );
  INV_X1 U11864 ( .A(n17188), .ZN(n10320) );
  NAND2_X1 U11865 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10192) );
  CLKBUF_X2 U11866 ( .A(n12787), .Z(n17499) );
  NAND2_X1 U11867 ( .A1(n18219), .A2(n18381), .ZN(n18169) );
  NOR2_X1 U11868 ( .A1(n9980), .A2(n18047), .ZN(n10305) );
  NAND2_X1 U11869 ( .A1(n10170), .A2(n18228), .ZN(n10169) );
  NOR2_X1 U11870 ( .A1(n10387), .A2(n9755), .ZN(n10386) );
  NOR2_X1 U11871 ( .A1(n10304), .A2(n18433), .ZN(n10387) );
  INV_X1 U11872 ( .A(n18571), .ZN(n18549) );
  INV_X1 U11873 ( .A(n19161), .ZN(n10271) );
  NAND2_X1 U11874 ( .A1(n19167), .A2(n19162), .ZN(n10269) );
  NAND2_X1 U11875 ( .A1(n18311), .A2(n12909), .ZN(n18304) );
  NAND2_X1 U11876 ( .A1(n12905), .A2(n18658), .ZN(n9997) );
  INV_X1 U11877 ( .A(n10279), .ZN(n9807) );
  NAND2_X1 U11878 ( .A1(n18353), .A2(n12853), .ZN(n10279) );
  AND2_X1 U11879 ( .A1(n9813), .A2(n9724), .ZN(n18363) );
  NOR2_X1 U11880 ( .A1(n12697), .A2(n18732), .ZN(n12951) );
  NAND2_X1 U11881 ( .A1(n9815), .A2(n9814), .ZN(n9813) );
  INV_X1 U11882 ( .A(n18373), .ZN(n9815) );
  INV_X1 U11883 ( .A(n18372), .ZN(n9814) );
  XNOR2_X1 U11884 ( .A(n17926), .B(n19320), .ZN(n18373) );
  NAND2_X1 U11885 ( .A1(n12959), .A2(n12952), .ZN(n19155) );
  INV_X1 U11886 ( .A(n19173), .ZN(n14230) );
  OR2_X1 U11887 ( .A1(n13381), .A2(n20288), .ZN(n14006) );
  OR3_X1 U11888 ( .A1(n16883), .A2(n13304), .A3(n20288), .ZN(n14007) );
  AND2_X1 U11889 ( .A1(n20345), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20369) );
  NAND2_X1 U11890 ( .A1(n11461), .A2(n11460), .ZN(n20396) );
  INV_X1 U11891 ( .A(n14976), .ZN(n10131) );
  INV_X1 U11892 ( .A(n13292), .ZN(n10136) );
  AOI21_X2 U11893 ( .B1(n11382), .B2(n11381), .A(n13293), .ZN(n15054) );
  INV_X1 U11894 ( .A(n16937), .ZN(n16921) );
  NAND2_X1 U11895 ( .A1(n15290), .A2(n20473), .ZN(n9875) );
  XNOR2_X1 U11896 ( .A(n10061), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15292) );
  OAI21_X1 U11897 ( .B1(n14351), .B2(n15048), .A(n14350), .ZN(n10061) );
  NAND2_X1 U11898 ( .A1(n10044), .A2(n13251), .ZN(n14351) );
  NAND2_X1 U11899 ( .A1(n13253), .A2(n13252), .ZN(n14350) );
  XNOR2_X1 U11900 ( .A(n15070), .B(n15317), .ZN(n15315) );
  NAND2_X1 U11901 ( .A1(n15069), .A2(n15068), .ZN(n15070) );
  OAI21_X1 U11902 ( .B1(n13251), .B2(n15265), .A(n15216), .ZN(n15068) );
  NOR2_X1 U11903 ( .A1(n15350), .A2(n15266), .ZN(n15326) );
  AND2_X1 U11904 ( .A1(n13738), .A2(n13729), .ZN(n20473) );
  INV_X1 U11905 ( .A(n20473), .ZN(n20486) );
  NOR2_X2 U11906 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20934) );
  NOR2_X1 U11907 ( .A1(n15560), .A2(n15562), .ZN(n20872) );
  OR2_X1 U11908 ( .A1(n20750), .A2(n20749), .ZN(n20772) );
  INV_X1 U11909 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21095) );
  NOR2_X1 U11910 ( .A1(n10064), .A2(n10065), .ZN(n13047) );
  INV_X1 U11911 ( .A(n16789), .ZN(n19412) );
  NOR2_X1 U11912 ( .A1(n19409), .A2(n16789), .ZN(n15964) );
  NOR2_X1 U11913 ( .A1(n9598), .A2(n9835), .ZN(n9843) );
  NAND2_X1 U11914 ( .A1(n10127), .A2(n10126), .ZN(n10125) );
  INV_X1 U11915 ( .A(n11854), .ZN(n10127) );
  INV_X1 U11916 ( .A(n10124), .ZN(n10126) );
  OR2_X1 U11917 ( .A1(n9598), .A2(n13517), .ZN(n16061) );
  XNOR2_X1 U11918 ( .A(n12562), .B(n12561), .ZN(n14369) );
  INV_X1 U11919 ( .A(n14623), .ZN(n14630) );
  INV_X1 U11920 ( .A(n15580), .ZN(n16068) );
  NAND2_X1 U11921 ( .A1(n10112), .A2(n10433), .ZN(n16062) );
  INV_X1 U11922 ( .A(n10113), .ZN(n10112) );
  INV_X2 U11923 ( .A(n16137), .ZN(n19431) );
  INV_X1 U11924 ( .A(n16171), .ZN(n19437) );
  NAND2_X1 U11925 ( .A1(n19479), .A2(n13434), .ZN(n19445) );
  OR2_X1 U11926 ( .A1(n19479), .A2(n13396), .ZN(n13433) );
  XNOR2_X1 U11927 ( .A(n12568), .B(n12567), .ZN(n14357) );
  XNOR2_X1 U11928 ( .A(n16191), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13025) );
  INV_X1 U11929 ( .A(n19383), .ZN(n10073) );
  AND2_X1 U11930 ( .A1(n16436), .A2(n13019), .ZN(n16433) );
  OR2_X1 U11931 ( .A1(n19383), .A2(n10064), .ZN(n16439) );
  INV_X1 U11932 ( .A(n16436), .ZN(n16410) );
  XNOR2_X1 U11933 ( .A(n10197), .B(n9661), .ZN(n14348) );
  NAND2_X1 U11934 ( .A1(n10198), .A2(n9707), .ZN(n10197) );
  NOR2_X1 U11935 ( .A1(n14360), .A2(n12048), .ZN(n12587) );
  NAND2_X1 U11936 ( .A1(n9952), .A2(n9796), .ZN(n12558) );
  NAND2_X1 U11937 ( .A1(n12313), .A2(n12568), .ZN(n16177) );
  OAI211_X1 U11938 ( .C1(n16191), .C2(n10463), .A(n10462), .B(n10460), .ZN(
        n10214) );
  NAND2_X1 U11939 ( .A1(n12741), .A2(n12738), .ZN(n10056) );
  NAND2_X1 U11940 ( .A1(n9889), .A2(n12741), .ZN(n16466) );
  OR2_X1 U11941 ( .A1(n16202), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9889) );
  NAND2_X1 U11942 ( .A1(n9865), .A2(n16255), .ZN(n9802) );
  INV_X1 U11943 ( .A(n16237), .ZN(n9803) );
  AOI21_X1 U11944 ( .B1(n16262), .B2(n16250), .A(n16249), .ZN(n16254) );
  XNOR2_X1 U11945 ( .A(n16290), .B(n16532), .ZN(n16552) );
  XNOR2_X1 U11946 ( .A(n10539), .B(n16277), .ZN(n16556) );
  AND2_X1 U11947 ( .A1(n10534), .A2(n16276), .ZN(n10533) );
  NAND2_X1 U11948 ( .A1(n9832), .A2(n16290), .ZN(n16563) );
  NAND2_X1 U11949 ( .A1(n9833), .A2(n12454), .ZN(n9832) );
  AND2_X1 U11950 ( .A1(n16565), .A2(n16724), .ZN(n10079) );
  NAND2_X1 U11951 ( .A1(n10259), .A2(n10263), .ZN(n16308) );
  AND2_X1 U11952 ( .A1(n10013), .A2(n10260), .ZN(n16306) );
  NAND2_X1 U11953 ( .A1(n12554), .A2(n12317), .ZN(n16669) );
  AND2_X1 U11954 ( .A1(n12554), .A2(n20276), .ZN(n16689) );
  INV_X1 U11955 ( .A(n16689), .ZN(n16721) );
  NAND2_X1 U11956 ( .A1(n12554), .A2(n12201), .ZN(n16708) );
  NAND2_X1 U11957 ( .A1(n13903), .A2(n10063), .ZN(n12200) );
  INV_X1 U11958 ( .A(n16669), .ZN(n16727) );
  INV_X1 U11959 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20034) );
  INV_X1 U11960 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20271) );
  NOR2_X2 U11961 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20258) );
  NAND2_X1 U11962 ( .A1(n13692), .A2(n13633), .ZN(n20264) );
  NAND2_X1 U11963 ( .A1(n19353), .A2(n19153), .ZN(n17971) );
  AND2_X1 U11964 ( .A1(n10326), .A2(n10321), .ZN(n17119) );
  OR2_X1 U11965 ( .A1(n17124), .A2(n17123), .ZN(n17125) );
  INV_X1 U11966 ( .A(n17485), .ZN(n17468) );
  NOR2_X1 U11967 ( .A1(n17589), .A2(n17590), .ZN(n17574) );
  NOR2_X1 U11968 ( .A1(n17728), .A2(n17697), .ZN(n17713) );
  INV_X1 U11969 ( .A(n17756), .ZN(n17753) );
  INV_X1 U11970 ( .A(n17760), .ZN(n17775) );
  NOR2_X1 U11971 ( .A1(n16896), .A2(n10570), .ZN(n17779) );
  CLKBUF_X1 U11972 ( .A(n18038), .Z(n18030) );
  NOR2_X1 U11973 ( .A1(n12889), .A2(n13038), .ZN(n13026) );
  AND2_X1 U11974 ( .A1(n13276), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10181) );
  INV_X1 U11975 ( .A(n10081), .ZN(n13275) );
  INV_X1 U11976 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18407) );
  AND2_X1 U11977 ( .A1(n18504), .A2(n10346), .ZN(n18463) );
  AOI21_X1 U11978 ( .B1(n18703), .B2(n10349), .A(n10347), .ZN(n10346) );
  NAND2_X1 U11979 ( .A1(n18487), .A2(n18448), .ZN(n10349) );
  NOR2_X1 U11980 ( .A1(n19177), .A2(n10348), .ZN(n10347) );
  OAI21_X1 U11981 ( .B1(n18469), .B2(n18567), .A(n10342), .ZN(n10341) );
  AOI21_X1 U11982 ( .B1(n18479), .B2(n18468), .A(n18467), .ZN(n10342) );
  NAND2_X1 U11983 ( .A1(n18466), .A2(n10345), .ZN(n10344) );
  NAND2_X1 U11984 ( .A1(n18684), .A2(n18464), .ZN(n10345) );
  INV_X1 U11985 ( .A(n10274), .ZN(n10273) );
  OR2_X1 U11986 ( .A1(n19199), .A2(n10277), .ZN(n10276) );
  OAI21_X1 U11987 ( .B1(n19200), .B2(n19198), .A(n9709), .ZN(n10274) );
  INV_X1 U11988 ( .A(n19353), .ZN(n19212) );
  INV_X1 U11989 ( .A(n11879), .ZN(n10250) );
  INV_X1 U11990 ( .A(n10864), .ZN(n10141) );
  OAI21_X1 U11991 ( .B1(n11402), .B2(n11403), .A(n11401), .ZN(n9873) );
  NAND2_X1 U11992 ( .A1(n19693), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n9897) );
  NAND2_X1 U11993 ( .A1(n19990), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n9896) );
  NAND2_X1 U11994 ( .A1(n9621), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n9898) );
  NAND2_X1 U11995 ( .A1(n19727), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n9892) );
  NAND2_X1 U11996 ( .A1(n19919), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n9893) );
  NAND2_X1 U11997 ( .A1(n10017), .A2(n10016), .ZN(n11857) );
  NOR2_X1 U11998 ( .A1(n11810), .A2(n11777), .ZN(n11772) );
  OAI21_X1 U11999 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n19325), .A(
        n12712), .ZN(n12713) );
  OR2_X1 U12000 ( .A1(n12716), .A2(n12717), .ZN(n12712) );
  AND2_X1 U12001 ( .A1(n20933), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11392) );
  NAND2_X1 U12002 ( .A1(n20524), .A2(n10818), .ZN(n10825) );
  CLKBUF_X1 U12003 ( .A(n13148), .Z(n11287) );
  AND3_X1 U12004 ( .A1(n10967), .A2(n10949), .A3(n9717), .ZN(n11040) );
  INV_X1 U12005 ( .A(n11019), .ZN(n10036) );
  NAND2_X1 U12006 ( .A1(n15247), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10227) );
  OR2_X1 U12007 ( .A1(n11036), .A2(n11035), .ZN(n13224) );
  AND2_X1 U12008 ( .A1(n10230), .A2(n10847), .ZN(n10850) );
  AND2_X1 U12009 ( .A1(n10907), .A2(n10906), .ZN(n10923) );
  AND2_X1 U12010 ( .A1(n13189), .A2(n10144), .ZN(n9885) );
  INV_X1 U12011 ( .A(n10823), .ZN(n10237) );
  NAND2_X1 U12012 ( .A1(n14671), .A2(n11442), .ZN(n11448) );
  OAI21_X1 U12013 ( .B1(n13712), .B2(n10818), .A(n20532), .ZN(n11437) );
  NAND2_X1 U12014 ( .A1(n10820), .A2(n10846), .ZN(n11444) );
  INV_X1 U12015 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9816) );
  OR2_X1 U12016 ( .A1(n10947), .A2(n10946), .ZN(n13201) );
  OAI21_X1 U12017 ( .B1(n13304), .B2(n10840), .A(n13728), .ZN(n9859) );
  NAND2_X1 U12018 ( .A1(n14010), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10936) );
  NAND2_X1 U12019 ( .A1(n13222), .A2(n11398), .ZN(n11419) );
  INV_X1 U12020 ( .A(n12471), .ZN(n12447) );
  AND2_X2 U12021 ( .A1(n9906), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10046) );
  INV_X1 U12022 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9906) );
  AOI21_X1 U12023 ( .B1(n14598), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A(n9767), .ZN(n14585) );
  AOI21_X1 U12024 ( .B1(n14607), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A(n9772), .ZN(n14580) );
  AOI21_X1 U12025 ( .B1(n14607), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A(n9768), .ZN(n14550) );
  AOI21_X1 U12026 ( .B1(n14607), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A(n9769), .ZN(n14544) );
  AND2_X1 U12027 ( .A1(n10427), .A2(n9774), .ZN(n10105) );
  AOI21_X1 U12028 ( .B1(n14607), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A(n9740), .ZN(n14513) );
  AOI21_X1 U12029 ( .B1(n14601), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A(n9779), .ZN(n14456) );
  AOI21_X1 U12030 ( .B1(n14601), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A(n9743), .ZN(n14449) );
  AOI21_X1 U12031 ( .B1(n14601), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A(n9777), .ZN(n14491) );
  AND2_X1 U12032 ( .A1(n10405), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11821) );
  INV_X1 U12033 ( .A(n16230), .ZN(n10219) );
  INV_X1 U12034 ( .A(n10545), .ZN(n10544) );
  NAND2_X1 U12035 ( .A1(n9827), .A2(n11863), .ZN(n9829) );
  AND2_X1 U12036 ( .A1(n11879), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n9827) );
  AOI21_X1 U12037 ( .B1(n19759), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A(n9678), .ZN(n11917) );
  NAND2_X1 U12038 ( .A1(n10068), .A2(n10066), .ZN(n11634) );
  NAND2_X1 U12039 ( .A1(n10069), .A2(n11742), .ZN(n10068) );
  AND2_X1 U12040 ( .A1(n11794), .A2(n11741), .ZN(n12322) );
  AND2_X1 U12041 ( .A1(n11778), .A2(n11785), .ZN(n11792) );
  INV_X1 U12042 ( .A(n11786), .ZN(n11791) );
  NAND2_X1 U12043 ( .A1(n11880), .A2(n9620), .ZN(n11908) );
  AND2_X1 U12044 ( .A1(n11565), .A2(n11839), .ZN(n11567) );
  INV_X1 U12045 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11630) );
  INV_X1 U12046 ( .A(n14236), .ZN(n10186) );
  OAI22_X1 U12047 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19197), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12713), .ZN(n12718) );
  NAND2_X1 U12048 ( .A1(n10502), .A2(n14692), .ZN(n10501) );
  INV_X1 U12049 ( .A(n14708), .ZN(n10502) );
  NOR2_X1 U12050 ( .A1(n14787), .A2(n14769), .ZN(n10505) );
  OR2_X1 U12051 ( .A1(n14810), .A2(n10150), .ZN(n10149) );
  INV_X1 U12052 ( .A(n10566), .ZN(n10150) );
  AND2_X1 U12053 ( .A1(n11161), .A2(n11160), .ZN(n14902) );
  OR2_X1 U12054 ( .A1(n11090), .A2(n14128), .ZN(n14131) );
  AND2_X1 U12055 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n10585), .ZN(
        n11042) );
  NAND2_X1 U12056 ( .A1(n11020), .A2(n11018), .ZN(n13167) );
  NAND2_X1 U12057 ( .A1(n14703), .A2(n10473), .ZN(n10472) );
  INV_X1 U12058 ( .A(n14693), .ZN(n10473) );
  NOR2_X1 U12059 ( .A1(n10477), .A2(n14831), .ZN(n10476) );
  INV_X1 U12060 ( .A(n14842), .ZN(n10477) );
  NOR2_X1 U12061 ( .A1(n10920), .A2(n10144), .ZN(n13164) );
  INV_X1 U12062 ( .A(n13237), .ZN(n9927) );
  INV_X1 U12063 ( .A(n11481), .ZN(n10479) );
  INV_X1 U12064 ( .A(n11018), .ZN(n9857) );
  INV_X1 U12065 ( .A(n11020), .ZN(n9858) );
  NAND2_X1 U12066 ( .A1(n10152), .A2(n10151), .ZN(n13187) );
  AND2_X1 U12067 ( .A1(n13189), .A2(n9939), .ZN(n9938) );
  OR2_X1 U12068 ( .A1(n10917), .A2(n10916), .ZN(n13182) );
  NAND2_X1 U12069 ( .A1(n10031), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10935) );
  AND4_X2 U12070 ( .A1(n10731), .A2(n10730), .A3(n10729), .A4(n10728), .ZN(
        n10819) );
  NOR2_X1 U12071 ( .A1(n10561), .A2(n10715), .ZN(n10731) );
  OAI21_X1 U12072 ( .B1(n21179), .B2(n16996), .A(n21186), .ZN(n20496) );
  NAND2_X1 U12073 ( .A1(n10937), .A2(n10936), .ZN(n11432) );
  NAND2_X1 U12074 ( .A1(n9869), .A2(n9868), .ZN(n9867) );
  NAND2_X1 U12075 ( .A1(n11429), .A2(n11428), .ZN(n13301) );
  MUX2_X1 U12076 ( .A(n11930), .B(n11747), .S(n11800), .Z(n12375) );
  OAI21_X1 U12077 ( .B1(n15645), .B2(n16750), .A(n16207), .ZN(n15610) );
  AND2_X1 U12078 ( .A1(n12516), .A2(n12279), .ZN(n10454) );
  INV_X1 U12079 ( .A(n10451), .ZN(n9912) );
  NAND2_X1 U12080 ( .A1(n9909), .A2(n12373), .ZN(n12390) );
  NAND2_X1 U12081 ( .A1(n12372), .A2(n12532), .ZN(n9909) );
  NOR2_X1 U12082 ( .A1(n16740), .A2(n15951), .ZN(n15940) );
  NAND2_X1 U12083 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12285) );
  NAND2_X1 U12084 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12267) );
  INV_X1 U12085 ( .A(n13007), .ZN(n10491) );
  AND2_X1 U12086 ( .A1(n12747), .A2(n15593), .ZN(n10492) );
  AOI21_X1 U12087 ( .B1(n14607), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A(n9770), .ZN(n14571) );
  AOI21_X1 U12088 ( .B1(n14607), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(n9771), .ZN(n14565) );
  CLKBUF_X1 U12089 ( .A(n14454), .Z(n14606) );
  AOI21_X1 U12090 ( .B1(n14607), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A(n9741), .ZN(n14530) );
  AOI21_X1 U12091 ( .B1(n14607), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A(n9742), .ZN(n14524) );
  NAND2_X1 U12092 ( .A1(n14502), .A2(n10426), .ZN(n10424) );
  OR2_X1 U12093 ( .A1(n14502), .A2(n14537), .ZN(n10425) );
  NAND2_X1 U12094 ( .A1(n14431), .A2(n10123), .ZN(n10122) );
  INV_X1 U12095 ( .A(n16028), .ZN(n10123) );
  NOR2_X1 U12096 ( .A1(n10369), .A2(n16173), .ZN(n10366) );
  INV_X1 U12097 ( .A(n10368), .ZN(n10367) );
  NAND2_X1 U12098 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10368) );
  INV_X1 U12099 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10369) );
  NOR2_X1 U12100 ( .A1(n13120), .A2(n13022), .ZN(n13122) );
  NAND2_X1 U12101 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12281) );
  NOR2_X1 U12102 ( .A1(n13105), .A2(n16837), .ZN(n10380) );
  NAND2_X1 U12103 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12271) );
  NAND2_X1 U12104 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12248) );
  NAND2_X1 U12105 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12244) );
  NAND2_X1 U12106 ( .A1(n10542), .A2(n12542), .ZN(n10446) );
  INV_X1 U12107 ( .A(n12536), .ZN(n10542) );
  NOR2_X1 U12108 ( .A1(n10545), .A2(n12537), .ZN(n10543) );
  OR2_X1 U12109 ( .A1(n15616), .A2(n12048), .ZN(n16192) );
  NAND2_X1 U12110 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10514) );
  NAND2_X1 U12111 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12297) );
  INV_X1 U12112 ( .A(n15622), .ZN(n10420) );
  INV_X1 U12113 ( .A(n15652), .ZN(n9961) );
  NAND2_X1 U12114 ( .A1(n16267), .A2(n10255), .ZN(n10254) );
  NAND2_X1 U12115 ( .A1(n16374), .A2(n11977), .ZN(n9899) );
  AND2_X1 U12116 ( .A1(n12359), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10510) );
  AND2_X1 U12117 ( .A1(n12258), .A2(n10407), .ZN(n15717) );
  AND2_X1 U12118 ( .A1(n9632), .A2(n9758), .ZN(n10407) );
  INV_X1 U12119 ( .A(n14037), .ZN(n10488) );
  OR2_X1 U12120 ( .A1(n15812), .A2(n12048), .ZN(n12470) );
  NAND2_X1 U12121 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12238) );
  NAND2_X1 U12122 ( .A1(n10509), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9946) );
  AND2_X1 U12123 ( .A1(n11957), .A2(n11961), .ZN(n10382) );
  AND2_X1 U12124 ( .A1(n12045), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10210) );
  NAND2_X1 U12125 ( .A1(n10074), .A2(n12331), .ZN(n11783) );
  NAND2_X1 U12126 ( .A1(n11903), .A2(n11902), .ZN(n10356) );
  INV_X1 U12127 ( .A(n10211), .ZN(n11918) );
  NOR2_X1 U12128 ( .A1(n11670), .A2(n11669), .ZN(n11671) );
  INV_X1 U12129 ( .A(n11667), .ZN(n11670) );
  INV_X1 U12130 ( .A(n11668), .ZN(n11669) );
  AOI21_X1 U12131 ( .B1(n10074), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12004) );
  INV_X1 U12132 ( .A(n12045), .ZN(n12195) );
  NAND2_X1 U12133 ( .A1(n14556), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13623) );
  OAI21_X1 U12134 ( .B1(n13627), .B2(n13630), .A(n13629), .ZN(n13690) );
  NAND2_X1 U12135 ( .A1(n14556), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13688) );
  AND2_X1 U12136 ( .A1(n9836), .A2(n11856), .ZN(n11875) );
  INV_X1 U12137 ( .A(n11883), .ZN(n19919) );
  NAND3_X1 U12138 ( .A1(n20258), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20102), 
        .ZN(n16770) );
  AND2_X1 U12139 ( .A1(n19754), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13694) );
  XNOR2_X1 U12140 ( .A(n11839), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11623) );
  NAND2_X1 U12141 ( .A1(n11593), .A2(n11592), .ZN(n11625) );
  NAND2_X1 U12142 ( .A1(n12876), .A2(n17972), .ZN(n14231) );
  INV_X1 U12143 ( .A(n18181), .ZN(n10310) );
  NOR2_X1 U12144 ( .A1(n18222), .A2(n10312), .ZN(n10311) );
  NAND2_X1 U12145 ( .A1(n10081), .A2(n18228), .ZN(n10084) );
  NAND2_X1 U12146 ( .A1(n13027), .A2(n12971), .ZN(n12930) );
  NAND2_X1 U12147 ( .A1(n18045), .A2(n10304), .ZN(n10303) );
  NAND2_X1 U12148 ( .A1(n10088), .A2(n9810), .ZN(n9988) );
  AND2_X1 U12149 ( .A1(n10398), .A2(n9734), .ZN(n10088) );
  INV_X1 U12150 ( .A(n12863), .ZN(n9987) );
  INV_X1 U12151 ( .A(n18316), .ZN(n10399) );
  NAND2_X1 U12152 ( .A1(n9808), .A2(n9806), .ZN(n12857) );
  NAND2_X1 U12153 ( .A1(n9982), .A2(n9663), .ZN(n9806) );
  NAND2_X1 U12154 ( .A1(n9981), .A2(n9663), .ZN(n9808) );
  OAI211_X1 U12155 ( .C1(n17700), .C2(n10293), .A(n10292), .B(n9712), .ZN(
        n10291) );
  INV_X1 U12156 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U12157 ( .A1(n17733), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10292) );
  NOR2_X1 U12158 ( .A1(n12888), .A2(n12887), .ZN(n12952) );
  NOR2_X1 U12159 ( .A1(n10298), .A2(n17972), .ZN(n10297) );
  AND2_X1 U12160 ( .A1(n12695), .A2(n19360), .ZN(n10270) );
  OAI21_X1 U12161 ( .B1(n14231), .B2(n12886), .A(n12877), .ZN(n19161) );
  NAND2_X1 U12162 ( .A1(n19167), .A2(n12708), .ZN(n19173) );
  AOI221_X1 U12163 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19214), .C1(n18707), 
        .C2(P3_STATE2_REG_1__SCAN_IN), .A(n19337), .ZN(n18719) );
  NAND2_X1 U12164 ( .A1(n14013), .A2(n14010), .ZN(n10843) );
  INV_X1 U12165 ( .A(n10961), .ZN(n11023) );
  INV_X1 U12166 ( .A(n10843), .ZN(n14008) );
  NAND2_X1 U12167 ( .A1(n11465), .A2(n11464), .ZN(n11468) );
  OR2_X1 U12168 ( .A1(n14671), .A2(n11463), .ZN(n11464) );
  OAI21_X1 U12169 ( .B1(n9613), .B2(P1_EBX_REG_1__SCAN_IN), .A(n11462), .ZN(
        n11463) );
  AND2_X1 U12170 ( .A1(n11498), .A2(n11497), .ZN(n14112) );
  INV_X1 U12171 ( .A(n15503), .ZN(n11494) );
  AND2_X1 U12172 ( .A1(n11468), .A2(n10482), .ZN(n13755) );
  NAND2_X1 U12173 ( .A1(n13509), .A2(n21355), .ZN(n10482) );
  OR2_X1 U12174 ( .A1(n11372), .A2(n15056), .ZN(n10596) );
  AND2_X1 U12175 ( .A1(n10594), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11358) );
  AOI21_X1 U12176 ( .B1(n15079), .B2(n13162), .A(n11357), .ZN(n14720) );
  AND2_X1 U12177 ( .A1(n10593), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11340) );
  CLKBUF_X1 U12178 ( .A(n14718), .Z(n14719) );
  CLKBUF_X1 U12179 ( .A(n14731), .Z(n14743) );
  AND2_X1 U12180 ( .A1(n10592), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11322) );
  OR2_X1 U12181 ( .A1(n15102), .A2(n11371), .ZN(n11332) );
  AND2_X1 U12182 ( .A1(n11300), .A2(n10503), .ZN(n14752) );
  NAND2_X1 U12183 ( .A1(n11300), .A2(n10505), .ZN(n14767) );
  NAND2_X1 U12184 ( .A1(n11300), .A2(n11299), .ZN(n14766) );
  CLKBUF_X1 U12185 ( .A(n14784), .Z(n14785) );
  OR2_X1 U12186 ( .A1(n11208), .A2(n10590), .ZN(n11226) );
  NAND2_X1 U12187 ( .A1(n10589), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11208) );
  INV_X1 U12188 ( .A(n11175), .ZN(n10589) );
  NAND2_X1 U12189 ( .A1(n11137), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11175) );
  AND2_X1 U12190 ( .A1(n14907), .A2(n14884), .ZN(n14885) );
  INV_X1 U12191 ( .A(n11075), .ZN(n10586) );
  NAND2_X1 U12192 ( .A1(n11082), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11075) );
  NAND2_X1 U12193 ( .A1(n11023), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11043) );
  NOR2_X1 U12194 ( .A1(n10563), .A2(n11025), .ZN(n11026) );
  INV_X1 U12195 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10584) );
  OAI21_X1 U12196 ( .B1(n13251), .B2(n15236), .A(n14352), .ZN(n9826) );
  AND2_X1 U12197 ( .A1(n11547), .A2(n11546), .ZN(n14721) );
  AND2_X1 U12198 ( .A1(n9634), .A2(n14748), .ZN(n10483) );
  OR2_X1 U12199 ( .A1(n15099), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9943) );
  AND2_X1 U12200 ( .A1(n15236), .A2(n15343), .ZN(n9942) );
  NAND2_X1 U12201 ( .A1(n10247), .A2(n10059), .ZN(n15106) );
  NOR2_X1 U12202 ( .A1(n9699), .A2(n10583), .ZN(n10059) );
  NAND2_X1 U12203 ( .A1(n14799), .A2(n14783), .ZN(n14782) );
  NAND2_X1 U12204 ( .A1(n13249), .A2(n10555), .ZN(n15117) );
  AND2_X1 U12205 ( .A1(n10234), .A2(n13246), .ZN(n13249) );
  NAND2_X1 U12206 ( .A1(n14859), .A2(n10476), .ZN(n14829) );
  NAND2_X1 U12207 ( .A1(n14859), .A2(n14842), .ZN(n14843) );
  INV_X1 U12208 ( .A(n14873), .ZN(n10481) );
  OR2_X1 U12209 ( .A1(n15236), .A2(n13244), .ZN(n15176) );
  NAND2_X1 U12210 ( .A1(n14939), .A2(n9627), .ZN(n14889) );
  INV_X1 U12211 ( .A(n9933), .ZN(n15187) );
  AND2_X1 U12212 ( .A1(n10057), .A2(n16922), .ZN(n16918) );
  NAND2_X1 U12213 ( .A1(n9852), .A2(n13212), .ZN(n16925) );
  NAND2_X1 U12214 ( .A1(n11482), .A2(n11481), .ZN(n16975) );
  AOI21_X1 U12215 ( .B1(n15478), .B2(n15477), .A(n20460), .ZN(n16969) );
  NOR2_X1 U12216 ( .A1(n15469), .A2(n13760), .ZN(n15478) );
  AND2_X1 U12217 ( .A1(n15467), .A2(n13752), .ZN(n15493) );
  NAND2_X1 U12218 ( .A1(n15556), .A2(n13222), .ZN(n13180) );
  OR2_X1 U12219 ( .A1(n13472), .A2(n14647), .ZN(n13721) );
  AND2_X1 U12220 ( .A1(n13719), .A2(n13718), .ZN(n13738) );
  OAI21_X1 U12221 ( .B1(n13304), .B2(n14013), .A(n13454), .ZN(n13720) );
  NAND2_X1 U12222 ( .A1(n10985), .A2(n10144), .ZN(n10982) );
  INV_X1 U12223 ( .A(n10863), .ZN(n9923) );
  NAND2_X1 U12224 ( .A1(n10879), .A2(n10863), .ZN(n10035) );
  NAND2_X1 U12225 ( .A1(n10995), .A2(n15561), .ZN(n10060) );
  INV_X1 U12226 ( .A(n13254), .ZN(n16846) );
  OR3_X1 U12227 ( .A1(n13479), .A2(n13478), .A3(n13477), .ZN(n16849) );
  AND2_X1 U12228 ( .A1(n20611), .A2(n20934), .ZN(n20613) );
  NAND2_X1 U12229 ( .A1(n15562), .A2(n15561), .ZN(n20750) );
  NAND2_X1 U12230 ( .A1(n11432), .A2(n13301), .ZN(n11433) );
  OR2_X1 U12231 ( .A1(n11641), .A2(n11640), .ZN(n11643) );
  XNOR2_X1 U12232 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11675) );
  OAI21_X1 U12233 ( .B1(n20279), .B2(n11771), .A(n11755), .ZN(n13014) );
  NAND2_X1 U12234 ( .A1(n20275), .A2(n10070), .ZN(n11755) );
  AND2_X1 U12235 ( .A1(n13913), .A2(n10063), .ZN(n10070) );
  NAND2_X1 U12236 ( .A1(n12584), .A2(n12527), .ZN(n12534) );
  AOI21_X1 U12237 ( .B1(n15661), .B2(n19409), .A(n16216), .ZN(n15645) );
  AND2_X1 U12238 ( .A1(n12451), .A2(n12456), .ZN(n15721) );
  AND2_X1 U12239 ( .A1(n15738), .A2(n16287), .ZN(n15719) );
  NOR2_X1 U12240 ( .A1(n15796), .A2(n16334), .ZN(n15783) );
  NOR2_X1 U12241 ( .A1(n15849), .A2(n16386), .ZN(n15835) );
  NOR2_X1 U12242 ( .A1(n15906), .A2(n15908), .ZN(n15891) );
  NAND2_X1 U12243 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12235) );
  OR2_X1 U12244 ( .A1(n12062), .A2(n12061), .ZN(n13818) );
  NOR2_X1 U12245 ( .A1(n12209), .A2(n9751), .ZN(n10205) );
  AND2_X1 U12246 ( .A1(n15631), .A2(n10489), .ZN(n12562) );
  AND2_X1 U12247 ( .A1(n9773), .A2(n10490), .ZN(n10489) );
  INV_X1 U12248 ( .A(n12197), .ZN(n10490) );
  AOI21_X1 U12249 ( .B1(n14598), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n9786), .ZN(n14599) );
  AOI22_X1 U12250 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n14598), .ZN(n14615) );
  NOR2_X1 U12251 ( .A1(n10433), .A2(n10431), .ZN(n10430) );
  INV_X1 U12252 ( .A(n10437), .ZN(n10431) );
  NAND2_X1 U12253 ( .A1(n15981), .A2(n10432), .ZN(n10434) );
  NOR2_X1 U12254 ( .A1(n10433), .A2(n15983), .ZN(n10432) );
  NOR2_X1 U12255 ( .A1(n16008), .A2(n10063), .ZN(n16016) );
  AND2_X1 U12256 ( .A1(n16017), .A2(n16016), .ZN(n16019) );
  NOR2_X1 U12257 ( .A1(n16033), .A2(n10122), .ZN(n16030) );
  NAND2_X1 U12258 ( .A1(n10439), .A2(n16044), .ZN(n10438) );
  INV_X1 U12259 ( .A(n10440), .ZN(n10439) );
  NAND2_X1 U12260 ( .A1(n10115), .A2(n9649), .ZN(n10114) );
  NAND2_X1 U12261 ( .A1(n13764), .A2(n9692), .ZN(n10116) );
  INV_X1 U12262 ( .A(n10117), .ZN(n10115) );
  NAND2_X1 U12263 ( .A1(n10405), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12564) );
  AND2_X1 U12264 ( .A1(n12304), .A2(n12303), .ZN(n12743) );
  NAND2_X1 U12265 ( .A1(n13116), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13118) );
  NOR2_X1 U12266 ( .A1(n13113), .A2(n13112), .ZN(n13116) );
  NAND2_X1 U12267 ( .A1(n10380), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13113) );
  AND2_X1 U12268 ( .A1(n12291), .A2(n12290), .ZN(n16023) );
  NAND2_X1 U12269 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12263) );
  AND2_X1 U12270 ( .A1(n12262), .A2(n12261), .ZN(n15767) );
  INV_X1 U12271 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16332) );
  INV_X1 U12272 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15815) );
  AND2_X1 U12273 ( .A1(n10377), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10376) );
  AND2_X1 U12274 ( .A1(n12227), .A2(n12226), .ZN(n14098) );
  INV_X1 U12275 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13069) );
  NAND3_X1 U12276 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13066) );
  NAND2_X1 U12277 ( .A1(n12583), .A2(n14632), .ZN(n12585) );
  NOR2_X1 U12278 ( .A1(n12570), .A2(n12569), .ZN(n9951) );
  INV_X1 U12279 ( .A(n9794), .ZN(n10053) );
  NAND2_X1 U12280 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12310) );
  AND2_X1 U12281 ( .A1(n13060), .A2(n10444), .ZN(n12579) );
  AND2_X1 U12282 ( .A1(n12412), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10444) );
  AND2_X1 U12283 ( .A1(n15581), .A2(n12544), .ZN(n12991) );
  NAND2_X1 U12284 ( .A1(n10464), .A2(n12738), .ZN(n10459) );
  INV_X1 U12285 ( .A(n16211), .ZN(n10008) );
  NAND2_X1 U12286 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12277) );
  NAND2_X1 U12287 ( .A1(n10579), .A2(n10421), .ZN(n15640) );
  NAND2_X1 U12288 ( .A1(n16219), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16213) );
  NAND2_X1 U12289 ( .A1(n16204), .A2(n16484), .ZN(n10155) );
  NAND2_X1 U12290 ( .A1(n16203), .A2(n16220), .ZN(n10156) );
  NAND2_X1 U12291 ( .A1(n9961), .A2(n12183), .ZN(n15635) );
  INV_X1 U12292 ( .A(n16238), .ZN(n9905) );
  AND2_X1 U12293 ( .A1(n12359), .A2(n16655), .ZN(n16509) );
  INV_X1 U12294 ( .A(n15686), .ZN(n12176) );
  INV_X1 U12295 ( .A(n16264), .ZN(n10215) );
  NAND2_X1 U12296 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12275) );
  INV_X1 U12297 ( .A(n13777), .ZN(n9963) );
  NAND2_X1 U12298 ( .A1(n10535), .A2(n10536), .ZN(n10534) );
  NAND2_X1 U12299 ( .A1(n16267), .A2(n9954), .ZN(n9833) );
  INV_X1 U12300 ( .A(n16288), .ZN(n9954) );
  NAND2_X1 U12301 ( .A1(n10515), .A2(n10518), .ZN(n10263) );
  NAND2_X1 U12302 ( .A1(n10519), .A2(n16322), .ZN(n10518) );
  INV_X1 U12303 ( .A(n10521), .ZN(n10519) );
  NAND2_X1 U12304 ( .A1(n10261), .A2(n16307), .ZN(n10260) );
  INV_X1 U12305 ( .A(n10263), .ZN(n10261) );
  AND2_X1 U12306 ( .A1(n10515), .A2(n16307), .ZN(n10262) );
  AND2_X1 U12307 ( .A1(n12256), .A2(n12255), .ZN(n14194) );
  NAND2_X1 U12308 ( .A1(n12258), .A2(n12257), .ZN(n14193) );
  NAND2_X1 U12309 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12251) );
  AND2_X1 U12310 ( .A1(n16655), .A2(n16629), .ZN(n16616) );
  INV_X1 U12311 ( .A(n13826), .ZN(n12242) );
  AND2_X1 U12312 ( .A1(n12109), .A2(n12108), .ZN(n13745) );
  NOR2_X1 U12313 ( .A1(n9967), .A2(n9757), .ZN(n9966) );
  INV_X1 U12314 ( .A(n10487), .ZN(n9967) );
  AND2_X1 U12315 ( .A1(n12234), .A2(n12233), .ZN(n13957) );
  NAND2_X1 U12316 ( .A1(n10405), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12232) );
  NAND2_X1 U12317 ( .A1(n12229), .A2(n12228), .ZN(n14100) );
  AND2_X1 U12318 ( .A1(n15861), .A2(n12437), .ZN(n16389) );
  INV_X1 U12319 ( .A(n10363), .ZN(n10362) );
  AND2_X1 U12320 ( .A1(n12221), .A2(n13836), .ZN(n10415) );
  NOR2_X1 U12321 ( .A1(n13971), .A2(n14076), .ZN(n14072) );
  NAND2_X1 U12322 ( .A1(n14072), .A2(n14071), .ZN(n14074) );
  NAND2_X1 U12323 ( .A1(n12212), .A2(n12213), .ZN(n13804) );
  NAND2_X1 U12324 ( .A1(n10416), .A2(n10417), .ZN(n13845) );
  INV_X1 U12325 ( .A(n13804), .ZN(n10416) );
  AND2_X1 U12326 ( .A1(n12345), .A2(n13657), .ZN(n16694) );
  NOR2_X1 U12327 ( .A1(n16729), .A2(n12356), .ZN(n16693) );
  OAI211_X1 U12328 ( .C1(n12011), .C2(n12162), .A(n12010), .B(n12023), .ZN(
        n13547) );
  AND2_X1 U12329 ( .A1(n14605), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11890) );
  NAND2_X1 U12330 ( .A1(n9837), .A2(n13522), .ZN(n10423) );
  NAND2_X1 U12331 ( .A1(n16714), .A2(n9838), .ZN(n9837) );
  XNOR2_X1 U12332 ( .A(n13690), .B(n13688), .ZN(n13631) );
  AND2_X1 U12333 ( .A1(n13871), .A2(n13870), .ZN(n16744) );
  INV_X1 U12334 ( .A(n19755), .ZN(n19759) );
  INV_X1 U12335 ( .A(n19993), .ZN(n19723) );
  AND2_X1 U12336 ( .A1(n19598), .A2(n19597), .ZN(n19792) );
  INV_X1 U12337 ( .A(n20043), .ZN(n20039) );
  NAND2_X1 U12338 ( .A1(n11697), .A2(n11839), .ZN(n11704) );
  NOR2_X2 U12339 ( .A1(n16771), .A2(n16770), .ZN(n19575) );
  INV_X1 U12340 ( .A(n19576), .ZN(n19571) );
  INV_X1 U12341 ( .A(n19575), .ZN(n19573) );
  NOR2_X1 U12342 ( .A1(n20264), .A2(n19523), .ZN(n20098) );
  AND2_X1 U12343 ( .A1(n13694), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20105) );
  NOR2_X1 U12344 ( .A1(n13911), .A2(n10071), .ZN(n13912) );
  NAND2_X1 U12345 ( .A1(n10064), .A2(n10072), .ZN(n10071) );
  INV_X1 U12346 ( .A(n16810), .ZN(n10072) );
  AND2_X1 U12347 ( .A1(n16742), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13352) );
  INV_X1 U12348 ( .A(n10314), .ZN(n17166) );
  OAI21_X1 U12350 ( .B1(n10319), .B2(n10316), .A(n10318), .ZN(n10315) );
  NAND2_X1 U12351 ( .A1(n10308), .A2(n10307), .ZN(n10306) );
  INV_X1 U12352 ( .A(n18124), .ZN(n10307) );
  NOR2_X1 U12353 ( .A1(n19270), .A2(n17254), .ZN(n17228) );
  NAND2_X1 U12354 ( .A1(n17327), .A2(n12590), .ZN(n17330) );
  INV_X1 U12355 ( .A(n18250), .ZN(n12590) );
  NAND2_X1 U12356 ( .A1(n17574), .A2(n9656), .ZN(n17539) );
  INV_X1 U12357 ( .A(n17617), .ZN(n10332) );
  NOR2_X1 U12358 ( .A1(n17999), .A2(n17997), .ZN(n10188) );
  NOR2_X1 U12359 ( .A1(n12676), .A2(n12675), .ZN(n17785) );
  NOR2_X1 U12360 ( .A1(n12818), .A2(n10086), .ZN(n10085) );
  NOR2_X1 U12361 ( .A1(n14229), .A2(n12710), .ZN(n10400) );
  NAND2_X1 U12362 ( .A1(n12812), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12806) );
  OAI21_X1 U12363 ( .B1(n16898), .B2(n16897), .A(n19353), .ZN(n16899) );
  NOR2_X1 U12364 ( .A1(n12697), .A2(n18749), .ZN(n19183) );
  AND2_X1 U12365 ( .A1(n10323), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10322) );
  INV_X1 U12366 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12596) );
  NOR2_X1 U12367 ( .A1(n18514), .A2(n18080), .ZN(n18428) );
  INV_X1 U12368 ( .A(n18205), .ZN(n18189) );
  NAND2_X1 U12369 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18250) );
  NOR2_X2 U12370 ( .A1(n18314), .A2(n18318), .ZN(n18286) );
  NOR2_X1 U12371 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18707), .ZN(n18219) );
  INV_X1 U12372 ( .A(n10084), .ZN(n12934) );
  NAND2_X1 U12373 ( .A1(n16888), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16887) );
  NAND2_X1 U12374 ( .A1(n12870), .A2(n9974), .ZN(n9973) );
  AND2_X1 U12375 ( .A1(n10304), .A2(n18047), .ZN(n9974) );
  NOR2_X1 U12376 ( .A1(n18069), .A2(n12919), .ZN(n18389) );
  NAND2_X1 U12377 ( .A1(n12870), .A2(n10304), .ZN(n18071) );
  NOR2_X1 U12378 ( .A1(n18449), .A2(n18461), .ZN(n10348) );
  OAI21_X1 U12379 ( .B1(n9616), .B2(n18512), .A(n9650), .ZN(n10177) );
  NAND2_X1 U12380 ( .A1(n18292), .A2(n9616), .ZN(n10178) );
  INV_X1 U12381 ( .A(n18261), .ZN(n12865) );
  XNOR2_X1 U12382 ( .A(n12910), .B(n12912), .ZN(n10000) );
  XNOR2_X1 U12383 ( .A(n9988), .B(n9987), .ZN(n18302) );
  INV_X1 U12384 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18306) );
  INV_X1 U12385 ( .A(n12907), .ZN(n10339) );
  NOR2_X1 U12386 ( .A1(n18324), .A2(n18647), .ZN(n18325) );
  NOR2_X1 U12387 ( .A1(n17785), .A2(n12947), .ZN(n12959) );
  OAI21_X1 U12388 ( .B1(n12721), .B2(n12881), .A(n12875), .ZN(n12950) );
  NAND2_X1 U12389 ( .A1(n19169), .A2(n19177), .ZN(n18684) );
  AND4_X1 U12390 ( .A1(n12847), .A2(n12846), .A3(n12845), .A4(n12844), .ZN(
        n12848) );
  INV_X2 U12391 ( .A(n12822), .ZN(n17738) );
  NOR2_X1 U12392 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18719), .ZN(n19010) );
  AOI22_X1 U12393 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12665) );
  AOI211_X1 U12394 ( .C1(n17570), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n12663), .B(n12662), .ZN(n12664) );
  NAND3_X1 U12395 ( .A1(n12656), .A2(n12655), .A3(n12654), .ZN(n18736) );
  AOI22_X1 U12396 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12843), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12655) );
  AOI211_X1 U12397 ( .C1(n17570), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n12684), .B(n12683), .ZN(n12685) );
  INV_X1 U12398 ( .A(n19010), .ZN(n19063) );
  OR2_X1 U12399 ( .A1(n19201), .A2(n19202), .ZN(n10275) );
  NAND2_X1 U12400 ( .A1(n10265), .A2(n19181), .ZN(n10264) );
  AND2_X1 U12401 ( .A1(n19200), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10277) );
  NOR3_X1 U12402 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19239), .A3(n19224), 
        .ZN(n19228) );
  INV_X1 U12403 ( .A(n13718), .ZN(n20288) );
  NAND2_X1 U12404 ( .A1(n14025), .A2(n14023), .ZN(n20354) );
  NOR2_X1 U12405 ( .A1(n20354), .A2(n14814), .ZN(n20308) );
  OR3_X1 U12406 ( .A1(n21173), .A2(n16962), .A3(n14014), .ZN(n20345) );
  XNOR2_X1 U12407 ( .A(n11468), .B(n13509), .ZN(n14041) );
  INV_X1 U12408 ( .A(n20369), .ZN(n20336) );
  NAND2_X1 U12409 ( .A1(n14799), .A2(n10485), .ZN(n14755) );
  INV_X1 U12410 ( .A(n15045), .ZN(n10133) );
  CLKBUF_X1 U12411 ( .A(n13319), .Z(n15018) );
  INV_X1 U12412 ( .A(n14973), .ZN(n15017) );
  INV_X1 U12413 ( .A(n15031), .ZN(n15041) );
  NOR2_X1 U12414 ( .A1(n15041), .A2(n13747), .ZN(n15043) );
  NAND2_X2 U12415 ( .A1(n15031), .A2(n13747), .ZN(n15045) );
  INV_X1 U12416 ( .A(n15043), .ZN(n15034) );
  OR2_X1 U12417 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16998), .ZN(n20410) );
  AND2_X1 U12418 ( .A1(n13557), .A2(n16874), .ZN(n20408) );
  OAI21_X1 U12419 ( .B1(n13556), .B2(n21184), .A(n13588), .ZN(n13557) );
  INV_X2 U12420 ( .A(n20410), .ZN(n21176) );
  XNOR2_X1 U12421 ( .A(n14004), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14353) );
  NOR2_X1 U12422 ( .A1(n14003), .A2(n14002), .ZN(n14004) );
  AOI21_X2 U12423 ( .B1(n14708), .B2(n14707), .A(n14691), .ZN(n15075) );
  INV_X1 U12424 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15143) );
  CLKBUF_X1 U12425 ( .A(n14827), .Z(n14828) );
  NOR2_X1 U12426 ( .A1(n15040), .A2(n15039), .ZN(n20384) );
  XNOR2_X1 U12427 ( .A(n14655), .B(n14654), .ZN(n15283) );
  NAND3_X1 U12428 ( .A1(n10467), .A2(n10466), .A3(n10468), .ZN(n14655) );
  NAND2_X1 U12429 ( .A1(n14352), .A2(n9703), .ZN(n10042) );
  OAI21_X1 U12430 ( .B1(n9710), .B2(n15080), .A(n15081), .ZN(n15082) );
  XNOR2_X1 U12431 ( .A(n9940), .B(n15327), .ZN(n15334) );
  NAND2_X1 U12432 ( .A1(n9944), .A2(n9941), .ZN(n9940) );
  OR2_X1 U12433 ( .A1(n15095), .A2(n15343), .ZN(n9944) );
  AOI21_X1 U12434 ( .B1(n9943), .B2(n10583), .A(n9942), .ZN(n9941) );
  XNOR2_X1 U12435 ( .A(n9856), .B(n15343), .ZN(n15335) );
  NAND2_X1 U12436 ( .A1(n10242), .A2(n10241), .ZN(n9856) );
  NAND3_X1 U12437 ( .A1(n10244), .A2(n10583), .A3(n10243), .ZN(n10242) );
  NAND2_X1 U12438 ( .A1(n15372), .A2(n15264), .ZN(n15350) );
  NAND2_X1 U12439 ( .A1(n15151), .A2(n13246), .ZN(n10390) );
  OAI21_X1 U12440 ( .B1(n9931), .B2(n10583), .A(n9929), .ZN(n15155) );
  NAND2_X1 U12441 ( .A1(n9931), .A2(n9930), .ZN(n9929) );
  OAI21_X1 U12442 ( .B1(n9933), .B2(n9932), .A(n15153), .ZN(n9931) );
  AND2_X1 U12443 ( .A1(n15467), .A2(n15259), .ZN(n15459) );
  INV_X1 U12444 ( .A(n15151), .ZN(n15217) );
  NOR2_X1 U12445 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20477), .ZN(
        n13760) );
  AND2_X1 U12446 ( .A1(n13738), .A2(n15526), .ZN(n20477) );
  INV_X1 U12447 ( .A(n10974), .ZN(n10976) );
  INV_X1 U12448 ( .A(n20934), .ZN(n21010) );
  OR2_X1 U12449 ( .A1(n16883), .A2(n20782), .ZN(n21186) );
  INV_X1 U12450 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n21245) );
  OAI22_X1 U12451 ( .A1(n20505), .A2(n20504), .B1(n20777), .B2(n20646), .ZN(
        n20536) );
  OAI21_X1 U12452 ( .B1(n20547), .B2(n20546), .A(n21018), .ZN(n20567) );
  OAI21_X1 U12453 ( .B1(n20646), .B2(n20976), .A(n20645), .ZN(n20666) );
  INV_X1 U12454 ( .A(n20697), .ZN(n20688) );
  INV_X1 U12455 ( .A(n20735), .ZN(n20693) );
  NAND2_X1 U12456 ( .A1(n20533), .A2(n10818), .ZN(n20729) );
  OAI22_X1 U12457 ( .A1(n20706), .A2(n20705), .B1(n20704), .B2(n20976), .ZN(
        n20737) );
  OAI211_X1 U12458 ( .C1(n20798), .C2(n20782), .A(n20842), .B(n20781), .ZN(
        n20800) );
  AND2_X1 U12459 ( .A1(n20872), .A2(n20977), .ZN(n20896) );
  OAI211_X1 U12460 ( .C1(n20907), .C2(n21074), .A(n20985), .B(n20906), .ZN(
        n20928) );
  OAI21_X1 U12461 ( .B1(n20938), .B2(n20937), .A(n21018), .ZN(n20971) );
  OAI211_X1 U12462 ( .C1(n21002), .C2(n20986), .A(n20985), .B(n20984), .ZN(
        n21004) );
  INV_X1 U12463 ( .A(n20698), .ZN(n21014) );
  INV_X1 U12464 ( .A(n20709), .ZN(n21025) );
  INV_X1 U12465 ( .A(n20713), .ZN(n21031) );
  INV_X1 U12466 ( .A(n20717), .ZN(n21037) );
  INV_X1 U12467 ( .A(n20721), .ZN(n21043) );
  INV_X1 U12468 ( .A(n20725), .ZN(n21049) );
  INV_X1 U12469 ( .A(n20729), .ZN(n21055) );
  NOR2_X2 U12470 ( .A1(n21017), .A2(n20749), .ZN(n21065) );
  INV_X1 U12471 ( .A(n20733), .ZN(n21063) );
  NOR2_X1 U12472 ( .A1(n21185), .A2(n21074), .ZN(n16996) );
  NOR2_X1 U12473 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21179) );
  INV_X1 U12474 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n21185) );
  INV_X1 U12475 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20782) );
  INV_X1 U12476 ( .A(n21157), .ZN(n21153) );
  NAND2_X1 U12477 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n21175) );
  NAND2_X1 U12478 ( .A1(n15976), .A2(n19414), .ZN(n10374) );
  NAND2_X1 U12479 ( .A1(n12519), .A2(n12518), .ZN(n12541) );
  OR2_X1 U12480 ( .A1(n9684), .A2(n12521), .ZN(n12523) );
  INV_X1 U12481 ( .A(n15964), .ZN(n16833) );
  INV_X1 U12482 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16837) );
  INV_X1 U12483 ( .A(n16257), .ZN(n10370) );
  NAND2_X1 U12484 ( .A1(n10222), .A2(n10221), .ZN(n12453) );
  NAND2_X1 U12485 ( .A1(n10223), .A2(n12543), .ZN(n10222) );
  NAND2_X1 U12486 ( .A1(n12463), .A2(n12532), .ZN(n10221) );
  NAND2_X1 U12487 ( .A1(n12482), .A2(n10224), .ZN(n12477) );
  INV_X1 U12488 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n21330) );
  AND2_X1 U12489 ( .A1(n9835), .A2(n19414), .ZN(n15956) );
  INV_X1 U12490 ( .A(n19424), .ZN(n15963) );
  NAND2_X1 U12491 ( .A1(n19409), .A2(n19412), .ZN(n15975) );
  OR2_X1 U12492 ( .A1(n12104), .A2(n12103), .ZN(n14186) );
  NAND2_X1 U12493 ( .A1(n10063), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13499) );
  AND2_X1 U12494 ( .A1(n9959), .A2(n15595), .ZN(n16443) );
  OR2_X1 U12495 ( .A1(n15594), .A2(n15593), .ZN(n9959) );
  NAND2_X1 U12496 ( .A1(n15989), .A2(n15988), .ZN(n15987) );
  NOR2_X1 U12497 ( .A1(n15994), .A2(n10063), .ZN(n15995) );
  OR2_X1 U12498 ( .A1(n19431), .A2(n13535), .ZN(n16138) );
  INV_X1 U12499 ( .A(n19441), .ZN(n14122) );
  NAND2_X1 U12500 ( .A1(n10118), .A2(n13765), .ZN(n13770) );
  AND2_X1 U12501 ( .A1(n16138), .A2(n14366), .ZN(n19441) );
  OAI21_X1 U12502 ( .B1(n13868), .B2(n13393), .A(n13392), .ZN(n13394) );
  INV_X1 U12503 ( .A(n19445), .ZN(n19477) );
  INV_X1 U12504 ( .A(n13434), .ZN(n19476) );
  INV_X2 U12505 ( .A(n13366), .ZN(n19518) );
  INV_X2 U12506 ( .A(n13392), .ZN(n19517) );
  OR2_X1 U12507 ( .A1(n12997), .A2(n12996), .ZN(n16185) );
  INV_X1 U12508 ( .A(n9833), .ZN(n16300) );
  NAND2_X1 U12509 ( .A1(n16593), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10364) );
  INV_X1 U12510 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n21303) );
  INV_X1 U12511 ( .A(n16449), .ZN(n9957) );
  NOR2_X1 U12512 ( .A1(n16450), .A2(n16669), .ZN(n9956) );
  NAND2_X1 U12513 ( .A1(n16443), .A2(n16724), .ZN(n9958) );
  NOR2_X1 U12514 ( .A1(n16471), .A2(n16484), .ZN(n10513) );
  AND2_X1 U12515 ( .A1(n10200), .A2(n10199), .ZN(n16241) );
  OAI21_X1 U12516 ( .B1(n16237), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n16231), .ZN(n16518) );
  INV_X1 U12517 ( .A(n10216), .ZN(n16261) );
  AND2_X1 U12518 ( .A1(n16301), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10164) );
  OAI21_X1 U12519 ( .B1(n16354), .B2(n10521), .A(n10520), .ZN(n16324) );
  INV_X1 U12520 ( .A(n16310), .ZN(n16317) );
  NAND2_X1 U12521 ( .A1(n10523), .A2(n10527), .ZN(n16328) );
  NAND2_X1 U12522 ( .A1(n16354), .A2(n10529), .ZN(n10523) );
  OR2_X1 U12523 ( .A1(n13777), .A2(n13852), .ZN(n13998) );
  NAND2_X1 U12524 ( .A1(n16381), .A2(n10206), .ZN(n16664) );
  NAND2_X1 U12525 ( .A1(n16289), .A2(n16654), .ZN(n10206) );
  INV_X1 U12526 ( .A(n16267), .ZN(n16289) );
  NAND2_X1 U12527 ( .A1(n13528), .A2(n13529), .ZN(n13638) );
  INV_X1 U12528 ( .A(n10252), .ZN(n14200) );
  NAND2_X1 U12529 ( .A1(n13661), .A2(n12029), .ZN(n13973) );
  OAI21_X1 U12530 ( .B1(n16669), .B2(n10020), .A(n14635), .ZN(n13666) );
  INV_X1 U12531 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16742) );
  NAND2_X1 U12532 ( .A1(n9839), .A2(n13890), .ZN(n16755) );
  NAND2_X1 U12533 ( .A1(n9835), .A2(n9840), .ZN(n9839) );
  AND2_X1 U12534 ( .A1(n13905), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16752) );
  NOR2_X1 U12535 ( .A1(n10020), .A2(n13891), .ZN(n13863) );
  NOR2_X1 U12536 ( .A1(n16810), .A2(n20253), .ZN(n10076) );
  OR2_X1 U12537 ( .A1(n19592), .A2(n19589), .ZN(n19620) );
  INV_X1 U12538 ( .A(n19631), .ZN(n19652) );
  OAI21_X1 U12539 ( .B1(n19699), .B2(n19695), .A(n19694), .ZN(n19718) );
  OAI21_X1 U12540 ( .B1(n19730), .B2(n19726), .A(n19725), .ZN(n19749) );
  AND2_X1 U12541 ( .A1(n19753), .A2(n19723), .ZN(n19747) );
  AND2_X1 U12542 ( .A1(n19726), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19746) );
  OR2_X1 U12543 ( .A1(n19789), .A2(n19786), .ZN(n19813) );
  OAI21_X1 U12544 ( .B1(n20257), .B2(n19791), .A(n19790), .ZN(n19816) );
  INV_X1 U12545 ( .A(n19883), .ZN(n19849) );
  OR2_X1 U12546 ( .A1(n19988), .A2(n19857), .ZN(n19895) );
  OAI21_X1 U12547 ( .B1(n19863), .B2(n19862), .A(n19861), .ZN(n19885) );
  NAND2_X1 U12548 ( .A1(n10024), .A2(n20102), .ZN(n19915) );
  OAI21_X1 U12549 ( .B1(n10026), .B2(n10251), .A(n10025), .ZN(n10024) );
  INV_X1 U12550 ( .A(n19912), .ZN(n10025) );
  OAI21_X1 U12551 ( .B1(n19893), .B2(n19892), .A(n19891), .ZN(n19913) );
  OR2_X1 U12552 ( .A1(n20031), .A2(n19657), .ZN(n19955) );
  AND2_X1 U12553 ( .A1(n19578), .A2(n11785), .ZN(n19958) );
  INV_X1 U12554 ( .A(n20124), .ZN(n19963) );
  AND2_X1 U12555 ( .A1(n19578), .A2(n19553), .ZN(n19968) );
  OAI22_X1 U12556 ( .A1(n19552), .A2(n19571), .B1(n19551), .B2(n19573), .ZN(
        n19969) );
  OAI22_X1 U12557 ( .A1(n19565), .A2(n19571), .B1(n19564), .B2(n19573), .ZN(
        n19977) );
  OAI21_X1 U12558 ( .B1(n16776), .B2(n19695), .A(n16775), .ZN(n19982) );
  INV_X1 U12559 ( .A(n20113), .ZN(n20006) );
  OAI21_X1 U12560 ( .B1(n19999), .B2(n19998), .A(n19997), .ZN(n20026) );
  AND2_X1 U12561 ( .A1(n20102), .A2(n16777), .ZN(n20048) );
  AND2_X1 U12562 ( .A1(n19578), .A2(n10063), .ZN(n20052) );
  AND2_X1 U12563 ( .A1(n20102), .A2(n19542), .ZN(n20057) );
  AND2_X1 U12564 ( .A1(n20102), .A2(n19548), .ZN(n20063) );
  AND2_X1 U12565 ( .A1(n20102), .A2(n19555), .ZN(n20069) );
  AND2_X1 U12566 ( .A1(n20102), .A2(n19561), .ZN(n20074) );
  AND2_X1 U12567 ( .A1(n20102), .A2(n19568), .ZN(n20081) );
  AND2_X1 U12568 ( .A1(n19578), .A2(n19577), .ZN(n20084) );
  OAI222_X1 U12569 ( .A1(n20047), .A2(n20046), .B1(n20078), .B2(n20045), .C1(
        n20044), .C2(n20043), .ZN(n20086) );
  AND2_X1 U12570 ( .A1(n20102), .A2(n19581), .ZN(n20087) );
  INV_X1 U12571 ( .A(n19894), .ZN(n20094) );
  INV_X1 U12572 ( .A(n20052), .ZN(n20110) );
  INV_X1 U12573 ( .A(n19958), .ZN(n20117) );
  INV_X1 U12574 ( .A(n19968), .ZN(n20131) );
  INV_X1 U12575 ( .A(n19969), .ZN(n20137) );
  INV_X1 U12576 ( .A(n19976), .ZN(n20145) );
  INV_X1 U12577 ( .A(n19977), .ZN(n20153) );
  INV_X1 U12578 ( .A(n20084), .ZN(n20154) );
  OR2_X1 U12579 ( .A1(n20100), .A2(n20093), .ZN(n20157) );
  INV_X1 U12580 ( .A(n20105), .ZN(n20155) );
  OAI22_X1 U12581 ( .A1(n19574), .A2(n19573), .B1(n19572), .B2(n19571), .ZN(
        n20159) );
  NAND2_X1 U12582 ( .A1(n13352), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19381) );
  AND3_X1 U12583 ( .A1(n13930), .A2(n15577), .A3(n13929), .ZN(n14057) );
  INV_X1 U12584 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20167) );
  OR2_X1 U12585 ( .A1(n17128), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n13270) );
  INV_X1 U12586 ( .A(n10326), .ZN(n17136) );
  NAND2_X1 U12587 ( .A1(n10320), .A2(n10321), .ZN(n17176) );
  INV_X1 U12588 ( .A(n17462), .ZN(n17474) );
  AOI21_X2 U12589 ( .B1(n10321), .B2(n17241), .A(n17266), .ZN(n17243) );
  NAND2_X1 U12590 ( .A1(n12723), .A2(n19372), .ZN(n17485) );
  INV_X1 U12591 ( .A(n17408), .ZN(n17482) );
  AND2_X1 U12592 ( .A1(n17574), .A2(n10329), .ZN(n17538) );
  AND2_X1 U12593 ( .A1(n9656), .A2(n10330), .ZN(n10329) );
  NOR2_X1 U12594 ( .A1(n17535), .A2(n17171), .ZN(n10330) );
  NOR2_X1 U12595 ( .A1(n17201), .A2(n17576), .ZN(n10331) );
  AND2_X1 U12596 ( .A1(n16802), .A2(n9792), .ZN(n17604) );
  NAND2_X1 U12597 ( .A1(n16802), .A2(n9657), .ZN(n17615) );
  NOR2_X1 U12598 ( .A1(n17321), .A2(n17671), .ZN(n16802) );
  NAND2_X1 U12599 ( .A1(n16802), .A2(P3_EBX_REG_13__SCAN_IN), .ZN(n17657) );
  NAND2_X1 U12600 ( .A1(n17753), .A2(n9654), .ZN(n17728) );
  AND2_X1 U12601 ( .A1(n17753), .A2(P3_EBX_REG_6__SCAN_IN), .ZN(n17749) );
  AND2_X1 U12602 ( .A1(n17779), .A2(n14225), .ZN(n17757) );
  INV_X1 U12603 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17763) );
  INV_X1 U12604 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17774) );
  NOR2_X1 U12605 ( .A1(n12644), .A2(n10191), .ZN(n10190) );
  AND2_X1 U12606 ( .A1(n17811), .A2(n9797), .ZN(n17792) );
  NAND2_X1 U12607 ( .A1(n17811), .A2(n9658), .ZN(n17799) );
  NAND2_X1 U12608 ( .A1(n17811), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n17807) );
  NOR2_X1 U12609 ( .A1(n17995), .A2(n17817), .ZN(n17811) );
  NOR3_X1 U12610 ( .A1(n17860), .A2(n17827), .A3(n17784), .ZN(n17822) );
  INV_X1 U12611 ( .A(n17839), .ZN(n17835) );
  NOR3_X1 U12612 ( .A1(n17826), .A2(n17860), .A3(n17979), .ZN(n17849) );
  NAND2_X1 U12613 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17867), .ZN(n17860) );
  NOR2_X1 U12614 ( .A1(n17871), .A2(n18042), .ZN(n17867) );
  NAND2_X1 U12615 ( .A1(n16900), .A2(n10193), .ZN(n17871) );
  AND2_X1 U12616 ( .A1(n17864), .A2(n9617), .ZN(n10193) );
  NOR2_X1 U12617 ( .A1(n18025), .A2(n17898), .ZN(n17895) );
  AND2_X1 U12618 ( .A1(n16900), .A2(n9617), .ZN(n17899) );
  INV_X1 U12619 ( .A(n12891), .ZN(n17912) );
  AND2_X1 U12620 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17919), .ZN(n17914) );
  NOR2_X1 U12621 ( .A1(n18013), .A2(n17924), .ZN(n17919) );
  NOR2_X1 U12622 ( .A1(n12696), .A2(n16899), .ZN(n17921) );
  NOR2_X1 U12623 ( .A1(n12792), .A2(n12791), .ZN(n12797) );
  INV_X2 U12624 ( .A(n17921), .ZN(n17930) );
  INV_X1 U12625 ( .A(n17917), .ZN(n17927) );
  INV_X1 U12626 ( .A(n17928), .ZN(n17920) );
  NAND2_X1 U12627 ( .A1(n19354), .A2(n17970), .ZN(n17950) );
  INV_X1 U12628 ( .A(n17936), .ZN(n17952) );
  NOR2_X1 U12629 ( .A1(n19360), .A2(n18030), .ZN(n18031) );
  OAI211_X1 U12630 ( .C1(n19360), .C2(n19361), .A(n17975), .B(n17974), .ZN(
        n18038) );
  AOI21_X1 U12632 ( .B1(n18062), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n18050), .ZN(n18051) );
  NOR2_X1 U12633 ( .A1(n18049), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n18050) );
  AND2_X1 U12634 ( .A1(n18053), .A2(n9788), .ZN(n10289) );
  INV_X1 U12635 ( .A(n18399), .ZN(n18052) );
  NOR2_X2 U12636 ( .A1(n19214), .A2(n18374), .ZN(n18140) );
  INV_X1 U12637 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18318) );
  NOR2_X2 U12638 ( .A1(n18339), .A2(n18347), .ZN(n18323) );
  NAND2_X1 U12639 ( .A1(n19010), .A2(n18781), .ZN(n19061) );
  NAND2_X1 U12640 ( .A1(n18239), .A2(n18169), .ZN(n18343) );
  INV_X1 U12641 ( .A(n19061), .ZN(n19036) );
  INV_X1 U12642 ( .A(n18343), .ZN(n18378) );
  INV_X1 U12643 ( .A(n18371), .ZN(n18385) );
  INV_X1 U12644 ( .A(n18375), .ZN(n18384) );
  AND2_X1 U12645 ( .A1(n10296), .A2(n19169), .ZN(n18608) );
  NOR2_X1 U12646 ( .A1(n18703), .A2(n10298), .ZN(n10296) );
  NAND2_X1 U12647 ( .A1(n9993), .A2(n18403), .ZN(n9992) );
  INV_X1 U12648 ( .A(n13027), .ZN(n9993) );
  AND2_X1 U12649 ( .A1(n13032), .A2(n9990), .ZN(n9989) );
  NAND2_X1 U12650 ( .A1(n16818), .A2(n19150), .ZN(n9990) );
  AND2_X1 U12651 ( .A1(n10169), .A2(n10386), .ZN(n10174) );
  NAND2_X1 U12652 ( .A1(n12870), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10175) );
  INV_X1 U12653 ( .A(n10170), .ZN(n18087) );
  NOR2_X1 U12654 ( .A1(n18121), .A2(n12973), .ZN(n18096) );
  AOI221_X1 U12655 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18145), 
        .C1(n18141), .C2(n18162), .A(n18133), .ZN(n18134) );
  AND2_X1 U12656 ( .A1(n10351), .A2(n10350), .ZN(n18504) );
  NAND2_X1 U12657 ( .A1(n18514), .A2(n18571), .ZN(n10350) );
  NAND2_X1 U12658 ( .A1(n18523), .A2(n19150), .ZN(n10351) );
  INV_X1 U12659 ( .A(n18567), .ZN(n18616) );
  AND2_X1 U12660 ( .A1(n9997), .A2(n9998), .ZN(n18327) );
  NAND2_X1 U12661 ( .A1(n10280), .A2(n10279), .ZN(n18341) );
  INV_X1 U12662 ( .A(n9981), .ZN(n10280) );
  NAND2_X1 U12663 ( .A1(n18352), .A2(n18353), .ZN(n18351) );
  INV_X1 U12664 ( .A(n10302), .ZN(n18352) );
  INV_X1 U12665 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18682) );
  AND2_X1 U12666 ( .A1(n9813), .A2(n9812), .ZN(n18683) );
  NAND2_X1 U12667 ( .A1(n18373), .A2(n18372), .ZN(n9812) );
  INV_X1 U12668 ( .A(n18700), .ZN(n18693) );
  INV_X1 U12669 ( .A(n12963), .ZN(n18702) );
  NOR2_X1 U12670 ( .A1(n19155), .A2(n18702), .ZN(n18700) );
  AND2_X1 U12671 ( .A1(n19370), .A2(n17100), .ZN(n19352) );
  NOR3_X1 U12672 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n19359), .ZN(n18781) );
  INV_X1 U12673 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19193) );
  INV_X1 U12674 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19197) );
  NOR2_X1 U12675 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19330) );
  INV_X1 U12676 ( .A(n19332), .ZN(n19340) );
  INV_X1 U12677 ( .A(n17431), .ZN(n19216) );
  AOI21_X1 U12678 ( .B1(n19205), .B2(n19206), .A(n19212), .ZN(n10272) );
  NAND2_X1 U12679 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19361) );
  AND2_X2 U12680 ( .A1(n13317), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20492)
         );
  NAND2_X1 U12682 ( .A1(n10134), .A2(n14683), .ZN(P1_U2810) );
  NAND2_X1 U12683 ( .A1(n10397), .A2(n20333), .ZN(n10134) );
  NAND2_X1 U12684 ( .A1(n10135), .A2(n14951), .ZN(P1_U2842) );
  NAND2_X1 U12685 ( .A1(n10397), .A2(n20392), .ZN(n10135) );
  AOI21_X1 U12686 ( .B1(n11561), .B2(n20391), .A(n11560), .ZN(n11562) );
  NAND2_X1 U12687 ( .A1(n10132), .A2(n10129), .ZN(P1_U2874) );
  NOR2_X1 U12688 ( .A1(n10131), .A2(n10130), .ZN(n10129) );
  NAND2_X1 U12689 ( .A1(n10397), .A2(n10133), .ZN(n10132) );
  INV_X1 U12690 ( .A(n14977), .ZN(n10130) );
  AOI21_X1 U12691 ( .B1(n10397), .B2(n16931), .A(n13263), .ZN(n10396) );
  AOI21_X1 U12692 ( .B1(n15054), .B2(n16931), .A(n15053), .ZN(n15055) );
  NAND2_X1 U12693 ( .A1(n9855), .A2(n9853), .ZN(P1_U2975) );
  INV_X1 U12694 ( .A(n9854), .ZN(n9853) );
  NAND2_X1 U12695 ( .A1(n15335), .A2(n16926), .ZN(n9855) );
  OAI21_X1 U12696 ( .B1(n15097), .B2(n20491), .A(n15096), .ZN(n9854) );
  NAND2_X1 U12697 ( .A1(n15288), .A2(n10045), .ZN(n9876) );
  OAI21_X1 U12698 ( .B1(n15315), .B2(n20481), .A(n10286), .ZN(P1_U3004) );
  AOI21_X1 U12699 ( .B1(n15318), .B2(n15317), .A(n15316), .ZN(n10286) );
  OAI21_X1 U12700 ( .B1(n14364), .B2(n15975), .A(n10372), .ZN(P2_U2824) );
  AOI21_X1 U12701 ( .B1(n10375), .B2(n13130), .A(n10373), .ZN(n10372) );
  NAND2_X1 U12702 ( .A1(n14363), .A2(n10374), .ZN(n10373) );
  INV_X1 U12703 ( .A(n14369), .ZN(n10375) );
  AOI211_X1 U12704 ( .C1(n19406), .C2(n13060), .A(n13059), .B(n13058), .ZN(
        n13133) );
  NAND2_X1 U12705 ( .A1(n14630), .A2(n13130), .ZN(n13131) );
  NOR2_X1 U12706 ( .A1(n10020), .A2(n15955), .ZN(n15946) );
  OAI21_X1 U12707 ( .B1(n16058), .B2(P2_EBX_REG_2__SCAN_IN), .A(n10021), .ZN(
        n13635) );
  NAND2_X1 U12708 ( .A1(n16058), .A2(n10020), .ZN(n10021) );
  INV_X1 U12709 ( .A(n9842), .ZN(n13527) );
  AOI21_X1 U12710 ( .B1(n9598), .B2(n12370), .A(n9843), .ZN(n9842) );
  AOI21_X1 U12711 ( .B1(n14630), .B2(n19433), .A(n14629), .ZN(n14631) );
  OR2_X1 U12712 ( .A1(n14628), .A2(n14627), .ZN(n14629) );
  INV_X1 U12713 ( .A(n10110), .ZN(n10109) );
  OAI21_X1 U12714 ( .B1(n16068), .B2(n16165), .A(n16067), .ZN(n10110) );
  INV_X1 U12715 ( .A(n14347), .ZN(n10195) );
  OAI21_X1 U12716 ( .B1(n14357), .B2(n16409), .A(n14346), .ZN(n14347) );
  NAND2_X1 U12717 ( .A1(n9681), .A2(n10213), .ZN(n10212) );
  INV_X1 U12718 ( .A(n16200), .ZN(n10213) );
  NOR2_X1 U12719 ( .A1(n16209), .A2(n16208), .ZN(n10392) );
  NAND2_X1 U12720 ( .A1(n16464), .A2(n16426), .ZN(n10393) );
  INV_X1 U12721 ( .A(n10029), .ZN(n16282) );
  OAI21_X1 U12722 ( .B1(n16552), .B2(n16429), .A(n10030), .ZN(n10029) );
  AOI21_X1 U12723 ( .B1(n16281), .B2(n10023), .A(n16280), .ZN(n10030) );
  INV_X1 U12724 ( .A(n9830), .ZN(n16293) );
  OAI21_X1 U12725 ( .B1(n16563), .B2(n16429), .A(n9831), .ZN(n9830) );
  AOI21_X1 U12726 ( .B1(n16292), .B2(n10023), .A(n16291), .ZN(n9831) );
  NAND2_X1 U12727 ( .A1(n10023), .A2(n11868), .ZN(n10022) );
  NAND2_X1 U12728 ( .A1(n10023), .A2(n9835), .ZN(n9841) );
  AND2_X1 U12729 ( .A1(n12578), .A2(n12577), .ZN(n12589) );
  NOR2_X1 U12730 ( .A1(n12366), .A2(n12365), .ZN(n12556) );
  NAND2_X1 U12731 ( .A1(n13011), .A2(n13010), .ZN(n13012) );
  OAI211_X1 U12732 ( .C1(n12751), .C2(n13015), .A(n10549), .B(n9890), .ZN(
        P2_U3019) );
  NAND2_X1 U12733 ( .A1(n12740), .A2(n12739), .ZN(n12751) );
  INV_X1 U12734 ( .A(n10056), .ZN(n13015) );
  NAND2_X1 U12735 ( .A1(n16464), .A2(n16689), .ZN(n9887) );
  NAND2_X1 U12736 ( .A1(n9834), .A2(n12739), .ZN(n16527) );
  INV_X1 U12737 ( .A(n10235), .ZN(n16555) );
  OAI21_X1 U12738 ( .B1(n16552), .B2(n16706), .A(n10236), .ZN(n10235) );
  NOR2_X1 U12739 ( .A1(n16553), .A2(n9680), .ZN(n10236) );
  OAI21_X1 U12740 ( .B1(n16566), .B2(n16721), .A(n10077), .ZN(P2_U3028) );
  NOR2_X1 U12741 ( .A1(n16564), .A2(n10079), .ZN(n10078) );
  OAI21_X1 U12742 ( .B1(n16568), .B2(n16721), .A(n9969), .ZN(n9882) );
  NOR2_X1 U12743 ( .A1(n16809), .A2(n10075), .ZN(n16811) );
  NAND2_X1 U12744 ( .A1(n10064), .A2(n10076), .ZN(n10075) );
  AOI21_X1 U12745 ( .B1(n17127), .B2(n17126), .A(n17125), .ZN(n17131) );
  NAND2_X1 U12746 ( .A1(n17574), .A2(P3_EBX_REG_21__SCAN_IN), .ZN(n17560) );
  NAND2_X1 U12747 ( .A1(n17753), .A2(n9652), .ZN(n17730) );
  INV_X1 U12748 ( .A(n17779), .ZN(n17780) );
  AOI21_X1 U12749 ( .B1(n13289), .B2(n13288), .A(n13287), .ZN(n13290) );
  OR2_X1 U12750 ( .A1(n13286), .A2(n13285), .ZN(n13287) );
  OR2_X1 U12751 ( .A1(n12926), .A2(n12925), .ZN(P3_U2802) );
  OR2_X1 U12752 ( .A1(n12924), .A2(n12923), .ZN(n12925) );
  NAND2_X1 U12753 ( .A1(n10290), .A2(n10287), .ZN(P3_U2803) );
  NAND2_X1 U12754 ( .A1(n18048), .A2(n18047), .ZN(n10290) );
  AOI21_X1 U12755 ( .B1(n18052), .B2(n18293), .A(n10288), .ZN(n10287) );
  NAND2_X1 U12756 ( .A1(n18051), .A2(n10289), .ZN(n10288) );
  OAI21_X1 U12757 ( .B1(n10343), .B2(n9787), .A(n10340), .ZN(P3_U2841) );
  NOR2_X1 U12758 ( .A1(n18471), .A2(n10344), .ZN(n10343) );
  INV_X1 U12759 ( .A(n10341), .ZN(n10340) );
  NOR2_X2 U12760 ( .A1(n12618), .A2(n19179), .ZN(n12786) );
  INV_X1 U12761 ( .A(n12835), .ZN(n12813) );
  AND2_X1 U12762 ( .A1(n9626), .A2(n16238), .ZN(n9615) );
  AND2_X1 U12763 ( .A1(n18261), .A2(n10179), .ZN(n9616) );
  INV_X1 U12764 ( .A(n17922), .ZN(n12850) );
  NAND2_X1 U12765 ( .A1(n10410), .A2(n10409), .ZN(n14160) );
  INV_X1 U12766 ( .A(n10574), .ZN(n9980) );
  AND3_X1 U12767 ( .A1(n9655), .A2(P3_EAX_REG_0__SCAN_IN), .A3(n9782), .ZN(
        n9617) );
  AND4_X1 U12768 ( .A1(n10332), .A2(P3_EBX_REG_13__SCAN_IN), .A3(
        P3_EBX_REG_17__SCAN_IN), .A4(P3_EBX_REG_16__SCAN_IN), .ZN(n9618) );
  NAND2_X1 U12769 ( .A1(n10390), .A2(n9698), .ZN(n15115) );
  INV_X1 U12770 ( .A(n17826), .ZN(n12696) );
  NAND2_X1 U12771 ( .A1(n9963), .A2(n9964), .ZN(n14334) );
  NOR2_X1 U12772 ( .A1(n13518), .A2(n11856), .ZN(n9620) );
  NAND2_X1 U12773 ( .A1(n10253), .A2(n10510), .ZN(n16231) );
  AND3_X1 U12774 ( .A1(n11999), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n12412), .ZN(n9622) );
  INV_X1 U12775 ( .A(n19598), .ZN(n10027) );
  NAND2_X1 U12776 ( .A1(n19409), .A2(n13104), .ZN(n15690) );
  AND2_X1 U12777 ( .A1(n9964), .A2(n9750), .ZN(n9623) );
  NAND2_X1 U12778 ( .A1(n10148), .A2(n10566), .ZN(n14809) );
  NAND2_X1 U12779 ( .A1(n15671), .A2(n15672), .ZN(n15652) );
  AND2_X1 U12780 ( .A1(n12246), .A2(n12245), .ZN(n14085) );
  NAND2_X1 U12781 ( .A1(n10102), .A2(n10101), .ZN(n15981) );
  INV_X1 U12782 ( .A(n17926), .ZN(n9983) );
  AND2_X1 U12783 ( .A1(n10399), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9624) );
  AND2_X1 U12784 ( .A1(n12447), .A2(n12441), .ZN(n9625) );
  AND2_X1 U12785 ( .A1(n12500), .A2(n9688), .ZN(n9626) );
  AND2_X1 U12786 ( .A1(n11505), .A2(n10480), .ZN(n9627) );
  AND2_X4 U12787 ( .A1(n10400), .A2(n12709), .ZN(n9628) );
  AND2_X1 U12788 ( .A1(n10311), .A2(n10310), .ZN(n9629) );
  AND2_X1 U12789 ( .A1(n12257), .A2(n10408), .ZN(n9630) );
  AND4_X1 U12790 ( .A1(n11940), .A2(n11939), .A3(n11938), .A4(n11937), .ZN(
        n9631) );
  INV_X1 U12791 ( .A(n16033), .ZN(n10121) );
  AND2_X1 U12792 ( .A1(n9630), .A2(n14332), .ZN(n9632) );
  OR2_X1 U12793 ( .A1(n15642), .A2(n12539), .ZN(n16210) );
  NAND2_X1 U12794 ( .A1(n13722), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10937) );
  AND2_X1 U12795 ( .A1(n9625), .A2(n9745), .ZN(n9633) );
  NAND2_X1 U12796 ( .A1(n12176), .A2(n12175), .ZN(n15687) );
  AND2_X1 U12797 ( .A1(n10485), .A2(n10484), .ZN(n9634) );
  OR2_X1 U12798 ( .A1(n13852), .A2(n13997), .ZN(n9635) );
  AND2_X1 U12799 ( .A1(n11801), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n9636) );
  INV_X1 U12800 ( .A(n16342), .ZN(n10165) );
  AND2_X1 U12801 ( .A1(n15236), .A2(n13240), .ZN(n9637) );
  AND2_X1 U12802 ( .A1(n12418), .A2(n12419), .ZN(n9638) );
  AND2_X1 U12803 ( .A1(n9963), .A2(n9623), .ZN(n9639) );
  AND2_X1 U12804 ( .A1(n9677), .A2(n13828), .ZN(n9640) );
  AND2_X1 U12805 ( .A1(n10297), .A2(n9744), .ZN(n9641) );
  AND2_X1 U12806 ( .A1(n11875), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n9642) );
  AND2_X1 U12807 ( .A1(n9629), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9643) );
  AND2_X1 U12808 ( .A1(n10166), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9644) );
  NOR2_X1 U12809 ( .A1(n16351), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9645) );
  INV_X1 U12810 ( .A(n19177), .ZN(n10298) );
  NAND2_X1 U12811 ( .A1(n10073), .A2(n10064), .ZN(n16429) );
  NOR2_X1 U12812 ( .A1(n16955), .A2(n9781), .ZN(n9646) );
  OR2_X1 U12813 ( .A1(n12330), .A2(n11781), .ZN(n9647) );
  INV_X1 U12814 ( .A(n15977), .ZN(n10433) );
  NOR3_X1 U12815 ( .A1(n13933), .A2(n14085), .A3(n14095), .ZN(n14094) );
  AND2_X1 U12816 ( .A1(n13820), .A2(n13824), .ZN(n9648) );
  AND2_X1 U12817 ( .A1(n9648), .A2(n9747), .ZN(n9649) );
  NAND2_X1 U12818 ( .A1(n18054), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12595) );
  OR2_X1 U12819 ( .A1(n18228), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9650) );
  AND2_X1 U12820 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9651) );
  AND2_X1 U12821 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .ZN(n9652) );
  AND2_X1 U12822 ( .A1(n9652), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n9653) );
  AND2_X1 U12823 ( .A1(n9653), .A2(P3_EBX_REG_9__SCAN_IN), .ZN(n9654) );
  AND4_X1 U12824 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n9655) );
  AND2_X1 U12825 ( .A1(n10331), .A2(P3_EBX_REG_23__SCAN_IN), .ZN(n9656) );
  AND2_X1 U12826 ( .A1(n9618), .A2(P3_EBX_REG_18__SCAN_IN), .ZN(n9657) );
  AND2_X1 U12827 ( .A1(n10188), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n9658) );
  NAND2_X1 U12828 ( .A1(n10879), .A2(n20541), .ZN(n13484) );
  INV_X1 U12829 ( .A(n12802), .ZN(n12784) );
  INV_X1 U12830 ( .A(n12784), .ZN(n16791) );
  NAND2_X1 U12831 ( .A1(n15542), .A2(n10866), .ZN(n13452) );
  INV_X1 U12832 ( .A(n10295), .ZN(n18294) );
  NAND2_X1 U12833 ( .A1(n18375), .A2(n17902), .ZN(n10295) );
  AOI21_X2 U12834 ( .B1(n12962), .B2(n12961), .A(n19212), .ZN(n12963) );
  AND4_X1 U12835 ( .A1(n10777), .A2(n10776), .A3(n10775), .A4(n10774), .ZN(
        n9659) );
  NOR2_X1 U12836 ( .A1(n14229), .A2(n19179), .ZN(n12785) );
  INV_X1 U12837 ( .A(n12785), .ZN(n12822) );
  AND2_X1 U12838 ( .A1(n16900), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n9660) );
  XNOR2_X1 U12839 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12587), .ZN(
        n9661) );
  OR2_X1 U12840 ( .A1(n12407), .A2(n10452), .ZN(n12414) );
  OR2_X1 U12841 ( .A1(n18133), .A2(n10283), .ZN(n18070) );
  NAND2_X1 U12842 ( .A1(n13821), .A2(n9648), .ZN(n14190) );
  INV_X1 U12843 ( .A(n10254), .ZN(n16219) );
  NAND2_X1 U12844 ( .A1(n12258), .A2(n9632), .ZN(n14331) );
  AND2_X1 U12845 ( .A1(n14607), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11942) );
  NAND2_X1 U12846 ( .A1(n18292), .A2(n18261), .ZN(n18195) );
  INV_X1 U12847 ( .A(n10823), .ZN(n10838) );
  AND2_X1 U12848 ( .A1(n11863), .A2(n9620), .ZN(n9662) );
  NAND2_X1 U12849 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12855), .ZN(
        n9663) );
  NAND2_X1 U12850 ( .A1(n9952), .A2(n10053), .ZN(n12741) );
  NAND2_X1 U12851 ( .A1(n12517), .A2(n10454), .ZN(n9664) );
  OR2_X1 U12852 ( .A1(n9635), .A2(n10488), .ZN(n9665) );
  AND2_X1 U12853 ( .A1(n10424), .A2(n10105), .ZN(n9666) );
  INV_X1 U12854 ( .A(n9809), .ZN(n18133) );
  OR2_X1 U12855 ( .A1(n18167), .A2(n10304), .ZN(n9809) );
  INV_X1 U12856 ( .A(n10512), .ZN(n16202) );
  INV_X1 U12857 ( .A(n11687), .ZN(n10067) );
  AND2_X1 U12858 ( .A1(n13088), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13092) );
  NOR2_X1 U12859 ( .A1(n13777), .A2(n9665), .ZN(n14036) );
  NOR2_X1 U12860 ( .A1(n14827), .A2(n10149), .ZN(n14794) );
  NOR2_X1 U12861 ( .A1(n14109), .A2(n10496), .ZN(n14840) );
  NAND2_X1 U12862 ( .A1(n14904), .A2(n11192), .ZN(n14854) );
  AND4_X1 U12863 ( .A1(n12809), .A2(n12808), .A3(n12807), .A4(n12806), .ZN(
        n9667) );
  AND2_X1 U12864 ( .A1(n10355), .A2(n10045), .ZN(n9668) );
  NAND2_X1 U12865 ( .A1(n13077), .A2(n10377), .ZN(n13081) );
  INV_X2 U12866 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11839) );
  NAND2_X1 U12867 ( .A1(n13077), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13079) );
  AND2_X1 U12868 ( .A1(n9900), .A2(n9899), .ZN(n9669) );
  AND2_X1 U12869 ( .A1(n9918), .A2(n9917), .ZN(n9670) );
  AND4_X1 U12870 ( .A1(n10782), .A2(n10781), .A3(n10780), .A4(n10779), .ZN(
        n9671) );
  AND4_X1 U12871 ( .A1(n11914), .A2(n11916), .A3(n11917), .A4(n11915), .ZN(
        n9672) );
  AND2_X1 U12872 ( .A1(n12258), .A2(n9630), .ZN(n9673) );
  XOR2_X1 U12873 ( .A(n12342), .B(n11926), .Z(n9674) );
  AND2_X1 U12874 ( .A1(n10421), .A2(n10420), .ZN(n9675) );
  NAND2_X1 U12875 ( .A1(n10333), .A2(n12410), .ZN(n16438) );
  AND2_X1 U12876 ( .A1(n13074), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13077) );
  AND2_X1 U12877 ( .A1(n13092), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13094) );
  INV_X1 U12878 ( .A(n12742), .ZN(n10445) );
  AND2_X1 U12879 ( .A1(n12228), .A2(n10413), .ZN(n9677) );
  NOR2_X1 U12880 ( .A1(n15687), .A2(n16112), .ZN(n15671) );
  NOR2_X1 U12881 ( .A1(n18133), .A2(n18120), .ZN(n18121) );
  INV_X1 U12882 ( .A(n12406), .ZN(n10452) );
  AND3_X1 U12883 ( .A1(n11871), .A2(n11880), .A3(
        P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n9678) );
  NAND2_X1 U12884 ( .A1(n12482), .A2(n9633), .ZN(n9679) );
  AND2_X1 U12885 ( .A1(n16554), .A2(n16724), .ZN(n9680) );
  NOR2_X1 U12886 ( .A1(n13089), .A2(n16332), .ZN(n13088) );
  OR2_X1 U12887 ( .A1(n16450), .A2(n16409), .ZN(n9681) );
  NAND2_X1 U12888 ( .A1(n10309), .A2(n10311), .ZN(n12607) );
  AND4_X1 U12889 ( .A1(n12643), .A2(n12642), .A3(n12641), .A4(n12640), .ZN(
        n9682) );
  INV_X1 U12890 ( .A(n16908), .ZN(n20333) );
  INV_X1 U12891 ( .A(n20252), .ZN(n19657) );
  AND2_X1 U12892 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13063) );
  AND4_X1 U12893 ( .A1(n11936), .A2(n11935), .A3(n11934), .A4(n11933), .ZN(
        n9683) );
  AND2_X1 U12894 ( .A1(n12517), .A2(n12516), .ZN(n9684) );
  AND2_X1 U12895 ( .A1(n10174), .A2(n10175), .ZN(n18060) );
  OR2_X1 U12896 ( .A1(n16580), .A2(n21336), .ZN(n9685) );
  OR2_X1 U12897 ( .A1(n18682), .A2(n12851), .ZN(n9686) );
  INV_X1 U12898 ( .A(n15146), .ZN(n10391) );
  AND2_X1 U12899 ( .A1(n15236), .A2(n15444), .ZN(n9687) );
  OR2_X1 U12900 ( .A1(n9645), .A2(n16362), .ZN(n9688) );
  AND3_X1 U12901 ( .A1(n11647), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11646), .ZN(n9689) );
  AND2_X1 U12902 ( .A1(n12029), .A2(n12034), .ZN(n9690) );
  INV_X1 U12903 ( .A(n14827), .ZN(n10148) );
  AND2_X1 U12904 ( .A1(n12318), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9691) );
  INV_X1 U12905 ( .A(n19522), .ZN(n19597) );
  NAND2_X1 U12906 ( .A1(n13624), .A2(n13500), .ZN(n19522) );
  AND2_X1 U12907 ( .A1(n13763), .A2(n9649), .ZN(n9692) );
  AND2_X1 U12908 ( .A1(n9912), .A2(n9911), .ZN(n12427) );
  INV_X1 U12909 ( .A(n12890), .ZN(n18204) );
  AND2_X1 U12910 ( .A1(n9925), .A2(n13238), .ZN(n9693) );
  OR2_X1 U12911 ( .A1(n15236), .A2(n13245), .ZN(n9694) );
  AND2_X1 U12912 ( .A1(n10424), .A2(n10095), .ZN(n9695) );
  NAND2_X1 U12913 ( .A1(n12482), .A2(n9625), .ZN(n12468) );
  AND2_X1 U12914 ( .A1(n10536), .A2(n16275), .ZN(n9696) );
  AND2_X1 U12915 ( .A1(n10256), .A2(n16374), .ZN(n9697) );
  AND2_X1 U12916 ( .A1(n10389), .A2(n15146), .ZN(n9698) );
  AND2_X1 U12917 ( .A1(n10248), .A2(n10388), .ZN(n9699) );
  AND2_X1 U12918 ( .A1(n10260), .A2(n14330), .ZN(n9700) );
  INV_X1 U12919 ( .A(n14787), .ZN(n11299) );
  AND2_X1 U12920 ( .A1(n10224), .A2(n12449), .ZN(n9701) );
  AND2_X1 U12921 ( .A1(n9627), .A2(n10481), .ZN(n9702) );
  AND2_X1 U12922 ( .A1(n9668), .A2(n15216), .ZN(n9703) );
  AND2_X1 U12923 ( .A1(n9879), .A2(n11433), .ZN(n9704) );
  AND3_X1 U12924 ( .A1(n16263), .A2(n16283), .A3(n16251), .ZN(n9705) );
  AND2_X1 U12925 ( .A1(n10058), .A2(n16922), .ZN(n9706) );
  NAND2_X1 U12926 ( .A1(n13068), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13071) );
  NAND2_X1 U12927 ( .A1(n10121), .A2(n14431), .ZN(n16027) );
  AND2_X1 U12928 ( .A1(n10443), .A2(n12580), .ZN(n9707) );
  OR2_X1 U12929 ( .A1(n13104), .A2(n10370), .ZN(n9708) );
  NOR2_X1 U12930 ( .A1(n19351), .A2(n10275), .ZN(n9709) );
  AND2_X1 U12931 ( .A1(n11509), .A2(n11508), .ZN(n14891) );
  NAND2_X1 U12932 ( .A1(n14107), .A2(n11108), .ZN(n14109) );
  AND2_X1 U12933 ( .A1(n15099), .A2(n15216), .ZN(n9710) );
  OR2_X1 U12934 ( .A1(n16259), .A2(n16258), .ZN(n9711) );
  INV_X1 U12935 ( .A(n10012), .ZN(n12323) );
  NAND2_X1 U12936 ( .A1(n11803), .A2(n12331), .ZN(n10012) );
  INV_X1 U12937 ( .A(n10547), .ZN(n10546) );
  OR2_X1 U12938 ( .A1(n17736), .A2(n17763), .ZN(n9712) );
  NOR2_X1 U12939 ( .A1(n17973), .A2(n19360), .ZN(n9713) );
  NAND2_X1 U12940 ( .A1(n17811), .A2(n10188), .ZN(n10189) );
  AND2_X1 U12941 ( .A1(n9973), .A2(n9971), .ZN(n13037) );
  AND2_X1 U12942 ( .A1(n9638), .A2(n12406), .ZN(n9714) );
  NAND2_X1 U12943 ( .A1(n10981), .A2(n10919), .ZN(n9715) );
  INV_X1 U12944 ( .A(n11908), .ZN(n11956) );
  OAI21_X1 U12945 ( .B1(n18178), .B2(n18080), .A(n12869), .ZN(n10089) );
  AND2_X1 U12946 ( .A1(n16438), .A2(n10564), .ZN(n9716) );
  OAI211_X1 U12947 ( .C1(n12315), .C2(n14059), .A(n10205), .B(n10204), .ZN(
        n11854) );
  NAND2_X1 U12948 ( .A1(n12482), .A2(n12441), .ZN(n12445) );
  AND2_X1 U12949 ( .A1(n10968), .A2(n10036), .ZN(n9717) );
  AND2_X1 U12950 ( .A1(n10968), .A2(n10037), .ZN(n9718) );
  AND3_X1 U12951 ( .A1(n12820), .A2(n12815), .A3(n10087), .ZN(n9719) );
  AND3_X1 U12952 ( .A1(n16250), .A2(n12481), .A3(n10335), .ZN(n9720) );
  OR3_X1 U12953 ( .A1(n12737), .A2(n12736), .A3(n12735), .ZN(P3_U2640) );
  AND3_X1 U12954 ( .A1(n12819), .A2(n12817), .A3(n9719), .ZN(n9722) );
  AND2_X1 U12955 ( .A1(n10156), .A2(n10155), .ZN(n9723) );
  AND2_X1 U12956 ( .A1(n15597), .A2(n15596), .ZN(n12994) );
  OR2_X1 U12957 ( .A1(n17926), .A2(n19320), .ZN(n9724) );
  INV_X1 U12958 ( .A(n13190), .ZN(n9939) );
  AND2_X1 U12959 ( .A1(n9668), .A2(n15303), .ZN(n9725) );
  AND2_X1 U12960 ( .A1(n10503), .A2(n14744), .ZN(n9726) );
  INV_X1 U12961 ( .A(n16899), .ZN(n16900) );
  AND2_X1 U12962 ( .A1(n10478), .A2(n14135), .ZN(n9727) );
  NOR2_X1 U12963 ( .A1(n12692), .A2(n10291), .ZN(n9728) );
  NOR2_X1 U12964 ( .A1(n15629), .A2(n10449), .ZN(n9729) );
  INV_X1 U12965 ( .A(n18379), .ZN(n16901) );
  NAND2_X1 U12966 ( .A1(n12849), .A2(n12848), .ZN(n18379) );
  INV_X1 U12967 ( .A(n10528), .ZN(n10527) );
  NOR2_X1 U12968 ( .A1(n10530), .A2(n14329), .ZN(n10528) );
  AND2_X1 U12969 ( .A1(n10830), .A2(n10837), .ZN(n9730) );
  AND2_X1 U12970 ( .A1(n11803), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9731) );
  AND2_X1 U12971 ( .A1(n9620), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n9732) );
  NAND2_X1 U12972 ( .A1(n13766), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n9733) );
  NAND2_X1 U12973 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12861), .ZN(
        n9734) );
  AND2_X1 U12974 ( .A1(n12406), .A2(n12415), .ZN(n9735) );
  INV_X1 U12975 ( .A(n10582), .ZN(n10154) );
  INV_X1 U12976 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15829) );
  INV_X1 U12977 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10225) );
  INV_X2 U12978 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n10144) );
  OR3_X1 U12979 ( .A1(n13120), .A2(n10368), .A3(n10369), .ZN(n9736) );
  NAND2_X1 U12980 ( .A1(n14939), .A2(n11505), .ZN(n14888) );
  NAND2_X1 U12981 ( .A1(n10116), .A2(n10114), .ZN(n14380) );
  NAND2_X1 U12982 ( .A1(n13821), .A2(n13820), .ZN(n13822) );
  NAND2_X1 U12984 ( .A1(n13884), .A2(n12323), .ZN(n12315) );
  AND2_X1 U12985 ( .A1(n14799), .A2(n9634), .ZN(n9737) );
  NAND2_X1 U12986 ( .A1(n15690), .A2(n16257), .ZN(n15691) );
  INV_X1 U12987 ( .A(n20391), .ZN(n14972) );
  AND2_X1 U12988 ( .A1(n20396), .A2(n14974), .ZN(n20391) );
  OR2_X1 U12989 ( .A1(n13933), .A2(n14085), .ZN(n9738) );
  AND2_X1 U12990 ( .A1(n16802), .A2(n9618), .ZN(n9739) );
  NOR2_X2 U12991 ( .A1(n12626), .A2(n12625), .ZN(n19360) );
  INV_X1 U12992 ( .A(n19360), .ZN(n17972) );
  NOR2_X1 U12993 ( .A1(n16056), .A2(n10440), .ZN(n16043) );
  NOR2_X1 U12994 ( .A1(n13098), .A2(n15725), .ZN(n13100) );
  OR2_X1 U12995 ( .A1(n13777), .A2(n9962), .ZN(n15686) );
  OR2_X1 U12996 ( .A1(n16056), .A2(n10442), .ZN(n16048) );
  INV_X1 U12997 ( .A(n16351), .ZN(n10532) );
  INV_X1 U12998 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n14059) );
  NAND2_X1 U12999 ( .A1(n13092), .A2(n9651), .ZN(n13096) );
  AND2_X1 U13000 ( .A1(n20524), .A2(n20508), .ZN(n13222) );
  AND2_X1 U13001 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n9740) );
  AND2_X1 U13002 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n9741) );
  AND2_X1 U13003 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n9742) );
  AND2_X1 U13004 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n9743) );
  AND3_X1 U13005 ( .A1(n12875), .A2(n12881), .A3(n12874), .ZN(n9744) );
  XNOR2_X1 U13006 ( .A(n13195), .B(n13649), .ZN(n13726) );
  OR2_X1 U13007 ( .A1(n12532), .A2(n12448), .ZN(n9745) );
  NAND2_X1 U13008 ( .A1(n12050), .A2(n12049), .ZN(n13528) );
  NOR3_X1 U13009 ( .A1(n13120), .A2(n10369), .A3(n13022), .ZN(n13121) );
  NAND2_X1 U13010 ( .A1(n14074), .A2(n12044), .ZN(n13540) );
  AND2_X1 U13011 ( .A1(n13100), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13102) );
  AND2_X1 U13012 ( .A1(n12229), .A2(n9677), .ZN(n13827) );
  NAND2_X1 U13013 ( .A1(n18507), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12968) );
  INV_X1 U13014 ( .A(n12968), .ZN(n10179) );
  AND2_X1 U13015 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n9746) );
  NAND2_X1 U13016 ( .A1(n13528), .A2(n10487), .ZN(n13636) );
  NAND2_X1 U13017 ( .A1(n13528), .A2(n9966), .ZN(n13675) );
  NAND2_X1 U13018 ( .A1(n13661), .A2(n9690), .ZN(n13971) );
  AND4_X1 U13019 ( .A1(n14189), .A2(n14188), .A3(n14187), .A4(n14186), .ZN(
        n9747) );
  NOR2_X1 U13020 ( .A1(n13777), .A2(n9635), .ZN(n13996) );
  AND4_X1 U13021 ( .A1(n12213), .A2(n12221), .A3(n12212), .A4(n10417), .ZN(
        n9748) );
  AND2_X1 U13022 ( .A1(n18054), .A2(n10324), .ZN(n12591) );
  NAND2_X1 U13023 ( .A1(n12242), .A2(n12241), .ZN(n13933) );
  INV_X1 U13024 ( .A(n13891), .ZN(n9840) );
  OR2_X1 U13025 ( .A1(n16220), .A2(n16484), .ZN(n9749) );
  NAND2_X1 U13026 ( .A1(n19167), .A2(n12880), .ZN(n18703) );
  NOR2_X1 U13027 ( .A1(n12171), .A2(n15728), .ZN(n9750) );
  AND2_X1 U13028 ( .A1(n13926), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n9751) );
  AND2_X1 U13029 ( .A1(n20503), .A2(n10862), .ZN(n9752) );
  AND2_X1 U13030 ( .A1(n17574), .A2(n10331), .ZN(n9753) );
  CLKBUF_X3 U13031 ( .A(n12008), .Z(n12532) );
  OR2_X1 U13032 ( .A1(n10572), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9754) );
  NOR2_X1 U13033 ( .A1(n14733), .A2(n14735), .ZN(n11543) );
  BUF_X1 U13034 ( .A(n10813), .Z(n20508) );
  NOR2_X1 U13035 ( .A1(n18228), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9755) );
  AND2_X1 U13036 ( .A1(n17176), .A2(n12611), .ZN(n9756) );
  INV_X1 U13037 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15736) );
  INV_X1 U13038 ( .A(n14095), .ZN(n10412) );
  AND2_X1 U13039 ( .A1(n12250), .A2(n12249), .ZN(n14095) );
  INV_X1 U13040 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17477) );
  OR2_X1 U13041 ( .A1(n13676), .A2(n13681), .ZN(n9757) );
  NAND2_X1 U13042 ( .A1(n12269), .A2(n12268), .ZN(n9758) );
  INV_X1 U13043 ( .A(n14559), .ZN(n10103) );
  INV_X1 U13044 ( .A(n10877), .ZN(n13176) );
  OR2_X1 U13045 ( .A1(n10876), .A2(n10875), .ZN(n10877) );
  NOR2_X1 U13046 ( .A1(n18325), .A2(n12859), .ZN(n9759) );
  AND2_X1 U13047 ( .A1(n10476), .A2(n10475), .ZN(n9760) );
  AND2_X1 U13048 ( .A1(n9977), .A2(n18047), .ZN(n9761) );
  AND2_X1 U13049 ( .A1(n10456), .A2(n10455), .ZN(n9762) );
  AND2_X1 U13050 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n9763) );
  AND2_X1 U13051 ( .A1(n9651), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9764) );
  INV_X1 U13052 ( .A(n10015), .ZN(n19860) );
  OR2_X1 U13053 ( .A1(n11622), .A2(n11621), .ZN(n11930) );
  AND2_X1 U13054 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n9765) );
  INV_X1 U13055 ( .A(n10537), .ZN(n10536) );
  NAND2_X1 U13056 ( .A1(n10540), .A2(n16283), .ZN(n10537) );
  INV_X1 U13057 ( .A(n10559), .ZN(n10357) );
  INV_X1 U13058 ( .A(n11380), .ZN(n11371) );
  INV_X1 U13059 ( .A(n11371), .ZN(n13162) );
  NOR2_X1 U13060 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11380) );
  INV_X1 U13061 ( .A(n19406), .ZN(n16838) );
  NAND2_X1 U13062 ( .A1(n18054), .A2(n10323), .ZN(n12592) );
  NOR2_X1 U13063 ( .A1(n10302), .A2(n9644), .ZN(n9981) );
  INV_X1 U13064 ( .A(n13630), .ZN(n9838) );
  NAND2_X1 U13065 ( .A1(n16436), .A2(n16733), .ZN(n16409) );
  INV_X1 U13066 ( .A(n16409), .ZN(n10023) );
  AND2_X1 U13067 ( .A1(n17753), .A2(n9653), .ZN(n9766) );
  NAND3_X1 U13068 ( .A1(n12762), .A2(n12761), .A3(n12760), .ZN(n13029) );
  INV_X1 U13069 ( .A(n13627), .ZN(n11868) );
  AND2_X1 U13070 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n9767) );
  AND2_X1 U13071 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n9768) );
  AND2_X1 U13072 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n9769) );
  AND2_X1 U13073 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n9770) );
  AND2_X1 U13074 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n9771) );
  AND2_X1 U13075 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n9772) );
  INV_X1 U13076 ( .A(n14671), .ZN(n14651) );
  XNOR2_X1 U13077 ( .A(n12857), .B(n12858), .ZN(n18324) );
  AND2_X1 U13078 ( .A1(n10492), .A2(n10491), .ZN(n9773) );
  AND2_X1 U13079 ( .A1(n14536), .A2(n14535), .ZN(n9774) );
  AND2_X1 U13080 ( .A1(n12183), .A2(n9960), .ZN(n9775) );
  NOR2_X1 U13081 ( .A1(n9982), .A2(n9981), .ZN(n9776) );
  INV_X1 U13082 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18647) );
  AND2_X1 U13083 ( .A1(n14447), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n9777) );
  AND2_X1 U13084 ( .A1(n14447), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n9778) );
  AND2_X1 U13085 ( .A1(n14447), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n9779) );
  NOR2_X1 U13086 ( .A1(n12973), .A2(n18098), .ZN(n10284) );
  INV_X1 U13087 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17731) );
  OR2_X1 U13088 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n10304), .ZN(
        n9780) );
  AND2_X1 U13089 ( .A1(n11482), .A2(n10478), .ZN(n9781) );
  INV_X1 U13090 ( .A(n16429), .ZN(n16383) );
  AND3_X1 U13091 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_1__SCAN_IN), .ZN(n9782) );
  AND2_X1 U13092 ( .A1(n12931), .A2(n12928), .ZN(n9783) );
  AND2_X1 U13093 ( .A1(n10255), .A2(n10513), .ZN(n9784) );
  NOR2_X1 U13094 ( .A1(n18217), .A2(n18222), .ZN(n17287) );
  OR2_X1 U13095 ( .A1(n21336), .A2(n16592), .ZN(n9785) );
  AND2_X1 U13096 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n9786) );
  OR2_X1 U13097 ( .A1(n18695), .A2(n18465), .ZN(n9787) );
  OR2_X1 U13099 ( .A1(n18701), .A2(n19289), .ZN(n9788) );
  INV_X1 U13100 ( .A(n20166), .ZN(n15574) );
  AND2_X1 U13101 ( .A1(READY12_REG_SCAN_IN), .A2(READY21_REG_SCAN_IN), .ZN(
        n20166) );
  INV_X1 U13102 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17237) );
  INV_X1 U13103 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10455) );
  INV_X1 U13104 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19189) );
  AND3_X1 U13105 ( .A1(n15327), .A2(n15337), .A3(n15343), .ZN(n9789) );
  AND2_X1 U13106 ( .A1(n15386), .A2(n15371), .ZN(n9790) );
  AND2_X1 U13107 ( .A1(n10309), .A2(n9629), .ZN(n9791) );
  AND2_X1 U13108 ( .A1(n9657), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n9792) );
  NOR2_X1 U13109 ( .A1(n9785), .A2(n16591), .ZN(n9793) );
  INV_X1 U13110 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17618) );
  INV_X1 U13111 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10045) );
  INV_X1 U13112 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n17437) );
  NAND2_X1 U13113 ( .A1(n13163), .A2(n20934), .ZN(n20491) );
  INV_X1 U13114 ( .A(n20491), .ZN(n16931) );
  INV_X1 U13115 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n9996) );
  INV_X1 U13116 ( .A(n15304), .ZN(n10403) );
  INV_X1 U13117 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n10065) );
  INV_X1 U13118 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10313) );
  OR2_X1 U13119 ( .A1(n16471), .A2(n10514), .ZN(n9794) );
  INV_X1 U13120 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10312) );
  OR2_X1 U13121 ( .A1(n9785), .A2(n10364), .ZN(n9795) );
  AND2_X1 U13122 ( .A1(n10053), .A2(n9951), .ZN(n9796) );
  INV_X1 U13123 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10378) );
  AND2_X1 U13124 ( .A1(n9658), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n9797) );
  OAI221_X1 U13125 ( .B1(n20667), .B2(n20782), .C1(n20667), .C2(n20650), .A(
        n20985), .ZN(n20669) );
  AOI22_X2 U13126 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20531), .B1(DATAI_29_), 
        .B2(n20493), .ZN(n21053) );
  AOI22_X2 U13127 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20531), .B1(DATAI_24_), 
        .B2(n20493), .ZN(n21023) );
  NOR2_X2 U13128 ( .A1(n20491), .A2(n20490), .ZN(n20531) );
  NAND2_X1 U13129 ( .A1(n9798), .A2(n11875), .ZN(n10015) );
  NAND2_X1 U13130 ( .A1(n9798), .A2(n9620), .ZN(n11883) );
  NAND2_X1 U13131 ( .A1(n9798), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10249) );
  NAND2_X1 U13132 ( .A1(n9642), .A2(n9798), .ZN(n10016) );
  NAND2_X1 U13133 ( .A1(n9732), .A2(n9798), .ZN(n9828) );
  AND2_X2 U13134 ( .A1(n13873), .A2(n13627), .ZN(n9798) );
  INV_X1 U13135 ( .A(n10356), .ZN(n9800) );
  AOI21_X2 U13136 ( .B1(n9672), .B2(n11919), .A(n10559), .ZN(n9801) );
  NAND2_X2 U13137 ( .A1(n9801), .A2(n9800), .ZN(n10541) );
  NAND2_X1 U13138 ( .A1(n9810), .A2(n10398), .ZN(n18315) );
  INV_X1 U13139 ( .A(n18324), .ZN(n9811) );
  NAND3_X1 U13140 ( .A1(n13208), .A2(n13944), .A3(n9818), .ZN(n9817) );
  NAND2_X1 U13141 ( .A1(n9819), .A2(n20461), .ZN(n9818) );
  INV_X1 U13142 ( .A(n13989), .ZN(n9819) );
  NAND2_X1 U13143 ( .A1(n13748), .A2(n13749), .ZN(n9820) );
  INV_X1 U13144 ( .A(n9821), .ZN(n10285) );
  NAND3_X1 U13145 ( .A1(n10967), .A2(n10968), .A3(n10949), .ZN(n11020) );
  XNOR2_X2 U13146 ( .A(n9823), .B(n10878), .ZN(n10968) );
  NAND2_X1 U13147 ( .A1(n10143), .A2(n10142), .ZN(n9823) );
  AND2_X2 U13148 ( .A1(n9824), .A2(n10168), .ZN(n10967) );
  NAND2_X1 U13149 ( .A1(n13181), .A2(n10974), .ZN(n9824) );
  INV_X1 U13150 ( .A(n9826), .ZN(n9825) );
  NAND2_X1 U13151 ( .A1(n15086), .A2(n10401), .ZN(n14352) );
  XNOR2_X2 U13152 ( .A(n11931), .B(n9850), .ZN(n14147) );
  AND2_X1 U13153 ( .A1(n9829), .A2(n9828), .ZN(n11916) );
  AND2_X2 U13154 ( .A1(n11868), .A2(n13873), .ZN(n11863) );
  CLKBUF_X1 U13155 ( .A(n16714), .Z(n9835) );
  AND2_X2 U13156 ( .A1(n13518), .A2(n16714), .ZN(n11879) );
  NOR2_X2 U13157 ( .A1(n16714), .A2(n9836), .ZN(n11871) );
  NAND3_X1 U13158 ( .A1(n13448), .A2(n13447), .A3(n9841), .ZN(P2_U3013) );
  AND2_X1 U13159 ( .A1(n11903), .A2(n9845), .ZN(n9847) );
  NAND2_X1 U13160 ( .A1(n9683), .A2(n9631), .ZN(n9846) );
  AND4_X2 U13161 ( .A1(n11911), .A2(n11909), .A3(n11912), .A4(n11910), .ZN(
        n11919) );
  NAND2_X2 U13162 ( .A1(n9945), .A2(n9848), .ZN(n14203) );
  NAND2_X1 U13163 ( .A1(n11954), .A2(n14208), .ZN(n10252) );
  INV_X1 U13164 ( .A(n11931), .ZN(n9849) );
  AND2_X1 U13165 ( .A1(n12204), .A2(n9851), .ZN(n12205) );
  NAND2_X1 U13166 ( .A1(n16933), .A2(n16932), .ZN(n9852) );
  XNOR2_X2 U13167 ( .A(n9860), .B(n10858), .ZN(n20607) );
  OAI21_X2 U13168 ( .B1(n13720), .B2(n9859), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10858) );
  NAND2_X1 U13169 ( .A1(n9730), .A2(n10238), .ZN(n13304) );
  OAI21_X2 U13170 ( .B1(n10032), .B2(n10599), .A(n10836), .ZN(n9860) );
  NAND2_X2 U13171 ( .A1(n9861), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10032) );
  NAND3_X1 U13172 ( .A1(n10832), .A2(n10833), .A3(n10834), .ZN(n9861) );
  NAND2_X2 U13173 ( .A1(n13250), .A2(n15236), .ZN(n15086) );
  AND2_X2 U13174 ( .A1(n10508), .A2(n9862), .ZN(n10163) );
  NAND2_X1 U13175 ( .A1(n9863), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9862) );
  NAND2_X1 U13176 ( .A1(n14202), .A2(n12368), .ZN(n16430) );
  NAND2_X1 U13177 ( .A1(n9864), .A2(n11974), .ZN(n10508) );
  NAND2_X1 U13178 ( .A1(n14203), .A2(n11975), .ZN(n9864) );
  AND2_X1 U13179 ( .A1(n16268), .A2(n9865), .ZN(n16544) );
  NAND2_X1 U13180 ( .A1(n16267), .A2(n16519), .ZN(n9865) );
  NAND3_X1 U13181 ( .A1(n9866), .A2(n10385), .A3(n9615), .ZN(n10011) );
  NAND3_X1 U13182 ( .A1(n9866), .A2(n10385), .A3(n9615), .ZN(n9903) );
  NAND3_X1 U13183 ( .A1(n9866), .A2(n10385), .A3(n9626), .ZN(n10200) );
  NAND2_X1 U13184 ( .A1(n9870), .A2(n9867), .ZN(n11418) );
  INV_X1 U13185 ( .A(n11406), .ZN(n9869) );
  NAND2_X1 U13186 ( .A1(n9871), .A2(n11405), .ZN(n9870) );
  NAND2_X1 U13187 ( .A1(n9873), .A2(n9872), .ZN(n9871) );
  NAND2_X1 U13188 ( .A1(n11402), .A2(n11403), .ZN(n9872) );
  INV_X1 U13189 ( .A(n13711), .ZN(n9879) );
  NAND2_X1 U13190 ( .A1(n9881), .A2(n11431), .ZN(n9880) );
  NAND2_X1 U13191 ( .A1(n11421), .A2(n11420), .ZN(n9881) );
  NAND3_X1 U13192 ( .A1(n14328), .A2(n14327), .A3(n10262), .ZN(n10013) );
  NAND2_X2 U13193 ( .A1(n9935), .A2(n13237), .ZN(n15218) );
  NAND2_X1 U13194 ( .A1(n10985), .A2(n9885), .ZN(n9883) );
  NAND2_X1 U13195 ( .A1(n16267), .A2(n9784), .ZN(n10512) );
  OAI21_X1 U13196 ( .B1(n15292), .B2(n20293), .A(n10396), .ZN(P1_U2969) );
  OAI211_X1 U13197 ( .C1(n16466), .C2(n16706), .A(n16465), .B(n9887), .ZN(
        P2_U3020) );
  NAND2_X1 U13198 ( .A1(n10010), .A2(n10009), .ZN(n9888) );
  OR2_X1 U13199 ( .A1(n13025), .A2(n16721), .ZN(n9890) );
  NAND3_X1 U13200 ( .A1(n9894), .A2(n9893), .A3(n9892), .ZN(n9891) );
  NAND3_X1 U13201 ( .A1(n9898), .A2(n9897), .A3(n9896), .ZN(n9895) );
  NAND3_X1 U13202 ( .A1(n9902), .A2(n9901), .A3(n9697), .ZN(n9900) );
  NAND2_X1 U13203 ( .A1(n12411), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16370) );
  NAND3_X1 U13204 ( .A1(n11973), .A2(n10257), .A3(n12367), .ZN(n9902) );
  OR2_X1 U13205 ( .A1(n10158), .A2(n9905), .ZN(n9904) );
  XNOR2_X2 U13206 ( .A(n12411), .B(n11977), .ZN(n10157) );
  OAI21_X1 U13207 ( .B1(n11901), .B2(n11800), .A(n11688), .ZN(n12372) );
  NAND2_X1 U13208 ( .A1(n12543), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n9908) );
  OR2_X2 U13209 ( .A1(n11900), .A2(n11899), .ZN(n12371) );
  AND2_X1 U13210 ( .A1(n14443), .A2(n10046), .ZN(n14475) );
  NOR2_X1 U13211 ( .A1(n12407), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n9911) );
  NAND2_X1 U13212 ( .A1(n13168), .A2(n13169), .ZN(n9913) );
  NAND2_X1 U13213 ( .A1(n9913), .A2(n13174), .ZN(n13989) );
  OAI21_X2 U13214 ( .B1(n15560), .B2(n13645), .A(n13205), .ZN(n13987) );
  NAND3_X1 U13215 ( .A1(n13987), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n9917) );
  NAND2_X1 U13216 ( .A1(n13989), .A2(n9919), .ZN(n9918) );
  XNOR2_X1 U13217 ( .A(n9935), .B(n15237), .ZN(n15516) );
  XNOR2_X1 U13218 ( .A(n9936), .B(n10895), .ZN(n10985) );
  OAI21_X2 U13219 ( .B1(n10032), .B2(n16848), .A(n10841), .ZN(n9936) );
  NAND2_X1 U13220 ( .A1(n9945), .A2(n11932), .ZN(n14199) );
  NAND2_X1 U13221 ( .A1(n10163), .A2(n9946), .ZN(n16400) );
  NAND3_X1 U13222 ( .A1(n11871), .A2(n11863), .A3(
        P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n9953) );
  OAI21_X1 U13223 ( .B1(n11904), .B2(n21270), .A(n9953), .ZN(n11858) );
  OR2_X1 U13224 ( .A1(n16563), .A2(n16706), .ZN(n10080) );
  NOR2_X4 U13225 ( .A1(n15632), .A2(n15633), .ZN(n15631) );
  NAND2_X1 U13226 ( .A1(n10362), .A2(n9968), .ZN(n16381) );
  NAND3_X1 U13227 ( .A1(n10361), .A2(n10163), .A3(n10162), .ZN(n9968) );
  NAND2_X1 U13228 ( .A1(n16310), .A2(n12739), .ZN(n9970) );
  NAND3_X1 U13229 ( .A1(n9975), .A2(n9972), .A3(n9761), .ZN(n9971) );
  XNOR2_X1 U13230 ( .A(n12850), .B(n9983), .ZN(n12851) );
  NAND2_X2 U13231 ( .A1(n9984), .A2(n12797), .ZN(n17926) );
  NOR2_X1 U13232 ( .A1(n9986), .A2(n9985), .ZN(n9984) );
  NAND2_X1 U13233 ( .A1(n12793), .A2(n12794), .ZN(n9985) );
  NAND2_X1 U13234 ( .A1(n12795), .A2(n12796), .ZN(n9986) );
  NOR2_X2 U13235 ( .A1(n12620), .A2(n19179), .ZN(n17732) );
  NAND2_X2 U13236 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19179) );
  AND2_X1 U13237 ( .A1(n9991), .A2(n9989), .ZN(n13044) );
  OR2_X1 U13238 ( .A1(n13026), .A2(n9992), .ZN(n9991) );
  NAND4_X1 U13239 ( .A1(n18208), .A2(n18561), .A3(n18196), .A4(n9996), .ZN(
        n9995) );
  OR2_X2 U13240 ( .A1(n16342), .A2(n9795), .ZN(n16309) );
  NAND2_X2 U13241 ( .A1(n16360), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16342) );
  INV_X2 U13243 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12709) );
  INV_X1 U13244 ( .A(n18335), .ZN(n9998) );
  NAND2_X1 U13245 ( .A1(n11999), .A2(n12412), .ZN(n11996) );
  AND2_X2 U13246 ( .A1(n11868), .A2(n13703), .ZN(n11880) );
  AND3_X2 U13247 ( .A1(n11861), .A2(n11859), .A3(n11860), .ZN(n13873) );
  NAND2_X2 U13248 ( .A1(n10002), .A2(n10001), .ZN(n10405) );
  NAND2_X1 U13249 ( .A1(n11813), .A2(n11812), .ZN(n11822) );
  INV_X1 U13250 ( .A(n10003), .ZN(n10002) );
  NAND2_X1 U13251 ( .A1(n10004), .A2(n12405), .ZN(n14204) );
  NAND2_X1 U13252 ( .A1(n13963), .A2(n12402), .ZN(n10004) );
  NAND2_X1 U13253 ( .A1(n10005), .A2(n15927), .ZN(n13963) );
  NAND3_X1 U13254 ( .A1(n11920), .A2(n12048), .A3(n10541), .ZN(n10005) );
  INV_X1 U13255 ( .A(n10155), .ZN(n10006) );
  AOI21_X1 U13256 ( .B1(n10006), .B2(n16210), .A(n10008), .ZN(n10010) );
  INV_X1 U13257 ( .A(n10156), .ZN(n10007) );
  NAND2_X1 U13258 ( .A1(n10007), .A2(n16210), .ZN(n10009) );
  NAND3_X1 U13259 ( .A1(n10159), .A2(n16230), .A3(n10011), .ZN(n12515) );
  NAND4_X1 U13260 ( .A1(n11811), .A2(n13534), .A3(n12323), .A4(n11773), .ZN(
        n11813) );
  CLKBUF_X1 U13261 ( .A(n10405), .Z(n10014) );
  NAND2_X1 U13262 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12208) );
  NAND2_X1 U13263 ( .A1(n10014), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12215) );
  NAND2_X1 U13264 ( .A1(n10405), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11836) );
  NAND2_X1 U13265 ( .A1(n10405), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11814) );
  NAND2_X1 U13266 ( .A1(n10405), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11832) );
  NAND2_X1 U13267 ( .A1(n11863), .A2(n10018), .ZN(n10017) );
  INV_X1 U13268 ( .A(n11781), .ZN(n10019) );
  AND3_X2 U13269 ( .A1(n10019), .A2(n9731), .A3(n11779), .ZN(n12209) );
  CLKBUF_X1 U13270 ( .A(n13627), .Z(n10020) );
  NAND3_X1 U13271 ( .A1(n14645), .A2(n14644), .A3(n10022), .ZN(P2_U3012) );
  XNOR2_X2 U13272 ( .A(n13764), .B(n13763), .ZN(n19598) );
  NAND2_X1 U13273 ( .A1(n10034), .A2(n10240), .ZN(n15186) );
  INV_X1 U13274 ( .A(n15199), .ZN(n10033) );
  INV_X1 U13275 ( .A(n15200), .ZN(n10034) );
  NAND2_X2 U13276 ( .A1(n20607), .A2(n10880), .ZN(n10879) );
  NAND3_X1 U13277 ( .A1(n10967), .A2(n10949), .A3(n9718), .ZN(n13166) );
  NAND3_X1 U13278 ( .A1(n10041), .A2(n10042), .A3(n10039), .ZN(n10354) );
  NAND3_X1 U13279 ( .A1(n10040), .A2(n14352), .A3(n13251), .ZN(n10039) );
  AND2_X4 U13280 ( .A1(n10046), .A2(n11564), .ZN(n11718) );
  AND2_X4 U13281 ( .A1(n10046), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11731) );
  NAND2_X1 U13282 ( .A1(n10048), .A2(n11839), .ZN(n10047) );
  NAND4_X1 U13283 ( .A1(n11710), .A2(n11712), .A3(n11709), .A4(n11711), .ZN(
        n10048) );
  NAND4_X1 U13284 ( .A1(n11705), .A2(n11708), .A3(n11707), .A4(n11706), .ZN(
        n10050) );
  NAND2_X1 U13285 ( .A1(n12319), .A2(n9691), .ZN(n11797) );
  NAND2_X1 U13286 ( .A1(n11789), .A2(n10051), .ZN(n12319) );
  NAND2_X1 U13287 ( .A1(n10052), .A2(n11788), .ZN(n10051) );
  NAND2_X1 U13288 ( .A1(n11804), .A2(n11786), .ZN(n10052) );
  NAND3_X1 U13289 ( .A1(n10055), .A2(n13024), .A3(n10054), .ZN(P2_U2987) );
  OR2_X1 U13290 ( .A1(n13025), .A2(n16439), .ZN(n10054) );
  NAND3_X1 U13291 ( .A1(n12740), .A2(n10056), .A3(n16383), .ZN(n10055) );
  AND2_X1 U13292 ( .A1(n12339), .A2(n10062), .ZN(n11765) );
  CLKBUF_X1 U13293 ( .A(n10074), .Z(n10063) );
  NAND3_X1 U13294 ( .A1(n12927), .A2(n10082), .A3(n10303), .ZN(n10081) );
  NAND3_X1 U13295 ( .A1(n12927), .A2(n10303), .A3(n13038), .ZN(n13276) );
  AND2_X1 U13296 ( .A1(n10084), .A2(n9783), .ZN(n12929) );
  NAND3_X1 U13297 ( .A1(n9722), .A2(n10085), .A3(n12814), .ZN(n12891) );
  NAND3_X1 U13298 ( .A1(n11784), .A2(n16778), .A3(n10090), .ZN(n11799) );
  NAND2_X1 U13299 ( .A1(n13884), .A2(n10090), .ZN(n13906) );
  NAND2_X1 U13300 ( .A1(n10092), .A2(n11839), .ZN(n10091) );
  NAND4_X1 U13301 ( .A1(n11600), .A2(n11601), .A3(n11598), .A4(n11599), .ZN(
        n10092) );
  NAND2_X1 U13302 ( .A1(n10094), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10093) );
  NAND4_X1 U13303 ( .A1(n11597), .A2(n11596), .A3(n11594), .A4(n11595), .ZN(
        n10094) );
  NAND2_X1 U13304 ( .A1(n15993), .A2(n10097), .ZN(n10101) );
  INV_X1 U13305 ( .A(n15996), .ZN(n10098) );
  NAND2_X1 U13306 ( .A1(n13626), .A2(n10106), .ZN(n20254) );
  NAND2_X1 U13307 ( .A1(n10423), .A2(n10107), .ZN(n10106) );
  INV_X1 U13308 ( .A(n13526), .ZN(n10107) );
  NAND2_X1 U13309 ( .A1(n10108), .A2(n13526), .ZN(n13626) );
  INV_X1 U13310 ( .A(n10423), .ZN(n10108) );
  NAND2_X1 U13311 ( .A1(n10111), .A2(n10109), .ZN(P2_U2890) );
  NAND3_X1 U13312 ( .A1(n16062), .A2(n19437), .A3(n15978), .ZN(n10111) );
  NAND2_X1 U13313 ( .A1(n10113), .A2(n15977), .ZN(n15978) );
  NAND4_X1 U13314 ( .A1(n11817), .A2(n11814), .A3(n11816), .A4(n11815), .ZN(
        n10124) );
  NAND2_X1 U13315 ( .A1(n14203), .A2(n11976), .ZN(n10509) );
  NAND2_X1 U13316 ( .A1(n10161), .A2(n10357), .ZN(n10128) );
  NAND2_X1 U13317 ( .A1(n10128), .A2(n10356), .ZN(n11920) );
  NAND2_X1 U13318 ( .A1(n10879), .A2(n10137), .ZN(n10139) );
  NAND2_X1 U13319 ( .A1(n10138), .A2(n10866), .ZN(n10143) );
  NAND2_X1 U13320 ( .A1(n10139), .A2(n10140), .ZN(n10138) );
  INV_X1 U13321 ( .A(n14827), .ZN(n10145) );
  NAND2_X1 U13322 ( .A1(n10145), .A2(n10146), .ZN(n14784) );
  XNOR2_X1 U13323 ( .A(n13199), .B(n13198), .ZN(n13749) );
  AND2_X2 U13324 ( .A1(n10152), .A2(n10154), .ZN(n13181) );
  NAND2_X1 U13325 ( .A1(n10157), .A2(n16438), .ZN(n16371) );
  XNOR2_X1 U13326 ( .A(n16438), .B(n10157), .ZN(n16703) );
  NAND2_X1 U13327 ( .A1(n9672), .A2(n11919), .ZN(n10161) );
  NAND2_X1 U13328 ( .A1(n10509), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10162) );
  NAND2_X1 U13329 ( .A1(n16574), .A2(n10164), .ZN(n14339) );
  AOI22_X1 U13330 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11647) );
  NAND2_X1 U13331 ( .A1(n10966), .A2(n10965), .ZN(n13982) );
  NOR2_X1 U13332 ( .A1(n14706), .A2(n14708), .ZN(n14691) );
  INV_X4 U13333 ( .A(n10813), .ZN(n14013) );
  NAND2_X1 U13334 ( .A1(n10240), .A2(n10239), .ZN(n15163) );
  NOR2_X1 U13335 ( .A1(n18305), .A2(n18304), .ZN(n18303) );
  NOR2_X2 U13336 ( .A1(n18393), .A2(n18392), .ZN(n18401) );
  AOI21_X1 U13337 ( .B1(n15163), .B2(n15154), .A(n13243), .ZN(n15153) );
  XNOR2_X1 U13338 ( .A(n10354), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15286) );
  NOR2_X1 U13339 ( .A1(n15200), .A2(n9687), .ZN(n10239) );
  OAI211_X1 U13340 ( .C1(n16466), .C2(n16429), .A(n10393), .B(n10392), .ZN(
        P2_U2988) );
  NAND2_X1 U13341 ( .A1(n10371), .A2(n16830), .ZN(n16842) );
  OR2_X2 U13342 ( .A1(n15707), .A2(n15710), .ZN(n13104) );
  AOI21_X2 U13343 ( .B1(n15587), .B2(n19409), .A(n15588), .ZN(n13126) );
  NAND2_X1 U13344 ( .A1(n10238), .A2(n10830), .ZN(n13467) );
  INV_X1 U13345 ( .A(n10500), .ZN(n11381) );
  INV_X2 U13346 ( .A(n14784), .ZN(n11300) );
  NOR2_X2 U13347 ( .A1(n10167), .A2(n14229), .ZN(n12842) );
  NAND2_X1 U13348 ( .A1(n12708), .A2(n10183), .ZN(n10182) );
  INV_X1 U13349 ( .A(n10189), .ZN(n17802) );
  NOR2_X2 U13350 ( .A1(n12699), .A2(n12696), .ZN(n12886) );
  NAND2_X2 U13351 ( .A1(n9682), .A2(n10190), .ZN(n17826) );
  NAND3_X1 U13352 ( .A1(n12645), .A2(n12646), .A3(n10192), .ZN(n10191) );
  INV_X1 U13353 ( .A(n11777), .ZN(n12369) );
  NAND2_X2 U13354 ( .A1(n11725), .A2(n11724), .ZN(n11777) );
  NAND2_X2 U13355 ( .A1(n10194), .A2(n11654), .ZN(n11778) );
  NAND3_X1 U13356 ( .A1(n11649), .A2(n9689), .A3(n11648), .ZN(n10194) );
  INV_X1 U13357 ( .A(n12383), .ZN(n12367) );
  OAI211_X1 U13358 ( .C1(n14349), .C2(n16429), .A(n10196), .B(n10195), .ZN(
        P2_U2983) );
  NAND2_X1 U13359 ( .A1(n14348), .A2(n16426), .ZN(n10196) );
  NAND2_X1 U13360 ( .A1(n12582), .A2(n12581), .ZN(n10198) );
  XNOR2_X2 U13361 ( .A(n12203), .B(n11835), .ZN(n13627) );
  INV_X2 U13362 ( .A(n12209), .ZN(n12218) );
  NAND2_X1 U13363 ( .A1(n11840), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10204) );
  AND2_X2 U13364 ( .A1(n11799), .A2(n11798), .ZN(n11840) );
  NOR2_X2 U13365 ( .A1(n12423), .A2(n12543), .ZN(n12475) );
  AND2_X4 U13366 ( .A1(n15518), .A2(n13457), .ZN(n10883) );
  NOR2_X4 U13367 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15518) );
  OAI21_X1 U13368 ( .B1(n10228), .B2(n11189), .A(n11026), .ZN(n14068) );
  NAND2_X1 U13369 ( .A1(n11022), .A2(n11021), .ZN(n10228) );
  INV_X1 U13370 ( .A(n11439), .ZN(n10229) );
  AND3_X2 U13371 ( .A1(n10229), .A2(n10846), .A3(n10820), .ZN(n10238) );
  INV_X2 U13372 ( .A(n10230), .ZN(n10846) );
  NAND2_X1 U13373 ( .A1(n11455), .A2(n20532), .ZN(n10230) );
  NAND2_X1 U13374 ( .A1(n10234), .A2(n10231), .ZN(n10352) );
  INV_X1 U13375 ( .A(n13249), .ZN(n15147) );
  NAND2_X1 U13376 ( .A1(n11973), .A2(n12367), .ZN(n11978) );
  NOR2_X2 U13377 ( .A1(n10818), .A2(n10237), .ZN(n11434) );
  NAND2_X1 U13378 ( .A1(n10238), .A2(n13255), .ZN(n13472) );
  NAND2_X1 U13379 ( .A1(n10968), .A2(n10967), .ZN(n10995) );
  INV_X1 U13380 ( .A(n10949), .ZN(n15561) );
  NAND2_X1 U13381 ( .A1(n15095), .A2(n15216), .ZN(n10241) );
  INV_X1 U13382 ( .A(n13247), .ZN(n10246) );
  NAND3_X1 U13383 ( .A1(n10246), .A2(n15218), .A3(n10245), .ZN(n10247) );
  NAND2_X1 U13384 ( .A1(n13247), .A2(n13246), .ZN(n10389) );
  OAI22_X1 U13385 ( .A1(n10249), .A2(n10250), .B1(n19696), .B2(n11872), .ZN(
        n11873) );
  OAI21_X1 U13386 ( .B1(n9621), .B2(n20044), .A(n20104), .ZN(n10251) );
  CLKBUF_X1 U13387 ( .A(n16267), .Z(n10253) );
  NAND3_X1 U13388 ( .A1(n14328), .A2(n14327), .A3(n10515), .ZN(n10259) );
  AND2_X1 U13389 ( .A1(n19194), .A2(n19195), .ZN(n19192) );
  NAND2_X1 U13390 ( .A1(n10264), .A2(n19190), .ZN(n19194) );
  INV_X2 U13391 ( .A(n19182), .ZN(n19169) );
  NAND2_X2 U13392 ( .A1(n10271), .A2(n10269), .ZN(n19182) );
  XNOR2_X1 U13393 ( .A(n12851), .B(n18682), .ZN(n18364) );
  NAND2_X2 U13394 ( .A1(n18618), .A2(n10304), .ZN(n18292) );
  AND2_X2 U13395 ( .A1(n10278), .A2(n18261), .ZN(n18618) );
  OAI21_X1 U13396 ( .B1(n18301), .B2(n12864), .A(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10278) );
  NAND3_X1 U13397 ( .A1(n10820), .A2(n10846), .A3(n13722), .ZN(n10845) );
  INV_X1 U13398 ( .A(n11434), .ZN(n13746) );
  INV_X2 U13399 ( .A(n10819), .ZN(n20520) );
  XNOR2_X1 U13400 ( .A(n10583), .B(n15427), .ZN(n15166) );
  NOR2_X2 U13401 ( .A1(n17104), .A2(n19360), .ZN(n18375) );
  NAND3_X1 U13402 ( .A1(n19184), .A2(n19169), .A3(n10297), .ZN(n18450) );
  NAND3_X1 U13403 ( .A1(n19184), .A2(n19169), .A3(n9641), .ZN(n10301) );
  OAI21_X1 U13404 ( .B1(n18363), .B2(n18364), .A(n9686), .ZN(n10302) );
  OR2_X2 U13405 ( .A1(n18302), .A2(n18306), .ZN(n10394) );
  INV_X1 U13406 ( .A(n10308), .ZN(n17209) );
  INV_X1 U13407 ( .A(n10306), .ZN(n17208) );
  NAND2_X1 U13409 ( .A1(n17217), .A2(n10321), .ZN(n10308) );
  NAND2_X1 U13411 ( .A1(n10309), .A2(n9643), .ZN(n12602) );
  NOR2_X1 U13412 ( .A1(n17189), .A2(n18095), .ZN(n17188) );
  AOI21_X1 U13413 ( .B1(n17189), .B2(n10321), .A(n10315), .ZN(n10314) );
  AND2_X2 U13414 ( .A1(n18054), .A2(n10322), .ZN(n12612) );
  NAND2_X1 U13416 ( .A1(n14204), .A2(n14205), .ZN(n10333) );
  NAND3_X1 U13417 ( .A1(n18379), .A2(n17926), .A3(n12850), .ZN(n10338) );
  NAND2_X1 U13418 ( .A1(n18361), .A2(n18362), .ZN(n18360) );
  XNOR2_X1 U13419 ( .A(n12902), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18361) );
  NAND2_X1 U13420 ( .A1(n11871), .A2(n11880), .ZN(n19696) );
  OR2_X1 U13421 ( .A1(n16778), .A2(n14561), .ZN(n10358) );
  NAND2_X4 U13422 ( .A1(n10360), .A2(n10359), .ZN(n16778) );
  NAND2_X1 U13423 ( .A1(n10367), .A2(n10366), .ZN(n10365) );
  NAND2_X1 U13424 ( .A1(n9596), .A2(n9708), .ZN(n10371) );
  OAI21_X1 U13425 ( .B1(n13126), .B2(n16750), .A(n13125), .ZN(n14364) );
  NAND2_X1 U13426 ( .A1(n13077), .A2(n10376), .ZN(n13084) );
  INV_X1 U13427 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10379) );
  NAND2_X1 U13428 ( .A1(n13092), .A2(n9764), .ZN(n13098) );
  NAND3_X1 U13429 ( .A1(n10383), .A2(n10382), .A3(n10381), .ZN(n10384) );
  NAND2_X1 U13430 ( .A1(n18379), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18372) );
  OAI21_X1 U13431 ( .B1(n12864), .B2(n18301), .A(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12890) );
  NOR2_X1 U13432 ( .A1(n12864), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10395) );
  NAND2_X1 U13433 ( .A1(n12859), .A2(n10399), .ZN(n10398) );
  INV_X2 U13434 ( .A(n10583), .ZN(n15216) );
  NAND2_X1 U13435 ( .A1(n10583), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15185) );
  INV_X2 U13436 ( .A(n12331), .ZN(n11785) );
  NAND2_X2 U13437 ( .A1(n10404), .A2(n11574), .ZN(n12331) );
  NAND3_X1 U13438 ( .A1(n11573), .A2(n11572), .A3(n10569), .ZN(n10404) );
  NAND2_X1 U13439 ( .A1(n12229), .A2(n9640), .ZN(n13826) );
  AND2_X1 U13440 ( .A1(n12994), .A2(n12995), .ZN(n12997) );
  NAND4_X1 U13441 ( .A1(n10415), .A2(n12213), .A3(n12212), .A4(n10417), .ZN(
        n13835) );
  AND2_X1 U13442 ( .A1(n10579), .A2(n15703), .ZN(n15637) );
  NAND3_X1 U13443 ( .A1(n10425), .A2(n10427), .A3(n10424), .ZN(n16003) );
  NOR2_X1 U13444 ( .A1(n14519), .A2(n10428), .ZN(n10426) );
  NAND2_X1 U13445 ( .A1(n14519), .A2(n10428), .ZN(n10427) );
  INV_X1 U13446 ( .A(n14501), .ZN(n10428) );
  NAND2_X1 U13447 ( .A1(n15989), .A2(n10437), .ZN(n10435) );
  NAND2_X1 U13448 ( .A1(n10434), .A2(n10429), .ZN(n14622) );
  AOI21_X1 U13449 ( .B1(n15989), .B2(n10430), .A(n14596), .ZN(n10429) );
  NOR2_X1 U13450 ( .A1(n16056), .A2(n10438), .ZN(n16039) );
  INV_X1 U13451 ( .A(n16056), .ZN(n16053) );
  INV_X1 U13452 ( .A(n10578), .ZN(n10442) );
  CLKBUF_X1 U13453 ( .A(n14447), .Z(n10447) );
  AOI21_X1 U13454 ( .B1(n14601), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A(n9746), .ZN(n14506) );
  NAND2_X1 U13455 ( .A1(n12519), .A2(n10448), .ZN(n12520) );
  OAI21_X1 U13456 ( .B1(n12541), .B2(n16838), .A(n10450), .ZN(n10449) );
  INV_X1 U13457 ( .A(n15630), .ZN(n10450) );
  NAND2_X1 U13458 ( .A1(n9638), .A2(n9735), .ZN(n10451) );
  NAND2_X1 U13459 ( .A1(n12517), .A2(n10453), .ZN(n12529) );
  AND2_X4 U13460 ( .A1(n10457), .A2(n11564), .ZN(n14509) );
  AND2_X1 U13461 ( .A1(n14443), .A2(n10457), .ZN(n14474) );
  AND2_X2 U13462 ( .A1(n11563), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10457) );
  AOI21_X1 U13463 ( .B1(n11823), .B2(n9636), .A(n9763), .ZN(n11818) );
  AOI21_X1 U13464 ( .B1(n12230), .B2(P2_REIP_REG_3__SCAN_IN), .A(n9765), .ZN(
        n11837) );
  OAI21_X1 U13465 ( .B1(n16195), .B2(n16197), .A(n10458), .ZN(n10462) );
  NAND2_X1 U13466 ( .A1(n16195), .A2(n10459), .ZN(n10458) );
  NAND2_X1 U13467 ( .A1(n16191), .A2(n10461), .ZN(n10460) );
  AND2_X1 U13468 ( .A1(n16197), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10461) );
  NAND2_X1 U13469 ( .A1(n16195), .A2(n10464), .ZN(n10463) );
  INV_X1 U13470 ( .A(n16197), .ZN(n10464) );
  AND2_X2 U13471 ( .A1(n10465), .A2(n10605), .ZN(n10705) );
  NAND2_X1 U13472 ( .A1(n14702), .A2(n10469), .ZN(n10466) );
  AND2_X1 U13473 ( .A1(n14702), .A2(n10470), .ZN(n11557) );
  NAND2_X1 U13474 ( .A1(n14702), .A2(n10471), .ZN(n14672) );
  NAND2_X1 U13475 ( .A1(n14702), .A2(n14703), .ZN(n14705) );
  AND2_X1 U13476 ( .A1(n10471), .A2(n14673), .ZN(n10469) );
  NAND2_X1 U13477 ( .A1(n11482), .A2(n9727), .ZN(n15504) );
  INV_X1 U13478 ( .A(n15504), .ZN(n11495) );
  NAND2_X1 U13479 ( .A1(n14799), .A2(n10483), .ZN(n14733) );
  NAND2_X1 U13480 ( .A1(n15631), .A2(n9773), .ZN(n13009) );
  NAND2_X1 U13481 ( .A1(n15631), .A2(n10492), .ZN(n15595) );
  AND2_X1 U13482 ( .A1(n15631), .A2(n12747), .ZN(n15594) );
  INV_X1 U13483 ( .A(n14109), .ZN(n10493) );
  NAND2_X1 U13484 ( .A1(n10493), .A2(n10494), .ZN(n14827) );
  NAND2_X1 U13485 ( .A1(n14718), .A2(n14720), .ZN(n14706) );
  NAND2_X1 U13486 ( .A1(n11300), .A2(n9726), .ZN(n14731) );
  NAND2_X1 U13487 ( .A1(n11920), .A2(n10541), .ZN(n10507) );
  NAND2_X1 U13488 ( .A1(n10507), .A2(n10506), .ZN(n13978) );
  INV_X1 U13489 ( .A(n13967), .ZN(n10506) );
  NAND2_X1 U13490 ( .A1(n10509), .A2(n10508), .ZN(n16431) );
  AND2_X1 U13491 ( .A1(n10253), .A2(n12359), .ZN(n16237) );
  AND2_X2 U13492 ( .A1(n16219), .A2(n10511), .ZN(n12987) );
  OAI21_X1 U13493 ( .B1(n16354), .B2(n16351), .A(n16352), .ZN(n16338) );
  AOI21_X1 U13494 ( .B1(n16351), .B2(n16352), .A(n10531), .ZN(n10530) );
  INV_X1 U13495 ( .A(n16339), .ZN(n10531) );
  OAI21_X1 U13496 ( .B1(n16248), .B2(n10537), .A(n10533), .ZN(n10539) );
  INV_X1 U13497 ( .A(n16247), .ZN(n10535) );
  INV_X1 U13498 ( .A(n16246), .ZN(n10540) );
  AND2_X2 U13499 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11581) );
  NAND2_X1 U13500 ( .A1(n16205), .A2(n12526), .ZN(n10545) );
  NAND2_X1 U13501 ( .A1(n12514), .A2(n9749), .ZN(n10547) );
  XNOR2_X1 U13502 ( .A(n12558), .B(n12557), .ZN(n14349) );
  NAND2_X1 U13503 ( .A1(n13017), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13075) );
  INV_X1 U13504 ( .A(n13071), .ZN(n13017) );
  NAND2_X1 U13505 ( .A1(n13115), .A2(n16224), .ZN(n15661) );
  AND2_X1 U13506 ( .A1(n14193), .A2(n14195), .ZN(n16583) );
  INV_X1 U13507 ( .A(n13181), .ZN(n10975) );
  OAI22_X1 U13508 ( .A1(n19325), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n19193), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12716) );
  INV_X4 U13509 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19325) );
  OR2_X1 U13510 ( .A1(n15216), .A2(n15512), .ZN(n13237) );
  OR2_X1 U13511 ( .A1(n15216), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15048) );
  INV_X1 U13512 ( .A(n16309), .ZN(n14323) );
  OR2_X1 U13513 ( .A1(n13632), .A2(n13631), .ZN(n13633) );
  CLKBUF_X1 U13514 ( .A(n16360), .Z(n16382) );
  INV_X1 U13515 ( .A(n12438), .ZN(n12440) );
  NOR2_X1 U13516 ( .A1(n10548), .A2(n13012), .ZN(n13013) );
  NAND2_X1 U13517 ( .A1(n11495), .A2(n11494), .ZN(n15506) );
  AND2_X2 U13518 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15519) );
  INV_X1 U13519 ( .A(n12987), .ZN(n12740) );
  XNOR2_X1 U13520 ( .A(n12987), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16453) );
  NAND4_X4 U13521 ( .A1(n10767), .A2(n10766), .A3(n10765), .A4(n10764), .ZN(
        n10813) );
  CLKBUF_X1 U13522 ( .A(n13467), .Z(n13707) );
  NAND2_X1 U13523 ( .A1(n11840), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11826) );
  INV_X1 U13524 ( .A(n11787), .ZN(n11788) );
  NAND2_X1 U13525 ( .A1(n16179), .A2(n16689), .ZN(n12555) );
  INV_X1 U13526 ( .A(n12517), .ZN(n15664) );
  AOI22_X1 U13527 ( .A1(n14447), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11733), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11719) );
  NAND2_X1 U13528 ( .A1(n11863), .A2(n11875), .ZN(n11905) );
  CLKBUF_X1 U13529 ( .A(n13873), .Z(n15933) );
  NAND2_X1 U13530 ( .A1(n13873), .A2(n9838), .ZN(n13697) );
  AOI22_X1 U13531 ( .A1(n12230), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11833) );
  NOR2_X1 U13532 ( .A1(n10842), .A2(n13361), .ZN(n13473) );
  CLKBUF_X1 U13533 ( .A(n11718), .Z(n14597) );
  AOI22_X1 U13534 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9604), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11707) );
  AND2_X1 U13535 ( .A1(n11773), .A2(n11772), .ZN(n11805) );
  AND2_X2 U13536 ( .A1(n13627), .A2(n13703), .ZN(n11876) );
  AND2_X1 U13537 ( .A1(n16188), .A2(n16689), .ZN(n10548) );
  AND2_X1 U13538 ( .A1(n14358), .A2(n13055), .ZN(n19404) );
  NOR2_X1 U13539 ( .A1(n12750), .A2(n10552), .ZN(n10549) );
  INV_X1 U13540 ( .A(n16706), .ZN(n12739) );
  AND2_X1 U13541 ( .A1(n11733), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10550) );
  NOR2_X1 U13542 ( .A1(n13259), .A2(n20833), .ZN(n10551) );
  AND2_X1 U13543 ( .A1(n16081), .A2(n16724), .ZN(n10552) );
  NOR2_X1 U13544 ( .A1(n20874), .A2(n20873), .ZN(n10553) );
  INV_X1 U13545 ( .A(n20061), .ZN(n20149) );
  OR2_X1 U13546 ( .A1(n20031), .A2(n20030), .ZN(n20061) );
  OR2_X1 U13547 ( .A1(n18239), .A2(n12920), .ZN(n10554) );
  AND2_X1 U13548 ( .A1(n15409), .A2(n15385), .ZN(n10555) );
  OR2_X1 U13549 ( .A1(n20508), .A2(n13346), .ZN(n10556) );
  OR2_X1 U13550 ( .A1(n11841), .A2(n20262), .ZN(n10557) );
  OR2_X1 U13551 ( .A1(n12532), .A2(n12450), .ZN(n10558) );
  AND2_X1 U13552 ( .A1(n11918), .A2(n10064), .ZN(n10559) );
  AND2_X1 U13553 ( .A1(n14454), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10560) );
  AND2_X1 U13554 ( .A1(n13148), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10561) );
  AND3_X1 U13555 ( .A1(n11651), .A2(n11839), .A3(n11650), .ZN(n10562) );
  NAND2_X1 U13556 ( .A1(n10829), .A2(n10828), .ZN(n10842) );
  INV_X1 U13557 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16437) );
  AND2_X1 U13558 ( .A1(n13338), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n16771)
         );
  AND2_X1 U13559 ( .A1(n11374), .A2(P1_EAX_REG_5__SCAN_IN), .ZN(n10563) );
  INV_X1 U13560 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12605) );
  AND3_X1 U13561 ( .A1(n16377), .A2(n16372), .A3(n16390), .ZN(n10564) );
  AND2_X1 U13562 ( .A1(n12480), .A2(n16307), .ZN(n10565) );
  AND2_X1 U13563 ( .A1(n11242), .A2(n11241), .ZN(n10566) );
  INV_X1 U13564 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12853) );
  INV_X1 U13565 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18288) );
  INV_X1 U13566 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18613) );
  INV_X1 U13567 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15778) );
  NOR2_X1 U13568 ( .A1(n16376), .A2(n16389), .ZN(n10567) );
  NAND2_X1 U13569 ( .A1(n13354), .A2(n13129), .ZN(n15936) );
  INV_X1 U13570 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11639) );
  OR2_X1 U13571 ( .A1(n19431), .A2(n19577), .ZN(n16165) );
  INV_X1 U13572 ( .A(n16165), .ZN(n19433) );
  AND2_X1 U13573 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10568) );
  INV_X1 U13574 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18413) );
  INV_X1 U13575 ( .A(n15994), .ZN(n14535) );
  INV_X1 U13576 ( .A(n15297), .ZN(n11561) );
  AND3_X1 U13577 ( .A1(n11571), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11570), .ZN(n10569) );
  INV_X1 U13578 ( .A(n13823), .ZN(n13824) );
  NAND2_X1 U13579 ( .A1(n10983), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11189) );
  INV_X1 U13580 ( .A(n11189), .ZN(n14127) );
  OR3_X1 U13581 ( .A1(n19360), .A2(n18721), .A3(n19212), .ZN(n10570) );
  INV_X1 U13582 ( .A(n20453), .ZN(n13552) );
  AND4_X1 U13583 ( .A1(n11666), .A2(n11665), .A3(n11664), .A4(n11663), .ZN(
        n10571) );
  NAND2_X1 U13584 ( .A1(n10144), .A2(n20496), .ZN(n20649) );
  AND2_X1 U13585 ( .A1(n20396), .A2(n20532), .ZN(n20392) );
  NAND2_X1 U13586 ( .A1(n14007), .A2(n14006), .ZN(n21173) );
  AND2_X1 U13587 ( .A1(n10835), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10572) );
  OR2_X1 U13588 ( .A1(n14007), .A2(n20508), .ZN(n13588) );
  AND3_X1 U13589 ( .A1(n14148), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n12403), .ZN(n10573) );
  OR2_X1 U13590 ( .A1(n18228), .A2(n18391), .ZN(n10574) );
  AND2_X1 U13591 ( .A1(n13038), .A2(n18616), .ZN(n10575) );
  OR2_X1 U13592 ( .A1(n13259), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14136) );
  INV_X1 U13593 ( .A(n14136), .ZN(n16962) );
  NOR2_X1 U13594 ( .A1(n13268), .A2(n13267), .ZN(n10576) );
  OR2_X1 U13595 ( .A1(n12605), .A2(n17471), .ZN(n10577) );
  INV_X1 U13596 ( .A(n13854), .ZN(n14611) );
  OR2_X1 U13597 ( .A1(n14390), .A2(n14389), .ZN(n10578) );
  AND2_X1 U13598 ( .A1(n13696), .A2(n13695), .ZN(n10580) );
  AND2_X1 U13599 ( .A1(n10907), .A2(n13183), .ZN(n10582) );
  INV_X1 U13600 ( .A(n14010), .ZN(n10812) );
  NOR2_X1 U13601 ( .A1(n20532), .A2(n21074), .ZN(n10986) );
  INV_X1 U13602 ( .A(n11390), .ZN(n11442) );
  AND2_X1 U13603 ( .A1(n11396), .A2(n11395), .ZN(n11402) );
  NAND2_X1 U13604 ( .A1(n11390), .A2(n20512), .ZN(n10824) );
  AND2_X1 U13605 ( .A1(n11424), .A2(n11412), .ZN(n11422) );
  OR2_X1 U13606 ( .A1(n11016), .A2(n11015), .ZN(n13215) );
  AOI22_X1 U13607 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n14463), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11620) );
  NAND2_X1 U13608 ( .A1(n20873), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11424) );
  NAND2_X1 U13609 ( .A1(n13254), .A2(n20516), .ZN(n10828) );
  OR2_X1 U13610 ( .A1(n11018), .A2(n11017), .ZN(n11019) );
  INV_X1 U13611 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n12516) );
  NAND2_X1 U13612 ( .A1(n11800), .A2(n11687), .ZN(n11688) );
  AND2_X1 U13613 ( .A1(n16211), .A2(n12525), .ZN(n12526) );
  AOI22_X1 U13614 ( .A1(n14454), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11733), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11709) );
  INV_X1 U13615 ( .A(n10826), .ZN(n10830) );
  INV_X1 U13616 ( .A(n11024), .ZN(n11025) );
  INV_X1 U13617 ( .A(n11262), .ZN(n10591) );
  OR2_X1 U13618 ( .A1(n10893), .A2(n10892), .ZN(n13183) );
  AND4_X1 U13619 ( .A1(n10727), .A2(n10726), .A3(n10725), .A4(n10724), .ZN(
        n10728) );
  AND2_X1 U13620 ( .A1(n16011), .A2(n16009), .ZN(n14499) );
  INV_X1 U13621 ( .A(n15689), .ZN(n12175) );
  NAND2_X1 U13622 ( .A1(n12842), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12788) );
  INV_X1 U13623 ( .A(n11419), .ZN(n11430) );
  NOR2_X1 U13624 ( .A1(n13453), .A2(n11451), .ZN(n13730) );
  INV_X1 U13625 ( .A(n11333), .ZN(n10593) );
  INV_X1 U13626 ( .A(n11301), .ZN(n10592) );
  AND2_X1 U13627 ( .A1(n10591), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11277) );
  AND2_X1 U13628 ( .A1(n14108), .A2(n14111), .ZN(n11108) );
  OR2_X1 U13629 ( .A1(n10959), .A2(n10958), .ZN(n13172) );
  NAND2_X1 U13630 ( .A1(n10935), .A2(n10934), .ZN(n20644) );
  AND2_X1 U13631 ( .A1(n12374), .A2(n12375), .ZN(n11690) );
  INV_X1 U13632 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n12449) );
  OR2_X1 U13633 ( .A1(n12532), .A2(n13634), .ZN(n12373) );
  AND2_X1 U13634 ( .A1(n14495), .A2(n14494), .ZN(n16007) );
  CLKBUF_X3 U13635 ( .A(n11942), .Z(n14462) );
  INV_X1 U13636 ( .A(n14160), .ZN(n12258) );
  INV_X1 U13637 ( .A(n11901), .ZN(n12022) );
  INV_X1 U13638 ( .A(n12412), .ZN(n12048) );
  AND2_X1 U13639 ( .A1(n11759), .A2(n11758), .ZN(n12337) );
  AOI21_X1 U13640 ( .B1(n12230), .B2(P2_REIP_REG_0__SCAN_IN), .A(n11802), .ZN(
        n11817) );
  INV_X1 U13641 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n21273) );
  OR2_X1 U13642 ( .A1(n10304), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12928) );
  INV_X1 U13643 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n21222) );
  INV_X1 U13644 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n21256) );
  NAND2_X1 U13645 ( .A1(n11277), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11301) );
  OR2_X1 U13646 ( .A1(n15138), .A2(n11371), .ZN(n11261) );
  INV_X1 U13647 ( .A(n11043), .ZN(n10585) );
  INV_X1 U13648 ( .A(n15047), .ZN(n13252) );
  OR2_X1 U13649 ( .A1(n10839), .A2(n13458), .ZN(n13728) );
  INV_X1 U13650 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15523) );
  INV_X1 U13651 ( .A(n20540), .ZN(n20609) );
  INV_X1 U13652 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20836) );
  AND3_X1 U13653 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n10144), .A3(n20496), 
        .ZN(n20533) );
  INV_X1 U13654 ( .A(n13772), .ZN(n12212) );
  INV_X1 U13655 ( .A(n13934), .ZN(n12241) );
  OR2_X1 U13656 ( .A1(n14555), .A2(n14560), .ZN(n14591) );
  OR2_X1 U13657 ( .A1(n14481), .A2(n14480), .ZN(n14497) );
  INV_X1 U13658 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16654) );
  INV_X1 U13659 ( .A(n12337), .ZN(n12341) );
  INV_X1 U13660 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13888) );
  NOR2_X1 U13661 ( .A1(n20038), .A2(n20037), .ZN(n20042) );
  INV_X1 U13662 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n17121) );
  NOR2_X1 U13663 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18122), .ZN(
        n18104) );
  OAI211_X1 U13664 ( .C1(n12717), .C2(n12716), .A(n12872), .B(n12715), .ZN(
        n12881) );
  NAND2_X1 U13665 ( .A1(n16985), .A2(n10144), .ZN(n13259) );
  INV_X1 U13666 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n14940) );
  NAND2_X1 U13667 ( .A1(n10998), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10961) );
  INV_X1 U13668 ( .A(n20350), .ZN(n20338) );
  AND2_X1 U13669 ( .A1(n11515), .A2(n11514), .ZN(n14860) );
  AND2_X1 U13670 ( .A1(n21074), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13810) );
  NAND2_X1 U13671 ( .A1(n11243), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11262) );
  AND3_X1 U13672 ( .A1(n14870), .A2(n14906), .A3(n14920), .ZN(n14907) );
  NAND2_X1 U13673 ( .A1(n10586), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11103) );
  INV_X1 U13674 ( .A(n14653), .ZN(n14654) );
  OR2_X1 U13675 ( .A1(n15400), .A2(n15276), .ZN(n15353) );
  AND2_X1 U13676 ( .A1(n11521), .A2(n11520), .ZN(n14831) );
  AND2_X1 U13677 ( .A1(n15197), .A2(n15196), .ZN(n15212) );
  INV_X1 U13678 ( .A(n15526), .ZN(n21184) );
  OR2_X1 U13679 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20743), .ZN(
        n20734) );
  INV_X1 U13680 ( .A(n20570), .ZN(n20495) );
  INV_X1 U13681 ( .A(n20978), .ZN(n21017) );
  INV_X1 U13682 ( .A(n14012), .ZN(n16874) );
  NOR2_X1 U13683 ( .A1(n20173), .A2(n20166), .ZN(n13916) );
  AND2_X1 U13684 ( .A1(n12299), .A2(n12298), .ZN(n15622) );
  INV_X1 U13685 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15725) );
  NAND2_X1 U13686 ( .A1(n11643), .A2(n11642), .ZN(n11743) );
  AND2_X1 U13687 ( .A1(n12240), .A2(n12239), .ZN(n13934) );
  AND2_X1 U13688 ( .A1(n13626), .A2(n13625), .ZN(n13632) );
  INV_X1 U13689 ( .A(n16138), .ZN(n16161) );
  OR2_X1 U13690 ( .A1(n14410), .A2(n14409), .ZN(n16044) );
  AND2_X1 U13691 ( .A1(n12080), .A2(n12079), .ZN(n13676) );
  AND2_X1 U13692 ( .A1(n16778), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13395) );
  AND2_X1 U13693 ( .A1(n12186), .A2(n12185), .ZN(n15633) );
  NOR2_X1 U13694 ( .A1(n14320), .A2(n14319), .ZN(n14321) );
  AND3_X1 U13695 ( .A1(n12136), .A2(n12135), .A3(n12134), .ZN(n13852) );
  NOR2_X1 U13696 ( .A1(n12341), .A2(n12340), .ZN(n13904) );
  NAND2_X1 U13697 ( .A1(n15573), .A2(n13503), .ZN(n13504) );
  INV_X1 U13698 ( .A(n19409), .ZN(n16750) );
  AND2_X1 U13699 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19628), .ZN(
        n19660) );
  AND2_X1 U13700 ( .A1(n19692), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19726) );
  OR2_X1 U13701 ( .A1(n19923), .A2(n19921), .ZN(n19950) );
  OR2_X1 U13702 ( .A1(n19995), .A2(n19991), .ZN(n20022) );
  AND2_X1 U13703 ( .A1(n20102), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19578) );
  INV_X1 U13704 ( .A(n20072), .ZN(n20138) );
  INV_X1 U13705 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20044) );
  AND2_X1 U13706 ( .A1(n17408), .A2(P3_EBX_REG_29__SCAN_IN), .ZN(n17123) );
  OR2_X1 U13707 ( .A1(n19284), .A2(n17183), .ZN(n12724) );
  INV_X1 U13708 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17361) );
  NAND2_X1 U13709 ( .A1(n19357), .A2(n17424), .ZN(n12731) );
  NOR2_X1 U13710 ( .A1(n13284), .A2(n17121), .ZN(n13285) );
  NOR2_X1 U13711 ( .A1(n18528), .A2(n18196), .ZN(n18507) );
  NOR2_X1 U13712 ( .A1(n17902), .A2(n12893), .ZN(n12912) );
  NAND2_X1 U13713 ( .A1(n19371), .A2(n14234), .ZN(n19177) );
  NOR2_X1 U13714 ( .A1(n12637), .A2(n12636), .ZN(n18721) );
  OR2_X1 U13715 ( .A1(n11157), .A2(n14940), .ZN(n11159) );
  INV_X1 U13716 ( .A(n20354), .ZN(n20327) );
  AND2_X1 U13717 ( .A1(n14025), .A2(n14019), .ZN(n20367) );
  NOR2_X1 U13718 ( .A1(n20396), .A2(n11559), .ZN(n11560) );
  INV_X1 U13719 ( .A(n20396), .ZN(n14968) );
  NAND2_X1 U13720 ( .A1(n11457), .A2(n11456), .ZN(n13306) );
  INV_X1 U13721 ( .A(n13553), .ZN(n20439) );
  NOR2_X1 U13722 ( .A1(n14169), .A2(n14168), .ZN(n20387) );
  INV_X1 U13723 ( .A(n20293), .ZN(n16926) );
  AND2_X1 U13724 ( .A1(n15328), .A2(n15279), .ZN(n15318) );
  NOR2_X1 U13725 ( .A1(n16968), .A2(n16945), .ZN(n16956) );
  INV_X1 U13726 ( .A(n15493), .ZN(n20458) );
  INV_X1 U13727 ( .A(n20481), .ZN(n16965) );
  NOR2_X1 U13728 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16985) );
  AND2_X1 U13729 ( .A1(n16880), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13718) );
  OAI211_X1 U13730 ( .C1(n20534), .C2(n20782), .A(n20842), .B(n20500), .ZN(
        n20537) );
  OAI22_X1 U13731 ( .A1(n20577), .A2(n20576), .B1(n20704), .B2(n20777), .ZN(
        n20601) );
  OAI22_X1 U13732 ( .A1(n20616), .A2(n20615), .B1(n21074), .B2(n20614), .ZN(
        n20639) );
  INV_X1 U13733 ( .A(n20663), .ZN(n20668) );
  OR2_X1 U13734 ( .A1(n15553), .A2(n20495), .ZN(n20900) );
  OR2_X1 U13735 ( .A1(n15553), .A2(n20570), .ZN(n20809) );
  INV_X1 U13736 ( .A(n20871), .ZN(n20749) );
  INV_X1 U13737 ( .A(n20772), .ZN(n20799) );
  AND2_X1 U13738 ( .A1(n20872), .A2(n20932), .ZN(n20865) );
  AND2_X1 U13739 ( .A1(n20875), .A2(n20981), .ZN(n20837) );
  OAI22_X1 U13740 ( .A1(n20911), .A2(n20910), .B1(n20976), .B2(n20909), .ZN(
        n20927) );
  NOR2_X2 U13741 ( .A1(n21017), .A2(n20900), .ZN(n20970) );
  INV_X1 U13742 ( .A(n21069), .ZN(n21003) );
  AND2_X1 U13743 ( .A1(n21185), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16880) );
  INV_X1 U13744 ( .A(n21175), .ZN(n21075) );
  INV_X1 U13745 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21092) );
  INV_X1 U13746 ( .A(n21141), .ZN(n21144) );
  AND2_X1 U13747 ( .A1(n14058), .A2(n14059), .ZN(n15573) );
  INV_X1 U13748 ( .A(n15936), .ZN(n13130) );
  AND2_X1 U13749 ( .A1(n13048), .A2(n13047), .ZN(n19406) );
  INV_X1 U13750 ( .A(n15955), .ZN(n19414) );
  OR2_X1 U13751 ( .A1(n12132), .A2(n12131), .ZN(n14185) );
  INV_X1 U13752 ( .A(n16061), .ZN(n16036) );
  AND2_X1 U13753 ( .A1(n12039), .A2(n12038), .ZN(n14076) );
  NAND2_X1 U13754 ( .A1(n14059), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13630) );
  AND3_X1 U13755 ( .A1(n11823), .A2(n13910), .A3(n13045), .ZN(n13348) );
  AOI21_X1 U13756 ( .B1(n15619), .B2(n10023), .A(n13023), .ZN(n13024) );
  INV_X1 U13757 ( .A(n16439), .ZN(n16426) );
  INV_X1 U13758 ( .A(n11853), .ZN(n11856) );
  AND2_X1 U13759 ( .A1(n14318), .A2(n13656), .ZN(n16729) );
  INV_X1 U13760 ( .A(n16708), .ZN(n16724) );
  NAND2_X1 U13761 ( .A1(n19532), .A2(n19531), .ZN(n19582) );
  AND2_X1 U13762 ( .A1(n20264), .A2(n19523), .ZN(n19820) );
  OAI21_X1 U13763 ( .B1(n19664), .B2(n19663), .A(n19662), .ZN(n19685) );
  AND2_X1 U13764 ( .A1(n19792), .A2(n20252), .ZN(n19719) );
  OAI21_X1 U13765 ( .B1(n19730), .B2(n19729), .A(n19728), .ZN(n19748) );
  AND2_X1 U13766 ( .A1(n19792), .A2(n19723), .ZN(n19780) );
  INV_X1 U13767 ( .A(n19854), .ZN(n19815) );
  NAND2_X1 U13768 ( .A1(n19830), .A2(n19829), .ZN(n19850) );
  INV_X1 U13769 ( .A(n19895), .ZN(n19914) );
  AND2_X1 U13770 ( .A1(n20264), .A2(n20254), .ZN(n20252) );
  NOR2_X2 U13771 ( .A1(n19988), .A2(n19657), .ZN(n19983) );
  NOR2_X2 U13772 ( .A1(n20031), .A2(n19993), .ZN(n20025) );
  AND2_X1 U13773 ( .A1(n20102), .A2(n19538), .ZN(n20053) );
  AND2_X1 U13774 ( .A1(n19578), .A2(n12532), .ZN(n20072) );
  OAI22_X1 U13775 ( .A1(n19536), .A2(n19571), .B1(n19535), .B2(n19573), .ZN(
        n20113) );
  OAI22_X1 U13776 ( .A1(n19559), .A2(n19571), .B1(n19558), .B2(n19573), .ZN(
        n20073) );
  NOR2_X2 U13777 ( .A1(n14365), .A2(n16770), .ZN(n19576) );
  INV_X1 U13778 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n21286) );
  NOR2_X1 U13779 ( .A1(n19152), .A2(n17971), .ZN(n19357) );
  NOR2_X1 U13780 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17150), .ZN(n17135) );
  INV_X1 U13781 ( .A(n17153), .ZN(n17142) );
  NOR2_X1 U13782 ( .A1(n17474), .A2(n12724), .ZN(n17169) );
  NOR2_X1 U13783 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17236), .ZN(n17220) );
  NOR2_X1 U13784 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17262), .ZN(n17244) );
  INV_X1 U13785 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18707) );
  NOR2_X1 U13786 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17336), .ZN(n17314) );
  NOR2_X1 U13787 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17343), .ZN(n17342) );
  INV_X1 U13788 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17410) );
  INV_X1 U13789 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17444) );
  INV_X1 U13790 ( .A(n17471), .ZN(n17460) );
  INV_X1 U13791 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17263) );
  INV_X1 U13792 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17697) );
  NOR2_X1 U13793 ( .A1(n17827), .A2(n17853), .ZN(n17843) );
  INV_X1 U13794 ( .A(n18219), .ZN(n18380) );
  INV_X1 U13795 ( .A(n17971), .ZN(n17974) );
  NAND2_X1 U13796 ( .A1(n12927), .A2(n18045), .ZN(n12889) );
  INV_X1 U13797 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18117) );
  INV_X1 U13798 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18298) );
  INV_X1 U13799 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18163) );
  NOR2_X1 U13800 ( .A1(n18562), .A2(n18561), .ZN(n18558) );
  INV_X1 U13801 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18561) );
  INV_X1 U13802 ( .A(n18685), .ZN(n18650) );
  NOR2_X1 U13803 ( .A1(n18450), .A2(n18702), .ZN(n18698) );
  NOR2_X1 U13804 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19335), .ZN(
        n19337) );
  INV_X1 U13805 ( .A(n18824), .ZN(n18817) );
  INV_X1 U13806 ( .A(n18846), .ZN(n18839) );
  INV_X1 U13807 ( .A(n18860), .ZN(n18865) );
  INV_X1 U13808 ( .A(n18892), .ZN(n18885) );
  INV_X1 U13809 ( .A(n18972), .ZN(n18979) );
  INV_X1 U13810 ( .A(n19005), .ZN(n18998) );
  NOR2_X1 U13811 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19196), .ZN(
        n18985) );
  INV_X1 U13812 ( .A(n19089), .ZN(n19080) );
  AND2_X1 U13813 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19036), .ZN(n19134) );
  INV_X1 U13814 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19215) );
  NOR2_X1 U13815 ( .A1(n19368), .A2(n19240), .ZN(n19239) );
  INV_X1 U13816 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20979) );
  AOI21_X1 U13817 ( .B1(n15283), .B2(n20367), .A(n14666), .ZN(n14667) );
  INV_X1 U13818 ( .A(n20367), .ZN(n20325) );
  INV_X1 U13819 ( .A(n20377), .ZN(n20360) );
  OAI211_X2 U13820 ( .C1(n13458), .C2(n13306), .A(n13305), .B(n13553), .ZN(
        n15031) );
  NAND2_X1 U13821 ( .A1(n20408), .A2(n10837), .ZN(n20397) );
  INV_X1 U13822 ( .A(n20408), .ZN(n20428) );
  OR3_X1 U13823 ( .A1(n14007), .A2(n14013), .A3(n21075), .ZN(n13553) );
  NAND2_X1 U13824 ( .A1(n16937), .A2(n13652), .ZN(n16929) );
  OR2_X1 U13825 ( .A1(n13556), .A2(n16864), .ZN(n20293) );
  OR2_X1 U13826 ( .A1(n16969), .A2(n15495), .ZN(n16968) );
  INV_X1 U13827 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20489) );
  OR2_X1 U13828 ( .A1(n20610), .A2(n20900), .ZN(n20563) );
  OR2_X1 U13829 ( .A1(n20610), .A2(n20809), .ZN(n20599) );
  OR2_X1 U13830 ( .A1(n20610), .A2(n20831), .ZN(n20643) );
  OR2_X1 U13831 ( .A1(n20610), .A2(n20749), .ZN(n20663) );
  OR2_X1 U13832 ( .A1(n20750), .A2(n20900), .ZN(n20697) );
  OR2_X1 U13833 ( .A1(n20750), .A2(n20809), .ZN(n20735) );
  OR2_X1 U13834 ( .A1(n20750), .A2(n20831), .ZN(n20765) );
  NAND2_X1 U13835 ( .A1(n20872), .A2(n20773), .ZN(n20829) );
  AOI22_X1 U13836 ( .A1(n20840), .A2(n20837), .B1(n20835), .B2(n20834), .ZN(
        n20870) );
  NAND2_X1 U13837 ( .A1(n20872), .A2(n20871), .ZN(n20931) );
  NAND2_X1 U13838 ( .A1(n20978), .A2(n20932), .ZN(n21007) );
  NAND2_X1 U13839 ( .A1(n20978), .A2(n20977), .ZN(n21069) );
  INV_X2 U13840 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21074) );
  NOR2_X1 U13841 ( .A1(n21172), .A2(n21082), .ZN(n21157) );
  INV_X1 U13842 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21086) );
  OR2_X1 U13843 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21086), .ZN(n21170) );
  OR2_X1 U13844 ( .A1(n13917), .A2(n19381), .ZN(n15576) );
  INV_X1 U13845 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20036) );
  NAND2_X1 U13846 ( .A1(n19489), .A2(n20036), .ZN(n15955) );
  OR2_X1 U13847 ( .A1(n19402), .A2(n20104), .ZN(n19424) );
  AND2_X1 U13848 ( .A1(n13516), .A2(n13532), .ZN(n16058) );
  INV_X1 U13849 ( .A(n20254), .ZN(n19523) );
  OR2_X1 U13850 ( .A1(n16019), .A2(n16018), .ZN(n16110) );
  OR2_X1 U13851 ( .A1(n19431), .A2(n11794), .ZN(n16171) );
  AND2_X1 U13852 ( .A1(n13533), .A2(n13532), .ZN(n16137) );
  AND2_X1 U13853 ( .A1(n16171), .A2(n16165), .ZN(n14084) );
  OR2_X1 U13854 ( .A1(n13630), .A2(n16742), .ZN(n13434) );
  NAND2_X1 U13855 ( .A1(n13394), .A2(n15568), .ZN(n19479) );
  OR2_X1 U13856 ( .A1(n19517), .A2(n19489), .ZN(n13366) );
  AND2_X1 U13857 ( .A1(n16153), .A2(n16152), .ZN(n19497) );
  NAND2_X1 U13858 ( .A1(n13348), .A2(n10064), .ZN(n13392) );
  INV_X1 U13859 ( .A(n19489), .ZN(n19520) );
  NOR2_X1 U13860 ( .A1(n16567), .A2(n14324), .ZN(n14341) );
  NAND2_X1 U13861 ( .A1(n12554), .A2(n20278), .ZN(n16706) );
  INV_X1 U13862 ( .A(n16814), .ZN(n16809) );
  NAND2_X1 U13863 ( .A1(n19820), .A2(n19753), .ZN(n19625) );
  NAND2_X1 U13864 ( .A1(n19753), .A2(n20252), .ZN(n19683) );
  INV_X1 U13865 ( .A(n19747), .ZN(n19745) );
  NAND2_X1 U13866 ( .A1(n20098), .A2(n19753), .ZN(n19819) );
  NAND2_X1 U13867 ( .A1(n19792), .A2(n20098), .ZN(n19854) );
  OR2_X1 U13868 ( .A1(n20031), .A2(n19857), .ZN(n19883) );
  AOI211_X2 U13869 ( .C1(n16769), .C2(n16768), .A(n16767), .B(n19996), .ZN(
        n19987) );
  INV_X1 U13870 ( .A(n20159), .ZN(n20029) );
  INV_X1 U13871 ( .A(n20073), .ZN(n20144) );
  INV_X1 U13872 ( .A(n20250), .ZN(n20165) );
  NAND2_X1 U13873 ( .A1(n20167), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20284) );
  INV_X1 U13874 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19359) );
  INV_X1 U13875 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17340) );
  NAND2_X1 U13876 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n19222), .ZN(n17431) );
  INV_X1 U13877 ( .A(n17766), .ZN(n17760) );
  NAND2_X1 U13878 ( .A1(n17779), .A2(n17826), .ZN(n17766) );
  INV_X1 U13879 ( .A(n17858), .ZN(n17842) );
  NOR2_X1 U13880 ( .A1(n18029), .A2(n17889), .ZN(n17886) );
  NOR2_X1 U13881 ( .A1(n12772), .A2(n12771), .ZN(n17909) );
  NAND2_X1 U13882 ( .A1(n19183), .A2(n16900), .ZN(n17917) );
  OR2_X1 U13883 ( .A1(n19214), .A2(n18380), .ZN(n19354) );
  OR2_X1 U13884 ( .A1(n17971), .A2(n17933), .ZN(n17970) );
  AND2_X1 U13885 ( .A1(n12945), .A2(n12944), .ZN(n12946) );
  NAND2_X1 U13886 ( .A1(n18375), .A2(n13029), .ZN(n18248) );
  INV_X1 U13887 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18347) );
  NAND2_X1 U13888 ( .A1(n12963), .A2(n18403), .ZN(n18567) );
  INV_X1 U13889 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18601) );
  INV_X1 U13890 ( .A(n18698), .ZN(n18677) );
  NAND2_X1 U13891 ( .A1(n18701), .A2(n18702), .ZN(n18685) );
  INV_X1 U13892 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19196) );
  INV_X1 U13893 ( .A(n19096), .ZN(n19039) );
  INV_X1 U13894 ( .A(n19085), .ZN(n19083) );
  INV_X1 U13895 ( .A(n19074), .ZN(n19124) );
  INV_X1 U13896 ( .A(n18978), .ZN(n19149) );
  INV_X1 U13897 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19335) );
  INV_X1 U13898 ( .A(n19310), .ZN(n19223) );
  INV_X1 U13899 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19237) );
  INV_X1 U13900 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19260) );
  NAND2_X1 U13901 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19237), .ZN(n19368) );
  NOR2_X1 U13902 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13339), .ZN(n17085)
         );
  INV_X1 U13903 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20189) );
  OAI21_X1 U13904 ( .B1(n14980), .B2(n14970), .A(n11562), .ZN(P1_U2843) );
  NAND2_X1 U13905 ( .A1(n13291), .A2(n13290), .ZN(P3_U2801) );
  NAND2_X1 U13906 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10997) );
  AND2_X2 U13907 ( .A1(n11042), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11082) );
  INV_X1 U13908 ( .A(n11103), .ZN(n10587) );
  NAND2_X1 U13909 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10588) );
  NOR2_X2 U13910 ( .A1(n11159), .A2(n10588), .ZN(n11137) );
  NAND2_X1 U13911 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10590) );
  INV_X1 U13912 ( .A(n11350), .ZN(n10594) );
  INV_X1 U13913 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15056) );
  INV_X1 U13914 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10595) );
  NAND2_X1 U13915 ( .A1(n10596), .A2(n10595), .ZN(n10597) );
  NAND2_X1 U13916 ( .A1(n14003), .A2(n10597), .ZN(n15052) );
  INV_X1 U13918 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10599) );
  AND2_X2 U13919 ( .A1(n10599), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10607) );
  AND2_X2 U13921 ( .A1(n10606), .A2(n13457), .ZN(n10768) );
  BUF_X4 U13922 ( .A(n10768), .Z(n11309) );
  AOI22_X1 U13923 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11309), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10604) );
  AND2_X2 U13924 ( .A1(n15518), .A2(n13485), .ZN(n10791) );
  AOI22_X1 U13925 ( .A1(n13139), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U13926 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10883), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10602) );
  INV_X1 U13927 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10600) );
  AOI22_X1 U13928 ( .A1(n10667), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9608), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10601) );
  NAND4_X1 U13929 ( .A1(n10604), .A2(n10603), .A3(n10602), .A4(n10601), .ZN(
        n10613) );
  AOI22_X1 U13930 ( .A1(n13149), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13141), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10611) );
  AND2_X2 U13931 ( .A1(n13485), .A2(n15519), .ZN(n10804) );
  AOI22_X1 U13932 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10610) );
  AND2_X2 U13933 ( .A1(n10606), .A2(n10607), .ZN(n10759) );
  AOI22_X1 U13934 ( .A1(n13138), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10609) );
  AND2_X2 U13935 ( .A1(n10607), .A2(n15519), .ZN(n10700) );
  AND2_X4 U13936 ( .A1(n13457), .A2(n15519), .ZN(n13148) );
  AOI22_X1 U13937 ( .A1(n11246), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10608) );
  NAND4_X1 U13938 ( .A1(n10611), .A2(n10610), .A3(n10609), .A4(n10608), .ZN(
        n10612) );
  NOR2_X1 U13939 ( .A1(n10613), .A2(n10612), .ZN(n11363) );
  AOI22_X1 U13940 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10617) );
  AOI22_X1 U13941 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10616) );
  AOI22_X1 U13942 ( .A1(n10799), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10883), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U13943 ( .A1(n13138), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10614) );
  NAND4_X1 U13944 ( .A1(n10617), .A2(n10616), .A3(n10615), .A4(n10614), .ZN(
        n10623) );
  AOI22_X1 U13945 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10667), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10621) );
  AOI22_X1 U13946 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11309), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U13947 ( .A1(n11246), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9608), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13948 ( .A1(n13149), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10618) );
  NAND4_X1 U13949 ( .A1(n10621), .A2(n10620), .A3(n10619), .A4(n10618), .ZN(
        n10622) );
  NOR2_X1 U13950 ( .A1(n10623), .A2(n10622), .ZN(n11344) );
  AOI22_X1 U13951 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n9593), .B1(
        n10667), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10629) );
  AOI22_X1 U13952 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10628) );
  BUF_X4 U13953 ( .A(n10759), .Z(n11302) );
  AOI22_X1 U13954 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n11302), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10627) );
  AOI22_X1 U13955 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11310), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10626) );
  NAND4_X1 U13956 ( .A1(n10629), .A2(n10628), .A3(n10627), .A4(n10626), .ZN(
        n10635) );
  AOI22_X1 U13957 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n11268), .B1(
        n11309), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10633) );
  BUF_X1 U13958 ( .A(n10672), .Z(n13141) );
  AOI22_X1 U13959 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13141), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10632) );
  AOI22_X1 U13960 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10631) );
  AOI22_X1 U13961 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10630) );
  NAND4_X1 U13962 ( .A1(n10633), .A2(n10632), .A3(n10631), .A4(n10630), .ZN(
        n10634) );
  NOR2_X1 U13963 ( .A1(n10635), .A2(n10634), .ZN(n11327) );
  AOI22_X1 U13964 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13139), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10639) );
  AOI22_X1 U13965 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10638) );
  BUF_X4 U13966 ( .A(n10768), .Z(n15522) );
  AOI22_X1 U13967 ( .A1(n15522), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10883), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10637) );
  AOI22_X1 U13968 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10636) );
  NAND4_X1 U13969 ( .A1(n10639), .A2(n10638), .A3(n10637), .A4(n10636), .ZN(
        n10645) );
  AOI22_X1 U13970 ( .A1(n10667), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10643) );
  AOI22_X1 U13971 ( .A1(n11268), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13141), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10642) );
  AOI22_X1 U13972 ( .A1(n11302), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10641) );
  AOI22_X1 U13973 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10640) );
  NAND4_X1 U13974 ( .A1(n10643), .A2(n10642), .A3(n10641), .A4(n10640), .ZN(
        n10644) );
  NOR2_X1 U13975 ( .A1(n10645), .A2(n10644), .ZN(n11326) );
  NOR2_X1 U13976 ( .A1(n11327), .A2(n11326), .ZN(n11335) );
  AOI22_X1 U13977 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10667), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10650) );
  AOI22_X1 U13978 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10649) );
  AOI22_X1 U13979 ( .A1(n11302), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U13980 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10647) );
  NAND4_X1 U13981 ( .A1(n10650), .A2(n10649), .A3(n10648), .A4(n10647), .ZN(
        n10656) );
  AOI22_X1 U13982 ( .A1(n11268), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15522), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10654) );
  AOI22_X1 U13983 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13984 ( .A1(n10799), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10883), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U13985 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10651) );
  NAND4_X1 U13986 ( .A1(n10654), .A2(n10653), .A3(n10652), .A4(n10651), .ZN(
        n10655) );
  OR2_X1 U13987 ( .A1(n10656), .A2(n10655), .ZN(n11336) );
  NAND2_X1 U13988 ( .A1(n11335), .A2(n11336), .ZN(n11345) );
  NOR2_X1 U13989 ( .A1(n11344), .A2(n11345), .ZN(n11351) );
  AOI22_X1 U13990 ( .A1(n13149), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11309), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10660) );
  AOI22_X1 U13991 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13140), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10659) );
  AOI22_X1 U13992 ( .A1(n10799), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U13993 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10657) );
  NAND4_X1 U13994 ( .A1(n10660), .A2(n10659), .A3(n10658), .A4(n10657), .ZN(
        n10666) );
  AOI22_X1 U13995 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10667), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U13996 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10663) );
  AOI22_X1 U13997 ( .A1(n11302), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10662) );
  AOI22_X1 U13998 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10661) );
  NAND4_X1 U13999 ( .A1(n10664), .A2(n10663), .A3(n10662), .A4(n10661), .ZN(
        n10665) );
  OR2_X1 U14000 ( .A1(n10666), .A2(n10665), .ZN(n11352) );
  NAND2_X1 U14001 ( .A1(n11351), .A2(n11352), .ZN(n11362) );
  NOR2_X1 U14002 ( .A1(n11363), .A2(n11362), .ZN(n11375) );
  AOI22_X1 U14003 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10667), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U14004 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10670) );
  AOI22_X1 U14005 ( .A1(n13138), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10669) );
  AOI22_X1 U14006 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10668) );
  NAND4_X1 U14007 ( .A1(n10671), .A2(n10670), .A3(n10669), .A4(n10668), .ZN(
        n10678) );
  AOI22_X1 U14008 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15522), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10676) );
  AOI22_X1 U14009 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13140), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10675) );
  BUF_X2 U14010 ( .A(n10672), .Z(n11304) );
  AOI22_X1 U14011 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10674) );
  AOI22_X1 U14012 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10673) );
  NAND4_X1 U14013 ( .A1(n10676), .A2(n10675), .A3(n10674), .A4(n10673), .ZN(
        n10677) );
  OR2_X1 U14014 ( .A1(n10678), .A2(n10677), .ZN(n11376) );
  NAND2_X1 U14015 ( .A1(n11375), .A2(n11376), .ZN(n13136) );
  AOI22_X1 U14016 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11302), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U14017 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U14018 ( .A1(n10791), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13140), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U14019 ( .A1(n10799), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10679) );
  NAND4_X1 U14020 ( .A1(n10682), .A2(n10681), .A3(n10680), .A4(n10679), .ZN(
        n10689) );
  AOI22_X1 U14021 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13146), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U14022 ( .A1(n11309), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11280), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U14023 ( .A1(n10667), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10700), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10685) );
  AOI22_X1 U14024 ( .A1(n13149), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10684) );
  NAND4_X1 U14025 ( .A1(n10687), .A2(n10686), .A3(n10685), .A4(n10684), .ZN(
        n10688) );
  NOR2_X1 U14026 ( .A1(n10689), .A2(n10688), .ZN(n13137) );
  XNOR2_X1 U14027 ( .A(n13136), .B(n13137), .ZN(n10745) );
  AOI22_X1 U14028 ( .A1(n10699), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10700), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U14029 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10732), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U14030 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9619), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U14031 ( .A1(n13138), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13140), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U14032 ( .A1(n10625), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10624), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10697) );
  AOI22_X1 U14033 ( .A1(n10683), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10791), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10696) );
  AOI22_X1 U14034 ( .A1(n10799), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10883), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10695) );
  AOI22_X1 U14035 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U14036 ( .A1(n10624), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10699), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10704) );
  AOI22_X1 U14037 ( .A1(n10625), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10700), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U14038 ( .A1(n13138), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10791), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10702) );
  NAND4_X1 U14039 ( .A1(n10704), .A2(n10703), .A3(n10702), .A4(n10701), .ZN(
        n10711) );
  AOI22_X1 U14040 ( .A1(n10705), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10768), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10709) );
  AOI22_X1 U14041 ( .A1(n10683), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10804), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10708) );
  AOI22_X1 U14042 ( .A1(n10799), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10883), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10707) );
  AOI22_X1 U14043 ( .A1(n10732), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10706) );
  NAND4_X1 U14044 ( .A1(n10709), .A2(n10708), .A3(n10707), .A4(n10706), .ZN(
        n10710) );
  OR2_X2 U14045 ( .A1(n10711), .A2(n10710), .ZN(n10823) );
  NAND2_X1 U14046 ( .A1(n13149), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10714) );
  NAND2_X1 U14047 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10713) );
  NAND2_X1 U14048 ( .A1(n13138), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10712) );
  NAND3_X1 U14049 ( .A1(n10714), .A2(n10713), .A3(n10712), .ZN(n10715) );
  NAND2_X1 U14050 ( .A1(n10625), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10719) );
  NAND2_X1 U14051 ( .A1(n10699), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10718) );
  NAND2_X1 U14052 ( .A1(n10799), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10717) );
  NAND2_X1 U14053 ( .A1(n10883), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10716) );
  NAND2_X1 U14054 ( .A1(n10683), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10723) );
  NAND2_X1 U14055 ( .A1(n10732), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10722) );
  NAND2_X1 U14056 ( .A1(n10791), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10721) );
  NAND2_X1 U14057 ( .A1(n11310), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10720) );
  NAND2_X1 U14058 ( .A1(n10624), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10727) );
  NAND2_X1 U14059 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10726) );
  NAND2_X1 U14060 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10725) );
  NAND2_X1 U14061 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10724) );
  AOI22_X1 U14062 ( .A1(n10625), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10624), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10736) );
  AOI22_X1 U14063 ( .A1(n15522), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10732), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10735) );
  AOI22_X1 U14064 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11304), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U14065 ( .A1(n13138), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13140), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10733) );
  NAND4_X1 U14066 ( .A1(n10736), .A2(n10735), .A3(n10734), .A4(n10733), .ZN(
        n10742) );
  AOI22_X1 U14067 ( .A1(n10699), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10700), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10740) );
  AOI22_X1 U14068 ( .A1(n10683), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10791), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10739) );
  AOI22_X1 U14069 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9619), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10738) );
  AOI22_X1 U14070 ( .A1(n10883), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10737) );
  NAND4_X1 U14071 ( .A1(n10740), .A2(n10739), .A3(n10738), .A4(n10737), .ZN(
        n10741) );
  OAI21_X1 U14072 ( .B1(n20979), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n21074), .ZN(n10744) );
  NAND2_X1 U14073 ( .A1(n11374), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n10743) );
  OAI211_X1 U14074 ( .C1(n10745), .C2(n11364), .A(n10744), .B(n10743), .ZN(
        n10746) );
  OAI21_X1 U14075 ( .B1(n15052), .B2(n11371), .A(n10746), .ZN(n11382) );
  NAND2_X1 U14076 ( .A1(n10683), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10750) );
  NAND2_X1 U14077 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10749) );
  NAND2_X1 U14078 ( .A1(n11310), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10748) );
  NAND2_X1 U14079 ( .A1(n10883), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10747) );
  AND4_X2 U14080 ( .A1(n10750), .A2(n10749), .A3(n10748), .A4(n10747), .ZN(
        n10767) );
  NAND2_X1 U14081 ( .A1(n10624), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10754) );
  NAND2_X1 U14082 ( .A1(n10625), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10753) );
  NAND2_X1 U14083 ( .A1(n10699), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10752) );
  NAND2_X1 U14084 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10751) );
  NAND2_X1 U14085 ( .A1(n13149), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10758) );
  NAND2_X1 U14086 ( .A1(n10732), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10757) );
  NAND2_X1 U14087 ( .A1(n10799), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10756) );
  NAND2_X1 U14088 ( .A1(n13148), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10755) );
  AND4_X2 U14089 ( .A1(n10758), .A2(n10757), .A3(n10756), .A4(n10755), .ZN(
        n10765) );
  NAND2_X1 U14090 ( .A1(n10759), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10763) );
  NAND2_X1 U14091 ( .A1(n10791), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10762) );
  NAND2_X1 U14092 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10761) );
  NAND2_X1 U14093 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10760) );
  AOI22_X1 U14094 ( .A1(n11268), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10768), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U14095 ( .A1(n10683), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13140), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10771) );
  AOI22_X1 U14096 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10883), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10770) );
  AOI22_X1 U14097 ( .A1(n10732), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10769) );
  AOI22_X1 U14098 ( .A1(n10624), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10699), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U14099 ( .A1(n10625), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10700), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10776) );
  AOI22_X1 U14100 ( .A1(n13138), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10791), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10775) );
  AOI22_X1 U14101 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9619), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10774) );
  AND2_X4 U14103 ( .A1(n10813), .A2(n11438), .ZN(n14671) );
  NAND2_X1 U14104 ( .A1(n13148), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10782) );
  NAND2_X1 U14105 ( .A1(n11310), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10781) );
  NAND2_X1 U14106 ( .A1(n10683), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10780) );
  NAND2_X1 U14107 ( .A1(n10732), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10779) );
  NAND2_X1 U14108 ( .A1(n10768), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10786) );
  NAND2_X1 U14109 ( .A1(n13149), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10785) );
  NAND2_X1 U14110 ( .A1(n10799), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10784) );
  NAND2_X1 U14111 ( .A1(n10883), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10783) );
  NAND2_X1 U14112 ( .A1(n10624), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10790) );
  NAND2_X1 U14113 ( .A1(n10699), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10789) );
  NAND2_X1 U14114 ( .A1(n9619), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10788) );
  NAND2_X1 U14115 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10787) );
  NAND2_X1 U14116 ( .A1(n10625), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10795) );
  NAND2_X1 U14117 ( .A1(n13138), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10794) );
  NAND2_X1 U14118 ( .A1(n10700), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10793) );
  NAND2_X1 U14119 ( .A1(n10791), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10792) );
  AND4_X4 U14120 ( .A1(n9671), .A2(n10798), .A3(n10797), .A4(n10796), .ZN(
        n14010) );
  AOI22_X1 U14121 ( .A1(n10683), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11309), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U14122 ( .A1(n10699), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10799), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10802) );
  AOI22_X1 U14123 ( .A1(n10624), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10791), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10801) );
  AOI22_X1 U14124 ( .A1(n10625), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10800) );
  NAND4_X1 U14125 ( .A1(n10803), .A2(n10802), .A3(n10801), .A4(n10800), .ZN(
        n10810) );
  AOI22_X1 U14126 ( .A1(n11302), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10700), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U14127 ( .A1(n10732), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10804), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U14128 ( .A1(n11268), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10883), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U14129 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9619), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10805) );
  NAND4_X1 U14130 ( .A1(n10808), .A2(n10807), .A3(n10806), .A4(n10805), .ZN(
        n10809) );
  OR2_X2 U14131 ( .A1(n10810), .A2(n10809), .ZN(n20512) );
  NAND2_X1 U14132 ( .A1(n10837), .A2(n20512), .ZN(n10811) );
  AND2_X2 U14133 ( .A1(n14013), .A2(n10812), .ZN(n10847) );
  NAND2_X1 U14134 ( .A1(n14010), .A2(n10813), .ZN(n14026) );
  INV_X1 U14135 ( .A(n14026), .ZN(n10814) );
  AOI21_X2 U14136 ( .B1(n10847), .B2(n20520), .A(n10814), .ZN(n10848) );
  NOR2_X2 U14137 ( .A1(n20512), .A2(n11438), .ZN(n11458) );
  INV_X1 U14138 ( .A(n11458), .ZN(n10817) );
  INV_X1 U14139 ( .A(n11438), .ZN(n10815) );
  AND2_X1 U14140 ( .A1(n10815), .A2(n20512), .ZN(n10816) );
  NAND4_X1 U14141 ( .A1(n10851), .A2(n10848), .A3(n10817), .A4(n13454), .ZN(
        n10822) );
  NAND2_X1 U14142 ( .A1(n10838), .A2(n10818), .ZN(n11455) );
  NOR2_X1 U14143 ( .A1(n10822), .A2(n10821), .ZN(n10834) );
  OAI21_X1 U14144 ( .B1(n10825), .B2(n20512), .A(n10824), .ZN(n10827) );
  NOR2_X1 U14145 ( .A1(n10827), .A2(n10830), .ZN(n10829) );
  NAND2_X1 U14146 ( .A1(n10842), .A2(n14010), .ZN(n10833) );
  INV_X1 U14147 ( .A(n13467), .ZN(n10831) );
  XNOR2_X1 U14148 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n10840) );
  INV_X1 U14149 ( .A(n10840), .ZN(n13346) );
  NAND2_X1 U14150 ( .A1(n10831), .A2(n10556), .ZN(n10832) );
  NAND2_X1 U14151 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10860) );
  OAI21_X1 U14152 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n10860), .ZN(n20833) );
  INV_X1 U14153 ( .A(n16880), .ZN(n10835) );
  INV_X1 U14154 ( .A(n13318), .ZN(n13708) );
  NAND2_X1 U14155 ( .A1(n13708), .A2(n10838), .ZN(n10839) );
  NAND2_X1 U14156 ( .A1(n11458), .A2(n14008), .ZN(n13458) );
  MUX2_X1 U14157 ( .A(n13259), .B(n16880), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n10841) );
  NAND3_X1 U14158 ( .A1(n13746), .A2(n14647), .A3(n20516), .ZN(n10844) );
  NAND2_X1 U14159 ( .A1(n10842), .A2(n10844), .ZN(n10857) );
  NAND3_X1 U14160 ( .A1(n10845), .A2(n13254), .A3(n20508), .ZN(n10856) );
  INV_X1 U14161 ( .A(n10848), .ZN(n10849) );
  NOR2_X1 U14162 ( .A1(n10850), .A2(n10849), .ZN(n10855) );
  INV_X1 U14163 ( .A(n10851), .ZN(n10853) );
  NAND2_X1 U14164 ( .A1(n11458), .A2(n10983), .ZN(n11449) );
  NAND3_X1 U14165 ( .A1(n11449), .A2(n16985), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10852) );
  NOR2_X1 U14166 ( .A1(n10853), .A2(n10852), .ZN(n10854) );
  NAND4_X1 U14167 ( .A1(n10857), .A2(n10856), .A3(n10855), .A4(n10854), .ZN(
        n10894) );
  INV_X1 U14168 ( .A(n10860), .ZN(n10859) );
  NAND2_X1 U14169 ( .A1(n10859), .A2(n20836), .ZN(n20874) );
  NAND2_X1 U14170 ( .A1(n10860), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10861) );
  NAND2_X1 U14171 ( .A1(n20874), .A2(n10861), .ZN(n20503) );
  INV_X1 U14172 ( .A(n13259), .ZN(n10862) );
  NAND2_X1 U14173 ( .A1(n10879), .A2(n10865), .ZN(n10866) );
  INV_X1 U14174 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n21304) );
  AOI22_X1 U14175 ( .A1(n13139), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10699), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U14176 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U14177 ( .A1(n11302), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U14178 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10867) );
  NAND4_X1 U14179 ( .A1(n10870), .A2(n10869), .A3(n10868), .A4(n10867), .ZN(
        n10876) );
  AOI22_X1 U14180 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11309), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10874) );
  AOI22_X1 U14181 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13140), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U14182 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10872) );
  AOI22_X1 U14183 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10871) );
  NAND4_X1 U14184 ( .A1(n10874), .A2(n10873), .A3(n10872), .A4(n10871), .ZN(
        n10875) );
  INV_X1 U14185 ( .A(n10936), .ZN(n10924) );
  AOI22_X1 U14186 ( .A1(n10924), .A2(n10877), .B1(n11398), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10878) );
  INV_X1 U14187 ( .A(n20607), .ZN(n10882) );
  INV_X1 U14188 ( .A(n10937), .ZN(n10907) );
  AOI22_X1 U14189 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13139), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10887) );
  AOI22_X1 U14190 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13149), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10886) );
  AOI22_X1 U14191 ( .A1(n10667), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13141), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10885) );
  AOI22_X1 U14192 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10883), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10884) );
  NAND4_X1 U14193 ( .A1(n10887), .A2(n10886), .A3(n10885), .A4(n10884), .ZN(
        n10893) );
  AOI22_X1 U14194 ( .A1(n11302), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10700), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U14195 ( .A1(n11303), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10890) );
  AOI22_X1 U14196 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10889) );
  AOI22_X1 U14197 ( .A1(n15522), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10888) );
  NAND4_X1 U14198 ( .A1(n10891), .A2(n10890), .A3(n10889), .A4(n10888), .ZN(
        n10892) );
  INV_X1 U14199 ( .A(n10894), .ZN(n10895) );
  AOI22_X1 U14200 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n9593), .B1(
        n10699), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10899) );
  AOI22_X1 U14201 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10700), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U14202 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11302), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U14203 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10896) );
  NAND4_X1 U14204 ( .A1(n10899), .A2(n10898), .A3(n10897), .A4(n10896), .ZN(
        n10905) );
  AOI22_X1 U14205 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n11268), .B1(
        n15522), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10903) );
  AOI22_X1 U14206 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13140), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10902) );
  AOI22_X1 U14207 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n13141), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10901) );
  AOI22_X1 U14208 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10900) );
  NAND4_X1 U14209 ( .A1(n10903), .A2(n10902), .A3(n10901), .A4(n10900), .ZN(
        n10904) );
  NAND2_X1 U14210 ( .A1(n13722), .A2(n13229), .ZN(n10920) );
  INV_X1 U14211 ( .A(n13229), .ZN(n10906) );
  AOI22_X1 U14212 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11302), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U14213 ( .A1(n13139), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10699), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U14214 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U14215 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10908) );
  NAND4_X1 U14216 ( .A1(n10911), .A2(n10910), .A3(n10909), .A4(n10908), .ZN(
        n10917) );
  AOI22_X1 U14217 ( .A1(n11309), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11280), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U14218 ( .A1(n11246), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10914) );
  AOI22_X1 U14219 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13140), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10913) );
  AOI22_X1 U14220 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10912) );
  NAND4_X1 U14221 ( .A1(n10915), .A2(n10914), .A3(n10913), .A4(n10912), .ZN(
        n10916) );
  MUX2_X1 U14222 ( .A(n13164), .B(n10923), .S(n13182), .Z(n10918) );
  INV_X1 U14223 ( .A(n13164), .ZN(n10919) );
  INV_X1 U14224 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10922) );
  AOI21_X1 U14225 ( .B1(n14010), .B2(n13182), .A(n10144), .ZN(n10921) );
  INV_X1 U14226 ( .A(n10923), .ZN(n10927) );
  NAND2_X1 U14227 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10926) );
  NAND2_X1 U14228 ( .A1(n10924), .A2(n13183), .ZN(n10925) );
  INV_X1 U14229 ( .A(n10928), .ZN(n10929) );
  NOR3_X1 U14230 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20836), .A3(
        n20901), .ZN(n20748) );
  NAND2_X1 U14231 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20748), .ZN(
        n20741) );
  NAND2_X1 U14232 ( .A1(n20873), .A2(n20741), .ZN(n10932) );
  NAND3_X1 U14233 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21015) );
  INV_X1 U14234 ( .A(n21015), .ZN(n10931) );
  NAND2_X1 U14235 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10931), .ZN(
        n21009) );
  NAND2_X1 U14236 ( .A1(n10932), .A2(n21009), .ZN(n20775) );
  OAI22_X1 U14237 ( .A1(n13259), .A2(n20775), .B1(n16880), .B2(n20873), .ZN(
        n10933) );
  INV_X1 U14238 ( .A(n10933), .ZN(n10934) );
  AOI22_X1 U14239 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13146), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U14240 ( .A1(n11309), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11280), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U14241 ( .A1(n10667), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10700), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U14242 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10938) );
  NAND4_X1 U14243 ( .A1(n10941), .A2(n10940), .A3(n10939), .A4(n10938), .ZN(
        n10947) );
  AOI22_X1 U14244 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13138), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10945) );
  AOI22_X1 U14245 ( .A1(n13139), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U14246 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U14247 ( .A1(n11303), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10942) );
  NAND4_X1 U14248 ( .A1(n10945), .A2(n10944), .A3(n10943), .A4(n10942), .ZN(
        n10946) );
  AOI22_X1 U14249 ( .A1(n11432), .A2(n13201), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n11398), .ZN(n10948) );
  AOI22_X1 U14250 ( .A1(n13139), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10699), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10953) );
  AOI22_X1 U14251 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10700), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10952) );
  AOI22_X1 U14252 ( .A1(n11302), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10951) );
  AOI22_X1 U14253 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10950) );
  NAND4_X1 U14254 ( .A1(n10953), .A2(n10952), .A3(n10951), .A4(n10950), .ZN(
        n10959) );
  AOI22_X1 U14255 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11309), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U14256 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10956) );
  AOI22_X1 U14257 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10955) );
  AOI22_X1 U14258 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10954) );
  NAND4_X1 U14259 ( .A1(n10957), .A2(n10956), .A3(n10955), .A4(n10954), .ZN(
        n10958) );
  AOI22_X1 U14260 ( .A1(n11432), .A2(n13172), .B1(
        P1_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n11398), .ZN(n11018) );
  NAND2_X1 U14261 ( .A1(n10960), .A2(n13167), .ZN(n10966) );
  OAI21_X1 U14262 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10998), .A(
        n10961), .ZN(n20359) );
  NAND2_X1 U14263 ( .A1(n13708), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10989) );
  OAI21_X1 U14264 ( .B1(n20979), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n21074), .ZN(n10963) );
  NAND2_X1 U14265 ( .A1(n11374), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n10962) );
  OAI211_X1 U14266 ( .C1(n10989), .C2(n21245), .A(n10963), .B(n10962), .ZN(
        n10964) );
  OAI21_X1 U14267 ( .B1(n11371), .B2(n20359), .A(n10964), .ZN(n10965) );
  NAND2_X1 U14268 ( .A1(n15556), .A2(n14127), .ZN(n10973) );
  INV_X1 U14269 ( .A(n10989), .ZN(n11004) );
  INV_X1 U14270 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n10970) );
  XNOR2_X1 U14271 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14018) );
  AOI21_X1 U14272 ( .B1(n13162), .B2(n14018), .A(n13810), .ZN(n10969) );
  OAI21_X1 U14273 ( .B1(n11368), .B2(n10970), .A(n10969), .ZN(n10971) );
  AOI21_X1 U14274 ( .B1(n11004), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10971), .ZN(n10972) );
  NAND2_X1 U14275 ( .A1(n10973), .A2(n10972), .ZN(n13808) );
  XNOR2_X2 U14276 ( .A(n10976), .B(n10975), .ZN(n15553) );
  NAND2_X1 U14277 ( .A1(n15553), .A2(n14127), .ZN(n10980) );
  INV_X1 U14278 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n10977) );
  INV_X1 U14279 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13949) );
  OAI22_X1 U14280 ( .A1(n11368), .A2(n10977), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13949), .ZN(n10978) );
  AOI21_X1 U14281 ( .B1(n11004), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n10978), .ZN(n10979) );
  NAND2_X1 U14282 ( .A1(n10980), .A2(n10979), .ZN(n13685) );
  NAND2_X1 U14283 ( .A1(n20570), .A2(n10983), .ZN(n10984) );
  NAND2_X1 U14284 ( .A1(n10984), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13511) );
  NAND2_X1 U14285 ( .A1(n21074), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10988) );
  NAND2_X1 U14286 ( .A1(n10986), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n10987) );
  OAI211_X1 U14287 ( .C1(n10989), .C2(n16848), .A(n10988), .B(n10987), .ZN(
        n10990) );
  AOI21_X1 U14288 ( .B1(n20606), .B2(n14127), .A(n10990), .ZN(n13510) );
  OR2_X1 U14289 ( .A1(n13511), .A2(n13510), .ZN(n13513) );
  INV_X1 U14290 ( .A(n13510), .ZN(n10991) );
  OR2_X1 U14291 ( .A1(n10991), .A2(n11371), .ZN(n10992) );
  NAND2_X1 U14292 ( .A1(n13513), .A2(n10992), .ZN(n13684) );
  NAND2_X1 U14293 ( .A1(n13685), .A2(n13684), .ZN(n13811) );
  NAND2_X1 U14294 ( .A1(n13810), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10993) );
  NAND2_X1 U14295 ( .A1(n13811), .A2(n10993), .ZN(n10994) );
  AND2_X2 U14296 ( .A1(n13808), .A2(n10994), .ZN(n13785) );
  INV_X1 U14297 ( .A(n15560), .ZN(n10996) );
  NAND2_X1 U14298 ( .A1(n10996), .A2(n14127), .ZN(n11006) );
  INV_X1 U14299 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n11002) );
  INV_X1 U14300 ( .A(n10997), .ZN(n11000) );
  INV_X1 U14301 ( .A(n10998), .ZN(n10999) );
  OAI21_X1 U14302 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11000), .A(
        n10999), .ZN(n20374) );
  AOI22_X1 U14303 ( .A1(n13162), .A2(n20374), .B1(n13810), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11001) );
  OAI21_X1 U14304 ( .B1(n11368), .B2(n11002), .A(n11001), .ZN(n11003) );
  AOI21_X1 U14305 ( .B1(n11004), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11003), .ZN(n11005) );
  AND3_X2 U14306 ( .A1(n13982), .A2(n13785), .A3(n13784), .ZN(n13983) );
  AOI22_X1 U14307 ( .A1(n13139), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10699), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11010) );
  AOI22_X1 U14308 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11009) );
  AOI22_X1 U14309 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11008) );
  AOI22_X1 U14310 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11007) );
  NAND4_X1 U14311 ( .A1(n11010), .A2(n11009), .A3(n11008), .A4(n11007), .ZN(
        n11016) );
  AOI22_X1 U14312 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11286), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11014) );
  AOI22_X1 U14313 ( .A1(n15522), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11013) );
  AOI22_X1 U14314 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11012) );
  AOI22_X1 U14315 ( .A1(n11302), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11011) );
  NAND4_X1 U14316 ( .A1(n11014), .A2(n11013), .A3(n11012), .A4(n11011), .ZN(
        n11015) );
  AOI22_X1 U14317 ( .A1(n11432), .A2(n13215), .B1(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .B2(n11398), .ZN(n11017) );
  NAND2_X1 U14318 ( .A1(n13169), .A2(n11017), .ZN(n11022) );
  INV_X1 U14319 ( .A(n11040), .ZN(n11021) );
  OAI21_X1 U14320 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11023), .A(
        n11043), .ZN(n20344) );
  AOI22_X1 U14321 ( .A1(n11380), .A2(n20344), .B1(n13810), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11024) );
  NAND2_X1 U14322 ( .A1(n13983), .A2(n14068), .ZN(n14066) );
  AOI22_X1 U14323 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10699), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11030) );
  AOI22_X1 U14324 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U14325 ( .A1(n11302), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10791), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11028) );
  AOI22_X1 U14326 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11027) );
  NAND4_X1 U14327 ( .A1(n11030), .A2(n11029), .A3(n11028), .A4(n11027), .ZN(
        n11036) );
  AOI22_X1 U14328 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15522), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11034) );
  AOI22_X1 U14329 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11033) );
  INV_X1 U14330 ( .A(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n21285) );
  AOI22_X1 U14331 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11032) );
  AOI22_X1 U14332 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11031) );
  NAND4_X1 U14333 ( .A1(n11034), .A2(n11033), .A3(n11032), .A4(n11031), .ZN(
        n11035) );
  NAND2_X1 U14334 ( .A1(n11432), .A2(n13224), .ZN(n11038) );
  NAND2_X1 U14335 ( .A1(n11398), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11037) );
  NAND2_X1 U14336 ( .A1(n11038), .A2(n11037), .ZN(n11039) );
  OR2_X1 U14337 ( .A1(n11040), .A2(n11039), .ZN(n11041) );
  NAND2_X1 U14338 ( .A1(n11041), .A2(n13166), .ZN(n13213) );
  INV_X1 U14339 ( .A(n11042), .ZN(n11084) );
  INV_X1 U14340 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11044) );
  NAND2_X1 U14341 ( .A1(n11044), .A2(n11043), .ZN(n11045) );
  NAND2_X1 U14342 ( .A1(n11084), .A2(n11045), .ZN(n20335) );
  AOI22_X1 U14343 ( .A1(n20335), .A2(n13162), .B1(n13810), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11047) );
  NAND2_X1 U14344 ( .A1(n11374), .A2(P1_EAX_REG_6__SCAN_IN), .ZN(n11046) );
  INV_X1 U14345 ( .A(n14125), .ZN(n11048) );
  INV_X1 U14346 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11050) );
  NAND2_X1 U14347 ( .A1(n11432), .A2(n13229), .ZN(n11049) );
  OAI21_X1 U14348 ( .B1(n11416), .B2(n11050), .A(n11049), .ZN(n11051) );
  INV_X1 U14349 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n14165) );
  AOI22_X1 U14350 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11309), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U14351 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13141), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U14352 ( .A1(n11246), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U14353 ( .A1(n13139), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11052) );
  NAND4_X1 U14354 ( .A1(n11055), .A2(n11054), .A3(n11053), .A4(n11052), .ZN(
        n11061) );
  AOI22_X1 U14355 ( .A1(n11302), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10699), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11059) );
  AOI22_X1 U14356 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11058) );
  AOI22_X1 U14357 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11057) );
  AOI22_X1 U14358 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11056) );
  NAND4_X1 U14359 ( .A1(n11059), .A2(n11058), .A3(n11057), .A4(n11056), .ZN(
        n11060) );
  OR2_X1 U14360 ( .A1(n11061), .A2(n11060), .ZN(n11062) );
  NAND2_X1 U14361 ( .A1(n14127), .A2(n11062), .ZN(n11064) );
  XNOR2_X1 U14362 ( .A(n11082), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15252) );
  AOI22_X1 U14363 ( .A1(n15252), .A2(n13162), .B1(n13810), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11063) );
  OAI211_X1 U14364 ( .C1(n11368), .C2(n14165), .A(n11064), .B(n11063), .ZN(
        n14134) );
  AND2_X1 U14365 ( .A1(n14127), .A2(n14134), .ZN(n14130) );
  AOI22_X1 U14366 ( .A1(n13139), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10699), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11068) );
  AOI22_X1 U14367 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11309), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U14368 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U14369 ( .A1(n11310), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11065) );
  NAND4_X1 U14370 ( .A1(n11068), .A2(n11067), .A3(n11066), .A4(n11065), .ZN(
        n11074) );
  AOI22_X1 U14371 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11280), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11072) );
  AOI22_X1 U14372 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11071) );
  AOI22_X1 U14373 ( .A1(n11302), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U14374 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11069) );
  NAND4_X1 U14375 ( .A1(n11072), .A2(n11071), .A3(n11070), .A4(n11069), .ZN(
        n11073) );
  OAI21_X1 U14376 ( .B1(n11074), .B2(n11073), .A(n14127), .ZN(n11079) );
  XNOR2_X1 U14377 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11075), .ZN(
        n20310) );
  INV_X1 U14378 ( .A(n20310), .ZN(n11076) );
  AOI22_X1 U14379 ( .A1(n13810), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n11380), .B2(n11076), .ZN(n11078) );
  NAND2_X1 U14380 ( .A1(n11374), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11077) );
  INV_X1 U14381 ( .A(n15037), .ZN(n11080) );
  AND2_X1 U14382 ( .A1(n14130), .A2(n11080), .ZN(n11081) );
  NAND2_X1 U14383 ( .A1(n14126), .A2(n11081), .ZN(n11092) );
  INV_X1 U14384 ( .A(n14134), .ZN(n11090) );
  INV_X1 U14385 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11088) );
  INV_X1 U14386 ( .A(n11082), .ZN(n11086) );
  INV_X1 U14387 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11083) );
  NAND2_X1 U14388 ( .A1(n11084), .A2(n11083), .ZN(n11085) );
  NAND2_X1 U14389 ( .A1(n11086), .A2(n11085), .ZN(n20319) );
  AOI22_X1 U14390 ( .A1(n20319), .A2(n13162), .B1(n13810), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11087) );
  OAI21_X1 U14391 ( .B1(n11368), .B2(n11088), .A(n11087), .ZN(n11089) );
  INV_X1 U14392 ( .A(n11089), .ZN(n14128) );
  NAND2_X1 U14393 ( .A1(n11092), .A2(n11091), .ZN(n14108) );
  AOI22_X1 U14394 ( .A1(n13139), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11096) );
  AOI22_X1 U14395 ( .A1(n10791), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11095) );
  AOI22_X1 U14396 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11094) );
  AOI22_X1 U14397 ( .A1(n13141), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11093) );
  NAND4_X1 U14398 ( .A1(n11096), .A2(n11095), .A3(n11094), .A4(n11093), .ZN(
        n11102) );
  AOI22_X1 U14399 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10699), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11100) );
  AOI22_X1 U14400 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11302), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11099) );
  AOI22_X1 U14401 ( .A1(n11309), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11280), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U14402 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11097) );
  NAND4_X1 U14403 ( .A1(n11100), .A2(n11099), .A3(n11098), .A4(n11097), .ZN(
        n11101) );
  OAI21_X1 U14404 ( .B1(n11102), .B2(n11101), .A(n14127), .ZN(n11107) );
  XNOR2_X1 U14405 ( .A(n11103), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16911) );
  OR2_X1 U14406 ( .A1(n16911), .A2(n11371), .ZN(n11106) );
  NAND2_X1 U14407 ( .A1(n11374), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11105) );
  NAND2_X1 U14408 ( .A1(n13810), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11104) );
  NAND4_X1 U14409 ( .A1(n11107), .A2(n11106), .A3(n11105), .A4(n11104), .ZN(
        n14111) );
  AOI22_X1 U14410 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11302), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U14411 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15522), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11111) );
  AOI22_X1 U14412 ( .A1(n10667), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11110) );
  AOI22_X1 U14413 ( .A1(n13141), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11109) );
  NAND4_X1 U14414 ( .A1(n11112), .A2(n11111), .A3(n11110), .A4(n11109), .ZN(
        n11118) );
  AOI22_X1 U14415 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11280), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11116) );
  AOI22_X1 U14416 ( .A1(n13139), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11115) );
  AOI22_X1 U14417 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11114) );
  AOI22_X1 U14418 ( .A1(n10791), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11113) );
  NAND4_X1 U14419 ( .A1(n11116), .A2(n11115), .A3(n11114), .A4(n11113), .ZN(
        n11117) );
  NOR2_X1 U14420 ( .A1(n11118), .A2(n11117), .ZN(n11121) );
  NAND2_X1 U14421 ( .A1(n11374), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11120) );
  NAND2_X1 U14422 ( .A1(n13810), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11119) );
  OAI211_X1 U14423 ( .C1(n11189), .C2(n11121), .A(n11120), .B(n11119), .ZN(
        n11122) );
  INV_X1 U14424 ( .A(n11122), .ZN(n11126) );
  INV_X1 U14425 ( .A(n11159), .ZN(n11123) );
  NAND2_X1 U14426 ( .A1(n11123), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11124) );
  INV_X1 U14427 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14914) );
  XNOR2_X1 U14428 ( .A(n11124), .B(n14914), .ZN(n15203) );
  NAND2_X1 U14429 ( .A1(n15203), .A2(n13162), .ZN(n11125) );
  NAND2_X1 U14430 ( .A1(n11126), .A2(n11125), .ZN(n14906) );
  AOI22_X1 U14431 ( .A1(n10667), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11280), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11130) );
  AOI22_X1 U14432 ( .A1(n11309), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13141), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11129) );
  AOI22_X1 U14433 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11128) );
  AOI22_X1 U14434 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11127) );
  NAND4_X1 U14435 ( .A1(n11130), .A2(n11129), .A3(n11128), .A4(n11127), .ZN(
        n11136) );
  AOI22_X1 U14436 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11134) );
  AOI22_X1 U14437 ( .A1(n11302), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11133) );
  AOI22_X1 U14438 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11132) );
  AOI22_X1 U14439 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11131) );
  NAND4_X1 U14440 ( .A1(n11134), .A2(n11133), .A3(n11132), .A4(n11131), .ZN(
        n11135) );
  NOR2_X1 U14441 ( .A1(n11136), .A2(n11135), .ZN(n11142) );
  INV_X1 U14442 ( .A(n11137), .ZN(n11138) );
  INV_X1 U14443 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n14892) );
  XNOR2_X1 U14444 ( .A(n11138), .B(n14892), .ZN(n15191) );
  NAND2_X1 U14445 ( .A1(n15191), .A2(n13162), .ZN(n11141) );
  INV_X1 U14446 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n15025) );
  INV_X1 U14447 ( .A(n13810), .ZN(n11220) );
  OAI22_X1 U14448 ( .A1(n11368), .A2(n15025), .B1(n11220), .B2(n14892), .ZN(
        n11139) );
  INV_X1 U14449 ( .A(n11139), .ZN(n11140) );
  OAI211_X1 U14450 ( .C1(n11142), .C2(n11189), .A(n11141), .B(n11140), .ZN(
        n14884) );
  AOI22_X1 U14451 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11302), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11146) );
  AOI22_X1 U14452 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10667), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11145) );
  AOI22_X1 U14453 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11144) );
  AOI22_X1 U14454 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11143) );
  NAND4_X1 U14455 ( .A1(n11146), .A2(n11145), .A3(n11144), .A4(n11143), .ZN(
        n11152) );
  AOI22_X1 U14456 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13141), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11150) );
  AOI22_X1 U14457 ( .A1(n11309), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11149) );
  AOI22_X1 U14458 ( .A1(n11246), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11148) );
  AOI22_X1 U14459 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11147) );
  NAND4_X1 U14460 ( .A1(n11150), .A2(n11149), .A3(n11148), .A4(n11147), .ZN(
        n11151) );
  NOR2_X1 U14461 ( .A1(n11152), .A2(n11151), .ZN(n11156) );
  INV_X1 U14462 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n15032) );
  INV_X1 U14463 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14922) );
  OAI22_X1 U14464 ( .A1(n11368), .A2(n15032), .B1(n11220), .B2(n14922), .ZN(
        n11153) );
  INV_X1 U14465 ( .A(n11153), .ZN(n11155) );
  XNOR2_X1 U14466 ( .A(n11159), .B(n14922), .ZN(n15208) );
  NAND2_X1 U14467 ( .A1(n15208), .A2(n13162), .ZN(n11154) );
  OAI211_X1 U14468 ( .C1(n11189), .C2(n11156), .A(n11155), .B(n11154), .ZN(
        n14920) );
  NAND2_X1 U14469 ( .A1(n11374), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11161) );
  NAND2_X1 U14470 ( .A1(n11157), .A2(n14940), .ZN(n11158) );
  NAND2_X1 U14471 ( .A1(n11159), .A2(n11158), .ZN(n15223) );
  AOI22_X1 U14472 ( .A1(n15223), .A2(n13162), .B1(n13810), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11160) );
  AOI22_X1 U14473 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11302), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11165) );
  AOI22_X1 U14474 ( .A1(n11268), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13141), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11164) );
  AOI22_X1 U14475 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11163) );
  AOI22_X1 U14476 ( .A1(n11309), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11162) );
  NAND4_X1 U14477 ( .A1(n11165), .A2(n11164), .A3(n11163), .A4(n11162), .ZN(
        n11171) );
  AOI22_X1 U14478 ( .A1(n13139), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10667), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11169) );
  AOI22_X1 U14479 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11168) );
  AOI22_X1 U14480 ( .A1(n11246), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11310), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11167) );
  AOI22_X1 U14481 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11166) );
  NAND4_X1 U14482 ( .A1(n11169), .A2(n11168), .A3(n11167), .A4(n11166), .ZN(
        n11170) );
  OR2_X1 U14483 ( .A1(n11171), .A2(n11170), .ZN(n11172) );
  NAND2_X1 U14484 ( .A1(n14127), .A2(n11172), .ZN(n14932) );
  NAND2_X1 U14485 ( .A1(n14902), .A2(n14932), .ZN(n11173) );
  NAND4_X1 U14486 ( .A1(n14906), .A2(n14884), .A3(n14920), .A4(n11173), .ZN(
        n11191) );
  INV_X1 U14487 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11174) );
  XNOR2_X1 U14488 ( .A(n11175), .B(n11174), .ZN(n15174) );
  AOI22_X1 U14489 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n13146), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11179) );
  AOI22_X1 U14490 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n11281), .B1(
        n11302), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11178) );
  AOI22_X1 U14491 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11280), .B1(
        n13141), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11177) );
  AOI22_X1 U14492 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11176) );
  NAND4_X1 U14493 ( .A1(n11179), .A2(n11178), .A3(n11177), .A4(n11176), .ZN(
        n11185) );
  AOI22_X1 U14494 ( .A1(n13139), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10667), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11183) );
  AOI22_X1 U14495 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10791), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11182) );
  AOI22_X1 U14496 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n11268), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11181) );
  AOI22_X1 U14497 ( .A1(n11309), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11180) );
  NAND4_X1 U14498 ( .A1(n11183), .A2(n11182), .A3(n11181), .A4(n11180), .ZN(
        n11184) );
  NOR2_X1 U14499 ( .A1(n11185), .A2(n11184), .ZN(n11188) );
  NAND2_X1 U14500 ( .A1(n11374), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11187) );
  NAND2_X1 U14501 ( .A1(n13810), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11186) );
  OAI211_X1 U14502 ( .C1(n11189), .C2(n11188), .A(n11187), .B(n11186), .ZN(
        n11190) );
  AOI21_X1 U14503 ( .B1(n15174), .B2(n13162), .A(n11190), .ZN(n14871) );
  XNOR2_X1 U14504 ( .A(n11208), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15170) );
  NAND2_X1 U14505 ( .A1(n15170), .A2(n13162), .ZN(n11207) );
  AOI22_X1 U14506 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11302), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11196) );
  AOI22_X1 U14507 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13149), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11195) );
  AOI22_X1 U14508 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11194) );
  AOI22_X1 U14509 ( .A1(n10791), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11310), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11193) );
  NAND4_X1 U14510 ( .A1(n11196), .A2(n11195), .A3(n11194), .A4(n11193), .ZN(
        n11202) );
  AOI22_X1 U14511 ( .A1(n15522), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11280), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11200) );
  AOI22_X1 U14512 ( .A1(n13141), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11199) );
  AOI22_X1 U14513 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U14514 ( .A1(n10667), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11197) );
  NAND4_X1 U14515 ( .A1(n11200), .A2(n11199), .A3(n11198), .A4(n11197), .ZN(
        n11201) );
  NOR2_X1 U14516 ( .A1(n11202), .A2(n11201), .ZN(n11205) );
  INV_X1 U14517 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15168) );
  AOI21_X1 U14518 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15168), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11203) );
  AOI21_X1 U14519 ( .B1(n11374), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11203), .ZN(
        n11204) );
  OAI21_X1 U14520 ( .B1(n11364), .B2(n11205), .A(n11204), .ZN(n11206) );
  NAND2_X1 U14521 ( .A1(n11207), .A2(n11206), .ZN(n14855) );
  OR2_X1 U14522 ( .A1(n11208), .A2(n15168), .ZN(n11209) );
  INV_X1 U14523 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14846) );
  XNOR2_X1 U14524 ( .A(n11209), .B(n14846), .ZN(n15159) );
  NAND2_X1 U14525 ( .A1(n15159), .A2(n13162), .ZN(n11225) );
  AOI22_X1 U14526 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10667), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11213) );
  AOI22_X1 U14527 ( .A1(n11268), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11309), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14528 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11211) );
  AOI22_X1 U14529 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11310), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11210) );
  NAND4_X1 U14530 ( .A1(n11213), .A2(n11212), .A3(n11211), .A4(n11210), .ZN(
        n11219) );
  AOI22_X1 U14531 ( .A1(n11302), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13141), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11217) );
  AOI22_X1 U14532 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11216) );
  AOI22_X1 U14533 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11215) );
  AOI22_X1 U14534 ( .A1(n13147), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11214) );
  NAND4_X1 U14535 ( .A1(n11217), .A2(n11216), .A3(n11215), .A4(n11214), .ZN(
        n11218) );
  OR2_X1 U14536 ( .A1(n11219), .A2(n11218), .ZN(n11223) );
  INV_X1 U14537 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n11221) );
  OAI22_X1 U14538 ( .A1(n11368), .A2(n11221), .B1(n11220), .B2(n14846), .ZN(
        n11222) );
  AOI21_X1 U14539 ( .B1(n13158), .B2(n11223), .A(n11222), .ZN(n11224) );
  NAND2_X1 U14540 ( .A1(n11225), .A2(n11224), .ZN(n14841) );
  XNOR2_X1 U14541 ( .A(n11226), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15145) );
  NAND2_X1 U14542 ( .A1(n15145), .A2(n11380), .ZN(n11242) );
  AOI22_X1 U14543 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11280), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11231) );
  AOI22_X1 U14544 ( .A1(n11302), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11230) );
  AOI22_X1 U14545 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11229) );
  AOI22_X1 U14546 ( .A1(n10791), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11227), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11228) );
  NAND4_X1 U14547 ( .A1(n11231), .A2(n11230), .A3(n11229), .A4(n11228), .ZN(
        n11237) );
  AOI22_X1 U14548 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10667), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11235) );
  AOI22_X1 U14549 ( .A1(n11268), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11309), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11234) );
  AOI22_X1 U14550 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11233) );
  AOI22_X1 U14551 ( .A1(n13141), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11232) );
  NAND4_X1 U14552 ( .A1(n11235), .A2(n11234), .A3(n11233), .A4(n11232), .ZN(
        n11236) );
  OAI21_X1 U14553 ( .B1(n11237), .B2(n11236), .A(n13158), .ZN(n11240) );
  NAND2_X1 U14554 ( .A1(n11374), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n11239) );
  NAND2_X1 U14555 ( .A1(n21074), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11238) );
  NAND4_X1 U14556 ( .A1(n11240), .A2(n11371), .A3(n11239), .A4(n11238), .ZN(
        n11241) );
  INV_X1 U14557 ( .A(n11243), .ZN(n11244) );
  INV_X1 U14558 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14818) );
  NAND2_X1 U14559 ( .A1(n11244), .A2(n14818), .ZN(n11245) );
  NAND2_X1 U14560 ( .A1(n11262), .A2(n11245), .ZN(n15138) );
  AOI22_X1 U14561 ( .A1(n13139), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10667), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11250) );
  AOI22_X1 U14562 ( .A1(n11302), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11249) );
  AOI22_X1 U14563 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11248) );
  AOI22_X1 U14564 ( .A1(n11310), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11247) );
  NAND4_X1 U14565 ( .A1(n11250), .A2(n11249), .A3(n11248), .A4(n11247), .ZN(
        n11256) );
  AOI22_X1 U14566 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11280), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14567 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15522), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11253) );
  AOI22_X1 U14568 ( .A1(n11268), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11252) );
  AOI22_X1 U14569 ( .A1(n13141), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11251) );
  NAND4_X1 U14570 ( .A1(n11254), .A2(n11253), .A3(n11252), .A4(n11251), .ZN(
        n11255) );
  OAI21_X1 U14571 ( .B1(n11256), .B2(n11255), .A(n13158), .ZN(n11259) );
  NAND2_X1 U14572 ( .A1(n11374), .A2(P1_EAX_REG_19__SCAN_IN), .ZN(n11258) );
  NAND2_X1 U14573 ( .A1(n21074), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11257) );
  NAND4_X1 U14574 ( .A1(n11259), .A2(n11371), .A3(n11258), .A4(n11257), .ZN(
        n11260) );
  NAND2_X1 U14575 ( .A1(n11261), .A2(n11260), .ZN(n14810) );
  XNOR2_X1 U14576 ( .A(n11262), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15127) );
  INV_X1 U14577 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15125) );
  AOI21_X1 U14578 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15125), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11263) );
  AOI21_X1 U14579 ( .B1(n11374), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11263), .ZN(
        n11276) );
  AOI22_X1 U14580 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10667), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11267) );
  AOI22_X1 U14581 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11266) );
  AOI22_X1 U14582 ( .A1(n11302), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11310), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11265) );
  AOI22_X1 U14583 ( .A1(n11280), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11264) );
  NAND4_X1 U14584 ( .A1(n11267), .A2(n11266), .A3(n11265), .A4(n11264), .ZN(
        n11274) );
  AOI22_X1 U14585 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11272) );
  AOI22_X1 U14586 ( .A1(n11246), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13141), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11271) );
  AOI22_X1 U14587 ( .A1(n11309), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11270) );
  AOI22_X1 U14588 ( .A1(n11268), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11269) );
  NAND4_X1 U14589 ( .A1(n11272), .A2(n11271), .A3(n11270), .A4(n11269), .ZN(
        n11273) );
  OAI21_X1 U14590 ( .B1(n11274), .B2(n11273), .A(n13158), .ZN(n11275) );
  AOI22_X1 U14591 ( .A1(n15127), .A2(n13162), .B1(n11276), .B2(n11275), .ZN(
        n14795) );
  INV_X1 U14592 ( .A(n11277), .ZN(n11278) );
  INV_X1 U14593 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15120) );
  NAND2_X1 U14594 ( .A1(n11278), .A2(n15120), .ZN(n11279) );
  NAND2_X1 U14595 ( .A1(n11301), .A2(n11279), .ZN(n15119) );
  AOI22_X1 U14596 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11280), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11285) );
  AOI22_X1 U14597 ( .A1(n11246), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11284) );
  AOI22_X1 U14598 ( .A1(n15522), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11283) );
  AOI22_X1 U14599 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11282) );
  NAND4_X1 U14600 ( .A1(n11285), .A2(n11284), .A3(n11283), .A4(n11282), .ZN(
        n11293) );
  AOI22_X1 U14601 ( .A1(n13139), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11302), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11291) );
  AOI22_X1 U14602 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10667), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11290) );
  AOI22_X1 U14603 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11289) );
  AOI22_X1 U14604 ( .A1(n13141), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11310), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11288) );
  NAND4_X1 U14605 ( .A1(n11291), .A2(n11290), .A3(n11289), .A4(n11288), .ZN(
        n11292) );
  OAI21_X1 U14606 ( .B1(n11293), .B2(n11292), .A(n13158), .ZN(n11296) );
  NAND2_X1 U14607 ( .A1(n11374), .A2(P1_EAX_REG_21__SCAN_IN), .ZN(n11295) );
  NAND2_X1 U14608 ( .A1(n21074), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11294) );
  NAND4_X1 U14609 ( .A1(n11296), .A2(n11371), .A3(n11295), .A4(n11294), .ZN(
        n11297) );
  NAND2_X1 U14610 ( .A1(n11298), .A2(n11297), .ZN(n14787) );
  XNOR2_X1 U14611 ( .A(n11301), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15109) );
  NAND2_X1 U14612 ( .A1(n15109), .A2(n13162), .ZN(n11321) );
  AOI22_X1 U14613 ( .A1(n13146), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13149), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11308) );
  AOI22_X1 U14614 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11302), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11307) );
  AOI22_X1 U14615 ( .A1(n11246), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11303), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11306) );
  AOI22_X1 U14616 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11305) );
  NAND4_X1 U14617 ( .A1(n11308), .A2(n11307), .A3(n11306), .A4(n11305), .ZN(
        n11316) );
  AOI22_X1 U14618 ( .A1(n13139), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10699), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11314) );
  AOI22_X1 U14619 ( .A1(n11309), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11280), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11313) );
  AOI22_X1 U14620 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11312) );
  AOI22_X1 U14621 ( .A1(n11310), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11311) );
  NAND4_X1 U14622 ( .A1(n11314), .A2(n11313), .A3(n11312), .A4(n11311), .ZN(
        n11315) );
  NOR2_X1 U14623 ( .A1(n11316), .A2(n11315), .ZN(n11319) );
  INV_X1 U14624 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15111) );
  AOI21_X1 U14625 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15111), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11317) );
  AOI21_X1 U14626 ( .B1(n11374), .B2(P1_EAX_REG_22__SCAN_IN), .A(n11317), .ZN(
        n11318) );
  OAI21_X1 U14627 ( .B1(n11364), .B2(n11319), .A(n11318), .ZN(n11320) );
  NAND2_X1 U14628 ( .A1(n11321), .A2(n11320), .ZN(n14769) );
  INV_X1 U14629 ( .A(n11322), .ZN(n11324) );
  INV_X1 U14630 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11323) );
  NAND2_X1 U14631 ( .A1(n11324), .A2(n11323), .ZN(n11325) );
  NAND2_X1 U14632 ( .A1(n11333), .A2(n11325), .ZN(n15102) );
  XNOR2_X1 U14633 ( .A(n11327), .B(n11326), .ZN(n11330) );
  OAI21_X1 U14634 ( .B1(n20979), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n21074), .ZN(n11329) );
  NAND2_X1 U14635 ( .A1(n11374), .A2(P1_EAX_REG_23__SCAN_IN), .ZN(n11328) );
  OAI211_X1 U14636 ( .C1(n11330), .C2(n11364), .A(n11329), .B(n11328), .ZN(
        n11331) );
  NAND2_X1 U14637 ( .A1(n11332), .A2(n11331), .ZN(n14753) );
  XNOR2_X1 U14638 ( .A(n11333), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15094) );
  INV_X1 U14639 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15092) );
  NOR2_X1 U14640 ( .A1(n15092), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11334) );
  AOI211_X1 U14641 ( .C1(n11374), .C2(P1_EAX_REG_24__SCAN_IN), .A(n13162), .B(
        n11334), .ZN(n11339) );
  XOR2_X1 U14642 ( .A(n11336), .B(n11335), .Z(n11337) );
  NAND2_X1 U14643 ( .A1(n11337), .A2(n13158), .ZN(n11338) );
  AOI22_X1 U14644 ( .A1(n15094), .A2(n11380), .B1(n11339), .B2(n11338), .ZN(
        n14744) );
  INV_X1 U14645 ( .A(n11340), .ZN(n11342) );
  INV_X1 U14646 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11341) );
  NAND2_X1 U14647 ( .A1(n11342), .A2(n11341), .ZN(n11343) );
  NAND2_X1 U14648 ( .A1(n11350), .A2(n11343), .ZN(n15088) );
  XNOR2_X1 U14649 ( .A(n11345), .B(n11344), .ZN(n11348) );
  OAI21_X1 U14650 ( .B1(n20979), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n21074), .ZN(n11347) );
  NAND2_X1 U14651 ( .A1(n11374), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n11346) );
  OAI211_X1 U14652 ( .C1(n11348), .C2(n11364), .A(n11347), .B(n11346), .ZN(
        n11349) );
  OAI21_X1 U14653 ( .B1(n15088), .B2(n11371), .A(n11349), .ZN(n14732) );
  NOR2_X2 U14654 ( .A1(n14731), .A2(n14732), .ZN(n14718) );
  XNOR2_X1 U14655 ( .A(n11350), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15079) );
  XOR2_X1 U14656 ( .A(n11352), .B(n11351), .Z(n11356) );
  INV_X1 U14657 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n11354) );
  NAND2_X1 U14658 ( .A1(n21074), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11353) );
  OAI211_X1 U14659 ( .C1(n11368), .C2(n11354), .A(n11371), .B(n11353), .ZN(
        n11355) );
  AOI21_X1 U14660 ( .B1(n11356), .B2(n13158), .A(n11355), .ZN(n11357) );
  INV_X1 U14661 ( .A(n11358), .ZN(n11360) );
  INV_X1 U14662 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11359) );
  NAND2_X1 U14663 ( .A1(n11360), .A2(n11359), .ZN(n11361) );
  NAND2_X1 U14664 ( .A1(n11372), .A2(n11361), .ZN(n15073) );
  XNOR2_X1 U14665 ( .A(n11363), .B(n11362), .ZN(n11365) );
  NOR2_X1 U14666 ( .A1(n11365), .A2(n11364), .ZN(n11370) );
  INV_X1 U14667 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n11367) );
  NAND2_X1 U14668 ( .A1(n21074), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11366) );
  OAI211_X1 U14669 ( .C1(n11368), .C2(n11367), .A(n11371), .B(n11366), .ZN(
        n11369) );
  OAI22_X1 U14670 ( .A1(n15073), .A2(n11371), .B1(n11370), .B2(n11369), .ZN(
        n14708) );
  XNOR2_X1 U14671 ( .A(n11372), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15058) );
  NOR2_X1 U14672 ( .A1(n15056), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11373) );
  AOI211_X1 U14673 ( .C1(n11374), .C2(P1_EAX_REG_28__SCAN_IN), .A(n11380), .B(
        n11373), .ZN(n11379) );
  XOR2_X1 U14674 ( .A(n11376), .B(n11375), .Z(n11377) );
  NAND2_X1 U14675 ( .A1(n11377), .A2(n13158), .ZN(n11378) );
  AOI22_X1 U14676 ( .A1(n15058), .A2(n11380), .B1(n11379), .B2(n11378), .ZN(
        n14692) );
  INV_X1 U14677 ( .A(n15054), .ZN(n14980) );
  NAND2_X1 U14678 ( .A1(n14013), .A2(n20524), .ZN(n11383) );
  XNOR2_X1 U14679 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11388) );
  NAND2_X1 U14680 ( .A1(n11392), .A2(n11388), .ZN(n11385) );
  NAND2_X1 U14681 ( .A1(n20901), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11384) );
  NAND2_X1 U14682 ( .A1(n11385), .A2(n11384), .ZN(n11409) );
  XNOR2_X1 U14683 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11408) );
  XNOR2_X1 U14684 ( .A(n11409), .B(n11408), .ZN(n13299) );
  INV_X1 U14685 ( .A(n13299), .ZN(n11404) );
  NAND2_X1 U14686 ( .A1(n11432), .A2(n11404), .ZN(n11406) );
  NAND2_X1 U14687 ( .A1(n11432), .A2(n20508), .ZN(n11387) );
  NAND2_X1 U14688 ( .A1(n10838), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11386) );
  NAND2_X1 U14689 ( .A1(n11387), .A2(n11386), .ZN(n11397) );
  OR2_X1 U14690 ( .A1(n11397), .A2(n14013), .ZN(n11389) );
  XNOR2_X1 U14691 ( .A(n11388), .B(n11392), .ZN(n13297) );
  NAND2_X1 U14692 ( .A1(n11389), .A2(n13297), .ZN(n11403) );
  AND2_X1 U14693 ( .A1(n16848), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11391) );
  NOR2_X1 U14694 ( .A1(n11392), .A2(n11391), .ZN(n11393) );
  OAI211_X1 U14695 ( .C1(n14010), .C2(n11390), .A(n11407), .B(n11393), .ZN(
        n11396) );
  NAND2_X1 U14696 ( .A1(n11432), .A2(n11393), .ZN(n11394) );
  INV_X1 U14697 ( .A(n11397), .ZN(n11400) );
  NAND2_X1 U14698 ( .A1(n11398), .A2(n13297), .ZN(n11399) );
  NAND2_X1 U14699 ( .A1(n11400), .A2(n11399), .ZN(n11401) );
  OAI211_X1 U14700 ( .C1(n11404), .C2(n11416), .A(n11406), .B(n11407), .ZN(
        n11405) );
  NAND2_X1 U14701 ( .A1(n11409), .A2(n11408), .ZN(n11411) );
  NAND2_X1 U14702 ( .A1(n20836), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11410) );
  NAND2_X1 U14703 ( .A1(n11411), .A2(n11410), .ZN(n11423) );
  NAND2_X1 U14704 ( .A1(n15523), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11412) );
  NAND2_X1 U14705 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n21245), .ZN(
        n11426) );
  INV_X1 U14706 ( .A(n11426), .ZN(n11413) );
  NAND2_X1 U14707 ( .A1(n11424), .A2(n11413), .ZN(n11414) );
  NAND2_X1 U14708 ( .A1(n11416), .A2(n13298), .ZN(n11417) );
  NAND2_X1 U14709 ( .A1(n11418), .A2(n11417), .ZN(n11421) );
  AOI22_X1 U14710 ( .A1(n11430), .A2(n13298), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n10144), .ZN(n11420) );
  NAND2_X1 U14711 ( .A1(n11423), .A2(n11422), .ZN(n11425) );
  NAND2_X1 U14712 ( .A1(n11425), .A2(n11424), .ZN(n11427) );
  NAND2_X1 U14713 ( .A1(n11427), .A2(n11426), .ZN(n11429) );
  NAND2_X1 U14714 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20489), .ZN(
        n11428) );
  NAND2_X1 U14715 ( .A1(n11430), .A2(n13301), .ZN(n11431) );
  NAND2_X1 U14716 ( .A1(n10842), .A2(n14008), .ZN(n11447) );
  NAND2_X1 U14717 ( .A1(n11434), .A2(n20508), .ZN(n11452) );
  AND2_X1 U14718 ( .A1(n11452), .A2(n10837), .ZN(n11435) );
  NAND2_X1 U14719 ( .A1(n10845), .A2(n11435), .ZN(n13475) );
  OAI21_X1 U14720 ( .B1(n11437), .B2(n11458), .A(n20508), .ZN(n11441) );
  OR2_X1 U14721 ( .A1(n11438), .A2(n14010), .ZN(n11466) );
  NAND2_X1 U14722 ( .A1(n14652), .A2(n11439), .ZN(n11440) );
  OAI211_X1 U14723 ( .C1(n11442), .C2(n14026), .A(n11441), .B(n11440), .ZN(
        n11443) );
  INV_X1 U14724 ( .A(n11443), .ZN(n11446) );
  NAND2_X1 U14725 ( .A1(n11444), .A2(n14671), .ZN(n11445) );
  NAND4_X1 U14726 ( .A1(n11447), .A2(n13475), .A3(n11446), .A4(n11445), .ZN(
        n13453) );
  MUX2_X1 U14727 ( .A(n11448), .B(n13712), .S(n10837), .Z(n11450) );
  NAND2_X1 U14728 ( .A1(n11450), .A2(n11449), .ZN(n11451) );
  INV_X1 U14729 ( .A(n11452), .ZN(n11453) );
  NOR2_X1 U14730 ( .A1(n13470), .A2(n20288), .ZN(n11454) );
  NAND2_X1 U14731 ( .A1(n16883), .A2(n11454), .ZN(n11461) );
  INV_X1 U14732 ( .A(n20532), .ZN(n14974) );
  AND3_X1 U14733 ( .A1(n14974), .A2(n13722), .A3(n13718), .ZN(n11457) );
  INV_X1 U14734 ( .A(n11455), .ZN(n11456) );
  INV_X1 U14735 ( .A(n13306), .ZN(n11459) );
  NAND3_X1 U14736 ( .A1(n11459), .A2(n11458), .A3(n21355), .ZN(n11460) );
  INV_X2 U14737 ( .A(n20392), .ZN(n14970) );
  INV_X1 U14738 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n21208) );
  NAND2_X1 U14739 ( .A1(n11555), .A2(n21208), .ZN(n11465) );
  INV_X1 U14740 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13727) );
  NAND2_X1 U14741 ( .A1(n11466), .A2(n13727), .ZN(n11462) );
  NAND2_X1 U14742 ( .A1(n11466), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11467) );
  OAI21_X1 U14743 ( .B1(n14671), .B2(P1_EBX_REG_0__SCAN_IN), .A(n11467), .ZN(
        n13509) );
  INV_X1 U14744 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13198) );
  NAND2_X1 U14745 ( .A1(n11466), .A2(n13198), .ZN(n11470) );
  OAI211_X1 U14746 ( .C1(n9614), .C2(P1_EBX_REG_2__SCAN_IN), .A(n11470), .B(
        n14651), .ZN(n11471) );
  OAI21_X1 U14747 ( .B1(n11556), .B2(P1_EBX_REG_2__SCAN_IN), .A(n11471), .ZN(
        n13754) );
  MUX2_X1 U14748 ( .A(n11548), .B(n14671), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n11473) );
  NOR2_X1 U14749 ( .A1(n14652), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11472) );
  NOR2_X1 U14750 ( .A1(n11473), .A2(n11472), .ZN(n13786) );
  INV_X1 U14751 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20395) );
  NAND2_X1 U14752 ( .A1(n11548), .A2(n20395), .ZN(n11476) );
  NAND2_X1 U14753 ( .A1(n14651), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11474) );
  OAI211_X1 U14754 ( .C1(n9613), .C2(P1_EBX_REG_5__SCAN_IN), .A(n11474), .B(
        n11466), .ZN(n11475) );
  NAND2_X1 U14755 ( .A1(n11476), .A2(n11475), .ZN(n16972) );
  INV_X1 U14756 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n11477) );
  NAND2_X1 U14757 ( .A1(n11555), .A2(n11477), .ZN(n11480) );
  INV_X1 U14758 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20461) );
  OAI21_X1 U14759 ( .B1(n14671), .B2(n20461), .A(n11466), .ZN(n11478) );
  OAI21_X1 U14760 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(n9613), .A(n11478), .ZN(
        n11479) );
  INV_X1 U14761 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20389) );
  NAND2_X1 U14762 ( .A1(n11548), .A2(n20389), .ZN(n11485) );
  NAND2_X1 U14763 ( .A1(n14651), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11483) );
  OAI211_X1 U14764 ( .C1(n9613), .C2(P1_EBX_REG_7__SCAN_IN), .A(n11483), .B(
        n11466), .ZN(n11484) );
  AND2_X1 U14765 ( .A1(n11485), .A2(n11484), .ZN(n16952) );
  INV_X1 U14766 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16945) );
  OAI21_X1 U14767 ( .B1(n14671), .B2(n16945), .A(n11466), .ZN(n11486) );
  OAI21_X1 U14768 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(n9613), .A(n11486), .ZN(
        n11487) );
  OAI21_X1 U14769 ( .B1(n11556), .B2(P1_EBX_REG_6__SCAN_IN), .A(n11487), .ZN(
        n16953) );
  NAND2_X1 U14770 ( .A1(n16952), .A2(n16953), .ZN(n11488) );
  INV_X1 U14771 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16951) );
  OAI21_X1 U14772 ( .B1(n14671), .B2(n16951), .A(n11466), .ZN(n11489) );
  OAI21_X1 U14773 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(n9614), .A(n11489), .ZN(
        n11490) );
  OAI21_X1 U14774 ( .B1(n11556), .B2(P1_EBX_REG_8__SCAN_IN), .A(n11490), .ZN(
        n14135) );
  INV_X1 U14775 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20386) );
  NAND2_X1 U14776 ( .A1(n11548), .A2(n20386), .ZN(n11493) );
  NAND2_X1 U14777 ( .A1(n14651), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11491) );
  OAI211_X1 U14778 ( .C1(n9614), .C2(P1_EBX_REG_9__SCAN_IN), .A(n11491), .B(
        n11466), .ZN(n11492) );
  NAND2_X1 U14779 ( .A1(n11493), .A2(n11492), .ZN(n15503) );
  INV_X1 U14780 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14114) );
  NAND2_X1 U14781 ( .A1(n11555), .A2(n14114), .ZN(n11498) );
  INV_X1 U14782 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15227) );
  NAND2_X1 U14783 ( .A1(n11466), .A2(n15227), .ZN(n11496) );
  OAI211_X1 U14784 ( .C1(n9613), .C2(P1_EBX_REG_10__SCAN_IN), .A(n11496), .B(
        n14651), .ZN(n11497) );
  MUX2_X1 U14785 ( .A(n11548), .B(n14671), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n11500) );
  NOR2_X1 U14786 ( .A1(n14652), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11499) );
  NOR2_X1 U14787 ( .A1(n11500), .A2(n11499), .ZN(n14936) );
  MUX2_X1 U14788 ( .A(n11548), .B(n14671), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n11502) );
  NOR2_X1 U14789 ( .A1(n14652), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11501) );
  NOR2_X1 U14790 ( .A1(n11502), .A2(n11501), .ZN(n14910) );
  INV_X1 U14791 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15471) );
  OAI21_X1 U14792 ( .B1(n14671), .B2(n15471), .A(n11466), .ZN(n11503) );
  OAI21_X1 U14793 ( .B1(P1_EBX_REG_12__SCAN_IN), .B2(n9614), .A(n11503), .ZN(
        n11504) );
  OAI21_X1 U14794 ( .B1(n11556), .B2(P1_EBX_REG_12__SCAN_IN), .A(n11504), .ZN(
        n14927) );
  AND2_X1 U14795 ( .A1(n14910), .A2(n14927), .ZN(n11505) );
  INV_X1 U14796 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n11506) );
  NAND2_X1 U14797 ( .A1(n11555), .A2(n11506), .ZN(n11509) );
  INV_X1 U14798 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15444) );
  NAND2_X1 U14799 ( .A1(n11466), .A2(n15444), .ZN(n11507) );
  OAI211_X1 U14800 ( .C1(n9614), .C2(P1_EBX_REG_14__SCAN_IN), .A(n11507), .B(
        n14651), .ZN(n11508) );
  MUX2_X1 U14801 ( .A(n11548), .B(n14671), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n11510) );
  INV_X1 U14802 ( .A(n11510), .ZN(n11512) );
  INV_X1 U14803 ( .A(n14652), .ZN(n11523) );
  INV_X1 U14804 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15429) );
  NAND2_X1 U14805 ( .A1(n11523), .A2(n15429), .ZN(n11511) );
  NAND2_X1 U14806 ( .A1(n11512), .A2(n11511), .ZN(n14873) );
  INV_X1 U14807 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14964) );
  NAND2_X1 U14808 ( .A1(n11555), .A2(n14964), .ZN(n11515) );
  INV_X1 U14809 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15427) );
  NAND2_X1 U14810 ( .A1(n11466), .A2(n15427), .ZN(n11513) );
  OAI211_X1 U14811 ( .C1(n9613), .C2(P1_EBX_REG_16__SCAN_IN), .A(n11513), .B(
        n14651), .ZN(n11514) );
  NOR2_X2 U14812 ( .A1(n14875), .A2(n14860), .ZN(n14859) );
  MUX2_X1 U14813 ( .A(n11548), .B(n14671), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n11517) );
  NOR2_X1 U14814 ( .A1(n14652), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11516) );
  NOR2_X1 U14815 ( .A1(n11517), .A2(n11516), .ZN(n14842) );
  INV_X1 U14816 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n11518) );
  NAND2_X1 U14817 ( .A1(n11555), .A2(n11518), .ZN(n11521) );
  INV_X1 U14818 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15409) );
  NAND2_X1 U14819 ( .A1(n11466), .A2(n15409), .ZN(n11519) );
  OAI211_X1 U14820 ( .C1(n9614), .C2(P1_EBX_REG_18__SCAN_IN), .A(n11519), .B(
        n14651), .ZN(n11520) );
  MUX2_X1 U14821 ( .A(n11548), .B(n14671), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n11522) );
  INV_X1 U14822 ( .A(n11522), .ZN(n11525) );
  INV_X1 U14823 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15385) );
  NAND2_X1 U14824 ( .A1(n11523), .A2(n15385), .ZN(n11524) );
  NAND2_X1 U14825 ( .A1(n11525), .A2(n11524), .ZN(n14812) );
  INV_X1 U14826 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15386) );
  OAI21_X1 U14827 ( .B1(n14671), .B2(n15386), .A(n11466), .ZN(n11526) );
  OAI21_X1 U14828 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(n9614), .A(n11526), .ZN(
        n11527) );
  OAI21_X1 U14829 ( .B1(n11556), .B2(P1_EBX_REG_20__SCAN_IN), .A(n11527), .ZN(
        n14797) );
  AND2_X2 U14830 ( .A1(n14796), .A2(n14797), .ZN(n14799) );
  MUX2_X1 U14831 ( .A(n11548), .B(n14671), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n11529) );
  NOR2_X1 U14832 ( .A1(n14652), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11528) );
  NOR2_X1 U14833 ( .A1(n11529), .A2(n11528), .ZN(n14783) );
  INV_X1 U14834 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14958) );
  NAND2_X1 U14835 ( .A1(n11555), .A2(n14958), .ZN(n11532) );
  INV_X1 U14836 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15361) );
  NAND2_X1 U14837 ( .A1(n11466), .A2(n15361), .ZN(n11530) );
  OAI211_X1 U14838 ( .C1(n9614), .C2(P1_EBX_REG_22__SCAN_IN), .A(n11530), .B(
        n14651), .ZN(n11531) );
  INV_X1 U14839 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n11533) );
  NAND2_X1 U14840 ( .A1(n11548), .A2(n11533), .ZN(n11536) );
  NAND2_X1 U14841 ( .A1(n14651), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11534) );
  OAI211_X1 U14842 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n9613), .A(n11534), .B(
        n11466), .ZN(n11535) );
  NAND2_X1 U14843 ( .A1(n11536), .A2(n11535), .ZN(n14754) );
  INV_X1 U14844 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15343) );
  NAND2_X1 U14845 ( .A1(n11466), .A2(n15343), .ZN(n11537) );
  OAI211_X1 U14846 ( .C1(n9613), .C2(P1_EBX_REG_24__SCAN_IN), .A(n11537), .B(
        n14651), .ZN(n11538) );
  OAI21_X1 U14847 ( .B1(n11556), .B2(P1_EBX_REG_24__SCAN_IN), .A(n11538), .ZN(
        n14748) );
  INV_X1 U14848 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n11539) );
  NAND2_X1 U14849 ( .A1(n11548), .A2(n11539), .ZN(n11542) );
  NAND2_X1 U14850 ( .A1(n14651), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11540) );
  OAI211_X1 U14851 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n9614), .A(n11540), .B(
        n11466), .ZN(n11541) );
  NAND2_X1 U14852 ( .A1(n11542), .A2(n11541), .ZN(n14735) );
  INV_X1 U14853 ( .A(n11543), .ZN(n14734) );
  INV_X1 U14854 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n11544) );
  NAND2_X1 U14855 ( .A1(n11555), .A2(n11544), .ZN(n11547) );
  INV_X1 U14856 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15059) );
  NAND2_X1 U14857 ( .A1(n11466), .A2(n15059), .ZN(n11545) );
  OAI211_X1 U14858 ( .C1(n9614), .C2(P1_EBX_REG_26__SCAN_IN), .A(n11545), .B(
        n14651), .ZN(n11546) );
  MUX2_X1 U14859 ( .A(n11548), .B(n14671), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n11550) );
  NOR2_X1 U14860 ( .A1(n14652), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11549) );
  NOR2_X1 U14861 ( .A1(n11550), .A2(n11549), .ZN(n14703) );
  INV_X1 U14862 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n11554) );
  INV_X1 U14863 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11552) );
  NOR2_X1 U14864 ( .A1(n9613), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n11551) );
  AOI211_X1 U14865 ( .C1(n11552), .C2(n11466), .A(n14671), .B(n11551), .ZN(
        n11553) );
  AOI21_X1 U14866 ( .B1(n11555), .B2(n11554), .A(n11553), .ZN(n14693) );
  OAI22_X1 U14867 ( .A1(n14652), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(n9613), .ZN(n14669) );
  OAI22_X1 U14868 ( .A1(n14669), .A2(n14671), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n11556), .ZN(n11558) );
  OAI21_X1 U14869 ( .B1(n11557), .B2(n11558), .A(n14672), .ZN(n15297) );
  INV_X1 U14870 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n11559) );
  NAND2_X2 U14871 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20287), .ZN(n20237) );
  NOR2_X1 U14872 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19380) );
  INV_X1 U14873 ( .A(n19380), .ZN(n20177) );
  NAND3_X1 U14874 ( .A1(n20167), .A2(n20237), .A3(n20177), .ZN(n20173) );
  NOR2_X4 U14875 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11579) );
  AND2_X4 U14876 ( .A1(n11579), .A2(n11564), .ZN(n14447) );
  AOI22_X1 U14877 ( .A1(n11731), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14447), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11569) );
  INV_X1 U14878 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U14879 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9604), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11568) );
  AND2_X2 U14880 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11580) );
  AND2_X4 U14881 ( .A1(n11580), .A2(n11564), .ZN(n14454) );
  AND2_X4 U14882 ( .A1(n11580), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11733) );
  AOI22_X1 U14883 ( .A1(n14454), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11733), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11565) );
  AND2_X4 U14884 ( .A1(n11579), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11732) );
  AOI22_X1 U14885 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14610), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11566) );
  NAND4_X1 U14886 ( .A1(n11569), .A2(n11568), .A3(n11567), .A4(n11566), .ZN(
        n11574) );
  AOI22_X1 U14887 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U14888 ( .A1(n14454), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11733), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14889 ( .A1(n14601), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14610), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U14890 ( .A1(n11731), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14447), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11572) );
  NAND2_X1 U14891 ( .A1(n13916), .A2(n11785), .ZN(n11660) );
  BUF_X4 U14892 ( .A(n11731), .Z(n14605) );
  AND2_X2 U14893 ( .A1(n11718), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11941) );
  AOI22_X1 U14894 ( .A1(n12122), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14895 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n14463), .B1(
        n12094), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11577) );
  AND2_X4 U14896 ( .A1(n14605), .A2(n11839), .ZN(n14464) );
  AOI22_X1 U14897 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11576) );
  AND2_X2 U14898 ( .A1(n9606), .A2(n11839), .ZN(n14465) );
  AOI22_X1 U14899 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11575) );
  NAND4_X1 U14900 ( .A1(n11578), .A2(n11577), .A3(n11576), .A4(n11575), .ZN(
        n11588) );
  AND2_X2 U14901 ( .A1(n14509), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11661) );
  AOI22_X1 U14902 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n14470), .ZN(n11586) );
  INV_X1 U14903 ( .A(n11733), .ZN(n13854) );
  AND2_X2 U14904 ( .A1(n11733), .A2(n11839), .ZN(n14471) );
  AOI22_X1 U14905 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n14471), .B1(
        n11662), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11585) );
  AND2_X2 U14906 ( .A1(n14443), .A2(n13887), .ZN(n14473) );
  INV_X1 U14907 ( .A(n11581), .ZN(n13859) );
  AOI22_X1 U14908 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14909 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n14475), .B1(
        n14474), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11583) );
  NAND4_X1 U14910 ( .A1(n11586), .A2(n11585), .A3(n11584), .A4(n11583), .ZN(
        n11587) );
  NAND2_X1 U14911 ( .A1(n20034), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11632) );
  INV_X1 U14912 ( .A(n11632), .ZN(n11589) );
  NAND2_X1 U14913 ( .A1(n11675), .A2(n11589), .ZN(n11591) );
  NAND2_X1 U14914 ( .A1(n20032), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11590) );
  NAND2_X1 U14915 ( .A1(n11591), .A2(n11590), .ZN(n11629) );
  NAND2_X1 U14916 ( .A1(n11629), .A2(n11628), .ZN(n11593) );
  NAND2_X1 U14917 ( .A1(n20271), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11592) );
  XNOR2_X1 U14918 ( .A(n11625), .B(n11623), .ZN(n11746) );
  AOI22_X1 U14919 ( .A1(n11731), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14447), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U14920 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9604), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U14921 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U14922 ( .A1(n14454), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11733), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U14923 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U14924 ( .A1(n11731), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14447), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U14925 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14610), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U14926 ( .A1(n14454), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11733), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U14927 ( .A1(n11731), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14610), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14928 ( .A1(n14454), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11733), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14929 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14930 ( .A1(n14447), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11732), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11602) );
  NAND4_X1 U14931 ( .A1(n11605), .A2(n11604), .A3(n11603), .A4(n11602), .ZN(
        n11606) );
  AOI22_X1 U14932 ( .A1(n11731), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14447), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U14933 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9604), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U14934 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14454), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11608) );
  AOI22_X1 U14935 ( .A1(n9606), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11733), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11607) );
  NAND4_X1 U14936 ( .A1(n11610), .A2(n11609), .A3(n11608), .A4(n11607), .ZN(
        n11611) );
  AOI22_X1 U14937 ( .A1(n12122), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11616) );
  AOI22_X1 U14938 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U14939 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11662), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11614) );
  AOI22_X1 U14940 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n14471), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11613) );
  NAND4_X1 U14941 ( .A1(n11616), .A2(n11615), .A3(n11614), .A4(n11613), .ZN(
        n11622) );
  AOI22_X1 U14942 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n14472), .ZN(n11619) );
  AOI22_X1 U14943 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14474), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14944 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n14475), .B1(
        n14470), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11617) );
  NAND4_X1 U14945 ( .A1(n11620), .A2(n11619), .A3(n11618), .A4(n11617), .ZN(
        n11621) );
  INV_X1 U14946 ( .A(n11623), .ZN(n11624) );
  NAND2_X1 U14947 ( .A1(n11625), .A2(n11624), .ZN(n11627) );
  INV_X1 U14948 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20262) );
  NAND2_X1 U14949 ( .A1(n20262), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11626) );
  NAND2_X1 U14950 ( .A1(n11627), .A2(n11626), .ZN(n11641) );
  OR2_X1 U14951 ( .A1(n11641), .A2(n11642), .ZN(n11747) );
  XNOR2_X1 U14952 ( .A(n11629), .B(n11628), .ZN(n11687) );
  NAND2_X1 U14953 ( .A1(n11630), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11631) );
  NAND2_X1 U14954 ( .A1(n11632), .A2(n11631), .ZN(n11674) );
  INV_X1 U14955 ( .A(n11674), .ZN(n11745) );
  XNOR2_X1 U14956 ( .A(n11675), .B(n11632), .ZN(n11742) );
  NAND2_X1 U14957 ( .A1(n11745), .A2(n11675), .ZN(n11633) );
  AOI22_X1 U14958 ( .A1(n11634), .A2(n11773), .B1(n11780), .B2(n11633), .ZN(
        n11637) );
  NOR2_X1 U14959 ( .A1(n13395), .A2(n10064), .ZN(n11635) );
  MUX2_X1 U14960 ( .A(n11635), .B(n11780), .S(n10067), .Z(n11636) );
  OAI211_X1 U14961 ( .C1(n11637), .C2(n11636), .A(n11746), .B(n11747), .ZN(
        n11638) );
  OAI21_X1 U14962 ( .B1(n11690), .B2(n11780), .A(n11638), .ZN(n11644) );
  NOR2_X1 U14963 ( .A1(n11639), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11640) );
  NAND2_X1 U14964 ( .A1(n11644), .A2(n11743), .ZN(n11645) );
  MUX2_X1 U14965 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n11645), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n11658) );
  NAND2_X1 U14966 ( .A1(n11658), .A2(n11773), .ZN(n11655) );
  AOI22_X1 U14967 ( .A1(n14454), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11733), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14968 ( .A1(n14601), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14610), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14969 ( .A1(n11731), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14447), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U14970 ( .A1(n11731), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14447), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14971 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14610), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14972 ( .A1(n14454), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11733), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14973 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11652) );
  NAND3_X1 U14974 ( .A1(n10562), .A2(n11653), .A3(n11652), .ZN(n11654) );
  INV_X1 U14975 ( .A(n11778), .ZN(n19553) );
  NAND2_X1 U14976 ( .A1(n11655), .A2(n19553), .ZN(n11659) );
  INV_X1 U14977 ( .A(n11743), .ZN(n11656) );
  NAND2_X1 U14978 ( .A1(n13395), .A2(n11656), .ZN(n11657) );
  MUX2_X1 U14979 ( .A(n11660), .B(n11659), .S(n13868), .Z(n11770) );
  AOI22_X1 U14980 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__0__SCAN_IN), .B2(n14475), .ZN(n11666) );
  AOI22_X1 U14981 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n11662), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11665) );
  AOI22_X1 U14982 ( .A1(n14474), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14983 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n14470), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U14984 ( .A1(n12122), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14464), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U14985 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n11676), .B1(
        n14463), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14986 ( .A1(n11941), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14987 ( .A1(n14462), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11668) );
  INV_X1 U14988 ( .A(n13428), .ZN(n12011) );
  MUX2_X1 U14989 ( .A(n12011), .B(n11674), .S(n11800), .Z(n12391) );
  INV_X1 U14990 ( .A(n11675), .ZN(n11689) );
  AOI22_X1 U14991 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14992 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n14463), .B1(
        n11676), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14993 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n14464), .B1(
        n12094), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14994 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n14471), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11677) );
  NAND4_X1 U14995 ( .A1(n11680), .A2(n11679), .A3(n11678), .A4(n11677), .ZN(
        n11686) );
  AOI22_X1 U14996 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n14475), .ZN(n11684) );
  AOI22_X1 U14997 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n14465), .B1(
        n11662), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14998 ( .A1(n14474), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U14999 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n14470), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11681) );
  NAND4_X1 U15000 ( .A1(n11684), .A2(n11683), .A3(n11682), .A4(n11681), .ZN(
        n11685) );
  OAI21_X1 U15001 ( .B1(n12391), .B2(n11689), .A(n12372), .ZN(n11691) );
  NAND2_X1 U15002 ( .A1(n11691), .A2(n11690), .ZN(n11692) );
  NAND2_X1 U15003 ( .A1(n11692), .A2(n11743), .ZN(n20279) );
  AOI22_X1 U15004 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9604), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U15005 ( .A1(n11731), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14447), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U15006 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U15007 ( .A1(n14454), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11733), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11693) );
  NAND4_X1 U15008 ( .A1(n11696), .A2(n11695), .A3(n11694), .A4(n11693), .ZN(
        n11697) );
  AOI22_X1 U15009 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11701) );
  AOI22_X1 U15010 ( .A1(n11731), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14447), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U15011 ( .A1(n14454), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11733), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U15012 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14610), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11698) );
  NAND4_X1 U15013 ( .A1(n11701), .A2(n11700), .A3(n11699), .A4(n11698), .ZN(
        n11702) );
  NAND2_X1 U15014 ( .A1(n11702), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11703) );
  AOI22_X1 U15015 ( .A1(n11731), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14447), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U15016 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14610), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11706) );
  NOR2_X1 U15017 ( .A1(n10550), .A2(n10560), .ZN(n11705) );
  AOI22_X1 U15018 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U15019 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14610), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U15020 ( .A1(n11731), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14447), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U15021 ( .A1(n11731), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9604), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U15022 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U15023 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14447), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U15024 ( .A1(n14454), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11733), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11713) );
  NAND4_X1 U15025 ( .A1(n11716), .A2(n11715), .A3(n11714), .A4(n11713), .ZN(
        n11717) );
  NAND2_X1 U15026 ( .A1(n11717), .A2(n11839), .ZN(n11725) );
  AOI22_X1 U15027 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11722) );
  AOI22_X1 U15028 ( .A1(n11731), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14454), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11721) );
  AOI22_X1 U15029 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9605), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11720) );
  NAND4_X1 U15030 ( .A1(n11722), .A2(n11721), .A3(n11720), .A4(n11719), .ZN(
        n11723) );
  NAND2_X1 U15031 ( .A1(n11723), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11724) );
  AOI22_X1 U15032 ( .A1(n11731), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14447), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11730) );
  AOI22_X1 U15033 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9604), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11729) );
  AOI22_X1 U15034 ( .A1(n14454), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11733), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11726) );
  AOI22_X1 U15035 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14610), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11727) );
  NAND4_X1 U15036 ( .A1(n11730), .A2(n11729), .A3(n11728), .A4(n11727), .ZN(
        n11740) );
  AOI22_X1 U15037 ( .A1(n11718), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U15038 ( .A1(n11731), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14447), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U15039 ( .A1(n11732), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9606), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U15040 ( .A1(n14454), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11733), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11734) );
  NAND4_X1 U15041 ( .A1(n11738), .A2(n11737), .A3(n11736), .A4(n11735), .ZN(
        n11739) );
  NAND2_X2 U15042 ( .A1(n11740), .A2(n11739), .ZN(n13517) );
  NAND2_X1 U15043 ( .A1(n13913), .A2(n13928), .ZN(n11771) );
  NAND4_X1 U15044 ( .A1(n11747), .A2(n11746), .A3(n10067), .A4(n11742), .ZN(
        n11744) );
  NAND4_X1 U15045 ( .A1(n11747), .A2(n11746), .A3(n10067), .A4(n11745), .ZN(
        n11748) );
  AND2_X1 U15046 ( .A1(n11748), .A2(n16742), .ZN(n11749) );
  NAND2_X1 U15047 ( .A1(n13910), .A2(n11749), .ZN(n11754) );
  INV_X1 U15048 ( .A(n11890), .ZN(n11750) );
  AOI21_X1 U15049 ( .B1(n11581), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16810) );
  NAND2_X1 U15050 ( .A1(n11750), .A2(n16810), .ZN(n11752) );
  INV_X1 U15051 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n11751) );
  NAND2_X1 U15052 ( .A1(n11752), .A2(n11751), .ZN(n11753) );
  NAND2_X1 U15053 ( .A1(n11753), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13501) );
  NAND2_X1 U15054 ( .A1(n11754), .A2(n13501), .ZN(n20275) );
  NOR2_X1 U15055 ( .A1(n13517), .A2(n19545), .ZN(n11790) );
  NAND4_X1 U15056 ( .A1(n11792), .A2(n11791), .A3(n11773), .A4(n11790), .ZN(
        n11812) );
  NAND2_X1 U15057 ( .A1(n11782), .A2(n12331), .ZN(n11756) );
  NAND2_X1 U15058 ( .A1(n13911), .A2(n11756), .ZN(n11759) );
  NOR2_X1 U15059 ( .A1(n11778), .A2(n14561), .ZN(n12338) );
  INV_X1 U15060 ( .A(n13517), .ZN(n19577) );
  OAI211_X1 U15061 ( .C1(n12338), .C2(n16778), .A(n19545), .B(n19577), .ZN(
        n11757) );
  NAND2_X1 U15062 ( .A1(n11757), .A2(n12331), .ZN(n11758) );
  INV_X1 U15063 ( .A(n11772), .ZN(n11760) );
  NAND2_X1 U15064 ( .A1(n11760), .A2(n11786), .ZN(n11762) );
  NAND2_X1 U15065 ( .A1(n11762), .A2(n19577), .ZN(n11761) );
  NAND2_X1 U15066 ( .A1(n11761), .A2(n13928), .ZN(n12339) );
  NOR2_X4 U15067 ( .A1(n12008), .A2(n13517), .ZN(n13534) );
  NAND3_X1 U15068 ( .A1(n11823), .A2(n13910), .A3(n13916), .ZN(n11764) );
  MUX2_X1 U15069 ( .A(n11823), .B(n11785), .S(n10064), .Z(n11766) );
  NAND3_X1 U15070 ( .A1(n11766), .A2(n13910), .A3(n15574), .ZN(n11767) );
  NAND2_X1 U15071 ( .A1(n13865), .A2(n11767), .ZN(n11768) );
  INV_X1 U15072 ( .A(n11771), .ZN(n20278) );
  INV_X1 U15073 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n21270) );
  NOR2_X1 U15074 ( .A1(n11778), .A2(n13517), .ZN(n11804) );
  INV_X1 U15075 ( .A(n11794), .ZN(n11774) );
  NAND2_X1 U15076 ( .A1(n11780), .A2(n12331), .ZN(n11781) );
  AOI21_X1 U15077 ( .B1(n19545), .B2(n11794), .A(n11785), .ZN(n11789) );
  NAND3_X1 U15078 ( .A1(n11792), .A2(n11791), .A3(n11790), .ZN(n12318) );
  NAND2_X1 U15079 ( .A1(n11793), .A2(n12322), .ZN(n11795) );
  AOI21_X1 U15080 ( .B1(n11795), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n13395), 
        .ZN(n11796) );
  NAND2_X1 U15081 ( .A1(n11797), .A2(n11796), .ZN(n11798) );
  NOR2_X1 U15082 ( .A1(n11800), .A2(n14059), .ZN(n11801) );
  INV_X1 U15083 ( .A(n13926), .ZN(n11841) );
  NAND2_X1 U15084 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13429) );
  NAND2_X1 U15085 ( .A1(n11841), .A2(n13429), .ZN(n11802) );
  INV_X1 U15086 ( .A(n11840), .ZN(n11816) );
  NAND2_X1 U15087 ( .A1(n12209), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n11815) );
  NAND2_X1 U15088 ( .A1(n13928), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11809) );
  AND3_X1 U15089 ( .A1(n11803), .A2(n12331), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n11806) );
  NAND4_X1 U15090 ( .A1(n12320), .A2(n11806), .A3(n11805), .A4(n11804), .ZN(
        n11807) );
  AND2_X1 U15091 ( .A1(n11741), .A2(n19566), .ZN(n11811) );
  NAND2_X1 U15092 ( .A1(n11819), .A2(n11818), .ZN(n11820) );
  NOR2_X2 U15093 ( .A1(n11821), .A2(n11820), .ZN(n11827) );
  INV_X1 U15094 ( .A(n11822), .ZN(n11824) );
  NAND2_X1 U15095 ( .A1(n11823), .A2(n16778), .ZN(n12199) );
  NAND2_X1 U15096 ( .A1(n11824), .A2(n12199), .ZN(n12314) );
  AOI22_X1 U15097 ( .A1(n12314), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n13926), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11825) );
  NAND2_X1 U15098 ( .A1(n11852), .A2(n11853), .ZN(n11831) );
  INV_X1 U15099 ( .A(n11827), .ZN(n11828) );
  NAND2_X2 U15100 ( .A1(n11831), .A2(n11830), .ZN(n12203) );
  INV_X1 U15101 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13634) );
  OAI21_X1 U15102 ( .B1(n20271), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16742), 
        .ZN(n11834) );
  INV_X1 U15103 ( .A(n12202), .ZN(n11847) );
  INV_X1 U15104 ( .A(n12209), .ZN(n11838) );
  INV_X1 U15105 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13702) );
  NAND2_X1 U15106 ( .A1(n11840), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11842) );
  NAND2_X1 U15107 ( .A1(n11842), .A2(n10557), .ZN(n11843) );
  INV_X1 U15108 ( .A(n11850), .ZN(n11845) );
  INV_X1 U15109 ( .A(n12204), .ZN(n11844) );
  NAND2_X1 U15110 ( .A1(n12202), .A2(n11844), .ZN(n11848) );
  NAND2_X1 U15111 ( .A1(n11845), .A2(n11848), .ZN(n11846) );
  OR2_X2 U15112 ( .A1(n12203), .A2(n11846), .ZN(n11861) );
  NAND2_X1 U15113 ( .A1(n11847), .A2(n12204), .ZN(n11849) );
  MUX2_X1 U15114 ( .A(n11849), .B(n11848), .S(n11850), .Z(n11860) );
  AND2_X1 U15115 ( .A1(n11850), .A2(n11849), .ZN(n11851) );
  NAND2_X1 U15116 ( .A1(n12203), .A2(n11851), .ZN(n11859) );
  INV_X1 U15117 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11855) );
  NOR2_X1 U15118 ( .A1(n11858), .A2(n11857), .ZN(n11889) );
  INV_X1 U15119 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n21194) );
  AND2_X2 U15120 ( .A1(n11876), .A2(n9620), .ZN(n19661) );
  NAND2_X1 U15121 ( .A1(n19661), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11862) );
  OAI211_X1 U15122 ( .C1(n20043), .C2(n21194), .A(n11862), .B(n14561), .ZN(
        n11867) );
  INV_X1 U15123 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11865) );
  INV_X1 U15124 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11864) );
  OAI22_X1 U15125 ( .A1(n11905), .A2(n11865), .B1(n19630), .B2(n11864), .ZN(
        n11866) );
  NOR2_X1 U15126 ( .A1(n11867), .A2(n11866), .ZN(n11888) );
  INV_X1 U15127 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11870) );
  INV_X1 U15128 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11869) );
  OAI22_X1 U15129 ( .A1(n11870), .A2(n11906), .B1(n11907), .B2(n11869), .ZN(
        n11874) );
  INV_X1 U15130 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11872) );
  NOR2_X1 U15131 ( .A1(n11874), .A2(n11873), .ZN(n11887) );
  INV_X1 U15132 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11878) );
  INV_X1 U15133 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11877) );
  OAI22_X1 U15134 ( .A1(n11878), .A2(n11913), .B1(n11908), .B2(n11877), .ZN(
        n11885) );
  INV_X1 U15135 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11882) );
  INV_X1 U15136 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11881) );
  OAI22_X1 U15137 ( .A1(n11883), .A2(n11882), .B1(n19755), .B2(n11881), .ZN(
        n11884) );
  NOR2_X1 U15138 ( .A1(n11885), .A2(n11884), .ZN(n11886) );
  NAND4_X1 U15139 ( .A1(n11889), .A2(n11888), .A3(n11887), .A4(n11886), .ZN(
        n11903) );
  AOI22_X1 U15140 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n11941), .B1(
        n14461), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U15141 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n14463), .B1(
        n12094), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U15142 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U15143 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11891) );
  NAND4_X1 U15144 ( .A1(n11894), .A2(n11893), .A3(n11892), .A4(n11891), .ZN(
        n11900) );
  AOI22_X1 U15145 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n14470), .ZN(n11898) );
  AOI22_X1 U15146 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n14471), .B1(
        n11662), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11897) );
  AOI22_X1 U15147 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11896) );
  AOI22_X1 U15148 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14475), .B1(
        n14474), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11895) );
  NAND4_X1 U15149 ( .A1(n11898), .A2(n11897), .A3(n11896), .A4(n11895), .ZN(
        n11899) );
  NAND3_X1 U15150 ( .A1(n10064), .A2(n13428), .A3(n12371), .ZN(n11925) );
  NAND2_X1 U15151 ( .A1(n11925), .A2(n12022), .ZN(n11902) );
  AOI22_X1 U15152 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19990), .B1(
        n9662), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U15153 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19627), .B1(
        n19530), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U15154 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19587), .B1(
        n19661), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U15155 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19860), .B1(
        n9621), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11914) );
  INV_X1 U15156 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12342) );
  INV_X1 U15157 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13427) );
  AOI21_X1 U15158 ( .B1(n10064), .B2(n13428), .A(n13427), .ZN(n13426) );
  INV_X1 U15159 ( .A(n13426), .ZN(n11922) );
  XNOR2_X1 U15160 ( .A(n13428), .B(n12371), .ZN(n11921) );
  NOR2_X1 U15161 ( .A1(n11922), .A2(n11921), .ZN(n11924) );
  INV_X1 U15162 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13440) );
  AOI21_X1 U15163 ( .B1(n11922), .B2(n11921), .A(n11924), .ZN(n11923) );
  INV_X1 U15164 ( .A(n11923), .ZN(n13441) );
  NOR2_X1 U15165 ( .A1(n13440), .A2(n13441), .ZN(n13439) );
  NOR2_X1 U15166 ( .A1(n11924), .A2(n13439), .ZN(n11926) );
  XNOR2_X1 U15167 ( .A(n11925), .B(n12022), .ZN(n13667) );
  NAND2_X1 U15168 ( .A1(n9674), .A2(n13667), .ZN(n14637) );
  OR2_X1 U15169 ( .A1(n11926), .A2(n12342), .ZN(n11927) );
  NAND2_X1 U15170 ( .A1(n14637), .A2(n11927), .ZN(n11928) );
  INV_X1 U15171 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14151) );
  XNOR2_X1 U15172 ( .A(n11928), .B(n14151), .ZN(n13967) );
  NAND2_X1 U15173 ( .A1(n11928), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11929) );
  INV_X1 U15174 ( .A(n11930), .ZN(n12035) );
  INV_X1 U15175 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14207) );
  AOI22_X1 U15176 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n9621), .B1(
        n19919), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11936) );
  AOI22_X1 U15177 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19990), .B1(
        n9662), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11935) );
  AOI22_X1 U15178 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19693), .B1(
        n19661), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11934) );
  AOI22_X1 U15179 ( .A1(n19828), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n19727), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U15180 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n16774), .B1(
        n20039), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11940) );
  AOI22_X1 U15181 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19530), .B1(
        n19587), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11939) );
  AOI22_X1 U15182 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19627), .B1(
        n19759), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U15183 ( .A1(n19860), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11956), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U15184 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11946) );
  AOI22_X1 U15185 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n14463), .B1(
        n14462), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U15186 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11944) );
  AOI22_X1 U15187 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11943) );
  NAND4_X1 U15188 ( .A1(n11946), .A2(n11945), .A3(n11944), .A4(n11943), .ZN(
        n11952) );
  AOI22_X1 U15189 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__5__SCAN_IN), .B2(n14470), .ZN(n11950) );
  AOI22_X1 U15190 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n11662), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U15191 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U15192 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n14475), .B1(
        n14474), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11947) );
  NAND4_X1 U15193 ( .A1(n11950), .A2(n11949), .A3(n11948), .A4(n11947), .ZN(
        n11951) );
  INV_X1 U15194 ( .A(n12379), .ZN(n12043) );
  NAND2_X1 U15195 ( .A1(n12043), .A2(n10064), .ZN(n11953) );
  INV_X1 U15196 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14208) );
  INV_X1 U15197 ( .A(n11954), .ZN(n11955) );
  NAND2_X1 U15198 ( .A1(n11955), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11975) );
  AOI22_X1 U15199 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19759), .B1(
        n11956), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U15200 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19627), .B1(
        n19661), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U15201 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19587), .B1(
        n19530), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U15202 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20039), .B1(
        n9662), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U15203 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19860), .B1(
        n19828), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11960) );
  AOI22_X1 U15204 ( .A1(n12122), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14464), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U15205 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n11941), .B1(
        n14463), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11964) );
  AOI22_X1 U15206 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U15207 ( .A1(n14462), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11962) );
  NAND4_X1 U15208 ( .A1(n11965), .A2(n11964), .A3(n11963), .A4(n11962), .ZN(
        n11971) );
  AOI22_X1 U15209 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n14472), .ZN(n11969) );
  AOI22_X1 U15210 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n14471), .B1(
        n11662), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11968) );
  AOI22_X1 U15211 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14474), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U15212 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n14475), .B1(
        n14470), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11966) );
  NAND4_X1 U15213 ( .A1(n11969), .A2(n11968), .A3(n11967), .A4(n11966), .ZN(
        n11970) );
  NAND2_X1 U15214 ( .A1(n12381), .A2(n10064), .ZN(n11972) );
  XNOR2_X1 U15215 ( .A(n12368), .B(n11978), .ZN(n11976) );
  INV_X1 U15216 ( .A(n11976), .ZN(n11974) );
  INV_X1 U15217 ( .A(n11975), .ZN(n14202) );
  INV_X1 U15218 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11977) );
  INV_X1 U15219 ( .A(n12368), .ZN(n11979) );
  NAND2_X1 U15220 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11983) );
  NAND2_X1 U15221 ( .A1(n12122), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11982) );
  NAND2_X1 U15222 ( .A1(n11941), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11981) );
  NAND2_X1 U15223 ( .A1(n14463), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11980) );
  AOI22_X1 U15224 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n14475), .B1(
        n14470), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11987) );
  NAND2_X1 U15225 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11986) );
  AOI22_X1 U15226 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14474), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11985) );
  NAND2_X1 U15227 ( .A1(n14472), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11984) );
  NAND2_X1 U15228 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11991) );
  NAND2_X1 U15229 ( .A1(n12094), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11990) );
  NAND2_X1 U15230 ( .A1(n11662), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11989) );
  NAND2_X1 U15231 ( .A1(n11612), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11988) );
  AOI22_X1 U15232 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n14465), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11992) );
  XNOR2_X1 U15233 ( .A(n11996), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16403) );
  INV_X1 U15234 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16681) );
  NAND2_X1 U15235 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16591) );
  INV_X1 U15236 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16361) );
  NOR3_X1 U15237 ( .A1(n16654), .A2(n9601), .A3(n16361), .ZN(n16629) );
  NAND2_X1 U15238 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16629), .ZN(
        n12000) );
  NOR2_X1 U15239 ( .A1(n16591), .A2(n12000), .ZN(n14316) );
  AND3_X1 U15240 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12001) );
  NAND2_X1 U15241 ( .A1(n14316), .A2(n12001), .ZN(n16288) );
  INV_X1 U15242 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12454) );
  OR2_X1 U15243 ( .A1(n16288), .A2(n12454), .ZN(n16534) );
  NAND2_X1 U15244 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12002) );
  NOR2_X1 U15245 ( .A1(n16534), .A2(n12002), .ZN(n16519) );
  INV_X1 U15246 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16255) );
  INV_X1 U15247 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16498) );
  INV_X1 U15248 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16471) );
  AND2_X1 U15249 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13002) );
  NAND2_X1 U15250 ( .A1(n13002), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12570) );
  XNOR2_X1 U15251 ( .A(n12988), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16181) );
  NAND2_X1 U15252 ( .A1(n12003), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12007) );
  NAND2_X1 U15253 ( .A1(n13517), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12005) );
  AND2_X1 U15254 ( .A1(n12005), .A2(n12004), .ZN(n12006) );
  NAND2_X1 U15255 ( .A1(n12007), .A2(n12006), .ZN(n13548) );
  NAND2_X2 U15256 ( .A1(n12009), .A2(n12532), .ZN(n12162) );
  MUX2_X1 U15257 ( .A(n19577), .B(n20034), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12010) );
  OR2_X1 U15258 ( .A1(n11794), .A2(n12193), .ZN(n12023) );
  NAND2_X1 U15259 ( .A1(n13548), .A2(n13547), .ZN(n12018) );
  INV_X1 U15260 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20184) );
  OR2_X1 U15261 ( .A1(n12189), .A2(n20184), .ZN(n12013) );
  AOI22_X1 U15262 ( .A1(n12045), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12559), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12012) );
  NAND2_X1 U15263 ( .A1(n12013), .A2(n12012), .ZN(n12019) );
  XNOR2_X1 U15264 ( .A(n12018), .B(n12019), .ZN(n13793) );
  NAND2_X1 U15265 ( .A1(n11794), .A2(n19577), .ZN(n12014) );
  MUX2_X1 U15266 ( .A(n12014), .B(n20032), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12017) );
  INV_X1 U15267 ( .A(n12371), .ZN(n12015) );
  OR2_X1 U15268 ( .A1(n12162), .A2(n12015), .ZN(n12016) );
  AND2_X1 U15269 ( .A1(n12017), .A2(n12016), .ZN(n13792) );
  INV_X1 U15270 ( .A(n12019), .ZN(n12020) );
  NAND2_X1 U15271 ( .A1(n12018), .A2(n12020), .ZN(n12021) );
  NAND2_X1 U15272 ( .A1(n13794), .A2(n12021), .ZN(n12028) );
  OR2_X1 U15273 ( .A1(n12162), .A2(n12022), .ZN(n12024) );
  OAI211_X1 U15274 ( .C1(n20104), .C2(n20271), .A(n12024), .B(n12023), .ZN(
        n12026) );
  XNOR2_X1 U15275 ( .A(n12028), .B(n12026), .ZN(n13659) );
  INV_X1 U15276 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19473) );
  OAI22_X1 U15277 ( .A1(n12195), .A2(n19473), .B1(n12193), .B2(n12342), .ZN(
        n12025) );
  AOI21_X1 U15278 ( .B1(n12003), .B2(P2_REIP_REG_2__SCAN_IN), .A(n12025), .ZN(
        n13658) );
  INV_X1 U15279 ( .A(n12026), .ZN(n12027) );
  NAND2_X1 U15280 ( .A1(n12028), .A2(n12027), .ZN(n12029) );
  INV_X1 U15281 ( .A(n12162), .ZN(n12030) );
  NAND2_X1 U15282 ( .A1(n12003), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U15283 ( .A1(n12559), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12031) );
  AOI22_X1 U15284 ( .A1(n12045), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12559), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12037) );
  OR2_X1 U15285 ( .A1(n12162), .A2(n12035), .ZN(n12036) );
  AND2_X1 U15286 ( .A1(n12037), .A2(n12036), .ZN(n12039) );
  NAND2_X1 U15287 ( .A1(n12003), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12038) );
  INV_X1 U15288 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n12040) );
  OR2_X1 U15289 ( .A1(n12189), .A2(n12040), .ZN(n12042) );
  AOI22_X1 U15290 ( .A1(n12045), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12559), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12041) );
  OAI211_X1 U15291 ( .C1(n12043), .C2(n12162), .A(n12042), .B(n12041), .ZN(
        n14071) );
  OR2_X1 U15292 ( .A1(n12162), .A2(n12381), .ZN(n12044) );
  INV_X1 U15293 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20193) );
  OR2_X1 U15294 ( .A1(n12189), .A2(n20193), .ZN(n12047) );
  AOI22_X1 U15295 ( .A1(n12045), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12559), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12046) );
  NAND2_X1 U15296 ( .A1(n12047), .A2(n12046), .ZN(n13541) );
  NAND2_X1 U15297 ( .A1(n13540), .A2(n13541), .ZN(n12050) );
  OR2_X1 U15298 ( .A1(n12162), .A2(n12048), .ZN(n12049) );
  INV_X1 U15299 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20195) );
  OR2_X1 U15300 ( .A1(n12189), .A2(n20195), .ZN(n12052) );
  AOI22_X1 U15301 ( .A1(n12045), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n12559), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12051) );
  NAND2_X1 U15302 ( .A1(n12052), .A2(n12051), .ZN(n13529) );
  INV_X1 U15303 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20197) );
  OR2_X1 U15304 ( .A1(n12189), .A2(n20197), .ZN(n12065) );
  AOI22_X1 U15305 ( .A1(n12045), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12559), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U15306 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14464), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12056) );
  AOI22_X1 U15307 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n11941), .B1(
        n14462), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12055) );
  AOI22_X1 U15308 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11662), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12054) );
  AOI22_X1 U15309 ( .A1(n14463), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12053) );
  NAND4_X1 U15310 ( .A1(n12056), .A2(n12055), .A3(n12054), .A4(n12053), .ZN(
        n12062) );
  AOI22_X1 U15311 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U15312 ( .A1(n14465), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U15313 ( .A1(n14474), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U15314 ( .A1(n14475), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14470), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12057) );
  NAND4_X1 U15315 ( .A1(n12060), .A2(n12059), .A3(n12058), .A4(n12057), .ZN(
        n12061) );
  INV_X1 U15316 ( .A(n13818), .ZN(n14103) );
  OR2_X1 U15317 ( .A1(n12162), .A2(n14103), .ZN(n12063) );
  AOI22_X1 U15318 ( .A1(n12045), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12559), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15319 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U15320 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n14464), .B1(
        n14462), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15321 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n11662), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U15322 ( .A1(n14463), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12067) );
  NAND4_X1 U15323 ( .A1(n12070), .A2(n12069), .A3(n12068), .A4(n12067), .ZN(
        n12076) );
  AOI22_X1 U15324 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n14472), .ZN(n12074) );
  AOI22_X1 U15325 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12073) );
  AOI22_X1 U15326 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n14474), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U15327 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n14475), .B1(
        n14470), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12071) );
  NAND4_X1 U15328 ( .A1(n12074), .A2(n12073), .A3(n12072), .A4(n12071), .ZN(
        n12075) );
  NOR2_X1 U15329 ( .A1(n12076), .A2(n12075), .ZN(n13823) );
  OR2_X1 U15330 ( .A1(n12162), .A2(n13823), .ZN(n12077) );
  AND2_X1 U15331 ( .A1(n12078), .A2(n12077), .ZN(n12080) );
  NAND2_X1 U15332 ( .A1(n12003), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12079) );
  INV_X1 U15333 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20199) );
  OR2_X1 U15334 ( .A1(n12189), .A2(n20199), .ZN(n12093) );
  AOI22_X1 U15335 ( .A1(n12045), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12559), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15336 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11941), .B1(
        n14461), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U15337 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n14463), .B1(
        n14462), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U15338 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15339 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12081) );
  NAND4_X1 U15340 ( .A1(n12084), .A2(n12083), .A3(n12082), .A4(n12081), .ZN(
        n12090) );
  AOI22_X1 U15341 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n14470), .ZN(n12088) );
  AOI22_X1 U15342 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11662), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12087) );
  AOI22_X1 U15343 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U15344 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n14475), .B1(
        n14474), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12085) );
  NAND4_X1 U15345 ( .A1(n12088), .A2(n12087), .A3(n12086), .A4(n12085), .ZN(
        n12089) );
  NOR2_X1 U15346 ( .A1(n12090), .A2(n12089), .ZN(n13955) );
  OR2_X1 U15347 ( .A1(n12162), .A2(n13955), .ZN(n12091) );
  AOI22_X1 U15348 ( .A1(n12045), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12559), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12107) );
  AOI22_X1 U15349 ( .A1(n12122), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U15350 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n14463), .B1(
        n12094), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U15351 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15352 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12095) );
  NAND4_X1 U15353 ( .A1(n12098), .A2(n12097), .A3(n12096), .A4(n12095), .ZN(
        n12104) );
  AOI22_X1 U15354 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n14470), .ZN(n12102) );
  AOI22_X1 U15355 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11662), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U15356 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U15357 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n14475), .B1(
        n14474), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12099) );
  NAND4_X1 U15358 ( .A1(n12102), .A2(n12101), .A3(n12100), .A4(n12099), .ZN(
        n12103) );
  INV_X1 U15359 ( .A(n14186), .ZN(n12105) );
  OR2_X1 U15360 ( .A1(n12162), .A2(n12105), .ZN(n12106) );
  AND2_X1 U15361 ( .A1(n12107), .A2(n12106), .ZN(n12109) );
  NAND2_X1 U15362 ( .A1(n12003), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15363 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12113) );
  AOI22_X1 U15364 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11676), .B1(
        n14462), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12112) );
  AOI22_X1 U15365 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12111) );
  AOI22_X1 U15366 ( .A1(n14463), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12110) );
  NAND4_X1 U15367 ( .A1(n12113), .A2(n12112), .A3(n12111), .A4(n12110), .ZN(
        n12119) );
  AOI22_X1 U15368 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n14472), .ZN(n12117) );
  AOI22_X1 U15369 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11662), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U15370 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n14474), .B1(
        n14470), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U15371 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14475), .B1(
        n14473), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12114) );
  NAND4_X1 U15372 ( .A1(n12117), .A2(n12116), .A3(n12115), .A4(n12114), .ZN(
        n12118) );
  OR2_X1 U15373 ( .A1(n12119), .A2(n12118), .ZN(n14184) );
  INV_X1 U15374 ( .A(n14184), .ZN(n14087) );
  INV_X1 U15375 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20205) );
  OR2_X1 U15376 ( .A1(n12189), .A2(n20205), .ZN(n12121) );
  AOI22_X1 U15377 ( .A1(n12045), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12559), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12120) );
  OAI211_X1 U15378 ( .C1(n14087), .C2(n12162), .A(n12121), .B(n12120), .ZN(
        n13778) );
  NAND2_X1 U15379 ( .A1(n13779), .A2(n13778), .ZN(n13777) );
  INV_X1 U15380 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n20207) );
  OR2_X1 U15381 ( .A1(n12189), .A2(n20207), .ZN(n12136) );
  AOI22_X1 U15382 ( .A1(n12045), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12559), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U15383 ( .A1(n12122), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12126) );
  AOI22_X1 U15384 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n14463), .B1(
        n14462), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12125) );
  AOI22_X1 U15385 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12124) );
  AOI22_X1 U15386 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12123) );
  NAND4_X1 U15387 ( .A1(n12126), .A2(n12125), .A3(n12124), .A4(n12123), .ZN(
        n12132) );
  AOI22_X1 U15388 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__5__SCAN_IN), .B2(n14470), .ZN(n12130) );
  AOI22_X1 U15389 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n11662), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15390 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12128) );
  AOI22_X1 U15391 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n14475), .B1(
        n14474), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12127) );
  NAND4_X1 U15392 ( .A1(n12130), .A2(n12129), .A3(n12128), .A4(n12127), .ZN(
        n12131) );
  INV_X1 U15393 ( .A(n14185), .ZN(n12133) );
  OR2_X1 U15394 ( .A1(n12162), .A2(n12133), .ZN(n12134) );
  INV_X1 U15395 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n21272) );
  OR2_X1 U15396 ( .A1(n12189), .A2(n21272), .ZN(n12149) );
  AOI22_X1 U15397 ( .A1(n12045), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12559), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15398 ( .A1(n12122), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12140) );
  AOI22_X1 U15399 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n14463), .B1(
        n14462), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U15400 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U15401 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12137) );
  NAND4_X1 U15402 ( .A1(n12140), .A2(n12139), .A3(n12138), .A4(n12137), .ZN(
        n12146) );
  AOI22_X1 U15403 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n14470), .ZN(n12144) );
  AOI22_X1 U15404 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11662), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12143) );
  AOI22_X1 U15405 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12142) );
  AOI22_X1 U15406 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14475), .B1(
        n14474), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12141) );
  NAND4_X1 U15407 ( .A1(n12144), .A2(n12143), .A3(n12142), .A4(n12141), .ZN(
        n12145) );
  OR2_X1 U15408 ( .A1(n12146), .A2(n12145), .ZN(n14187) );
  INV_X1 U15409 ( .A(n14187), .ZN(n14181) );
  OR2_X1 U15410 ( .A1(n12162), .A2(n14181), .ZN(n12147) );
  AOI22_X1 U15411 ( .A1(n12122), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U15412 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n14463), .B1(
        n14462), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15413 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U15414 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12150) );
  NAND4_X1 U15415 ( .A1(n12153), .A2(n12152), .A3(n12151), .A4(n12150), .ZN(
        n12159) );
  AOI22_X1 U15416 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n14470), .ZN(n12157) );
  AOI22_X1 U15417 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11662), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U15418 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12155) );
  AOI22_X1 U15419 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14475), .B1(
        n14474), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12154) );
  NAND4_X1 U15420 ( .A1(n12157), .A2(n12156), .A3(n12155), .A4(n12154), .ZN(
        n12158) );
  NOR2_X1 U15421 ( .A1(n12159), .A2(n12158), .ZN(n14183) );
  INV_X1 U15422 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20210) );
  OR2_X1 U15423 ( .A1(n12189), .A2(n20210), .ZN(n12161) );
  AOI22_X1 U15424 ( .A1(n12045), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12559), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12160) );
  OAI211_X1 U15425 ( .C1(n14183), .C2(n12162), .A(n12161), .B(n12160), .ZN(
        n14037) );
  INV_X1 U15426 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n12163) );
  OR2_X1 U15427 ( .A1(n12189), .A2(n12163), .ZN(n12165) );
  AOI22_X1 U15428 ( .A1(n12045), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12559), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12164) );
  NAND2_X1 U15429 ( .A1(n12165), .A2(n12164), .ZN(n15762) );
  INV_X1 U15430 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20217) );
  OR2_X1 U15431 ( .A1(n12189), .A2(n20217), .ZN(n12167) );
  AOI22_X1 U15432 ( .A1(n12045), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12559), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12166) );
  NAND2_X1 U15433 ( .A1(n12167), .A2(n12166), .ZN(n15729) );
  INV_X1 U15434 ( .A(n15729), .ZN(n12171) );
  INV_X1 U15435 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n12168) );
  OAI22_X1 U15436 ( .A1(n12195), .A2(n12168), .B1(n12193), .B2(n12454), .ZN(
        n12169) );
  AOI21_X1 U15437 ( .B1(n12003), .B2(P2_REIP_REG_18__SCAN_IN), .A(n12169), 
        .ZN(n15746) );
  INV_X1 U15438 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13413) );
  INV_X1 U15439 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16301) );
  OAI22_X1 U15440 ( .A1(n12195), .A2(n13413), .B1(n12193), .B2(n16301), .ZN(
        n12170) );
  AOI21_X1 U15441 ( .B1(n12003), .B2(P2_REIP_REG_17__SCAN_IN), .A(n12170), 
        .ZN(n14336) );
  OR2_X1 U15442 ( .A1(n15746), .A2(n14336), .ZN(n15728) );
  INV_X1 U15443 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20219) );
  OR2_X1 U15444 ( .A1(n12189), .A2(n20219), .ZN(n12173) );
  AOI22_X1 U15445 ( .A1(n12045), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12559), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12172) );
  NAND2_X1 U15446 ( .A1(n12173), .A2(n12172), .ZN(n15701) );
  INV_X1 U15447 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13408) );
  OAI22_X1 U15448 ( .A1(n12195), .A2(n13408), .B1(n12193), .B2(n16255), .ZN(
        n12174) );
  AOI21_X1 U15449 ( .B1(n12003), .B2(P2_REIP_REG_21__SCAN_IN), .A(n12174), 
        .ZN(n15689) );
  INV_X1 U15450 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n12177) );
  INV_X1 U15451 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12507) );
  OAI22_X1 U15452 ( .A1(n12195), .A2(n12177), .B1(n12193), .B2(n12507), .ZN(
        n12178) );
  AOI21_X1 U15453 ( .B1(n12003), .B2(P2_REIP_REG_22__SCAN_IN), .A(n12178), 
        .ZN(n16112) );
  INV_X1 U15454 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20225) );
  OR2_X1 U15455 ( .A1(n12189), .A2(n20225), .ZN(n12180) );
  AOI22_X1 U15456 ( .A1(n12045), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12559), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12179) );
  NAND2_X1 U15457 ( .A1(n12180), .A2(n12179), .ZN(n15672) );
  INV_X1 U15458 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n12181) );
  INV_X1 U15459 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16484) );
  OAI22_X1 U15460 ( .A1(n12195), .A2(n12181), .B1(n12193), .B2(n16484), .ZN(
        n12182) );
  AOI21_X1 U15461 ( .B1(n12003), .B2(P2_REIP_REG_24__SCAN_IN), .A(n12182), 
        .ZN(n15653) );
  INV_X1 U15462 ( .A(n15653), .ZN(n12183) );
  INV_X1 U15463 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13419) );
  OAI22_X1 U15464 ( .A1(n12195), .A2(n13419), .B1(n12193), .B2(n16471), .ZN(
        n12184) );
  AOI21_X1 U15465 ( .B1(n12003), .B2(P2_REIP_REG_25__SCAN_IN), .A(n12184), 
        .ZN(n15636) );
  INV_X1 U15466 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20230) );
  OR2_X1 U15467 ( .A1(n12189), .A2(n20230), .ZN(n12186) );
  AOI22_X1 U15468 ( .A1(n12045), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12559), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12185) );
  INV_X1 U15469 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20233) );
  OR2_X1 U15470 ( .A1(n12189), .A2(n20233), .ZN(n12188) );
  AOI22_X1 U15471 ( .A1(n12045), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12559), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12187) );
  NAND2_X1 U15472 ( .A1(n12188), .A2(n12187), .ZN(n12747) );
  INV_X1 U15473 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20234) );
  OR2_X1 U15474 ( .A1(n12189), .A2(n20234), .ZN(n12191) );
  AOI22_X1 U15475 ( .A1(n12045), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12559), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12190) );
  NAND2_X1 U15476 ( .A1(n12191), .A2(n12190), .ZN(n15593) );
  INV_X1 U15477 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13424) );
  INV_X1 U15478 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13001) );
  OAI22_X1 U15479 ( .A1(n12195), .A2(n13424), .B1(n12193), .B2(n13001), .ZN(
        n12192) );
  AOI21_X1 U15480 ( .B1(n12003), .B2(P2_REIP_REG_29__SCAN_IN), .A(n12192), 
        .ZN(n13007) );
  INV_X1 U15481 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12194) );
  INV_X1 U15482 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12569) );
  OAI22_X1 U15483 ( .A1(n12195), .A2(n12194), .B1(n12193), .B2(n12569), .ZN(
        n12196) );
  AOI21_X1 U15484 ( .B1(n12003), .B2(P2_REIP_REG_30__SCAN_IN), .A(n12196), 
        .ZN(n12197) );
  AND2_X1 U15485 ( .A1(n13009), .A2(n12197), .ZN(n12198) );
  NAND2_X1 U15486 ( .A1(n12199), .A2(n13911), .ZN(n13903) );
  NAND2_X1 U15487 ( .A1(n13906), .A2(n12200), .ZN(n12201) );
  NOR2_X1 U15488 ( .A1(n14623), .A2(n16708), .ZN(n12366) );
  NAND2_X1 U15489 ( .A1(n12203), .A2(n12202), .ZN(n12206) );
  NAND2_X1 U15490 ( .A1(n12206), .A2(n12205), .ZN(n13773) );
  AOI22_X1 U15491 ( .A1(n12230), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12207) );
  AND2_X1 U15492 ( .A1(n12208), .A2(n12207), .ZN(n12211) );
  NAND2_X1 U15493 ( .A1(n12302), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n12210) );
  AND2_X1 U15494 ( .A1(n12211), .A2(n12210), .ZN(n13772) );
  AOI22_X1 U15495 ( .A1(n12230), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12214) );
  AND2_X1 U15496 ( .A1(n12215), .A2(n12214), .ZN(n12217) );
  NAND2_X1 U15497 ( .A1(n12302), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n12216) );
  AND2_X1 U15498 ( .A1(n12217), .A2(n12216), .ZN(n13803) );
  AOI22_X1 U15499 ( .A1(n12230), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12220) );
  OAI211_X1 U15500 ( .C1(n12218), .C2(n21330), .A(n12220), .B(n12219), .ZN(
        n12221) );
  INV_X1 U15501 ( .A(n12221), .ZN(n13844) );
  INV_X1 U15502 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U15503 ( .A1(n12230), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12223) );
  OAI211_X1 U15504 ( .C1(n12218), .C2(n12413), .A(n12223), .B(n12222), .ZN(
        n13836) );
  AOI22_X1 U15505 ( .A1(n12230), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12224) );
  AND2_X1 U15506 ( .A1(n12225), .A2(n12224), .ZN(n12227) );
  NAND2_X1 U15507 ( .A1(n12302), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15508 ( .A1(n12563), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12231) );
  AND2_X1 U15509 ( .A1(n12232), .A2(n12231), .ZN(n12234) );
  NAND2_X1 U15510 ( .A1(n12302), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12233) );
  INV_X1 U15511 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U15512 ( .A1(n12563), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n12236) );
  OAI211_X1 U15513 ( .C1(n12218), .C2(n12426), .A(n12236), .B(n12235), .ZN(
        n13828) );
  AOI22_X1 U15514 ( .A1(n12563), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n12237) );
  AND2_X1 U15515 ( .A1(n12238), .A2(n12237), .ZN(n12240) );
  NAND2_X1 U15516 ( .A1(n12302), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U15517 ( .A1(n12563), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n12243) );
  AND2_X1 U15518 ( .A1(n12244), .A2(n12243), .ZN(n12246) );
  NAND2_X1 U15519 ( .A1(n12302), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U15520 ( .A1(n12563), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n12247) );
  AND2_X1 U15521 ( .A1(n12248), .A2(n12247), .ZN(n12250) );
  NAND2_X1 U15522 ( .A1(n12302), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12249) );
  INV_X1 U15523 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n12448) );
  AOI22_X1 U15524 ( .A1(n12563), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n12252) );
  OAI211_X1 U15525 ( .C1(n12218), .C2(n12448), .A(n12252), .B(n12251), .ZN(
        n14161) );
  AOI22_X1 U15526 ( .A1(n12563), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n12253) );
  AND2_X1 U15527 ( .A1(n12254), .A2(n12253), .ZN(n12256) );
  NAND2_X1 U15528 ( .A1(n12302), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U15529 ( .A1(n12563), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n12259) );
  AND2_X1 U15530 ( .A1(n12260), .A2(n12259), .ZN(n12262) );
  NAND2_X1 U15531 ( .A1(n12302), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12261) );
  INV_X1 U15532 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15533 ( .A1(n12563), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n12264) );
  OAI211_X1 U15534 ( .C1(n12218), .C2(n12265), .A(n12264), .B(n12263), .ZN(
        n14332) );
  AOI22_X1 U15535 ( .A1(n12563), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n12266) );
  AND2_X1 U15536 ( .A1(n12267), .A2(n12266), .ZN(n12269) );
  NAND2_X1 U15537 ( .A1(n12302), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15538 ( .A1(n12563), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n12270) );
  AND2_X1 U15539 ( .A1(n12271), .A2(n12270), .ZN(n12273) );
  NAND2_X1 U15540 ( .A1(n12302), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15541 ( .A1(n12563), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n12276) );
  OAI211_X1 U15542 ( .C1(n12218), .C2(n10455), .A(n12276), .B(n12275), .ZN(
        n15703) );
  INV_X1 U15543 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n12279) );
  AOI22_X1 U15544 ( .A1(n12563), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n12278) );
  OAI211_X1 U15545 ( .C1(n12218), .C2(n12279), .A(n12278), .B(n12277), .ZN(
        n15641) );
  AOI22_X1 U15546 ( .A1(n12563), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n12280) );
  AND2_X1 U15547 ( .A1(n12281), .A2(n12280), .ZN(n12283) );
  NAND2_X1 U15548 ( .A1(n12302), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12282) );
  AND2_X1 U15549 ( .A1(n12283), .A2(n12282), .ZN(n15657) );
  AOI22_X1 U15550 ( .A1(n12563), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n12284) );
  AND2_X1 U15551 ( .A1(n12285), .A2(n12284), .ZN(n12287) );
  NAND2_X1 U15552 ( .A1(n12302), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12286) );
  AND2_X1 U15553 ( .A1(n12287), .A2(n12286), .ZN(n15674) );
  AOI22_X1 U15554 ( .A1(n12563), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n12288) );
  AND2_X1 U15555 ( .A1(n12289), .A2(n12288), .ZN(n12291) );
  NAND2_X1 U15556 ( .A1(n12302), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12290) );
  NOR2_X1 U15557 ( .A1(n15657), .A2(n15656), .ZN(n15638) );
  AND2_X1 U15558 ( .A1(n15641), .A2(n15638), .ZN(n12294) );
  INV_X1 U15559 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U15560 ( .A1(n12563), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n12293) );
  OAI211_X1 U15561 ( .C1(n12218), .C2(n12459), .A(n12293), .B(n12292), .ZN(
        n15695) );
  AND2_X1 U15562 ( .A1(n12294), .A2(n15695), .ZN(n12295) );
  AOI22_X1 U15563 ( .A1(n12563), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n12296) );
  AND2_X1 U15564 ( .A1(n12297), .A2(n12296), .ZN(n12299) );
  NAND2_X1 U15565 ( .A1(n12302), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15566 ( .A1(n12563), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12300) );
  AND2_X1 U15567 ( .A1(n12301), .A2(n12300), .ZN(n12304) );
  NAND2_X1 U15568 ( .A1(n12302), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12303) );
  INV_X1 U15569 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n12531) );
  AOI22_X1 U15570 ( .A1(n12563), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12306) );
  OAI211_X1 U15571 ( .C1(n12218), .C2(n12531), .A(n12306), .B(n12305), .ZN(
        n15596) );
  INV_X1 U15572 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U15573 ( .A1(n12563), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12308) );
  OAI211_X1 U15574 ( .C1(n12218), .C2(n12309), .A(n12308), .B(n12307), .ZN(
        n12995) );
  INV_X1 U15575 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n14632) );
  AOI22_X1 U15576 ( .A1(n12563), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12311) );
  OAI211_X1 U15577 ( .C1(n12218), .C2(n14632), .A(n12311), .B(n12310), .ZN(
        n12312) );
  OR2_X1 U15578 ( .A1(n12997), .A2(n12312), .ZN(n12313) );
  NAND2_X1 U15579 ( .A1(n13892), .A2(n10064), .ZN(n12316) );
  NAND2_X1 U15580 ( .A1(n12316), .A2(n12315), .ZN(n12317) );
  NAND3_X1 U15581 ( .A1(n12319), .A2(n11773), .A3(n12318), .ZN(n12327) );
  NAND2_X1 U15582 ( .A1(n10012), .A2(n11778), .ZN(n12321) );
  INV_X1 U15583 ( .A(n12320), .ZN(n13357) );
  AOI22_X1 U15584 ( .A1(n12321), .A2(n13357), .B1(n11785), .B2(n16778), .ZN(
        n12326) );
  INV_X1 U15585 ( .A(n12322), .ZN(n12324) );
  NAND3_X1 U15586 ( .A1(n12324), .A2(n12323), .A3(n11793), .ZN(n12325) );
  AND3_X1 U15587 ( .A1(n12327), .A2(n12326), .A3(n12325), .ZN(n12335) );
  NAND2_X1 U15588 ( .A1(n13885), .A2(n12339), .ZN(n12329) );
  NAND2_X1 U15589 ( .A1(n12329), .A2(n19545), .ZN(n12334) );
  INV_X1 U15590 ( .A(n12330), .ZN(n12333) );
  AND3_X1 U15591 ( .A1(n10064), .A2(n11773), .A3(n12331), .ZN(n12332) );
  NAND2_X1 U15592 ( .A1(n12333), .A2(n12332), .ZN(n13531) );
  AND3_X1 U15593 ( .A1(n12335), .A2(n12334), .A3(n13531), .ZN(n13891) );
  NAND2_X1 U15594 ( .A1(n13891), .A2(n9647), .ZN(n12336) );
  NAND2_X1 U15595 ( .A1(n12554), .A2(n12336), .ZN(n14318) );
  NAND2_X1 U15596 ( .A1(n12339), .A2(n12338), .ZN(n12340) );
  NAND2_X1 U15597 ( .A1(n12554), .A2(n13904), .ZN(n13656) );
  NAND2_X1 U15598 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16715) );
  NAND2_X1 U15599 ( .A1(n12342), .A2(n16715), .ZN(n12354) );
  OR2_X1 U15600 ( .A1(n13656), .A2(n12354), .ZN(n13669) );
  OAI21_X1 U15601 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n14318), .A(
        n13669), .ZN(n12343) );
  INV_X1 U15602 ( .A(n12343), .ZN(n12345) );
  INV_X1 U15603 ( .A(n16715), .ZN(n12353) );
  OR2_X1 U15604 ( .A1(n14318), .A2(n12353), .ZN(n12344) );
  NOR2_X1 U15605 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16754) );
  NOR2_X1 U15606 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13340) );
  NAND2_X1 U15607 ( .A1(n16754), .A2(n13340), .ZN(n16394) );
  INV_X2 U15608 ( .A(n16394), .ZN(n16434) );
  OR2_X1 U15609 ( .A1(n12554), .A2(n16434), .ZN(n16728) );
  AND2_X1 U15610 ( .A1(n12344), .A2(n16728), .ZN(n13657) );
  NAND2_X1 U15611 ( .A1(n16694), .A2(n16729), .ZN(n12572) );
  NOR3_X1 U15612 ( .A1(n14151), .A2(n14208), .A3(n14207), .ZN(n16695) );
  NAND3_X1 U15613 ( .A1(n16694), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n16695), .ZN(n12346) );
  NAND2_X1 U15614 ( .A1(n12572), .A2(n12346), .ZN(n16682) );
  INV_X1 U15615 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16674) );
  NOR2_X1 U15616 ( .A1(n16674), .A2(n16681), .ZN(n12358) );
  OR2_X1 U15617 ( .A1(n16729), .A2(n12358), .ZN(n12347) );
  NAND2_X1 U15618 ( .A1(n16682), .A2(n12347), .ZN(n16660) );
  AND2_X1 U15619 ( .A1(n16519), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12359) );
  NOR2_X1 U15620 ( .A1(n16729), .A2(n12359), .ZN(n12348) );
  NOR2_X1 U15621 ( .A1(n16660), .A2(n12348), .ZN(n16520) );
  AND2_X1 U15622 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16494) );
  OR2_X1 U15623 ( .A1(n16729), .A2(n16494), .ZN(n12349) );
  AND2_X1 U15624 ( .A1(n16520), .A2(n12349), .ZN(n16485) );
  AND3_X1 U15625 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12360) );
  OR2_X1 U15626 ( .A1(n16729), .A2(n12360), .ZN(n12350) );
  NAND2_X1 U15627 ( .A1(n16485), .A2(n12350), .ZN(n12745) );
  INV_X1 U15628 ( .A(n12570), .ZN(n12351) );
  NOR2_X1 U15629 ( .A1(n16729), .A2(n12351), .ZN(n12352) );
  OR3_X1 U15630 ( .A1(n12745), .A2(n12352), .A3(n12569), .ZN(n12573) );
  INV_X1 U15631 ( .A(n13656), .ZN(n14315) );
  AND2_X1 U15632 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12353), .ZN(
        n12355) );
  OAI21_X1 U15633 ( .B1(n14315), .B2(n12355), .A(n12354), .ZN(n12356) );
  NAND2_X1 U15634 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12357), .ZN(
        n16680) );
  INV_X1 U15635 ( .A(n12358), .ZN(n16665) );
  NOR2_X2 U15636 ( .A1(n16680), .A2(n16665), .ZN(n16655) );
  NAND2_X1 U15637 ( .A1(n16509), .A2(n16494), .ZN(n16455) );
  INV_X1 U15638 ( .A(n12360), .ZN(n12361) );
  OAI21_X1 U15639 ( .B1(n13000), .B2(n12570), .A(n12569), .ZN(n12363) );
  NAND2_X1 U15640 ( .A1(n16434), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n16172) );
  INV_X1 U15641 ( .A(n16172), .ZN(n12362) );
  AOI21_X1 U15642 ( .B1(n12573), .B2(n12363), .A(n12362), .ZN(n12364) );
  OAI21_X1 U15643 ( .B1(n16177), .B2(n16669), .A(n12364), .ZN(n12365) );
  INV_X1 U15644 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n12370) );
  NAND2_X1 U15645 ( .A1(n12543), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n12392) );
  INV_X1 U15646 ( .A(n12384), .ZN(n12378) );
  INV_X1 U15647 ( .A(n12375), .ZN(n12376) );
  MUX2_X1 U15648 ( .A(n12376), .B(P2_EBX_REG_4__SCAN_IN), .S(n12543), .Z(
        n12400) );
  INV_X1 U15649 ( .A(n12400), .ZN(n12377) );
  INV_X1 U15650 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n12380) );
  MUX2_X1 U15651 ( .A(n12380), .B(n12379), .S(n12532), .Z(n12406) );
  INV_X1 U15652 ( .A(n12381), .ZN(n12382) );
  MUX2_X1 U15653 ( .A(n21330), .B(n12382), .S(n12532), .Z(n12418) );
  XNOR2_X1 U15654 ( .A(n12414), .B(n12418), .ZN(n19407) );
  INV_X1 U15655 ( .A(n12385), .ZN(n12388) );
  INV_X1 U15656 ( .A(n12386), .ZN(n12387) );
  NAND2_X1 U15657 ( .A1(n12388), .A2(n12387), .ZN(n12389) );
  NAND2_X1 U15658 ( .A1(n12384), .A2(n12389), .ZN(n15927) );
  XNOR2_X1 U15659 ( .A(n12395), .B(n12390), .ZN(n15945) );
  XNOR2_X1 U15660 ( .A(n15945), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13664) );
  OAI21_X1 U15661 ( .B1(n12391), .B2(n12543), .A(n12392), .ZN(n15965) );
  NAND2_X1 U15662 ( .A1(n15965), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13443) );
  INV_X1 U15663 ( .A(n12392), .ZN(n12393) );
  NAND2_X1 U15664 ( .A1(n12393), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n12394) );
  AND2_X1 U15665 ( .A1(n12395), .A2(n12394), .ZN(n13442) );
  NAND2_X1 U15666 ( .A1(n13442), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12397) );
  INV_X1 U15667 ( .A(n13442), .ZN(n15954) );
  AND2_X1 U15668 ( .A1(n15954), .A2(n13440), .ZN(n12396) );
  AOI21_X1 U15669 ( .B1(n13443), .B2(n12397), .A(n12396), .ZN(n13663) );
  NAND2_X1 U15670 ( .A1(n13664), .A2(n13663), .ZN(n13662) );
  INV_X1 U15671 ( .A(n15945), .ZN(n12398) );
  NAND2_X1 U15672 ( .A1(n12398), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12399) );
  NAND2_X1 U15673 ( .A1(n13662), .A2(n12399), .ZN(n14148) );
  XNOR2_X1 U15674 ( .A(n12400), .B(n12384), .ZN(n15914) );
  NAND2_X1 U15675 ( .A1(n15914), .A2(n14207), .ZN(n12403) );
  OAI21_X1 U15676 ( .B1(n14148), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n12403), .ZN(n12401) );
  INV_X1 U15677 ( .A(n12401), .ZN(n12402) );
  NOR2_X1 U15678 ( .A1(n15914), .A2(n14207), .ZN(n12404) );
  NOR2_X1 U15679 ( .A1(n10573), .A2(n12404), .ZN(n12405) );
  XNOR2_X1 U15680 ( .A(n12407), .B(n12406), .ZN(n12408) );
  NAND2_X1 U15681 ( .A1(n12408), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12410) );
  INV_X1 U15682 ( .A(n12408), .ZN(n15898) );
  NAND2_X1 U15683 ( .A1(n15898), .A2(n14208), .ZN(n12409) );
  AND2_X1 U15684 ( .A1(n12410), .A2(n12409), .ZN(n14205) );
  MUX2_X1 U15685 ( .A(n12413), .B(n12412), .S(n12532), .Z(n12419) );
  NAND2_X1 U15686 ( .A1(n12543), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12415) );
  INV_X1 U15687 ( .A(n12415), .ZN(n12416) );
  NAND2_X1 U15688 ( .A1(n12423), .A2(n12416), .ZN(n12417) );
  NAND2_X1 U15689 ( .A1(n12434), .A2(n12417), .ZN(n15866) );
  NOR2_X1 U15690 ( .A1(n15866), .A2(n12048), .ZN(n12430) );
  NAND2_X1 U15691 ( .A1(n12430), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16405) );
  INV_X1 U15692 ( .A(n12418), .ZN(n12421) );
  INV_X1 U15693 ( .A(n12419), .ZN(n12420) );
  OAI21_X1 U15694 ( .B1(n12414), .B2(n12421), .A(n12420), .ZN(n12422) );
  AND2_X1 U15695 ( .A1(n12422), .A2(n12423), .ZN(n15886) );
  NAND2_X1 U15696 ( .A1(n15886), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16423) );
  AND2_X1 U15697 ( .A1(n16405), .A2(n16423), .ZN(n16374) );
  INV_X1 U15698 ( .A(n12427), .ZN(n12425) );
  NOR2_X1 U15699 ( .A1(n12532), .A2(n12426), .ZN(n12424) );
  AOI21_X1 U15700 ( .B1(n12425), .B2(n12424), .A(n12475), .ZN(n12428) );
  NAND2_X1 U15701 ( .A1(n12427), .A2(n12426), .ZN(n12438) );
  NAND2_X1 U15702 ( .A1(n12428), .A2(n12438), .ZN(n15842) );
  OR2_X1 U15703 ( .A1(n15842), .A2(n12048), .ZN(n12429) );
  NAND2_X1 U15704 ( .A1(n12429), .A2(n9601), .ZN(n16377) );
  INV_X1 U15705 ( .A(n12430), .ZN(n12431) );
  NAND2_X1 U15706 ( .A1(n12431), .A2(n16674), .ZN(n16404) );
  INV_X1 U15707 ( .A(n15886), .ZN(n12432) );
  NAND2_X1 U15708 ( .A1(n12432), .A2(n16681), .ZN(n16422) );
  AND2_X1 U15709 ( .A1(n16404), .A2(n16422), .ZN(n16372) );
  NAND2_X1 U15710 ( .A1(n12543), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12433) );
  XNOR2_X1 U15711 ( .A(n12434), .B(n12433), .ZN(n15861) );
  NAND2_X1 U15712 ( .A1(n15861), .A2(n12412), .ZN(n12435) );
  NAND2_X1 U15713 ( .A1(n12435), .A2(n16654), .ZN(n16390) );
  NAND2_X1 U15714 ( .A1(n12412), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12436) );
  NOR2_X1 U15715 ( .A1(n15842), .A2(n12436), .ZN(n16376) );
  AND2_X1 U15716 ( .A1(n12412), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12437) );
  INV_X1 U15717 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n12439) );
  NAND2_X1 U15718 ( .A1(n12440), .A2(n12439), .ZN(n12443) );
  INV_X2 U15719 ( .A(n12475), .ZN(n12522) );
  NAND2_X1 U15720 ( .A1(n12543), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12441) );
  INV_X1 U15721 ( .A(n12441), .ZN(n12442) );
  NAND2_X1 U15722 ( .A1(n12443), .A2(n12442), .ZN(n12444) );
  NAND2_X1 U15723 ( .A1(n12445), .A2(n12444), .ZN(n15812) );
  INV_X1 U15724 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16615) );
  NOR2_X1 U15725 ( .A1(n12470), .A2(n16615), .ZN(n16351) );
  INV_X1 U15726 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12446) );
  NOR2_X1 U15727 ( .A1(n12532), .A2(n12446), .ZN(n12471) );
  NAND2_X1 U15728 ( .A1(n12543), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12466) );
  NAND2_X1 U15729 ( .A1(n12543), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12464) );
  NAND3_X1 U15730 ( .A1(n12452), .A2(n12543), .A3(P2_EBX_REG_19__SCAN_IN), 
        .ZN(n12451) );
  NOR2_X1 U15731 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(P2_EBX_REG_18__SCAN_IN), 
        .ZN(n12450) );
  NAND2_X1 U15732 ( .A1(n15721), .A2(n12412), .ZN(n12485) );
  INV_X1 U15733 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16532) );
  NAND2_X1 U15734 ( .A1(n12485), .A2(n16532), .ZN(n16274) );
  NAND2_X1 U15735 ( .A1(n15743), .A2(n12412), .ZN(n12455) );
  NAND2_X1 U15736 ( .A1(n12455), .A2(n12454), .ZN(n16276) );
  NAND2_X1 U15737 ( .A1(n12456), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12457) );
  MUX2_X1 U15738 ( .A(n12457), .B(n12456), .S(n12532), .Z(n12458) );
  INV_X1 U15739 ( .A(n12460), .ZN(n12461) );
  NAND2_X1 U15740 ( .A1(n12458), .A2(n12461), .ZN(n15712) );
  INV_X1 U15741 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16535) );
  OAI21_X1 U15742 ( .B1(n15712), .B2(n12048), .A(n16535), .ZN(n16264) );
  NAND2_X1 U15743 ( .A1(n12460), .A2(n12459), .ZN(n12504) );
  NAND2_X1 U15744 ( .A1(n12504), .A2(n12522), .ZN(n12501) );
  AND3_X1 U15745 ( .A1(n12461), .A2(n12543), .A3(P2_EBX_REG_21__SCAN_IN), .ZN(
        n12462) );
  OR2_X1 U15746 ( .A1(n12501), .A2(n12462), .ZN(n12483) );
  OAI21_X1 U15747 ( .B1(n12483), .B2(n12048), .A(n16255), .ZN(n16252) );
  OAI21_X1 U15748 ( .B1(n12465), .B2(n12464), .A(n12463), .ZN(n15753) );
  OR2_X1 U15749 ( .A1(n15753), .A2(n12048), .ZN(n12487) );
  NAND2_X1 U15750 ( .A1(n12487), .A2(n16301), .ZN(n14325) );
  XNOR2_X1 U15751 ( .A(n9679), .B(n12466), .ZN(n15780) );
  NAND2_X1 U15752 ( .A1(n15780), .A2(n12412), .ZN(n12467) );
  INV_X1 U15753 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21336) );
  NAND2_X1 U15754 ( .A1(n12467), .A2(n21336), .ZN(n16323) );
  XNOR2_X1 U15755 ( .A(n12468), .B(n9745), .ZN(n15793) );
  NAND2_X1 U15756 ( .A1(n15793), .A2(n12412), .ZN(n12469) );
  INV_X1 U15757 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16592) );
  NAND2_X1 U15758 ( .A1(n12469), .A2(n16592), .ZN(n16330) );
  NAND2_X1 U15759 ( .A1(n12470), .A2(n16615), .ZN(n16352) );
  NAND2_X1 U15760 ( .A1(n12445), .A2(n12471), .ZN(n12472) );
  NAND2_X1 U15761 ( .A1(n12468), .A2(n12472), .ZN(n15807) );
  INV_X1 U15762 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12473) );
  OAI21_X1 U15763 ( .B1(n15807), .B2(n12048), .A(n12473), .ZN(n16340) );
  AND4_X1 U15764 ( .A1(n16323), .A2(n16330), .A3(n16352), .A4(n16340), .ZN(
        n12474) );
  AND2_X1 U15765 ( .A1(n14325), .A2(n12474), .ZN(n12480) );
  NOR2_X1 U15766 ( .A1(n12532), .A2(n12449), .ZN(n12476) );
  AOI21_X1 U15767 ( .B1(n12477), .B2(n12476), .A(n12475), .ZN(n12479) );
  NAND2_X1 U15768 ( .A1(n12479), .A2(n12478), .ZN(n15768) );
  XNOR2_X1 U15769 ( .A(n12488), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16307) );
  AND2_X1 U15770 ( .A1(n16252), .A2(n10565), .ZN(n12481) );
  OR2_X1 U15771 ( .A1(n12482), .A2(n12048), .ZN(n16362) );
  INV_X1 U15772 ( .A(n12483), .ZN(n15698) );
  AND2_X1 U15773 ( .A1(n12412), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12484) );
  NAND2_X1 U15774 ( .A1(n15698), .A2(n12484), .ZN(n16251) );
  INV_X1 U15775 ( .A(n12485), .ZN(n12486) );
  NAND2_X1 U15776 ( .A1(n12486), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16275) );
  NOR2_X1 U15777 ( .A1(n12487), .A2(n16301), .ZN(n16246) );
  INV_X1 U15778 ( .A(n12488), .ZN(n12489) );
  NAND2_X1 U15779 ( .A1(n12489), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14330) );
  INV_X1 U15780 ( .A(n15780), .ZN(n12490) );
  INV_X1 U15781 ( .A(n15807), .ZN(n12492) );
  AND2_X1 U15782 ( .A1(n12412), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12491) );
  NAND2_X1 U15783 ( .A1(n12492), .A2(n12491), .ZN(n16339) );
  AND2_X1 U15784 ( .A1(n12412), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12493) );
  NAND2_X1 U15785 ( .A1(n15793), .A2(n12493), .ZN(n16329) );
  NAND4_X1 U15786 ( .A1(n14330), .A2(n16322), .A3(n16339), .A4(n16329), .ZN(
        n12494) );
  NOR2_X1 U15787 ( .A1(n16246), .A2(n12494), .ZN(n12495) );
  AND2_X1 U15788 ( .A1(n16275), .A2(n12495), .ZN(n12499) );
  INV_X1 U15789 ( .A(n15712), .ZN(n12497) );
  AND2_X1 U15790 ( .A1(n12412), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12496) );
  NAND2_X1 U15791 ( .A1(n12497), .A2(n12496), .ZN(n16263) );
  AND2_X1 U15792 ( .A1(n12412), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12498) );
  NAND2_X1 U15793 ( .A1(n15743), .A2(n12498), .ZN(n16283) );
  NAND2_X1 U15794 ( .A1(n12543), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12502) );
  NAND2_X1 U15795 ( .A1(n12501), .A2(n12502), .ZN(n12509) );
  INV_X1 U15796 ( .A(n12502), .ZN(n12503) );
  NAND2_X1 U15797 ( .A1(n12504), .A2(n12503), .ZN(n12505) );
  NAND2_X1 U15798 ( .A1(n12509), .A2(n12505), .ZN(n16839) );
  OR2_X1 U15799 ( .A1(n16839), .A2(n12048), .ZN(n12506) );
  NAND2_X1 U15800 ( .A1(n12506), .A2(n12507), .ZN(n16239) );
  OR3_X1 U15801 ( .A1(n16839), .A2(n12048), .A3(n12507), .ZN(n16238) );
  INV_X1 U15802 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12508) );
  NOR2_X1 U15803 ( .A1(n12532), .A2(n12508), .ZN(n12510) );
  NOR2_X2 U15804 ( .A1(n12509), .A2(n12510), .ZN(n12517) );
  NAND2_X1 U15805 ( .A1(n12509), .A2(n12510), .ZN(n12511) );
  NAND2_X1 U15806 ( .A1(n15664), .A2(n12511), .ZN(n15682) );
  OR2_X1 U15807 ( .A1(n15682), .A2(n12048), .ZN(n12512) );
  XNOR2_X1 U15808 ( .A(n12512), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16230) );
  NAND2_X1 U15809 ( .A1(n12412), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12513) );
  OR2_X1 U15810 ( .A1(n15682), .A2(n12513), .ZN(n12514) );
  NAND2_X1 U15811 ( .A1(n12522), .A2(n12412), .ZN(n16220) );
  INV_X1 U15812 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n15999) );
  INV_X1 U15813 ( .A(n12584), .ZN(n12519) );
  NAND3_X1 U15814 ( .A1(n9664), .A2(n12543), .A3(P2_EBX_REG_26__SCAN_IN), .ZN(
        n12518) );
  XNOR2_X1 U15815 ( .A(n12520), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16205) );
  NAND2_X1 U15816 ( .A1(n12543), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12521) );
  NAND3_X1 U15817 ( .A1(n12523), .A2(n9664), .A3(n12522), .ZN(n15642) );
  OR2_X1 U15818 ( .A1(n15642), .A2(n12048), .ZN(n12524) );
  NAND2_X1 U15819 ( .A1(n12524), .A2(n16471), .ZN(n16211) );
  NAND2_X1 U15820 ( .A1(n16220), .A2(n16484), .ZN(n12525) );
  NAND2_X1 U15821 ( .A1(n12543), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12527) );
  INV_X1 U15822 ( .A(n12527), .ZN(n12528) );
  NAND2_X1 U15823 ( .A1(n12529), .A2(n12528), .ZN(n12530) );
  NAND2_X1 U15824 ( .A1(n12534), .A2(n12530), .ZN(n15616) );
  INV_X1 U15825 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12738) );
  AND2_X1 U15826 ( .A1(n16192), .A2(n12738), .ZN(n12537) );
  NOR2_X1 U15827 ( .A1(n12532), .A2(n12531), .ZN(n12533) );
  NAND2_X1 U15828 ( .A1(n12534), .A2(n12533), .ZN(n12535) );
  NAND2_X1 U15829 ( .A1(n12547), .A2(n12535), .ZN(n15601) );
  NOR2_X1 U15830 ( .A1(n15601), .A2(n12048), .ZN(n16196) );
  OAI21_X1 U15831 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n16196), .ZN(n12536) );
  INV_X1 U15832 ( .A(n16196), .ZN(n12538) );
  INV_X1 U15833 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12998) );
  NAND2_X1 U15834 ( .A1(n12538), .A2(n12998), .ZN(n12542) );
  NAND2_X1 U15835 ( .A1(n12412), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12540) );
  NAND2_X1 U15836 ( .A1(n12412), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12539) );
  OAI21_X1 U15837 ( .B1(n12541), .B2(n12540), .A(n16210), .ZN(n12742) );
  NAND2_X1 U15838 ( .A1(n12543), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12545) );
  XNOR2_X1 U15839 ( .A(n12547), .B(n12545), .ZN(n15581) );
  AOI21_X1 U15840 ( .B1(n15581), .B2(n12412), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12992) );
  AND2_X1 U15841 ( .A1(n12412), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12544) );
  NOR2_X1 U15842 ( .A1(n12582), .A2(n12991), .ZN(n12553) );
  INV_X1 U15843 ( .A(n12545), .ZN(n12546) );
  INV_X1 U15844 ( .A(n12583), .ZN(n12549) );
  NOR2_X1 U15845 ( .A1(n12532), .A2(n14632), .ZN(n12548) );
  OAI21_X1 U15846 ( .B1(n12550), .B2(n12048), .A(n12569), .ZN(n12581) );
  INV_X1 U15847 ( .A(n12581), .ZN(n12551) );
  INV_X1 U15848 ( .A(n12550), .ZN(n13060) );
  NOR2_X1 U15849 ( .A1(n12551), .A2(n12579), .ZN(n12552) );
  XNOR2_X1 U15850 ( .A(n12553), .B(n12552), .ZN(n16179) );
  AND2_X1 U15851 ( .A1(n13913), .A2(n11780), .ZN(n20276) );
  OAI211_X1 U15852 ( .C1(n16706), .C2(n16181), .A(n12556), .B(n12555), .ZN(
        P2_U3016) );
  INV_X1 U15853 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12557) );
  AOI222_X1 U15854 ( .A1(n12003), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12045), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), 
        .C2(n12559), .ZN(n12560) );
  INV_X1 U15855 ( .A(n12560), .ZN(n12561) );
  AOI22_X1 U15856 ( .A1(n12563), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12565) );
  OAI211_X1 U15857 ( .C1(n12218), .C2(n10065), .A(n12565), .B(n12564), .ZN(
        n12566) );
  INV_X1 U15858 ( .A(n12566), .ZN(n12567) );
  NOR4_X1 U15859 ( .A1(n13000), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12570), .A4(n12569), .ZN(n12571) );
  AND2_X1 U15860 ( .A1(n16434), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14343) );
  NOR2_X1 U15861 ( .A1(n12571), .A2(n14343), .ZN(n12575) );
  NAND3_X1 U15862 ( .A1(n12573), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12572), .ZN(n12574) );
  OAI211_X1 U15863 ( .C1(n14357), .C2(n16669), .A(n12575), .B(n12574), .ZN(
        n12576) );
  INV_X1 U15864 ( .A(n12576), .ZN(n12577) );
  MUX2_X1 U15865 ( .A(n12585), .B(n12584), .S(n12532), .Z(n14360) );
  NAND2_X1 U15866 ( .A1(n14348), .A2(n16689), .ZN(n12588) );
  OAI211_X1 U15867 ( .C1(n14349), .C2(n16706), .A(n12589), .B(n12588), .ZN(
        P2_U3015) );
  NAND2_X1 U15868 ( .A1(n18323), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18314) );
  NAND2_X1 U15869 ( .A1(n18286), .A2(n18252), .ZN(n18217) );
  NAND2_X1 U15870 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18222) );
  NAND2_X1 U15871 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18181) );
  NAND2_X1 U15872 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18149) );
  NOR2_X2 U15873 ( .A1(n12602), .A2(n18149), .ZN(n18135) );
  NAND2_X1 U15874 ( .A1(n18135), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n18108) );
  NAND2_X1 U15875 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18113) );
  NAND2_X1 U15876 ( .A1(n12600), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12597) );
  NAND2_X1 U15877 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18076) );
  NOR2_X4 U15878 ( .A1(n12597), .A2(n18076), .ZN(n18054) );
  XOR2_X1 U15879 ( .A(n12612), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n17009) );
  INV_X1 U15880 ( .A(n12591), .ZN(n12594) );
  INV_X1 U15881 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17147) );
  NOR2_X1 U15882 ( .A1(n12594), .A2(n17147), .ZN(n12593) );
  OAI21_X1 U15883 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n12593), .A(
        n12592), .ZN(n12920) );
  INV_X1 U15884 ( .A(n12920), .ZN(n17138) );
  AOI21_X1 U15885 ( .B1(n12594), .B2(n17147), .A(n12593), .ZN(n18044) );
  AOI21_X1 U15886 ( .B1(n12595), .B2(n12596), .A(n12591), .ZN(n18059) );
  NOR2_X1 U15887 ( .A1(n17477), .A2(n12597), .ZN(n12610) );
  AND2_X1 U15888 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n12610), .ZN(
        n12598) );
  OAI21_X1 U15889 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n12598), .A(
        n12595), .ZN(n12599) );
  INV_X1 U15890 ( .A(n12599), .ZN(n18067) );
  INV_X1 U15891 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12601) );
  NAND2_X1 U15892 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n12600), .ZN(
        n18091) );
  AOI21_X1 U15893 ( .B1(n12601), .B2(n18091), .A(n12610), .ZN(n18095) );
  INV_X1 U15894 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17202) );
  INV_X1 U15895 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17221) );
  NOR2_X1 U15896 ( .A1(n17477), .A2(n12602), .ZN(n18148) );
  INV_X1 U15897 ( .A(n18148), .ZN(n12603) );
  NOR2_X1 U15898 ( .A1(n18149), .A2(n12603), .ZN(n17229) );
  INV_X1 U15899 ( .A(n17229), .ZN(n18111) );
  NOR2_X1 U15900 ( .A1(n17221), .A2(n18111), .ZN(n12608) );
  NAND2_X1 U15901 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12608), .ZN(
        n12604) );
  INV_X1 U15902 ( .A(n18091), .ZN(n18065) );
  AOI21_X1 U15903 ( .B1(n17202), .B2(n12604), .A(n18065), .ZN(n18112) );
  XOR2_X1 U15904 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n12608), .Z(
        n18124) );
  NAND2_X1 U15905 ( .A1(n12612), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12606) );
  XNOR2_X2 U15906 ( .A(n12606), .B(n12605), .ZN(n10319) );
  NAND2_X1 U15907 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18148), .ZN(
        n17241) );
  NOR2_X1 U15908 ( .A1(n17477), .A2(n12607), .ZN(n18180) );
  NAND2_X1 U15909 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18180), .ZN(
        n17276) );
  NOR2_X1 U15910 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17276), .ZN(
        n17275) );
  NOR2_X1 U15911 ( .A1(n17275), .A2(n10319), .ZN(n17266) );
  OAI21_X1 U15912 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17434), .A(
        n17243), .ZN(n17219) );
  AOI21_X1 U15913 ( .B1(n17221), .B2(n18111), .A(n12608), .ZN(n18139) );
  OR2_X2 U15914 ( .A1(n17219), .A2(n18139), .ZN(n17217) );
  NOR2_X1 U15915 ( .A1(n17198), .A2(n17434), .ZN(n17189) );
  XOR2_X1 U15916 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n12610), .Z(
        n18081) );
  INV_X1 U15917 ( .A(n18081), .ZN(n12611) );
  NOR2_X2 U15918 ( .A1(n18067), .A2(n17166), .ZN(n17165) );
  NOR2_X1 U15919 ( .A1(n17165), .A2(n17434), .ZN(n17156) );
  NOR2_X1 U15921 ( .A1(n17155), .A2(n17434), .ZN(n17146) );
  AOI21_X1 U15922 ( .B1(n12592), .B2(n17121), .A(n12612), .ZN(n17118) );
  NOR2_X1 U15923 ( .A1(n17120), .A2(n10319), .ZN(n13265) );
  NOR3_X1 U15924 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n19222) );
  NAND2_X1 U15925 ( .A1(n10321), .A2(n19216), .ZN(n17472) );
  NOR3_X1 U15926 ( .A1(n17009), .A2(n13265), .A3(n17472), .ZN(n12737) );
  INV_X1 U15927 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19240) );
  NOR2_X1 U15928 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n19224) );
  INV_X2 U15929 ( .A(n17563), .ZN(n17701) );
  AOI22_X1 U15930 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12616) );
  AOI22_X1 U15931 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14270), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12615) );
  AOI22_X1 U15932 ( .A1(n12812), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12614) );
  AOI22_X1 U15933 ( .A1(n17734), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12613) );
  NAND4_X1 U15934 ( .A1(n12616), .A2(n12615), .A3(n12614), .A4(n12613), .ZN(
        n12626) );
  INV_X4 U15935 ( .A(n17578), .ZN(n17721) );
  AOI22_X1 U15936 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17738), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12624) );
  AOI22_X1 U15937 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12623) );
  AOI22_X1 U15938 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12622) );
  INV_X2 U15939 ( .A(n12784), .ZN(n17720) );
  AOI22_X1 U15940 ( .A1(n17720), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12621) );
  NAND4_X1 U15941 ( .A1(n12624), .A2(n12623), .A3(n12622), .A4(n12621), .ZN(
        n12625) );
  OAI211_X1 U15942 ( .C1(n19228), .C2(n17972), .A(n19361), .B(n19359), .ZN(
        n12727) );
  AOI22_X1 U15943 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U15944 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17738), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12630) );
  INV_X2 U15945 ( .A(n17489), .ZN(n17737) );
  AOI22_X1 U15946 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12629) );
  AOI22_X1 U15947 ( .A1(n17676), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12628) );
  NAND4_X1 U15948 ( .A1(n12631), .A2(n12630), .A3(n12629), .A4(n12628), .ZN(
        n12637) );
  AOI22_X1 U15949 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12812), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12635) );
  AOI22_X1 U15950 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12836), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12634) );
  AOI22_X1 U15951 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12843), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12633) );
  AOI22_X1 U15952 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12632) );
  NAND4_X1 U15953 ( .A1(n12635), .A2(n12634), .A3(n12633), .A4(n12632), .ZN(
        n12636) );
  AOI22_X1 U15954 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17643), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17676), .ZN(n12646) );
  AOI22_X1 U15955 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17720), .ZN(n12645) );
  AOI22_X1 U15956 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n14305), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17733), .ZN(n12638) );
  OAI21_X1 U15957 ( .B1(n12822), .B2(n21273), .A(n12638), .ZN(n12644) );
  AOI22_X1 U15958 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12836), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12643) );
  AOI22_X1 U15959 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9611), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12642) );
  AOI22_X1 U15960 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17719), .ZN(n12641) );
  INV_X1 U15961 ( .A(n9628), .ZN(n17700) );
  AOI22_X1 U15962 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n9628), .B1(
        n12812), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12640) );
  NAND2_X1 U15963 ( .A1(n18721), .A2(n17826), .ZN(n12698) );
  AOI22_X1 U15964 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12656) );
  AOI22_X1 U15965 ( .A1(n12812), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12647) );
  OAI21_X1 U15966 ( .B1(n17489), .B2(n21222), .A(n12647), .ZN(n12653) );
  AOI22_X1 U15967 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12651) );
  AOI22_X1 U15968 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12836), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12650) );
  AOI22_X1 U15969 ( .A1(n17714), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12649) );
  AOI22_X1 U15970 ( .A1(n17720), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12648) );
  NAND4_X1 U15971 ( .A1(n12651), .A2(n12650), .A3(n12649), .A4(n12648), .ZN(
        n12652) );
  AOI211_X1 U15972 ( .C1(n9597), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n12653), .B(n12652), .ZN(n12654) );
  AOI22_X1 U15973 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12666) );
  AOI22_X1 U15974 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12843), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12657) );
  OAI21_X1 U15975 ( .B1(n17736), .B2(n17774), .A(n12657), .ZN(n12663) );
  AOI22_X1 U15976 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17738), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12661) );
  AOI22_X1 U15977 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12660) );
  AOI22_X1 U15978 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17734), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12659) );
  AOI22_X1 U15979 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12658) );
  NAND4_X1 U15980 ( .A1(n12661), .A2(n12660), .A3(n12659), .A4(n12658), .ZN(
        n12662) );
  AOI22_X1 U15981 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12670) );
  AOI22_X1 U15982 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12836), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12669) );
  AOI22_X1 U15983 ( .A1(n17714), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16791), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12668) );
  AOI22_X1 U15984 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12667) );
  NAND4_X1 U15985 ( .A1(n12670), .A2(n12669), .A3(n12668), .A4(n12667), .ZN(
        n12676) );
  AOI22_X1 U15986 ( .A1(n12812), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12674) );
  AOI22_X1 U15987 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12673) );
  AOI22_X1 U15988 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12672) );
  AOI22_X1 U15989 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12671) );
  NAND4_X1 U15990 ( .A1(n12674), .A2(n12673), .A3(n12672), .A4(n12671), .ZN(
        n12675) );
  AOI22_X1 U15991 ( .A1(n17714), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12687) );
  AOI22_X1 U15992 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12686) );
  AOI22_X1 U15993 ( .A1(n12812), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12836), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12677) );
  OAI21_X1 U15994 ( .B1(n12678), .B2(n21256), .A(n12677), .ZN(n12684) );
  AOI22_X1 U15995 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12682) );
  AOI22_X1 U15996 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12681) );
  AOI22_X1 U15997 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12680) );
  AOI22_X1 U15998 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16791), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12679) );
  NAND4_X1 U15999 ( .A1(n12682), .A2(n12681), .A3(n12680), .A4(n12679), .ZN(
        n12683) );
  NOR2_X1 U16000 ( .A1(n17785), .A2(n18745), .ZN(n12884) );
  NOR2_X1 U16001 ( .A1(n12698), .A2(n14223), .ZN(n12695) );
  AOI22_X1 U16002 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17734), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12694) );
  AOI22_X1 U16003 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12693) );
  AOI22_X1 U16004 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12691) );
  AOI22_X1 U16005 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17738), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12690) );
  AOI22_X1 U16006 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16791), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12689) );
  AOI22_X1 U16007 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12688) );
  NAND4_X1 U16008 ( .A1(n12691), .A2(n12690), .A3(n12689), .A4(n12688), .ZN(
        n12692) );
  NAND3_X1 U16009 ( .A1(n12694), .A2(n12693), .A3(n9728), .ZN(n14224) );
  NOR2_X1 U16010 ( .A1(n19360), .A2(n17424), .ZN(n12879) );
  NAND2_X1 U16011 ( .A1(n18745), .A2(n18749), .ZN(n12701) );
  NOR4_X2 U16012 ( .A1(n18736), .A2(n14224), .A3(n12698), .A4(n12701), .ZN(
        n12707) );
  NAND2_X1 U16013 ( .A1(n12707), .A2(n18732), .ZN(n12953) );
  NAND2_X1 U16014 ( .A1(n17973), .A2(n12953), .ZN(n17103) );
  NAND2_X1 U16015 ( .A1(n12879), .A2(n17103), .ZN(n12876) );
  INV_X1 U16016 ( .A(n19167), .ZN(n19170) );
  NOR2_X1 U16017 ( .A1(n18721), .A2(n17972), .ZN(n12878) );
  OAI21_X1 U16018 ( .B1(n12696), .B2(n19183), .A(n12878), .ZN(n12956) );
  OAI21_X1 U16019 ( .B1(n12951), .B2(n12702), .A(n12956), .ZN(n12706) );
  INV_X1 U16020 ( .A(n14224), .ZN(n18742) );
  AOI22_X1 U16021 ( .A1(n12699), .A2(n12698), .B1(n18742), .B2(n19183), .ZN(
        n12705) );
  OR2_X1 U16022 ( .A1(n18732), .A2(n12879), .ZN(n12888) );
  AOI21_X1 U16023 ( .B1(n17826), .B2(n12701), .A(n18742), .ZN(n12700) );
  AOI21_X1 U16024 ( .B1(n12701), .B2(n12888), .A(n12700), .ZN(n12704) );
  AND2_X1 U16025 ( .A1(n18749), .A2(n12951), .ZN(n12960) );
  OAI21_X1 U16026 ( .B1(n12702), .B2(n12960), .A(n18721), .ZN(n12703) );
  NAND3_X1 U16027 ( .A1(n12705), .A2(n12704), .A3(n12703), .ZN(n12954) );
  NAND2_X1 U16028 ( .A1(n12707), .A2(n12877), .ZN(n12880) );
  INV_X1 U16029 ( .A(n12880), .ZN(n12708) );
  XNOR2_X1 U16030 ( .A(n12871), .B(n12873), .ZN(n12721) );
  NOR2_X1 U16031 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19197), .ZN(
        n12714) );
  NAND2_X1 U16032 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12713), .ZN(
        n12719) );
  AOI22_X1 U16033 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12718), .B1(
        n12714), .B2(n12719), .ZN(n12872) );
  NAND2_X1 U16034 ( .A1(n12717), .A2(n12716), .ZN(n12715) );
  AOI21_X1 U16035 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12719), .A(
        n12718), .ZN(n12720) );
  INV_X1 U16036 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19284) );
  INV_X1 U16037 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19279) );
  INV_X1 U16038 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19277) );
  INV_X1 U16039 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19270) );
  INV_X1 U16040 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19263) );
  INV_X1 U16041 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19254) );
  INV_X1 U16042 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19249) );
  INV_X1 U16043 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19244) );
  NAND2_X1 U16044 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17461) );
  NOR2_X1 U16045 ( .A1(n19244), .A2(n17461), .ZN(n17423) );
  NAND3_X1 U16046 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .A3(n17423), .ZN(n17382) );
  NOR2_X1 U16047 ( .A1(n19249), .A2(n17382), .ZN(n17384) );
  NAND2_X1 U16048 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n17384), .ZN(n17373) );
  NOR2_X1 U16049 ( .A1(n19254), .A2(n17373), .ZN(n17341) );
  NAND4_X1 U16050 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n17341), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n17301) );
  NOR2_X1 U16051 ( .A1(n19260), .A2(n17301), .ZN(n17302) );
  NAND2_X1 U16052 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17302), .ZN(n17293) );
  NOR2_X1 U16053 ( .A1(n19263), .A2(n17293), .ZN(n17270) );
  NAND3_X1 U16054 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(n17270), .ZN(n17254) );
  NAND4_X1 U16055 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n17228), .A3(
        P3_REIP_REG_19__SCAN_IN), .A4(P3_REIP_REG_18__SCAN_IN), .ZN(n17200) );
  NOR3_X1 U16056 ( .A1(n19279), .A2(n19277), .A3(n17200), .ZN(n17185) );
  NAND2_X1 U16057 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n17185), .ZN(n17183) );
  INV_X1 U16058 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19287) );
  INV_X1 U16059 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19285) );
  NOR2_X1 U16060 ( .A1(n19287), .A2(n19285), .ZN(n12722) );
  NAND2_X1 U16061 ( .A1(n17169), .A2(n12722), .ZN(n17153) );
  INV_X1 U16062 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19291) );
  INV_X1 U16063 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19289) );
  NOR2_X1 U16064 ( .A1(n19291), .A2(n19289), .ZN(n17134) );
  NAND3_X1 U16065 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17142), .A3(n17134), 
        .ZN(n12728) );
  NOR2_X1 U16066 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n12728), .ZN(n13267) );
  INV_X1 U16067 ( .A(n13267), .ZN(n12726) );
  NAND2_X1 U16068 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17134), .ZN(n12725) );
  INV_X1 U16069 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19214) );
  NOR2_X2 U16070 ( .A1(n19335), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19091) );
  NAND2_X1 U16071 ( .A1(n19214), .A2(n19091), .ZN(n19208) );
  INV_X1 U16072 ( .A(n19208), .ZN(n19204) );
  AOI211_X1 U16073 ( .C1(P3_STATE2_REG_0__SCAN_IN), .C2(n19204), .A(n19216), 
        .B(n18695), .ZN(n12723) );
  INV_X1 U16074 ( .A(n19357), .ZN(n19372) );
  NOR2_X1 U16075 ( .A1(n17468), .A2(n12724), .ZN(n17163) );
  NAND3_X1 U16076 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n17163), .ZN(n17133) );
  NAND2_X1 U16077 ( .A1(n17474), .A2(n17485), .ZN(n17483) );
  OAI21_X1 U16078 ( .B1(n12725), .B2(n17133), .A(n17483), .ZN(n17132) );
  INV_X1 U16079 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19297) );
  AOI21_X1 U16080 ( .B1(n12726), .B2(n17132), .A(n19297), .ZN(n12736) );
  INV_X1 U16081 ( .A(n12727), .ZN(n19206) );
  AOI211_X4 U16082 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n17972), .A(n19206), .B(
        n12731), .ZN(n17408) );
  INV_X1 U16083 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19299) );
  NOR3_X1 U16084 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19299), .A3(n12728), 
        .ZN(n12729) );
  AOI21_X1 U16085 ( .B1(n17408), .B2(P3_EBX_REG_31__SCAN_IN), .A(n12729), .ZN(
        n12734) );
  NAND2_X1 U16086 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n17972), .ZN(n12730) );
  AOI211_X4 U16087 ( .C1(n19359), .C2(n19361), .A(n12731), .B(n12730), .ZN(
        n17470) );
  NOR3_X1 U16088 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17448) );
  NAND2_X1 U16089 ( .A1(n17448), .A2(n17444), .ZN(n17443) );
  NOR2_X2 U16090 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17443), .ZN(n17419) );
  NAND2_X1 U16091 ( .A1(n17419), .A2(n17410), .ZN(n17409) );
  NOR2_X2 U16092 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17409), .ZN(n17392) );
  INV_X1 U16093 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17386) );
  NAND2_X1 U16094 ( .A1(n17392), .A2(n17386), .ZN(n17385) );
  NOR2_X2 U16095 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17385), .ZN(n17358) );
  NAND2_X1 U16096 ( .A1(n17358), .A2(n17361), .ZN(n17343) );
  INV_X1 U16097 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17337) );
  NAND2_X1 U16098 ( .A1(n17342), .A2(n17337), .ZN(n17336) );
  INV_X1 U16099 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17308) );
  NAND2_X1 U16100 ( .A1(n17314), .A2(n17308), .ZN(n17307) );
  NOR2_X2 U16101 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17307), .ZN(n17288) );
  INV_X1 U16102 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17279) );
  NAND2_X1 U16103 ( .A1(n17288), .A2(n17279), .ZN(n17278) );
  NOR2_X2 U16104 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17278), .ZN(n17267) );
  NAND2_X1 U16105 ( .A1(n17267), .A2(n17263), .ZN(n17262) );
  NAND2_X1 U16106 ( .A1(n17244), .A2(n17237), .ZN(n17236) );
  INV_X1 U16107 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17576) );
  NAND2_X1 U16108 ( .A1(n17220), .A2(n17576), .ZN(n17213) );
  NOR2_X2 U16109 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17213), .ZN(n17197) );
  INV_X1 U16110 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17186) );
  NAND2_X1 U16111 ( .A1(n17197), .A2(n17186), .ZN(n17192) );
  NOR2_X2 U16112 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17192), .ZN(n17175) );
  INV_X1 U16113 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17171) );
  NAND2_X1 U16114 ( .A1(n17175), .A2(n17171), .ZN(n17170) );
  NOR2_X2 U16115 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17170), .ZN(n17154) );
  INV_X1 U16116 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17528) );
  NAND2_X1 U16117 ( .A1(n17154), .A2(n17528), .ZN(n17150) );
  INV_X1 U16118 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17515) );
  NAND2_X1 U16119 ( .A1(n17135), .A2(n17515), .ZN(n13269) );
  NOR2_X1 U16120 ( .A1(n17481), .A2(n13269), .ZN(n13266) );
  INV_X1 U16121 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n12732) );
  NAND2_X1 U16122 ( .A1(n13266), .A2(n12732), .ZN(n12733) );
  NAND3_X1 U16123 ( .A1(n12734), .A2(n12733), .A3(n10577), .ZN(n12735) );
  AOI21_X1 U16124 ( .B1(n12743), .B2(n15624), .A(n15597), .ZN(n15619) );
  INV_X1 U16125 ( .A(n15619), .ZN(n15990) );
  NAND2_X1 U16126 ( .A1(n16434), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n13020) );
  INV_X1 U16127 ( .A(n13000), .ZN(n13003) );
  NOR2_X1 U16128 ( .A1(n13000), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12744) );
  OR2_X1 U16129 ( .A1(n12745), .A2(n12744), .ZN(n16448) );
  OAI21_X1 U16130 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13003), .A(
        n16448), .ZN(n12746) );
  OAI211_X1 U16131 ( .C1(n15990), .C2(n16669), .A(n13020), .B(n12746), .ZN(
        n12750) );
  INV_X1 U16132 ( .A(n12747), .ZN(n12749) );
  INV_X1 U16133 ( .A(n15631), .ZN(n12748) );
  AOI21_X1 U16134 ( .B1(n12749), .B2(n12748), .A(n15594), .ZN(n16081) );
  AOI22_X1 U16135 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17684), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12762) );
  AOI22_X1 U16136 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17721), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12761) );
  AOI22_X1 U16137 ( .A1(n17733), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12753) );
  OAI21_X1 U16138 ( .B1(n21273), .B2(n17700), .A(n12753), .ZN(n12759) );
  AOI22_X1 U16139 ( .A1(n17714), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12757) );
  AOI22_X1 U16140 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9611), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U16141 ( .A1(n17734), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14305), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U16142 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12754) );
  NAND4_X1 U16143 ( .A1(n12757), .A2(n12756), .A3(n12755), .A4(n12754), .ZN(
        n12758) );
  AOI211_X1 U16144 ( .C1(n17720), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n12759), .B(n12758), .ZN(n12760) );
  AOI22_X1 U16145 ( .A1(n17676), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12766) );
  AOI22_X1 U16146 ( .A1(n17738), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17734), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12765) );
  AOI22_X1 U16147 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12764) );
  AOI22_X1 U16148 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12763) );
  NAND4_X1 U16149 ( .A1(n12766), .A2(n12765), .A3(n12764), .A4(n12763), .ZN(
        n12772) );
  AOI22_X1 U16150 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12812), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12770) );
  AOI22_X1 U16151 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16791), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U16152 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12768) );
  AOI22_X1 U16153 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12767) );
  NAND4_X1 U16154 ( .A1(n12770), .A2(n12769), .A3(n12768), .A4(n12767), .ZN(
        n12771) );
  AOI22_X1 U16155 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12776) );
  AOI22_X1 U16156 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14305), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12775) );
  AOI22_X1 U16157 ( .A1(n12752), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12774) );
  AOI22_X1 U16158 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16791), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12773) );
  NAND4_X1 U16159 ( .A1(n12776), .A2(n12775), .A3(n12774), .A4(n12773), .ZN(
        n12782) );
  AOI22_X1 U16160 ( .A1(n17738), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12780) );
  AOI22_X1 U16161 ( .A1(n12842), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12836), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12779) );
  AOI22_X1 U16162 ( .A1(n12812), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12778) );
  AOI22_X1 U16163 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12777) );
  NAND4_X1 U16164 ( .A1(n12780), .A2(n12779), .A3(n12778), .A4(n12777), .ZN(
        n12781) );
  INV_X1 U16165 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n21308) );
  AOI22_X1 U16166 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n9595), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12783) );
  OAI21_X1 U16167 ( .B1(n12784), .B2(n21308), .A(n12783), .ZN(n12792) );
  AOI22_X1 U16168 ( .A1(n12812), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12785), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12790) );
  AOI22_X1 U16169 ( .A1(n12787), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12786), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12789) );
  NAND3_X1 U16170 ( .A1(n12790), .A2(n12789), .A3(n12788), .ZN(n12791) );
  AOI22_X1 U16171 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14305), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12796) );
  AOI22_X1 U16172 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12843), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12795) );
  AOI22_X1 U16173 ( .A1(n12752), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12794) );
  AOI22_X1 U16174 ( .A1(n9628), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12793) );
  AOI22_X1 U16175 ( .A1(n12752), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12801) );
  AOI22_X1 U16176 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12843), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12800) );
  AOI22_X1 U16177 ( .A1(n12842), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9597), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12799) );
  AOI22_X1 U16178 ( .A1(n17676), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12798) );
  AOI22_X1 U16179 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12802), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12804) );
  OAI21_X1 U16180 ( .B1(n12822), .B2(n17774), .A(n12804), .ZN(n12805) );
  INV_X1 U16181 ( .A(n12805), .ZN(n12809) );
  AOI22_X1 U16182 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12808) );
  AOI22_X1 U16183 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14305), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12807) );
  AOI22_X1 U16184 ( .A1(n12752), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12843), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12820) );
  AOI22_X1 U16185 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14305), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12819) );
  AOI22_X1 U16186 ( .A1(n12836), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12811) );
  OAI21_X1 U16187 ( .B1(n12822), .B2(n17763), .A(n12811), .ZN(n12818) );
  AOI22_X1 U16188 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14270), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12817) );
  AOI22_X1 U16189 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16791), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12816) );
  AOI22_X1 U16190 ( .A1(n12812), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12815) );
  AOI22_X1 U16191 ( .A1(n17676), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12814) );
  NAND2_X1 U16192 ( .A1(n12854), .A2(n12891), .ZN(n12856) );
  NOR2_X1 U16193 ( .A1(n17909), .A2(n12856), .ZN(n12860) );
  AOI22_X1 U16194 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12843), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12831) );
  AOI22_X1 U16195 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14270), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12830) );
  INV_X1 U16196 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17755) );
  AOI22_X1 U16197 ( .A1(n17734), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12821) );
  OAI21_X1 U16198 ( .B1(n12822), .B2(n17755), .A(n12821), .ZN(n12828) );
  AOI22_X1 U16199 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12826) );
  AOI22_X1 U16200 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14305), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12825) );
  AOI22_X1 U16201 ( .A1(n12812), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12824) );
  AOI22_X1 U16202 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16791), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12823) );
  NAND4_X1 U16203 ( .A1(n12826), .A2(n12825), .A3(n12824), .A4(n12823), .ZN(
        n12827) );
  AOI211_X1 U16204 ( .C1(n17737), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n12828), .B(n12827), .ZN(n12829) );
  NAND3_X1 U16205 ( .A1(n12831), .A2(n12830), .A3(n12829), .ZN(n12892) );
  NOR2_X1 U16206 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18228), .ZN(
        n12832) );
  AOI21_X1 U16207 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18228), .A(
        n12832), .ZN(n13038) );
  INV_X1 U16208 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n21267) );
  AOI22_X1 U16209 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12834) );
  OAI21_X1 U16210 ( .B1(n12835), .B2(n21267), .A(n12834), .ZN(n12841) );
  AOI22_X1 U16211 ( .A1(n12836), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14305), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12839) );
  AOI22_X1 U16212 ( .A1(n12812), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12838) );
  NAND3_X1 U16213 ( .A1(n12839), .A2(n12838), .A3(n12837), .ZN(n12840) );
  NOR2_X1 U16214 ( .A1(n12841), .A2(n12840), .ZN(n12849) );
  AOI22_X1 U16215 ( .A1(n12842), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12847) );
  AOI22_X1 U16216 ( .A1(n12785), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12802), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12846) );
  AOI22_X1 U16217 ( .A1(n12752), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12843), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12845) );
  AOI22_X1 U16218 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12844) );
  INV_X1 U16219 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19320) );
  XNOR2_X1 U16220 ( .A(n12854), .B(n17912), .ZN(n12855) );
  XNOR2_X1 U16221 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n12855), .ZN(
        n18342) );
  XNOR2_X1 U16222 ( .A(n12856), .B(n17909), .ZN(n12858) );
  NOR2_X1 U16223 ( .A1(n12857), .A2(n12858), .ZN(n12859) );
  INV_X1 U16224 ( .A(n12892), .ZN(n17906) );
  XNOR2_X1 U16225 ( .A(n12860), .B(n17906), .ZN(n12861) );
  XNOR2_X1 U16226 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n12861), .ZN(
        n18316) );
  OAI21_X1 U16227 ( .B1(n12862), .B2(n13029), .A(n18228), .ZN(n12863) );
  INV_X1 U16228 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18583) );
  NOR2_X1 U16229 ( .A1(n18601), .A2(n18583), .ZN(n18265) );
  NAND2_X1 U16230 ( .A1(n18265), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18562) );
  NAND2_X1 U16231 ( .A1(n18558), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18528) );
  INV_X1 U16232 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18196) );
  INV_X1 U16233 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18512) );
  NAND2_X1 U16234 ( .A1(n18601), .A2(n18583), .ZN(n18255) );
  NOR3_X1 U16235 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n18255), .ZN(n18208) );
  NAND2_X1 U16236 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18489) );
  INV_X1 U16237 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18465) );
  NAND2_X1 U16238 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18464) );
  NOR3_X1 U16239 ( .A1(n18163), .A2(n18465), .A3(n18464), .ZN(n12867) );
  NAND2_X1 U16240 ( .A1(n12867), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12973) );
  INV_X1 U16241 ( .A(n18489), .ZN(n18161) );
  NAND2_X1 U16242 ( .A1(n18161), .A2(n12867), .ZN(n18453) );
  NOR2_X1 U16243 ( .A1(n18453), .A2(n18117), .ZN(n18410) );
  NAND2_X1 U16244 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18410), .ZN(
        n18080) );
  NAND2_X1 U16245 ( .A1(n18228), .A2(n18163), .ZN(n18162) );
  NOR2_X1 U16246 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18162), .ZN(
        n12868) );
  INV_X1 U16247 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18451) );
  NAND2_X1 U16248 ( .A1(n12868), .A2(n18451), .ZN(n18122) );
  INV_X1 U16249 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18098) );
  NAND3_X1 U16250 ( .A1(n18104), .A2(n18098), .A3(n18117), .ZN(n12869) );
  INV_X1 U16251 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18433) );
  NOR2_X1 U16252 ( .A1(n18413), .A2(n18407), .ZN(n18391) );
  INV_X1 U16253 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n18047) );
  NAND2_X1 U16254 ( .A1(n13037), .A2(n18228), .ZN(n12927) );
  AOI21_X1 U16255 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n12709), .A(
        n12871), .ZN(n12882) );
  NAND3_X1 U16256 ( .A1(n12873), .A2(n12872), .A3(n12882), .ZN(n12874) );
  NOR2_X1 U16257 ( .A1(n12879), .A2(n12878), .ZN(n19371) );
  NOR2_X1 U16258 ( .A1(n18749), .A2(n18742), .ZN(n19163) );
  INV_X1 U16259 ( .A(n12881), .ZN(n12883) );
  AOI21_X1 U16260 ( .B1(n12883), .B2(n12882), .A(n12950), .ZN(n19154) );
  INV_X1 U16261 ( .A(n18732), .ZN(n12948) );
  NAND2_X1 U16262 ( .A1(n12948), .A2(n17972), .ZN(n12947) );
  INV_X1 U16263 ( .A(n12884), .ZN(n12885) );
  OAI211_X1 U16264 ( .C1(n18742), .C2(n19183), .A(n12886), .B(n12885), .ZN(
        n12887) );
  AOI211_X1 U16265 ( .C1(n13038), .C2(n12889), .A(n13026), .B(n18248), .ZN(
        n12926) );
  NOR2_X1 U16266 ( .A1(n18294), .A2(n18371), .ZN(n18142) );
  NAND2_X1 U16267 ( .A1(n18204), .A2(n18507), .ZN(n18205) );
  NAND2_X1 U16268 ( .A1(n18428), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18069) );
  INV_X1 U16269 ( .A(n18391), .ZN(n12919) );
  INV_X1 U16270 ( .A(n13029), .ZN(n17902) );
  NOR2_X1 U16271 ( .A1(n17916), .A2(n12898), .ZN(n12897) );
  NAND2_X1 U16272 ( .A1(n12897), .A2(n12891), .ZN(n12895) );
  NOR2_X1 U16273 ( .A1(n17909), .A2(n12895), .ZN(n12894) );
  NAND2_X1 U16274 ( .A1(n12894), .A2(n12892), .ZN(n12893) );
  XNOR2_X1 U16275 ( .A(n13029), .B(n12893), .ZN(n18305) );
  XNOR2_X1 U16276 ( .A(n17906), .B(n12894), .ZN(n12907) );
  XOR2_X1 U16277 ( .A(n17909), .B(n12895), .Z(n12896) );
  NAND2_X1 U16278 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12896), .ZN(
        n12906) );
  XNOR2_X1 U16279 ( .A(n18647), .B(n12896), .ZN(n18328) );
  INV_X1 U16280 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18658) );
  XNOR2_X1 U16281 ( .A(n17912), .B(n12897), .ZN(n18337) );
  XOR2_X1 U16282 ( .A(n17916), .B(n12898), .Z(n12899) );
  NAND2_X1 U16283 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12899), .ZN(
        n12904) );
  XNOR2_X1 U16284 ( .A(n12853), .B(n12899), .ZN(n18350) );
  OR2_X1 U16285 ( .A1(n18682), .A2(n12902), .ZN(n12903) );
  AOI21_X1 U16286 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17926), .A(
        n18379), .ZN(n12901) );
  INV_X1 U16287 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18687) );
  NOR2_X1 U16288 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17926), .ZN(
        n12900) );
  AOI221_X1 U16289 ( .B1(n18379), .B2(n17926), .C1(n12901), .C2(n18687), .A(
        n12900), .ZN(n18362) );
  NAND2_X1 U16290 ( .A1(n12903), .A2(n18360), .ZN(n18349) );
  NAND2_X1 U16291 ( .A1(n18350), .A2(n18349), .ZN(n18348) );
  NAND2_X1 U16292 ( .A1(n12904), .A2(n18348), .ZN(n18336) );
  NAND2_X1 U16293 ( .A1(n18337), .A2(n18336), .ZN(n12905) );
  NOR2_X1 U16294 ( .A1(n18337), .A2(n18336), .ZN(n18335) );
  NAND2_X1 U16295 ( .A1(n12907), .A2(n12908), .ZN(n12909) );
  NAND2_X1 U16296 ( .A1(n12912), .A2(n12910), .ZN(n12913) );
  NAND2_X1 U16297 ( .A1(n18305), .A2(n18304), .ZN(n12911) );
  NAND2_X1 U16298 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18285), .ZN(
        n18284) );
  NAND2_X2 U16299 ( .A1(n12913), .A2(n18284), .ZN(n18544) );
  NOR2_X2 U16300 ( .A1(n18080), .A2(n18523), .ZN(n18427) );
  NAND2_X1 U16301 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18427), .ZN(
        n18068) );
  NOR2_X2 U16302 ( .A1(n12919), .A2(n18068), .ZN(n18388) );
  OAI22_X1 U16303 ( .A1(n18389), .A2(n10295), .B1(n18388), .B2(n18385), .ZN(
        n18062) );
  NOR2_X1 U16304 ( .A1(n18047), .A2(n18062), .ZN(n12915) );
  INV_X1 U16305 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12914) );
  NOR3_X1 U16306 ( .A1(n18142), .A2(n12915), .A3(n12914), .ZN(n12924) );
  INV_X1 U16307 ( .A(n19330), .ZN(n19370) );
  NAND2_X1 U16308 ( .A1(n18707), .A2(n19335), .ZN(n17100) );
  AND2_X1 U16309 ( .A1(n18054), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12939) );
  NAND2_X1 U16310 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16805) );
  OAI21_X1 U16311 ( .B1(n12939), .B2(n16805), .A(n18381), .ZN(n12916) );
  AOI21_X1 U16312 ( .B1(n18219), .B2(n12595), .A(n12916), .ZN(n18056) );
  OAI21_X1 U16313 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18169), .A(
        n18056), .ZN(n18043) );
  INV_X1 U16314 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12917) );
  OAI21_X1 U16315 ( .B1(n17477), .B2(n18169), .A(n19061), .ZN(n18075) );
  NAND2_X1 U16316 ( .A1(n12939), .A2(n18075), .ZN(n18049) );
  AOI221_X1 U16317 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C1(n17147), .C2(n12917), .A(
        n18049), .ZN(n12918) );
  NOR2_X1 U16318 ( .A1(n18701), .A2(n19291), .ZN(n13034) );
  AOI211_X1 U16319 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n18043), .A(
        n12918), .B(n13034), .ZN(n12922) );
  NOR2_X2 U16320 ( .A1(n18283), .A2(n12968), .ZN(n18174) );
  NAND2_X1 U16321 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18408) );
  NOR2_X1 U16322 ( .A1(n12919), .A2(n18408), .ZN(n12972) );
  NAND3_X1 U16323 ( .A1(n18410), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n12972), .ZN(n12976) );
  NOR2_X1 U16324 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n12976), .ZN(
        n13036) );
  NAND2_X1 U16325 ( .A1(n18174), .A2(n13036), .ZN(n12921) );
  NAND3_X1 U16326 ( .A1(n12922), .A2(n12921), .A3(n10554), .ZN(n12923) );
  NAND2_X1 U16327 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12970) );
  INV_X1 U16328 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16889) );
  NOR2_X1 U16329 ( .A1(n12970), .A2(n16889), .ZN(n12971) );
  NAND2_X1 U16330 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n10304), .ZN(
        n12931) );
  NAND2_X1 U16331 ( .A1(n16887), .A2(n12929), .ZN(n12936) );
  INV_X1 U16332 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17000) );
  OAI21_X1 U16333 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n17000), .A(
        n12930), .ZN(n12933) );
  OAI22_X1 U16334 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n10304), .B1(
        n12931), .B2(n17000), .ZN(n12932) );
  OAI21_X1 U16335 ( .B1(n12934), .B2(n12933), .A(n12932), .ZN(n12935) );
  NAND2_X1 U16336 ( .A1(n12936), .A2(n12935), .ZN(n12986) );
  INV_X1 U16337 ( .A(n12970), .ZN(n17011) );
  NAND2_X1 U16338 ( .A1(n18389), .A2(n17011), .ZN(n13028) );
  INV_X1 U16339 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19319) );
  NAND3_X1 U16340 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n19319), .ZN(n12966) );
  NAND2_X1 U16341 ( .A1(n18389), .A2(n12971), .ZN(n16820) );
  OAI21_X1 U16342 ( .B1(n17000), .B2(n16820), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12937) );
  OAI21_X1 U16343 ( .B1(n13028), .B2(n12966), .A(n12937), .ZN(n12964) );
  NAND2_X1 U16344 ( .A1(n17011), .A2(n18388), .ZN(n16818) );
  NAND2_X1 U16345 ( .A1(n12971), .A2(n18388), .ZN(n16821) );
  OAI21_X1 U16346 ( .B1(n17000), .B2(n16821), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12938) );
  OAI21_X1 U16347 ( .B1(n12966), .B2(n16818), .A(n12938), .ZN(n12965) );
  AOI22_X1 U16348 ( .A1(n18294), .A2(n12964), .B1(n18371), .B2(n12965), .ZN(
        n12945) );
  NOR2_X1 U16349 ( .A1(n19297), .A2(n18701), .ZN(n12980) );
  NAND3_X1 U16350 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(n12939), .ZN(n13281) );
  NOR2_X1 U16351 ( .A1(n17121), .A2(n13281), .ZN(n12940) );
  NAND2_X1 U16352 ( .A1(n12940), .A2(n18075), .ZN(n17006) );
  XOR2_X1 U16353 ( .A(n12605), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n12942) );
  NOR2_X1 U16354 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18169), .ZN(
        n13279) );
  INV_X1 U16355 ( .A(n12592), .ZN(n12941) );
  OR2_X1 U16356 ( .A1(n19061), .A2(n12940), .ZN(n13282) );
  OAI211_X1 U16357 ( .C1(n12941), .C2(n18380), .A(n18381), .B(n13282), .ZN(
        n13283) );
  NOR2_X1 U16358 ( .A1(n13279), .A2(n13283), .ZN(n17004) );
  OAI22_X1 U16359 ( .A1(n17006), .A2(n12942), .B1(n17004), .B2(n12605), .ZN(
        n12943) );
  AOI211_X1 U16360 ( .C1(n18140), .C2(n10321), .A(n12980), .B(n12943), .ZN(
        n12944) );
  OAI21_X1 U16361 ( .B1(n12986), .B2(n18248), .A(n12946), .ZN(P3_U2799) );
  OAI21_X1 U16362 ( .B1(n12948), .B2(n17972), .A(n12947), .ZN(n12949) );
  OAI21_X1 U16363 ( .B1(n19228), .B2(n12949), .A(n19361), .ZN(n17102) );
  NOR3_X1 U16364 ( .A1(n12951), .A2(n12950), .A3(n17102), .ZN(n12958) );
  INV_X1 U16365 ( .A(n12952), .ZN(n12955) );
  OAI21_X1 U16366 ( .B1(n12955), .B2(n12954), .A(n12953), .ZN(n12957) );
  NAND2_X1 U16367 ( .A1(n12957), .A2(n12956), .ZN(n14233) );
  AOI211_X1 U16368 ( .C1(n12959), .C2(n19154), .A(n12958), .B(n14233), .ZN(
        n12962) );
  OAI21_X1 U16369 ( .B1(n12960), .B2(n14224), .A(n9744), .ZN(n12961) );
  NOR2_X1 U16370 ( .A1(n17902), .A2(n19155), .ZN(n18403) );
  NOR2_X1 U16371 ( .A1(n13029), .A2(n18693), .ZN(n18617) );
  AOI22_X1 U16372 ( .A1(n18698), .A2(n12965), .B1(n18617), .B2(n12964), .ZN(
        n12984) );
  INV_X1 U16373 ( .A(n12966), .ZN(n12982) );
  NOR3_X1 U16374 ( .A1(n18658), .A2(n12853), .A3(n18647), .ZN(n18607) );
  INV_X1 U16375 ( .A(n18607), .ZN(n18622) );
  NAND2_X1 U16376 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18609) );
  OR2_X1 U16377 ( .A1(n18622), .A2(n18609), .ZN(n12967) );
  OR2_X1 U16378 ( .A1(n18613), .A2(n12967), .ZN(n18515) );
  AOI21_X1 U16379 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18603) );
  OR2_X1 U16380 ( .A1(n18515), .A2(n18603), .ZN(n18548) );
  NOR2_X1 U16381 ( .A1(n12968), .A2(n18548), .ZN(n12974) );
  NOR3_X1 U16382 ( .A1(n18682), .A2(n19320), .A3(n12967), .ZN(n18594) );
  NAND2_X1 U16383 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18594), .ZN(
        n18546) );
  NOR2_X1 U16384 ( .A1(n12968), .A2(n18546), .ZN(n18487) );
  OAI21_X1 U16385 ( .B1(n19169), .B2(n18687), .A(n19184), .ZN(n18671) );
  AOI22_X1 U16386 ( .A1(n10298), .A2(n12974), .B1(n18487), .B2(n18671), .ZN(
        n13033) );
  NAND2_X1 U16387 ( .A1(n18410), .A2(n12972), .ZN(n12969) );
  NOR4_X1 U16388 ( .A1(n13033), .A2(n18702), .A3(n12970), .A4(n12969), .ZN(
        n16815) );
  NOR2_X1 U16389 ( .A1(n18608), .A2(n18702), .ZN(n18651) );
  INV_X1 U16390 ( .A(n12971), .ZN(n12979) );
  INV_X1 U16391 ( .A(n12972), .ZN(n18387) );
  INV_X1 U16392 ( .A(n12973), .ZN(n12975) );
  INV_X1 U16393 ( .A(n12974), .ZN(n18449) );
  OAI21_X1 U16394 ( .B1(n18489), .B2(n18449), .A(n10298), .ZN(n18490) );
  OAI21_X1 U16395 ( .B1(n12975), .B2(n19177), .A(n18490), .ZN(n18432) );
  AOI21_X1 U16396 ( .B1(n10298), .B2(n18387), .A(n18432), .ZN(n18390) );
  NOR2_X1 U16397 ( .A1(n18687), .A2(n18546), .ZN(n18593) );
  NAND2_X1 U16398 ( .A1(n10179), .A2(n18593), .ZN(n18505) );
  OAI21_X1 U16399 ( .B1(n18505), .B2(n12976), .A(n19182), .ZN(n12978) );
  NAND2_X1 U16400 ( .A1(n18410), .A2(n18487), .ZN(n18424) );
  OAI21_X1 U16401 ( .B1(n18387), .B2(n18424), .A(n18703), .ZN(n12977) );
  NAND4_X1 U16402 ( .A1(n18390), .A2(n18685), .A3(n12978), .A4(n12977), .ZN(
        n13030) );
  AOI22_X1 U16403 ( .A1(n18651), .A2(n12979), .B1(n18701), .B2(n13030), .ZN(
        n16891) );
  INV_X1 U16404 ( .A(n18651), .ZN(n18686) );
  AOI221_X1 U16405 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16891), 
        .C1(n18686), .C2(n16891), .A(n19319), .ZN(n12981) );
  AOI211_X1 U16406 ( .C1(n12982), .C2(n16815), .A(n12981), .B(n12980), .ZN(
        n12983) );
  AND2_X1 U16407 ( .A1(n12984), .A2(n12983), .ZN(n12985) );
  OAI21_X1 U16408 ( .B1(n12986), .B2(n18567), .A(n12985), .ZN(P3_U2831) );
  AOI21_X1 U16409 ( .B1(n12987), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12989) );
  NOR2_X1 U16410 ( .A1(n12992), .A2(n12991), .ZN(n12993) );
  XNOR2_X1 U16411 ( .A(n12990), .B(n12993), .ZN(n16188) );
  NOR2_X1 U16412 ( .A1(n12994), .A2(n12995), .ZN(n12996) );
  INV_X1 U16413 ( .A(n16185), .ZN(n15586) );
  NAND2_X1 U16414 ( .A1(n12998), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12999) );
  NOR2_X1 U16415 ( .A1(n13000), .A2(n12999), .ZN(n16446) );
  OAI21_X1 U16416 ( .B1(n16448), .B2(n16446), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13005) );
  NAND2_X1 U16417 ( .A1(n16434), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n16183) );
  NAND3_X1 U16418 ( .A1(n13003), .A2(n13002), .A3(n13001), .ZN(n13004) );
  NAND3_X1 U16419 ( .A1(n13005), .A2(n16183), .A3(n13004), .ZN(n13006) );
  AOI21_X1 U16420 ( .B1(n15586), .B2(n16727), .A(n13006), .ZN(n13011) );
  NAND2_X1 U16421 ( .A1(n15595), .A2(n13007), .ZN(n13008) );
  NAND2_X1 U16422 ( .A1(n15580), .A2(n16724), .ZN(n13010) );
  OAI21_X1 U16423 ( .B1(n16190), .B2(n16706), .A(n13013), .ZN(P2_U3017) );
  INV_X1 U16424 ( .A(n19381), .ZN(n13532) );
  AND2_X1 U16425 ( .A1(n16778), .A2(n13532), .ZN(n13045) );
  OR2_X1 U16426 ( .A1(n20258), .A2(n16754), .ZN(n20255) );
  NAND2_X1 U16427 ( .A1(n20255), .A2(n14059), .ZN(n13016) );
  AND2_X1 U16428 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n16733) );
  INV_X1 U16429 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13022) );
  NAND2_X1 U16430 ( .A1(n13086), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13089) );
  NAND2_X1 U16431 ( .A1(n13102), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13105) );
  INV_X1 U16432 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13108) );
  INV_X1 U16433 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13112) );
  INV_X1 U16434 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15626) );
  OR2_X2 U16435 ( .A1(n13118), .A2(n15626), .ZN(n13120) );
  AND2_X1 U16436 ( .A1(n13120), .A2(n13022), .ZN(n13018) );
  NOR2_X1 U16437 ( .A1(n13122), .A2(n13018), .ZN(n15611) );
  NAND2_X1 U16438 ( .A1(n20036), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13049) );
  NAND2_X1 U16439 ( .A1(n13630), .A2(n13049), .ZN(n13019) );
  NAND2_X1 U16440 ( .A1(n15611), .A2(n16433), .ZN(n13021) );
  OAI211_X1 U16441 ( .C1(n13022), .C2(n16436), .A(n13021), .B(n13020), .ZN(
        n13023) );
  INV_X1 U16442 ( .A(n18450), .ZN(n19150) );
  INV_X1 U16443 ( .A(n13028), .ZN(n16816) );
  NOR2_X1 U16444 ( .A1(n13029), .A2(n19155), .ZN(n18571) );
  OR2_X1 U16445 ( .A1(n16816), .A2(n18549), .ZN(n13031) );
  NAND2_X1 U16446 ( .A1(n19184), .A2(n19177), .ZN(n18547) );
  AOI21_X1 U16447 ( .B1(n18047), .B2(n18547), .A(n13030), .ZN(n16819) );
  AND2_X1 U16448 ( .A1(n13031), .A2(n16819), .ZN(n13032) );
  NAND2_X1 U16449 ( .A1(n18701), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13043) );
  INV_X1 U16450 ( .A(n13033), .ZN(n18409) );
  OAI22_X1 U16451 ( .A1(n18450), .A2(n18523), .B1(n18514), .B2(n18549), .ZN(
        n18486) );
  NOR2_X1 U16452 ( .A1(n18409), .A2(n18486), .ZN(n18386) );
  NOR2_X1 U16453 ( .A1(n18386), .A2(n18702), .ZN(n18479) );
  NOR4_X1 U16454 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18228), .A3(
        n18045), .A4(n18693), .ZN(n13035) );
  AOI211_X1 U16455 ( .C1(n18479), .C2(n13036), .A(n13035), .B(n13034), .ZN(
        n13041) );
  INV_X1 U16456 ( .A(n13037), .ZN(n13039) );
  NAND2_X1 U16457 ( .A1(n13039), .A2(n10575), .ZN(n13040) );
  OAI21_X1 U16458 ( .B1(n13044), .B2(n13043), .A(n13042), .ZN(P3_U2834) );
  NAND2_X1 U16459 ( .A1(n15574), .A2(n20036), .ZN(n13046) );
  NAND2_X1 U16460 ( .A1(n13348), .A2(n13046), .ZN(n13054) );
  INV_X1 U16461 ( .A(n13054), .ZN(n13048) );
  NAND2_X1 U16462 ( .A1(n13903), .A2(n13910), .ZN(n13917) );
  INV_X1 U16463 ( .A(n13049), .ZN(n13050) );
  NAND2_X1 U16464 ( .A1(n13050), .A2(n13340), .ZN(n16789) );
  NAND2_X1 U16465 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20044), .ZN(n19785) );
  INV_X1 U16466 ( .A(n19785), .ZN(n13051) );
  NAND2_X1 U16467 ( .A1(n13352), .A2(n13051), .ZN(n14061) );
  NAND2_X1 U16468 ( .A1(n16789), .A2(n14061), .ZN(n13052) );
  NOR2_X1 U16469 ( .A1(n13052), .A2(n16434), .ZN(n13053) );
  AND2_X2 U16470 ( .A1(n15576), .A2(n13053), .ZN(n19402) );
  INV_X1 U16471 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16173) );
  AND2_X1 U16472 ( .A1(n13916), .A2(n20036), .ZN(n13927) );
  OR2_X1 U16473 ( .A1(n13392), .A2(n13927), .ZN(n14358) );
  OR2_X1 U16474 ( .A1(n13054), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n13055) );
  AOI22_X1 U16475 ( .A1(n19402), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n16835), 
        .B2(P2_EBX_REG_30__SCAN_IN), .ZN(n13056) );
  OAI21_X1 U16476 ( .B1(n19424), .B2(n16173), .A(n13056), .ZN(n13059) );
  INV_X1 U16477 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13061) );
  XNOR2_X1 U16478 ( .A(n13062), .B(n13061), .ZN(n14342) );
  MUX2_X2 U16479 ( .A(n14342), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n19409) );
  MUX2_X1 U16480 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n16740) );
  INV_X1 U16481 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15960) );
  MUX2_X1 U16482 ( .A(n15960), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n15951) );
  INV_X1 U16483 ( .A(n13063), .ZN(n13065) );
  INV_X1 U16484 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14636) );
  NAND2_X1 U16485 ( .A1(n15960), .A2(n14636), .ZN(n13064) );
  NAND2_X1 U16486 ( .A1(n13065), .A2(n13064), .ZN(n15941) );
  NAND2_X1 U16487 ( .A1(n15940), .A2(n15941), .ZN(n15922) );
  OAI21_X1 U16488 ( .B1(n13063), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13066), .ZN(n15924) );
  INV_X1 U16489 ( .A(n15924), .ZN(n13067) );
  OR2_X1 U16490 ( .A1(n15922), .A2(n13067), .ZN(n15906) );
  AND2_X1 U16491 ( .A1(n13066), .A2(n13069), .ZN(n13070) );
  NOR2_X1 U16492 ( .A1(n13068), .A2(n13070), .ZN(n15908) );
  OR2_X1 U16493 ( .A1(n13068), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13072) );
  NAND2_X1 U16494 ( .A1(n13071), .A2(n13072), .ZN(n15893) );
  NAND2_X1 U16495 ( .A1(n15891), .A2(n15893), .ZN(n19408) );
  NAND2_X1 U16496 ( .A1(n13071), .A2(n16437), .ZN(n13073) );
  AND2_X1 U16497 ( .A1(n13075), .A2(n13073), .ZN(n19411) );
  AND2_X1 U16498 ( .A1(n13075), .A2(n21303), .ZN(n13076) );
  NOR2_X1 U16499 ( .A1(n13074), .A2(n13076), .ZN(n16419) );
  NOR2_X1 U16500 ( .A1(n13074), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13078) );
  OR2_X1 U16501 ( .A1(n13077), .A2(n13078), .ZN(n16412) );
  NAND2_X1 U16502 ( .A1(n15874), .A2(n16412), .ZN(n15856) );
  OR2_X1 U16503 ( .A1(n13077), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13080) );
  AND2_X1 U16504 ( .A1(n13079), .A2(n13080), .ZN(n16395) );
  OR2_X1 U16505 ( .A1(n15856), .A2(n16395), .ZN(n15849) );
  NAND2_X1 U16506 ( .A1(n13079), .A2(n10379), .ZN(n13082) );
  AND2_X1 U16507 ( .A1(n13081), .A2(n13082), .ZN(n16386) );
  NAND2_X1 U16508 ( .A1(n13081), .A2(n15829), .ZN(n13083) );
  NAND2_X1 U16509 ( .A1(n13084), .A2(n13083), .ZN(n16366) );
  AND2_X1 U16510 ( .A1(n15835), .A2(n16366), .ZN(n15820) );
  AND2_X1 U16511 ( .A1(n13084), .A2(n15815), .ZN(n13085) );
  OR2_X1 U16512 ( .A1(n13085), .A2(n13086), .ZN(n16356) );
  NAND2_X1 U16513 ( .A1(n15820), .A2(n16356), .ZN(n15802) );
  OR2_X1 U16514 ( .A1(n13086), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13087) );
  AND2_X1 U16515 ( .A1(n13087), .A2(n13089), .ZN(n16345) );
  OR2_X1 U16516 ( .A1(n15802), .A2(n16345), .ZN(n15796) );
  INV_X1 U16517 ( .A(n13088), .ZN(n13091) );
  NAND2_X1 U16518 ( .A1(n13089), .A2(n16332), .ZN(n13090) );
  AND2_X1 U16519 ( .A1(n13091), .A2(n13090), .ZN(n16334) );
  AND2_X1 U16520 ( .A1(n13091), .A2(n15778), .ZN(n13093) );
  OR2_X1 U16521 ( .A1(n13093), .A2(n13092), .ZN(n16320) );
  NAND2_X1 U16522 ( .A1(n15783), .A2(n16320), .ZN(n15763) );
  NOR2_X1 U16523 ( .A1(n13092), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13095) );
  OR2_X1 U16524 ( .A1(n13094), .A2(n13095), .ZN(n16312) );
  INV_X1 U16525 ( .A(n16312), .ZN(n15765) );
  OR2_X1 U16526 ( .A1(n13094), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13097) );
  AND2_X1 U16527 ( .A1(n13096), .A2(n13097), .ZN(n16297) );
  NAND2_X1 U16528 ( .A1(n13096), .A2(n15736), .ZN(n13099) );
  NAND2_X1 U16529 ( .A1(n13098), .A2(n13099), .ZN(n16287) );
  AND2_X1 U16530 ( .A1(n13098), .A2(n15725), .ZN(n13101) );
  OR2_X1 U16531 ( .A1(n13101), .A2(n13100), .ZN(n16279) );
  NAND2_X1 U16532 ( .A1(n15719), .A2(n16279), .ZN(n15707) );
  NOR2_X1 U16533 ( .A1(n13100), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13103) );
  OR2_X1 U16534 ( .A1(n13102), .A2(n13103), .ZN(n16270) );
  INV_X1 U16535 ( .A(n16270), .ZN(n15710) );
  OR2_X1 U16536 ( .A1(n13102), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13106) );
  NAND2_X1 U16537 ( .A1(n13105), .A2(n13106), .ZN(n16257) );
  NAND2_X1 U16538 ( .A1(n13105), .A2(n16837), .ZN(n13107) );
  NAND2_X1 U16539 ( .A1(n13109), .A2(n13107), .ZN(n16830) );
  NAND2_X1 U16540 ( .A1(n16842), .A2(n19409), .ZN(n13111) );
  NAND2_X1 U16541 ( .A1(n13109), .A2(n13108), .ZN(n13110) );
  NAND2_X1 U16542 ( .A1(n13113), .A2(n13110), .ZN(n16233) );
  NAND2_X1 U16543 ( .A1(n13111), .A2(n16233), .ZN(n15660) );
  NAND2_X1 U16544 ( .A1(n15660), .A2(n19409), .ZN(n13115) );
  AND2_X1 U16545 ( .A1(n13113), .A2(n13112), .ZN(n13114) );
  OR2_X1 U16546 ( .A1(n13114), .A2(n13116), .ZN(n16224) );
  OR2_X1 U16547 ( .A1(n13116), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13117) );
  AND2_X1 U16548 ( .A1(n13117), .A2(n13118), .ZN(n16216) );
  NAND2_X1 U16549 ( .A1(n13118), .A2(n15626), .ZN(n13119) );
  NAND2_X1 U16550 ( .A1(n13120), .A2(n13119), .ZN(n16207) );
  NOR2_X1 U16551 ( .A1(n13122), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13123) );
  OR2_X1 U16552 ( .A1(n13121), .A2(n13123), .ZN(n16199) );
  OAI21_X2 U16553 ( .B1(n15602), .B2(n16750), .A(n16199), .ZN(n15587) );
  OR2_X1 U16554 ( .A1(n13121), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13124) );
  NAND2_X1 U16555 ( .A1(n9736), .A2(n13124), .ZN(n16184) );
  INV_X1 U16556 ( .A(n16184), .ZN(n15588) );
  INV_X1 U16557 ( .A(n13126), .ZN(n15589) );
  XNOR2_X1 U16558 ( .A(n9736), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16175) );
  AOI21_X1 U16559 ( .B1(n15589), .B2(n16175), .A(n16789), .ZN(n13127) );
  INV_X1 U16560 ( .A(n16175), .ZN(n13125) );
  OAI21_X1 U16561 ( .B1(n15964), .B2(n13127), .A(n14364), .ZN(n13132) );
  INV_X1 U16562 ( .A(n15576), .ZN(n13354) );
  INV_X1 U16563 ( .A(n13927), .ZN(n13128) );
  INV_X1 U16564 ( .A(n13928), .ZN(n15567) );
  NOR2_X1 U16565 ( .A1(n13128), .A2(n15567), .ZN(n13129) );
  NAND3_X1 U16566 ( .A1(n13133), .A2(n13132), .A3(n13131), .ZN(P2_U2825) );
  INV_X1 U16567 ( .A(n14003), .ZN(n13134) );
  XOR2_X1 U16568 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n13134), .Z(
        n14677) );
  INV_X1 U16569 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14002) );
  AOI21_X1 U16570 ( .B1(n14002), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13135) );
  AOI21_X1 U16571 ( .B1(n11374), .B2(P1_EAX_REG_30__SCAN_IN), .A(n13135), .ZN(
        n13161) );
  NOR2_X1 U16572 ( .A1(n13137), .A2(n13136), .ZN(n13157) );
  AOI22_X1 U16573 ( .A1(n13139), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13138), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13145) );
  AOI22_X1 U16574 ( .A1(n11281), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10700), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13144) );
  AOI22_X1 U16575 ( .A1(n10667), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10646), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13143) );
  AOI22_X1 U16576 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n13141), .B1(
        n13140), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13142) );
  NAND4_X1 U16577 ( .A1(n13145), .A2(n13144), .A3(n13143), .A4(n13142), .ZN(
        n13155) );
  AOI22_X1 U16578 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n13146), .B1(
        n10732), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13153) );
  AOI22_X1 U16579 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n15522), .B1(
        n13147), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13152) );
  AOI22_X1 U16580 ( .A1(n10791), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9608), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13151) );
  AOI22_X1 U16581 ( .A1(n13149), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13148), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13150) );
  NAND4_X1 U16582 ( .A1(n13153), .A2(n13152), .A3(n13151), .A4(n13150), .ZN(
        n13154) );
  NOR2_X1 U16583 ( .A1(n13155), .A2(n13154), .ZN(n13156) );
  XNOR2_X1 U16584 ( .A(n13157), .B(n13156), .ZN(n13159) );
  NAND2_X1 U16585 ( .A1(n13159), .A2(n13158), .ZN(n13160) );
  AOI22_X1 U16586 ( .A1(n14677), .A2(n13162), .B1(n13161), .B2(n13160), .ZN(
        n13292) );
  NAND3_X1 U16587 ( .A1(n10144), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16990) );
  INV_X1 U16588 ( .A(n16990), .ZN(n13163) );
  AND2_X1 U16589 ( .A1(n13164), .A2(n13222), .ZN(n13165) );
  INV_X1 U16590 ( .A(n13222), .ZN(n13645) );
  AND2_X1 U16591 ( .A1(n13167), .A2(n13222), .ZN(n13168) );
  NAND2_X1 U16592 ( .A1(n13183), .A2(n13182), .ZN(n13175) );
  NAND2_X1 U16593 ( .A1(n13175), .A2(n13176), .ZN(n13203) );
  NAND2_X1 U16594 ( .A1(n13203), .A2(n13201), .ZN(n13171) );
  INV_X1 U16595 ( .A(n13171), .ZN(n13173) );
  INV_X1 U16596 ( .A(n13172), .ZN(n13170) );
  OR2_X1 U16597 ( .A1(n13171), .A2(n13170), .ZN(n13214) );
  OAI211_X1 U16598 ( .C1(n13173), .C2(n13172), .A(n10847), .B(n13214), .ZN(
        n13174) );
  OAI21_X1 U16599 ( .B1(n13176), .B2(n13175), .A(n13203), .ZN(n13178) );
  NAND2_X1 U16600 ( .A1(n14010), .A2(n20516), .ZN(n13647) );
  INV_X1 U16601 ( .A(n13647), .ZN(n13177) );
  AOI21_X1 U16602 ( .B1(n13178), .B2(n10847), .A(n13177), .ZN(n13179) );
  NAND2_X1 U16603 ( .A1(n13180), .A2(n13179), .ZN(n13748) );
  INV_X1 U16604 ( .A(n13182), .ZN(n13188) );
  XNOR2_X1 U16605 ( .A(n13188), .B(n13183), .ZN(n13185) );
  NAND2_X1 U16606 ( .A1(n13712), .A2(n20524), .ZN(n13184) );
  AOI21_X1 U16607 ( .B1(n13185), .B2(n10847), .A(n13184), .ZN(n13186) );
  NAND2_X1 U16608 ( .A1(n13187), .A2(n13186), .ZN(n13195) );
  NAND2_X1 U16609 ( .A1(n10847), .A2(n13188), .ZN(n13646) );
  NAND2_X1 U16610 ( .A1(n13646), .A2(n13647), .ZN(n13190) );
  OR2_X1 U16611 ( .A1(n13190), .A2(n13189), .ZN(n13192) );
  INV_X1 U16612 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13732) );
  AOI21_X1 U16613 ( .B1(n9939), .B2(n13645), .A(n13732), .ZN(n13191) );
  NAND2_X1 U16614 ( .A1(n13726), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13197) );
  INV_X1 U16615 ( .A(n13649), .ZN(n13194) );
  NAND2_X1 U16616 ( .A1(n13195), .A2(n13194), .ZN(n13196) );
  NAND2_X1 U16617 ( .A1(n13199), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13200) );
  INV_X1 U16618 ( .A(n13201), .ZN(n13202) );
  XNOR2_X1 U16619 ( .A(n13203), .B(n13202), .ZN(n13204) );
  NAND2_X1 U16620 ( .A1(n13204), .A2(n10847), .ZN(n13205) );
  INV_X1 U16621 ( .A(n13987), .ZN(n13207) );
  INV_X1 U16622 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13206) );
  NAND2_X1 U16623 ( .A1(n13207), .A2(n13206), .ZN(n13208) );
  XNOR2_X1 U16624 ( .A(n13214), .B(n13215), .ZN(n13209) );
  NAND2_X1 U16625 ( .A1(n13209), .A2(n10847), .ZN(n13210) );
  INV_X1 U16626 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16979) );
  NAND2_X1 U16627 ( .A1(n13211), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13212) );
  OR2_X1 U16628 ( .A1(n13213), .A2(n13645), .ZN(n13219) );
  INV_X1 U16629 ( .A(n13214), .ZN(n13216) );
  NAND2_X1 U16630 ( .A1(n13216), .A2(n13215), .ZN(n13223) );
  XNOR2_X1 U16631 ( .A(n13223), .B(n13224), .ZN(n13217) );
  NAND2_X1 U16632 ( .A1(n13217), .A2(n10847), .ZN(n13218) );
  NAND2_X1 U16633 ( .A1(n13219), .A2(n13218), .ZN(n13221) );
  INV_X1 U16634 ( .A(n13221), .ZN(n13220) );
  NAND2_X1 U16635 ( .A1(n13220), .A2(n16945), .ZN(n16923) );
  NAND2_X1 U16636 ( .A1(n13221), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16922) );
  NAND2_X1 U16637 ( .A1(n14126), .A2(n13222), .ZN(n13228) );
  INV_X1 U16638 ( .A(n13223), .ZN(n13225) );
  NAND2_X1 U16639 ( .A1(n13225), .A2(n13224), .ZN(n13231) );
  XNOR2_X1 U16640 ( .A(n13231), .B(n13229), .ZN(n13226) );
  NAND2_X1 U16641 ( .A1(n13226), .A2(n10847), .ZN(n13227) );
  NAND2_X1 U16642 ( .A1(n13228), .A2(n13227), .ZN(n16916) );
  NAND2_X1 U16643 ( .A1(n10847), .A2(n13229), .ZN(n13230) );
  OR2_X1 U16644 ( .A1(n13231), .A2(n13230), .ZN(n13232) );
  OAI21_X1 U16645 ( .B1(n16916), .B2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13235) );
  INV_X1 U16646 ( .A(n15247), .ZN(n13234) );
  INV_X1 U16647 ( .A(n16916), .ZN(n15244) );
  NOR2_X1 U16648 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13233) );
  AOI22_X1 U16649 ( .A1(n13235), .A2(n13234), .B1(n15244), .B2(n13233), .ZN(
        n13236) );
  INV_X1 U16650 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15512) );
  NAND2_X1 U16651 ( .A1(n15236), .A2(n15512), .ZN(n13238) );
  INV_X1 U16652 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15457) );
  NAND2_X1 U16653 ( .A1(n15236), .A2(n15457), .ZN(n13239) );
  NAND2_X1 U16654 ( .A1(n15185), .A2(n13239), .ZN(n15200) );
  NAND2_X1 U16655 ( .A1(n15216), .A2(n15471), .ZN(n15199) );
  NAND2_X1 U16656 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13240) );
  NOR2_X1 U16657 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13241) );
  OR2_X1 U16658 ( .A1(n15236), .A2(n13241), .ZN(n13242) );
  AND2_X1 U16659 ( .A1(n15179), .A2(n13242), .ZN(n15154) );
  NAND2_X1 U16660 ( .A1(n15236), .A2(n15429), .ZN(n15178) );
  NAND2_X1 U16661 ( .A1(n15166), .A2(n15178), .ZN(n13243) );
  OAI21_X1 U16662 ( .B1(n10583), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15153), .ZN(n13247) );
  NOR2_X1 U16663 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15152) );
  AND4_X1 U16664 ( .A1(n15152), .A2(n15444), .A3(n15457), .A4(n15471), .ZN(
        n13244) );
  NOR2_X1 U16665 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13245) );
  XNOR2_X1 U16666 ( .A(n15236), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15146) );
  AND2_X1 U16667 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15262) );
  NAND2_X1 U16668 ( .A1(n15262), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15362) );
  INV_X1 U16669 ( .A(n15362), .ZN(n13248) );
  INV_X1 U16670 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15371) );
  INV_X1 U16671 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15327) );
  INV_X1 U16672 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15337) );
  NOR2_X1 U16673 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15303) );
  AND2_X1 U16674 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15277) );
  NAND2_X1 U16675 ( .A1(n15277), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15265) );
  AND2_X1 U16676 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15304) );
  NAND2_X1 U16677 ( .A1(n15236), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15047) );
  NAND2_X1 U16678 ( .A1(n13254), .A2(n14010), .ZN(n13255) );
  NAND2_X1 U16679 ( .A1(n21010), .A2(n13259), .ZN(n21174) );
  NAND2_X1 U16680 ( .A1(n21174), .A2(n10144), .ZN(n13256) );
  NAND2_X1 U16681 ( .A1(n10144), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13258) );
  NAND2_X1 U16682 ( .A1(n20979), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13257) );
  NAND2_X1 U16683 ( .A1(n13258), .A2(n13257), .ZN(n13652) );
  NAND2_X1 U16684 ( .A1(n14677), .A2(n15241), .ZN(n13262) );
  NAND2_X1 U16685 ( .A1(n16962), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15289) );
  OAI21_X1 U16686 ( .B1(n16937), .B2(n14002), .A(n15289), .ZN(n13260) );
  INV_X1 U16687 ( .A(n13260), .ZN(n13261) );
  NAND2_X1 U16688 ( .A1(n13262), .A2(n13261), .ZN(n13263) );
  INV_X1 U16689 ( .A(n17009), .ZN(n13264) );
  XNOR2_X1 U16690 ( .A(n13265), .B(n13264), .ZN(n13273) );
  OAI21_X1 U16691 ( .B1(n17408), .B2(n13266), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n13271) );
  INV_X1 U16692 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17005) );
  OAI22_X1 U16693 ( .A1(n17005), .A2(n17471), .B1(n19299), .B2(n17132), .ZN(
        n13268) );
  NAND2_X1 U16694 ( .A1(n17470), .A2(n13269), .ZN(n17128) );
  NAND3_X1 U16695 ( .A1(n13271), .A2(n10576), .A3(n13270), .ZN(n13272) );
  AOI21_X1 U16696 ( .B1(n13273), .B2(n19216), .A(n13272), .ZN(n13274) );
  INV_X1 U16697 ( .A(n13274), .ZN(P3_U2641) );
  NOR2_X1 U16698 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16816), .ZN(
        n13277) );
  NAND2_X1 U16699 ( .A1(n18294), .A2(n16820), .ZN(n17001) );
  OAI22_X1 U16700 ( .A1(n16826), .A2(n18248), .B1(n13277), .B2(n17001), .ZN(
        n13278) );
  INV_X1 U16701 ( .A(n13278), .ZN(n13291) );
  NAND2_X1 U16702 ( .A1(n18371), .A2(n16821), .ZN(n17002) );
  INV_X1 U16703 ( .A(n17002), .ZN(n13289) );
  NAND2_X1 U16704 ( .A1(n16818), .A2(n16889), .ZN(n13288) );
  INV_X2 U16705 ( .A(n18701), .ZN(n18695) );
  NAND2_X1 U16706 ( .A1(n18695), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16824) );
  OAI21_X1 U16707 ( .B1(n18140), .B2(n13279), .A(n17118), .ZN(n13280) );
  OAI211_X1 U16708 ( .C1(n13282), .C2(n13281), .A(n16824), .B(n13280), .ZN(
        n13286) );
  INV_X1 U16709 ( .A(n13283), .ZN(n13284) );
  NAND2_X1 U16710 ( .A1(n13293), .A2(n13292), .ZN(n13296) );
  AOI22_X1 U16711 ( .A1(n11374), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n13810), .ZN(n13294) );
  INV_X1 U16712 ( .A(n13294), .ZN(n13295) );
  OR2_X1 U16713 ( .A1(n16883), .A2(n13721), .ZN(n13303) );
  INV_X1 U16714 ( .A(n13454), .ZN(n15544) );
  NOR3_X1 U16715 ( .A1(n13299), .A2(n13298), .A3(n13297), .ZN(n13300) );
  OR2_X1 U16716 ( .A1(n13301), .A2(n13300), .ZN(n13386) );
  NOR2_X1 U16717 ( .A1(n13386), .A2(n21075), .ZN(n13706) );
  NAND2_X1 U16718 ( .A1(n15544), .A2(n13706), .ZN(n13302) );
  NAND2_X1 U16719 ( .A1(n13303), .A2(n13302), .ZN(n13478) );
  NAND2_X1 U16720 ( .A1(n13478), .A2(n13718), .ZN(n13305) );
  AND2_X1 U16721 ( .A1(n15031), .A2(n14974), .ZN(n13307) );
  NAND2_X1 U16722 ( .A1(n14650), .A2(n13307), .ZN(n13324) );
  NOR4_X1 U16723 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_15__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_13__SCAN_IN), .ZN(n13311) );
  NOR4_X1 U16724 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_19__SCAN_IN), .A3(P1_ADDRESS_REG_18__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n13310) );
  NOR4_X1 U16725 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13309) );
  NOR4_X1 U16726 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(
        P1_ADDRESS_REG_11__SCAN_IN), .A3(P1_ADDRESS_REG_10__SCAN_IN), .A4(
        P1_ADDRESS_REG_9__SCAN_IN), .ZN(n13308) );
  AND4_X1 U16727 ( .A1(n13311), .A2(n13310), .A3(n13309), .A4(n13308), .ZN(
        n13316) );
  NOR4_X1 U16728 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_6__SCAN_IN), .ZN(n13314) );
  NOR4_X1 U16729 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(
        P1_ADDRESS_REG_23__SCAN_IN), .A3(P1_ADDRESS_REG_22__SCAN_IN), .A4(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n13313) );
  NOR4_X1 U16730 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_25__SCAN_IN), .ZN(n13312) );
  AND4_X1 U16731 ( .A1(n13314), .A2(n13313), .A3(n13312), .A4(n21095), .ZN(
        n13315) );
  NAND2_X1 U16732 ( .A1(n13316), .A2(n13315), .ZN(n13317) );
  NAND3_X1 U16733 ( .A1(n15031), .A2(n13708), .A3(n20492), .ZN(n14973) );
  INV_X1 U16734 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n17018) );
  NOR2_X1 U16735 ( .A1(n14973), .A2(n17018), .ZN(n13322) );
  NOR3_X1 U16736 ( .A1(n15041), .A2(n20492), .A3(n13318), .ZN(n13319) );
  AOI22_X1 U16737 ( .A1(n15018), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15041), .ZN(n13320) );
  INV_X1 U16738 ( .A(n13320), .ZN(n13321) );
  NOR2_X1 U16739 ( .A1(n13322), .A2(n13321), .ZN(n13323) );
  NAND2_X1 U16740 ( .A1(n13324), .A2(n13323), .ZN(P1_U2873) );
  NOR2_X1 U16741 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13326) );
  NOR4_X1 U16742 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13325) );
  NAND4_X1 U16743 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13326), .A4(n13325), .ZN(n13339) );
  INV_X1 U16744 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21171) );
  NOR3_X1 U16745 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n21171), .ZN(n13328) );
  NOR4_X1 U16746 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_2__SCAN_IN), 
        .A3(P1_BE_N_REG_3__SCAN_IN), .A4(P1_D_C_N_REG_SCAN_IN), .ZN(n13327) );
  NAND4_X1 U16747 ( .A1(n20492), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13328), .A4(
        n13327), .ZN(U214) );
  NOR4_X1 U16748 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13332) );
  NOR4_X1 U16749 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n13331) );
  NOR4_X1 U16750 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13330) );
  NOR4_X1 U16751 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13329) );
  AND4_X1 U16752 ( .A1(n13332), .A2(n13331), .A3(n13330), .A4(n13329), .ZN(
        n13337) );
  NOR4_X1 U16753 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n13335) );
  NOR4_X1 U16754 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13334) );
  NOR4_X1 U16755 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13333) );
  AND4_X1 U16756 ( .A1(n13335), .A2(n13334), .A3(n13333), .A4(n20189), .ZN(
        n13336) );
  NAND2_X1 U16757 ( .A1(n13337), .A2(n13336), .ZN(n13338) );
  NOR2_X1 U16758 ( .A1(n14365), .A2(n13339), .ZN(n17017) );
  NAND2_X1 U16759 ( .A1(n17017), .A2(U214), .ZN(U212) );
  NAND2_X1 U16760 ( .A1(n20044), .A2(n16742), .ZN(n14058) );
  NAND2_X1 U16761 ( .A1(n20036), .A2(n13340), .ZN(n13341) );
  NAND2_X1 U16762 ( .A1(n14058), .A2(n13341), .ZN(n13342) );
  NAND2_X1 U16763 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n13503) );
  NOR2_X1 U16764 ( .A1(n13503), .A2(n14059), .ZN(n16743) );
  OR2_X1 U16765 ( .A1(n13342), .A2(n16743), .ZN(n13344) );
  NOR2_X1 U16766 ( .A1(n14059), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13343) );
  AND2_X1 U16767 ( .A1(n13343), .A2(n20166), .ZN(n16783) );
  NOR2_X1 U16768 ( .A1(n13344), .A2(n16783), .ZN(P2_U3178) );
  INV_X1 U16769 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21080) );
  INV_X1 U16770 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21083) );
  NOR2_X1 U16771 ( .A1(n21080), .A2(n21083), .ZN(n13345) );
  INV_X1 U16772 ( .A(HOLD), .ZN(n21090) );
  OAI222_X1 U16773 ( .A1(n13345), .A2(P1_STATE_REG_1__SCAN_IN), .B1(n13345), 
        .B2(HOLD), .C1(n21090), .C2(n21092), .ZN(n13347) );
  NAND2_X1 U16774 ( .A1(n13346), .A2(n21080), .ZN(n14012) );
  OAI211_X1 U16775 ( .C1(n21175), .C2(n21086), .A(n13347), .B(n14012), .ZN(
        P1_U3195) );
  NOR2_X1 U16776 ( .A1(n13911), .A2(n19381), .ZN(n13391) );
  NAND2_X1 U16777 ( .A1(n13391), .A2(n13910), .ZN(n15969) );
  INV_X1 U16778 ( .A(n15969), .ZN(n13351) );
  INV_X1 U16779 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n20286) );
  INV_X1 U16780 ( .A(n13348), .ZN(n13350) );
  INV_X1 U16781 ( .A(n20258), .ZN(n20037) );
  NOR2_X1 U16782 ( .A1(n20037), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13355) );
  INV_X1 U16783 ( .A(n13355), .ZN(n13349) );
  OAI211_X1 U16784 ( .C1(n13351), .C2(n20286), .A(n13350), .B(n13349), .ZN(
        P2_U2814) );
  INV_X1 U16785 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n13353) );
  INV_X1 U16786 ( .A(n13352), .ZN(n16785) );
  OAI22_X1 U16787 ( .A1(n13354), .A2(n13353), .B1(n16785), .B2(n20037), .ZN(
        P2_U2816) );
  OAI21_X1 U16788 ( .B1(P2_READREQUEST_REG_SCAN_IN), .B2(n13355), .A(n15576), 
        .ZN(n13356) );
  OAI21_X1 U16789 ( .B1(n13357), .B2(n15576), .A(n13356), .ZN(P2_U3612) );
  INV_X1 U16790 ( .A(P2_UWORD_REG_9__SCAN_IN), .ZN(n13418) );
  INV_X1 U16791 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n17049) );
  OR2_X1 U16792 ( .A1(n14365), .A2(n17049), .ZN(n13359) );
  INV_X2 U16793 ( .A(n16771), .ZN(n14365) );
  NAND2_X1 U16794 ( .A1(n14365), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13358) );
  NAND2_X1 U16795 ( .A1(n13359), .A2(n13358), .ZN(n16092) );
  NAND2_X1 U16796 ( .A1(n19489), .A2(n16092), .ZN(n13367) );
  NAND2_X1 U16797 ( .A1(n19517), .A2(P2_EAX_REG_25__SCAN_IN), .ZN(n13360) );
  OAI211_X1 U16798 ( .C1(n13366), .C2(n13418), .A(n13367), .B(n13360), .ZN(
        P2_U2961) );
  OR2_X1 U16799 ( .A1(n11390), .A2(n10837), .ZN(n13361) );
  INV_X1 U16800 ( .A(n13386), .ZN(n13362) );
  NAND2_X1 U16801 ( .A1(n13473), .A2(n13362), .ZN(n13381) );
  NAND2_X1 U16802 ( .A1(n20934), .A2(n21185), .ZN(n20291) );
  INV_X1 U16803 ( .A(n20291), .ZN(n14646) );
  AOI21_X1 U16804 ( .B1(n14006), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n14646), 
        .ZN(n13363) );
  NAND2_X1 U16805 ( .A1(n14007), .A2(n13363), .ZN(P1_U2801) );
  INV_X1 U16806 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13401) );
  INV_X1 U16807 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n17064) );
  OR2_X1 U16808 ( .A1(n14365), .A2(n17064), .ZN(n13365) );
  NAND2_X1 U16809 ( .A1(n14365), .A2(BUF2_REG_0__SCAN_IN), .ZN(n13364) );
  AND2_X1 U16810 ( .A1(n13365), .A2(n13364), .ZN(n19495) );
  INV_X1 U16811 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13402) );
  OAI222_X1 U16812 ( .A1(n13366), .A2(n13401), .B1(n19520), .B2(n19495), .C1(
        n13392), .C2(n13402), .ZN(P2_U2952) );
  INV_X1 U16813 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19459) );
  NAND2_X1 U16814 ( .A1(n19518), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13368) );
  OAI211_X1 U16815 ( .C1(n19459), .C2(n13392), .A(n13368), .B(n13367), .ZN(
        P2_U2976) );
  NAND2_X1 U16816 ( .A1(n19518), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13372) );
  INV_X1 U16817 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n13369) );
  OR2_X1 U16818 ( .A1(n14365), .A2(n13369), .ZN(n13371) );
  NAND2_X1 U16819 ( .A1(n14365), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13370) );
  NAND2_X1 U16820 ( .A1(n13371), .A2(n13370), .ZN(n14624) );
  NAND2_X1 U16821 ( .A1(n19489), .A2(n14624), .ZN(n13373) );
  OAI211_X1 U16822 ( .C1(n12194), .C2(n13392), .A(n13372), .B(n13373), .ZN(
        P2_U2966) );
  INV_X1 U16823 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19449) );
  NAND2_X1 U16824 ( .A1(n19518), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13374) );
  OAI211_X1 U16825 ( .C1(n19449), .C2(n13392), .A(n13374), .B(n13373), .ZN(
        P2_U2981) );
  INV_X1 U16826 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19457) );
  NAND2_X1 U16827 ( .A1(n19518), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13378) );
  INV_X1 U16828 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n13375) );
  OR2_X1 U16829 ( .A1(n14365), .A2(n13375), .ZN(n13377) );
  NAND2_X1 U16830 ( .A1(n14365), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13376) );
  NAND2_X1 U16831 ( .A1(n13377), .A2(n13376), .ZN(n16084) );
  NAND2_X1 U16832 ( .A1(n19489), .A2(n16084), .ZN(n13379) );
  OAI211_X1 U16833 ( .C1(n19457), .C2(n13392), .A(n13378), .B(n13379), .ZN(
        P2_U2977) );
  INV_X1 U16834 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13416) );
  NAND2_X1 U16835 ( .A1(n19518), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13380) );
  OAI211_X1 U16836 ( .C1(n13416), .C2(n13392), .A(n13380), .B(n13379), .ZN(
        P2_U2962) );
  NAND2_X1 U16837 ( .A1(n16883), .A2(n14647), .ZN(n13383) );
  NAND2_X1 U16838 ( .A1(n13381), .A2(n13304), .ZN(n13382) );
  NAND2_X1 U16839 ( .A1(n13383), .A2(n13382), .ZN(n20289) );
  NAND2_X1 U16840 ( .A1(n9613), .A2(n14012), .ZN(n13468) );
  INV_X1 U16841 ( .A(n13468), .ZN(n13384) );
  AOI21_X1 U16842 ( .B1(n13384), .B2(n14647), .A(n21075), .ZN(n21177) );
  OR2_X1 U16843 ( .A1(n20289), .A2(n21177), .ZN(n16866) );
  AND2_X1 U16844 ( .A1(n16866), .A2(n13718), .ZN(n20294) );
  INV_X1 U16845 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13390) );
  AND3_X1 U16846 ( .A1(n13304), .A2(n16864), .A3(n13721), .ZN(n13385) );
  MUX2_X1 U16847 ( .A(n13470), .B(n13385), .S(n16883), .Z(n13388) );
  NAND2_X1 U16848 ( .A1(n13473), .A2(n13386), .ZN(n13387) );
  NAND2_X1 U16849 ( .A1(n13388), .A2(n13387), .ZN(n16867) );
  NAND2_X1 U16850 ( .A1(n20294), .A2(n16867), .ZN(n13389) );
  OAI21_X1 U16851 ( .B1(n20294), .B2(n13390), .A(n13389), .ZN(P1_U3484) );
  INV_X1 U16852 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13398) );
  INV_X1 U16853 ( .A(n13391), .ZN(n13393) );
  INV_X1 U16854 ( .A(n20173), .ZN(n15568) );
  INV_X1 U16855 ( .A(n13395), .ZN(n13396) );
  INV_X1 U16856 ( .A(P2_UWORD_REG_14__SCAN_IN), .ZN(n13397) );
  OAI222_X1 U16857 ( .A1(n13398), .A2(n19445), .B1(n13433), .B2(n12194), .C1(
        n13434), .C2(n13397), .ZN(P2_U2921) );
  INV_X1 U16858 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n13400) );
  INV_X1 U16859 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n13399) );
  OAI222_X1 U16860 ( .A1(n13400), .A2(n19445), .B1(n13433), .B2(n12168), .C1(
        n13434), .C2(n13399), .ZN(P2_U2933) );
  INV_X1 U16861 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n13403) );
  OAI222_X1 U16862 ( .A1(n13403), .A2(n19445), .B1(n13433), .B2(n13402), .C1(
        n13434), .C2(n13401), .ZN(P2_U2935) );
  INV_X1 U16863 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n13406) );
  INV_X1 U16864 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13405) );
  INV_X1 U16865 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n13404) );
  OAI222_X1 U16866 ( .A1(n13406), .A2(n19445), .B1(n13433), .B2(n13405), .C1(
        n13434), .C2(n13404), .ZN(P2_U2931) );
  INV_X1 U16867 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n13409) );
  INV_X1 U16868 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n13407) );
  OAI222_X1 U16869 ( .A1(n13409), .A2(n19445), .B1(n13433), .B2(n13408), .C1(
        n13434), .C2(n13407), .ZN(P2_U2930) );
  INV_X1 U16870 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n13411) );
  INV_X1 U16871 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n13410) );
  OAI222_X1 U16872 ( .A1(n13411), .A2(n19445), .B1(n13433), .B2(n12177), .C1(
        n13434), .C2(n13410), .ZN(P2_U2929) );
  INV_X1 U16873 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n13414) );
  INV_X1 U16874 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n13412) );
  OAI222_X1 U16875 ( .A1(n13414), .A2(n19445), .B1(n13433), .B2(n13413), .C1(
        n13434), .C2(n13412), .ZN(P2_U2934) );
  INV_X1 U16876 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n13417) );
  INV_X1 U16877 ( .A(P2_UWORD_REG_10__SCAN_IN), .ZN(n13415) );
  OAI222_X1 U16878 ( .A1(n13417), .A2(n19445), .B1(n13433), .B2(n13416), .C1(
        n13434), .C2(n13415), .ZN(P2_U2925) );
  INV_X1 U16879 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n13420) );
  OAI222_X1 U16880 ( .A1(n13420), .A2(n19445), .B1(n13433), .B2(n13419), .C1(
        n13434), .C2(n13418), .ZN(P2_U2926) );
  INV_X1 U16881 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13422) );
  INV_X1 U16882 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n21288) );
  INV_X1 U16883 ( .A(P2_UWORD_REG_12__SCAN_IN), .ZN(n13421) );
  OAI222_X1 U16884 ( .A1(n13422), .A2(n19445), .B1(n13433), .B2(n21288), .C1(
        n13434), .C2(n13421), .ZN(P2_U2923) );
  INV_X1 U16885 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n13425) );
  INV_X1 U16886 ( .A(P2_UWORD_REG_13__SCAN_IN), .ZN(n13423) );
  OAI222_X1 U16887 ( .A1(n13425), .A2(n19445), .B1(n13433), .B2(n13424), .C1(
        n13434), .C2(n13423), .ZN(P2_U2922) );
  OAI21_X1 U16888 ( .B1(n15965), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13443), .ZN(n16720) );
  AOI21_X1 U16889 ( .B1(n13428), .B2(n13427), .A(n13426), .ZN(n16726) );
  INV_X1 U16890 ( .A(n13429), .ZN(n13430) );
  INV_X1 U16891 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19395) );
  NOR2_X1 U16892 ( .A1(n16394), .A2(n19395), .ZN(n16723) );
  AOI211_X1 U16893 ( .C1(n16383), .C2(n16726), .A(n13430), .B(n16723), .ZN(
        n13432) );
  OAI21_X1 U16894 ( .B1(n16410), .B2(n9838), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13431) );
  OAI211_X1 U16895 ( .C1(n16720), .C2(n16439), .A(n13432), .B(n13431), .ZN(
        P2_U3014) );
  INV_X1 U16896 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n16136) );
  INV_X1 U16897 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n17083) );
  INV_X1 U16898 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n21331) );
  OAI222_X1 U16899 ( .A1(n13433), .A2(n16136), .B1(n19445), .B2(n17083), .C1(
        n13434), .C2(n21331), .ZN(P2_U2932) );
  INV_X1 U16900 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n13436) );
  INV_X1 U16901 ( .A(n13433), .ZN(n19443) );
  AOI22_X1 U16902 ( .A1(n19443), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n19476), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13435) );
  OAI21_X1 U16903 ( .B1(n19445), .B2(n13436), .A(n13435), .ZN(P2_U2928) );
  INV_X1 U16904 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n13438) );
  AOI22_X1 U16905 ( .A1(n19443), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n19476), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13437) );
  OAI21_X1 U16906 ( .B1(n19445), .B2(n13438), .A(n13437), .ZN(P2_U2924) );
  AND2_X1 U16907 ( .A1(n16434), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n16711) );
  AOI21_X1 U16908 ( .B1(n13441), .B2(n13440), .A(n13439), .ZN(n16713) );
  INV_X1 U16909 ( .A(n16713), .ZN(n13445) );
  XNOR2_X1 U16910 ( .A(n13442), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13444) );
  XNOR2_X1 U16911 ( .A(n13444), .B(n13443), .ZN(n16709) );
  OAI22_X1 U16912 ( .A1(n13445), .A2(n16429), .B1(n16439), .B2(n16709), .ZN(
        n13446) );
  AOI211_X1 U16913 ( .C1(n16410), .C2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n16711), .B(n13446), .ZN(n13448) );
  NAND2_X1 U16914 ( .A1(n16433), .A2(n15960), .ZN(n13447) );
  INV_X1 U16915 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13451) );
  NOR2_X1 U16916 ( .A1(n10847), .A2(n21175), .ZN(n13449) );
  OR2_X2 U16917 ( .A1(n14007), .A2(n13449), .ZN(n20453) );
  INV_X1 U16918 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20403) );
  MUX2_X1 U16919 ( .A(DATAI_15_), .B(BUF1_REG_15__SCAN_IN), .S(n20492), .Z(
        n15023) );
  INV_X1 U16920 ( .A(n15023), .ZN(n13450) );
  OAI222_X1 U16921 ( .A1(n13588), .A2(n13451), .B1(n13552), .B2(n20403), .C1(
        n13553), .C2(n13450), .ZN(P1_U2967) );
  INV_X1 U16922 ( .A(n13453), .ZN(n13456) );
  AND3_X1 U16923 ( .A1(n13454), .A2(n20524), .A3(n10851), .ZN(n13455) );
  NAND2_X1 U16924 ( .A1(n13456), .A2(n13455), .ZN(n16847) );
  INV_X1 U16925 ( .A(n16847), .ZN(n13487) );
  NAND2_X1 U16926 ( .A1(n13470), .A2(n13721), .ZN(n15531) );
  XNOR2_X1 U16927 ( .A(n13457), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13464) );
  AND2_X1 U16928 ( .A1(n13473), .A2(n20508), .ZN(n15526) );
  XNOR2_X1 U16929 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13460) );
  INV_X1 U16930 ( .A(n13458), .ZN(n13459) );
  NAND2_X1 U16931 ( .A1(n13459), .A2(n16846), .ZN(n15528) );
  OAI22_X1 U16932 ( .A1(n21184), .A2(n13460), .B1(n15528), .B2(n13464), .ZN(
        n13461) );
  AOI21_X1 U16933 ( .B1(n15531), .B2(n13464), .A(n13461), .ZN(n13462) );
  OAI21_X1 U16934 ( .B1(n13452), .B2(n13487), .A(n13462), .ZN(n15536) );
  INV_X1 U16935 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13463) );
  AOI22_X1 U16936 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13727), .B2(n13463), .ZN(
        n13491) );
  NOR2_X1 U16937 ( .A1(n21185), .A2(n13732), .ZN(n13489) );
  INV_X1 U16938 ( .A(n13464), .ZN(n13466) );
  INV_X1 U16939 ( .A(n21186), .ZN(n13465) );
  AOI222_X1 U16940 ( .A1(n15536), .A2(n16985), .B1(n13491), .B2(n13489), .C1(
        n13466), .C2(n13465), .ZN(n13483) );
  OAI211_X1 U16941 ( .C1(n15526), .C2(n10831), .A(n13468), .B(n21175), .ZN(
        n13469) );
  INV_X1 U16942 ( .A(n13469), .ZN(n13471) );
  INV_X1 U16943 ( .A(n13470), .ZN(n13733) );
  MUX2_X1 U16944 ( .A(n13471), .B(n13733), .S(n16883), .Z(n13479) );
  INV_X1 U16945 ( .A(n13472), .ZN(n13474) );
  OR2_X1 U16946 ( .A1(n13474), .A2(n13473), .ZN(n13476) );
  OAI21_X1 U16947 ( .B1(n20512), .B2(n14026), .A(n13716), .ZN(n13477) );
  INV_X1 U16948 ( .A(n16996), .ZN(n16998) );
  NOR2_X1 U16949 ( .A1(n10144), .A2(n16998), .ZN(n15549) );
  AND2_X1 U16950 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n15549), .ZN(n13480) );
  AOI21_X1 U16951 ( .B1(n16849), .B2(n13718), .A(n13480), .ZN(n16988) );
  NAND2_X1 U16952 ( .A1(n10144), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13481) );
  NAND2_X1 U16953 ( .A1(n16988), .A2(n13481), .ZN(n21192) );
  INV_X1 U16954 ( .A(n21192), .ZN(n13496) );
  NAND2_X1 U16955 ( .A1(n13496), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13482) );
  OAI21_X1 U16956 ( .B1(n13483), .B2(n13496), .A(n13482), .ZN(P1_U3472) );
  NOR2_X1 U16957 ( .A1(n13485), .A2(n13457), .ZN(n13488) );
  AOI22_X1 U16958 ( .A1(n15526), .A2(n10600), .B1(n13488), .B2(n16846), .ZN(
        n13486) );
  OAI21_X1 U16959 ( .B1(n13484), .B2(n13487), .A(n13486), .ZN(n16850) );
  INV_X1 U16960 ( .A(n13488), .ZN(n13492) );
  INV_X1 U16961 ( .A(n13489), .ZN(n13490) );
  OAI22_X1 U16962 ( .A1(n21186), .A2(n13492), .B1(n13491), .B2(n13490), .ZN(
        n13493) );
  AOI21_X1 U16963 ( .B1(n16850), .B2(n16985), .A(n13493), .ZN(n13495) );
  NAND2_X1 U16964 ( .A1(n13496), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13494) );
  OAI21_X1 U16965 ( .B1(n13496), .B2(n13495), .A(n13494), .ZN(P1_U3473) );
  NAND2_X1 U16966 ( .A1(n19566), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13497) );
  AOI22_X1 U16967 ( .A1(n13693), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20258), .B2(n20034), .ZN(n13498) );
  NAND4_X1 U16968 ( .A1(n13524), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13499), 
        .A4(n20104), .ZN(n13500) );
  OAI22_X1 U16969 ( .A1(n13501), .A2(n20044), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20104), .ZN(n13502) );
  AOI21_X1 U16970 ( .B1(n19597), .B2(n20255), .A(n13502), .ZN(n13507) );
  INV_X1 U16971 ( .A(n16743), .ZN(n13931) );
  AOI21_X1 U16972 ( .B1(n20275), .B2(n11751), .A(n13931), .ZN(n13506) );
  NOR2_X1 U16973 ( .A1(n20102), .A2(n13506), .ZN(n20272) );
  INV_X1 U16974 ( .A(n20272), .ZN(n20269) );
  MUX2_X1 U16975 ( .A(n20034), .B(n13507), .S(n20269), .Z(n13508) );
  INV_X1 U16976 ( .A(n13508), .ZN(P2_U3605) );
  OAI21_X1 U16977 ( .B1(n14652), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13509), .ZN(n20487) );
  INV_X1 U16978 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13514) );
  NAND2_X1 U16979 ( .A1(n13511), .A2(n13510), .ZN(n13512) );
  NAND2_X1 U16980 ( .A1(n13513), .A2(n13512), .ZN(n14055) );
  OAI222_X1 U16981 ( .A1(n20487), .A2(n14972), .B1(n20396), .B2(n13514), .C1(
        n14055), .C2(n14970), .ZN(P1_U2872) );
  INV_X1 U16982 ( .A(n13905), .ZN(n13515) );
  INV_X1 U16983 ( .A(n13906), .ZN(n13857) );
  NAND2_X1 U16984 ( .A1(n13515), .A2(n13857), .ZN(n13866) );
  NAND2_X1 U16985 ( .A1(n13866), .A2(n9647), .ZN(n13516) );
  NOR2_X1 U16986 ( .A1(n9598), .A2(n13518), .ZN(n13519) );
  AOI21_X1 U16987 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n9598), .A(n13519), .ZN(
        n13520) );
  OAI21_X1 U16988 ( .B1(n16061), .B2(n19522), .A(n13520), .ZN(P2_U2887) );
  NAND2_X1 U16989 ( .A1(n20032), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19855) );
  NAND2_X1 U16990 ( .A1(n20034), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13521) );
  NAND2_X1 U16991 ( .A1(n19855), .A2(n13521), .ZN(n19690) );
  AND2_X1 U16992 ( .A1(n19690), .A2(n20258), .ZN(n19889) );
  AOI21_X1 U16993 ( .B1(n13693), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19889), .ZN(n13522) );
  OAI21_X1 U16994 ( .B1(n19523), .B2(n16061), .A(n13527), .ZN(P2_U2886) );
  XNOR2_X1 U16995 ( .A(n13528), .B(n13529), .ZN(n16687) );
  NAND2_X1 U16996 ( .A1(n12320), .A2(n15574), .ZN(n13914) );
  NOR2_X1 U16997 ( .A1(n13917), .A2(n13914), .ZN(n13530) );
  AOI21_X1 U16998 ( .B1(n13905), .B2(n13904), .A(n13530), .ZN(n13867) );
  NAND2_X1 U16999 ( .A1(n13867), .A2(n13531), .ZN(n13533) );
  INV_X1 U17000 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19463) );
  INV_X1 U17001 ( .A(n13534), .ZN(n13535) );
  NAND2_X1 U17002 ( .A1(n19577), .A2(n19566), .ZN(n13536) );
  INV_X1 U17003 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13537) );
  OR2_X1 U17004 ( .A1(n14365), .A2(n13537), .ZN(n13539) );
  NAND2_X1 U17005 ( .A1(n14365), .A2(BUF2_REG_7__SCAN_IN), .ZN(n13538) );
  AND2_X1 U17006 ( .A1(n13539), .A2(n13538), .ZN(n19508) );
  OAI222_X1 U17007 ( .A1(n16687), .A2(n14084), .B1(n19463), .B2(n16137), .C1(
        n19441), .C2(n19508), .ZN(P2_U2912) );
  INV_X1 U17008 ( .A(n13541), .ZN(n13542) );
  XNOR2_X1 U17009 ( .A(n13540), .B(n13542), .ZN(n19416) );
  INV_X1 U17010 ( .A(n19416), .ZN(n13546) );
  INV_X1 U17011 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19465) );
  INV_X1 U17012 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n13543) );
  OR2_X1 U17013 ( .A1(n14365), .A2(n13543), .ZN(n13545) );
  NAND2_X1 U17014 ( .A1(n14365), .A2(BUF2_REG_6__SCAN_IN), .ZN(n13544) );
  AND2_X1 U17015 ( .A1(n13545), .A2(n13544), .ZN(n19506) );
  OAI222_X1 U17016 ( .A1(n13546), .A2(n14084), .B1(n19465), .B2(n16137), .C1(
        n19441), .C2(n19506), .ZN(P2_U2913) );
  OAI21_X1 U17017 ( .B1(n13548), .B2(n13547), .A(n12018), .ZN(n13549) );
  INV_X1 U17018 ( .A(n13549), .ZN(n16725) );
  NAND2_X1 U17019 ( .A1(n19597), .A2(n16725), .ZN(n19435) );
  OAI211_X1 U17020 ( .C1(n19597), .C2(n16725), .A(n19435), .B(n19437), .ZN(
        n13551) );
  AOI22_X1 U17021 ( .A1(n19433), .A2(n16725), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19431), .ZN(n13550) );
  OAI211_X1 U17022 ( .C1(n19495), .C2(n19441), .A(n13551), .B(n13550), .ZN(
        P2_U2919) );
  AOI22_X1 U17023 ( .A1(n20454), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20453), .ZN(n13554) );
  MUX2_X1 U17024 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n20492), .Z(
        n15028) );
  NAND2_X1 U17025 ( .A1(n20439), .A2(n15028), .ZN(n20451) );
  NAND2_X1 U17026 ( .A1(n13554), .A2(n20451), .ZN(P1_U2950) );
  AOI22_X1 U17027 ( .A1(n20454), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20453), .ZN(n13555) );
  MUX2_X1 U17028 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n20492), .Z(
        n15042) );
  NAND2_X1 U17029 ( .A1(n20439), .A2(n15042), .ZN(n20443) );
  NAND2_X1 U17030 ( .A1(n13555), .A2(n20443), .ZN(P1_U2946) );
  INV_X1 U17031 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13559) );
  NOR2_X4 U17032 ( .A1(n20408), .A2(n21176), .ZN(n20426) );
  AOI22_X1 U17033 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13558) );
  OAI21_X1 U17034 ( .B1(n13559), .B2(n20397), .A(n13558), .ZN(P1_U2918) );
  INV_X1 U17035 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13561) );
  AOI22_X1 U17036 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13560) );
  OAI21_X1 U17037 ( .B1(n13561), .B2(n20397), .A(n13560), .ZN(P1_U2920) );
  INV_X1 U17038 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13563) );
  AOI22_X1 U17039 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13562) );
  OAI21_X1 U17040 ( .B1(n13563), .B2(n20397), .A(n13562), .ZN(P1_U2911) );
  INV_X1 U17041 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13565) );
  AOI22_X1 U17042 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13564) );
  OAI21_X1 U17043 ( .B1(n13565), .B2(n20397), .A(n13564), .ZN(P1_U2915) );
  INV_X1 U17044 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13567) );
  AOI22_X1 U17045 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13566) );
  OAI21_X1 U17046 ( .B1(n13567), .B2(n20397), .A(n13566), .ZN(P1_U2912) );
  INV_X1 U17047 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13569) );
  AOI22_X1 U17048 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13568) );
  OAI21_X1 U17049 ( .B1(n13569), .B2(n20397), .A(n13568), .ZN(P1_U2906) );
  INV_X1 U17050 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13571) );
  AOI22_X1 U17051 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13570) );
  OAI21_X1 U17052 ( .B1(n13571), .B2(n20397), .A(n13570), .ZN(P1_U2914) );
  AOI22_X1 U17053 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13572) );
  OAI21_X1 U17054 ( .B1(n11221), .B2(n20397), .A(n13572), .ZN(P1_U2919) );
  AOI22_X1 U17055 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13573) );
  OAI21_X1 U17056 ( .B1(n11367), .B2(n20397), .A(n13573), .ZN(P1_U2909) );
  INV_X1 U17057 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13575) );
  AOI22_X1 U17058 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13574) );
  OAI21_X1 U17059 ( .B1(n13575), .B2(n20397), .A(n13574), .ZN(P1_U2913) );
  INV_X1 U17060 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13577) );
  AOI22_X1 U17061 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13576) );
  OAI21_X1 U17062 ( .B1(n13577), .B2(n20397), .A(n13576), .ZN(P1_U2908) );
  INV_X1 U17063 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13579) );
  AOI22_X1 U17064 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13578) );
  OAI21_X1 U17065 ( .B1(n13579), .B2(n20397), .A(n13578), .ZN(P1_U2907) );
  INV_X1 U17066 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13581) );
  AOI22_X1 U17067 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13580) );
  OAI21_X1 U17068 ( .B1(n13581), .B2(n20397), .A(n13580), .ZN(P1_U2917) );
  AOI22_X1 U17069 ( .A1(n20454), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20453), .ZN(n13584) );
  INV_X1 U17070 ( .A(DATAI_6_), .ZN(n13583) );
  NAND2_X1 U17071 ( .A1(n20492), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13582) );
  OAI21_X1 U17072 ( .B1(n20492), .B2(n13583), .A(n13582), .ZN(n14997) );
  NAND2_X1 U17073 ( .A1(n20439), .A2(n14997), .ZN(n13589) );
  NAND2_X1 U17074 ( .A1(n13584), .A2(n13589), .ZN(P1_U2943) );
  AOI22_X1 U17075 ( .A1(n20454), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20453), .ZN(n13587) );
  INV_X1 U17076 ( .A(DATAI_2_), .ZN(n13586) );
  NAND2_X1 U17077 ( .A1(n20492), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13585) );
  OAI21_X1 U17078 ( .B1(n20492), .B2(n13586), .A(n13585), .ZN(n15011) );
  NAND2_X1 U17079 ( .A1(n20439), .A2(n15011), .ZN(n13605) );
  NAND2_X1 U17080 ( .A1(n13587), .A2(n13605), .ZN(P1_U2939) );
  INV_X2 U17081 ( .A(n13588), .ZN(n20454) );
  AOI22_X1 U17082 ( .A1(n20454), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20453), .ZN(n13590) );
  NAND2_X1 U17083 ( .A1(n13590), .A2(n13589), .ZN(P1_U2958) );
  AOI22_X1 U17084 ( .A1(n20454), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20453), .ZN(n13593) );
  INV_X1 U17085 ( .A(DATAI_3_), .ZN(n13592) );
  NAND2_X1 U17086 ( .A1(n20492), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13591) );
  OAI21_X1 U17087 ( .B1(n20492), .B2(n13592), .A(n13591), .ZN(n15008) );
  NAND2_X1 U17088 ( .A1(n20439), .A2(n15008), .ZN(n13609) );
  NAND2_X1 U17089 ( .A1(n13593), .A2(n13609), .ZN(P1_U2940) );
  AOI22_X1 U17090 ( .A1(n20454), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20453), .ZN(n13596) );
  INV_X1 U17091 ( .A(DATAI_7_), .ZN(n13595) );
  NAND2_X1 U17092 ( .A1(n20492), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13594) );
  OAI21_X1 U17093 ( .B1(n20492), .B2(n13595), .A(n13594), .ZN(n14993) );
  NAND2_X1 U17094 ( .A1(n20439), .A2(n14993), .ZN(n13597) );
  NAND2_X1 U17095 ( .A1(n13596), .A2(n13597), .ZN(P1_U2959) );
  AOI22_X1 U17096 ( .A1(n20454), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20453), .ZN(n13598) );
  NAND2_X1 U17097 ( .A1(n13598), .A2(n13597), .ZN(P1_U2944) );
  AOI22_X1 U17098 ( .A1(n20454), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20453), .ZN(n13601) );
  INV_X1 U17099 ( .A(DATAI_0_), .ZN(n13600) );
  NAND2_X1 U17100 ( .A1(n20492), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13599) );
  OAI21_X1 U17101 ( .B1(n20492), .B2(n13600), .A(n13599), .ZN(n15019) );
  NAND2_X1 U17102 ( .A1(n20439), .A2(n15019), .ZN(n13621) );
  NAND2_X1 U17103 ( .A1(n13601), .A2(n13621), .ZN(P1_U2952) );
  AOI22_X1 U17104 ( .A1(n20454), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20453), .ZN(n13604) );
  INV_X1 U17105 ( .A(DATAI_1_), .ZN(n13603) );
  NAND2_X1 U17106 ( .A1(n20492), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13602) );
  OAI21_X1 U17107 ( .B1(n20492), .B2(n13603), .A(n13602), .ZN(n15014) );
  NAND2_X1 U17108 ( .A1(n20439), .A2(n15014), .ZN(n13607) );
  NAND2_X1 U17109 ( .A1(n13604), .A2(n13607), .ZN(P1_U2953) );
  AOI22_X1 U17110 ( .A1(n20454), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20453), .ZN(n13606) );
  NAND2_X1 U17111 ( .A1(n13606), .A2(n13605), .ZN(P1_U2954) );
  AOI22_X1 U17112 ( .A1(n20454), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20453), .ZN(n13608) );
  NAND2_X1 U17113 ( .A1(n13608), .A2(n13607), .ZN(P1_U2938) );
  AOI22_X1 U17114 ( .A1(n20454), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20453), .ZN(n13610) );
  NAND2_X1 U17115 ( .A1(n13610), .A2(n13609), .ZN(P1_U2955) );
  AOI22_X1 U17116 ( .A1(n20454), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20453), .ZN(n13613) );
  INV_X1 U17117 ( .A(DATAI_4_), .ZN(n13612) );
  NAND2_X1 U17118 ( .A1(n20492), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13611) );
  OAI21_X1 U17119 ( .B1(n20492), .B2(n13612), .A(n13611), .ZN(n15005) );
  NAND2_X1 U17120 ( .A1(n20439), .A2(n15005), .ZN(n13617) );
  NAND2_X1 U17121 ( .A1(n13613), .A2(n13617), .ZN(P1_U2956) );
  AOI22_X1 U17122 ( .A1(n20454), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20453), .ZN(n13616) );
  INV_X1 U17123 ( .A(DATAI_5_), .ZN(n13615) );
  NAND2_X1 U17124 ( .A1(n20492), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13614) );
  OAI21_X1 U17125 ( .B1(n20492), .B2(n13615), .A(n13614), .ZN(n15001) );
  NAND2_X1 U17126 ( .A1(n20439), .A2(n15001), .ZN(n13619) );
  NAND2_X1 U17127 ( .A1(n13616), .A2(n13619), .ZN(P1_U2942) );
  AOI22_X1 U17128 ( .A1(n20454), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20453), .ZN(n13618) );
  NAND2_X1 U17129 ( .A1(n13618), .A2(n13617), .ZN(P1_U2941) );
  AOI22_X1 U17130 ( .A1(n20454), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20453), .ZN(n13620) );
  NAND2_X1 U17131 ( .A1(n13620), .A2(n13619), .ZN(P1_U2957) );
  AOI22_X1 U17132 ( .A1(n20454), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20453), .ZN(n13622) );
  NAND2_X1 U17133 ( .A1(n13622), .A2(n13621), .ZN(P1_U2937) );
  NAND2_X1 U17134 ( .A1(n13624), .A2(n13623), .ZN(n13625) );
  AOI21_X1 U17135 ( .B1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13628) );
  NOR2_X1 U17136 ( .A1(n13694), .A2(n13628), .ZN(n19697) );
  AND2_X1 U17137 ( .A1(n19697), .A2(n20258), .ZN(n16773) );
  AOI21_X1 U17138 ( .B1(n13693), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n16773), .ZN(n13629) );
  NAND2_X1 U17139 ( .A1(n13632), .A2(n13631), .ZN(n13692) );
  OAI21_X1 U17140 ( .B1(n20264), .B2(n16061), .A(n13635), .ZN(P2_U2885) );
  NAND2_X1 U17141 ( .A1(n13638), .A2(n13637), .ZN(n13639) );
  AND2_X1 U17142 ( .A1(n13636), .A2(n13639), .ZN(n16672) );
  INV_X1 U17143 ( .A(n16672), .ZN(n13644) );
  INV_X1 U17144 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n13640) );
  OR2_X1 U17145 ( .A1(n14365), .A2(n13640), .ZN(n13642) );
  NAND2_X1 U17146 ( .A1(n14365), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13641) );
  NAND2_X1 U17147 ( .A1(n13642), .A2(n13641), .ZN(n19488) );
  AOI22_X1 U17148 ( .A1(n14122), .A2(n19488), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n19431), .ZN(n13643) );
  OAI21_X1 U17149 ( .B1(n13644), .B2(n14084), .A(n13643), .ZN(P2_U2911) );
  OR2_X1 U17150 ( .A1(n20570), .A2(n13645), .ZN(n13648) );
  NAND4_X1 U17151 ( .A1(n13648), .A2(n13647), .A3(n13646), .A4(n13732), .ZN(
        n13650) );
  NAND2_X1 U17152 ( .A1(n13650), .A2(n13649), .ZN(n20482) );
  INV_X1 U17153 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13651) );
  OR2_X1 U17154 ( .A1(n20348), .A2(n13651), .ZN(n20484) );
  OAI21_X1 U17155 ( .B1(n16921), .B2(n13652), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13653) );
  OAI211_X1 U17156 ( .C1(n20482), .C2(n20293), .A(n20484), .B(n13653), .ZN(
        n13654) );
  INV_X1 U17157 ( .A(n13654), .ZN(n13655) );
  OAI21_X1 U17158 ( .B1(n20491), .B2(n14055), .A(n13655), .ZN(P1_U2999) );
  MUX2_X1 U17159 ( .A(n14318), .B(n13656), .S(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n13674) );
  INV_X1 U17160 ( .A(n13657), .ZN(n13672) );
  OR2_X1 U17161 ( .A1(n13659), .A2(n13658), .ZN(n13660) );
  NAND2_X1 U17162 ( .A1(n13661), .A2(n13660), .ZN(n20268) );
  NAND2_X1 U17163 ( .A1(n16434), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n14635) );
  INV_X1 U17164 ( .A(n13662), .ZN(n14643) );
  NOR2_X1 U17165 ( .A1(n13664), .A2(n13663), .ZN(n14642) );
  NOR3_X1 U17166 ( .A1(n16721), .A2(n14643), .A3(n14642), .ZN(n13665) );
  AOI211_X1 U17167 ( .C1(n16724), .C2(n20268), .A(n13666), .B(n13665), .ZN(
        n13670) );
  OR2_X1 U17168 ( .A1(n9674), .A2(n13667), .ZN(n14638) );
  NAND3_X1 U17169 ( .A1(n12739), .A2(n14637), .A3(n14638), .ZN(n13668) );
  NAND3_X1 U17170 ( .A1(n13670), .A2(n13669), .A3(n13668), .ZN(n13671) );
  AOI21_X1 U17171 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n13672), .A(
        n13671), .ZN(n13673) );
  OAI21_X1 U17172 ( .B1(n16715), .B2(n13674), .A(n13673), .ZN(P2_U3044) );
  OR2_X1 U17173 ( .A1(n13636), .A2(n13681), .ZN(n13679) );
  NAND2_X1 U17174 ( .A1(n13679), .A2(n13676), .ZN(n13677) );
  NAND2_X1 U17175 ( .A1(n13675), .A2(n13677), .ZN(n16642) );
  AOI22_X1 U17176 ( .A1(n14122), .A2(n16084), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n19431), .ZN(n13678) );
  OAI21_X1 U17177 ( .B1(n16642), .B2(n14084), .A(n13678), .ZN(P2_U2909) );
  INV_X1 U17178 ( .A(n13679), .ZN(n13680) );
  AOI21_X1 U17179 ( .B1(n13681), .B2(n13636), .A(n13680), .ZN(n16652) );
  INV_X1 U17180 ( .A(n16652), .ZN(n13683) );
  AOI22_X1 U17181 ( .A1(n14122), .A2(n16092), .B1(P2_EAX_REG_9__SCAN_IN), .B2(
        n19431), .ZN(n13682) );
  OAI21_X1 U17182 ( .B1(n13683), .B2(n14084), .A(n13682), .ZN(P2_U2910) );
  OAI21_X1 U17183 ( .B1(n13685), .B2(n13684), .A(n13811), .ZN(n14049) );
  XNOR2_X1 U17184 ( .A(n14041), .B(n9613), .ZN(n13737) );
  INV_X1 U17185 ( .A(n13737), .ZN(n13686) );
  AOI22_X1 U17186 ( .A1(n20391), .A2(n13686), .B1(n14968), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13687) );
  OAI21_X1 U17187 ( .B1(n14049), .B2(n14970), .A(n13687), .ZN(P1_U2871) );
  INV_X1 U17188 ( .A(n13688), .ZN(n13689) );
  NAND2_X1 U17189 ( .A1(n13690), .A2(n13689), .ZN(n13691) );
  NAND2_X1 U17190 ( .A1(n13692), .A2(n13691), .ZN(n13764) );
  NAND2_X1 U17191 ( .A1(n13693), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13696) );
  OAI211_X1 U17192 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n13694), .A(
        n20155), .B(n20258), .ZN(n13695) );
  INV_X1 U17193 ( .A(n13766), .ZN(n13698) );
  NAND2_X1 U17194 ( .A1(n14556), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13699) );
  NAND2_X1 U17195 ( .A1(n13698), .A2(n13699), .ZN(n13701) );
  INV_X1 U17196 ( .A(n13699), .ZN(n13700) );
  NAND2_X1 U17197 ( .A1(n13766), .A2(n13700), .ZN(n13767) );
  MUX2_X1 U17198 ( .A(n13703), .B(n13702), .S(n9598), .Z(n13704) );
  OAI21_X1 U17199 ( .B1(n19598), .B2(n16061), .A(n13704), .ZN(P2_U2884) );
  NAND2_X1 U17200 ( .A1(n20508), .A2(n14012), .ZN(n13705) );
  NAND2_X1 U17201 ( .A1(n13706), .A2(n13705), .ZN(n13714) );
  OAI21_X1 U17202 ( .B1(n13707), .B2(n21075), .A(n10837), .ZN(n13710) );
  NAND2_X1 U17203 ( .A1(n10847), .A2(n14012), .ZN(n13709) );
  AOI21_X1 U17204 ( .B1(n13710), .B2(n13709), .A(n13708), .ZN(n13711) );
  MUX2_X1 U17205 ( .A(n13714), .B(n13713), .S(n13712), .Z(n13717) );
  NAND3_X1 U17206 ( .A1(n16883), .A2(n16846), .A3(n20508), .ZN(n13715) );
  NAND3_X1 U17207 ( .A1(n13717), .A2(n13716), .A3(n13715), .ZN(n13719) );
  INV_X1 U17208 ( .A(n13738), .ZN(n13725) );
  OAI211_X1 U17209 ( .C1(n13722), .C2(n13728), .A(n13721), .B(n16864), .ZN(
        n13723) );
  NOR2_X1 U17210 ( .A1(n13720), .A2(n13723), .ZN(n13724) );
  XNOR2_X1 U17211 ( .A(n13726), .B(n13727), .ZN(n13952) );
  OR2_X1 U17212 ( .A1(n13304), .A2(n20508), .ZN(n16877) );
  OAI21_X1 U17213 ( .B1(n13728), .B2(n20520), .A(n16877), .ZN(n13729) );
  NOR2_X1 U17214 ( .A1(n13738), .A2(n16962), .ZN(n20478) );
  INV_X1 U17215 ( .A(n13730), .ZN(n13731) );
  NAND2_X1 U17216 ( .A1(n15382), .A2(n13732), .ZN(n13750) );
  OR2_X1 U17217 ( .A1(n16939), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13734) );
  NAND2_X1 U17218 ( .A1(n13750), .A2(n13734), .ZN(n20476) );
  OAI21_X1 U17219 ( .B1(n20478), .B2(n20476), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13736) );
  INV_X1 U17220 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21162) );
  NOR2_X1 U17221 ( .A1(n20348), .A2(n21162), .ZN(n13951) );
  INV_X1 U17222 ( .A(n13951), .ZN(n13735) );
  OAI211_X1 U17223 ( .C1(n20486), .C2(n13737), .A(n13736), .B(n13735), .ZN(
        n13740) );
  INV_X1 U17224 ( .A(n16944), .ZN(n15269) );
  NOR3_X1 U17225 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n15269), .A3(
        n13760), .ZN(n13739) );
  AOI211_X1 U17226 ( .C1(n16965), .C2(n13952), .A(n13740), .B(n13739), .ZN(
        n13741) );
  INV_X1 U17227 ( .A(n13741), .ZN(P1_U3030) );
  INV_X1 U17228 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19455) );
  INV_X1 U17229 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13742) );
  OR2_X1 U17230 ( .A1(n14365), .A2(n13742), .ZN(n13744) );
  NAND2_X1 U17231 ( .A1(n14365), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13743) );
  AND2_X1 U17232 ( .A1(n13744), .A2(n13743), .ZN(n19512) );
  XNOR2_X1 U17233 ( .A(n13675), .B(n13745), .ZN(n16628) );
  OAI222_X1 U17234 ( .A1(n16137), .A2(n19455), .B1(n19512), .B2(n19441), .C1(
        n16628), .C2(n14084), .ZN(P2_U2908) );
  NAND2_X1 U17235 ( .A1(n13746), .A2(n20532), .ZN(n13747) );
  INV_X1 U17236 ( .A(n15014), .ZN(n20509) );
  OAI222_X1 U17237 ( .A1(n14049), .A2(n15045), .B1(n15034), .B2(n20509), .C1(
        n15031), .C2(n10977), .ZN(P1_U2903) );
  INV_X1 U17238 ( .A(n15019), .ZN(n20501) );
  INV_X1 U17239 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20429) );
  OAI222_X1 U17240 ( .A1(n14055), .A2(n15045), .B1(n15034), .B2(n20501), .C1(
        n15031), .C2(n20429), .ZN(P1_U2904) );
  XNOR2_X1 U17241 ( .A(n13749), .B(n13748), .ZN(n13943) );
  NAND2_X1 U17242 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13753) );
  INV_X1 U17243 ( .A(n20478), .ZN(n13751) );
  NAND2_X1 U17244 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15476) );
  NAND2_X1 U17245 ( .A1(n16942), .A2(n15476), .ZN(n13752) );
  OAI21_X1 U17246 ( .B1(n16939), .B2(n13753), .A(n15493), .ZN(n13759) );
  AND2_X1 U17247 ( .A1(n16962), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n13758) );
  AOI21_X1 U17248 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20459) );
  INV_X1 U17249 ( .A(n20459), .ZN(n16970) );
  NOR2_X1 U17250 ( .A1(n13755), .A2(n13754), .ZN(n13756) );
  OR2_X1 U17251 ( .A1(n13787), .A2(n13756), .ZN(n14020) );
  OAI22_X1 U17252 ( .A1(n16939), .A2(n16970), .B1(n20486), .B2(n14020), .ZN(
        n13757) );
  AOI211_X1 U17253 ( .C1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n13759), .A(
        n13758), .B(n13757), .ZN(n13762) );
  INV_X1 U17254 ( .A(n15478), .ZN(n16943) );
  OR3_X1 U17255 ( .A1(n13727), .A2(n16943), .A3(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13761) );
  OAI211_X1 U17256 ( .C1(n20481), .C2(n13943), .A(n13762), .B(n13761), .ZN(
        P1_U3029) );
  NAND2_X1 U17257 ( .A1(n19566), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13765) );
  AND2_X1 U17258 ( .A1(n14556), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13768) );
  NAND2_X1 U17259 ( .A1(n13821), .A2(n13768), .ZN(n13841) );
  INV_X1 U17260 ( .A(n13767), .ZN(n13769) );
  OR3_X1 U17261 ( .A1(n13770), .A2(n13769), .A3(n13768), .ZN(n13771) );
  NAND2_X1 U17262 ( .A1(n13841), .A2(n13771), .ZN(n15921) );
  NAND2_X1 U17263 ( .A1(n13773), .A2(n13772), .ZN(n13774) );
  AND2_X1 U17264 ( .A1(n13804), .A2(n13774), .ZN(n15918) );
  INV_X1 U17265 ( .A(n15918), .ZN(n14157) );
  NOR2_X1 U17266 ( .A1(n14157), .A2(n9598), .ZN(n13775) );
  AOI21_X1 U17267 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n9598), .A(n13775), .ZN(
        n13776) );
  OAI21_X1 U17268 ( .B1(n15921), .B2(n16061), .A(n13776), .ZN(P2_U2883) );
  OR2_X1 U17269 ( .A1(n13779), .A2(n13778), .ZN(n13780) );
  NAND2_X1 U17270 ( .A1(n13777), .A2(n13780), .ZN(n16623) );
  INV_X1 U17271 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19453) );
  INV_X1 U17272 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n13781) );
  OR2_X1 U17273 ( .A1(n14365), .A2(n13781), .ZN(n13783) );
  NAND2_X1 U17274 ( .A1(n14365), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13782) );
  AND2_X1 U17275 ( .A1(n13783), .A2(n13782), .ZN(n19514) );
  OAI222_X1 U17276 ( .A1(n16623), .A2(n14084), .B1(n16137), .B2(n19453), .C1(
        n19441), .C2(n19514), .ZN(P2_U2907) );
  NAND2_X1 U17277 ( .A1(n13785), .A2(n13784), .ZN(n13985) );
  OAI21_X1 U17278 ( .B1(n13785), .B2(n13784), .A(n13985), .ZN(n13945) );
  OR2_X1 U17279 ( .A1(n13787), .A2(n13786), .ZN(n13788) );
  AND2_X1 U17280 ( .A1(n16974), .A2(n13788), .ZN(n20472) );
  AOI22_X1 U17281 ( .A1(n20391), .A2(n20472), .B1(n14968), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n13789) );
  OAI21_X1 U17282 ( .B1(n13945), .B2(n14970), .A(n13789), .ZN(P1_U2869) );
  INV_X1 U17283 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n17058) );
  OR2_X1 U17284 ( .A1(n14365), .A2(n17058), .ZN(n13791) );
  NAND2_X1 U17285 ( .A1(n14365), .A2(BUF2_REG_2__SCAN_IN), .ZN(n13790) );
  AND2_X1 U17286 ( .A1(n13791), .A2(n13790), .ZN(n19499) );
  XNOR2_X1 U17287 ( .A(n20264), .B(n20268), .ZN(n13799) );
  OR2_X1 U17288 ( .A1(n13793), .A2(n13792), .ZN(n13795) );
  NAND2_X1 U17289 ( .A1(n13795), .A2(n13794), .ZN(n19432) );
  NOR2_X1 U17290 ( .A1(n20254), .A2(n19432), .ZN(n13796) );
  AOI21_X1 U17291 ( .B1(n20254), .B2(n19432), .A(n13796), .ZN(n19436) );
  NAND2_X1 U17292 ( .A1(n19436), .A2(n19435), .ZN(n19434) );
  INV_X1 U17293 ( .A(n13796), .ZN(n13797) );
  NAND2_X1 U17294 ( .A1(n19434), .A2(n13797), .ZN(n13798) );
  NAND2_X1 U17295 ( .A1(n13798), .A2(n13799), .ZN(n14075) );
  OAI21_X1 U17296 ( .B1(n13799), .B2(n13798), .A(n14075), .ZN(n13800) );
  NAND2_X1 U17297 ( .A1(n13800), .A2(n19437), .ZN(n13802) );
  AOI22_X1 U17298 ( .A1(n19433), .A2(n20268), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19431), .ZN(n13801) );
  OAI211_X1 U17299 ( .C1(n19441), .C2(n19499), .A(n13802), .B(n13801), .ZN(
        P2_U2917) );
  XOR2_X1 U17300 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13841), .Z(n13807)
         );
  NAND2_X1 U17301 ( .A1(n13804), .A2(n13803), .ZN(n13805) );
  NAND2_X1 U17302 ( .A1(n13845), .A2(n13805), .ZN(n15894) );
  MUX2_X1 U17303 ( .A(n15894), .B(n12380), .S(n9598), .Z(n13806) );
  OAI21_X1 U17304 ( .B1(n13807), .B2(n16061), .A(n13806), .ZN(P2_U2882) );
  INV_X1 U17305 ( .A(n15008), .ZN(n20517) );
  OAI222_X1 U17306 ( .A1(n13945), .A2(n15045), .B1(n15034), .B2(n20517), .C1(
        n15031), .C2(n11002), .ZN(P1_U2901) );
  INV_X1 U17307 ( .A(n13808), .ZN(n13809) );
  AOI21_X1 U17308 ( .B1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n13810), .A(
        n13809), .ZN(n13814) );
  INV_X1 U17309 ( .A(n13811), .ZN(n13813) );
  NAND2_X1 U17310 ( .A1(n13814), .A2(n13813), .ZN(n13812) );
  OAI21_X1 U17311 ( .B1(n13814), .B2(n13813), .A(n13812), .ZN(n14035) );
  INV_X1 U17312 ( .A(n14020), .ZN(n13815) );
  AOI22_X1 U17313 ( .A1(n20391), .A2(n13815), .B1(n14968), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13816) );
  OAI21_X1 U17314 ( .B1(n14035), .B2(n14970), .A(n13816), .ZN(P1_U2870) );
  AND2_X1 U17315 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13833) );
  NAND3_X1 U17316 ( .A1(n13833), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13817) );
  NOR2_X1 U17317 ( .A1(n13955), .A2(n13817), .ZN(n13819) );
  AND3_X1 U17318 ( .A1(n14556), .A2(n13819), .A3(n13818), .ZN(n13820) );
  INV_X1 U17319 ( .A(n13822), .ZN(n13825) );
  OAI211_X1 U17320 ( .C1(n13825), .C2(n13824), .A(n16036), .B(n14190), .ZN(
        n13832) );
  OR2_X1 U17321 ( .A1(n13827), .A2(n13828), .ZN(n13829) );
  NAND2_X1 U17322 ( .A1(n13826), .A2(n13829), .ZN(n16646) );
  INV_X1 U17323 ( .A(n16646), .ZN(n13830) );
  NAND2_X1 U17324 ( .A1(n13830), .A2(n16058), .ZN(n13831) );
  OAI211_X1 U17325 ( .C1(n16058), .C2(n12426), .A(n13832), .B(n13831), .ZN(
        P2_U2877) );
  INV_X1 U17326 ( .A(n13833), .ZN(n13834) );
  NOR2_X1 U17327 ( .A1(n13841), .A2(n13834), .ZN(n13954) );
  XNOR2_X1 U17328 ( .A(n13954), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13840) );
  OR2_X1 U17329 ( .A1(n9748), .A2(n13836), .ZN(n13837) );
  AND2_X1 U17330 ( .A1(n13835), .A2(n13837), .ZN(n16685) );
  NOR2_X1 U17331 ( .A1(n16058), .A2(n12413), .ZN(n13838) );
  AOI21_X1 U17332 ( .B1(n16685), .B2(n16058), .A(n13838), .ZN(n13839) );
  OAI21_X1 U17333 ( .B1(n13840), .B2(n16061), .A(n13839), .ZN(P2_U2880) );
  INV_X1 U17334 ( .A(n15011), .ZN(n20513) );
  OAI222_X1 U17335 ( .A1(n14035), .A2(n15045), .B1(n15034), .B2(n20513), .C1(
        n15031), .C2(n10970), .ZN(P1_U2902) );
  INV_X1 U17336 ( .A(n13841), .ZN(n13842) );
  AOI21_X1 U17337 ( .B1(n13842), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13843) );
  NOR3_X1 U17338 ( .A1(n13843), .A2(n13954), .A3(n16061), .ZN(n13848) );
  AND2_X1 U17339 ( .A1(n13845), .A2(n13844), .ZN(n13846) );
  NOR2_X1 U17340 ( .A1(n9748), .A2(n13846), .ZN(n19415) );
  MUX2_X1 U17341 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n19415), .S(n16058), .Z(
        n13847) );
  OR2_X1 U17342 ( .A1(n13848), .A2(n13847), .ZN(P2_U2881) );
  INV_X1 U17343 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19451) );
  INV_X1 U17344 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13849) );
  OR2_X1 U17345 ( .A1(n14365), .A2(n13849), .ZN(n13851) );
  NAND2_X1 U17346 ( .A1(n14365), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13850) );
  AND2_X1 U17347 ( .A1(n13851), .A2(n13850), .ZN(n19516) );
  XOR2_X1 U17348 ( .A(n13777), .B(n13852), .Z(n16611) );
  INV_X1 U17349 ( .A(n16611), .ZN(n13853) );
  OAI222_X1 U17350 ( .A1(n16137), .A2(n19451), .B1(n19516), .B2(n19441), .C1(
        n13853), .C2(n14084), .ZN(P2_U2906) );
  NAND2_X1 U17351 ( .A1(n9647), .A2(n12315), .ZN(n13858) );
  NAND2_X1 U17352 ( .A1(n13858), .A2(n13854), .ZN(n13856) );
  NAND2_X1 U17353 ( .A1(n13892), .A2(n13859), .ZN(n13855) );
  NAND2_X1 U17354 ( .A1(n13856), .A2(n13855), .ZN(n13877) );
  NOR2_X1 U17355 ( .A1(n13887), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13876) );
  OR2_X1 U17356 ( .A1(n13857), .A2(n13904), .ZN(n13875) );
  OAI21_X1 U17357 ( .B1(n14611), .B2(n13876), .A(n13875), .ZN(n13862) );
  NAND3_X1 U17358 ( .A1(n13858), .A2(n13887), .A3(n13854), .ZN(n13861) );
  NAND3_X1 U17359 ( .A1(n13892), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        n13859), .ZN(n13860) );
  NAND3_X1 U17360 ( .A1(n13862), .A2(n13861), .A3(n13860), .ZN(n13864) );
  AOI211_X1 U17361 ( .C1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(n13877), .A(
        n13864), .B(n13863), .ZN(n16758) );
  INV_X1 U17362 ( .A(n16758), .ZN(n13872) );
  AND3_X1 U17363 ( .A1(n13867), .A2(n13866), .A3(n13865), .ZN(n13871) );
  INV_X1 U17364 ( .A(n13868), .ZN(n13869) );
  INV_X1 U17365 ( .A(n13911), .ZN(n16812) );
  NAND3_X1 U17366 ( .A1(n13869), .A2(n16812), .A3(n13916), .ZN(n13870) );
  MUX2_X1 U17367 ( .A(n13872), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n16744), .Z(n13923) );
  INV_X1 U17368 ( .A(n13923), .ZN(n13899) );
  NAND2_X1 U17369 ( .A1(n15933), .A2(n9840), .ZN(n13883) );
  INV_X1 U17370 ( .A(n13876), .ZN(n13874) );
  AOI22_X1 U17371 ( .A1(n13875), .A2(n13874), .B1(n11581), .B2(n13892), .ZN(
        n13879) );
  NOR2_X1 U17372 ( .A1(n13877), .A2(n13876), .ZN(n13878) );
  MUX2_X1 U17373 ( .A(n13879), .B(n13878), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13881) );
  INV_X1 U17374 ( .A(n14471), .ZN(n13880) );
  AND2_X1 U17375 ( .A1(n13881), .A2(n13880), .ZN(n13882) );
  NAND2_X1 U17376 ( .A1(n13883), .A2(n13882), .ZN(n16762) );
  MUX2_X1 U17377 ( .A(n16762), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n16744), .Z(n13922) );
  INV_X1 U17378 ( .A(n13922), .ZN(n13898) );
  OAI21_X1 U17379 ( .B1(n13899), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n13898), .ZN(n13902) );
  INV_X1 U17380 ( .A(n13884), .ZN(n13886) );
  NAND2_X1 U17381 ( .A1(n13886), .A2(n13885), .ZN(n13893) );
  NOR2_X1 U17382 ( .A1(n11579), .A2(n13887), .ZN(n13889) );
  AOI22_X1 U17383 ( .A1(n13893), .A2(n13889), .B1(n13888), .B2(n13892), .ZN(
        n13890) );
  INV_X1 U17384 ( .A(n16755), .ZN(n13895) );
  MUX2_X1 U17385 ( .A(n13893), .B(n13892), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n13894) );
  AOI21_X1 U17386 ( .B1(n9836), .B2(n9840), .A(n13894), .ZN(n16741) );
  OAI211_X1 U17387 ( .C1(n13895), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16741), .ZN(n13896) );
  INV_X1 U17388 ( .A(n16744), .ZN(n13920) );
  OAI211_X1 U17389 ( .C1(n20032), .C2(n16755), .A(n13896), .B(n13920), .ZN(
        n13897) );
  AOI21_X1 U17390 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13898), .A(
        n13897), .ZN(n13901) );
  NAND2_X1 U17391 ( .A1(n13899), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13900) );
  AOI22_X1 U17392 ( .A1(n13902), .A2(n20262), .B1(n13901), .B2(n13900), .ZN(
        n13925) );
  INV_X1 U17393 ( .A(n13903), .ZN(n13909) );
  INV_X1 U17394 ( .A(n13904), .ZN(n13907) );
  MUX2_X1 U17395 ( .A(n13907), .B(n13906), .S(n13905), .Z(n13908) );
  OAI21_X1 U17396 ( .B1(n13910), .B2(n13909), .A(n13908), .ZN(n20274) );
  AOI21_X1 U17397 ( .B1(n13913), .B2(n16778), .A(n13912), .ZN(n13919) );
  INV_X1 U17398 ( .A(n13914), .ZN(n13915) );
  NOR3_X1 U17399 ( .A1(n13917), .A2(n13916), .A3(n13915), .ZN(n19382) );
  OAI21_X1 U17400 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n19382), .ZN(n13918) );
  OAI211_X1 U17401 ( .C1(n13920), .C2(n11639), .A(n13919), .B(n13918), .ZN(
        n13921) );
  AOI211_X1 U17402 ( .C1(n13923), .C2(n13922), .A(n20274), .B(n13921), .ZN(
        n13924) );
  OAI21_X1 U17403 ( .B1(n13925), .B2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n13924), .ZN(n14056) );
  OAI21_X1 U17404 ( .B1(n14056), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n13930) );
  NOR2_X1 U17405 ( .A1(n13926), .A2(n20044), .ZN(n15577) );
  NAND3_X1 U17406 ( .A1(n11823), .A2(n13928), .A3(n13927), .ZN(n13929) );
  OAI21_X1 U17407 ( .B1(n14057), .B2(n14059), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13932) );
  NAND2_X1 U17408 ( .A1(n13932), .A2(n13931), .ZN(P2_U3593) );
  NAND2_X1 U17409 ( .A1(n13826), .A2(n13934), .ZN(n13935) );
  NAND2_X1 U17410 ( .A1(n13933), .A2(n13935), .ZN(n16635) );
  INV_X1 U17411 ( .A(n14190), .ZN(n13936) );
  NAND2_X1 U17412 ( .A1(n13936), .A2(n14186), .ZN(n14088) );
  OAI211_X1 U17413 ( .C1(n13936), .C2(n14186), .A(n14088), .B(n16036), .ZN(
        n13938) );
  NAND2_X1 U17414 ( .A1(n9598), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n13937) );
  OAI211_X1 U17415 ( .C1(n16635), .C2(n9598), .A(n13938), .B(n13937), .ZN(
        P2_U2876) );
  INV_X1 U17416 ( .A(n14035), .ZN(n13941) );
  AOI22_X1 U17417 ( .A1(n16921), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n16962), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13939) );
  OAI21_X1 U17418 ( .B1(n14018), .B2(n16929), .A(n13939), .ZN(n13940) );
  AOI21_X1 U17419 ( .B1(n13941), .B2(n16931), .A(n13940), .ZN(n13942) );
  OAI21_X1 U17420 ( .B1(n20293), .B2(n13943), .A(n13942), .ZN(P1_U2997) );
  XOR2_X1 U17421 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n13944), .Z(
        n13988) );
  XNOR2_X1 U17422 ( .A(n13988), .B(n13987), .ZN(n20469) );
  INV_X1 U17423 ( .A(n13945), .ZN(n20378) );
  AOI22_X1 U17424 ( .A1(n16921), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n16962), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n13946) );
  OAI21_X1 U17425 ( .B1(n20374), .B2(n16929), .A(n13946), .ZN(n13947) );
  AOI21_X1 U17426 ( .B1(n20378), .B2(n16931), .A(n13947), .ZN(n13948) );
  OAI21_X1 U17427 ( .B1(n20293), .B2(n20469), .A(n13948), .ZN(P1_U2996) );
  MUX2_X1 U17428 ( .A(n16921), .B(n15241), .S(n13949), .Z(n13950) );
  AOI211_X1 U17429 ( .C1(n13952), .C2(n16926), .A(n13951), .B(n13950), .ZN(
        n13953) );
  OAI21_X1 U17430 ( .B1(n20491), .B2(n14049), .A(n13953), .ZN(P1_U2998) );
  INV_X1 U17431 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n13962) );
  NAND2_X1 U17432 ( .A1(n13954), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14102) );
  NOR2_X1 U17433 ( .A1(n14102), .A2(n14103), .ZN(n14101) );
  INV_X1 U17434 ( .A(n13955), .ZN(n13956) );
  OAI211_X1 U17435 ( .C1(n14101), .C2(n13956), .A(n16036), .B(n13822), .ZN(
        n13961) );
  AND2_X1 U17436 ( .A1(n14100), .A2(n13957), .ZN(n13958) );
  OR2_X1 U17437 ( .A1(n13958), .A2(n13827), .ZN(n16658) );
  INV_X1 U17438 ( .A(n16658), .ZN(n13959) );
  NAND2_X1 U17439 ( .A1(n13959), .A2(n16058), .ZN(n13960) );
  OAI211_X1 U17440 ( .C1(n16058), .C2(n13962), .A(n13961), .B(n13960), .ZN(
        P2_U2878) );
  XNOR2_X1 U17441 ( .A(n14148), .B(n14151), .ZN(n13964) );
  XNOR2_X1 U17442 ( .A(n14149), .B(n13964), .ZN(n13981) );
  AOI22_X1 U17443 ( .A1(n16410), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_REIP_REG_3__SCAN_IN), .B2(n16434), .ZN(n13965) );
  OAI21_X1 U17444 ( .B1(n16413), .B2(n15924), .A(n13965), .ZN(n13966) );
  AOI21_X1 U17445 ( .B1(n15933), .B2(n10023), .A(n13966), .ZN(n13970) );
  NAND3_X1 U17446 ( .A1(n13978), .A2(n16383), .A3(n13968), .ZN(n13969) );
  OAI211_X1 U17447 ( .C1(n13981), .C2(n16439), .A(n13970), .B(n13969), .ZN(
        P2_U3011) );
  NAND2_X1 U17448 ( .A1(n13973), .A2(n13972), .ZN(n13974) );
  NAND2_X1 U17449 ( .A1(n13971), .A2(n13974), .ZN(n15937) );
  INV_X1 U17450 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n20188) );
  OAI22_X1 U17451 ( .A1(n16708), .A2(n15937), .B1(n20188), .B2(n16394), .ZN(
        n13977) );
  INV_X1 U17452 ( .A(n16694), .ZN(n13975) );
  MUX2_X1 U17453 ( .A(n13975), .B(n16693), .S(n14151), .Z(n13976) );
  AOI211_X1 U17454 ( .C1(n16727), .C2(n15933), .A(n13977), .B(n13976), .ZN(
        n13980) );
  NAND3_X1 U17455 ( .A1(n13978), .A2(n12739), .A3(n13968), .ZN(n13979) );
  OAI211_X1 U17456 ( .C1(n13981), .C2(n16721), .A(n13980), .B(n13979), .ZN(
        P2_U3043) );
  INV_X1 U17457 ( .A(n13982), .ZN(n13984) );
  AOI21_X1 U17458 ( .B1(n13985), .B2(n13984), .A(n13983), .ZN(n13994) );
  INV_X1 U17459 ( .A(n13994), .ZN(n20361) );
  XOR2_X1 U17460 ( .A(n16973), .B(n16974), .Z(n20465) );
  AOI22_X1 U17461 ( .A1(n20465), .A2(n20391), .B1(n14968), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n13986) );
  OAI21_X1 U17462 ( .B1(n20361), .B2(n14970), .A(n13986), .ZN(P1_U2868) );
  AOI22_X1 U17463 ( .A1(n13988), .A2(n13987), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13944), .ZN(n13991) );
  XNOR2_X1 U17464 ( .A(n13989), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13990) );
  XNOR2_X1 U17465 ( .A(n13991), .B(n13990), .ZN(n20462) );
  INV_X1 U17466 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21097) );
  NOR2_X1 U17467 ( .A1(n20348), .A2(n21097), .ZN(n20464) );
  AOI21_X1 U17468 ( .B1(n16921), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20464), .ZN(n13992) );
  OAI21_X1 U17469 ( .B1(n20359), .B2(n16929), .A(n13992), .ZN(n13993) );
  AOI21_X1 U17470 ( .B1(n13994), .B2(n16931), .A(n13993), .ZN(n13995) );
  OAI21_X1 U17471 ( .B1(n20462), .B2(n20293), .A(n13995), .ZN(P1_U2995) );
  AND2_X1 U17472 ( .A1(n13998), .A2(n13997), .ZN(n13999) );
  NOR2_X1 U17473 ( .A1(n13996), .A2(n13999), .ZN(n16599) );
  INV_X1 U17474 ( .A(n16599), .ZN(n14001) );
  AOI22_X1 U17475 ( .A1(n14122), .A2(n14624), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19431), .ZN(n14000) );
  OAI21_X1 U17476 ( .B1(n14001), .B2(n14084), .A(n14000), .ZN(P2_U2905) );
  INV_X1 U17477 ( .A(n15005), .ZN(n20521) );
  INV_X1 U17478 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20422) );
  OAI222_X1 U17479 ( .A1(n20361), .A2(n15045), .B1(n15034), .B2(n20521), .C1(
        n20422), .C2(n15031), .ZN(P1_U2900) );
  AND2_X1 U17480 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n10144), .ZN(n14005) );
  NAND2_X1 U17481 ( .A1(n11380), .A2(n14005), .ZN(n14016) );
  INV_X1 U17482 ( .A(n21173), .ZN(n14027) );
  NAND2_X1 U17483 ( .A1(n21173), .A2(n14008), .ZN(n14009) );
  NAND2_X1 U17484 ( .A1(n16908), .A2(n14009), .ZN(n20377) );
  NOR2_X1 U17485 ( .A1(n14027), .A2(n14010), .ZN(n14025) );
  AND2_X1 U17486 ( .A1(n21175), .A2(n20979), .ZN(n16873) );
  INV_X1 U17487 ( .A(n16873), .ZN(n14011) );
  AOI21_X1 U17488 ( .B1(n14013), .B2(n14012), .A(n14011), .ZN(n14023) );
  NOR2_X1 U17489 ( .A1(n20354), .A2(n21162), .ZN(n20366) );
  NOR2_X1 U17490 ( .A1(n20354), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n14045) );
  NAND2_X1 U17491 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21179), .ZN(n16992) );
  OAI21_X1 U17492 ( .B1(n16992), .B2(n10144), .A(n14016), .ZN(n14014) );
  NAND2_X1 U17493 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n20345), .ZN(n14015) );
  OAI22_X1 U17494 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n20366), .B1(n14045), 
        .B2(n14015), .ZN(n14034) );
  INV_X1 U17495 ( .A(n14016), .ZN(n14017) );
  AND2_X2 U17496 ( .A1(n14353), .A2(n14017), .ZN(n20375) );
  INV_X1 U17497 ( .A(n14018), .ZN(n14032) );
  NAND2_X1 U17498 ( .A1(n20508), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14021) );
  NOR2_X1 U17499 ( .A1(n14021), .A2(n16873), .ZN(n14019) );
  NOR2_X1 U17500 ( .A1(n20325), .A2(n14020), .ZN(n14031) );
  INV_X1 U17501 ( .A(n14021), .ZN(n14022) );
  NOR2_X1 U17502 ( .A1(n14023), .A2(n14022), .ZN(n14024) );
  AND2_X2 U17503 ( .A1(n14025), .A2(n14024), .ZN(n20350) );
  INV_X1 U17504 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n14029) );
  NOR2_X1 U17505 ( .A1(n14027), .A2(n14026), .ZN(n20368) );
  INV_X1 U17506 ( .A(n13452), .ZN(n20499) );
  AOI22_X1 U17507 ( .A1(n20368), .A2(n20499), .B1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20369), .ZN(n14028) );
  OAI21_X1 U17508 ( .B1(n20338), .B2(n14029), .A(n14028), .ZN(n14030) );
  AOI211_X1 U17509 ( .C1(n20375), .C2(n14032), .A(n14031), .B(n14030), .ZN(
        n14033) );
  OAI211_X1 U17510 ( .C1(n14035), .C2(n20360), .A(n14034), .B(n14033), .ZN(
        P1_U2838) );
  NOR2_X1 U17511 ( .A1(n13996), .A2(n14037), .ZN(n14038) );
  OR2_X1 U17512 ( .A1(n14036), .A2(n14038), .ZN(n16585) );
  INV_X1 U17513 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19447) );
  INV_X1 U17514 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14039) );
  NOR2_X1 U17515 ( .A1(n14365), .A2(n14039), .ZN(n14040) );
  AOI21_X1 U17516 ( .B1(BUF2_REG_15__SCAN_IN), .B2(n14365), .A(n14040), .ZN(
        n19521) );
  OAI222_X1 U17517 ( .A1(n16585), .A2(n14084), .B1(n16137), .B2(n19447), .C1(
        n19521), .C2(n19441), .ZN(P2_U2904) );
  MUX2_X1 U17518 ( .A(n20375), .B(n20369), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n14047) );
  AND2_X1 U17519 ( .A1(n20367), .A2(n14041), .ZN(n14046) );
  NAND2_X1 U17520 ( .A1(n20350), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n14043) );
  INV_X1 U17521 ( .A(n20345), .ZN(n20326) );
  AOI22_X1 U17522 ( .A1(n20368), .A2(n20981), .B1(n20326), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14042) );
  NAND2_X1 U17523 ( .A1(n14043), .A2(n14042), .ZN(n14044) );
  NOR4_X1 U17524 ( .A1(n14047), .A2(n14046), .A3(n14045), .A4(n14044), .ZN(
        n14048) );
  OAI21_X1 U17525 ( .B1(n20360), .B2(n14049), .A(n14048), .ZN(P1_U2839) );
  NAND2_X1 U17526 ( .A1(n20358), .A2(n20336), .ZN(n14053) );
  AOI22_X1 U17527 ( .A1(n20350), .A2(P1_EBX_REG_0__SCAN_IN), .B1(n20606), .B2(
        n20368), .ZN(n14051) );
  NAND2_X1 U17528 ( .A1(n20354), .A2(n20345), .ZN(n20346) );
  NAND2_X1 U17529 ( .A1(n20346), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n14050) );
  OAI211_X1 U17530 ( .C1(n20325), .C2(n20487), .A(n14051), .B(n14050), .ZN(
        n14052) );
  AOI21_X1 U17531 ( .B1(n14053), .B2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n14052), .ZN(n14054) );
  OAI21_X1 U17532 ( .B1(n20360), .B2(n14055), .A(n14054), .ZN(P1_U2840) );
  INV_X1 U17533 ( .A(n14056), .ZN(n14065) );
  INV_X1 U17534 ( .A(n14057), .ZN(n16787) );
  INV_X1 U17535 ( .A(n16752), .ZN(n16764) );
  NAND2_X1 U17536 ( .A1(n14057), .A2(n20166), .ZN(n16782) );
  OAI21_X1 U17537 ( .B1(n16764), .B2(n14058), .A(n16782), .ZN(n14060) );
  MUX2_X1 U17538 ( .A(n16787), .B(n14060), .S(n14059), .Z(n14064) );
  INV_X1 U17539 ( .A(n14061), .ZN(n14062) );
  AOI211_X1 U17540 ( .C1(n20275), .C2(n16743), .A(n16783), .B(n14062), .ZN(
        n14063) );
  OAI211_X1 U17541 ( .C1(n14065), .C2(n19381), .A(n14064), .B(n14063), .ZN(
        P2_U3176) );
  INV_X1 U17542 ( .A(n14066), .ZN(n14067) );
  NOR2_X1 U17543 ( .A1(n13983), .A2(n14068), .ZN(n14069) );
  NOR2_X1 U17544 ( .A1(n14067), .A2(n14069), .ZN(n20393) );
  INV_X1 U17545 ( .A(n20393), .ZN(n14070) );
  INV_X1 U17546 ( .A(n15001), .ZN(n20525) );
  INV_X1 U17547 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20420) );
  OAI222_X1 U17548 ( .A1(n14070), .A2(n15045), .B1(n15034), .B2(n20525), .C1(
        n15031), .C2(n20420), .ZN(P1_U2899) );
  OR2_X1 U17549 ( .A1(n14072), .A2(n14071), .ZN(n14073) );
  NAND2_X1 U17550 ( .A1(n14074), .A2(n14073), .ZN(n15899) );
  INV_X1 U17551 ( .A(n15937), .ZN(n20259) );
  XOR2_X1 U17552 ( .A(n15937), .B(n19598), .Z(n19427) );
  OAI21_X1 U17553 ( .B1(n16766), .B2(n20268), .A(n14075), .ZN(n19426) );
  NAND2_X1 U17554 ( .A1(n19427), .A2(n19426), .ZN(n19425) );
  OAI21_X1 U17555 ( .B1(n20259), .B2(n10027), .A(n19425), .ZN(n14077) );
  XNOR2_X1 U17556 ( .A(n13971), .B(n14076), .ZN(n15915) );
  NAND2_X1 U17557 ( .A1(n14077), .A2(n15915), .ZN(n14118) );
  INV_X1 U17558 ( .A(n15921), .ZN(n14078) );
  NAND3_X1 U17559 ( .A1(n14118), .A2(n14078), .A3(n19437), .ZN(n14083) );
  INV_X1 U17560 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n14079) );
  OR2_X1 U17561 ( .A1(n14365), .A2(n14079), .ZN(n14081) );
  NAND2_X1 U17562 ( .A1(n14365), .A2(BUF2_REG_5__SCAN_IN), .ZN(n14080) );
  AND2_X1 U17563 ( .A1(n14081), .A2(n14080), .ZN(n19504) );
  INV_X1 U17564 ( .A(n19504), .ZN(n19561) );
  AOI22_X1 U17565 ( .A1(n14122), .A2(n19561), .B1(n19431), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n14082) );
  OAI211_X1 U17566 ( .C1(n14084), .C2(n15899), .A(n14083), .B(n14082), .ZN(
        P2_U2914) );
  NAND2_X1 U17567 ( .A1(n13933), .A2(n14085), .ZN(n14086) );
  NAND2_X1 U17568 ( .A1(n9738), .A2(n14086), .ZN(n16619) );
  INV_X1 U17569 ( .A(n14088), .ZN(n14090) );
  NOR2_X1 U17570 ( .A1(n14088), .A2(n14087), .ZN(n14093) );
  INV_X1 U17571 ( .A(n14093), .ZN(n14089) );
  OAI211_X1 U17572 ( .C1(n14090), .C2(n14184), .A(n14089), .B(n16036), .ZN(
        n14092) );
  NAND2_X1 U17573 ( .A1(n9598), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14091) );
  OAI211_X1 U17574 ( .C1(n16619), .C2(n9598), .A(n14092), .B(n14091), .ZN(
        P2_U2875) );
  NAND2_X1 U17575 ( .A1(n14093), .A2(n14185), .ZN(n14182) );
  OAI211_X1 U17576 ( .C1(n14093), .C2(n14185), .A(n14182), .B(n16036), .ZN(
        n14097) );
  AOI21_X1 U17577 ( .B1(n14095), .B2(n9738), .A(n14094), .ZN(n16605) );
  NAND2_X1 U17578 ( .A1(n16605), .A2(n16058), .ZN(n14096) );
  OAI211_X1 U17579 ( .C1(n16058), .C2(n12446), .A(n14097), .B(n14096), .ZN(
        P2_U2874) );
  NAND2_X1 U17580 ( .A1(n13835), .A2(n14098), .ZN(n14099) );
  NAND2_X1 U17581 ( .A1(n14100), .A2(n14099), .ZN(n16670) );
  NOR2_X1 U17582 ( .A1(n16670), .A2(n9598), .ZN(n14105) );
  AOI211_X1 U17583 ( .C1(n14103), .C2(n14102), .A(n16061), .B(n14101), .ZN(
        n14104) );
  AOI211_X1 U17584 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n9598), .A(n14105), .B(
        n14104), .ZN(n14106) );
  INV_X1 U17585 ( .A(n14106), .ZN(P2_U2879) );
  AND2_X1 U17586 ( .A1(n14107), .A2(n14108), .ZN(n15040) );
  OAI21_X1 U17588 ( .B1(n15040), .B2(n14111), .A(n14110), .ZN(n16909) );
  AND2_X1 U17589 ( .A1(n15506), .A2(n14112), .ZN(n14113) );
  OR2_X1 U17590 ( .A1(n14113), .A2(n14937), .ZN(n16914) );
  OAI22_X1 U17591 ( .A1(n16914), .A2(n14972), .B1(n14114), .B2(n20396), .ZN(
        n14115) );
  INV_X1 U17592 ( .A(n14115), .ZN(n14116) );
  OAI21_X1 U17593 ( .B1(n16909), .B2(n14970), .A(n14116), .ZN(P1_U2862) );
  MUX2_X1 U17594 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n20492), .Z(
        n20432) );
  AOI22_X1 U17595 ( .A1(n15043), .A2(n20432), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15041), .ZN(n14117) );
  OAI21_X1 U17596 ( .B1(n16909), .B2(n15045), .A(n14117), .ZN(P1_U2894) );
  XNOR2_X1 U17597 ( .A(n14118), .B(n15921), .ZN(n14119) );
  NAND2_X1 U17598 ( .A1(n14119), .A2(n19437), .ZN(n14124) );
  INV_X1 U17599 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n17055) );
  OR2_X1 U17600 ( .A1(n14365), .A2(n17055), .ZN(n14121) );
  NAND2_X1 U17601 ( .A1(n14365), .A2(BUF2_REG_4__SCAN_IN), .ZN(n14120) );
  AND2_X1 U17602 ( .A1(n14121), .A2(n14120), .ZN(n19502) );
  INV_X1 U17603 ( .A(n19502), .ZN(n19555) );
  AOI22_X1 U17604 ( .A1(n14122), .A2(n19555), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19431), .ZN(n14123) );
  OAI211_X1 U17605 ( .C1(n15915), .C2(n16165), .A(n14124), .B(n14123), .ZN(
        P2_U2915) );
  XOR2_X1 U17606 ( .A(n14125), .B(n14067), .Z(n20332) );
  INV_X1 U17607 ( .A(n20332), .ZN(n14171) );
  INV_X1 U17608 ( .A(n14997), .ZN(n20528) );
  INV_X1 U17609 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20418) );
  OAI222_X1 U17610 ( .A1(n15045), .A2(n14171), .B1(n15034), .B2(n20528), .C1(
        n15031), .C2(n20418), .ZN(P1_U2898) );
  NAND2_X1 U17611 ( .A1(n14126), .A2(n14127), .ZN(n14129) );
  NAND2_X1 U17612 ( .A1(n14129), .A2(n14128), .ZN(n14167) );
  AND2_X1 U17613 ( .A1(n14107), .A2(n14167), .ZN(n14169) );
  NAND2_X1 U17614 ( .A1(n14126), .A2(n14130), .ZN(n14132) );
  NAND2_X1 U17615 ( .A1(n14132), .A2(n14131), .ZN(n14133) );
  NAND2_X1 U17616 ( .A1(n14133), .A2(n14107), .ZN(n15038) );
  OAI21_X1 U17617 ( .B1(n14169), .B2(n14134), .A(n15038), .ZN(n15250) );
  INV_X1 U17618 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21225) );
  NAND4_X1 U17619 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_3__SCAN_IN), .ZN(n20351)
         );
  NAND2_X1 U17620 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20315) );
  NOR3_X1 U17621 ( .A1(n21225), .A2(n20351), .A3(n20315), .ZN(n14137) );
  INV_X1 U17622 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21103) );
  NAND3_X1 U17623 ( .A1(n20327), .A2(n14137), .A3(n21103), .ZN(n14146) );
  INV_X1 U17624 ( .A(n15252), .ZN(n14144) );
  OAI21_X1 U17625 ( .B1(n9781), .B2(n14135), .A(n15504), .ZN(n16947) );
  NOR2_X1 U17626 ( .A1(n20325), .A2(n16947), .ZN(n14143) );
  INV_X1 U17627 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14141) );
  AOI21_X1 U17628 ( .B1(n20369), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16962), .ZN(n14140) );
  INV_X1 U17629 ( .A(n20346), .ZN(n14822) );
  NAND2_X1 U17630 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14137), .ZN(n14814) );
  INV_X1 U17631 ( .A(n14814), .ZN(n14138) );
  AND2_X1 U17632 ( .A1(n20345), .A2(n14138), .ZN(n14934) );
  NOR2_X1 U17633 ( .A1(n14822), .A2(n14934), .ZN(n20309) );
  NAND2_X1 U17634 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20309), .ZN(n14139) );
  OAI211_X1 U17635 ( .C1(n20338), .C2(n14141), .A(n14140), .B(n14139), .ZN(
        n14142) );
  AOI211_X1 U17636 ( .C1(n20375), .C2(n14144), .A(n14143), .B(n14142), .ZN(
        n14145) );
  OAI211_X1 U17637 ( .C1(n15250), .C2(n16908), .A(n14146), .B(n14145), .ZN(
        P1_U2832) );
  XNOR2_X1 U17638 ( .A(n14147), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14180) );
  INV_X1 U17639 ( .A(n14149), .ZN(n14152) );
  OAI21_X1 U17640 ( .B1(n14149), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n14148), .ZN(n14150) );
  OAI21_X1 U17641 ( .B1(n14152), .B2(n14151), .A(n14150), .ZN(n14154) );
  XNOR2_X1 U17642 ( .A(n15914), .B(n14207), .ZN(n14153) );
  XNOR2_X1 U17643 ( .A(n14154), .B(n14153), .ZN(n14178) );
  AOI22_X1 U17644 ( .A1(n16410), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n16434), .ZN(n14156) );
  NAND2_X1 U17645 ( .A1(n16433), .A2(n15908), .ZN(n14155) );
  OAI211_X1 U17646 ( .C1(n14157), .C2(n16409), .A(n14156), .B(n14155), .ZN(
        n14158) );
  AOI21_X1 U17647 ( .B1(n14178), .B2(n16426), .A(n14158), .ZN(n14159) );
  OAI21_X1 U17648 ( .B1(n14180), .B2(n16429), .A(n14159), .ZN(P2_U3010) );
  XNOR2_X1 U17649 ( .A(n14182), .B(n14181), .ZN(n14164) );
  OR2_X1 U17650 ( .A1(n14094), .A2(n14161), .ZN(n14162) );
  NAND2_X1 U17651 ( .A1(n14160), .A2(n14162), .ZN(n16596) );
  MUX2_X1 U17652 ( .A(n16596), .B(n12448), .S(n9598), .Z(n14163) );
  OAI21_X1 U17653 ( .B1(n14164), .B2(n16061), .A(n14163), .ZN(P2_U2873) );
  MUX2_X1 U17654 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n20492), .Z(
        n20430) );
  INV_X1 U17655 ( .A(n20430), .ZN(n14166) );
  OAI222_X1 U17656 ( .A1(n15250), .A2(n15045), .B1(n15034), .B2(n14166), .C1(
        n14165), .C2(n15031), .ZN(P1_U2896) );
  NOR2_X1 U17657 ( .A1(n14107), .A2(n14167), .ZN(n14168) );
  INV_X1 U17658 ( .A(n20387), .ZN(n14170) );
  INV_X1 U17659 ( .A(n14993), .ZN(n20535) );
  OAI222_X1 U17660 ( .A1(n14170), .A2(n15045), .B1(n15034), .B2(n20535), .C1(
        n15031), .C2(n11088), .ZN(P1_U2897) );
  INV_X1 U17661 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n14172) );
  XNOR2_X1 U17662 ( .A(n16975), .B(n16953), .ZN(n16961) );
  INV_X1 U17663 ( .A(n16961), .ZN(n20324) );
  OAI222_X1 U17664 ( .A1(n14172), .A2(n20396), .B1(n14972), .B2(n20324), .C1(
        n14970), .C2(n14171), .ZN(P1_U2866) );
  NOR2_X1 U17665 ( .A1(n15915), .A2(n16708), .ZN(n14177) );
  INV_X1 U17666 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n20190) );
  NAND2_X1 U17667 ( .A1(n15918), .A2(n16727), .ZN(n14175) );
  NAND2_X1 U17668 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16693), .ZN(
        n14206) );
  OAI21_X1 U17669 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16729), .A(
        n16694), .ZN(n14211) );
  INV_X1 U17670 ( .A(n14211), .ZN(n14173) );
  MUX2_X1 U17671 ( .A(n14206), .B(n14173), .S(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n14174) );
  OAI211_X1 U17672 ( .C1(n20190), .C2(n16394), .A(n14175), .B(n14174), .ZN(
        n14176) );
  AOI211_X1 U17673 ( .C1(n14178), .C2(n16689), .A(n14177), .B(n14176), .ZN(
        n14179) );
  OAI21_X1 U17674 ( .B1(n14180), .B2(n16706), .A(n14179), .ZN(P2_U3042) );
  OAI222_X1 U17675 ( .A1(n16947), .A2(n14972), .B1(n20396), .B2(n14141), .C1(
        n14970), .C2(n15250), .ZN(P1_U2864) );
  INV_X1 U17676 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n14198) );
  OAI21_X1 U17677 ( .B1(n14182), .B2(n14181), .A(n14183), .ZN(n14192) );
  INV_X1 U17678 ( .A(n14183), .ZN(n14189) );
  AND2_X1 U17679 ( .A1(n14185), .A2(n14184), .ZN(n14188) );
  INV_X1 U17680 ( .A(n14380), .ZN(n14191) );
  NAND3_X1 U17681 ( .A1(n14192), .A2(n16036), .A3(n14191), .ZN(n14197) );
  NAND2_X1 U17682 ( .A1(n14160), .A2(n14194), .ZN(n14195) );
  NAND2_X1 U17683 ( .A1(n16583), .A2(n16058), .ZN(n14196) );
  OAI211_X1 U17684 ( .C1(n16058), .C2(n14198), .A(n14197), .B(n14196), .ZN(
        P2_U2872) );
  OAI21_X1 U17685 ( .B1(n14202), .B2(n14200), .A(n14199), .ZN(n14201) );
  OAI21_X1 U17686 ( .B1(n14203), .B2(n14202), .A(n14201), .ZN(n14221) );
  XOR2_X1 U17687 ( .A(n14204), .B(n14205), .Z(n14219) );
  NOR2_X1 U17688 ( .A1(n15894), .A2(n16669), .ZN(n14214) );
  AOI221_X1 U17689 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n14208), .C2(n14207), .A(
        n14206), .ZN(n14210) );
  NOR2_X1 U17690 ( .A1(n16394), .A2(n12040), .ZN(n14209) );
  AOI211_X1 U17691 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n14211), .A(
        n14210), .B(n14209), .ZN(n14212) );
  OAI21_X1 U17692 ( .B1(n15899), .B2(n16708), .A(n14212), .ZN(n14213) );
  AOI211_X1 U17693 ( .C1(n14219), .C2(n16689), .A(n14214), .B(n14213), .ZN(
        n14215) );
  OAI21_X1 U17694 ( .B1(n14221), .B2(n16706), .A(n14215), .ZN(P2_U3041) );
  NOR2_X1 U17695 ( .A1(n15894), .A2(n16409), .ZN(n14218) );
  AOI22_X1 U17696 ( .A1(n16410), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        P2_REIP_REG_5__SCAN_IN), .B2(n16434), .ZN(n14216) );
  OAI21_X1 U17697 ( .B1(n16413), .B2(n15893), .A(n14216), .ZN(n14217) );
  AOI211_X1 U17698 ( .C1(n14219), .C2(n16426), .A(n14218), .B(n14217), .ZN(
        n14220) );
  OAI21_X1 U17699 ( .B1(n14221), .B2(n16429), .A(n14220), .ZN(P2_U3009) );
  AND2_X1 U17700 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n14239) );
  INV_X1 U17701 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n17535) );
  INV_X1 U17702 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17201) );
  NOR4_X1 U17703 ( .A1(n17171), .A2(n17535), .A3(n17201), .A4(n17576), .ZN(
        n14222) );
  NAND4_X1 U17704 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(n14239), .A4(n14222), .ZN(n17523) );
  INV_X1 U17705 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17321) );
  NAND4_X1 U17706 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .A4(P3_EBX_REG_2__SCAN_IN), .ZN(n17761) );
  INV_X1 U17707 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n17426) );
  NOR2_X1 U17708 ( .A1(n17761), .A2(n17426), .ZN(n14225) );
  NAND2_X1 U17709 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17757), .ZN(n17756) );
  NAND2_X1 U17710 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17713), .ZN(n17671) );
  NAND2_X1 U17711 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .ZN(n17617) );
  NAND2_X1 U17712 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17604), .ZN(n17561) );
  NOR3_X1 U17713 ( .A1(n17515), .A2(n17523), .A3(n17561), .ZN(n17512) );
  NAND2_X1 U17714 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17512), .ZN(n14226) );
  NOR2_X1 U17715 ( .A1(n17826), .A2(n14226), .ZN(n14228) );
  NAND2_X1 U17716 ( .A1(n17775), .A2(n14226), .ZN(n17513) );
  INV_X1 U17717 ( .A(n17513), .ZN(n14227) );
  MUX2_X1 U17718 ( .A(n14228), .B(n14227), .S(P3_EBX_REG_31__SCAN_IN), .Z(
        P3_U2672) );
  INV_X1 U17719 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19203) );
  OAI21_X1 U17720 ( .B1(n14229), .B2(n12710), .A(n19203), .ZN(n16806) );
  NAND2_X1 U17721 ( .A1(n14230), .A2(n16806), .ZN(n19158) );
  NOR2_X1 U17722 ( .A1(n19370), .A2(n19158), .ZN(n14238) );
  NAND2_X1 U17723 ( .A1(n19153), .A2(n19361), .ZN(n14236) );
  NAND3_X1 U17724 ( .A1(n19228), .A2(n14232), .A3(n14231), .ZN(n17933) );
  AOI211_X1 U17725 ( .C1(n14234), .C2(n9744), .A(n16898), .B(n14233), .ZN(
        n14235) );
  OAI21_X1 U17726 ( .B1(n14236), .B2(n17933), .A(n14235), .ZN(n19181) );
  INV_X1 U17727 ( .A(n19181), .ZN(n19191) );
  NAND2_X1 U17728 ( .A1(n19215), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18720) );
  NAND3_X1 U17729 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19311)
         );
  INV_X1 U17730 ( .A(n19311), .ZN(n19220) );
  NAND2_X1 U17731 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n19220), .ZN(n14237) );
  OAI211_X1 U17732 ( .C1(n19212), .C2(n19191), .A(n18720), .B(n14237), .ZN(
        n19332) );
  MUX2_X1 U17733 ( .A(n14238), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19340), .Z(P3_U3284) );
  NAND2_X1 U17734 ( .A1(n12696), .A2(n17779), .ZN(n17782) );
  NAND2_X1 U17735 ( .A1(n17604), .A2(n12696), .ZN(n17589) );
  INV_X1 U17736 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17590) );
  NAND2_X1 U17737 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17538), .ZN(n17529) );
  NAND2_X1 U17738 ( .A1(n17775), .A2(n17529), .ZN(n17527) );
  OAI21_X1 U17739 ( .B1(n14239), .B2(n17782), .A(n17527), .ZN(n17520) );
  AOI22_X1 U17740 ( .A1(n17684), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9610), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14243) );
  AOI22_X1 U17741 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14242) );
  AOI22_X1 U17742 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17738), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14241) );
  AOI22_X1 U17743 ( .A1(n9628), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14240) );
  NAND4_X1 U17744 ( .A1(n14243), .A2(n14242), .A3(n14241), .A4(n14240), .ZN(
        n14249) );
  AOI22_X1 U17745 ( .A1(n12813), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14247) );
  AOI22_X1 U17746 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17734), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14246) );
  AOI22_X1 U17747 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14305), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14245) );
  AOI22_X1 U17748 ( .A1(n17720), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14244) );
  NAND4_X1 U17749 ( .A1(n14247), .A2(n14246), .A3(n14245), .A4(n14244), .ZN(
        n14248) );
  NOR2_X1 U17750 ( .A1(n14249), .A2(n14248), .ZN(n17525) );
  AOI22_X1 U17751 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17721), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14253) );
  AOI22_X1 U17752 ( .A1(n17684), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14252) );
  AOI22_X1 U17753 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14251) );
  AOI22_X1 U17754 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14250) );
  NAND4_X1 U17755 ( .A1(n14253), .A2(n14252), .A3(n14251), .A4(n14250), .ZN(
        n14259) );
  AOI22_X1 U17756 ( .A1(n17734), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14257) );
  AOI22_X1 U17757 ( .A1(n17714), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16791), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14256) );
  AOI22_X1 U17758 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12813), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14255) );
  AOI22_X1 U17759 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14254) );
  NAND4_X1 U17760 ( .A1(n14257), .A2(n14256), .A3(n14255), .A4(n14254), .ZN(
        n14258) );
  NOR2_X1 U17761 ( .A1(n14259), .A2(n14258), .ZN(n17536) );
  AOI22_X1 U17762 ( .A1(n17720), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14263) );
  AOI22_X1 U17763 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14262) );
  AOI22_X1 U17764 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17738), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14261) );
  AOI22_X1 U17765 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14260) );
  NAND4_X1 U17766 ( .A1(n14263), .A2(n14262), .A3(n14261), .A4(n14260), .ZN(
        n14269) );
  AOI22_X1 U17767 ( .A1(n12842), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17684), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14267) );
  AOI22_X1 U17768 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14266) );
  AOI22_X1 U17769 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14265) );
  AOI22_X1 U17770 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12836), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14264) );
  NAND4_X1 U17771 ( .A1(n14267), .A2(n14266), .A3(n14265), .A4(n14264), .ZN(
        n14268) );
  NOR2_X1 U17772 ( .A1(n14269), .A2(n14268), .ZN(n17546) );
  AOI22_X1 U17773 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17643), .B1(
        n14270), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14274) );
  AOI22_X1 U17774 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17701), .ZN(n14273) );
  AOI22_X1 U17775 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17684), .B1(
        n17738), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14272) );
  AOI22_X1 U17776 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n9628), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17719), .ZN(n14271) );
  NAND4_X1 U17777 ( .A1(n14274), .A2(n14273), .A3(n14272), .A4(n14271), .ZN(
        n14280) );
  AOI22_X1 U17778 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n17733), .ZN(n14278) );
  AOI22_X1 U17779 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n9591), .ZN(n14277) );
  AOI22_X1 U17780 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17720), .B1(
        n17734), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14276) );
  AOI22_X1 U17781 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17676), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14275) );
  NAND4_X1 U17782 ( .A1(n14278), .A2(n14277), .A3(n14276), .A4(n14275), .ZN(
        n14279) );
  NOR2_X1 U17783 ( .A1(n14280), .A2(n14279), .ZN(n17545) );
  NOR2_X1 U17784 ( .A1(n17546), .A2(n17545), .ZN(n17542) );
  AOI22_X1 U17785 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9597), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14290) );
  AOI22_X1 U17786 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14289) );
  AOI22_X1 U17787 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n16791), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14281) );
  OAI21_X1 U17788 ( .B1(n17736), .B2(n21308), .A(n14281), .ZN(n14287) );
  AOI22_X1 U17789 ( .A1(n12842), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14285) );
  AOI22_X1 U17790 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17734), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14284) );
  AOI22_X1 U17791 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17738), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14283) );
  AOI22_X1 U17792 ( .A1(n12813), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14282) );
  NAND4_X1 U17793 ( .A1(n14285), .A2(n14284), .A3(n14283), .A4(n14282), .ZN(
        n14286) );
  AOI211_X1 U17794 ( .C1(n9611), .C2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n14287), .B(n14286), .ZN(n14288) );
  NAND3_X1 U17795 ( .A1(n14290), .A2(n14289), .A3(n14288), .ZN(n17541) );
  NAND2_X1 U17796 ( .A1(n17542), .A2(n17541), .ZN(n17540) );
  NOR2_X1 U17797 ( .A1(n17536), .A2(n17540), .ZN(n17532) );
  AOI22_X1 U17798 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14305), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14300) );
  AOI22_X1 U17799 ( .A1(n12842), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12836), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14299) );
  AOI22_X1 U17800 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(n9591), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14291) );
  OAI21_X1 U17801 ( .B1(n12627), .B2(n21222), .A(n14291), .ZN(n14297) );
  AOI22_X1 U17802 ( .A1(n12813), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14295) );
  AOI22_X1 U17803 ( .A1(n17684), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16791), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14294) );
  AOI22_X1 U17804 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14293) );
  AOI22_X1 U17805 ( .A1(n17738), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14292) );
  NAND4_X1 U17806 ( .A1(n14295), .A2(n14294), .A3(n14293), .A4(n14292), .ZN(
        n14296) );
  AOI211_X1 U17807 ( .C1(n9597), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n14297), .B(n14296), .ZN(n14298) );
  NAND3_X1 U17808 ( .A1(n14300), .A2(n14299), .A3(n14298), .ZN(n17531) );
  NAND2_X1 U17809 ( .A1(n17532), .A2(n17531), .ZN(n17530) );
  NOR2_X1 U17810 ( .A1(n17525), .A2(n17530), .ZN(n17524) );
  AOI22_X1 U17811 ( .A1(n17738), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14304) );
  AOI22_X1 U17812 ( .A1(n17643), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16791), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14303) );
  AOI22_X1 U17813 ( .A1(n12813), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14302) );
  AOI22_X1 U17814 ( .A1(n12842), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14301) );
  NAND4_X1 U17815 ( .A1(n14304), .A2(n14303), .A3(n14302), .A4(n14301), .ZN(
        n14311) );
  AOI22_X1 U17816 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9597), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14309) );
  AOI22_X1 U17817 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14308) );
  AOI22_X1 U17818 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17734), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14307) );
  AOI22_X1 U17819 ( .A1(n17684), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14305), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14306) );
  NAND4_X1 U17820 ( .A1(n14309), .A2(n14308), .A3(n14307), .A4(n14306), .ZN(
        n14310) );
  NOR2_X1 U17821 ( .A1(n14311), .A2(n14310), .ZN(n17516) );
  XNOR2_X1 U17822 ( .A(n17524), .B(n17516), .ZN(n17798) );
  AOI22_X1 U17823 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17520), .B1(n17760), 
        .B2(n17798), .ZN(n14314) );
  INV_X1 U17824 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14312) );
  INV_X1 U17825 ( .A(n17529), .ZN(n17534) );
  NAND3_X1 U17826 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14312), .A3(n17534), 
        .ZN(n14313) );
  NAND2_X1 U17827 ( .A1(n14314), .A2(n14313), .ZN(P3_U2675) );
  NOR2_X1 U17828 ( .A1(n12739), .A2(n14315), .ZN(n14322) );
  INV_X1 U17829 ( .A(n14316), .ZN(n14317) );
  INV_X1 U17830 ( .A(n16729), .ZN(n16716) );
  AOI21_X1 U17831 ( .B1(n14317), .B2(n16716), .A(n16660), .ZN(n16578) );
  INV_X1 U17832 ( .A(n16578), .ZN(n14320) );
  NOR2_X1 U17833 ( .A1(n14318), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14319) );
  OAI21_X1 U17834 ( .B1(n14323), .B2(n14322), .A(n14321), .ZN(n16567) );
  INV_X1 U17835 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16576) );
  AND2_X1 U17836 ( .A1(n16716), .A2(n16576), .ZN(n14324) );
  INV_X1 U17837 ( .A(n14325), .ZN(n14326) );
  NOR2_X1 U17838 ( .A1(n16246), .A2(n14326), .ZN(n16247) );
  INV_X1 U17839 ( .A(n16340), .ZN(n14329) );
  XOR2_X1 U17840 ( .A(n16247), .B(n16248), .Z(n16304) );
  OR2_X1 U17841 ( .A1(n9673), .A2(n14332), .ZN(n14333) );
  NAND2_X1 U17842 ( .A1(n14331), .A2(n14333), .ZN(n16299) );
  OR2_X1 U17843 ( .A1(n14334), .A2(n14336), .ZN(n15745) );
  INV_X1 U17844 ( .A(n15745), .ZN(n14335) );
  AOI21_X1 U17845 ( .B1(n14336), .B2(n14334), .A(n14335), .ZN(n16158) );
  NAND2_X1 U17846 ( .A1(n16158), .A2(n16724), .ZN(n14337) );
  NAND2_X1 U17847 ( .A1(n16434), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n16294) );
  OAI211_X1 U17848 ( .C1(n16669), .C2(n16299), .A(n14337), .B(n16294), .ZN(
        n14338) );
  AOI21_X1 U17849 ( .B1(n16304), .B2(n16689), .A(n14338), .ZN(n14340) );
  INV_X1 U17850 ( .A(n16591), .ZN(n16593) );
  NAND3_X1 U17851 ( .A1(n16616), .A2(n16593), .A3(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16580) );
  OAI211_X1 U17852 ( .C1(n14341), .C2(n16301), .A(n14340), .B(n14339), .ZN(
        P2_U3029) );
  NAND2_X1 U17853 ( .A1(n14342), .A2(n16433), .ZN(n14345) );
  AOI21_X1 U17854 ( .B1(n16410), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14343), .ZN(n14344) );
  NAND2_X1 U17855 ( .A1(n14650), .A2(n16931), .ZN(n14356) );
  INV_X1 U17856 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n14665) );
  NOR2_X1 U17857 ( .A1(n20348), .A2(n14665), .ZN(n15281) );
  NOR2_X1 U17858 ( .A1(n14353), .A2(n16929), .ZN(n14354) );
  AOI211_X1 U17859 ( .C1(n16921), .C2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15281), .B(n14354), .ZN(n14355) );
  OAI211_X1 U17860 ( .C1(n15286), .C2(n20293), .A(n14356), .B(n14355), .ZN(
        P1_U2968) );
  INV_X1 U17861 ( .A(n14357), .ZN(n15976) );
  INV_X1 U17862 ( .A(n19402), .ZN(n15968) );
  INV_X1 U17863 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n14359) );
  OAI22_X1 U17864 ( .A1(n15968), .A2(n14359), .B1(n10065), .B2(n14358), .ZN(
        n14362) );
  NOR2_X1 U17865 ( .A1(n14360), .A2(n16838), .ZN(n14361) );
  AOI211_X1 U17866 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n15963), .A(
        n14362), .B(n14361), .ZN(n14363) );
  NOR2_X2 U17867 ( .A1(n14366), .A2(n14365), .ZN(n16162) );
  AOI22_X1 U17868 ( .A1(n16162), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19431), .ZN(n14368) );
  NOR2_X2 U17869 ( .A1(n14366), .A2(n16771), .ZN(n16168) );
  NAND2_X1 U17870 ( .A1(n16168), .A2(BUF2_REG_31__SCAN_IN), .ZN(n14367) );
  OAI211_X1 U17871 ( .C1(n14369), .C2(n16165), .A(n14368), .B(n14367), .ZN(
        P2_U2888) );
  AOI22_X1 U17872 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14373) );
  AOI22_X1 U17873 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n14462), .B1(
        n14463), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14372) );
  AOI22_X1 U17874 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14371) );
  AOI22_X1 U17875 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14370) );
  NAND4_X1 U17876 ( .A1(n14373), .A2(n14372), .A3(n14371), .A4(n14370), .ZN(
        n14379) );
  AOI22_X1 U17877 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__0__SCAN_IN), .B2(n14470), .ZN(n14377) );
  AOI22_X1 U17878 ( .A1(n11662), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14376) );
  AOI22_X1 U17879 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14375) );
  AOI22_X1 U17880 ( .A1(n14475), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14474), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14374) );
  NAND4_X1 U17881 ( .A1(n14377), .A2(n14376), .A3(n14375), .A4(n14374), .ZN(
        n14378) );
  OR2_X1 U17882 ( .A1(n14379), .A2(n14378), .ZN(n16057) );
  NAND2_X1 U17883 ( .A1(n14380), .A2(n16057), .ZN(n16056) );
  AOI22_X1 U17884 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n14461), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14384) );
  AOI22_X1 U17885 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n14463), .B1(
        n14462), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14383) );
  AOI22_X1 U17886 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14382) );
  AOI22_X1 U17887 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14381) );
  NAND4_X1 U17888 ( .A1(n14384), .A2(n14383), .A3(n14382), .A4(n14381), .ZN(
        n14390) );
  AOI22_X1 U17889 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n14470), .ZN(n14388) );
  AOI22_X1 U17890 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11662), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14387) );
  AOI22_X1 U17891 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14386) );
  AOI22_X1 U17892 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n14475), .B1(
        n14474), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14385) );
  NAND4_X1 U17893 ( .A1(n14388), .A2(n14387), .A3(n14386), .A4(n14385), .ZN(
        n14389) );
  AOI22_X1 U17894 ( .A1(n12122), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14394) );
  AOI22_X1 U17895 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n14463), .B1(
        n14462), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14393) );
  AOI22_X1 U17896 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14392) );
  AOI22_X1 U17897 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14391) );
  NAND4_X1 U17898 ( .A1(n14394), .A2(n14393), .A3(n14392), .A4(n14391), .ZN(
        n14400) );
  AOI22_X1 U17899 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__2__SCAN_IN), .B2(n14470), .ZN(n14398) );
  AOI22_X1 U17900 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11662), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14397) );
  AOI22_X1 U17901 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14396) );
  AOI22_X1 U17902 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n14475), .B1(
        n14474), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14395) );
  NAND4_X1 U17903 ( .A1(n14398), .A2(n14397), .A3(n14396), .A4(n14395), .ZN(
        n14399) );
  NOR2_X1 U17904 ( .A1(n14400), .A2(n14399), .ZN(n16049) );
  AOI22_X1 U17905 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14404) );
  AOI22_X1 U17906 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n14463), .B1(
        n14462), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14403) );
  AOI22_X1 U17907 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14402) );
  AOI22_X1 U17908 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14401) );
  NAND4_X1 U17909 ( .A1(n14404), .A2(n14403), .A3(n14402), .A4(n14401), .ZN(
        n14410) );
  AOI22_X1 U17910 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__3__SCAN_IN), .B2(n14470), .ZN(n14408) );
  AOI22_X1 U17911 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11662), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14407) );
  AOI22_X1 U17912 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14406) );
  AOI22_X1 U17913 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n14475), .B1(
        n14474), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14405) );
  NAND4_X1 U17914 ( .A1(n14408), .A2(n14407), .A3(n14406), .A4(n14405), .ZN(
        n14409) );
  AOI22_X1 U17915 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14414) );
  AOI22_X1 U17916 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n14463), .B1(
        n14462), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14413) );
  AOI22_X1 U17917 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14412) );
  AOI22_X1 U17918 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14411) );
  NAND4_X1 U17919 ( .A1(n14414), .A2(n14413), .A3(n14412), .A4(n14411), .ZN(
        n14420) );
  AOI22_X1 U17920 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(n14470), .ZN(n14418) );
  AOI22_X1 U17921 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11662), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14417) );
  AOI22_X1 U17922 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14416) );
  AOI22_X1 U17923 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n14475), .B1(
        n14474), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14415) );
  NAND4_X1 U17924 ( .A1(n14418), .A2(n14417), .A3(n14416), .A4(n14415), .ZN(
        n14419) );
  OR2_X1 U17925 ( .A1(n14420), .A2(n14419), .ZN(n16040) );
  NAND2_X1 U17926 ( .A1(n16039), .A2(n16040), .ZN(n16033) );
  AOI22_X1 U17927 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14424) );
  AOI22_X1 U17928 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n14463), .B1(
        n11942), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14423) );
  AOI22_X1 U17929 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14422) );
  AOI22_X1 U17930 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14421) );
  NAND4_X1 U17931 ( .A1(n14424), .A2(n14423), .A3(n14422), .A4(n14421), .ZN(
        n14430) );
  AOI22_X1 U17932 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__5__SCAN_IN), .B2(n14470), .ZN(n14428) );
  AOI22_X1 U17933 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n11662), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14427) );
  AOI22_X1 U17934 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14426) );
  AOI22_X1 U17935 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n14475), .B1(
        n14474), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14425) );
  NAND4_X1 U17936 ( .A1(n14428), .A2(n14427), .A3(n14426), .A4(n14425), .ZN(
        n14429) );
  NOR2_X1 U17937 ( .A1(n14430), .A2(n14429), .ZN(n16035) );
  INV_X1 U17938 ( .A(n16035), .ZN(n14431) );
  AOI22_X1 U17939 ( .A1(n12122), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14435) );
  AOI22_X1 U17940 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n14463), .B1(
        n14462), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14434) );
  AOI22_X1 U17941 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14433) );
  AOI22_X1 U17942 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14432) );
  NAND4_X1 U17943 ( .A1(n14435), .A2(n14434), .A3(n14433), .A4(n14432), .ZN(
        n14442) );
  AOI22_X1 U17944 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n14470), .ZN(n14440) );
  AOI22_X1 U17945 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11662), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14439) );
  AOI22_X1 U17946 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14438) );
  AOI22_X1 U17947 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n14475), .B1(
        n14474), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14437) );
  NAND4_X1 U17948 ( .A1(n14440), .A2(n14439), .A3(n14438), .A4(n14437), .ZN(
        n14441) );
  NOR2_X1 U17949 ( .A1(n14442), .A2(n14441), .ZN(n16028) );
  AOI22_X1 U17950 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14605), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14451) );
  NAND2_X1 U17951 ( .A1(n14509), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n14446) );
  AND2_X1 U17952 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14444) );
  OR2_X1 U17953 ( .A1(n14444), .A2(n14443), .ZN(n14612) );
  NAND2_X1 U17954 ( .A1(n14611), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n14445) );
  AND3_X1 U17955 ( .A1(n14446), .A2(n14612), .A3(n14445), .ZN(n14450) );
  AOI22_X1 U17956 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14598), .B1(
        n14606), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14448) );
  NAND4_X1 U17957 ( .A1(n14451), .A2(n14450), .A3(n14449), .A4(n14448), .ZN(
        n14460) );
  AOI22_X1 U17958 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14605), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14458) );
  NAND2_X1 U17959 ( .A1(n14509), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n14453) );
  INV_X1 U17960 ( .A(n14612), .ZN(n14577) );
  NAND2_X1 U17961 ( .A1(n14611), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n14452) );
  AND3_X1 U17962 ( .A1(n14453), .A2(n14577), .A3(n14452), .ZN(n14457) );
  AOI22_X1 U17963 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14606), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14455) );
  NAND4_X1 U17964 ( .A1(n14458), .A2(n14457), .A3(n14456), .A4(n14455), .ZN(
        n14459) );
  NAND2_X1 U17965 ( .A1(n14460), .A2(n14459), .ZN(n14500) );
  AOI22_X1 U17966 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11941), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14469) );
  AOI22_X1 U17967 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n14463), .B1(
        n14462), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14468) );
  AOI22_X1 U17968 ( .A1(n14464), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11612), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14467) );
  AOI22_X1 U17969 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14465), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14466) );
  NAND4_X1 U17970 ( .A1(n14469), .A2(n14468), .A3(n14467), .A4(n14466), .ZN(
        n14481) );
  AOI22_X1 U17971 ( .A1(n11661), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n14470), .ZN(n14479) );
  AOI22_X1 U17972 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11662), .B1(
        n14471), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14478) );
  AOI22_X1 U17973 ( .A1(n14473), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14472), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14477) );
  AOI22_X1 U17974 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n14475), .B1(
        n14474), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14476) );
  NAND4_X1 U17975 ( .A1(n14479), .A2(n14478), .A3(n14477), .A4(n14476), .ZN(
        n14480) );
  AOI22_X1 U17976 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14605), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14487) );
  NAND2_X1 U17977 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n14483) );
  NAND2_X1 U17978 ( .A1(n14611), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n14482) );
  AND3_X1 U17979 ( .A1(n14483), .A2(n14612), .A3(n14482), .ZN(n14486) );
  AOI22_X1 U17980 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14606), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14484) );
  NAND4_X1 U17981 ( .A1(n14487), .A2(n14486), .A3(n14485), .A4(n14484), .ZN(
        n14495) );
  AOI22_X1 U17982 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14605), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14493) );
  NAND2_X1 U17983 ( .A1(n9603), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n14489) );
  NAND2_X1 U17984 ( .A1(n14611), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14488) );
  AND3_X1 U17985 ( .A1(n14489), .A2(n14577), .A3(n14488), .ZN(n14492) );
  AOI22_X1 U17986 ( .A1(n14610), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14606), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14490) );
  NAND4_X1 U17987 ( .A1(n14493), .A2(n14492), .A3(n14491), .A4(n14490), .ZN(
        n14494) );
  NAND2_X1 U17988 ( .A1(n14497), .A2(n16007), .ZN(n14496) );
  INV_X1 U17989 ( .A(n14556), .ZN(n14539) );
  NOR2_X1 U17990 ( .A1(n14496), .A2(n14500), .ZN(n14518) );
  AOI211_X1 U17991 ( .C1(n14500), .C2(n14496), .A(n14539), .B(n14518), .ZN(
        n16011) );
  NAND2_X1 U17992 ( .A1(n14561), .A2(n16007), .ZN(n14498) );
  XNOR2_X1 U17993 ( .A(n14498), .B(n14497), .ZN(n16009) );
  NOR2_X1 U17994 ( .A1(n14561), .A2(n14500), .ZN(n16010) );
  NAND3_X1 U17995 ( .A1(n16009), .A2(n16007), .A3(n16010), .ZN(n14501) );
  AOI22_X1 U17996 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14605), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14508) );
  NAND2_X1 U17997 ( .A1(n14509), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n14504) );
  NAND2_X1 U17998 ( .A1(n14611), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n14503) );
  AND3_X1 U17999 ( .A1(n14504), .A2(n14612), .A3(n14503), .ZN(n14507) );
  AOI22_X1 U18000 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14606), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14505) );
  NAND4_X1 U18001 ( .A1(n14508), .A2(n14507), .A3(n14506), .A4(n14505), .ZN(
        n14517) );
  AOI22_X1 U18002 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14605), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14515) );
  NAND2_X1 U18003 ( .A1(n14509), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n14511) );
  NAND2_X1 U18004 ( .A1(n14611), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14510) );
  AND3_X1 U18005 ( .A1(n14511), .A2(n14577), .A3(n14510), .ZN(n14514) );
  AOI22_X1 U18006 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14606), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14512) );
  NAND4_X1 U18007 ( .A1(n14515), .A2(n14514), .A3(n14513), .A4(n14512), .ZN(
        n14516) );
  AND2_X1 U18008 ( .A1(n14517), .A2(n14516), .ZN(n14520) );
  NAND2_X1 U18009 ( .A1(n14518), .A2(n14520), .ZN(n14540) );
  OAI211_X1 U18010 ( .C1(n14518), .C2(n14520), .A(n14556), .B(n14540), .ZN(
        n14537) );
  INV_X1 U18011 ( .A(n14537), .ZN(n14519) );
  NAND2_X1 U18012 ( .A1(n10064), .A2(n14520), .ZN(n16002) );
  INV_X1 U18013 ( .A(n16002), .ZN(n14536) );
  AOI22_X1 U18014 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14605), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14526) );
  NAND2_X1 U18015 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n14522) );
  NAND2_X1 U18016 ( .A1(n14611), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n14521) );
  AND3_X1 U18017 ( .A1(n14522), .A2(n14612), .A3(n14521), .ZN(n14525) );
  AOI22_X1 U18018 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14606), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14523) );
  NAND4_X1 U18019 ( .A1(n14526), .A2(n14525), .A3(n14524), .A4(n14523), .ZN(
        n14534) );
  AOI22_X1 U18020 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14605), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14532) );
  NAND2_X1 U18021 ( .A1(n9603), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n14528) );
  NAND2_X1 U18022 ( .A1(n14611), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14527) );
  AND3_X1 U18023 ( .A1(n14528), .A2(n14577), .A3(n14527), .ZN(n14531) );
  AOI22_X1 U18024 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14606), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14529) );
  NAND4_X1 U18025 ( .A1(n14532), .A2(n14531), .A3(n14530), .A4(n14529), .ZN(
        n14533) );
  NAND2_X1 U18026 ( .A1(n14534), .A2(n14533), .ZN(n15994) );
  INV_X1 U18027 ( .A(n14540), .ZN(n14538) );
  AND2_X1 U18028 ( .A1(n14538), .A2(n14535), .ZN(n14558) );
  AOI211_X1 U18029 ( .C1(n15994), .C2(n14540), .A(n14539), .B(n14558), .ZN(
        n15996) );
  AOI22_X1 U18030 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14605), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14546) );
  NAND2_X1 U18031 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n14542) );
  NAND2_X1 U18032 ( .A1(n14611), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n14541) );
  AND3_X1 U18033 ( .A1(n14542), .A2(n14612), .A3(n14541), .ZN(n14545) );
  AOI22_X1 U18034 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14606), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14543) );
  NAND4_X1 U18035 ( .A1(n14546), .A2(n14545), .A3(n14544), .A4(n14543), .ZN(
        n14554) );
  AOI22_X1 U18036 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14605), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14552) );
  NAND2_X1 U18037 ( .A1(n9603), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n14548) );
  NAND2_X1 U18038 ( .A1(n14611), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14547) );
  AND3_X1 U18039 ( .A1(n14548), .A2(n14577), .A3(n14547), .ZN(n14551) );
  AOI22_X1 U18040 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14606), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14549) );
  NAND4_X1 U18041 ( .A1(n14552), .A2(n14551), .A3(n14550), .A4(n14549), .ZN(
        n14553) );
  NAND2_X1 U18042 ( .A1(n14554), .A2(n14553), .ZN(n14560) );
  INV_X1 U18043 ( .A(n14560), .ZN(n14557) );
  INV_X1 U18044 ( .A(n14558), .ZN(n14555) );
  OAI211_X1 U18045 ( .C1(n14558), .C2(n14557), .A(n14556), .B(n14591), .ZN(
        n14559) );
  NOR2_X1 U18046 ( .A1(n14561), .A2(n14560), .ZN(n15988) );
  AOI22_X1 U18047 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14605), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14567) );
  NAND2_X1 U18048 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n14563) );
  NAND2_X1 U18049 ( .A1(n14611), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n14562) );
  AND3_X1 U18050 ( .A1(n14563), .A2(n14612), .A3(n14562), .ZN(n14566) );
  AOI22_X1 U18051 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14606), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14564) );
  NAND4_X1 U18052 ( .A1(n14567), .A2(n14566), .A3(n14565), .A4(n14564), .ZN(
        n14575) );
  AOI22_X1 U18053 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14605), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14573) );
  NAND2_X1 U18054 ( .A1(n9604), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n14569) );
  NAND2_X1 U18055 ( .A1(n14611), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n14568) );
  AND3_X1 U18056 ( .A1(n14569), .A2(n14577), .A3(n14568), .ZN(n14572) );
  AOI22_X1 U18057 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14606), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14570) );
  NAND4_X1 U18058 ( .A1(n14573), .A2(n14572), .A3(n14571), .A4(n14570), .ZN(
        n14574) );
  NAND2_X1 U18059 ( .A1(n14575), .A2(n14574), .ZN(n15983) );
  AOI22_X1 U18060 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14605), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14582) );
  NAND2_X1 U18061 ( .A1(n9603), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n14578) );
  NAND2_X1 U18062 ( .A1(n14606), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n14576) );
  AND3_X1 U18063 ( .A1(n14578), .A2(n14577), .A3(n14576), .ZN(n14581) );
  AOI22_X1 U18064 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14611), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14579) );
  NAND4_X1 U18065 ( .A1(n14582), .A2(n14581), .A3(n14580), .A4(n14579), .ZN(
        n14590) );
  AOI22_X1 U18066 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14605), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14588) );
  NAND2_X1 U18067 ( .A1(n14509), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n14584) );
  NAND2_X1 U18068 ( .A1(n14611), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n14583) );
  AND3_X1 U18069 ( .A1(n14584), .A2(n14612), .A3(n14583), .ZN(n14587) );
  AOI22_X1 U18070 ( .A1(n14601), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14606), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14586) );
  NAND4_X1 U18071 ( .A1(n14588), .A2(n14587), .A3(n14586), .A4(n14585), .ZN(
        n14589) );
  NAND2_X1 U18072 ( .A1(n14590), .A2(n14589), .ZN(n14595) );
  INV_X1 U18073 ( .A(n14591), .ZN(n15982) );
  INV_X1 U18074 ( .A(n15983), .ZN(n14592) );
  NAND2_X1 U18075 ( .A1(n15982), .A2(n14593), .ZN(n14594) );
  NOR2_X1 U18076 ( .A1(n14594), .A2(n14595), .ZN(n14596) );
  AOI21_X1 U18077 ( .B1(n14595), .B2(n14594), .A(n14596), .ZN(n15977) );
  AOI22_X1 U18078 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14605), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14600) );
  NAND2_X1 U18079 ( .A1(n14600), .A2(n14599), .ZN(n14619) );
  INV_X1 U18080 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14604) );
  AOI21_X1 U18081 ( .B1(n9604), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n14612), .ZN(n14603) );
  AOI22_X1 U18082 ( .A1(n14601), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14606), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14602) );
  OAI211_X1 U18083 ( .C1(n13854), .C2(n14604), .A(n14603), .B(n14602), .ZN(
        n14618) );
  AOI22_X1 U18084 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14605), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14609) );
  AOI22_X1 U18085 ( .A1(n14607), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14606), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14608) );
  NAND2_X1 U18086 ( .A1(n14609), .A2(n14608), .ZN(n14617) );
  NAND2_X1 U18087 ( .A1(n14509), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n14614) );
  NAND2_X1 U18088 ( .A1(n14611), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n14613) );
  NAND4_X1 U18089 ( .A1(n14615), .A2(n14614), .A3(n14613), .A4(n14612), .ZN(
        n14616) );
  OAI22_X1 U18090 ( .A1(n14619), .A2(n14618), .B1(n14617), .B2(n14616), .ZN(
        n14620) );
  INV_X1 U18091 ( .A(n14620), .ZN(n14621) );
  XNOR2_X1 U18092 ( .A(n14622), .B(n14621), .ZN(n14634) );
  AOI22_X1 U18093 ( .A1(n16161), .A2(n14624), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n19431), .ZN(n14626) );
  NAND2_X1 U18094 ( .A1(n16168), .A2(BUF2_REG_30__SCAN_IN), .ZN(n14625) );
  NAND2_X1 U18095 ( .A1(n14626), .A2(n14625), .ZN(n14628) );
  AND2_X1 U18096 ( .A1(n16162), .A2(BUF1_REG_30__SCAN_IN), .ZN(n14627) );
  OAI21_X1 U18097 ( .B1(n14634), .B2(n16171), .A(n14631), .ZN(P2_U2889) );
  MUX2_X1 U18098 ( .A(n16177), .B(n14632), .S(n9598), .Z(n14633) );
  OAI21_X1 U18099 ( .B1(n14634), .B2(n16061), .A(n14633), .ZN(P2_U2857) );
  INV_X1 U18100 ( .A(n15941), .ZN(n14641) );
  OAI21_X1 U18101 ( .B1(n16436), .B2(n14636), .A(n14635), .ZN(n14640) );
  AND3_X1 U18102 ( .A1(n14638), .A2(n16383), .A3(n14637), .ZN(n14639) );
  AOI211_X1 U18103 ( .C1(n14641), .C2(n16433), .A(n14640), .B(n14639), .ZN(
        n14645) );
  OR3_X1 U18104 ( .A1(n14643), .A2(n14642), .A3(n16439), .ZN(n14644) );
  OR2_X1 U18105 ( .A1(n14646), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n14649) );
  NAND2_X1 U18106 ( .A1(n14651), .A2(n14647), .ZN(n14648) );
  MUX2_X1 U18107 ( .A(n14649), .B(n14648), .S(n21173), .Z(P1_U3487) );
  INV_X1 U18108 ( .A(n14650), .ZN(n14668) );
  AOI22_X1 U18109 ( .A1(n14652), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n9614), .ZN(n14673) );
  AOI22_X1 U18110 ( .A1(n14652), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n9614), .ZN(n14653) );
  INV_X1 U18111 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21140) );
  INV_X1 U18112 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21131) );
  AND4_X1 U18113 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(P1_REIP_REG_10__SCAN_IN), .A4(P1_REIP_REG_9__SCAN_IN), .ZN(n14820)
         );
  INV_X1 U18114 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21117) );
  INV_X1 U18115 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21115) );
  NOR2_X1 U18116 ( .A1(n21117), .A2(n21115), .ZN(n14863) );
  NAND4_X1 U18117 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .A3(P1_REIP_REG_13__SCAN_IN), .A4(n14863), .ZN(n14815) );
  INV_X1 U18118 ( .A(n14815), .ZN(n14821) );
  NAND2_X1 U18119 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14816) );
  INV_X1 U18120 ( .A(n14816), .ZN(n14656) );
  NAND3_X1 U18121 ( .A1(n14820), .A2(n14821), .A3(n14656), .ZN(n14657) );
  NOR2_X1 U18122 ( .A1(n14814), .A2(n14657), .ZN(n14770) );
  INV_X1 U18123 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21126) );
  INV_X1 U18124 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21124) );
  NOR2_X1 U18125 ( .A1(n21126), .A2(n21124), .ZN(n14773) );
  NAND2_X1 U18126 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n14773), .ZN(n14758) );
  INV_X1 U18127 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n15100) );
  NOR2_X1 U18128 ( .A1(n14758), .A2(n15100), .ZN(n14658) );
  NAND2_X1 U18129 ( .A1(n14770), .A2(n14658), .ZN(n14745) );
  NOR2_X1 U18130 ( .A1(n21131), .A2(n14745), .ZN(n14737) );
  NAND3_X1 U18131 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .A3(n14737), .ZN(n14711) );
  INV_X1 U18132 ( .A(n14711), .ZN(n14659) );
  AND2_X1 U18133 ( .A1(n20345), .A2(n14659), .ZN(n14709) );
  NAND2_X1 U18134 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n14709), .ZN(n14694) );
  OR2_X1 U18135 ( .A1(n21140), .A2(n14694), .ZN(n14660) );
  NAND2_X1 U18136 ( .A1(n20346), .A2(n14660), .ZN(n14698) );
  NAND2_X1 U18137 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14661) );
  NAND2_X1 U18138 ( .A1(n20346), .A2(n14661), .ZN(n14662) );
  AND2_X1 U18139 ( .A1(n14698), .A2(n14662), .ZN(n14681) );
  AOI22_X1 U18140 ( .A1(n20350), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20369), .ZN(n14664) );
  OR3_X1 U18141 ( .A1(n20354), .A2(n14694), .A3(n21140), .ZN(n14685) );
  INV_X1 U18142 ( .A(n14685), .ZN(n14676) );
  NAND4_X1 U18143 ( .A1(n14676), .A2(P1_REIP_REG_30__SCAN_IN), .A3(
        P1_REIP_REG_29__SCAN_IN), .A4(n14665), .ZN(n14663) );
  OAI211_X1 U18144 ( .C1(n14681), .C2(n14665), .A(n14664), .B(n14663), .ZN(
        n14666) );
  OAI21_X1 U18145 ( .B1(n14668), .B2(n16908), .A(n14667), .ZN(P1_U2809) );
  INV_X1 U18146 ( .A(n14669), .ZN(n14670) );
  AOI22_X1 U18147 ( .A1(n14672), .A2(n14671), .B1(n14670), .B2(n11557), .ZN(
        n14675) );
  INV_X1 U18148 ( .A(n14673), .ZN(n14674) );
  XNOR2_X1 U18149 ( .A(n14675), .B(n14674), .ZN(n15290) );
  AOI21_X1 U18150 ( .B1(n14676), .B2(P1_REIP_REG_29__SCAN_IN), .A(
        P1_REIP_REG_30__SCAN_IN), .ZN(n14680) );
  NAND2_X1 U18151 ( .A1(n20375), .A2(n14677), .ZN(n14679) );
  AOI22_X1 U18152 ( .A1(n20350), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20369), .ZN(n14678) );
  OAI211_X1 U18153 ( .C1(n14681), .C2(n14680), .A(n14679), .B(n14678), .ZN(
        n14682) );
  AOI21_X1 U18154 ( .B1(n15290), .B2(n20367), .A(n14682), .ZN(n14683) );
  NAND2_X1 U18155 ( .A1(n15054), .A2(n20333), .ZN(n14690) );
  INV_X1 U18156 ( .A(n14698), .ZN(n14688) );
  AOI22_X1 U18157 ( .A1(n20350), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20369), .ZN(n14684) );
  OAI21_X1 U18158 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(n14685), .A(n14684), 
        .ZN(n14687) );
  NOR2_X1 U18159 ( .A1(n20358), .A2(n15052), .ZN(n14686) );
  AOI211_X1 U18160 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n14688), .A(n14687), 
        .B(n14686), .ZN(n14689) );
  OAI211_X1 U18161 ( .C1(n15297), .C2(n20325), .A(n14690), .B(n14689), .ZN(
        P1_U2811) );
  OAI21_X1 U18162 ( .B1(n14691), .B2(n14692), .A(n11381), .ZN(n15066) );
  AOI21_X1 U18163 ( .B1(n14693), .B2(n14705), .A(n11557), .ZN(n15301) );
  INV_X1 U18164 ( .A(n14694), .ZN(n14695) );
  NOR2_X1 U18165 ( .A1(n14695), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14699) );
  NAND2_X1 U18166 ( .A1(n20375), .A2(n15058), .ZN(n14697) );
  AOI22_X1 U18167 ( .A1(n20350), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20369), .ZN(n14696) );
  OAI211_X1 U18168 ( .C1(n14699), .C2(n14698), .A(n14697), .B(n14696), .ZN(
        n14700) );
  AOI21_X1 U18169 ( .B1(n15301), .B2(n20367), .A(n14700), .ZN(n14701) );
  OAI21_X1 U18170 ( .B1(n15066), .B2(n16908), .A(n14701), .ZN(P1_U2812) );
  OR2_X1 U18171 ( .A1(n14702), .A2(n14703), .ZN(n14704) );
  NAND2_X1 U18172 ( .A1(n14705), .A2(n14704), .ZN(n15314) );
  BUF_X1 U18173 ( .A(n14706), .Z(n14707) );
  NAND2_X1 U18174 ( .A1(n15075), .A2(n20333), .ZN(n14717) );
  INV_X1 U18175 ( .A(n15073), .ZN(n14715) );
  INV_X1 U18176 ( .A(n14709), .ZN(n14710) );
  NAND2_X1 U18177 ( .A1(n20346), .A2(n14710), .ZN(n14723) );
  INV_X1 U18178 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n15071) );
  AOI22_X1 U18179 ( .A1(n20350), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20369), .ZN(n14713) );
  OR3_X1 U18180 ( .A1(n20354), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14711), .ZN(
        n14712) );
  OAI211_X1 U18181 ( .C1(n14723), .C2(n15071), .A(n14713), .B(n14712), .ZN(
        n14714) );
  AOI21_X1 U18182 ( .B1(n20375), .B2(n14715), .A(n14714), .ZN(n14716) );
  OAI211_X1 U18183 ( .C1(n15314), .C2(n20325), .A(n14717), .B(n14716), .ZN(
        P1_U2813) );
  OAI21_X1 U18184 ( .B1(n14719), .B2(n14720), .A(n14707), .ZN(n15085) );
  AOI21_X1 U18185 ( .B1(n14721), .B2(n14734), .A(n14702), .ZN(n15321) );
  INV_X1 U18186 ( .A(n15079), .ZN(n14728) );
  AOI22_X1 U18187 ( .A1(n20350), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20369), .ZN(n14727) );
  NAND2_X1 U18188 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n14737), .ZN(n14722) );
  NOR2_X1 U18189 ( .A1(n20354), .A2(n14722), .ZN(n14725) );
  INV_X1 U18190 ( .A(n14723), .ZN(n14724) );
  OAI21_X1 U18191 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n14725), .A(n14724), 
        .ZN(n14726) );
  OAI211_X1 U18192 ( .C1(n20358), .C2(n14728), .A(n14727), .B(n14726), .ZN(
        n14729) );
  AOI21_X1 U18193 ( .B1(n15321), .B2(n20367), .A(n14729), .ZN(n14730) );
  OAI21_X1 U18194 ( .B1(n15085), .B2(n16908), .A(n14730), .ZN(P1_U2814) );
  AOI21_X1 U18195 ( .B1(n14732), .B2(n14743), .A(n14719), .ZN(n15090) );
  INV_X1 U18196 ( .A(n15090), .ZN(n14990) );
  AOI21_X1 U18197 ( .B1(n14735), .B2(n14733), .A(n11543), .ZN(n15332) );
  NOR2_X1 U18198 ( .A1(n20358), .A2(n15088), .ZN(n14741) );
  OAI21_X1 U18199 ( .B1(n20326), .B2(n14745), .A(n20346), .ZN(n14759) );
  INV_X1 U18200 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21133) );
  AOI22_X1 U18201 ( .A1(n20350), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20369), .ZN(n14739) );
  NAND2_X1 U18202 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14736) );
  OAI211_X1 U18203 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14737), .A(n20327), 
        .B(n14736), .ZN(n14738) );
  OAI211_X1 U18204 ( .C1(n14759), .C2(n21133), .A(n14739), .B(n14738), .ZN(
        n14740) );
  AOI211_X1 U18205 ( .C1(n15332), .C2(n20367), .A(n14741), .B(n14740), .ZN(
        n14742) );
  OAI21_X1 U18206 ( .B1(n14990), .B2(n16908), .A(n14742), .ZN(P1_U2815) );
  OAI21_X1 U18207 ( .B1(n14752), .B2(n14744), .A(n14743), .ZN(n15097) );
  AOI22_X1 U18208 ( .A1(n20350), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20369), .ZN(n14747) );
  OR3_X1 U18209 ( .A1(n20354), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n14745), .ZN(
        n14746) );
  OAI211_X1 U18210 ( .C1(n14759), .C2(n21131), .A(n14747), .B(n14746), .ZN(
        n14750) );
  OAI21_X1 U18211 ( .B1(n9737), .B2(n14748), .A(n14733), .ZN(n15336) );
  NOR2_X1 U18212 ( .A1(n15336), .A2(n20325), .ZN(n14749) );
  AOI211_X1 U18213 ( .C1(n20375), .C2(n15094), .A(n14750), .B(n14749), .ZN(
        n14751) );
  OAI21_X1 U18214 ( .B1(n15097), .B2(n16908), .A(n14751), .ZN(P1_U2816) );
  AOI21_X1 U18215 ( .B1(n14753), .B2(n14767), .A(n14752), .ZN(n15104) );
  INV_X1 U18216 ( .A(n15104), .ZN(n14996) );
  AND2_X1 U18217 ( .A1(n14755), .A2(n14754), .ZN(n14756) );
  NOR2_X1 U18218 ( .A1(n9737), .A2(n14756), .ZN(n15348) );
  AOI22_X1 U18219 ( .A1(n20350), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20369), .ZN(n14763) );
  INV_X1 U18220 ( .A(n14770), .ZN(n14757) );
  OR2_X1 U18221 ( .A1(n20354), .A2(n14757), .ZN(n14772) );
  NOR2_X1 U18222 ( .A1(n14772), .A2(n14758), .ZN(n14761) );
  INV_X1 U18223 ( .A(n14759), .ZN(n14760) );
  OAI21_X1 U18224 ( .B1(n14761), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14760), 
        .ZN(n14762) );
  OAI211_X1 U18225 ( .C1(n20358), .C2(n15102), .A(n14763), .B(n14762), .ZN(
        n14764) );
  AOI21_X1 U18226 ( .B1(n15348), .B2(n20367), .A(n14764), .ZN(n14765) );
  OAI21_X1 U18227 ( .B1(n14996), .B2(n16908), .A(n14765), .ZN(P1_U2817) );
  INV_X1 U18228 ( .A(n14767), .ZN(n14768) );
  AOI21_X1 U18229 ( .B1(n14769), .B2(n14766), .A(n14768), .ZN(n15113) );
  INV_X1 U18230 ( .A(n15113), .ZN(n15000) );
  NAND3_X1 U18231 ( .A1(n20345), .A2(n14770), .A3(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n14771) );
  NAND2_X1 U18232 ( .A1(n20346), .A2(n14771), .ZN(n14800) );
  OAI21_X1 U18233 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n20354), .A(n14800), 
        .ZN(n14780) );
  INV_X1 U18234 ( .A(n15109), .ZN(n14776) );
  AOI22_X1 U18235 ( .A1(n20350), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20369), .ZN(n14775) );
  INV_X1 U18236 ( .A(n14772), .ZN(n14802) );
  INV_X1 U18237 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21128) );
  NAND3_X1 U18238 ( .A1(n14802), .A2(n14773), .A3(n21128), .ZN(n14774) );
  OAI211_X1 U18239 ( .C1(n20358), .C2(n14776), .A(n14775), .B(n14774), .ZN(
        n14779) );
  XNOR2_X1 U18240 ( .A(n14782), .B(n14777), .ZN(n15357) );
  NOR2_X1 U18241 ( .A1(n15357), .A2(n20325), .ZN(n14778) );
  AOI211_X1 U18242 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n14780), .A(n14779), 
        .B(n14778), .ZN(n14781) );
  OAI21_X1 U18243 ( .B1(n15000), .B2(n16908), .A(n14781), .ZN(P1_U2818) );
  OAI21_X1 U18244 ( .B1(n14799), .B2(n14783), .A(n14782), .ZN(n15369) );
  INV_X1 U18245 ( .A(n14766), .ZN(n14786) );
  AOI21_X1 U18246 ( .B1(n14787), .B2(n14785), .A(n14786), .ZN(n15123) );
  NAND2_X1 U18247 ( .A1(n15123), .A2(n20333), .ZN(n14793) );
  INV_X1 U18248 ( .A(n15119), .ZN(n14791) );
  NAND3_X1 U18249 ( .A1(n14802), .A2(P1_REIP_REG_20__SCAN_IN), .A3(n21126), 
        .ZN(n14789) );
  AOI22_X1 U18250 ( .A1(n20350), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20369), .ZN(n14788) );
  OAI211_X1 U18251 ( .C1(n14800), .C2(n21126), .A(n14789), .B(n14788), .ZN(
        n14790) );
  AOI21_X1 U18252 ( .B1(n20375), .B2(n14791), .A(n14790), .ZN(n14792) );
  OAI211_X1 U18253 ( .C1(n15369), .C2(n20325), .A(n14793), .B(n14792), .ZN(
        P1_U2819) );
  OAI21_X1 U18254 ( .B1(n14794), .B2(n14795), .A(n14785), .ZN(n15135) );
  NOR2_X1 U18255 ( .A1(n14796), .A2(n14797), .ZN(n14798) );
  OR2_X1 U18256 ( .A1(n14799), .A2(n14798), .ZN(n15380) );
  INV_X1 U18257 ( .A(n15380), .ZN(n14807) );
  NAND2_X1 U18258 ( .A1(n20375), .A2(n15127), .ZN(n14805) );
  AOI22_X1 U18259 ( .A1(n20350), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20369), .ZN(n14804) );
  INV_X1 U18260 ( .A(n14800), .ZN(n14801) );
  OAI21_X1 U18261 ( .B1(n14802), .B2(P1_REIP_REG_20__SCAN_IN), .A(n14801), 
        .ZN(n14803) );
  NAND3_X1 U18262 ( .A1(n14805), .A2(n14804), .A3(n14803), .ZN(n14806) );
  AOI21_X1 U18263 ( .B1(n14807), .B2(n20367), .A(n14806), .ZN(n14808) );
  OAI21_X1 U18264 ( .B1(n15135), .B2(n16908), .A(n14808), .ZN(P1_U2820) );
  AND2_X1 U18265 ( .A1(n14809), .A2(n14810), .ZN(n14811) );
  OR2_X1 U18266 ( .A1(n14811), .A2(n14794), .ZN(n15142) );
  AND2_X1 U18267 ( .A1(n14829), .A2(n14812), .ZN(n14813) );
  NOR2_X1 U18268 ( .A1(n14796), .A2(n14813), .ZN(n15395) );
  NAND2_X1 U18269 ( .A1(n20308), .A2(n14820), .ZN(n14909) );
  NOR2_X1 U18270 ( .A1(n14815), .A2(n14909), .ZN(n14832) );
  OAI211_X1 U18271 ( .C1(P1_REIP_REG_19__SCAN_IN), .C2(P1_REIP_REG_18__SCAN_IN), .A(n14832), .B(n14816), .ZN(n14817) );
  INV_X2 U18272 ( .A(n16962), .ZN(n20348) );
  OAI211_X1 U18273 ( .C1(n20336), .C2(n14818), .A(n14817), .B(n20348), .ZN(
        n14819) );
  AOI21_X1 U18274 ( .B1(n20350), .B2(P1_EBX_REG_19__SCAN_IN), .A(n14819), .ZN(
        n14824) );
  NAND2_X1 U18275 ( .A1(n14934), .A2(n14820), .ZN(n14857) );
  NAND2_X1 U18276 ( .A1(n20346), .A2(n14857), .ZN(n14923) );
  OAI21_X1 U18277 ( .B1(n14822), .B2(n14821), .A(n14923), .ZN(n14845) );
  NAND2_X1 U18278 ( .A1(n14845), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n14823) );
  OAI211_X1 U18279 ( .C1(n20358), .C2(n15138), .A(n14824), .B(n14823), .ZN(
        n14825) );
  AOI21_X1 U18280 ( .B1(n15395), .B2(n20367), .A(n14825), .ZN(n14826) );
  OAI21_X1 U18281 ( .B1(n15142), .B2(n16908), .A(n14826), .ZN(P1_U2821) );
  OAI21_X1 U18282 ( .B1(n10148), .B2(n10566), .A(n14809), .ZN(n15150) );
  INV_X1 U18283 ( .A(n14829), .ZN(n14830) );
  AOI21_X1 U18284 ( .B1(n14831), .B2(n14843), .A(n14830), .ZN(n15408) );
  INV_X1 U18285 ( .A(n15145), .ZN(n14837) );
  INV_X1 U18286 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21120) );
  AOI21_X1 U18287 ( .B1(n14832), .B2(n21120), .A(n16962), .ZN(n14833) );
  OAI21_X1 U18288 ( .B1(n15143), .B2(n20336), .A(n14833), .ZN(n14834) );
  AOI21_X1 U18289 ( .B1(n20350), .B2(P1_EBX_REG_18__SCAN_IN), .A(n14834), .ZN(
        n14836) );
  NAND2_X1 U18290 ( .A1(n14845), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14835) );
  OAI211_X1 U18291 ( .C1(n20358), .C2(n14837), .A(n14836), .B(n14835), .ZN(
        n14838) );
  AOI21_X1 U18292 ( .B1(n15408), .B2(n20367), .A(n14838), .ZN(n14839) );
  OAI21_X1 U18293 ( .B1(n15150), .B2(n16908), .A(n14839), .ZN(P1_U2822) );
  OAI21_X1 U18294 ( .B1(n14840), .B2(n14841), .A(n14828), .ZN(n15156) );
  OR2_X1 U18295 ( .A1(n14859), .A2(n14842), .ZN(n14844) );
  AND2_X1 U18296 ( .A1(n14844), .A2(n14843), .ZN(n15420) );
  INV_X1 U18297 ( .A(n14845), .ZN(n14851) );
  INV_X1 U18298 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21112) );
  INV_X1 U18299 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21111) );
  NOR3_X1 U18300 ( .A1(n21112), .A2(n21111), .A3(n14909), .ZN(n14881) );
  AOI21_X1 U18301 ( .B1(n14863), .B2(n14881), .A(P1_REIP_REG_17__SCAN_IN), 
        .ZN(n14850) );
  OAI21_X1 U18302 ( .B1(n20336), .B2(n14846), .A(n20348), .ZN(n14848) );
  NOR2_X1 U18303 ( .A1(n20358), .A2(n15159), .ZN(n14847) );
  AOI211_X1 U18304 ( .C1(P1_EBX_REG_17__SCAN_IN), .C2(n20350), .A(n14848), .B(
        n14847), .ZN(n14849) );
  OAI21_X1 U18305 ( .B1(n14851), .B2(n14850), .A(n14849), .ZN(n14852) );
  AOI21_X1 U18306 ( .B1(n20367), .B2(n15420), .A(n14852), .ZN(n14853) );
  OAI21_X1 U18307 ( .B1(n15156), .B2(n16908), .A(n14853), .ZN(P1_U2823) );
  AND2_X1 U18308 ( .A1(n14854), .A2(n14855), .ZN(n14856) );
  OR2_X1 U18309 ( .A1(n14856), .A2(n14840), .ZN(n15173) );
  NAND2_X1 U18310 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n14858) );
  OAI21_X1 U18311 ( .B1(n14858), .B2(n14857), .A(n20346), .ZN(n14896) );
  INV_X1 U18312 ( .A(n14896), .ZN(n14880) );
  AOI21_X1 U18313 ( .B1(n14860), .B2(n14875), .A(n14859), .ZN(n14861) );
  INV_X1 U18314 ( .A(n14861), .ZN(n15424) );
  OAI21_X1 U18315 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n14881), .ZN(n14864) );
  NAND2_X1 U18316 ( .A1(n20369), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14862) );
  OAI211_X1 U18317 ( .C1(n14864), .C2(n14863), .A(n20348), .B(n14862), .ZN(
        n14865) );
  AOI21_X1 U18318 ( .B1(n20350), .B2(P1_EBX_REG_16__SCAN_IN), .A(n14865), .ZN(
        n14867) );
  NAND2_X1 U18319 ( .A1(n20375), .A2(n15170), .ZN(n14866) );
  OAI211_X1 U18320 ( .C1(n15424), .C2(n20325), .A(n14867), .B(n14866), .ZN(
        n14868) );
  AOI21_X1 U18321 ( .B1(n14880), .B2(P1_REIP_REG_16__SCAN_IN), .A(n14868), 
        .ZN(n14869) );
  OAI21_X1 U18322 ( .B1(n15173), .B2(n16908), .A(n14869), .ZN(P1_U2824) );
  OAI21_X1 U18323 ( .B1(n14932), .B2(n14110), .A(n14905), .ZN(n14870) );
  INV_X1 U18324 ( .A(n14871), .ZN(n14872) );
  OAI21_X1 U18325 ( .B1(n14885), .B2(n14872), .A(n14854), .ZN(n15184) );
  NAND2_X1 U18326 ( .A1(n14889), .A2(n14873), .ZN(n14874) );
  NAND2_X1 U18327 ( .A1(n14875), .A2(n14874), .ZN(n15439) );
  NOR2_X1 U18328 ( .A1(n15439), .A2(n20325), .ZN(n14879) );
  AOI21_X1 U18329 ( .B1(n20369), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16962), .ZN(n14877) );
  NAND2_X1 U18330 ( .A1(n20350), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n14876) );
  OAI211_X1 U18331 ( .C1(n20358), .C2(n15174), .A(n14877), .B(n14876), .ZN(
        n14878) );
  AOI211_X1 U18332 ( .C1(n14880), .C2(P1_REIP_REG_15__SCAN_IN), .A(n14879), 
        .B(n14878), .ZN(n14883) );
  NAND2_X1 U18333 ( .A1(n14881), .A2(n21115), .ZN(n14882) );
  OAI211_X1 U18334 ( .C1(n15184), .C2(n16908), .A(n14883), .B(n14882), .ZN(
        P1_U2825) );
  INV_X1 U18335 ( .A(n14884), .ZN(n14887) );
  INV_X1 U18336 ( .A(n14907), .ZN(n14886) );
  AOI21_X1 U18337 ( .B1(n14887), .B2(n14886), .A(n14885), .ZN(n15193) );
  INV_X1 U18338 ( .A(n15193), .ZN(n15027) );
  INV_X1 U18339 ( .A(n15191), .ZN(n14900) );
  INV_X1 U18340 ( .A(n14889), .ZN(n14890) );
  AOI21_X1 U18341 ( .B1(n14891), .B2(n14888), .A(n14890), .ZN(n15449) );
  INV_X1 U18342 ( .A(n15449), .ZN(n14895) );
  OAI21_X1 U18343 ( .B1(n20336), .B2(n14892), .A(n20348), .ZN(n14893) );
  AOI21_X1 U18344 ( .B1(n20350), .B2(P1_EBX_REG_14__SCAN_IN), .A(n14893), .ZN(
        n14894) );
  OAI21_X1 U18345 ( .B1(n14895), .B2(n20325), .A(n14894), .ZN(n14899) );
  OR2_X1 U18346 ( .A1(n21111), .A2(n14909), .ZN(n14897) );
  AOI21_X1 U18347 ( .B1(n14897), .B2(n21112), .A(n14896), .ZN(n14898) );
  AOI211_X1 U18348 ( .C1(n20375), .C2(n14900), .A(n14899), .B(n14898), .ZN(
        n14901) );
  OAI21_X1 U18349 ( .B1(n15027), .B2(n16908), .A(n14901), .ZN(P1_U2826) );
  INV_X1 U18350 ( .A(n14110), .ZN(n14904) );
  INV_X1 U18351 ( .A(n14902), .ZN(n14903) );
  OAI21_X1 U18352 ( .B1(n14904), .B2(n14903), .A(n14905), .ZN(n14931) );
  OAI21_X1 U18353 ( .B1(n14931), .B2(n14932), .A(n14905), .ZN(n14921) );
  NAND2_X1 U18354 ( .A1(n14921), .A2(n14920), .ZN(n14919) );
  INV_X1 U18355 ( .A(n14906), .ZN(n14908) );
  AOI21_X1 U18356 ( .B1(n14919), .B2(n14908), .A(n14907), .ZN(n15205) );
  INV_X1 U18357 ( .A(n15205), .ZN(n15030) );
  MUX2_X1 U18358 ( .A(n14923), .B(n14909), .S(n21111), .Z(n14918) );
  INV_X1 U18359 ( .A(n14888), .ZN(n14912) );
  AOI21_X1 U18360 ( .B1(n14939), .B2(n14927), .A(n14910), .ZN(n14911) );
  NOR2_X1 U18361 ( .A1(n14912), .A2(n14911), .ZN(n15453) );
  NAND2_X1 U18362 ( .A1(n20350), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n14913) );
  OAI211_X1 U18363 ( .C1(n20336), .C2(n14914), .A(n14913), .B(n20348), .ZN(
        n14916) );
  NOR2_X1 U18364 ( .A1(n20358), .A2(n15203), .ZN(n14915) );
  AOI211_X1 U18365 ( .C1(n15453), .C2(n20367), .A(n14916), .B(n14915), .ZN(
        n14917) );
  OAI211_X1 U18366 ( .C1(n15030), .C2(n16908), .A(n14918), .B(n14917), .ZN(
        P1_U2827) );
  OAI21_X1 U18367 ( .B1(n14921), .B2(n14920), .A(n14919), .ZN(n15215) );
  OAI21_X1 U18368 ( .B1(n20336), .B2(n14922), .A(n20348), .ZN(n14926) );
  NAND4_X1 U18369 ( .A1(n20308), .A2(P1_REIP_REG_10__SCAN_IN), .A3(
        P1_REIP_REG_11__SCAN_IN), .A4(P1_REIP_REG_9__SCAN_IN), .ZN(n14924) );
  INV_X1 U18370 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15207) );
  AOI21_X1 U18371 ( .B1(n14924), .B2(n15207), .A(n14923), .ZN(n14925) );
  AOI211_X1 U18372 ( .C1(P1_EBX_REG_12__SCAN_IN), .C2(n20350), .A(n14926), .B(
        n14925), .ZN(n14930) );
  INV_X1 U18373 ( .A(n15208), .ZN(n14928) );
  XOR2_X1 U18374 ( .A(n14927), .B(n14939), .Z(n15475) );
  AOI22_X1 U18375 ( .A1(n20375), .A2(n14928), .B1(n15475), .B2(n20367), .ZN(
        n14929) );
  OAI211_X1 U18376 ( .C1(n15215), .C2(n16908), .A(n14930), .B(n14929), .ZN(
        P1_U2828) );
  XOR2_X1 U18377 ( .A(n14932), .B(n14931), .Z(n15225) );
  NAND2_X1 U18378 ( .A1(n15225), .A2(n20333), .ZN(n14948) );
  NAND2_X1 U18379 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14943) );
  INV_X1 U18380 ( .A(n14943), .ZN(n14933) );
  NAND2_X1 U18381 ( .A1(n14934), .A2(n14933), .ZN(n14935) );
  AND2_X1 U18382 ( .A1(n20346), .A2(n14935), .ZN(n16906) );
  NOR2_X1 U18383 ( .A1(n14937), .A2(n14936), .ZN(n14938) );
  OR2_X1 U18384 ( .A1(n14939), .A2(n14938), .ZN(n15483) );
  OAI21_X1 U18385 ( .B1(n20336), .B2(n14940), .A(n20348), .ZN(n14941) );
  AOI21_X1 U18386 ( .B1(n20350), .B2(P1_EBX_REG_11__SCAN_IN), .A(n14941), .ZN(
        n14942) );
  OAI21_X1 U18387 ( .B1(n15483), .B2(n20325), .A(n14942), .ZN(n14946) );
  INV_X1 U18388 ( .A(n20308), .ZN(n14944) );
  NOR3_X1 U18389 ( .A1(n14944), .A2(P1_REIP_REG_11__SCAN_IN), .A3(n14943), 
        .ZN(n14945) );
  AOI211_X1 U18390 ( .C1(n16906), .C2(P1_REIP_REG_11__SCAN_IN), .A(n14946), 
        .B(n14945), .ZN(n14947) );
  OAI211_X1 U18391 ( .C1(n20358), .C2(n15223), .A(n14948), .B(n14947), .ZN(
        P1_U2829) );
  INV_X1 U18392 ( .A(n15283), .ZN(n14950) );
  INV_X1 U18393 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14949) );
  OAI22_X1 U18394 ( .A1(n14950), .A2(n14972), .B1(n14949), .B2(n20396), .ZN(
        P1_U2841) );
  AOI22_X1 U18395 ( .A1(n15290), .A2(n20391), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n14968), .ZN(n14951) );
  AOI22_X1 U18396 ( .A1(n15301), .A2(n20391), .B1(n14968), .B2(
        P1_EBX_REG_28__SCAN_IN), .ZN(n14952) );
  OAI21_X1 U18397 ( .B1(n15066), .B2(n14970), .A(n14952), .ZN(P1_U2844) );
  INV_X1 U18398 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14953) );
  INV_X1 U18399 ( .A(n15075), .ZN(n14985) );
  OAI222_X1 U18400 ( .A1(n15314), .A2(n14972), .B1(n14953), .B2(n20396), .C1(
        n14985), .C2(n14970), .ZN(P1_U2845) );
  AOI22_X1 U18401 ( .A1(n15321), .A2(n20391), .B1(n14968), .B2(
        P1_EBX_REG_26__SCAN_IN), .ZN(n14954) );
  OAI21_X1 U18402 ( .B1(n15085), .B2(n14970), .A(n14954), .ZN(P1_U2846) );
  AOI22_X1 U18403 ( .A1(n15332), .A2(n20391), .B1(n14968), .B2(
        P1_EBX_REG_25__SCAN_IN), .ZN(n14955) );
  OAI21_X1 U18404 ( .B1(n14990), .B2(n14970), .A(n14955), .ZN(P1_U2847) );
  INV_X1 U18405 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14956) );
  OAI222_X1 U18406 ( .A1(n15336), .A2(n14972), .B1(n14956), .B2(n20396), .C1(
        n15097), .C2(n14970), .ZN(P1_U2848) );
  AOI22_X1 U18407 ( .A1(n15348), .A2(n20391), .B1(n14968), .B2(
        P1_EBX_REG_23__SCAN_IN), .ZN(n14957) );
  OAI21_X1 U18408 ( .B1(n14996), .B2(n14970), .A(n14957), .ZN(P1_U2849) );
  OAI222_X1 U18409 ( .A1(n15000), .A2(n14970), .B1(n14972), .B2(n15357), .C1(
        n20396), .C2(n14958), .ZN(P1_U2850) );
  INV_X1 U18410 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14959) );
  INV_X1 U18411 ( .A(n15123), .ZN(n15004) );
  OAI222_X1 U18412 ( .A1(n15369), .A2(n14972), .B1(n14959), .B2(n20396), .C1(
        n15004), .C2(n14970), .ZN(P1_U2851) );
  INV_X1 U18413 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14960) );
  OAI222_X1 U18414 ( .A1(n15380), .A2(n14972), .B1(n14960), .B2(n20396), .C1(
        n15135), .C2(n14970), .ZN(P1_U2852) );
  AOI22_X1 U18415 ( .A1(n15395), .A2(n20391), .B1(n14968), .B2(
        P1_EBX_REG_19__SCAN_IN), .ZN(n14961) );
  OAI21_X1 U18416 ( .B1(n15142), .B2(n14970), .A(n14961), .ZN(P1_U2853) );
  AOI22_X1 U18417 ( .A1(n15408), .A2(n20391), .B1(n14968), .B2(
        P1_EBX_REG_18__SCAN_IN), .ZN(n14962) );
  OAI21_X1 U18418 ( .B1(n15150), .B2(n14970), .A(n14962), .ZN(P1_U2854) );
  AOI22_X1 U18419 ( .A1(n15420), .A2(n20391), .B1(n14968), .B2(
        P1_EBX_REG_17__SCAN_IN), .ZN(n14963) );
  OAI21_X1 U18420 ( .B1(n15156), .B2(n14970), .A(n14963), .ZN(P1_U2855) );
  OAI222_X1 U18421 ( .A1(n15424), .A2(n14972), .B1(n14964), .B2(n20396), .C1(
        n15173), .C2(n14970), .ZN(P1_U2856) );
  INV_X1 U18422 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14965) );
  OAI222_X1 U18423 ( .A1(n15439), .A2(n14972), .B1(n14965), .B2(n20396), .C1(
        n15184), .C2(n14970), .ZN(P1_U2857) );
  AOI22_X1 U18424 ( .A1(n15449), .A2(n20391), .B1(n14968), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n14966) );
  OAI21_X1 U18425 ( .B1(n15027), .B2(n14970), .A(n14966), .ZN(P1_U2858) );
  AOI22_X1 U18426 ( .A1(n15453), .A2(n20391), .B1(n14968), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14967) );
  OAI21_X1 U18427 ( .B1(n15030), .B2(n14970), .A(n14967), .ZN(P1_U2859) );
  AOI22_X1 U18428 ( .A1(n15475), .A2(n20391), .B1(n14968), .B2(
        P1_EBX_REG_12__SCAN_IN), .ZN(n14969) );
  OAI21_X1 U18429 ( .B1(n15215), .B2(n14970), .A(n14969), .ZN(P1_U2860) );
  INV_X1 U18430 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14971) );
  INV_X1 U18431 ( .A(n15225), .ZN(n15036) );
  OAI222_X1 U18432 ( .A1(n15483), .A2(n14972), .B1(n14971), .B2(n20396), .C1(
        n15036), .C2(n14970), .ZN(P1_U2861) );
  AOI22_X1 U18433 ( .A1(n15017), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n15041), .ZN(n14977) );
  NOR3_X1 U18434 ( .A1(n15041), .A2(n14974), .A3(n20524), .ZN(n14975) );
  MUX2_X1 U18435 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n20492), .Z(
        n20438) );
  AOI22_X1 U18436 ( .A1(n15020), .A2(n20438), .B1(n15018), .B2(DATAI_30_), 
        .ZN(n14976) );
  AOI22_X1 U18437 ( .A1(n15017), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n15041), .ZN(n14979) );
  AOI22_X1 U18438 ( .A1(n15020), .A2(n15028), .B1(n15018), .B2(DATAI_29_), 
        .ZN(n14978) );
  OAI211_X1 U18439 ( .C1(n14980), .C2(n15045), .A(n14979), .B(n14978), .ZN(
        P1_U2875) );
  AOI22_X1 U18440 ( .A1(n15017), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n15041), .ZN(n14982) );
  MUX2_X1 U18441 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n20492), .Z(
        n20436) );
  AOI22_X1 U18442 ( .A1(n15020), .A2(n20436), .B1(n15018), .B2(DATAI_28_), 
        .ZN(n14981) );
  OAI211_X1 U18443 ( .C1(n15066), .C2(n15045), .A(n14982), .B(n14981), .ZN(
        P1_U2876) );
  AOI22_X1 U18444 ( .A1(n15017), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n15041), .ZN(n14984) );
  MUX2_X1 U18445 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n20492), .Z(
        n20434) );
  AOI22_X1 U18446 ( .A1(n15020), .A2(n20434), .B1(n15018), .B2(DATAI_27_), 
        .ZN(n14983) );
  OAI211_X1 U18447 ( .C1(n14985), .C2(n15045), .A(n14984), .B(n14983), .ZN(
        P1_U2877) );
  AOI22_X1 U18448 ( .A1(n15017), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n15041), .ZN(n14987) );
  AOI22_X1 U18449 ( .A1(n15020), .A2(n20432), .B1(n15018), .B2(DATAI_26_), 
        .ZN(n14986) );
  OAI211_X1 U18450 ( .C1(n15085), .C2(n15045), .A(n14987), .B(n14986), .ZN(
        P1_U2878) );
  AOI22_X1 U18451 ( .A1(n15017), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n15041), .ZN(n14989) );
  AOI22_X1 U18452 ( .A1(n15020), .A2(n15042), .B1(n15018), .B2(DATAI_25_), 
        .ZN(n14988) );
  OAI211_X1 U18453 ( .C1(n14990), .C2(n15045), .A(n14989), .B(n14988), .ZN(
        P1_U2879) );
  AOI22_X1 U18454 ( .A1(n15017), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n15041), .ZN(n14992) );
  AOI22_X1 U18455 ( .A1(n15020), .A2(n20430), .B1(n15018), .B2(DATAI_24_), 
        .ZN(n14991) );
  OAI211_X1 U18456 ( .C1(n15097), .C2(n15045), .A(n14992), .B(n14991), .ZN(
        P1_U2880) );
  AOI22_X1 U18457 ( .A1(n15017), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n15041), .ZN(n14995) );
  AOI22_X1 U18458 ( .A1(n15020), .A2(n14993), .B1(n15018), .B2(DATAI_23_), 
        .ZN(n14994) );
  OAI211_X1 U18459 ( .C1(n14996), .C2(n15045), .A(n14995), .B(n14994), .ZN(
        P1_U2881) );
  AOI22_X1 U18460 ( .A1(n15017), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n15041), .ZN(n14999) );
  AOI22_X1 U18461 ( .A1(n15020), .A2(n14997), .B1(n15018), .B2(DATAI_22_), 
        .ZN(n14998) );
  OAI211_X1 U18462 ( .C1(n15000), .C2(n15045), .A(n14999), .B(n14998), .ZN(
        P1_U2882) );
  AOI22_X1 U18463 ( .A1(n15017), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n15041), .ZN(n15003) );
  AOI22_X1 U18464 ( .A1(n15020), .A2(n15001), .B1(n15018), .B2(DATAI_21_), 
        .ZN(n15002) );
  OAI211_X1 U18465 ( .C1(n15004), .C2(n15045), .A(n15003), .B(n15002), .ZN(
        P1_U2883) );
  AOI22_X1 U18466 ( .A1(n15017), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n15041), .ZN(n15007) );
  AOI22_X1 U18467 ( .A1(n15020), .A2(n15005), .B1(n15018), .B2(DATAI_20_), 
        .ZN(n15006) );
  OAI211_X1 U18468 ( .C1(n15135), .C2(n15045), .A(n15007), .B(n15006), .ZN(
        P1_U2884) );
  AOI22_X1 U18469 ( .A1(n15017), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n15041), .ZN(n15010) );
  AOI22_X1 U18470 ( .A1(n15020), .A2(n15008), .B1(n15018), .B2(DATAI_19_), 
        .ZN(n15009) );
  OAI211_X1 U18471 ( .C1(n15142), .C2(n15045), .A(n15010), .B(n15009), .ZN(
        P1_U2885) );
  AOI22_X1 U18472 ( .A1(n15017), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n15041), .ZN(n15013) );
  AOI22_X1 U18473 ( .A1(n15020), .A2(n15011), .B1(n15018), .B2(DATAI_18_), 
        .ZN(n15012) );
  OAI211_X1 U18474 ( .C1(n15150), .C2(n15045), .A(n15013), .B(n15012), .ZN(
        P1_U2886) );
  AOI22_X1 U18475 ( .A1(n15017), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n15041), .ZN(n15016) );
  AOI22_X1 U18476 ( .A1(n15020), .A2(n15014), .B1(n15018), .B2(DATAI_17_), 
        .ZN(n15015) );
  OAI211_X1 U18477 ( .C1(n15156), .C2(n15045), .A(n15016), .B(n15015), .ZN(
        P1_U2887) );
  AOI22_X1 U18478 ( .A1(n15017), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n15041), .ZN(n15022) );
  AOI22_X1 U18479 ( .A1(n15020), .A2(n15019), .B1(n15018), .B2(DATAI_16_), 
        .ZN(n15021) );
  OAI211_X1 U18480 ( .C1(n15173), .C2(n15045), .A(n15022), .B(n15021), .ZN(
        P1_U2888) );
  AOI22_X1 U18481 ( .A1(n15043), .A2(n15023), .B1(P1_EAX_REG_15__SCAN_IN), 
        .B2(n15041), .ZN(n15024) );
  OAI21_X1 U18482 ( .B1(n15184), .B2(n15045), .A(n15024), .ZN(P1_U2889) );
  INV_X1 U18483 ( .A(n20438), .ZN(n15026) );
  OAI222_X1 U18484 ( .A1(n15027), .A2(n15045), .B1(n15034), .B2(n15026), .C1(
        n15025), .C2(n15031), .ZN(P1_U2890) );
  AOI22_X1 U18485 ( .A1(n15043), .A2(n15028), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15041), .ZN(n15029) );
  OAI21_X1 U18486 ( .B1(n15030), .B2(n15045), .A(n15029), .ZN(P1_U2891) );
  INV_X1 U18487 ( .A(n20436), .ZN(n15033) );
  OAI222_X1 U18488 ( .A1(n15215), .A2(n15045), .B1(n15034), .B2(n15033), .C1(
        n15032), .C2(n15031), .ZN(P1_U2892) );
  AOI22_X1 U18489 ( .A1(n15043), .A2(n20434), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n15041), .ZN(n15035) );
  OAI21_X1 U18490 ( .B1(n15036), .B2(n15045), .A(n15035), .ZN(P1_U2893) );
  AND2_X1 U18491 ( .A1(n15038), .A2(n15037), .ZN(n15039) );
  INV_X1 U18492 ( .A(n20384), .ZN(n15046) );
  AOI22_X1 U18493 ( .A1(n15043), .A2(n15042), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15041), .ZN(n15044) );
  OAI21_X1 U18494 ( .B1(n15046), .B2(n15045), .A(n15044), .ZN(P1_U2895) );
  NAND2_X1 U18495 ( .A1(n15048), .A2(n15047), .ZN(n15049) );
  XNOR2_X1 U18496 ( .A(n15050), .B(n15049), .ZN(n15300) );
  INV_X1 U18497 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21138) );
  NOR2_X1 U18498 ( .A1(n20348), .A2(n21138), .ZN(n15295) );
  AOI21_X1 U18499 ( .B1(n16921), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15295), .ZN(n15051) );
  OAI21_X1 U18500 ( .B1(n15052), .B2(n16929), .A(n15051), .ZN(n15053) );
  OAI21_X1 U18501 ( .B1(n20293), .B2(n15300), .A(n15055), .ZN(P1_U2970) );
  NOR2_X1 U18502 ( .A1(n20348), .A2(n21140), .ZN(n15307) );
  NOR2_X1 U18503 ( .A1(n16937), .A2(n15056), .ZN(n15057) );
  AOI211_X1 U18504 ( .C1(n15058), .C2(n15241), .A(n15307), .B(n15057), .ZN(
        n15065) );
  NAND2_X1 U18505 ( .A1(n15080), .A2(n15059), .ZN(n15067) );
  NAND2_X1 U18506 ( .A1(n15216), .A2(n15265), .ZN(n15081) );
  NAND3_X1 U18507 ( .A1(n15099), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15081), .ZN(n15060) );
  NAND2_X1 U18508 ( .A1(n15067), .A2(n15060), .ZN(n15062) );
  INV_X1 U18509 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15317) );
  MUX2_X1 U18510 ( .A(n15317), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n15236), .Z(n15061) );
  NAND2_X1 U18511 ( .A1(n15062), .A2(n15061), .ZN(n15063) );
  XNOR2_X1 U18512 ( .A(n15063), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15302) );
  NAND2_X1 U18513 ( .A1(n15302), .A2(n16926), .ZN(n15064) );
  OAI211_X1 U18514 ( .C1(n15066), .C2(n20491), .A(n15065), .B(n15064), .ZN(
        P1_U2971) );
  NAND2_X1 U18515 ( .A1(n15067), .A2(n10583), .ZN(n15069) );
  NOR2_X1 U18516 ( .A1(n20348), .A2(n15071), .ZN(n15311) );
  AOI21_X1 U18517 ( .B1(n16921), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15311), .ZN(n15072) );
  OAI21_X1 U18518 ( .B1(n15073), .B2(n16929), .A(n15072), .ZN(n15074) );
  AOI21_X1 U18519 ( .B1(n15075), .B2(n16931), .A(n15074), .ZN(n15076) );
  OAI21_X1 U18520 ( .B1(n20293), .B2(n15315), .A(n15076), .ZN(P1_U2972) );
  INV_X1 U18521 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21135) );
  NOR2_X1 U18522 ( .A1(n20348), .A2(n21135), .ZN(n15320) );
  INV_X1 U18523 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15077) );
  NOR2_X1 U18524 ( .A1(n16937), .A2(n15077), .ZN(n15078) );
  AOI211_X1 U18525 ( .C1(n15241), .C2(n15079), .A(n15320), .B(n15078), .ZN(
        n15084) );
  XNOR2_X1 U18526 ( .A(n15082), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15319) );
  NAND2_X1 U18527 ( .A1(n15319), .A2(n16926), .ZN(n15083) );
  OAI211_X1 U18528 ( .C1(n15085), .C2(n20491), .A(n15084), .B(n15083), .ZN(
        P1_U2973) );
  NOR2_X1 U18529 ( .A1(n20348), .A2(n21133), .ZN(n15331) );
  AOI21_X1 U18530 ( .B1(n16921), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15331), .ZN(n15087) );
  OAI21_X1 U18531 ( .B1(n15088), .B2(n16929), .A(n15087), .ZN(n15089) );
  AOI21_X1 U18532 ( .B1(n15090), .B2(n16931), .A(n15089), .ZN(n15091) );
  OAI21_X1 U18533 ( .B1(n20293), .B2(n15334), .A(n15091), .ZN(P1_U2974) );
  NOR2_X1 U18534 ( .A1(n20348), .A2(n21131), .ZN(n15341) );
  NOR2_X1 U18535 ( .A1(n16937), .A2(n15092), .ZN(n15093) );
  AOI211_X1 U18536 ( .C1(n15241), .C2(n15094), .A(n15341), .B(n15093), .ZN(
        n15096) );
  XNOR2_X1 U18537 ( .A(n15236), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15098) );
  XNOR2_X1 U18538 ( .A(n15099), .B(n15098), .ZN(n15356) );
  NOR2_X1 U18539 ( .A1(n20348), .A2(n15100), .ZN(n15349) );
  AOI21_X1 U18540 ( .B1(n16921), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15349), .ZN(n15101) );
  OAI21_X1 U18541 ( .B1(n15102), .B2(n16929), .A(n15101), .ZN(n15103) );
  AOI21_X1 U18542 ( .B1(n15104), .B2(n16931), .A(n15103), .ZN(n15105) );
  OAI21_X1 U18543 ( .B1(n15356), .B2(n20293), .A(n15105), .ZN(P1_U2976) );
  NAND2_X1 U18544 ( .A1(n15107), .A2(n15106), .ZN(n15108) );
  XNOR2_X1 U18545 ( .A(n15108), .B(n15361), .ZN(n15368) );
  NAND2_X1 U18546 ( .A1(n15241), .A2(n15109), .ZN(n15110) );
  NAND2_X1 U18547 ( .A1(n16962), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15358) );
  OAI211_X1 U18548 ( .C1(n16937), .C2(n15111), .A(n15110), .B(n15358), .ZN(
        n15112) );
  AOI21_X1 U18549 ( .B1(n15113), .B2(n16931), .A(n15112), .ZN(n15114) );
  OAI21_X1 U18550 ( .B1(n20293), .B2(n15368), .A(n15114), .ZN(P1_U2977) );
  INV_X1 U18551 ( .A(n15115), .ZN(n15116) );
  NAND3_X1 U18552 ( .A1(n15116), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15216), .ZN(n15132) );
  NOR2_X1 U18553 ( .A1(n15117), .A2(n15236), .ZN(n15128) );
  NAND2_X1 U18554 ( .A1(n15128), .A2(n15386), .ZN(n15130) );
  OAI21_X1 U18555 ( .B1(n15132), .B2(n15386), .A(n15130), .ZN(n15118) );
  XNOR2_X1 U18556 ( .A(n15118), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15378) );
  NOR2_X1 U18557 ( .A1(n16929), .A2(n15119), .ZN(n15122) );
  OR2_X1 U18558 ( .A1(n20348), .A2(n21126), .ZN(n15370) );
  OAI21_X1 U18559 ( .B1(n16937), .B2(n15120), .A(n15370), .ZN(n15121) );
  AOI211_X1 U18560 ( .C1(n15123), .C2(n16931), .A(n15122), .B(n15121), .ZN(
        n15124) );
  OAI21_X1 U18561 ( .B1(n15378), .B2(n20293), .A(n15124), .ZN(P1_U2978) );
  NOR2_X1 U18562 ( .A1(n20348), .A2(n21124), .ZN(n15390) );
  NOR2_X1 U18563 ( .A1(n16937), .A2(n15125), .ZN(n15126) );
  AOI211_X1 U18564 ( .C1(n15241), .C2(n15127), .A(n15390), .B(n15126), .ZN(
        n15134) );
  INV_X1 U18565 ( .A(n15128), .ZN(n15129) );
  NAND3_X1 U18566 ( .A1(n15129), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n15132), .ZN(n15131) );
  OAI211_X1 U18567 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15132), .A(
        n15131), .B(n15130), .ZN(n15379) );
  NAND2_X1 U18568 ( .A1(n15379), .A2(n16926), .ZN(n15133) );
  OAI211_X1 U18569 ( .C1(n15135), .C2(n20491), .A(n15134), .B(n15133), .ZN(
        P1_U2979) );
  NOR2_X1 U18570 ( .A1(n15236), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15136) );
  MUX2_X1 U18571 ( .A(n15216), .B(n15136), .S(n15115), .Z(n15137) );
  XNOR2_X1 U18572 ( .A(n15137), .B(n15385), .ZN(n15402) );
  NAND2_X1 U18573 ( .A1(n15402), .A2(n16926), .ZN(n15141) );
  INV_X1 U18574 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21121) );
  NOR2_X1 U18575 ( .A1(n20348), .A2(n21121), .ZN(n15396) );
  NOR2_X1 U18576 ( .A1(n16929), .A2(n15138), .ZN(n15139) );
  AOI211_X1 U18577 ( .C1(n16921), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15396), .B(n15139), .ZN(n15140) );
  OAI211_X1 U18578 ( .C1(n20491), .C2(n15142), .A(n15141), .B(n15140), .ZN(
        P1_U2980) );
  NOR2_X1 U18579 ( .A1(n20348), .A2(n21120), .ZN(n15407) );
  NOR2_X1 U18580 ( .A1(n16937), .A2(n15143), .ZN(n15144) );
  AOI211_X1 U18581 ( .C1(n15241), .C2(n15145), .A(n15407), .B(n15144), .ZN(
        n15149) );
  OR2_X1 U18582 ( .A1(n15147), .A2(n15146), .ZN(n15404) );
  NAND3_X1 U18583 ( .A1(n15404), .A2(n15115), .A3(n16926), .ZN(n15148) );
  OAI211_X1 U18584 ( .C1(n15150), .C2(n20491), .A(n15149), .B(n15148), .ZN(
        P1_U2981) );
  NOR2_X1 U18585 ( .A1(n15236), .A2(n15152), .ZN(n15195) );
  NOR2_X1 U18586 ( .A1(n15236), .A2(n15471), .ZN(n15198) );
  XNOR2_X1 U18587 ( .A(n15155), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15422) );
  INV_X1 U18588 ( .A(n15156), .ZN(n15161) );
  INV_X1 U18589 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n15157) );
  NOR2_X1 U18590 ( .A1(n20348), .A2(n15157), .ZN(n15419) );
  AOI21_X1 U18591 ( .B1(n16921), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15419), .ZN(n15158) );
  OAI21_X1 U18592 ( .B1(n15159), .B2(n16929), .A(n15158), .ZN(n15160) );
  AOI21_X1 U18593 ( .B1(n15161), .B2(n16931), .A(n15160), .ZN(n15162) );
  OAI21_X1 U18594 ( .B1(n15422), .B2(n20293), .A(n15162), .ZN(P1_U2982) );
  OR2_X1 U18595 ( .A1(n15151), .A2(n15163), .ZN(n15177) );
  INV_X1 U18596 ( .A(n15177), .ZN(n15165) );
  OAI21_X1 U18597 ( .B1(n15165), .B2(n15164), .A(n15178), .ZN(n15167) );
  XNOR2_X1 U18598 ( .A(n15167), .B(n15166), .ZN(n15423) );
  NAND2_X1 U18599 ( .A1(n15423), .A2(n16926), .ZN(n15172) );
  NOR2_X1 U18600 ( .A1(n20348), .A2(n21117), .ZN(n15425) );
  NOR2_X1 U18601 ( .A1(n16937), .A2(n15168), .ZN(n15169) );
  AOI211_X1 U18602 ( .C1(n15241), .C2(n15170), .A(n15425), .B(n15169), .ZN(
        n15171) );
  OAI211_X1 U18603 ( .C1(n20491), .C2(n15173), .A(n15172), .B(n15171), .ZN(
        P1_U2983) );
  NOR2_X1 U18604 ( .A1(n20348), .A2(n21115), .ZN(n15435) );
  NOR2_X1 U18605 ( .A1(n16929), .A2(n15174), .ZN(n15175) );
  AOI211_X1 U18606 ( .C1(n16921), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15435), .B(n15175), .ZN(n15183) );
  NAND2_X1 U18607 ( .A1(n15177), .A2(n15176), .ZN(n15181) );
  NAND2_X1 U18608 ( .A1(n15179), .A2(n15178), .ZN(n15180) );
  XNOR2_X1 U18609 ( .A(n15181), .B(n15180), .ZN(n15442) );
  NAND2_X1 U18610 ( .A1(n15442), .A2(n16926), .ZN(n15182) );
  OAI211_X1 U18611 ( .C1(n15184), .C2(n20491), .A(n15183), .B(n15182), .ZN(
        P1_U2984) );
  OAI21_X1 U18612 ( .B1(n15187), .B2(n15186), .A(n15185), .ZN(n15189) );
  XNOR2_X1 U18613 ( .A(n15236), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15188) );
  XNOR2_X1 U18614 ( .A(n15189), .B(n15188), .ZN(n15451) );
  NOR2_X1 U18615 ( .A1(n20348), .A2(n21112), .ZN(n15448) );
  AOI21_X1 U18616 ( .B1(n16921), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15448), .ZN(n15190) );
  OAI21_X1 U18617 ( .B1(n15191), .B2(n16929), .A(n15190), .ZN(n15192) );
  AOI21_X1 U18618 ( .B1(n15193), .B2(n16931), .A(n15192), .ZN(n15194) );
  OAI21_X1 U18619 ( .B1(n15451), .B2(n20293), .A(n15194), .ZN(P1_U2985) );
  OR2_X1 U18620 ( .A1(n15151), .A2(n9637), .ZN(n15197) );
  INV_X1 U18621 ( .A(n15195), .ZN(n15196) );
  NOR2_X1 U18622 ( .A1(n15198), .A2(n10033), .ZN(n15211) );
  NAND2_X1 U18623 ( .A1(n15212), .A2(n15211), .ZN(n15210) );
  NAND2_X1 U18624 ( .A1(n15210), .A2(n15199), .ZN(n15201) );
  XNOR2_X1 U18625 ( .A(n15201), .B(n15200), .ZN(n15462) );
  NOR2_X1 U18626 ( .A1(n20348), .A2(n21111), .ZN(n15452) );
  AOI21_X1 U18627 ( .B1(n16921), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15452), .ZN(n15202) );
  OAI21_X1 U18628 ( .B1(n15203), .B2(n16929), .A(n15202), .ZN(n15204) );
  AOI21_X1 U18629 ( .B1(n15205), .B2(n16931), .A(n15204), .ZN(n15206) );
  OAI21_X1 U18630 ( .B1(n20293), .B2(n15462), .A(n15206), .ZN(P1_U2986) );
  NOR2_X1 U18631 ( .A1(n20348), .A2(n15207), .ZN(n15474) );
  NOR2_X1 U18632 ( .A1(n16929), .A2(n15208), .ZN(n15209) );
  AOI211_X1 U18633 ( .C1(n16921), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15474), .B(n15209), .ZN(n15214) );
  OAI21_X1 U18634 ( .B1(n15212), .B2(n15211), .A(n15210), .ZN(n15463) );
  NAND2_X1 U18635 ( .A1(n15463), .A2(n16926), .ZN(n15213) );
  OAI211_X1 U18636 ( .C1(n15215), .C2(n20491), .A(n15214), .B(n15213), .ZN(
        P1_U2987) );
  NAND3_X1 U18637 ( .A1(n15217), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15216), .ZN(n15220) );
  INV_X1 U18638 ( .A(n15218), .ZN(n15219) );
  NAND3_X1 U18639 ( .A1(n15219), .A2(n10583), .A3(n15227), .ZN(n15230) );
  NAND2_X1 U18640 ( .A1(n15220), .A2(n15230), .ZN(n15221) );
  XNOR2_X1 U18641 ( .A(n15221), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15491) );
  INV_X1 U18642 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21108) );
  NOR2_X1 U18643 ( .A1(n20348), .A2(n21108), .ZN(n15485) );
  AOI21_X1 U18644 ( .B1(n16921), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n15485), .ZN(n15222) );
  OAI21_X1 U18645 ( .B1(n15223), .B2(n16929), .A(n15222), .ZN(n15224) );
  AOI21_X1 U18646 ( .B1(n15225), .B2(n16931), .A(n15224), .ZN(n15226) );
  OAI21_X1 U18647 ( .B1(n15491), .B2(n20293), .A(n15226), .ZN(P1_U2988) );
  NAND2_X1 U18648 ( .A1(n15218), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15229) );
  XNOR2_X1 U18649 ( .A(n15151), .B(n15227), .ZN(n15228) );
  MUX2_X1 U18650 ( .A(n15229), .B(n15228), .S(n15216), .Z(n15231) );
  NAND2_X1 U18651 ( .A1(n15231), .A2(n15230), .ZN(n15492) );
  NAND2_X1 U18652 ( .A1(n15492), .A2(n16926), .ZN(n15235) );
  INV_X1 U18653 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15232) );
  NAND2_X1 U18654 ( .A1(n16962), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n15498) );
  OAI21_X1 U18655 ( .B1(n16937), .B2(n15232), .A(n15498), .ZN(n15233) );
  AOI21_X1 U18656 ( .B1(n15241), .B2(n16911), .A(n15233), .ZN(n15234) );
  OAI211_X1 U18657 ( .C1(n20491), .C2(n16909), .A(n15235), .B(n15234), .ZN(
        P1_U2989) );
  XNOR2_X1 U18658 ( .A(n15236), .B(n15512), .ZN(n15237) );
  NAND2_X1 U18659 ( .A1(n20384), .A2(n16931), .ZN(n15243) );
  INV_X1 U18660 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n15238) );
  NOR2_X1 U18661 ( .A1(n20348), .A2(n15238), .ZN(n15509) );
  INV_X1 U18662 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15239) );
  NOR2_X1 U18663 ( .A1(n16937), .A2(n15239), .ZN(n15240) );
  AOI211_X1 U18664 ( .C1(n15241), .C2(n20310), .A(n15509), .B(n15240), .ZN(
        n15242) );
  OAI211_X1 U18665 ( .C1(n15516), .C2(n20293), .A(n15243), .B(n15242), .ZN(
        P1_U2990) );
  INV_X1 U18666 ( .A(n16918), .ZN(n15246) );
  INV_X1 U18667 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16915) );
  AOI21_X1 U18668 ( .B1(n16918), .B2(n16915), .A(n15244), .ZN(n15245) );
  AOI21_X1 U18669 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15246), .A(
        n15245), .ZN(n15249) );
  XNOR2_X1 U18670 ( .A(n15247), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15248) );
  XNOR2_X1 U18671 ( .A(n15249), .B(n15248), .ZN(n16946) );
  INV_X1 U18672 ( .A(n15250), .ZN(n15254) );
  AOI22_X1 U18673 ( .A1(n16921), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16962), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n15251) );
  OAI21_X1 U18674 ( .B1(n15252), .B2(n16929), .A(n15251), .ZN(n15253) );
  AOI21_X1 U18675 ( .B1(n15254), .B2(n16931), .A(n15253), .ZN(n15255) );
  OAI21_X1 U18676 ( .B1(n16946), .B2(n20293), .A(n15255), .ZN(P1_U2991) );
  NAND2_X1 U18677 ( .A1(n15269), .A2(n15467), .ZN(n15263) );
  INV_X1 U18678 ( .A(n15263), .ZN(n15496) );
  NOR2_X1 U18679 ( .A1(n15496), .A2(n13463), .ZN(n15282) );
  NOR2_X1 U18680 ( .A1(n20461), .A2(n13206), .ZN(n16938) );
  NAND2_X1 U18681 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16938), .ZN(
        n15256) );
  NOR2_X1 U18682 ( .A1(n15476), .A2(n15256), .ZN(n15464) );
  AND2_X1 U18683 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15487) );
  NAND2_X1 U18684 ( .A1(n15487), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15494) );
  NAND2_X1 U18685 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15488) );
  NOR2_X1 U18686 ( .A1(n15494), .A2(n15488), .ZN(n15465) );
  NAND2_X1 U18687 ( .A1(n15465), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15479) );
  NOR2_X1 U18688 ( .A1(n15471), .A2(n15479), .ZN(n15381) );
  NAND2_X1 U18689 ( .A1(n15464), .A2(n15381), .ZN(n15454) );
  NOR2_X1 U18690 ( .A1(n15457), .A2(n15454), .ZN(n15270) );
  INV_X1 U18691 ( .A(n15270), .ZN(n15258) );
  NOR2_X1 U18692 ( .A1(n15256), .A2(n20459), .ZN(n16940) );
  AND2_X1 U18693 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15381), .ZN(
        n15257) );
  NAND2_X1 U18694 ( .A1(n16940), .A2(n15257), .ZN(n15271) );
  AOI22_X1 U18695 ( .A1(n16942), .A2(n15258), .B1(n20460), .B2(n15271), .ZN(
        n15259) );
  NAND2_X1 U18696 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15414) );
  NAND2_X1 U18697 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15260) );
  NOR2_X1 U18698 ( .A1(n15414), .A2(n15260), .ZN(n15410) );
  NAND2_X1 U18699 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15410), .ZN(
        n15274) );
  NAND2_X1 U18700 ( .A1(n16944), .A2(n15274), .ZN(n15261) );
  NAND2_X1 U18701 ( .A1(n15459), .A2(n15261), .ZN(n15397) );
  INV_X1 U18702 ( .A(n15262), .ZN(n15373) );
  NAND2_X1 U18703 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15364) );
  NAND2_X1 U18704 ( .A1(n16944), .A2(n15364), .ZN(n15264) );
  AND2_X1 U18705 ( .A1(n16944), .A2(n15265), .ZN(n15266) );
  AND2_X1 U18706 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15279) );
  INV_X1 U18707 ( .A(n15279), .ZN(n15267) );
  NAND2_X1 U18708 ( .A1(n16944), .A2(n15267), .ZN(n15268) );
  NAND2_X1 U18709 ( .A1(n15326), .A2(n15268), .ZN(n15312) );
  AOI21_X1 U18710 ( .B1(n10403), .B2(n16944), .A(n15312), .ZN(n15293) );
  OAI211_X1 U18711 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15269), .A(
        n15293), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15287) );
  NAND2_X1 U18712 ( .A1(n15478), .A2(n15270), .ZN(n15273) );
  OR2_X1 U18713 ( .A1(n16939), .A2(n15271), .ZN(n15272) );
  NAND2_X1 U18714 ( .A1(n15273), .A2(n15272), .ZN(n15445) );
  INV_X1 U18715 ( .A(n15274), .ZN(n15275) );
  NAND2_X1 U18716 ( .A1(n15445), .A2(n15275), .ZN(n15400) );
  NAND2_X1 U18717 ( .A1(n13248), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15276) );
  INV_X1 U18718 ( .A(n15277), .ZN(n15278) );
  NOR2_X1 U18719 ( .A1(n15353), .A2(n15278), .ZN(n15328) );
  NAND3_X1 U18720 ( .A1(n15318), .A2(n15304), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15288) );
  NOR3_X1 U18721 ( .A1(n15288), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n10045), .ZN(n15280) );
  AOI211_X1 U18722 ( .C1(n15282), .C2(n15287), .A(n15281), .B(n15280), .ZN(
        n15285) );
  NAND2_X1 U18723 ( .A1(n15283), .A2(n20473), .ZN(n15284) );
  OAI211_X1 U18724 ( .C1(n15286), .C2(n20481), .A(n15285), .B(n15284), .ZN(
        P1_U3000) );
  OAI21_X1 U18725 ( .B1(n15292), .B2(n20481), .A(n15291), .ZN(P1_U3001) );
  INV_X1 U18726 ( .A(n15293), .ZN(n15296) );
  INV_X1 U18727 ( .A(n15318), .ZN(n15305) );
  NOR3_X1 U18728 ( .A1(n15305), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n10403), .ZN(n15294) );
  AOI211_X1 U18729 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15296), .A(
        n15295), .B(n15294), .ZN(n15299) );
  NAND2_X1 U18730 ( .A1(n11561), .A2(n20473), .ZN(n15298) );
  OAI211_X1 U18731 ( .C1(n15300), .C2(n20481), .A(n15299), .B(n15298), .ZN(
        P1_U3002) );
  INV_X1 U18732 ( .A(n15301), .ZN(n15310) );
  NAND2_X1 U18733 ( .A1(n15302), .A2(n16965), .ZN(n15309) );
  NOR3_X1 U18734 ( .A1(n15305), .A2(n15304), .A3(n15303), .ZN(n15306) );
  AOI211_X1 U18735 ( .C1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15312), .A(
        n15307), .B(n15306), .ZN(n15308) );
  OAI211_X1 U18736 ( .C1(n20486), .C2(n15310), .A(n15309), .B(n15308), .ZN(
        P1_U3003) );
  AOI21_X1 U18737 ( .B1(n15312), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15311), .ZN(n15313) );
  OAI21_X1 U18738 ( .B1(n15314), .B2(n20486), .A(n15313), .ZN(n15316) );
  INV_X1 U18739 ( .A(n15319), .ZN(n15325) );
  AOI21_X1 U18740 ( .B1(n15321), .B2(n20473), .A(n15320), .ZN(n15324) );
  NAND2_X1 U18741 ( .A1(n15328), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15322) );
  MUX2_X1 U18742 ( .A(n15322), .B(n15326), .S(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n15323) );
  OAI211_X1 U18743 ( .C1(n15325), .C2(n20481), .A(n15324), .B(n15323), .ZN(
        P1_U3005) );
  INV_X1 U18744 ( .A(n15326), .ZN(n15329) );
  MUX2_X1 U18745 ( .A(n15329), .B(n15328), .S(n15327), .Z(n15330) );
  AOI211_X1 U18746 ( .C1(n15332), .C2(n20473), .A(n15331), .B(n15330), .ZN(
        n15333) );
  OAI21_X1 U18747 ( .B1(n15334), .B2(n20481), .A(n15333), .ZN(P1_U3006) );
  INV_X1 U18748 ( .A(n15335), .ZN(n15347) );
  INV_X1 U18749 ( .A(n15336), .ZN(n15342) );
  NAND2_X1 U18750 ( .A1(n16939), .A2(n16943), .ZN(n15338) );
  AOI21_X1 U18751 ( .B1(n15338), .B2(n15337), .A(n15350), .ZN(n15339) );
  NOR2_X1 U18752 ( .A1(n15339), .A2(n15343), .ZN(n15340) );
  AOI211_X1 U18753 ( .C1(n15342), .C2(n20473), .A(n15341), .B(n15340), .ZN(
        n15346) );
  INV_X1 U18754 ( .A(n15353), .ZN(n15344) );
  NAND3_X1 U18755 ( .A1(n15344), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n15343), .ZN(n15345) );
  OAI211_X1 U18756 ( .C1(n15347), .C2(n20481), .A(n15346), .B(n15345), .ZN(
        P1_U3007) );
  NAND2_X1 U18757 ( .A1(n15348), .A2(n20473), .ZN(n15352) );
  AOI21_X1 U18758 ( .B1(n15350), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15349), .ZN(n15351) );
  OAI211_X1 U18759 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n15353), .A(
        n15352), .B(n15351), .ZN(n15354) );
  INV_X1 U18760 ( .A(n15354), .ZN(n15355) );
  OAI21_X1 U18761 ( .B1(n15356), .B2(n20481), .A(n15355), .ZN(P1_U3008) );
  INV_X1 U18762 ( .A(n15357), .ZN(n15360) );
  OAI21_X1 U18763 ( .B1(n15372), .B2(n15361), .A(n15358), .ZN(n15359) );
  AOI21_X1 U18764 ( .B1(n15360), .B2(n20473), .A(n15359), .ZN(n15367) );
  INV_X1 U18765 ( .A(n15400), .ZN(n15365) );
  NAND2_X1 U18766 ( .A1(n15362), .A2(n15361), .ZN(n15363) );
  NAND3_X1 U18767 ( .A1(n15365), .A2(n15364), .A3(n15363), .ZN(n15366) );
  OAI211_X1 U18768 ( .C1(n15368), .C2(n20481), .A(n15367), .B(n15366), .ZN(
        P1_U3009) );
  INV_X1 U18769 ( .A(n15369), .ZN(n15376) );
  OAI21_X1 U18770 ( .B1(n15372), .B2(n15371), .A(n15370), .ZN(n15375) );
  NOR3_X1 U18771 ( .A1(n15400), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15373), .ZN(n15374) );
  AOI211_X1 U18772 ( .C1(n20473), .C2(n15376), .A(n15375), .B(n15374), .ZN(
        n15377) );
  OAI21_X1 U18773 ( .B1(n15378), .B2(n20481), .A(n15377), .ZN(P1_U3010) );
  INV_X1 U18774 ( .A(n15379), .ZN(n15394) );
  NOR3_X1 U18775 ( .A1(n15400), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n15385), .ZN(n15392) );
  NOR2_X1 U18776 ( .A1(n15380), .A2(n20486), .ZN(n15391) );
  INV_X1 U18777 ( .A(n15397), .ZN(n15388) );
  NAND2_X1 U18778 ( .A1(n16940), .A2(n15381), .ZN(n15384) );
  NAND2_X1 U18779 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15382), .ZN(
        n15383) );
  OAI22_X1 U18780 ( .A1(n16939), .A2(n15384), .B1(n15383), .B2(n15454), .ZN(
        n15455) );
  OAI21_X1 U18781 ( .B1(n15455), .B2(n20477), .A(n15385), .ZN(n15387) );
  AOI21_X1 U18782 ( .B1(n15388), .B2(n15387), .A(n15386), .ZN(n15389) );
  NOR4_X1 U18783 ( .A1(n15392), .A2(n15391), .A3(n15390), .A4(n15389), .ZN(
        n15393) );
  OAI21_X1 U18784 ( .B1(n15394), .B2(n20481), .A(n15393), .ZN(P1_U3011) );
  NAND2_X1 U18785 ( .A1(n15395), .A2(n20473), .ZN(n15399) );
  AOI21_X1 U18786 ( .B1(n15397), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15396), .ZN(n15398) );
  OAI211_X1 U18787 ( .C1(n15400), .C2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15399), .B(n15398), .ZN(n15401) );
  AOI21_X1 U18788 ( .B1(n15402), .B2(n16965), .A(n15401), .ZN(n15403) );
  INV_X1 U18789 ( .A(n15403), .ZN(P1_U3012) );
  NAND3_X1 U18790 ( .A1(n15404), .A2(n15115), .A3(n16965), .ZN(n15413) );
  INV_X1 U18791 ( .A(n15410), .ZN(n15405) );
  INV_X1 U18792 ( .A(n15459), .ZN(n15446) );
  AOI21_X1 U18793 ( .B1(n16944), .B2(n15405), .A(n15446), .ZN(n15416) );
  NOR2_X1 U18794 ( .A1(n15416), .A2(n15409), .ZN(n15406) );
  AOI211_X1 U18795 ( .C1(n15408), .C2(n20473), .A(n15407), .B(n15406), .ZN(
        n15412) );
  NAND3_X1 U18796 ( .A1(n15445), .A2(n15410), .A3(n15409), .ZN(n15411) );
  NAND3_X1 U18797 ( .A1(n15413), .A2(n15412), .A3(n15411), .ZN(P1_U3013) );
  INV_X1 U18798 ( .A(n15445), .ZN(n15415) );
  NOR2_X1 U18799 ( .A1(n15415), .A2(n15414), .ZN(n15428) );
  AOI21_X1 U18800 ( .B1(n15428), .B2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15417) );
  NOR2_X1 U18801 ( .A1(n15417), .A2(n15416), .ZN(n15418) );
  AOI211_X1 U18802 ( .C1(n20473), .C2(n15420), .A(n15419), .B(n15418), .ZN(
        n15421) );
  OAI21_X1 U18803 ( .B1(n15422), .B2(n20481), .A(n15421), .ZN(P1_U3014) );
  INV_X1 U18804 ( .A(n15423), .ZN(n15434) );
  NOR2_X1 U18805 ( .A1(n15424), .A2(n20486), .ZN(n15426) );
  AOI211_X1 U18806 ( .C1(n15428), .C2(n15427), .A(n15426), .B(n15425), .ZN(
        n15433) );
  AND2_X1 U18807 ( .A1(n15429), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15430) );
  AND2_X1 U18808 ( .A1(n15445), .A2(n15430), .ZN(n15441) );
  NAND2_X1 U18809 ( .A1(n16944), .A2(n15444), .ZN(n15431) );
  NAND2_X1 U18810 ( .A1(n15459), .A2(n15431), .ZN(n15436) );
  OAI21_X1 U18811 ( .B1(n15441), .B2(n15436), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15432) );
  OAI211_X1 U18812 ( .C1(n15434), .C2(n20481), .A(n15433), .B(n15432), .ZN(
        P1_U3015) );
  INV_X1 U18813 ( .A(n15435), .ZN(n15438) );
  NAND2_X1 U18814 ( .A1(n15436), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15437) );
  OAI211_X1 U18815 ( .C1(n15439), .C2(n20486), .A(n15438), .B(n15437), .ZN(
        n15440) );
  AOI211_X1 U18816 ( .C1(n15442), .C2(n16965), .A(n15441), .B(n15440), .ZN(
        n15443) );
  INV_X1 U18817 ( .A(n15443), .ZN(P1_U3016) );
  MUX2_X1 U18818 ( .A(n15446), .B(n15445), .S(n15444), .Z(n15447) );
  AOI211_X1 U18819 ( .C1(n20473), .C2(n15449), .A(n15448), .B(n15447), .ZN(
        n15450) );
  OAI21_X1 U18820 ( .B1(n15451), .B2(n20481), .A(n15450), .ZN(P1_U3017) );
  AOI21_X1 U18821 ( .B1(n15453), .B2(n20473), .A(n15452), .ZN(n15461) );
  INV_X1 U18822 ( .A(n15454), .ZN(n15456) );
  AOI21_X1 U18823 ( .B1(n20477), .B2(n15456), .A(n15455), .ZN(n15458) );
  MUX2_X1 U18824 ( .A(n15459), .B(n15458), .S(n15457), .Z(n15460) );
  OAI211_X1 U18825 ( .C1(n15462), .C2(n20481), .A(n15461), .B(n15460), .ZN(
        P1_U3018) );
  INV_X1 U18826 ( .A(n15463), .ZN(n15482) );
  INV_X1 U18827 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15470) );
  AND2_X1 U18828 ( .A1(n15465), .A2(n15464), .ZN(n15468) );
  INV_X1 U18829 ( .A(n16940), .ZN(n15495) );
  OAI21_X1 U18830 ( .B1(n15495), .B2(n15479), .A(n20460), .ZN(n15466) );
  OAI211_X1 U18831 ( .C1(n15469), .C2(n15468), .A(n15467), .B(n15466), .ZN(
        n15486) );
  AOI21_X1 U18832 ( .B1(n15478), .B2(n15470), .A(n15486), .ZN(n15472) );
  NOR2_X1 U18833 ( .A1(n15472), .A2(n15471), .ZN(n15473) );
  AOI211_X1 U18834 ( .C1(n20473), .C2(n15475), .A(n15474), .B(n15473), .ZN(
        n15481) );
  INV_X1 U18835 ( .A(n15476), .ZN(n15477) );
  OR3_X1 U18836 ( .A1(n16968), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n15479), .ZN(n15480) );
  OAI211_X1 U18837 ( .C1(n15482), .C2(n20481), .A(n15481), .B(n15480), .ZN(
        P1_U3019) );
  NOR2_X1 U18838 ( .A1(n15483), .A2(n20486), .ZN(n15484) );
  AOI211_X1 U18839 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15486), .A(
        n15485), .B(n15484), .ZN(n15490) );
  NAND2_X1 U18840 ( .A1(n16956), .A2(n15487), .ZN(n15511) );
  OR3_X1 U18841 ( .A1(n15511), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n15488), .ZN(n15489) );
  OAI211_X1 U18842 ( .C1(n15491), .C2(n20481), .A(n15490), .B(n15489), .ZN(
        P1_U3020) );
  XNOR2_X1 U18843 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15502) );
  NAND2_X1 U18844 ( .A1(n15492), .A2(n16965), .ZN(n15501) );
  NOR3_X1 U18845 ( .A1(n20458), .A2(n15495), .A3(n15494), .ZN(n15497) );
  NOR2_X1 U18846 ( .A1(n15497), .A2(n15496), .ZN(n15510) );
  OAI21_X1 U18847 ( .B1(n16914), .B2(n20486), .A(n15498), .ZN(n15499) );
  AOI21_X1 U18848 ( .B1(n15510), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n15499), .ZN(n15500) );
  OAI211_X1 U18849 ( .C1(n15511), .C2(n15502), .A(n15501), .B(n15500), .ZN(
        P1_U3021) );
  NAND2_X1 U18850 ( .A1(n15504), .A2(n15503), .ZN(n15505) );
  AND2_X1 U18851 ( .A1(n15506), .A2(n15505), .ZN(n20383) );
  INV_X1 U18852 ( .A(n20383), .ZN(n15507) );
  NOR2_X1 U18853 ( .A1(n20486), .A2(n15507), .ZN(n15508) );
  AOI211_X1 U18854 ( .C1(n15510), .C2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15509), .B(n15508), .ZN(n15515) );
  INV_X1 U18855 ( .A(n15511), .ZN(n15513) );
  NAND2_X1 U18856 ( .A1(n15513), .A2(n15512), .ZN(n15514) );
  OAI211_X1 U18857 ( .C1(n15516), .C2(n20481), .A(n15515), .B(n15514), .ZN(
        P1_U3022) );
  NAND2_X1 U18858 ( .A1(n20774), .A2(n16847), .ZN(n15533) );
  MUX2_X1 U18859 ( .A(n15518), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n13457), .Z(n15520) );
  NOR2_X1 U18860 ( .A1(n15520), .A2(n15519), .ZN(n15530) );
  AOI21_X1 U18861 ( .B1(n13457), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n15523), .ZN(n15521) );
  NOR2_X1 U18862 ( .A1(n15522), .A2(n15521), .ZN(n21159) );
  XNOR2_X1 U18863 ( .A(n15524), .B(n15523), .ZN(n15525) );
  NAND2_X1 U18864 ( .A1(n15526), .A2(n15525), .ZN(n15527) );
  OAI21_X1 U18865 ( .B1(n21159), .B2(n15528), .A(n15527), .ZN(n15529) );
  AOI21_X1 U18866 ( .B1(n15531), .B2(n15530), .A(n15529), .ZN(n15532) );
  NAND2_X1 U18867 ( .A1(n15533), .A2(n15532), .ZN(n21158) );
  MUX2_X1 U18868 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n21158), .S(
        n16849), .Z(n16858) );
  NAND2_X1 U18869 ( .A1(n16858), .A2(n21185), .ZN(n15535) );
  NOR2_X1 U18870 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n21185), .ZN(n15537) );
  NAND2_X1 U18871 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n15537), .ZN(
        n15534) );
  NAND2_X1 U18872 ( .A1(n15535), .A2(n15534), .ZN(n15540) );
  MUX2_X1 U18873 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15536), .S(
        n16849), .Z(n16854) );
  AOI22_X1 U18874 ( .A1(n15537), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n21185), .B2(n16854), .ZN(n15538) );
  INV_X1 U18875 ( .A(n15538), .ZN(n15539) );
  NAND2_X1 U18876 ( .A1(n15540), .A2(n15539), .ZN(n16869) );
  INV_X1 U18877 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n15541) );
  NAND2_X1 U18878 ( .A1(n15541), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n15546) );
  INV_X1 U18879 ( .A(n20644), .ZN(n20904) );
  OR2_X1 U18880 ( .A1(n15542), .A2(n20904), .ZN(n15543) );
  XNOR2_X1 U18881 ( .A(n15543), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20356) );
  NAND2_X1 U18882 ( .A1(n20356), .A2(n15544), .ZN(n16986) );
  AND2_X1 U18883 ( .A1(n16849), .A2(n21185), .ZN(n15545) );
  MUX2_X1 U18884 ( .A(n15546), .B(n16986), .S(n15545), .Z(n16871) );
  OAI21_X1 U18885 ( .B1(n16869), .B2(n13485), .A(n16871), .ZN(n15550) );
  NOR2_X1 U18886 ( .A1(n15550), .A2(n16998), .ZN(n16878) );
  INV_X1 U18887 ( .A(n16878), .ZN(n15548) );
  NAND2_X1 U18888 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20782), .ZN(n15563) );
  NAND2_X1 U18889 ( .A1(n20606), .A2(n15563), .ZN(n15547) );
  OAI211_X1 U18890 ( .C1(n20570), .C2(n21010), .A(n15548), .B(n15547), .ZN(
        n15552) );
  OAI21_X1 U18891 ( .B1(n15550), .B2(P1_FLUSH_REG_SCAN_IN), .A(n15549), .ZN(
        n15551) );
  INV_X1 U18892 ( .A(n20649), .ZN(n20497) );
  NAND2_X1 U18893 ( .A1(n15551), .A2(n20649), .ZN(n20488) );
  MUX2_X1 U18894 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15552), .S(
        n20488), .Z(P1_U3478) );
  INV_X1 U18895 ( .A(n15563), .ZN(n15557) );
  NAND2_X1 U18896 ( .A1(n15553), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20877) );
  OAI211_X1 U18897 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n15553), .A(n20877), 
        .B(n20934), .ZN(n15554) );
  OAI21_X1 U18898 ( .B1(n15557), .B2(n13484), .A(n15554), .ZN(n15555) );
  MUX2_X1 U18899 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15555), .S(
        n20488), .Z(P1_U3477) );
  INV_X1 U18900 ( .A(n15562), .ZN(n20494) );
  XNOR2_X1 U18901 ( .A(n20494), .B(n20877), .ZN(n15558) );
  OAI22_X1 U18902 ( .A1(n15558), .A2(n21010), .B1(n13452), .B2(n15557), .ZN(
        n15559) );
  MUX2_X1 U18903 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n15559), .S(
        n20488), .Z(P1_U3476) );
  NOR2_X1 U18904 ( .A1(n20750), .A2(n20877), .ZN(n20744) );
  AOI211_X1 U18905 ( .C1(n10996), .C2(n20979), .A(n20872), .B(n20744), .ZN(
        n15565) );
  OR2_X1 U18906 ( .A1(n15553), .A2(n20979), .ZN(n20806) );
  NOR2_X1 U18907 ( .A1(n20806), .A2(n21010), .ZN(n20543) );
  AND2_X1 U18908 ( .A1(n20978), .A2(n20543), .ZN(n20937) );
  AOI21_X1 U18909 ( .B1(n15563), .B2(n20774), .A(n20937), .ZN(n15564) );
  OAI21_X1 U18910 ( .B1(n15565), .B2(n21010), .A(n15564), .ZN(n15566) );
  MUX2_X1 U18911 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15566), .S(
        n20488), .Z(P1_U3475) );
  NOR2_X1 U18912 ( .A1(n20166), .A2(n20044), .ZN(n15572) );
  AOI21_X1 U18913 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n15568), .A(n15567), 
        .ZN(n15570) );
  NOR3_X1 U18914 ( .A1(n15568), .A2(n10064), .A3(n16778), .ZN(n15569) );
  OAI21_X1 U18915 ( .B1(n15570), .B2(n15569), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n15571) );
  OAI21_X1 U18916 ( .B1(n15573), .B2(n15572), .A(n15571), .ZN(n15579) );
  NAND2_X1 U18917 ( .A1(n19476), .A2(n15574), .ZN(n15575) );
  OAI211_X1 U18918 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n15577), .A(n15576), 
        .B(n15575), .ZN(n15578) );
  MUX2_X1 U18919 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n15579), .S(n15578), 
        .Z(P2_U3610) );
  INV_X1 U18920 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15584) );
  NAND2_X1 U18921 ( .A1(n15581), .A2(n19406), .ZN(n15583) );
  INV_X2 U18922 ( .A(n19404), .ZN(n16835) );
  AOI22_X1 U18923 ( .A1(n19402), .A2(P2_REIP_REG_29__SCAN_IN), .B1(n16835), 
        .B2(P2_EBX_REG_29__SCAN_IN), .ZN(n15582) );
  OAI211_X1 U18924 ( .C1(n19424), .C2(n15584), .A(n15583), .B(n15582), .ZN(
        n15585) );
  AOI21_X1 U18925 ( .B1(n15586), .B2(n19414), .A(n15585), .ZN(n15592) );
  AOI21_X1 U18926 ( .B1(n15587), .B2(n15588), .A(n16789), .ZN(n15590) );
  OAI21_X1 U18927 ( .B1(n15964), .B2(n15590), .A(n15589), .ZN(n15591) );
  OAI211_X1 U18928 ( .C1(n15936), .C2(n16068), .A(n15592), .B(n15591), .ZN(
        P2_U2826) );
  INV_X1 U18929 ( .A(n16443), .ZN(n15609) );
  NOR2_X1 U18930 ( .A1(n15597), .A2(n15596), .ZN(n15598) );
  OR2_X1 U18931 ( .A1(n12994), .A2(n15598), .ZN(n16450) );
  INV_X1 U18932 ( .A(n16450), .ZN(n15607) );
  AOI22_X1 U18933 ( .A1(n19402), .A2(P2_REIP_REG_28__SCAN_IN), .B1(n16835), 
        .B2(P2_EBX_REG_28__SCAN_IN), .ZN(n15600) );
  NAND2_X1 U18934 ( .A1(n15963), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15599) );
  OAI211_X1 U18935 ( .C1(n15601), .C2(n16838), .A(n15600), .B(n15599), .ZN(
        n15606) );
  OAI21_X1 U18936 ( .B1(n15602), .B2(n16199), .A(n19412), .ZN(n15604) );
  INV_X1 U18937 ( .A(n15587), .ZN(n15603) );
  AOI21_X1 U18938 ( .B1(n16833), .B2(n15604), .A(n15603), .ZN(n15605) );
  OAI21_X1 U18939 ( .B1(n15609), .B2(n15936), .A(n15608), .ZN(P2_U2827) );
  INV_X1 U18940 ( .A(n16081), .ZN(n15621) );
  INV_X1 U18941 ( .A(n15610), .ZN(n15627) );
  INV_X1 U18942 ( .A(n15611), .ZN(n15612) );
  OAI21_X1 U18943 ( .B1(n15627), .B2(n15612), .A(n19412), .ZN(n15613) );
  AOI21_X1 U18944 ( .B1(n16833), .B2(n15613), .A(n15602), .ZN(n15618) );
  AOI22_X1 U18945 ( .A1(n19402), .A2(P2_REIP_REG_27__SCAN_IN), .B1(n16835), 
        .B2(P2_EBX_REG_27__SCAN_IN), .ZN(n15615) );
  NAND2_X1 U18946 ( .A1(n15963), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15614) );
  OAI211_X1 U18947 ( .C1(n15616), .C2(n16838), .A(n15615), .B(n15614), .ZN(
        n15617) );
  AOI211_X1 U18948 ( .C1(n15619), .C2(n19414), .A(n15618), .B(n15617), .ZN(
        n15620) );
  OAI21_X1 U18949 ( .B1(n15621), .B2(n15936), .A(n15620), .ZN(P2_U2828) );
  NAND2_X1 U18950 ( .A1(n15640), .A2(n15622), .ZN(n15623) );
  NAND2_X1 U18951 ( .A1(n15624), .A2(n15623), .ZN(n16460) );
  AOI22_X1 U18952 ( .A1(n19402), .A2(P2_REIP_REG_26__SCAN_IN), .B1(n16835), 
        .B2(P2_EBX_REG_26__SCAN_IN), .ZN(n15625) );
  OAI21_X1 U18953 ( .B1(n19424), .B2(n15626), .A(n15625), .ZN(n15630) );
  OAI21_X1 U18954 ( .B1(n15645), .B2(n16207), .A(n19412), .ZN(n15628) );
  AOI21_X1 U18955 ( .B1(n16833), .B2(n15628), .A(n15627), .ZN(n15629) );
  AOI21_X1 U18956 ( .B1(n15633), .B2(n15632), .A(n15631), .ZN(n16463) );
  NAND2_X1 U18957 ( .A1(n16463), .A2(n13130), .ZN(n15634) );
  OAI211_X1 U18958 ( .C1(n15955), .C2(n16460), .A(n9729), .B(n15634), .ZN(
        P2_U2829) );
  XOR2_X1 U18959 ( .A(n15636), .B(n15635), .Z(n16476) );
  INV_X1 U18960 ( .A(n16476), .ZN(n16098) );
  AND2_X1 U18961 ( .A1(n15637), .A2(n15695), .ZN(n15639) );
  AND2_X1 U18962 ( .A1(n15639), .A2(n15638), .ZN(n15655) );
  OAI21_X1 U18963 ( .B1(n15655), .B2(n15641), .A(n15640), .ZN(n16473) );
  INV_X1 U18964 ( .A(n16473), .ZN(n15650) );
  NOR2_X1 U18965 ( .A1(n15642), .A2(n16838), .ZN(n15649) );
  INV_X1 U18966 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n21315) );
  NAND2_X1 U18967 ( .A1(n15661), .A2(n16216), .ZN(n15643) );
  AOI21_X1 U18968 ( .B1(n15643), .B2(n19412), .A(n15964), .ZN(n15644) );
  OR2_X1 U18969 ( .A1(n15645), .A2(n15644), .ZN(n15647) );
  AOI22_X1 U18970 ( .A1(n19402), .A2(P2_REIP_REG_25__SCAN_IN), .B1(n16835), 
        .B2(P2_EBX_REG_25__SCAN_IN), .ZN(n15646) );
  OAI211_X1 U18971 ( .C1(n19424), .C2(n21315), .A(n15647), .B(n15646), .ZN(
        n15648) );
  AOI211_X1 U18972 ( .C1(n15650), .C2(n19414), .A(n15649), .B(n15648), .ZN(
        n15651) );
  OAI21_X1 U18973 ( .B1(n16098), .B2(n15936), .A(n15651), .ZN(P2_U2830) );
  NAND2_X1 U18974 ( .A1(n15652), .A2(n15653), .ZN(n15654) );
  NAND2_X1 U18975 ( .A1(n15635), .A2(n15654), .ZN(n16489) );
  INV_X1 U18976 ( .A(n15655), .ZN(n15659) );
  NAND2_X1 U18977 ( .A1(n15637), .A2(n15695), .ZN(n16024) );
  OR2_X1 U18978 ( .A1(n16024), .A2(n15656), .ZN(n15676) );
  NAND2_X1 U18979 ( .A1(n15676), .A2(n15657), .ZN(n15658) );
  NAND2_X1 U18980 ( .A1(n15659), .A2(n15658), .ZN(n16225) );
  INV_X1 U18981 ( .A(n16225), .ZN(n16487) );
  INV_X1 U18982 ( .A(n15660), .ZN(n15678) );
  OAI21_X1 U18983 ( .B1(n15678), .B2(n16224), .A(n19412), .ZN(n15663) );
  INV_X1 U18984 ( .A(n15661), .ZN(n15662) );
  AOI21_X1 U18985 ( .B1(n16833), .B2(n15663), .A(n15662), .ZN(n15669) );
  XNOR2_X1 U18986 ( .A(n15664), .B(P2_EBX_REG_24__SCAN_IN), .ZN(n15667) );
  AOI22_X1 U18987 ( .A1(n19402), .A2(P2_REIP_REG_24__SCAN_IN), .B1(n16835), 
        .B2(P2_EBX_REG_24__SCAN_IN), .ZN(n15666) );
  NAND2_X1 U18988 ( .A1(n15963), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15665) );
  OAI211_X1 U18989 ( .C1(n15667), .C2(n16838), .A(n15666), .B(n15665), .ZN(
        n15668) );
  AOI211_X1 U18990 ( .C1(n16487), .C2(n19414), .A(n15669), .B(n15668), .ZN(
        n15670) );
  OAI21_X1 U18991 ( .B1(n16489), .B2(n15936), .A(n15670), .ZN(P2_U2831) );
  OR2_X1 U18992 ( .A1(n15671), .A2(n15672), .ZN(n15673) );
  NAND2_X1 U18993 ( .A1(n15652), .A2(n15673), .ZN(n16501) );
  OR2_X1 U18994 ( .A1(n16024), .A2(n16023), .ZN(n16026) );
  NAND2_X1 U18995 ( .A1(n16026), .A2(n15674), .ZN(n15675) );
  NAND2_X1 U18996 ( .A1(n15676), .A2(n15675), .ZN(n16020) );
  INV_X1 U18997 ( .A(n16020), .ZN(n16500) );
  INV_X1 U18998 ( .A(n16842), .ZN(n15677) );
  OAI21_X1 U18999 ( .B1(n15677), .B2(n16233), .A(n19412), .ZN(n15679) );
  AOI21_X1 U19000 ( .B1(n16833), .B2(n15679), .A(n15678), .ZN(n15684) );
  AOI22_X1 U19001 ( .A1(n19402), .A2(P2_REIP_REG_23__SCAN_IN), .B1(n16835), 
        .B2(P2_EBX_REG_23__SCAN_IN), .ZN(n15681) );
  NAND2_X1 U19002 ( .A1(n15963), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15680) );
  OAI211_X1 U19003 ( .C1(n15682), .C2(n16838), .A(n15681), .B(n15680), .ZN(
        n15683) );
  AOI211_X1 U19004 ( .C1(n16500), .C2(n19414), .A(n15684), .B(n15683), .ZN(
        n15685) );
  OAI21_X1 U19005 ( .B1(n16501), .B2(n15936), .A(n15685), .ZN(P2_U2832) );
  INV_X1 U19006 ( .A(n15687), .ZN(n15688) );
  AOI21_X1 U19007 ( .B1(n15689), .B2(n15686), .A(n15688), .ZN(n16526) );
  INV_X1 U19008 ( .A(n16526), .ZN(n15700) );
  OAI211_X1 U19009 ( .C1(n15690), .C2(n16257), .A(n15691), .B(n19412), .ZN(
        n15694) );
  AOI22_X1 U19010 ( .A1(n19402), .A2(P2_REIP_REG_21__SCAN_IN), .B1(n16835), 
        .B2(P2_EBX_REG_21__SCAN_IN), .ZN(n15693) );
  NAND2_X1 U19011 ( .A1(n15963), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15692) );
  NAND3_X1 U19012 ( .A1(n15694), .A2(n15693), .A3(n15692), .ZN(n15697) );
  OAI21_X1 U19013 ( .B1(n15637), .B2(n15695), .A(n16024), .ZN(n16524) );
  NOR2_X1 U19014 ( .A1(n16524), .A2(n15955), .ZN(n15696) );
  AOI211_X1 U19015 ( .C1(n19406), .C2(n15698), .A(n15697), .B(n15696), .ZN(
        n15699) );
  OAI21_X1 U19016 ( .B1(n15700), .B2(n15936), .A(n15699), .ZN(P2_U2834) );
  OR2_X1 U19017 ( .A1(n9639), .A2(n15701), .ZN(n15702) );
  AND2_X1 U19018 ( .A1(n15686), .A2(n15702), .ZN(n16530) );
  INV_X1 U19019 ( .A(n16530), .ZN(n15716) );
  NOR2_X1 U19020 ( .A1(n10579), .A2(n15703), .ZN(n15704) );
  OR2_X1 U19021 ( .A1(n15637), .A2(n15704), .ZN(n16542) );
  INV_X1 U19022 ( .A(n16542), .ZN(n15714) );
  INV_X1 U19023 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15706) );
  AOI22_X1 U19024 ( .A1(n19402), .A2(P2_REIP_REG_20__SCAN_IN), .B1(n16835), 
        .B2(P2_EBX_REG_20__SCAN_IN), .ZN(n15705) );
  OAI21_X1 U19025 ( .B1(n19424), .B2(n15706), .A(n15705), .ZN(n15709) );
  AOI211_X1 U19026 ( .C1(n15710), .C2(n15707), .A(n16789), .B(n15690), .ZN(
        n15708) );
  AOI211_X1 U19027 ( .C1(n15964), .C2(n15710), .A(n15709), .B(n15708), .ZN(
        n15711) );
  OAI21_X1 U19028 ( .B1(n15712), .B2(n16838), .A(n15711), .ZN(n15713) );
  AOI21_X1 U19029 ( .B1(n15714), .B2(n19414), .A(n15713), .ZN(n15715) );
  OAI21_X1 U19030 ( .B1(n15716), .B2(n15936), .A(n15715), .ZN(P2_U2835) );
  INV_X1 U19031 ( .A(n15717), .ZN(n15732) );
  AOI21_X1 U19032 ( .B1(n15718), .B2(n15732), .A(n10579), .ZN(n16281) );
  INV_X1 U19033 ( .A(n16281), .ZN(n16551) );
  NOR2_X1 U19034 ( .A1(n16750), .A2(n15719), .ZN(n15720) );
  XNOR2_X1 U19035 ( .A(n15720), .B(n16279), .ZN(n15727) );
  NAND2_X1 U19036 ( .A1(n15721), .A2(n19406), .ZN(n15724) );
  OAI21_X1 U19037 ( .B1(n15968), .B2(n20217), .A(n16394), .ZN(n15722) );
  AOI21_X1 U19038 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n16835), .A(n15722), .ZN(
        n15723) );
  OAI211_X1 U19039 ( .C1(n19424), .C2(n15725), .A(n15724), .B(n15723), .ZN(
        n15726) );
  AOI21_X1 U19040 ( .B1(n15727), .B2(n19412), .A(n15726), .ZN(n15731) );
  NOR2_X1 U19041 ( .A1(n14334), .A2(n15728), .ZN(n15744) );
  XOR2_X1 U19042 ( .A(n15729), .B(n15744), .Z(n16554) );
  NAND2_X1 U19043 ( .A1(n16554), .A2(n13130), .ZN(n15730) );
  OAI211_X1 U19044 ( .C1(n16551), .C2(n15955), .A(n15731), .B(n15730), .ZN(
        P2_U2836) );
  INV_X1 U19045 ( .A(n14331), .ZN(n15733) );
  OAI21_X1 U19046 ( .B1(n15733), .B2(n9758), .A(n15732), .ZN(n16562) );
  INV_X1 U19047 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20215) );
  OAI21_X1 U19048 ( .B1(n15968), .B2(n20215), .A(n16394), .ZN(n15734) );
  AOI21_X1 U19049 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n16835), .A(n15734), .ZN(
        n15735) );
  OAI21_X1 U19050 ( .B1(n15736), .B2(n19424), .A(n15735), .ZN(n15742) );
  NAND2_X1 U19051 ( .A1(n15738), .A2(n19412), .ZN(n15737) );
  NAND2_X1 U19052 ( .A1(n16833), .A2(n15737), .ZN(n15740) );
  NOR2_X1 U19053 ( .A1(n15975), .A2(n15738), .ZN(n15739) );
  MUX2_X1 U19054 ( .A(n15740), .B(n15739), .S(n16287), .Z(n15741) );
  AOI211_X1 U19055 ( .C1(n19406), .C2(n15743), .A(n15742), .B(n15741), .ZN(
        n15748) );
  AOI21_X1 U19056 ( .B1(n15746), .B2(n15745), .A(n15744), .ZN(n16565) );
  NAND2_X1 U19057 ( .A1(n16565), .A2(n13130), .ZN(n15747) );
  OAI211_X1 U19058 ( .C1(n15955), .C2(n16562), .A(n15748), .B(n15747), .ZN(
        P2_U2837) );
  INV_X1 U19059 ( .A(n16158), .ZN(n15761) );
  INV_X1 U19060 ( .A(n15750), .ZN(n15749) );
  NOR2_X1 U19061 ( .A1(n15975), .A2(n15749), .ZN(n15752) );
  OAI21_X1 U19062 ( .B1(n16789), .B2(n15750), .A(n16833), .ZN(n15751) );
  MUX2_X1 U19063 ( .A(n15752), .B(n15751), .S(n16297), .Z(n15759) );
  NOR2_X1 U19064 ( .A1(n16299), .A2(n15955), .ZN(n15758) );
  NOR2_X1 U19065 ( .A1(n15753), .A2(n16838), .ZN(n15757) );
  INV_X1 U19066 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16295) );
  AOI21_X1 U19067 ( .B1(n19402), .B2(P2_REIP_REG_17__SCAN_IN), .A(n16434), 
        .ZN(n15755) );
  NAND2_X1 U19068 ( .A1(n16835), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15754) );
  OAI211_X1 U19069 ( .C1(n19424), .C2(n16295), .A(n15755), .B(n15754), .ZN(
        n15756) );
  NOR4_X1 U19070 ( .A1(n15759), .A2(n15758), .A3(n15757), .A4(n15756), .ZN(
        n15760) );
  OAI21_X1 U19071 ( .B1(n15761), .B2(n15936), .A(n15760), .ZN(P2_U2838) );
  OAI21_X1 U19072 ( .B1(n14036), .B2(n15762), .A(n14334), .ZN(n16572) );
  INV_X1 U19073 ( .A(n15975), .ZN(n15905) );
  NAND2_X1 U19074 ( .A1(n15905), .A2(n15763), .ZN(n15784) );
  NOR2_X1 U19075 ( .A1(n15763), .A2(n16789), .ZN(n15764) );
  NOR2_X1 U19076 ( .A1(n15964), .A2(n15764), .ZN(n15766) );
  MUX2_X1 U19077 ( .A(n15784), .B(n15766), .S(n15765), .Z(n15775) );
  AOI21_X1 U19078 ( .B1(n15767), .B2(n14193), .A(n9673), .ZN(n16569) );
  NOR2_X1 U19079 ( .A1(n15768), .A2(n16838), .ZN(n15773) );
  INV_X1 U19080 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15771) );
  AOI21_X1 U19081 ( .B1(n19402), .B2(P2_REIP_REG_16__SCAN_IN), .A(n16434), 
        .ZN(n15770) );
  NAND2_X1 U19082 ( .A1(n16835), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n15769) );
  OAI211_X1 U19083 ( .C1(n19424), .C2(n15771), .A(n15770), .B(n15769), .ZN(
        n15772) );
  AOI211_X1 U19084 ( .C1(n16569), .C2(n19414), .A(n15773), .B(n15772), .ZN(
        n15774) );
  OAI211_X1 U19085 ( .C1(n15936), .C2(n16572), .A(n15775), .B(n15774), .ZN(
        P2_U2839) );
  INV_X1 U19086 ( .A(n16320), .ZN(n15786) );
  NAND2_X1 U19087 ( .A1(n15964), .A2(n15786), .ZN(n15782) );
  AOI21_X1 U19088 ( .B1(n19402), .B2(P2_REIP_REG_15__SCAN_IN), .A(n16434), 
        .ZN(n15777) );
  NAND2_X1 U19089 ( .A1(n16835), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n15776) );
  OAI211_X1 U19090 ( .C1(n19424), .C2(n15778), .A(n15777), .B(n15776), .ZN(
        n15779) );
  AOI21_X1 U19091 ( .B1(n15780), .B2(n19406), .A(n15779), .ZN(n15781) );
  NAND2_X1 U19092 ( .A1(n15782), .A2(n15781), .ZN(n15788) );
  INV_X1 U19093 ( .A(n15783), .ZN(n15785) );
  AOI21_X1 U19094 ( .B1(n15786), .B2(n15785), .A(n15784), .ZN(n15787) );
  AOI211_X1 U19095 ( .C1(n19414), .C2(n16583), .A(n15788), .B(n15787), .ZN(
        n15789) );
  OAI21_X1 U19096 ( .B1(n16585), .B2(n15936), .A(n15789), .ZN(P2_U2840) );
  AOI21_X1 U19097 ( .B1(n19402), .B2(P2_REIP_REG_14__SCAN_IN), .A(n16434), 
        .ZN(n15791) );
  NAND2_X1 U19098 ( .A1(n16835), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15790) );
  OAI211_X1 U19099 ( .C1(n19424), .C2(n16332), .A(n15791), .B(n15790), .ZN(
        n15792) );
  AOI21_X1 U19100 ( .B1(n15793), .B2(n19406), .A(n15792), .ZN(n15794) );
  OAI21_X1 U19101 ( .B1(n16596), .B2(n15955), .A(n15794), .ZN(n15800) );
  INV_X1 U19102 ( .A(n15796), .ZN(n15795) );
  NOR2_X1 U19103 ( .A1(n15975), .A2(n15795), .ZN(n15798) );
  OAI21_X1 U19104 ( .B1(n16789), .B2(n15796), .A(n16833), .ZN(n15797) );
  MUX2_X1 U19105 ( .A(n15798), .B(n15797), .S(n16334), .Z(n15799) );
  AOI211_X1 U19106 ( .C1(n13130), .C2(n16599), .A(n15800), .B(n15799), .ZN(
        n15801) );
  INV_X1 U19107 ( .A(n15801), .ZN(P2_U2841) );
  NAND2_X1 U19108 ( .A1(n19409), .A2(n15802), .ZN(n15803) );
  XOR2_X1 U19109 ( .A(n15803), .B(n16345), .Z(n15811) );
  AOI21_X1 U19110 ( .B1(n19402), .B2(P2_REIP_REG_13__SCAN_IN), .A(n16434), 
        .ZN(n15804) );
  OAI21_X1 U19111 ( .B1(n19404), .B2(n12446), .A(n15804), .ZN(n15805) );
  AOI21_X1 U19112 ( .B1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n15963), .A(
        n15805), .ZN(n15806) );
  OAI21_X1 U19113 ( .B1(n15807), .B2(n16838), .A(n15806), .ZN(n15808) );
  AOI21_X1 U19114 ( .B1(n16605), .B2(n19414), .A(n15808), .ZN(n15810) );
  NAND2_X1 U19115 ( .A1(n16611), .A2(n13130), .ZN(n15809) );
  OAI211_X1 U19116 ( .C1(n15811), .C2(n16789), .A(n15810), .B(n15809), .ZN(
        P2_U2842) );
  INV_X1 U19117 ( .A(n16623), .ZN(n15825) );
  INV_X1 U19118 ( .A(n15812), .ZN(n15817) );
  AOI21_X1 U19119 ( .B1(n19402), .B2(P2_REIP_REG_12__SCAN_IN), .A(n16434), 
        .ZN(n15814) );
  NAND2_X1 U19120 ( .A1(n16835), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n15813) );
  OAI211_X1 U19121 ( .C1(n19424), .C2(n15815), .A(n15814), .B(n15813), .ZN(
        n15816) );
  AOI21_X1 U19122 ( .B1(n15817), .B2(n19406), .A(n15816), .ZN(n15818) );
  OAI21_X1 U19123 ( .B1(n16619), .B2(n15955), .A(n15818), .ZN(n15824) );
  NAND2_X1 U19124 ( .A1(n15820), .A2(n19412), .ZN(n15819) );
  NAND2_X1 U19125 ( .A1(n16833), .A2(n15819), .ZN(n15822) );
  NOR2_X1 U19126 ( .A1(n15975), .A2(n15820), .ZN(n15821) );
  MUX2_X1 U19127 ( .A(n15822), .B(n15821), .S(n16356), .Z(n15823) );
  AOI211_X1 U19128 ( .C1(n13130), .C2(n15825), .A(n15824), .B(n15823), .ZN(
        n15826) );
  INV_X1 U19129 ( .A(n15826), .ZN(P2_U2843) );
  INV_X1 U19130 ( .A(n16628), .ZN(n15840) );
  INV_X1 U19131 ( .A(n12482), .ZN(n15832) );
  AOI21_X1 U19132 ( .B1(n12438), .B2(P2_EBX_REG_11__SCAN_IN), .A(n16838), .ZN(
        n15831) );
  AOI21_X1 U19133 ( .B1(n19402), .B2(P2_REIP_REG_11__SCAN_IN), .A(n16434), 
        .ZN(n15828) );
  NAND2_X1 U19134 ( .A1(n16835), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n15827) );
  OAI211_X1 U19135 ( .C1(n19424), .C2(n15829), .A(n15828), .B(n15827), .ZN(
        n15830) );
  AOI21_X1 U19136 ( .B1(n15832), .B2(n15831), .A(n15830), .ZN(n15833) );
  OAI21_X1 U19137 ( .B1(n16635), .B2(n15955), .A(n15833), .ZN(n15839) );
  NAND2_X1 U19138 ( .A1(n15835), .A2(n19412), .ZN(n15834) );
  NAND2_X1 U19139 ( .A1(n16833), .A2(n15834), .ZN(n15837) );
  NOR2_X1 U19140 ( .A1(n15975), .A2(n15835), .ZN(n15836) );
  MUX2_X1 U19141 ( .A(n15837), .B(n15836), .S(n16366), .Z(n15838) );
  AOI211_X1 U19142 ( .C1(n13130), .C2(n15840), .A(n15839), .B(n15838), .ZN(
        n15841) );
  INV_X1 U19143 ( .A(n15841), .ZN(P2_U2844) );
  INV_X1 U19144 ( .A(n16642), .ZN(n15854) );
  INV_X1 U19145 ( .A(n15842), .ZN(n15846) );
  AOI21_X1 U19146 ( .B1(n19402), .B2(P2_REIP_REG_10__SCAN_IN), .A(n16434), 
        .ZN(n15844) );
  NAND2_X1 U19147 ( .A1(n16835), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n15843) );
  OAI211_X1 U19148 ( .C1(n19424), .C2(n10379), .A(n15844), .B(n15843), .ZN(
        n15845) );
  AOI21_X1 U19149 ( .B1(n15846), .B2(n19406), .A(n15845), .ZN(n15847) );
  OAI21_X1 U19150 ( .B1(n16646), .B2(n15955), .A(n15847), .ZN(n15853) );
  INV_X1 U19151 ( .A(n15849), .ZN(n15848) );
  NOR2_X1 U19152 ( .A1(n15975), .A2(n15848), .ZN(n15851) );
  OAI21_X1 U19153 ( .B1(n16789), .B2(n15849), .A(n16833), .ZN(n15850) );
  MUX2_X1 U19154 ( .A(n15851), .B(n15850), .S(n16386), .Z(n15852) );
  AOI211_X1 U19155 ( .C1(n15854), .C2(n13130), .A(n15853), .B(n15852), .ZN(
        n15855) );
  INV_X1 U19156 ( .A(n15855), .ZN(P2_U2845) );
  NAND2_X1 U19157 ( .A1(n19409), .A2(n15856), .ZN(n15857) );
  XOR2_X1 U19158 ( .A(n15857), .B(n16395), .Z(n15865) );
  AOI21_X1 U19159 ( .B1(n19402), .B2(P2_REIP_REG_9__SCAN_IN), .A(n16434), .ZN(
        n15859) );
  NAND2_X1 U19160 ( .A1(n16835), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n15858) );
  OAI211_X1 U19161 ( .C1(n19424), .C2(n10378), .A(n15859), .B(n15858), .ZN(
        n15860) );
  AOI21_X1 U19162 ( .B1(n15861), .B2(n19406), .A(n15860), .ZN(n15862) );
  OAI21_X1 U19163 ( .B1(n16658), .B2(n15955), .A(n15862), .ZN(n15863) );
  AOI21_X1 U19164 ( .B1(n16652), .B2(n13130), .A(n15863), .ZN(n15864) );
  OAI21_X1 U19165 ( .B1(n15865), .B2(n16789), .A(n15864), .ZN(P2_U2846) );
  INV_X1 U19166 ( .A(n15866), .ZN(n15871) );
  INV_X1 U19167 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15869) );
  AOI21_X1 U19168 ( .B1(n19402), .B2(P2_REIP_REG_8__SCAN_IN), .A(n16434), .ZN(
        n15868) );
  NAND2_X1 U19169 ( .A1(n16835), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n15867) );
  OAI211_X1 U19170 ( .C1(n19424), .C2(n15869), .A(n15868), .B(n15867), .ZN(
        n15870) );
  AOI21_X1 U19171 ( .B1(n15871), .B2(n19406), .A(n15870), .ZN(n15872) );
  OAI21_X1 U19172 ( .B1(n16670), .B2(n15955), .A(n15872), .ZN(n15878) );
  NAND2_X1 U19173 ( .A1(n15874), .A2(n19412), .ZN(n15873) );
  NAND2_X1 U19174 ( .A1(n16833), .A2(n15873), .ZN(n15876) );
  NOR2_X1 U19175 ( .A1(n15975), .A2(n15874), .ZN(n15875) );
  MUX2_X1 U19176 ( .A(n15876), .B(n15875), .S(n16412), .Z(n15877) );
  AOI211_X1 U19177 ( .C1(n13130), .C2(n16672), .A(n15878), .B(n15877), .ZN(
        n15879) );
  INV_X1 U19178 ( .A(n15879), .ZN(P2_U2847) );
  INV_X1 U19179 ( .A(n19413), .ZN(n15880) );
  NOR2_X1 U19180 ( .A1(n15975), .A2(n15880), .ZN(n15882) );
  OAI21_X1 U19181 ( .B1(n16789), .B2(n19413), .A(n16833), .ZN(n15881) );
  MUX2_X1 U19182 ( .A(n15882), .B(n15881), .S(n16419), .Z(n15890) );
  AOI21_X1 U19183 ( .B1(n19402), .B2(P2_REIP_REG_7__SCAN_IN), .A(n16434), .ZN(
        n15884) );
  NAND2_X1 U19184 ( .A1(n16835), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n15883) );
  OAI211_X1 U19185 ( .C1(n19424), .C2(n21303), .A(n15884), .B(n15883), .ZN(
        n15885) );
  AOI21_X1 U19186 ( .B1(n15886), .B2(n19406), .A(n15885), .ZN(n15888) );
  NAND2_X1 U19187 ( .A1(n16685), .A2(n19414), .ZN(n15887) );
  OAI211_X1 U19188 ( .C1(n16687), .C2(n15936), .A(n15888), .B(n15887), .ZN(
        n15889) );
  OR2_X1 U19189 ( .A1(n15890), .A2(n15889), .ZN(P2_U2848) );
  NOR2_X1 U19190 ( .A1(n16750), .A2(n15891), .ZN(n15892) );
  XOR2_X1 U19191 ( .A(n15893), .B(n15892), .Z(n15904) );
  INV_X1 U19192 ( .A(n15894), .ZN(n15902) );
  NAND2_X1 U19193 ( .A1(n16835), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n15895) );
  OAI211_X1 U19194 ( .C1(n15968), .C2(n12040), .A(n16394), .B(n15895), .ZN(
        n15896) );
  AOI21_X1 U19195 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n15963), .A(
        n15896), .ZN(n15897) );
  OAI21_X1 U19196 ( .B1(n15898), .B2(n16838), .A(n15897), .ZN(n15901) );
  NOR2_X1 U19197 ( .A1(n15899), .A2(n15936), .ZN(n15900) );
  AOI211_X1 U19198 ( .C1(n15902), .C2(n19414), .A(n15901), .B(n15900), .ZN(
        n15903) );
  OAI21_X1 U19199 ( .B1(n15904), .B2(n16789), .A(n15903), .ZN(P2_U2850) );
  NAND2_X1 U19200 ( .A1(n15905), .A2(n15906), .ZN(n15910) );
  NOR2_X1 U19201 ( .A1(n15906), .A2(n16789), .ZN(n15907) );
  NOR2_X1 U19202 ( .A1(n15964), .A2(n15907), .ZN(n15909) );
  MUX2_X1 U19203 ( .A(n15910), .B(n15909), .S(n15908), .Z(n15920) );
  NAND2_X1 U19204 ( .A1(n16835), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n15911) );
  OAI211_X1 U19205 ( .C1(n15968), .C2(n20190), .A(n16394), .B(n15911), .ZN(
        n15912) );
  AOI21_X1 U19206 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n15963), .A(
        n15912), .ZN(n15913) );
  OAI21_X1 U19207 ( .B1(n15914), .B2(n16838), .A(n15913), .ZN(n15917) );
  NOR2_X1 U19208 ( .A1(n15915), .A2(n15936), .ZN(n15916) );
  AOI211_X1 U19209 ( .C1(n15918), .C2(n19414), .A(n15917), .B(n15916), .ZN(
        n15919) );
  OAI211_X1 U19210 ( .C1(n15921), .C2(n15969), .A(n15920), .B(n15919), .ZN(
        P2_U2851) );
  OAI21_X1 U19211 ( .B1(n16789), .B2(n15922), .A(n16833), .ZN(n15926) );
  INV_X1 U19212 ( .A(n15922), .ZN(n15923) );
  NOR2_X1 U19213 ( .A1(n15975), .A2(n15923), .ZN(n15925) );
  MUX2_X1 U19214 ( .A(n15926), .B(n15925), .S(n15924), .Z(n15939) );
  OR2_X1 U19215 ( .A1(n19598), .A2(n15969), .ZN(n15935) );
  INV_X1 U19216 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15931) );
  AOI22_X1 U19217 ( .A1(n19402), .A2(P2_REIP_REG_3__SCAN_IN), .B1(n16835), 
        .B2(P2_EBX_REG_3__SCAN_IN), .ZN(n15930) );
  INV_X1 U19218 ( .A(n15927), .ZN(n15928) );
  NAND2_X1 U19219 ( .A1(n15928), .A2(n19406), .ZN(n15929) );
  OAI211_X1 U19220 ( .C1(n19424), .C2(n15931), .A(n15930), .B(n15929), .ZN(
        n15932) );
  AOI21_X1 U19221 ( .B1(n15933), .B2(n19414), .A(n15932), .ZN(n15934) );
  OAI211_X1 U19222 ( .C1(n15937), .C2(n15936), .A(n15935), .B(n15934), .ZN(
        n15938) );
  OR2_X1 U19223 ( .A1(n15939), .A2(n15938), .ZN(P2_U2852) );
  XOR2_X1 U19224 ( .A(n15950), .B(n15941), .Z(n15942) );
  NAND2_X1 U19225 ( .A1(n15942), .A2(n19412), .ZN(n15949) );
  NAND2_X1 U19226 ( .A1(n15963), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n15944) );
  AOI22_X1 U19227 ( .A1(n19402), .A2(P2_REIP_REG_2__SCAN_IN), .B1(n16835), 
        .B2(P2_EBX_REG_2__SCAN_IN), .ZN(n15943) );
  OAI211_X1 U19228 ( .C1(n15945), .C2(n16838), .A(n15944), .B(n15943), .ZN(
        n15947) );
  AOI211_X1 U19229 ( .C1(n13130), .C2(n20268), .A(n15947), .B(n15946), .ZN(
        n15948) );
  OAI211_X1 U19230 ( .C1(n15969), .C2(n20264), .A(n15949), .B(n15948), .ZN(
        P2_U2853) );
  AOI21_X1 U19231 ( .B1(n16740), .B2(n15951), .A(n15950), .ZN(n16749) );
  INV_X1 U19232 ( .A(n16749), .ZN(n15962) );
  AOI22_X1 U19233 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19402), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n15963), .ZN(n15953) );
  NAND2_X1 U19234 ( .A1(n16835), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n15952) );
  OAI211_X1 U19235 ( .C1(n16838), .C2(n15954), .A(n15953), .B(n15952), .ZN(
        n15957) );
  AOI211_X1 U19236 ( .C1(n13130), .C2(n19432), .A(n15957), .B(n15956), .ZN(
        n15958) );
  OAI21_X1 U19237 ( .B1(n19523), .B2(n15969), .A(n15958), .ZN(n15959) );
  AOI21_X1 U19238 ( .B1(n15964), .B2(n15960), .A(n15959), .ZN(n15961) );
  OAI21_X1 U19239 ( .B1(n15962), .B2(n16789), .A(n15961), .ZN(P2_U2854) );
  INV_X1 U19240 ( .A(n16740), .ZN(n15974) );
  OAI21_X1 U19241 ( .B1(n15964), .B2(n15963), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15973) );
  AOI22_X1 U19242 ( .A1(n13130), .A2(n16725), .B1(n19406), .B2(n15965), .ZN(
        n15967) );
  NAND2_X1 U19243 ( .A1(n16835), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n15966) );
  OAI211_X1 U19244 ( .C1(n15968), .C2(n19395), .A(n15967), .B(n15966), .ZN(
        n15971) );
  NOR2_X1 U19245 ( .A1(n19522), .A2(n15969), .ZN(n15970) );
  AOI211_X1 U19246 ( .C1(n19414), .C2(n9836), .A(n15971), .B(n15970), .ZN(
        n15972) );
  OAI211_X1 U19247 ( .C1(n15975), .C2(n15974), .A(n15973), .B(n15972), .ZN(
        P2_U2855) );
  MUX2_X1 U19248 ( .A(n15976), .B(P2_EBX_REG_31__SCAN_IN), .S(n9598), .Z(
        P2_U2856) );
  NAND3_X1 U19249 ( .A1(n16062), .A2(n15978), .A3(n16036), .ZN(n15980) );
  NAND2_X1 U19250 ( .A1(n9598), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15979) );
  OAI211_X1 U19251 ( .C1(n9598), .C2(n16185), .A(n15980), .B(n15979), .ZN(
        P2_U2858) );
  NOR2_X1 U19252 ( .A1(n15981), .A2(n15982), .ZN(n15984) );
  XNOR2_X1 U19253 ( .A(n15984), .B(n15983), .ZN(n16075) );
  NOR2_X1 U19254 ( .A1(n16450), .A2(n9598), .ZN(n15985) );
  AOI21_X1 U19255 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n9598), .A(n15985), .ZN(
        n15986) );
  OAI21_X1 U19256 ( .B1(n16075), .B2(n16061), .A(n15986), .ZN(P2_U2859) );
  OAI21_X1 U19257 ( .B1(n15989), .B2(n15988), .A(n15987), .ZN(n16083) );
  NOR2_X1 U19258 ( .A1(n15990), .A2(n9598), .ZN(n15991) );
  AOI21_X1 U19259 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n9598), .A(n15991), .ZN(
        n15992) );
  OAI21_X1 U19260 ( .B1(n16083), .B2(n16061), .A(n15992), .ZN(P2_U2860) );
  NOR2_X1 U19261 ( .A1(n16003), .A2(n16002), .ZN(n16001) );
  NOR2_X1 U19262 ( .A1(n16001), .A2(n15993), .ZN(n15998) );
  XNOR2_X1 U19263 ( .A(n15996), .B(n15995), .ZN(n15997) );
  XNOR2_X1 U19264 ( .A(n15998), .B(n15997), .ZN(n16090) );
  MUX2_X1 U19265 ( .A(n16460), .B(n15999), .S(n9598), .Z(n16000) );
  OAI21_X1 U19266 ( .B1(n16090), .B2(n16061), .A(n16000), .ZN(P2_U2861) );
  AOI21_X1 U19267 ( .B1(n16003), .B2(n16002), .A(n16001), .ZN(n16091) );
  NAND2_X1 U19268 ( .A1(n16091), .A2(n16036), .ZN(n16005) );
  NAND2_X1 U19269 ( .A1(n9598), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n16004) );
  OAI211_X1 U19270 ( .C1(n16473), .C2(n9598), .A(n16005), .B(n16004), .ZN(
        P2_U2862) );
  INV_X1 U19271 ( .A(n16009), .ZN(n16006) );
  XNOR2_X1 U19272 ( .A(n16030), .B(n16006), .ZN(n16017) );
  INV_X1 U19273 ( .A(n16007), .ZN(n16008) );
  AOI21_X1 U19274 ( .B1(n16030), .B2(n16009), .A(n16019), .ZN(n16013) );
  XNOR2_X1 U19275 ( .A(n16011), .B(n16010), .ZN(n16012) );
  XNOR2_X1 U19276 ( .A(n16013), .B(n16012), .ZN(n16104) );
  NOR2_X1 U19277 ( .A1(n16225), .A2(n9598), .ZN(n16014) );
  AOI21_X1 U19278 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n9598), .A(n16014), .ZN(
        n16015) );
  OAI21_X1 U19279 ( .B1(n16104), .B2(n16061), .A(n16015), .ZN(P2_U2863) );
  NOR2_X1 U19280 ( .A1(n16017), .A2(n16016), .ZN(n16018) );
  NOR2_X1 U19281 ( .A1(n16020), .A2(n9598), .ZN(n16021) );
  AOI21_X1 U19282 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n9598), .A(n16021), .ZN(
        n16022) );
  OAI21_X1 U19283 ( .B1(n16061), .B2(n16110), .A(n16022), .ZN(P2_U2864) );
  NAND2_X1 U19284 ( .A1(n16024), .A2(n16023), .ZN(n16025) );
  NAND2_X1 U19285 ( .A1(n16026), .A2(n16025), .ZN(n16827) );
  AND2_X1 U19286 ( .A1(n16027), .A2(n16028), .ZN(n16029) );
  NOR2_X1 U19287 ( .A1(n16030), .A2(n16029), .ZN(n16111) );
  NAND2_X1 U19288 ( .A1(n16111), .A2(n16036), .ZN(n16032) );
  NAND2_X1 U19289 ( .A1(n9598), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n16031) );
  OAI211_X1 U19290 ( .C1(n16827), .C2(n9598), .A(n16032), .B(n16031), .ZN(
        P2_U2865) );
  INV_X1 U19291 ( .A(n16027), .ZN(n16034) );
  AOI21_X1 U19292 ( .B1(n16035), .B2(n16033), .A(n16034), .ZN(n16120) );
  NAND2_X1 U19293 ( .A1(n16120), .A2(n16036), .ZN(n16038) );
  NAND2_X1 U19294 ( .A1(n9598), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n16037) );
  OAI211_X1 U19295 ( .C1(n16524), .C2(n9598), .A(n16038), .B(n16037), .ZN(
        P2_U2866) );
  OAI21_X1 U19296 ( .B1(n16039), .B2(n16040), .A(n16033), .ZN(n16132) );
  NOR2_X1 U19297 ( .A1(n16542), .A2(n9598), .ZN(n16041) );
  AOI21_X1 U19298 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n9598), .A(n16041), .ZN(
        n16042) );
  OAI21_X1 U19299 ( .B1(n16061), .B2(n16132), .A(n16042), .ZN(P2_U2867) );
  NOR2_X1 U19300 ( .A1(n16043), .A2(n16044), .ZN(n16045) );
  OR2_X1 U19301 ( .A1(n16039), .A2(n16045), .ZN(n16144) );
  NOR2_X1 U19302 ( .A1(n16551), .A2(n9598), .ZN(n16046) );
  AOI21_X1 U19303 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n9598), .A(n16046), .ZN(
        n16047) );
  OAI21_X1 U19304 ( .B1(n16061), .B2(n16144), .A(n16047), .ZN(P2_U2868) );
  AND2_X1 U19305 ( .A1(n16048), .A2(n16049), .ZN(n16050) );
  OR2_X1 U19306 ( .A1(n16050), .A2(n16043), .ZN(n16150) );
  NOR2_X1 U19307 ( .A1(n16562), .A2(n9598), .ZN(n16051) );
  AOI21_X1 U19308 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n9598), .A(n16051), .ZN(
        n16052) );
  OAI21_X1 U19309 ( .B1(n16061), .B2(n16150), .A(n16052), .ZN(P2_U2869) );
  OAI21_X1 U19310 ( .B1(n16053), .B2(n10578), .A(n16048), .ZN(n16160) );
  NOR2_X1 U19311 ( .A1(n16299), .A2(n9598), .ZN(n16054) );
  AOI21_X1 U19312 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n9598), .A(n16054), .ZN(
        n16055) );
  OAI21_X1 U19313 ( .B1(n16061), .B2(n16160), .A(n16055), .ZN(P2_U2870) );
  OAI21_X1 U19314 ( .B1(n14380), .B2(n16057), .A(n16056), .ZN(n16170) );
  NAND2_X1 U19315 ( .A1(n16569), .A2(n16058), .ZN(n16060) );
  NAND2_X1 U19316 ( .A1(n9598), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n16059) );
  OAI211_X1 U19317 ( .C1(n16170), .C2(n16061), .A(n16060), .B(n16059), .ZN(
        P2_U2871) );
  NAND2_X1 U19318 ( .A1(n16162), .A2(BUF1_REG_29__SCAN_IN), .ZN(n16066) );
  NAND2_X1 U19319 ( .A1(n16168), .A2(BUF2_REG_29__SCAN_IN), .ZN(n16065) );
  INV_X1 U19320 ( .A(n19516), .ZN(n16063) );
  AOI22_X1 U19321 ( .A1(n16161), .A2(n16063), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n19431), .ZN(n16064) );
  AND3_X1 U19322 ( .A1(n16066), .A2(n16065), .A3(n16064), .ZN(n16067) );
  NAND2_X1 U19323 ( .A1(n16168), .A2(BUF2_REG_28__SCAN_IN), .ZN(n16072) );
  NAND2_X1 U19324 ( .A1(n16162), .A2(BUF1_REG_28__SCAN_IN), .ZN(n16071) );
  INV_X1 U19325 ( .A(n19514), .ZN(n16069) );
  AOI22_X1 U19326 ( .A1(n16161), .A2(n16069), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n19431), .ZN(n16070) );
  NAND3_X1 U19327 ( .A1(n16072), .A2(n16071), .A3(n16070), .ZN(n16073) );
  AOI21_X1 U19328 ( .B1(n16443), .B2(n19433), .A(n16073), .ZN(n16074) );
  OAI21_X1 U19329 ( .B1(n16075), .B2(n16171), .A(n16074), .ZN(P2_U2891) );
  NAND2_X1 U19330 ( .A1(n16168), .A2(BUF2_REG_27__SCAN_IN), .ZN(n16079) );
  NAND2_X1 U19331 ( .A1(n16162), .A2(BUF1_REG_27__SCAN_IN), .ZN(n16078) );
  INV_X1 U19332 ( .A(n19512), .ZN(n16076) );
  AOI22_X1 U19333 ( .A1(n16161), .A2(n16076), .B1(P2_EAX_REG_27__SCAN_IN), 
        .B2(n19431), .ZN(n16077) );
  NAND3_X1 U19334 ( .A1(n16079), .A2(n16078), .A3(n16077), .ZN(n16080) );
  AOI21_X1 U19335 ( .B1(n16081), .B2(n19433), .A(n16080), .ZN(n16082) );
  OAI21_X1 U19336 ( .B1(n16083), .B2(n16171), .A(n16082), .ZN(P2_U2892) );
  NAND2_X1 U19337 ( .A1(n16162), .A2(BUF1_REG_26__SCAN_IN), .ZN(n16087) );
  NAND2_X1 U19338 ( .A1(n16168), .A2(BUF2_REG_26__SCAN_IN), .ZN(n16086) );
  AOI22_X1 U19339 ( .A1(n16161), .A2(n16084), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n19431), .ZN(n16085) );
  NAND3_X1 U19340 ( .A1(n16087), .A2(n16086), .A3(n16085), .ZN(n16088) );
  AOI21_X1 U19341 ( .B1(n16463), .B2(n19433), .A(n16088), .ZN(n16089) );
  OAI21_X1 U19342 ( .B1(n16090), .B2(n16171), .A(n16089), .ZN(P2_U2893) );
  NAND2_X1 U19343 ( .A1(n16091), .A2(n19437), .ZN(n16097) );
  NAND2_X1 U19344 ( .A1(n16162), .A2(BUF1_REG_25__SCAN_IN), .ZN(n16095) );
  NAND2_X1 U19345 ( .A1(n16168), .A2(BUF2_REG_25__SCAN_IN), .ZN(n16094) );
  AOI22_X1 U19346 ( .A1(n16161), .A2(n16092), .B1(P2_EAX_REG_25__SCAN_IN), 
        .B2(n19431), .ZN(n16093) );
  AND3_X1 U19347 ( .A1(n16095), .A2(n16094), .A3(n16093), .ZN(n16096) );
  OAI211_X1 U19348 ( .C1(n16098), .C2(n16165), .A(n16097), .B(n16096), .ZN(
        P2_U2894) );
  AOI22_X1 U19349 ( .A1(n16161), .A2(n19488), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n19431), .ZN(n16100) );
  NAND2_X1 U19350 ( .A1(n16162), .A2(BUF1_REG_24__SCAN_IN), .ZN(n16099) );
  NAND2_X1 U19351 ( .A1(n16100), .A2(n16099), .ZN(n16102) );
  NOR2_X1 U19352 ( .A1(n16489), .A2(n16165), .ZN(n16101) );
  AOI211_X1 U19353 ( .C1(n16168), .C2(BUF2_REG_24__SCAN_IN), .A(n16102), .B(
        n16101), .ZN(n16103) );
  OAI21_X1 U19354 ( .B1(n16104), .B2(n16171), .A(n16103), .ZN(P2_U2895) );
  INV_X1 U19355 ( .A(n19508), .ZN(n19581) );
  AOI22_X1 U19356 ( .A1(n16161), .A2(n19581), .B1(P2_EAX_REG_23__SCAN_IN), 
        .B2(n19431), .ZN(n16106) );
  NAND2_X1 U19357 ( .A1(n16162), .A2(BUF1_REG_23__SCAN_IN), .ZN(n16105) );
  NAND2_X1 U19358 ( .A1(n16106), .A2(n16105), .ZN(n16108) );
  NOR2_X1 U19359 ( .A1(n16501), .A2(n16165), .ZN(n16107) );
  AOI211_X1 U19360 ( .C1(n16168), .C2(BUF2_REG_23__SCAN_IN), .A(n16108), .B(
        n16107), .ZN(n16109) );
  OAI21_X1 U19361 ( .B1(n16171), .B2(n16110), .A(n16109), .ZN(P2_U2896) );
  INV_X1 U19362 ( .A(n16111), .ZN(n16119) );
  AND2_X1 U19363 ( .A1(n15687), .A2(n16112), .ZN(n16113) );
  OR2_X1 U19364 ( .A1(n16113), .A2(n15671), .ZN(n16508) );
  INV_X1 U19365 ( .A(n16508), .ZN(n16829) );
  NAND2_X1 U19366 ( .A1(n16168), .A2(BUF2_REG_22__SCAN_IN), .ZN(n16116) );
  NAND2_X1 U19367 ( .A1(n16162), .A2(BUF1_REG_22__SCAN_IN), .ZN(n16115) );
  INV_X1 U19368 ( .A(n19506), .ZN(n19568) );
  AOI22_X1 U19369 ( .A1(n16161), .A2(n19568), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19431), .ZN(n16114) );
  NAND3_X1 U19370 ( .A1(n16116), .A2(n16115), .A3(n16114), .ZN(n16117) );
  AOI21_X1 U19371 ( .B1(n16829), .B2(n19433), .A(n16117), .ZN(n16118) );
  OAI21_X1 U19372 ( .B1(n16171), .B2(n16119), .A(n16118), .ZN(P2_U2897) );
  INV_X1 U19373 ( .A(n16120), .ZN(n16126) );
  NAND2_X1 U19374 ( .A1(n16168), .A2(BUF2_REG_21__SCAN_IN), .ZN(n16123) );
  NAND2_X1 U19375 ( .A1(n16162), .A2(BUF1_REG_21__SCAN_IN), .ZN(n16122) );
  AOI22_X1 U19376 ( .A1(n16161), .A2(n19561), .B1(P2_EAX_REG_21__SCAN_IN), 
        .B2(n19431), .ZN(n16121) );
  NAND3_X1 U19377 ( .A1(n16123), .A2(n16122), .A3(n16121), .ZN(n16124) );
  AOI21_X1 U19378 ( .B1(n16526), .B2(n19433), .A(n16124), .ZN(n16125) );
  OAI21_X1 U19379 ( .B1(n16171), .B2(n16126), .A(n16125), .ZN(P2_U2898) );
  NAND2_X1 U19380 ( .A1(n16168), .A2(BUF2_REG_20__SCAN_IN), .ZN(n16129) );
  NAND2_X1 U19381 ( .A1(n16162), .A2(BUF1_REG_20__SCAN_IN), .ZN(n16128) );
  AOI22_X1 U19382 ( .A1(n16161), .A2(n19555), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19431), .ZN(n16127) );
  NAND3_X1 U19383 ( .A1(n16129), .A2(n16128), .A3(n16127), .ZN(n16130) );
  AOI21_X1 U19384 ( .B1(n16530), .B2(n19433), .A(n16130), .ZN(n16131) );
  OAI21_X1 U19385 ( .B1(n16171), .B2(n16132), .A(n16131), .ZN(P2_U2899) );
  NAND2_X1 U19386 ( .A1(n16554), .A2(n19433), .ZN(n16143) );
  INV_X1 U19387 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16133) );
  OR2_X1 U19388 ( .A1(n14365), .A2(n16133), .ZN(n16135) );
  NAND2_X1 U19389 ( .A1(n14365), .A2(BUF2_REG_3__SCAN_IN), .ZN(n16134) );
  AND2_X1 U19390 ( .A1(n16135), .A2(n16134), .ZN(n19547) );
  OAI22_X1 U19391 ( .A1(n19547), .A2(n16138), .B1(n16137), .B2(n16136), .ZN(
        n16141) );
  INV_X1 U19392 ( .A(n16168), .ZN(n16139) );
  NOR2_X1 U19393 ( .A1(n16139), .A2(n18738), .ZN(n16140) );
  AOI211_X1 U19394 ( .C1(BUF1_REG_19__SCAN_IN), .C2(n16162), .A(n16141), .B(
        n16140), .ZN(n16142) );
  OAI211_X1 U19395 ( .C1(n16171), .C2(n16144), .A(n16143), .B(n16142), .ZN(
        P2_U2900) );
  NAND2_X1 U19396 ( .A1(n16168), .A2(BUF2_REG_18__SCAN_IN), .ZN(n16147) );
  NAND2_X1 U19397 ( .A1(n16162), .A2(BUF1_REG_18__SCAN_IN), .ZN(n16146) );
  INV_X1 U19398 ( .A(n19499), .ZN(n19542) );
  AOI22_X1 U19399 ( .A1(n16161), .A2(n19542), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19431), .ZN(n16145) );
  NAND3_X1 U19400 ( .A1(n16147), .A2(n16146), .A3(n16145), .ZN(n16148) );
  AOI21_X1 U19401 ( .B1(n16565), .B2(n19433), .A(n16148), .ZN(n16149) );
  OAI21_X1 U19402 ( .B1(n16171), .B2(n16150), .A(n16149), .ZN(P2_U2901) );
  NAND2_X1 U19403 ( .A1(n16168), .A2(BUF2_REG_17__SCAN_IN), .ZN(n16156) );
  NAND2_X1 U19404 ( .A1(n16162), .A2(BUF1_REG_17__SCAN_IN), .ZN(n16155) );
  INV_X1 U19405 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16151) );
  OR2_X1 U19406 ( .A1(n14365), .A2(n16151), .ZN(n16153) );
  NAND2_X1 U19407 ( .A1(n14365), .A2(BUF2_REG_1__SCAN_IN), .ZN(n16152) );
  INV_X1 U19408 ( .A(n19497), .ZN(n19538) );
  AOI22_X1 U19409 ( .A1(n16161), .A2(n19538), .B1(P2_EAX_REG_17__SCAN_IN), 
        .B2(n19431), .ZN(n16154) );
  NAND3_X1 U19410 ( .A1(n16156), .A2(n16155), .A3(n16154), .ZN(n16157) );
  AOI21_X1 U19411 ( .B1(n16158), .B2(n19433), .A(n16157), .ZN(n16159) );
  OAI21_X1 U19412 ( .B1(n16171), .B2(n16160), .A(n16159), .ZN(P2_U2902) );
  INV_X1 U19413 ( .A(n19495), .ZN(n16777) );
  AOI22_X1 U19414 ( .A1(n16161), .A2(n16777), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19431), .ZN(n16164) );
  NAND2_X1 U19415 ( .A1(n16162), .A2(BUF1_REG_16__SCAN_IN), .ZN(n16163) );
  NAND2_X1 U19416 ( .A1(n16164), .A2(n16163), .ZN(n16167) );
  NOR2_X1 U19417 ( .A1(n16572), .A2(n16165), .ZN(n16166) );
  AOI211_X1 U19418 ( .C1(n16168), .C2(BUF2_REG_16__SCAN_IN), .A(n16167), .B(
        n16166), .ZN(n16169) );
  OAI21_X1 U19419 ( .B1(n16171), .B2(n16170), .A(n16169), .ZN(P2_U2903) );
  OAI21_X1 U19420 ( .B1(n16436), .B2(n16173), .A(n16172), .ZN(n16174) );
  AOI21_X1 U19421 ( .B1(n16175), .B2(n16433), .A(n16174), .ZN(n16176) );
  OAI21_X1 U19422 ( .B1(n16177), .B2(n16409), .A(n16176), .ZN(n16178) );
  AOI21_X1 U19423 ( .B1(n16179), .B2(n16426), .A(n16178), .ZN(n16180) );
  OAI21_X1 U19424 ( .B1(n16181), .B2(n16429), .A(n16180), .ZN(P2_U2984) );
  NAND2_X1 U19425 ( .A1(n16410), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16182) );
  OAI211_X1 U19426 ( .C1(n16184), .C2(n16413), .A(n16183), .B(n16182), .ZN(
        n16187) );
  NOR2_X1 U19427 ( .A1(n16185), .A2(n16409), .ZN(n16186) );
  AOI211_X1 U19428 ( .C1(n16426), .C2(n16188), .A(n16187), .B(n16186), .ZN(
        n16189) );
  OAI21_X1 U19429 ( .B1(n16190), .B2(n16429), .A(n16189), .ZN(P2_U2985) );
  INV_X1 U19430 ( .A(n16192), .ZN(n16193) );
  NAND2_X1 U19431 ( .A1(n16194), .A2(n16193), .ZN(n16195) );
  XNOR2_X1 U19432 ( .A(n16196), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16197) );
  NAND2_X1 U19433 ( .A1(n16434), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n16444) );
  NAND2_X1 U19434 ( .A1(n16410), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16198) );
  OAI211_X1 U19435 ( .C1(n16199), .C2(n16413), .A(n16444), .B(n16198), .ZN(
        n16200) );
  OAI21_X1 U19436 ( .B1(n16453), .B2(n16429), .A(n16201), .ZN(P2_U2986) );
  INV_X1 U19437 ( .A(n16222), .ZN(n16204) );
  NAND2_X1 U19438 ( .A1(n16222), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16203) );
  NOR2_X1 U19439 ( .A1(n16460), .A2(n16409), .ZN(n16209) );
  NAND2_X1 U19440 ( .A1(n16434), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n16458) );
  NAND2_X1 U19441 ( .A1(n16410), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16206) );
  OAI211_X1 U19442 ( .C1(n16207), .C2(n16413), .A(n16458), .B(n16206), .ZN(
        n16208) );
  NAND2_X1 U19443 ( .A1(n16211), .A2(n16210), .ZN(n16212) );
  XOR2_X1 U19444 ( .A(n16212), .B(n9723), .Z(n16479) );
  NAND2_X1 U19445 ( .A1(n16213), .A2(n16471), .ZN(n16467) );
  NAND3_X1 U19446 ( .A1(n10512), .A2(n16383), .A3(n16467), .ZN(n16218) );
  NAND2_X1 U19447 ( .A1(n16434), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n16470) );
  OAI21_X1 U19448 ( .B1(n16436), .B2(n21315), .A(n16470), .ZN(n16215) );
  NOR2_X1 U19449 ( .A1(n16473), .A2(n16409), .ZN(n16214) );
  AOI211_X1 U19450 ( .C1(n16433), .C2(n16216), .A(n16215), .B(n16214), .ZN(
        n16217) );
  OAI211_X1 U19451 ( .C1(n16439), .C2(n16479), .A(n16218), .B(n16217), .ZN(
        P2_U2989) );
  OAI21_X1 U19452 ( .B1(n9952), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16213), .ZN(n16480) );
  XNOR2_X1 U19453 ( .A(n16220), .B(n16484), .ZN(n16221) );
  XNOR2_X1 U19454 ( .A(n16222), .B(n16221), .ZN(n16488) );
  NAND2_X1 U19455 ( .A1(n16434), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n16482) );
  NAND2_X1 U19456 ( .A1(n16410), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16223) );
  OAI211_X1 U19457 ( .C1(n16224), .C2(n16413), .A(n16482), .B(n16223), .ZN(
        n16227) );
  NOR2_X1 U19458 ( .A1(n16225), .A2(n16409), .ZN(n16226) );
  AOI211_X1 U19459 ( .C1(n16426), .C2(n16488), .A(n16227), .B(n16226), .ZN(
        n16228) );
  OAI21_X1 U19460 ( .B1(n16480), .B2(n16429), .A(n16228), .ZN(P2_U2990) );
  XNOR2_X1 U19461 ( .A(n16229), .B(n16230), .ZN(n16504) );
  AOI21_X1 U19462 ( .B1(n16498), .B2(n16231), .A(n9952), .ZN(n16506) );
  NAND2_X1 U19463 ( .A1(n16506), .A2(n16383), .ZN(n16236) );
  NAND2_X1 U19464 ( .A1(n16434), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n16497) );
  NAND2_X1 U19465 ( .A1(n16410), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16232) );
  OAI211_X1 U19466 ( .C1(n16233), .C2(n16413), .A(n16497), .B(n16232), .ZN(
        n16234) );
  AOI21_X1 U19467 ( .B1(n16500), .B2(n10023), .A(n16234), .ZN(n16235) );
  OAI211_X1 U19468 ( .C1(n16504), .C2(n16439), .A(n16236), .B(n16235), .ZN(
        P2_U2991) );
  NAND2_X1 U19469 ( .A1(n16239), .A2(n16238), .ZN(n16240) );
  XNOR2_X1 U19470 ( .A(n16241), .B(n16240), .ZN(n16515) );
  NAND2_X1 U19471 ( .A1(n16434), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n16512) );
  NAND2_X1 U19472 ( .A1(n16410), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16242) );
  OAI211_X1 U19473 ( .C1(n16830), .C2(n16413), .A(n16512), .B(n16242), .ZN(
        n16244) );
  NOR2_X1 U19474 ( .A1(n16827), .A2(n16409), .ZN(n16243) );
  AOI211_X1 U19475 ( .C1(n16426), .C2(n16515), .A(n16244), .B(n16243), .ZN(
        n16245) );
  OAI21_X1 U19476 ( .B1(n16518), .B2(n16429), .A(n16245), .ZN(P2_U2992) );
  INV_X1 U19477 ( .A(n16263), .ZN(n16249) );
  NAND2_X1 U19478 ( .A1(n16252), .A2(n16251), .ZN(n16253) );
  XNOR2_X1 U19479 ( .A(n16254), .B(n16253), .ZN(n16529) );
  NOR2_X1 U19480 ( .A1(n16524), .A2(n16409), .ZN(n16259) );
  NAND2_X1 U19481 ( .A1(n16434), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n16523) );
  NAND2_X1 U19482 ( .A1(n16410), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16256) );
  OAI211_X1 U19483 ( .C1(n16257), .C2(n16413), .A(n16523), .B(n16256), .ZN(
        n16258) );
  OAI21_X1 U19484 ( .B1(n16529), .B2(n16439), .A(n16260), .ZN(P2_U2993) );
  NAND2_X1 U19485 ( .A1(n16262), .A2(n16261), .ZN(n16266) );
  NAND2_X1 U19486 ( .A1(n16264), .A2(n16263), .ZN(n16265) );
  XNOR2_X1 U19487 ( .A(n16266), .B(n16265), .ZN(n16546) );
  INV_X1 U19488 ( .A(n16534), .ZN(n16536) );
  OAI21_X1 U19489 ( .B1(n16290), .B2(n16532), .A(n16535), .ZN(n16268) );
  NOR2_X1 U19490 ( .A1(n16542), .A2(n16409), .ZN(n16272) );
  NAND2_X1 U19491 ( .A1(n16434), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n16538) );
  NAND2_X1 U19492 ( .A1(n16410), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16269) );
  OAI211_X1 U19493 ( .C1(n16270), .C2(n16413), .A(n16538), .B(n16269), .ZN(
        n16271) );
  AOI211_X1 U19494 ( .C1(n16544), .C2(n16383), .A(n16272), .B(n16271), .ZN(
        n16273) );
  OAI21_X1 U19495 ( .B1(n16546), .B2(n16439), .A(n16273), .ZN(P2_U2994) );
  NAND2_X1 U19496 ( .A1(n16275), .A2(n16274), .ZN(n16277) );
  NAND2_X1 U19497 ( .A1(n16434), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n16547) );
  NAND2_X1 U19498 ( .A1(n16410), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16278) );
  OAI211_X1 U19499 ( .C1(n16279), .C2(n16413), .A(n16547), .B(n16278), .ZN(
        n16280) );
  OAI21_X1 U19500 ( .B1(n16556), .B2(n16439), .A(n16282), .ZN(P2_U2995) );
  NAND2_X1 U19501 ( .A1(n16276), .A2(n16283), .ZN(n16284) );
  XNOR2_X1 U19502 ( .A(n16285), .B(n16284), .ZN(n16566) );
  INV_X1 U19503 ( .A(n16562), .ZN(n16292) );
  AND2_X1 U19504 ( .A1(n16434), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n16559) );
  AOI21_X1 U19505 ( .B1(n16410), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16559), .ZN(n16286) );
  OAI21_X1 U19506 ( .B1(n16287), .B2(n16413), .A(n16286), .ZN(n16291) );
  OAI21_X1 U19507 ( .B1(n16566), .B2(n16439), .A(n16293), .ZN(P2_U2996) );
  OAI21_X1 U19508 ( .B1(n16436), .B2(n16295), .A(n16294), .ZN(n16296) );
  AOI21_X1 U19509 ( .B1(n16297), .B2(n16433), .A(n16296), .ZN(n16298) );
  OAI21_X1 U19510 ( .B1(n16299), .B2(n16409), .A(n16298), .ZN(n16303) );
  AOI211_X1 U19511 ( .C1(n16309), .C2(n16301), .A(n16300), .B(n16429), .ZN(
        n16302) );
  AOI211_X1 U19512 ( .C1(n16426), .C2(n16304), .A(n16303), .B(n16302), .ZN(
        n16305) );
  INV_X1 U19513 ( .A(n16305), .ZN(P2_U2997) );
  OAI21_X1 U19514 ( .B1(n16308), .B2(n16307), .A(n16306), .ZN(n16568) );
  OAI211_X1 U19515 ( .C1(n16310), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n16309), .B(n16383), .ZN(n16315) );
  NAND2_X1 U19516 ( .A1(n16434), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n16570) );
  NAND2_X1 U19517 ( .A1(n16410), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16311) );
  OAI211_X1 U19518 ( .C1(n16413), .C2(n16312), .A(n16570), .B(n16311), .ZN(
        n16313) );
  AOI21_X1 U19519 ( .B1(n16569), .B2(n10023), .A(n16313), .ZN(n16314) );
  OAI211_X1 U19520 ( .C1(n16568), .C2(n16439), .A(n16315), .B(n16314), .ZN(
        P2_U2998) );
  INV_X1 U19521 ( .A(n16316), .ZN(n16318) );
  OAI21_X1 U19522 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16318), .A(
        n16317), .ZN(n16589) );
  NAND2_X1 U19523 ( .A1(n16434), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n16579) );
  NAND2_X1 U19524 ( .A1(n16410), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16319) );
  OAI211_X1 U19525 ( .C1(n16413), .C2(n16320), .A(n16579), .B(n16319), .ZN(
        n16321) );
  AOI21_X1 U19526 ( .B1(n16583), .B2(n10023), .A(n16321), .ZN(n16327) );
  NAND2_X1 U19527 ( .A1(n16323), .A2(n16322), .ZN(n16325) );
  XOR2_X1 U19528 ( .A(n16325), .B(n16324), .Z(n16587) );
  NAND2_X1 U19529 ( .A1(n16587), .A2(n16426), .ZN(n16326) );
  OAI211_X1 U19530 ( .C1(n16589), .C2(n16429), .A(n16327), .B(n16326), .ZN(
        P2_U2999) );
  OAI21_X1 U19531 ( .B1(n16343), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16316), .ZN(n16603) );
  NAND2_X1 U19532 ( .A1(n16330), .A2(n16329), .ZN(n16331) );
  XNOR2_X1 U19533 ( .A(n16328), .B(n16331), .ZN(n16600) );
  NAND2_X1 U19534 ( .A1(n16434), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n16595) );
  OAI21_X1 U19535 ( .B1(n16436), .B2(n16332), .A(n16595), .ZN(n16333) );
  AOI21_X1 U19536 ( .B1(n16433), .B2(n16334), .A(n16333), .ZN(n16335) );
  OAI21_X1 U19537 ( .B1(n16596), .B2(n16409), .A(n16335), .ZN(n16336) );
  AOI21_X1 U19538 ( .B1(n16600), .B2(n16426), .A(n16336), .ZN(n16337) );
  OAI21_X1 U19539 ( .B1(n16603), .B2(n16429), .A(n16337), .ZN(P2_U3000) );
  NAND2_X1 U19540 ( .A1(n16340), .A2(n16339), .ZN(n16341) );
  XNOR2_X1 U19541 ( .A(n16338), .B(n16341), .ZN(n16614) );
  AOI21_X1 U19542 ( .B1(n10165), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16344) );
  NOR2_X1 U19543 ( .A1(n16344), .A2(n16343), .ZN(n16604) );
  NAND2_X1 U19544 ( .A1(n16604), .A2(n16383), .ZN(n16350) );
  INV_X1 U19545 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16347) );
  NAND2_X1 U19546 ( .A1(n16433), .A2(n16345), .ZN(n16346) );
  NAND2_X1 U19547 ( .A1(n16434), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n16606) );
  OAI211_X1 U19548 ( .C1(n16347), .C2(n16436), .A(n16346), .B(n16606), .ZN(
        n16348) );
  AOI21_X1 U19549 ( .B1(n16605), .B2(n10023), .A(n16348), .ZN(n16349) );
  OAI211_X1 U19550 ( .C1(n16439), .C2(n16614), .A(n16350), .B(n16349), .ZN(
        P2_U3001) );
  XNOR2_X1 U19551 ( .A(n16342), .B(n16615), .ZN(n16627) );
  NAND2_X1 U19552 ( .A1(n10532), .A2(n16352), .ZN(n16353) );
  XNOR2_X1 U19553 ( .A(n16354), .B(n16353), .ZN(n16625) );
  NOR2_X1 U19554 ( .A1(n16619), .A2(n16409), .ZN(n16358) );
  NAND2_X1 U19555 ( .A1(n16434), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n16618) );
  NAND2_X1 U19556 ( .A1(n16410), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16355) );
  OAI211_X1 U19557 ( .C1(n16413), .C2(n16356), .A(n16618), .B(n16355), .ZN(
        n16357) );
  AOI211_X1 U19558 ( .C1(n16625), .C2(n16426), .A(n16358), .B(n16357), .ZN(
        n16359) );
  OAI21_X1 U19559 ( .B1(n16627), .B2(n16429), .A(n16359), .ZN(P2_U3002) );
  OAI21_X1 U19560 ( .B1(n16382), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16342), .ZN(n16640) );
  XNOR2_X1 U19561 ( .A(n16362), .B(n16361), .ZN(n16363) );
  XNOR2_X1 U19562 ( .A(n16364), .B(n16363), .ZN(n16638) );
  NOR2_X1 U19563 ( .A1(n16635), .A2(n16409), .ZN(n16368) );
  NAND2_X1 U19564 ( .A1(n16434), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n16634) );
  NAND2_X1 U19565 ( .A1(n16410), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16365) );
  OAI211_X1 U19566 ( .C1(n16413), .C2(n16366), .A(n16634), .B(n16365), .ZN(
        n16367) );
  AOI211_X1 U19567 ( .C1(n16638), .C2(n16426), .A(n16368), .B(n16367), .ZN(
        n16369) );
  OAI21_X1 U19568 ( .B1(n16640), .B2(n16429), .A(n16369), .ZN(P2_U3003) );
  NAND2_X1 U19569 ( .A1(n16371), .A2(n16370), .ZN(n16425) );
  INV_X1 U19570 ( .A(n16425), .ZN(n16375) );
  INV_X1 U19571 ( .A(n16372), .ZN(n16373) );
  AOI21_X1 U19572 ( .B1(n16375), .B2(n16374), .A(n16373), .ZN(n16393) );
  AOI21_X1 U19573 ( .B1(n16393), .B2(n16390), .A(n16389), .ZN(n16380) );
  INV_X1 U19574 ( .A(n16376), .ZN(n16378) );
  NAND2_X1 U19575 ( .A1(n16378), .A2(n16377), .ZN(n16379) );
  XNOR2_X1 U19576 ( .A(n16380), .B(n16379), .ZN(n16651) );
  AOI21_X1 U19577 ( .B1(n9601), .B2(n16381), .A(n16382), .ZN(n16641) );
  NAND2_X1 U19578 ( .A1(n16641), .A2(n16383), .ZN(n16388) );
  NAND2_X1 U19579 ( .A1(n16434), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n16645) );
  OAI21_X1 U19580 ( .B1(n16436), .B2(n10379), .A(n16645), .ZN(n16385) );
  NOR2_X1 U19581 ( .A1(n16646), .A2(n16409), .ZN(n16384) );
  AOI211_X1 U19582 ( .C1(n16386), .C2(n16433), .A(n16385), .B(n16384), .ZN(
        n16387) );
  OAI211_X1 U19583 ( .C1(n16651), .C2(n16439), .A(n16388), .B(n16387), .ZN(
        P2_U3004) );
  INV_X1 U19584 ( .A(n16389), .ZN(n16391) );
  NAND2_X1 U19585 ( .A1(n16391), .A2(n16390), .ZN(n16392) );
  XNOR2_X1 U19586 ( .A(n16393), .B(n16392), .ZN(n16661) );
  NOR2_X1 U19587 ( .A1(n16394), .A2(n20199), .ZN(n16653) );
  AOI21_X1 U19588 ( .B1(n16410), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16653), .ZN(n16397) );
  NAND2_X1 U19589 ( .A1(n16433), .A2(n16395), .ZN(n16396) );
  OAI211_X1 U19590 ( .C1(n16658), .C2(n16409), .A(n16397), .B(n16396), .ZN(
        n16398) );
  AOI21_X1 U19591 ( .B1(n16661), .B2(n16426), .A(n16398), .ZN(n16399) );
  OAI21_X1 U19592 ( .B1(n16664), .B2(n16429), .A(n16399), .ZN(P2_U3005) );
  XNOR2_X1 U19593 ( .A(n16401), .B(n16681), .ZN(n16418) );
  AOI22_X1 U19594 ( .A1(n16418), .A2(n16417), .B1(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16401), .ZN(n16402) );
  XOR2_X1 U19595 ( .A(n16403), .B(n16402), .Z(n16678) );
  NAND2_X1 U19596 ( .A1(n16405), .A2(n16404), .ZN(n16408) );
  INV_X1 U19597 ( .A(n16423), .ZN(n16406) );
  AOI21_X1 U19598 ( .B1(n16425), .B2(n16422), .A(n16406), .ZN(n16407) );
  XOR2_X1 U19599 ( .A(n16408), .B(n16407), .Z(n16676) );
  NOR2_X1 U19600 ( .A1(n16670), .A2(n16409), .ZN(n16415) );
  NAND2_X1 U19601 ( .A1(n16434), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n16668) );
  NAND2_X1 U19602 ( .A1(n16410), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16411) );
  OAI211_X1 U19603 ( .C1(n16413), .C2(n16412), .A(n16668), .B(n16411), .ZN(
        n16414) );
  AOI211_X1 U19604 ( .C1(n16676), .C2(n16426), .A(n16415), .B(n16414), .ZN(
        n16416) );
  OAI21_X1 U19605 ( .B1(n16678), .B2(n16429), .A(n16416), .ZN(P2_U3006) );
  XNOR2_X1 U19606 ( .A(n16418), .B(n16417), .ZN(n16692) );
  NAND2_X1 U19607 ( .A1(n16433), .A2(n16419), .ZN(n16420) );
  NAND2_X1 U19608 ( .A1(n16434), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n16679) );
  OAI211_X1 U19609 ( .C1(n21303), .C2(n16436), .A(n16420), .B(n16679), .ZN(
        n16421) );
  AOI21_X1 U19610 ( .B1(n16685), .B2(n10023), .A(n16421), .ZN(n16428) );
  NAND2_X1 U19611 ( .A1(n16423), .A2(n16422), .ZN(n16424) );
  XNOR2_X1 U19612 ( .A(n16425), .B(n16424), .ZN(n16690) );
  NAND2_X1 U19613 ( .A1(n16690), .A2(n16426), .ZN(n16427) );
  OAI211_X1 U19614 ( .C1(n16692), .C2(n16429), .A(n16428), .B(n16427), .ZN(
        P2_U3007) );
  NAND2_X1 U19615 ( .A1(n16431), .A2(n16430), .ZN(n16432) );
  XNOR2_X1 U19616 ( .A(n16432), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16707) );
  NAND2_X1 U19617 ( .A1(n16433), .A2(n19411), .ZN(n16435) );
  NAND2_X1 U19618 ( .A1(n16434), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n16699) );
  OAI211_X1 U19619 ( .C1(n16437), .C2(n16436), .A(n16435), .B(n16699), .ZN(
        n16441) );
  NOR2_X1 U19620 ( .A1(n16703), .A2(n16439), .ZN(n16440) );
  AOI211_X1 U19621 ( .C1(n10023), .C2(n19415), .A(n16441), .B(n16440), .ZN(
        n16442) );
  OAI21_X1 U19622 ( .B1(n16707), .B2(n16429), .A(n16442), .ZN(P2_U3008) );
  INV_X1 U19623 ( .A(n16444), .ZN(n16445) );
  OR2_X1 U19624 ( .A1(n16446), .A2(n16445), .ZN(n16447) );
  AOI21_X1 U19625 ( .B1(n16448), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16447), .ZN(n16449) );
  OAI21_X1 U19626 ( .B1(n16453), .B2(n16706), .A(n16452), .ZN(P2_U3018) );
  INV_X1 U19627 ( .A(n16485), .ZN(n16454) );
  NOR2_X1 U19628 ( .A1(n16455), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16481) );
  NOR2_X1 U19629 ( .A1(n16454), .A2(n16481), .ZN(n16472) );
  INV_X1 U19630 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16459) );
  INV_X1 U19631 ( .A(n16455), .ZN(n16468) );
  OAI21_X1 U19632 ( .B1(n16484), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16456) );
  OAI211_X1 U19633 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n16468), .B(n16456), .ZN(
        n16457) );
  OAI211_X1 U19634 ( .C1(n16472), .C2(n16459), .A(n16458), .B(n16457), .ZN(
        n16462) );
  NOR2_X1 U19635 ( .A1(n16460), .A2(n16669), .ZN(n16461) );
  AOI211_X1 U19636 ( .C1(n16463), .C2(n16724), .A(n16462), .B(n16461), .ZN(
        n16465) );
  NAND3_X1 U19637 ( .A1(n10512), .A2(n12739), .A3(n16467), .ZN(n16478) );
  NAND3_X1 U19638 ( .A1(n16468), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n16471), .ZN(n16469) );
  OAI211_X1 U19639 ( .C1(n16472), .C2(n16471), .A(n16470), .B(n16469), .ZN(
        n16475) );
  NOR2_X1 U19640 ( .A1(n16473), .A2(n16669), .ZN(n16474) );
  AOI211_X1 U19641 ( .C1(n16724), .C2(n16476), .A(n16475), .B(n16474), .ZN(
        n16477) );
  OAI211_X1 U19642 ( .C1(n16479), .C2(n16721), .A(n16478), .B(n16477), .ZN(
        P2_U3021) );
  OR2_X1 U19643 ( .A1(n16480), .A2(n16706), .ZN(n16493) );
  INV_X1 U19644 ( .A(n16481), .ZN(n16483) );
  OAI211_X1 U19645 ( .C1(n16485), .C2(n16484), .A(n16483), .B(n16482), .ZN(
        n16486) );
  AOI21_X1 U19646 ( .B1(n16487), .B2(n16727), .A(n16486), .ZN(n16492) );
  NAND2_X1 U19647 ( .A1(n16488), .A2(n16689), .ZN(n16491) );
  OR2_X1 U19648 ( .A1(n16489), .A2(n16708), .ZN(n16490) );
  NAND4_X1 U19649 ( .A1(n16493), .A2(n16492), .A3(n16491), .A4(n16490), .ZN(
        P2_U3022) );
  INV_X1 U19650 ( .A(n16494), .ZN(n16495) );
  OAI211_X1 U19651 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16509), .B(n16495), .ZN(
        n16496) );
  OAI211_X1 U19652 ( .C1(n16520), .C2(n16498), .A(n16497), .B(n16496), .ZN(
        n16499) );
  AOI21_X1 U19653 ( .B1(n16500), .B2(n16727), .A(n16499), .ZN(n16503) );
  OR2_X1 U19654 ( .A1(n16501), .A2(n16708), .ZN(n16502) );
  OAI211_X1 U19655 ( .C1(n16504), .C2(n16721), .A(n16503), .B(n16502), .ZN(
        n16505) );
  AOI21_X1 U19656 ( .B1(n16506), .B2(n12739), .A(n16505), .ZN(n16507) );
  INV_X1 U19657 ( .A(n16507), .ZN(P2_U3023) );
  NOR2_X1 U19658 ( .A1(n16508), .A2(n16708), .ZN(n16514) );
  INV_X1 U19659 ( .A(n16509), .ZN(n16510) );
  MUX2_X1 U19660 ( .A(n16510), .B(n16520), .S(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n16511) );
  OAI211_X1 U19661 ( .C1(n16827), .C2(n16669), .A(n16512), .B(n16511), .ZN(
        n16513) );
  NOR2_X1 U19662 ( .A1(n16514), .A2(n16513), .ZN(n16517) );
  NAND2_X1 U19663 ( .A1(n16515), .A2(n16689), .ZN(n16516) );
  OAI211_X1 U19664 ( .C1(n16518), .C2(n16706), .A(n16517), .B(n16516), .ZN(
        P2_U3024) );
  NAND2_X1 U19665 ( .A1(n16519), .A2(n16655), .ZN(n16521) );
  MUX2_X1 U19666 ( .A(n16521), .B(n16520), .S(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .Z(n16522) );
  OAI211_X1 U19667 ( .C1(n16524), .C2(n16669), .A(n16523), .B(n16522), .ZN(
        n16525) );
  AOI21_X1 U19668 ( .B1(n16526), .B2(n16724), .A(n16525), .ZN(n16528) );
  OAI211_X1 U19669 ( .C1(n16529), .C2(n16721), .A(n16528), .B(n16527), .ZN(
        P2_U3025) );
  NAND2_X1 U19670 ( .A1(n16530), .A2(n16724), .ZN(n16541) );
  NOR2_X1 U19671 ( .A1(n16729), .A2(n16536), .ZN(n16531) );
  OR2_X1 U19672 ( .A1(n16660), .A2(n16531), .ZN(n16560) );
  NAND2_X1 U19673 ( .A1(n16655), .A2(n16532), .ZN(n16533) );
  NOR2_X1 U19674 ( .A1(n16534), .A2(n16533), .ZN(n16549) );
  OAI21_X1 U19675 ( .B1(n16560), .B2(n16549), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16539) );
  NAND4_X1 U19676 ( .A1(n16536), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n16655), .A4(n16535), .ZN(n16537) );
  AND3_X1 U19677 ( .A1(n16539), .A2(n16538), .A3(n16537), .ZN(n16540) );
  OAI211_X1 U19678 ( .C1(n16542), .C2(n16669), .A(n16541), .B(n16540), .ZN(
        n16543) );
  AOI21_X1 U19679 ( .B1(n16544), .B2(n12739), .A(n16543), .ZN(n16545) );
  OAI21_X1 U19680 ( .B1(n16546), .B2(n16721), .A(n16545), .ZN(P2_U3026) );
  INV_X1 U19681 ( .A(n16547), .ZN(n16548) );
  AOI211_X1 U19682 ( .C1(n16560), .C2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n16549), .B(n16548), .ZN(n16550) );
  OAI21_X1 U19683 ( .B1(n16551), .B2(n16669), .A(n16550), .ZN(n16553) );
  OAI21_X1 U19684 ( .B1(n16556), .B2(n16721), .A(n16555), .ZN(P2_U3027) );
  NAND3_X1 U19685 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16557) );
  NOR3_X1 U19686 ( .A1(n16580), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n16557), .ZN(n16558) );
  AOI211_X1 U19687 ( .C1(n16560), .C2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n16559), .B(n16558), .ZN(n16561) );
  OAI21_X1 U19688 ( .B1(n16562), .B2(n16669), .A(n16561), .ZN(n16564) );
  INV_X1 U19689 ( .A(n16567), .ZN(n16577) );
  NAND2_X1 U19690 ( .A1(n16569), .A2(n16727), .ZN(n16571) );
  OAI211_X1 U19691 ( .C1(n16572), .C2(n16708), .A(n16571), .B(n16570), .ZN(
        n16573) );
  OAI21_X1 U19692 ( .B1(n16577), .B2(n16576), .A(n16575), .ZN(P2_U3030) );
  NOR2_X1 U19693 ( .A1(n16578), .A2(n21336), .ZN(n16582) );
  OAI21_X1 U19694 ( .B1(n16580), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16579), .ZN(n16581) );
  AOI211_X1 U19695 ( .C1(n16583), .C2(n16727), .A(n16582), .B(n16581), .ZN(
        n16584) );
  OAI21_X1 U19696 ( .B1(n16708), .B2(n16585), .A(n16584), .ZN(n16586) );
  AOI21_X1 U19697 ( .B1(n16587), .B2(n16689), .A(n16586), .ZN(n16588) );
  OAI21_X1 U19698 ( .B1(n16589), .B2(n16706), .A(n16588), .ZN(P2_U3031) );
  NOR2_X1 U19699 ( .A1(n16729), .A2(n16629), .ZN(n16590) );
  OR2_X1 U19700 ( .A1(n16660), .A2(n16590), .ZN(n16621) );
  AOI21_X1 U19701 ( .B1(n16616), .B2(n16591), .A(n16621), .ZN(n16609) );
  NOR2_X1 U19702 ( .A1(n16609), .A2(n16592), .ZN(n16598) );
  NAND3_X1 U19703 ( .A1(n16616), .A2(n16593), .A3(n16592), .ZN(n16594) );
  OAI211_X1 U19704 ( .C1(n16596), .C2(n16669), .A(n16595), .B(n16594), .ZN(
        n16597) );
  AOI211_X1 U19705 ( .C1(n16599), .C2(n16724), .A(n16598), .B(n16597), .ZN(
        n16602) );
  NAND2_X1 U19706 ( .A1(n16600), .A2(n16689), .ZN(n16601) );
  OAI211_X1 U19707 ( .C1(n16603), .C2(n16706), .A(n16602), .B(n16601), .ZN(
        P2_U3032) );
  NAND2_X1 U19708 ( .A1(n16604), .A2(n12739), .ZN(n16613) );
  AOI21_X1 U19709 ( .B1(n16616), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16608) );
  NAND2_X1 U19710 ( .A1(n16605), .A2(n16727), .ZN(n16607) );
  OAI211_X1 U19711 ( .C1(n16609), .C2(n16608), .A(n16607), .B(n16606), .ZN(
        n16610) );
  AOI21_X1 U19712 ( .B1(n16724), .B2(n16611), .A(n16610), .ZN(n16612) );
  OAI211_X1 U19713 ( .C1(n16614), .C2(n16721), .A(n16613), .B(n16612), .ZN(
        P2_U3033) );
  NAND2_X1 U19714 ( .A1(n16616), .A2(n16615), .ZN(n16617) );
  OAI211_X1 U19715 ( .C1(n16619), .C2(n16669), .A(n16618), .B(n16617), .ZN(
        n16620) );
  AOI21_X1 U19716 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16621), .A(
        n16620), .ZN(n16622) );
  OAI21_X1 U19717 ( .B1(n16708), .B2(n16623), .A(n16622), .ZN(n16624) );
  AOI21_X1 U19718 ( .B1(n16625), .B2(n16689), .A(n16624), .ZN(n16626) );
  OAI21_X1 U19719 ( .B1(n16627), .B2(n16706), .A(n16626), .ZN(P2_U3034) );
  NOR2_X1 U19720 ( .A1(n16628), .A2(n16708), .ZN(n16637) );
  INV_X1 U19721 ( .A(n16655), .ZN(n16630) );
  NOR2_X1 U19722 ( .A1(n16630), .A2(n16629), .ZN(n16632) );
  NOR3_X1 U19723 ( .A1(n16630), .A2(n16654), .A3(n9601), .ZN(n16631) );
  OAI22_X1 U19724 ( .A1(n16660), .A2(n16632), .B1(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16631), .ZN(n16633) );
  OAI211_X1 U19725 ( .C1(n16635), .C2(n16669), .A(n16634), .B(n16633), .ZN(
        n16636) );
  AOI211_X1 U19726 ( .C1(n16638), .C2(n16689), .A(n16637), .B(n16636), .ZN(
        n16639) );
  OAI21_X1 U19727 ( .B1(n16640), .B2(n16706), .A(n16639), .ZN(P2_U3035) );
  NAND2_X1 U19728 ( .A1(n16641), .A2(n12739), .ZN(n16650) );
  NOR2_X1 U19729 ( .A1(n16642), .A2(n16708), .ZN(n16648) );
  XNOR2_X1 U19730 ( .A(n16654), .B(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16643) );
  NAND2_X1 U19731 ( .A1(n16655), .A2(n16643), .ZN(n16644) );
  OAI211_X1 U19732 ( .C1(n16646), .C2(n16669), .A(n16645), .B(n16644), .ZN(
        n16647) );
  AOI211_X1 U19733 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n16660), .A(
        n16648), .B(n16647), .ZN(n16649) );
  OAI211_X1 U19734 ( .C1(n16651), .C2(n16721), .A(n16650), .B(n16649), .ZN(
        P2_U3036) );
  NAND2_X1 U19735 ( .A1(n16652), .A2(n16724), .ZN(n16657) );
  AOI21_X1 U19736 ( .B1(n16655), .B2(n16654), .A(n16653), .ZN(n16656) );
  OAI211_X1 U19737 ( .C1(n16669), .C2(n16658), .A(n16657), .B(n16656), .ZN(
        n16659) );
  AOI21_X1 U19738 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16660), .A(
        n16659), .ZN(n16663) );
  NAND2_X1 U19739 ( .A1(n16661), .A2(n16689), .ZN(n16662) );
  OAI211_X1 U19740 ( .C1(n16664), .C2(n16706), .A(n16663), .B(n16662), .ZN(
        P2_U3037) );
  INV_X1 U19741 ( .A(n16680), .ZN(n16666) );
  OAI211_X1 U19742 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16666), .B(n16665), .ZN(n16667) );
  OAI211_X1 U19743 ( .C1(n16670), .C2(n16669), .A(n16668), .B(n16667), .ZN(
        n16671) );
  AOI21_X1 U19744 ( .B1(n16724), .B2(n16672), .A(n16671), .ZN(n16673) );
  OAI21_X1 U19745 ( .B1(n16674), .B2(n16682), .A(n16673), .ZN(n16675) );
  AOI21_X1 U19746 ( .B1(n16676), .B2(n16689), .A(n16675), .ZN(n16677) );
  OAI21_X1 U19747 ( .B1(n16678), .B2(n16706), .A(n16677), .ZN(P2_U3038) );
  OAI21_X1 U19748 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16680), .A(
        n16679), .ZN(n16684) );
  NOR2_X1 U19749 ( .A1(n16682), .A2(n16681), .ZN(n16683) );
  AOI211_X1 U19750 ( .C1(n16727), .C2(n16685), .A(n16684), .B(n16683), .ZN(
        n16686) );
  OAI21_X1 U19751 ( .B1(n16708), .B2(n16687), .A(n16686), .ZN(n16688) );
  AOI21_X1 U19752 ( .B1(n16690), .B2(n16689), .A(n16688), .ZN(n16691) );
  OAI21_X1 U19753 ( .B1(n16692), .B2(n16706), .A(n16691), .ZN(P2_U3039) );
  NAND3_X1 U19754 ( .A1(n16695), .A2(n16693), .A3(n11977), .ZN(n16698) );
  OAI21_X1 U19755 ( .B1(n16729), .B2(n16695), .A(n16694), .ZN(n16696) );
  NAND2_X1 U19756 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16696), .ZN(
        n16697) );
  NAND3_X1 U19757 ( .A1(n16699), .A2(n16698), .A3(n16697), .ZN(n16700) );
  AOI21_X1 U19758 ( .B1(n19415), .B2(n16727), .A(n16700), .ZN(n16702) );
  NAND2_X1 U19759 ( .A1(n19416), .A2(n16724), .ZN(n16701) );
  OAI211_X1 U19760 ( .C1(n16703), .C2(n16721), .A(n16702), .B(n16701), .ZN(
        n16704) );
  INV_X1 U19761 ( .A(n16704), .ZN(n16705) );
  OAI21_X1 U19762 ( .B1(n16707), .B2(n16706), .A(n16705), .ZN(P2_U3040) );
  INV_X1 U19763 ( .A(n16728), .ZN(n16712) );
  INV_X1 U19764 ( .A(n19432), .ZN(n16738) );
  OAI22_X1 U19765 ( .A1(n16721), .A2(n16709), .B1(n16738), .B2(n16708), .ZN(
        n16710) );
  AOI211_X1 U19766 ( .C1(n16712), .C2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n16711), .B(n16710), .ZN(n16719) );
  AOI22_X1 U19767 ( .A1(n9835), .A2(n16727), .B1(n12739), .B2(n16713), .ZN(
        n16718) );
  OAI211_X1 U19768 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n16716), .B(n16715), .ZN(n16717) );
  NAND3_X1 U19769 ( .A1(n16719), .A2(n16718), .A3(n16717), .ZN(P2_U3045) );
  NOR2_X1 U19770 ( .A1(n16721), .A2(n16720), .ZN(n16722) );
  AOI211_X1 U19771 ( .C1(n16725), .C2(n16724), .A(n16723), .B(n16722), .ZN(
        n16732) );
  AOI22_X1 U19772 ( .A1(n9836), .A2(n16727), .B1(n12739), .B2(n16726), .ZN(
        n16731) );
  MUX2_X1 U19773 ( .A(n16729), .B(n16728), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n16730) );
  NAND3_X1 U19774 ( .A1(n16732), .A2(n16731), .A3(n16730), .ZN(P2_U3046) );
  AND2_X1 U19775 ( .A1(n20258), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20251) );
  INV_X1 U19776 ( .A(n20251), .ZN(n16736) );
  INV_X1 U19777 ( .A(n16733), .ZN(n16734) );
  NAND2_X1 U19778 ( .A1(n20255), .A2(n16734), .ZN(n16735) );
  MUX2_X1 U19779 ( .A(n16736), .B(n16735), .S(n20254), .Z(n16737) );
  OAI21_X1 U19780 ( .B1(n16738), .B2(n20104), .A(n16737), .ZN(n16739) );
  MUX2_X1 U19781 ( .A(n16739), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        n20272), .Z(P2_U3604) );
  MUX2_X1 U19782 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n16740), .S(
        n19409), .Z(n16751) );
  INV_X1 U19783 ( .A(n16754), .ZN(n20253) );
  OAI222_X1 U19784 ( .A1(n16764), .A2(n13525), .B1(n16742), .B2(n16751), .C1(
        n20253), .C2(n16741), .ZN(n16748) );
  NAND2_X1 U19785 ( .A1(n16743), .A2(P2_FLUSH_REG_SCAN_IN), .ZN(n16747) );
  OAI22_X1 U19786 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20104), .B1(n16744), 
        .B2(n19381), .ZN(n16745) );
  INV_X1 U19787 ( .A(n16745), .ZN(n16746) );
  NAND2_X1 U19788 ( .A1(n16747), .A2(n16746), .ZN(n16814) );
  MUX2_X1 U19789 ( .A(n16748), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n16809), .Z(P2_U3601) );
  AOI21_X1 U19790 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n16750), .A(
        n16749), .ZN(n16759) );
  NAND2_X1 U19791 ( .A1(n16751), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16760) );
  INV_X1 U19792 ( .A(n16760), .ZN(n16753) );
  AOI222_X1 U19793 ( .A1(n16755), .A2(n16754), .B1(n16759), .B2(n16753), .C1(
        n20254), .C2(n16752), .ZN(n16757) );
  NAND2_X1 U19794 ( .A1(n16809), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n16756) );
  OAI21_X1 U19795 ( .B1(n16757), .B2(n16809), .A(n16756), .ZN(P2_U3600) );
  OAI222_X1 U19796 ( .A1(n20264), .A2(n16764), .B1(n16760), .B2(n16759), .C1(
        n20253), .C2(n16758), .ZN(n16761) );
  MUX2_X1 U19797 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16761), .S(
        n16814), .Z(P2_U3599) );
  INV_X1 U19798 ( .A(n16762), .ZN(n16763) );
  OAI22_X1 U19799 ( .A1(n19598), .A2(n16764), .B1(n16763), .B2(n20253), .ZN(
        n16765) );
  MUX2_X1 U19800 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16765), .S(
        n16814), .Z(P2_U3596) );
  OAI21_X1 U19801 ( .B1(n19983), .B2(n20025), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n16769) );
  NOR2_X1 U19802 ( .A1(n19690), .A2(n20262), .ZN(n16772) );
  NAND2_X1 U19803 ( .A1(n19697), .A2(n16772), .ZN(n16768) );
  NAND2_X1 U19804 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20033) );
  NOR2_X1 U19805 ( .A1(n20033), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19998) );
  AND2_X1 U19806 ( .A1(n19998), .A2(n20034), .ZN(n19981) );
  AOI211_X1 U19807 ( .C1(n16774), .C2(n20104), .A(n20258), .B(n19981), .ZN(
        n16767) );
  INV_X1 U19808 ( .A(n20102), .ZN(n19996) );
  INV_X1 U19809 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16781) );
  AOI22_X1 U19810 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19576), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19575), .ZN(n20051) );
  INV_X1 U19811 ( .A(n20051), .ZN(n20106) );
  AOI22_X2 U19812 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19576), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19575), .ZN(n20109) );
  INV_X1 U19813 ( .A(n20109), .ZN(n19928) );
  AOI22_X1 U19814 ( .A1(n19983), .A2(n20106), .B1(n20025), .B2(n19928), .ZN(
        n16780) );
  INV_X1 U19815 ( .A(n16772), .ZN(n16776) );
  INV_X1 U19816 ( .A(n16773), .ZN(n19695) );
  OAI21_X1 U19817 ( .B1(n16774), .B2(n19981), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16775) );
  AND2_X1 U19818 ( .A1(n19578), .A2(n16778), .ZN(n19894) );
  AOI22_X1 U19819 ( .A1(n19982), .A2(n20048), .B1(n19981), .B2(n19894), .ZN(
        n16779) );
  OAI211_X1 U19820 ( .C1(n19987), .C2(n16781), .A(n16780), .B(n16779), .ZN(
        P2_U3144) );
  INV_X1 U19821 ( .A(n16782), .ZN(n16784) );
  OAI21_X1 U19822 ( .B1(n16784), .B2(n16783), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n16790) );
  OAI21_X1 U19823 ( .B1(n16785), .B2(n20166), .A(n19381), .ZN(n16786) );
  NAND3_X1 U19824 ( .A1(n16787), .A2(n19785), .A3(n16786), .ZN(n16788) );
  NAND3_X1 U19825 ( .A1(n16790), .A2(n16789), .A3(n16788), .ZN(P2_U3177) );
  AOI22_X1 U19826 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17721), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16801) );
  AOI22_X1 U19827 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16791), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16800) );
  AOI22_X1 U19828 ( .A1(n9628), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16792) );
  OAI21_X1 U19829 ( .B1(n12627), .B2(n21256), .A(n16792), .ZN(n16798) );
  AOI22_X1 U19830 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16796) );
  AOI22_X1 U19831 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12836), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16795) );
  AOI22_X1 U19832 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16794) );
  AOI22_X1 U19833 ( .A1(n17684), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12813), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16793) );
  NAND4_X1 U19834 ( .A1(n16796), .A2(n16795), .A3(n16794), .A4(n16793), .ZN(
        n16797) );
  AOI211_X1 U19835 ( .C1(n17738), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n16798), .B(n16797), .ZN(n16799) );
  NAND3_X1 U19836 ( .A1(n16801), .A2(n16800), .A3(n16799), .ZN(n17875) );
  INV_X1 U19837 ( .A(n17875), .ZN(n16804) );
  OAI21_X1 U19838 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n16802), .A(n17657), .ZN(
        n16803) );
  AOI22_X1 U19839 ( .A1(n17760), .A2(n16804), .B1(n16803), .B2(n17766), .ZN(
        P3_U2690) );
  INV_X1 U19840 ( .A(n16805), .ZN(n18334) );
  NOR2_X1 U19841 ( .A1(n18334), .A2(n19352), .ZN(n18712) );
  INV_X1 U19842 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19188) );
  NOR2_X1 U19843 ( .A1(n19188), .A2(n19335), .ZN(n18724) );
  OR2_X1 U19844 ( .A1(n16806), .A2(n17721), .ZN(n18708) );
  NOR2_X1 U19845 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18708), .ZN(n16807) );
  OAI21_X1 U19846 ( .B1(n16807), .B2(n19311), .A(n19063), .ZN(n18718) );
  OAI21_X1 U19847 ( .B1(n18712), .B2(n18724), .A(n18718), .ZN(n18713) );
  NAND2_X1 U19848 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19188), .ZN(n18760) );
  NAND2_X1 U19849 ( .A1(n18760), .A2(n18718), .ZN(n18711) );
  OAI21_X1 U19850 ( .B1(n18711), .B2(n18781), .A(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n16808) );
  OAI21_X1 U19851 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18713), .A(
        n16808), .ZN(P3_U2864) );
  NAND2_X1 U19852 ( .A1(n16812), .A2(n16811), .ZN(n16813) );
  OAI21_X1 U19853 ( .B1(n16814), .B2(n11639), .A(n16813), .ZN(P2_U3595) );
  AOI21_X1 U19854 ( .B1(n18617), .B2(n16816), .A(n16815), .ZN(n16817) );
  OAI21_X1 U19855 ( .B1(n16818), .B2(n18677), .A(n16817), .ZN(n16893) );
  AOI221_X1 U19856 ( .B1(n18608), .B2(n16819), .C1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n16819), .A(n18695), .ZN(
        n16823) );
  AOI22_X1 U19857 ( .A1(n18698), .A2(n16821), .B1(n18617), .B2(n16820), .ZN(
        n16890) );
  NAND2_X1 U19858 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16890), .ZN(
        n16822) );
  OAI22_X1 U19859 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16893), .B1(
        n16823), .B2(n16822), .ZN(n16825) );
  OAI211_X1 U19860 ( .C1(n16826), .C2(n18567), .A(n16825), .B(n16824), .ZN(
        P3_U2833) );
  INV_X1 U19861 ( .A(n16827), .ZN(n16828) );
  AOI22_X1 U19862 ( .A1(n16829), .A2(n13130), .B1(n16828), .B2(n19414), .ZN(
        n16845) );
  INV_X1 U19863 ( .A(n16830), .ZN(n16831) );
  NAND2_X1 U19864 ( .A1(n15691), .A2(n16831), .ZN(n16832) );
  NAND2_X1 U19865 ( .A1(n16832), .A2(n19412), .ZN(n16834) );
  NAND2_X1 U19866 ( .A1(n16834), .A2(n16833), .ZN(n16843) );
  AOI22_X1 U19867 ( .A1(n19402), .A2(P2_REIP_REG_22__SCAN_IN), .B1(n16835), 
        .B2(P2_EBX_REG_22__SCAN_IN), .ZN(n16836) );
  OAI21_X1 U19868 ( .B1(n19424), .B2(n16837), .A(n16836), .ZN(n16841) );
  NOR2_X1 U19869 ( .A1(n16839), .A2(n16838), .ZN(n16840) );
  AOI211_X1 U19870 ( .C1(n16843), .C2(n16842), .A(n16841), .B(n16840), .ZN(
        n16844) );
  NAND2_X1 U19871 ( .A1(n16845), .A2(n16844), .ZN(P2_U2833) );
  AOI22_X1 U19872 ( .A1(n20606), .A2(n16847), .B1(n16846), .B2(n16848), .ZN(
        n21190) );
  OAI211_X1 U19873 ( .C1(n16848), .C2(n21184), .A(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n21190), .ZN(n16851) );
  OAI211_X1 U19874 ( .C1(n20901), .C2(n16851), .A(n16850), .B(n16849), .ZN(
        n16853) );
  NAND2_X1 U19875 ( .A1(n20901), .A2(n16851), .ZN(n16852) );
  NAND2_X1 U19876 ( .A1(n16853), .A2(n16852), .ZN(n16855) );
  INV_X1 U19877 ( .A(n16855), .ZN(n16857) );
  AOI21_X1 U19878 ( .B1(n16855), .B2(n20836), .A(n16854), .ZN(n16856) );
  AOI21_X1 U19879 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16857), .A(
        n16856), .ZN(n16859) );
  INV_X1 U19880 ( .A(n16859), .ZN(n16862) );
  INV_X1 U19881 ( .A(n16858), .ZN(n16861) );
  OAI21_X1 U19882 ( .B1(n16859), .B2(n16858), .A(n20873), .ZN(n16860) );
  OAI21_X1 U19883 ( .B1(n16862), .B2(n16861), .A(n16860), .ZN(n16863) );
  NAND2_X1 U19884 ( .A1(n16863), .A2(n20489), .ZN(n16872) );
  NOR2_X1 U19885 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n16865) );
  OAI21_X1 U19886 ( .B1(n16866), .B2(n16865), .A(n16864), .ZN(n16868) );
  NOR2_X1 U19887 ( .A1(n16868), .A2(n16867), .ZN(n16870) );
  NAND4_X1 U19888 ( .A1(n16872), .A2(n16871), .A3(n16870), .A4(n16869), .ZN(
        n16879) );
  NAND2_X1 U19889 ( .A1(n16874), .A2(n16873), .ZN(n16876) );
  NOR3_X1 U19890 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21074), .A3(n21175), 
        .ZN(n16875) );
  OAI22_X1 U19891 ( .A1(n16877), .A2(n16876), .B1(n16880), .B2(n16875), .ZN(
        n16995) );
  AOI221_X1 U19892 ( .B1(n10144), .B2(n21185), .C1(n16879), .C2(n21185), .A(
        n16995), .ZN(n16997) );
  AOI21_X1 U19893 ( .B1(n16880), .B2(n16879), .A(n16878), .ZN(n16881) );
  OAI211_X1 U19894 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21175), .A(n16881), 
        .B(n16992), .ZN(n16882) );
  NOR2_X1 U19895 ( .A1(n16997), .A2(n16882), .ZN(n16886) );
  OR2_X1 U19896 ( .A1(n16992), .A2(n16883), .ZN(n16884) );
  NAND2_X1 U19897 ( .A1(n10144), .A2(n16884), .ZN(n16885) );
  OAI22_X1 U19898 ( .A1(n16886), .A2(n10144), .B1(n16997), .B2(n16885), .ZN(
        P1_U3161) );
  OAI21_X1 U19899 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16888), .A(
        n16887), .ZN(n17014) );
  NOR2_X1 U19900 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16889), .ZN(
        n17010) );
  AOI21_X1 U19901 ( .B1(n16891), .B2(n16890), .A(n17000), .ZN(n16892) );
  AOI21_X1 U19902 ( .B1(n17010), .B2(n16893), .A(n16892), .ZN(n16894) );
  NAND2_X1 U19903 ( .A1(n18695), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n17003) );
  OAI211_X1 U19904 ( .C1(n18567), .C2(n17014), .A(n16894), .B(n17003), .ZN(
        P3_U2832) );
  INV_X1 U19905 ( .A(n20426), .ZN(n20399) );
  INV_X1 U19906 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n17091) );
  NOR2_X1 U19907 ( .A1(n20399), .A2(n17091), .ZN(P1_U2905) );
  INV_X1 U19908 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16895) );
  NOR2_X1 U19909 ( .A1(n16895), .A2(n20269), .ZN(P2_U3047) );
  INV_X1 U19910 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18723) );
  NOR3_X1 U19911 ( .A1(n16896), .A2(n17424), .A3(n17972), .ZN(n16897) );
  NOR2_X1 U19912 ( .A1(n19183), .A2(n17930), .ZN(n17928) );
  NOR2_X1 U19913 ( .A1(n17826), .A2(n16899), .ZN(n17828) );
  NOR2_X1 U19914 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17828), .ZN(n16902) );
  OAI222_X1 U19915 ( .A1(n18723), .A2(n17920), .B1(n9660), .B2(n16902), .C1(
        n17917), .C2(n16901), .ZN(P3_U2735) );
  NAND2_X1 U19916 ( .A1(n20350), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n16904) );
  AOI21_X1 U19917 ( .B1(n20369), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16962), .ZN(n16903) );
  NAND2_X1 U19918 ( .A1(n16904), .A2(n16903), .ZN(n16905) );
  AOI21_X1 U19919 ( .B1(n16906), .B2(P1_REIP_REG_10__SCAN_IN), .A(n16905), 
        .ZN(n16907) );
  OAI21_X1 U19920 ( .B1(n16909), .B2(n16908), .A(n16907), .ZN(n16910) );
  AOI21_X1 U19921 ( .B1(n16911), .B2(n20375), .A(n16910), .ZN(n16913) );
  INV_X1 U19922 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21106) );
  NAND3_X1 U19923 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n20308), .A3(n21106), 
        .ZN(n16912) );
  OAI211_X1 U19924 ( .C1(n16914), .C2(n20325), .A(n16913), .B(n16912), .ZN(
        P1_U2830) );
  AOI22_X1 U19925 ( .A1(n16921), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16962), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16920) );
  XNOR2_X1 U19926 ( .A(n16916), .B(n16915), .ZN(n16917) );
  XNOR2_X1 U19927 ( .A(n16918), .B(n16917), .ZN(n16957) );
  AOI22_X1 U19928 ( .A1(n16957), .A2(n16926), .B1(n16931), .B2(n20387), .ZN(
        n16919) );
  OAI211_X1 U19929 ( .C1(n16929), .C2(n20319), .A(n16920), .B(n16919), .ZN(
        P1_U2992) );
  AOI22_X1 U19930 ( .A1(n16921), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n16962), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16928) );
  NAND2_X1 U19931 ( .A1(n16923), .A2(n16922), .ZN(n16924) );
  XNOR2_X1 U19932 ( .A(n16925), .B(n16924), .ZN(n16964) );
  AOI22_X1 U19933 ( .A1(n16926), .A2(n16964), .B1(n20332), .B2(n16931), .ZN(
        n16927) );
  OAI211_X1 U19934 ( .C1(n16929), .C2(n20335), .A(n16928), .B(n16927), .ZN(
        P1_U2993) );
  INV_X1 U19935 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20337) );
  NOR2_X1 U19936 ( .A1(n16929), .A2(n20344), .ZN(n16930) );
  AOI21_X1 U19937 ( .B1(n20393), .B2(n16931), .A(n16930), .ZN(n16935) );
  XNOR2_X1 U19938 ( .A(n16933), .B(n16932), .ZN(n16978) );
  OR2_X1 U19939 ( .A1(n16978), .A2(n20293), .ZN(n16934) );
  AND2_X1 U19940 ( .A1(n16935), .A2(n16934), .ZN(n16936) );
  NAND2_X1 U19941 ( .A1(n16962), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n16977) );
  OAI211_X1 U19942 ( .C1(n20337), .C2(n16937), .A(n16936), .B(n16977), .ZN(
        P1_U2994) );
  NAND2_X1 U19943 ( .A1(n16938), .A2(n16979), .ZN(n16984) );
  INV_X1 U19944 ( .A(n16938), .ZN(n20457) );
  NOR2_X1 U19945 ( .A1(n16940), .A2(n16939), .ZN(n16941) );
  AOI211_X1 U19946 ( .C1(n16942), .C2(n20457), .A(n16941), .B(n20458), .ZN(
        n16980) );
  OAI21_X1 U19947 ( .B1(n16943), .B2(n16984), .A(n16980), .ZN(n16963) );
  AOI21_X1 U19948 ( .B1(n16945), .B2(n16944), .A(n16963), .ZN(n16960) );
  OAI222_X1 U19949 ( .A1(n16947), .A2(n20486), .B1(n20348), .B2(n21103), .C1(
        n20481), .C2(n16946), .ZN(n16948) );
  INV_X1 U19950 ( .A(n16948), .ZN(n16950) );
  OAI221_X1 U19951 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16951), .C2(n16915), .A(
        n16956), .ZN(n16949) );
  OAI211_X1 U19952 ( .C1(n16960), .C2(n16951), .A(n16950), .B(n16949), .ZN(
        P1_U3023) );
  INV_X1 U19953 ( .A(n16975), .ZN(n16954) );
  AOI21_X1 U19954 ( .B1(n16954), .B2(n16953), .A(n16952), .ZN(n16955) );
  AOI22_X1 U19955 ( .A1(n16962), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n20473), 
        .B2(n9646), .ZN(n16959) );
  AOI22_X1 U19956 ( .A1(n16957), .A2(n16965), .B1(n16915), .B2(n16956), .ZN(
        n16958) );
  OAI211_X1 U19957 ( .C1(n16960), .C2(n16915), .A(n16959), .B(n16958), .ZN(
        P1_U3024) );
  AOI22_X1 U19958 ( .A1(n16962), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n20473), 
        .B2(n16961), .ZN(n16967) );
  AOI22_X1 U19959 ( .A1(n16965), .A2(n16964), .B1(n16963), .B2(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16966) );
  OAI211_X1 U19960 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16968), .A(
        n16967), .B(n16966), .ZN(P1_U3025) );
  INV_X1 U19961 ( .A(n16969), .ZN(n16971) );
  NAND2_X1 U19962 ( .A1(n16971), .A2(n16970), .ZN(n20468) );
  OAI21_X1 U19963 ( .B1(n16974), .B2(n16973), .A(n16972), .ZN(n16976) );
  AND2_X1 U19964 ( .A1(n16976), .A2(n16975), .ZN(n20390) );
  INV_X1 U19965 ( .A(n16977), .ZN(n16982) );
  OAI22_X1 U19966 ( .A1(n16980), .A2(n16979), .B1(n20481), .B2(n16978), .ZN(
        n16981) );
  AOI211_X1 U19967 ( .C1(n20473), .C2(n20390), .A(n16982), .B(n16981), .ZN(
        n16983) );
  OAI21_X1 U19968 ( .B1(n16984), .B2(n20468), .A(n16983), .ZN(P1_U3026) );
  INV_X1 U19969 ( .A(n16985), .ZN(n21189) );
  OR2_X1 U19970 ( .A1(n16986), .A2(n21189), .ZN(n16987) );
  OAI22_X1 U19971 ( .A1(n16988), .A2(n16987), .B1(n21245), .B2(n21192), .ZN(
        P1_U3468) );
  NAND4_X1 U19972 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .A3(n21074), .A4(n21175), .ZN(n16989) );
  NAND2_X1 U19973 ( .A1(n16990), .A2(n16989), .ZN(n21071) );
  INV_X1 U19974 ( .A(n21179), .ZN(n16993) );
  OAI21_X1 U19975 ( .B1(n16997), .B2(n10144), .A(n21185), .ZN(n16991) );
  OAI211_X1 U19976 ( .C1(n16993), .C2(n21175), .A(n16992), .B(n16991), .ZN(
        n16994) );
  AOI221_X1 U19977 ( .B1(n16996), .B2(n16995), .C1(n21071), .C2(n16995), .A(
        n16994), .ZN(P1_U3162) );
  NOR2_X1 U19978 ( .A1(n16997), .A2(n10144), .ZN(n16999) );
  OAI22_X1 U19979 ( .A1(n20782), .A2(n16999), .B1(n16998), .B2(n10144), .ZN(
        P1_U3466) );
  AOI21_X1 U19980 ( .B1(n17002), .B2(n17001), .A(n17000), .ZN(n17008) );
  OAI221_X1 U19981 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n17006), .C1(
        n17005), .C2(n17004), .A(n17003), .ZN(n17007) );
  AOI211_X1 U19982 ( .C1(n18140), .C2(n17009), .A(n17008), .B(n17007), .ZN(
        n17013) );
  NAND2_X1 U19983 ( .A1(n18410), .A2(n18174), .ZN(n18103) );
  NOR2_X1 U19984 ( .A1(n18387), .A2(n18103), .ZN(n18048) );
  NAND3_X1 U19985 ( .A1(n17011), .A2(n17010), .A3(n18048), .ZN(n17012) );
  OAI211_X1 U19986 ( .C1(n17014), .C2(n18248), .A(n17013), .B(n17012), .ZN(
        P3_U2800) );
  NOR3_X1 U19987 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n17016) );
  NOR4_X1 U19988 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17015) );
  NAND4_X1 U19989 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17016), .A3(n17015), .A4(
        U215), .ZN(U213) );
  INV_X2 U19990 ( .A(U214), .ZN(n17060) );
  NOR2_X1 U19991 ( .A1(n17060), .A2(n17017), .ZN(n17035) );
  INV_X1 U19992 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19442) );
  OAI222_X1 U19993 ( .A1(U214), .A2(n17091), .B1(n17063), .B2(n17018), .C1(
        U212), .C2(n19442), .ZN(U216) );
  INV_X1 U19994 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n17020) );
  INV_X2 U19995 ( .A(U212), .ZN(n17061) );
  AOI22_X1 U19996 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n17060), .ZN(n17019) );
  OAI21_X1 U19997 ( .B1(n17020), .B2(n17063), .A(n17019), .ZN(U217) );
  INV_X1 U19998 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n17022) );
  AOI22_X1 U19999 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n17060), .ZN(n17021) );
  OAI21_X1 U20000 ( .B1(n17022), .B2(n17063), .A(n17021), .ZN(U218) );
  INV_X1 U20001 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n17024) );
  AOI22_X1 U20002 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n17060), .ZN(n17023) );
  OAI21_X1 U20003 ( .B1(n17024), .B2(n17063), .A(n17023), .ZN(U219) );
  INV_X1 U20004 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n17026) );
  AOI22_X1 U20005 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n17060), .ZN(n17025) );
  OAI21_X1 U20006 ( .B1(n17026), .B2(n17063), .A(n17025), .ZN(U220) );
  AOI222_X1 U20007 ( .A1(n17061), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(n17035), 
        .B2(BUF1_REG_26__SCAN_IN), .C1(n17060), .C2(P1_DATAO_REG_26__SCAN_IN), 
        .ZN(n17027) );
  INV_X1 U20008 ( .A(n17027), .ZN(U221) );
  INV_X1 U20009 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U20010 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n17060), .ZN(n17028) );
  OAI21_X1 U20011 ( .B1(n17029), .B2(n17063), .A(n17028), .ZN(U222) );
  AOI222_X1 U20012 ( .A1(n17060), .A2(P1_DATAO_REG_24__SCAN_IN), .B1(n17035), 
        .B2(BUF1_REG_24__SCAN_IN), .C1(n17061), .C2(P2_DATAO_REG_24__SCAN_IN), 
        .ZN(n17030) );
  INV_X1 U20013 ( .A(n17030), .ZN(U223) );
  INV_X1 U20014 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n19572) );
  AOI22_X1 U20015 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n17060), .ZN(n17031) );
  OAI21_X1 U20016 ( .B1(n19572), .B2(n17063), .A(n17031), .ZN(U224) );
  INV_X1 U20017 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n19565) );
  AOI22_X1 U20018 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n17060), .ZN(n17032) );
  OAI21_X1 U20019 ( .B1(n19565), .B2(n17063), .A(n17032), .ZN(U225) );
  INV_X1 U20020 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n19559) );
  AOI22_X1 U20021 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n17060), .ZN(n17033) );
  OAI21_X1 U20022 ( .B1(n19559), .B2(n17063), .A(n17033), .ZN(U226) );
  INV_X1 U20023 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n19552) );
  AOI22_X1 U20024 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n17060), .ZN(n17034) );
  OAI21_X1 U20025 ( .B1(n19552), .B2(n17063), .A(n17034), .ZN(U227) );
  AOI222_X1 U20026 ( .A1(n17060), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n17035), 
        .B2(BUF1_REG_19__SCAN_IN), .C1(n17061), .C2(P2_DATAO_REG_19__SCAN_IN), 
        .ZN(n17036) );
  INV_X1 U20027 ( .A(n17036), .ZN(U228) );
  INV_X1 U20028 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20029 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n17060), .ZN(n17037) );
  OAI21_X1 U20030 ( .B1(n17038), .B2(n17063), .A(n17037), .ZN(U229) );
  INV_X1 U20031 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n19536) );
  AOI22_X1 U20032 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n17060), .ZN(n17039) );
  OAI21_X1 U20033 ( .B1(n19536), .B2(n17063), .A(n17039), .ZN(U230) );
  INV_X1 U20034 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20035 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n17060), .ZN(n17040) );
  OAI21_X1 U20036 ( .B1(n17041), .B2(n17063), .A(n17040), .ZN(U231) );
  AOI22_X1 U20037 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n17060), .ZN(n17042) );
  OAI21_X1 U20038 ( .B1(n14039), .B2(n17063), .A(n17042), .ZN(U232) );
  AOI22_X1 U20039 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n17060), .ZN(n17043) );
  OAI21_X1 U20040 ( .B1(n13369), .B2(n17063), .A(n17043), .ZN(U233) );
  AOI22_X1 U20041 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n17060), .ZN(n17044) );
  OAI21_X1 U20042 ( .B1(n13849), .B2(n17063), .A(n17044), .ZN(U234) );
  AOI22_X1 U20043 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n17060), .ZN(n17045) );
  OAI21_X1 U20044 ( .B1(n13781), .B2(n17063), .A(n17045), .ZN(U235) );
  AOI22_X1 U20045 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n17060), .ZN(n17046) );
  OAI21_X1 U20046 ( .B1(n13742), .B2(n17063), .A(n17046), .ZN(U236) );
  AOI22_X1 U20047 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n17060), .ZN(n17047) );
  OAI21_X1 U20048 ( .B1(n13375), .B2(n17063), .A(n17047), .ZN(U237) );
  AOI22_X1 U20049 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n17060), .ZN(n17048) );
  OAI21_X1 U20050 ( .B1(n17049), .B2(n17063), .A(n17048), .ZN(U238) );
  AOI22_X1 U20051 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n17060), .ZN(n17050) );
  OAI21_X1 U20052 ( .B1(n13640), .B2(n17063), .A(n17050), .ZN(U239) );
  AOI22_X1 U20053 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n17060), .ZN(n17051) );
  OAI21_X1 U20054 ( .B1(n13537), .B2(n17063), .A(n17051), .ZN(U240) );
  AOI22_X1 U20055 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n17060), .ZN(n17052) );
  OAI21_X1 U20056 ( .B1(n13543), .B2(n17063), .A(n17052), .ZN(U241) );
  AOI22_X1 U20057 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n17060), .ZN(n17053) );
  OAI21_X1 U20058 ( .B1(n14079), .B2(n17063), .A(n17053), .ZN(U242) );
  AOI22_X1 U20059 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n17060), .ZN(n17054) );
  OAI21_X1 U20060 ( .B1(n17055), .B2(n17063), .A(n17054), .ZN(U243) );
  AOI22_X1 U20061 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n17060), .ZN(n17056) );
  OAI21_X1 U20062 ( .B1(n16133), .B2(n17063), .A(n17056), .ZN(U244) );
  AOI22_X1 U20063 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n17060), .ZN(n17057) );
  OAI21_X1 U20064 ( .B1(n17058), .B2(n17063), .A(n17057), .ZN(U245) );
  AOI22_X1 U20065 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n17060), .ZN(n17059) );
  OAI21_X1 U20066 ( .B1(n16151), .B2(n17063), .A(n17059), .ZN(U246) );
  AOI22_X1 U20067 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n17061), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n17060), .ZN(n17062) );
  OAI21_X1 U20068 ( .B1(n17064), .B2(n17063), .A(n17062), .ZN(U247) );
  INV_X1 U20069 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n17065) );
  AOI22_X1 U20070 ( .A1(n17090), .A2(n17065), .B1(n18723), .B2(U215), .ZN(U251) );
  OAI22_X1 U20071 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n17090), .ZN(n17066) );
  INV_X1 U20072 ( .A(n17066), .ZN(U252) );
  INV_X1 U20073 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n17067) );
  INV_X1 U20074 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18733) );
  AOI22_X1 U20075 ( .A1(n17090), .A2(n17067), .B1(n18733), .B2(U215), .ZN(U253) );
  INV_X1 U20076 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n17068) );
  INV_X1 U20077 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18737) );
  AOI22_X1 U20078 ( .A1(n17090), .A2(n17068), .B1(n18737), .B2(U215), .ZN(U254) );
  INV_X1 U20079 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n17069) );
  INV_X1 U20080 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18741) );
  AOI22_X1 U20081 ( .A1(n17085), .A2(n17069), .B1(n18741), .B2(U215), .ZN(U255) );
  INV_X1 U20082 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n17070) );
  INV_X1 U20083 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18746) );
  AOI22_X1 U20084 ( .A1(n17090), .A2(n17070), .B1(n18746), .B2(U215), .ZN(U256) );
  INV_X1 U20085 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n17071) );
  INV_X1 U20086 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18751) );
  AOI22_X1 U20087 ( .A1(n17090), .A2(n17071), .B1(n18751), .B2(U215), .ZN(U257) );
  INV_X1 U20088 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n17072) );
  INV_X1 U20089 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n21237) );
  AOI22_X1 U20090 ( .A1(n17085), .A2(n17072), .B1(n21237), .B2(U215), .ZN(U258) );
  OAI22_X1 U20091 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n17085), .ZN(n17073) );
  INV_X1 U20092 ( .A(n17073), .ZN(U259) );
  INV_X1 U20093 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n17074) );
  INV_X1 U20094 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17896) );
  AOI22_X1 U20095 ( .A1(n17090), .A2(n17074), .B1(n17896), .B2(U215), .ZN(U260) );
  OAI22_X1 U20096 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n17090), .ZN(n17075) );
  INV_X1 U20097 ( .A(n17075), .ZN(U261) );
  INV_X1 U20098 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n17076) );
  INV_X1 U20099 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17887) );
  AOI22_X1 U20100 ( .A1(n17085), .A2(n17076), .B1(n17887), .B2(U215), .ZN(U262) );
  INV_X1 U20101 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n17077) );
  INV_X1 U20102 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17882) );
  AOI22_X1 U20103 ( .A1(n17085), .A2(n17077), .B1(n17882), .B2(U215), .ZN(U263) );
  OAI22_X1 U20104 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n17090), .ZN(n17078) );
  INV_X1 U20105 ( .A(n17078), .ZN(U264) );
  OAI22_X1 U20106 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17090), .ZN(n17079) );
  INV_X1 U20107 ( .A(n17079), .ZN(U265) );
  INV_X1 U20108 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n17080) );
  INV_X1 U20109 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n17868) );
  AOI22_X1 U20110 ( .A1(n17090), .A2(n17080), .B1(n17868), .B2(U215), .ZN(U266) );
  OAI22_X1 U20111 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17090), .ZN(n17081) );
  INV_X1 U20112 ( .A(n17081), .ZN(U267) );
  INV_X1 U20113 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n19535) );
  AOI22_X1 U20114 ( .A1(n17085), .A2(n13414), .B1(n19535), .B2(U215), .ZN(U268) );
  OAI22_X1 U20115 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17090), .ZN(n17082) );
  INV_X1 U20116 ( .A(n17082), .ZN(U269) );
  INV_X1 U20117 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n18738) );
  AOI22_X1 U20118 ( .A1(n17090), .A2(n17083), .B1(n18738), .B2(U215), .ZN(U270) );
  INV_X1 U20119 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n19551) );
  AOI22_X1 U20120 ( .A1(n17085), .A2(n13406), .B1(n19551), .B2(U215), .ZN(U271) );
  INV_X1 U20121 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n19558) );
  AOI22_X1 U20122 ( .A1(n17085), .A2(n13409), .B1(n19558), .B2(U215), .ZN(U272) );
  INV_X1 U20123 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19564) );
  AOI22_X1 U20124 ( .A1(n17090), .A2(n13411), .B1(n19564), .B2(U215), .ZN(U273) );
  INV_X1 U20125 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n19574) );
  AOI22_X1 U20126 ( .A1(n17090), .A2(n13436), .B1(n19574), .B2(U215), .ZN(U274) );
  INV_X1 U20127 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n21339) );
  INV_X1 U20128 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18727) );
  AOI22_X1 U20129 ( .A1(n17090), .A2(n21339), .B1(n18727), .B2(U215), .ZN(U275) );
  OAI22_X1 U20130 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17085), .ZN(n17084) );
  INV_X1 U20131 ( .A(n17084), .ZN(U276) );
  OAI22_X1 U20132 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17085), .ZN(n17086) );
  INV_X1 U20133 ( .A(n17086), .ZN(U277) );
  OAI22_X1 U20134 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17090), .ZN(n17087) );
  INV_X1 U20135 ( .A(n17087), .ZN(U278) );
  INV_X1 U20136 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n21246) );
  AOI22_X1 U20137 ( .A1(n17090), .A2(n13422), .B1(n21246), .B2(U215), .ZN(U279) );
  OAI22_X1 U20138 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17090), .ZN(n17088) );
  INV_X1 U20139 ( .A(n17088), .ZN(U280) );
  OAI22_X1 U20140 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17090), .ZN(n17089) );
  INV_X1 U20141 ( .A(n17089), .ZN(U281) );
  INV_X1 U20142 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18754) );
  AOI22_X1 U20143 ( .A1(n17090), .A2(n19442), .B1(n18754), .B2(U215), .ZN(U282) );
  INV_X1 U20144 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17934) );
  AOI222_X1 U20145 ( .A1(n17934), .A2(P3_DATAO_REG_30__SCAN_IN), .B1(n19442), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17091), .C2(
        P1_DATAO_REG_30__SCAN_IN), .ZN(n17092) );
  INV_X2 U20146 ( .A(n17095), .ZN(n17094) );
  INV_X1 U20147 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19258) );
  INV_X1 U20148 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20202) );
  AOI22_X1 U20149 ( .A1(n17094), .A2(n19258), .B1(n20202), .B2(n17095), .ZN(
        U347) );
  INV_X1 U20150 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19256) );
  INV_X1 U20151 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20200) );
  AOI22_X1 U20152 ( .A1(n17092), .A2(n19256), .B1(n20200), .B2(n17095), .ZN(
        U348) );
  INV_X1 U20153 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19253) );
  INV_X1 U20154 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20198) );
  AOI22_X1 U20155 ( .A1(n17094), .A2(n19253), .B1(n20198), .B2(n17095), .ZN(
        U349) );
  INV_X1 U20156 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19252) );
  INV_X1 U20157 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20196) );
  AOI22_X1 U20158 ( .A1(n17094), .A2(n19252), .B1(n20196), .B2(n17095), .ZN(
        U350) );
  INV_X1 U20159 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19250) );
  INV_X1 U20160 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20194) );
  AOI22_X1 U20161 ( .A1(n17094), .A2(n19250), .B1(n20194), .B2(n17095), .ZN(
        U351) );
  INV_X1 U20162 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19248) );
  INV_X1 U20163 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20192) );
  AOI22_X1 U20164 ( .A1(n17094), .A2(n19248), .B1(n20192), .B2(n17095), .ZN(
        U352) );
  INV_X1 U20165 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19247) );
  INV_X1 U20166 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20191) );
  AOI22_X1 U20167 ( .A1(n17094), .A2(n19247), .B1(n20191), .B2(n17095), .ZN(
        U353) );
  INV_X1 U20168 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19245) );
  AOI22_X1 U20169 ( .A1(n17094), .A2(n19245), .B1(n20189), .B2(n17095), .ZN(
        U354) );
  INV_X1 U20170 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19298) );
  INV_X1 U20171 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20239) );
  AOI22_X1 U20172 ( .A1(n17094), .A2(n19298), .B1(n20239), .B2(n17095), .ZN(
        U355) );
  INV_X1 U20173 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19294) );
  INV_X1 U20174 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20236) );
  AOI22_X1 U20175 ( .A1(n17094), .A2(n19294), .B1(n20236), .B2(n17095), .ZN(
        U356) );
  INV_X1 U20176 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19292) );
  INV_X1 U20177 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n21252) );
  AOI22_X1 U20178 ( .A1(n17094), .A2(n19292), .B1(n21252), .B2(n17095), .ZN(
        U357) );
  INV_X1 U20179 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19290) );
  INV_X1 U20180 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20232) );
  AOI22_X1 U20181 ( .A1(n17094), .A2(n19290), .B1(n20232), .B2(n17095), .ZN(
        U358) );
  INV_X1 U20182 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19288) );
  INV_X1 U20183 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20231) );
  AOI22_X1 U20184 ( .A1(n17094), .A2(n19288), .B1(n20231), .B2(n17095), .ZN(
        U359) );
  INV_X1 U20185 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19286) );
  INV_X1 U20186 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n21239) );
  AOI22_X1 U20187 ( .A1(n17094), .A2(n19286), .B1(n21239), .B2(n17095), .ZN(
        U360) );
  INV_X1 U20188 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19283) );
  INV_X1 U20189 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20228) );
  AOI22_X1 U20190 ( .A1(n17094), .A2(n19283), .B1(n20228), .B2(n17095), .ZN(
        U361) );
  INV_X1 U20191 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19282) );
  INV_X1 U20192 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20226) );
  AOI22_X1 U20193 ( .A1(n17094), .A2(n19282), .B1(n20226), .B2(n17095), .ZN(
        U362) );
  INV_X1 U20194 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19280) );
  INV_X1 U20195 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20224) );
  AOI22_X1 U20196 ( .A1(n17094), .A2(n19280), .B1(n20224), .B2(n17095), .ZN(
        U363) );
  INV_X1 U20197 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19278) );
  INV_X1 U20198 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20222) );
  AOI22_X1 U20199 ( .A1(n17094), .A2(n19278), .B1(n20222), .B2(n17095), .ZN(
        U364) );
  INV_X1 U20200 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19243) );
  INV_X1 U20201 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20187) );
  AOI22_X1 U20202 ( .A1(n17094), .A2(n19243), .B1(n20187), .B2(n17095), .ZN(
        U365) );
  INV_X1 U20203 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19276) );
  INV_X1 U20204 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n17093) );
  AOI22_X1 U20205 ( .A1(n17094), .A2(n19276), .B1(n17093), .B2(n17095), .ZN(
        U366) );
  INV_X1 U20206 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19274) );
  INV_X1 U20207 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20218) );
  AOI22_X1 U20208 ( .A1(n17094), .A2(n19274), .B1(n20218), .B2(n17095), .ZN(
        U367) );
  INV_X1 U20209 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19272) );
  INV_X1 U20210 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20216) );
  AOI22_X1 U20211 ( .A1(n17094), .A2(n19272), .B1(n20216), .B2(n17095), .ZN(
        U368) );
  INV_X1 U20212 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19269) );
  INV_X1 U20213 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20214) );
  AOI22_X1 U20214 ( .A1(n17094), .A2(n19269), .B1(n20214), .B2(n17095), .ZN(
        U369) );
  INV_X1 U20215 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19268) );
  INV_X1 U20216 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20212) );
  AOI22_X1 U20217 ( .A1(n17094), .A2(n19268), .B1(n20212), .B2(n17095), .ZN(
        U370) );
  INV_X1 U20218 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19266) );
  INV_X1 U20219 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20211) );
  AOI22_X1 U20220 ( .A1(n17092), .A2(n19266), .B1(n20211), .B2(n17095), .ZN(
        U371) );
  INV_X1 U20221 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19264) );
  INV_X1 U20222 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20209) );
  AOI22_X1 U20223 ( .A1(n17092), .A2(n19264), .B1(n20209), .B2(n17095), .ZN(
        U372) );
  INV_X1 U20224 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19262) );
  INV_X1 U20225 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20208) );
  AOI22_X1 U20226 ( .A1(n17094), .A2(n19262), .B1(n20208), .B2(n17095), .ZN(
        U373) );
  INV_X1 U20227 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19261) );
  INV_X1 U20228 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20206) );
  AOI22_X1 U20229 ( .A1(n17094), .A2(n19261), .B1(n20206), .B2(n17095), .ZN(
        U374) );
  INV_X1 U20230 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n21291) );
  INV_X1 U20231 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20204) );
  AOI22_X1 U20232 ( .A1(n17092), .A2(n21291), .B1(n20204), .B2(n17095), .ZN(
        U375) );
  INV_X1 U20233 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19241) );
  INV_X1 U20234 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20185) );
  AOI22_X1 U20235 ( .A1(n17094), .A2(n19241), .B1(n20185), .B2(n17095), .ZN(
        U376) );
  INV_X1 U20236 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n17096) );
  NAND2_X1 U20237 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19240), .ZN(n19230) );
  AOI22_X1 U20238 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19230), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n19237), .ZN(n19310) );
  OAI21_X1 U20239 ( .B1(n19237), .B2(n17096), .A(n19223), .ZN(P3_U2633) );
  NAND2_X1 U20240 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19214), .ZN(n17099) );
  INV_X1 U20241 ( .A(n17103), .ZN(n17097) );
  OAI21_X1 U20242 ( .B1(n17097), .B2(n17971), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17098) );
  OAI21_X1 U20243 ( .B1(n17100), .B2(n17099), .A(n17098), .ZN(P3_U2634) );
  INV_X2 U20244 ( .A(n19368), .ZN(n19349) );
  AOI21_X1 U20245 ( .B1(n19237), .B2(n19240), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n17101) );
  AOI22_X1 U20246 ( .A1(n19349), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n17101), 
        .B2(n19368), .ZN(P3_U2635) );
  OAI21_X1 U20247 ( .B1(n19224), .B2(BS16), .A(n19310), .ZN(n19308) );
  OAI21_X1 U20248 ( .B1(n19310), .B2(n19359), .A(n19308), .ZN(P3_U2636) );
  AND3_X1 U20249 ( .A1(n19153), .A2(n17103), .A3(n17102), .ZN(n19156) );
  NOR2_X1 U20250 ( .A1(n19156), .A2(n19212), .ZN(n19350) );
  INV_X1 U20251 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n21320) );
  OAI21_X1 U20252 ( .B1(n19350), .B2(n21320), .A(n17104), .ZN(P3_U2637) );
  NOR4_X1 U20253 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17108) );
  NOR4_X1 U20254 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17107) );
  NOR4_X1 U20255 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17106) );
  NOR4_X1 U20256 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17105) );
  NAND4_X1 U20257 ( .A1(n17108), .A2(n17107), .A3(n17106), .A4(n17105), .ZN(
        n17114) );
  NOR4_X1 U20258 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17112) );
  AOI211_X1 U20259 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_30__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17111) );
  NOR4_X1 U20260 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17110) );
  NOR4_X1 U20261 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17109) );
  NAND4_X1 U20262 ( .A1(n17112), .A2(n17111), .A3(n17110), .A4(n17109), .ZN(
        n17113) );
  NOR2_X1 U20263 ( .A1(n17114), .A2(n17113), .ZN(n19347) );
  INV_X1 U20264 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19305) );
  NOR3_X1 U20265 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n17116) );
  OAI21_X1 U20266 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17116), .A(n19347), .ZN(
        n17115) );
  OAI21_X1 U20267 ( .B1(n19347), .B2(n19305), .A(n17115), .ZN(P3_U2638) );
  INV_X1 U20268 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19342) );
  INV_X1 U20269 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19309) );
  AOI21_X1 U20270 ( .B1(n19342), .B2(n19309), .A(n17116), .ZN(n17117) );
  INV_X1 U20271 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19302) );
  INV_X1 U20272 ( .A(n19347), .ZN(n19345) );
  AOI22_X1 U20273 ( .A1(n19347), .A2(n17117), .B1(n19302), .B2(n19345), .ZN(
        P3_U2639) );
  INV_X1 U20274 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19293) );
  AOI21_X1 U20275 ( .B1(n17119), .B2(n17118), .A(n17431), .ZN(n17127) );
  INV_X1 U20276 ( .A(n17120), .ZN(n17126) );
  NAND2_X1 U20277 ( .A1(n17142), .A2(n17134), .ZN(n17122) );
  OAI22_X1 U20278 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17122), .B1(n17121), 
        .B2(n17471), .ZN(n17124) );
  INV_X1 U20279 ( .A(n17128), .ZN(n17129) );
  OAI21_X1 U20280 ( .B1(n17135), .B2(n17515), .A(n17129), .ZN(n17130) );
  OAI211_X1 U20281 ( .C1(n17132), .C2(n19293), .A(n17131), .B(n17130), .ZN(
        P3_U2642) );
  NAND2_X1 U20282 ( .A1(n17483), .A2(n17133), .ZN(n17161) );
  AOI22_X1 U20283 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17460), .B1(
        n17408), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17144) );
  AOI21_X1 U20284 ( .B1(n19291), .B2(n19289), .A(n17134), .ZN(n17141) );
  AOI211_X1 U20285 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17150), .A(n17135), .B(
        n17481), .ZN(n17140) );
  AOI211_X1 U20286 ( .C1(n17138), .C2(n17137), .A(n17136), .B(n17431), .ZN(
        n17139) );
  OAI211_X1 U20288 ( .C1(n19291), .C2(n17161), .A(n17144), .B(n17143), .ZN(
        P3_U2643) );
  AOI211_X1 U20289 ( .C1(n18044), .C2(n17146), .A(n17145), .B(n17431), .ZN(
        n17149) );
  OAI22_X1 U20290 ( .A1(n17147), .A2(n17471), .B1(n19289), .B2(n17161), .ZN(
        n17148) );
  AOI211_X1 U20291 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n17408), .A(n17149), .B(
        n17148), .ZN(n17152) );
  OAI211_X1 U20292 ( .C1(n17154), .C2(n17528), .A(n17470), .B(n17150), .ZN(
        n17151) );
  OAI211_X1 U20293 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n17153), .A(n17152), 
        .B(n17151), .ZN(P3_U2644) );
  AOI21_X1 U20294 ( .B1(n17169), .B2(P3_REIP_REG_25__SCAN_IN), .A(
        P3_REIP_REG_26__SCAN_IN), .ZN(n17162) );
  AOI22_X1 U20295 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17460), .B1(
        n17408), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n17160) );
  AOI211_X1 U20296 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17170), .A(n17154), .B(
        n17481), .ZN(n17158) );
  AOI211_X1 U20297 ( .C1(n18059), .C2(n17156), .A(n17155), .B(n17431), .ZN(
        n17157) );
  NOR2_X1 U20298 ( .A1(n17158), .A2(n17157), .ZN(n17159) );
  OAI211_X1 U20299 ( .C1(n17162), .C2(n17161), .A(n17160), .B(n17159), .ZN(
        P3_U2645) );
  AOI22_X1 U20300 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17460), .B1(
        n17408), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n17174) );
  INV_X1 U20301 ( .A(n17483), .ZN(n17164) );
  NOR2_X1 U20302 ( .A1(n17164), .A2(n17163), .ZN(n17168) );
  AOI211_X1 U20303 ( .C1(n18067), .C2(n17166), .A(n17165), .B(n17431), .ZN(
        n17167) );
  AOI221_X1 U20304 ( .B1(n17169), .B2(n19285), .C1(n17168), .C2(
        P3_REIP_REG_25__SCAN_IN), .A(n17167), .ZN(n17173) );
  OAI211_X1 U20305 ( .C1(n17175), .C2(n17171), .A(n17470), .B(n17170), .ZN(
        n17172) );
  NAND3_X1 U20306 ( .A1(n17174), .A2(n17173), .A3(n17172), .ZN(P3_U2646) );
  AOI21_X1 U20307 ( .B1(n17462), .B2(n17183), .A(n17468), .ZN(n17195) );
  AOI211_X1 U20308 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17192), .A(n17175), .B(
        n17481), .ZN(n17181) );
  INV_X1 U20309 ( .A(n17176), .ZN(n17177) );
  AOI211_X1 U20310 ( .C1(n18081), .C2(n17177), .A(n9756), .B(n17431), .ZN(
        n17180) );
  NOR3_X1 U20311 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17474), .A3(n17183), 
        .ZN(n17179) );
  INV_X1 U20312 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18085) );
  OAI22_X1 U20313 ( .A1(n18085), .A2(n17471), .B1(n17482), .B2(n17535), .ZN(
        n17178) );
  NOR4_X1 U20314 ( .A1(n17181), .A2(n17180), .A3(n17179), .A4(n17178), .ZN(
        n17182) );
  OAI21_X1 U20315 ( .B1(n17195), .B2(n19284), .A(n17182), .ZN(P3_U2647) );
  INV_X1 U20316 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19281) );
  AND2_X1 U20317 ( .A1(n17183), .A2(n17462), .ZN(n17184) );
  AOI22_X1 U20318 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17460), .B1(
        n17185), .B2(n17184), .ZN(n17194) );
  NOR2_X1 U20319 ( .A1(n17197), .A2(n17186), .ZN(n17187) );
  OAI22_X1 U20320 ( .A1(n17481), .A2(n17187), .B1(n17482), .B2(n17186), .ZN(
        n17191) );
  AOI211_X1 U20321 ( .C1(n18095), .C2(n17189), .A(n17188), .B(n17431), .ZN(
        n17190) );
  AOI21_X1 U20322 ( .B1(n17192), .B2(n17191), .A(n17190), .ZN(n17193) );
  OAI211_X1 U20323 ( .C1(n17195), .C2(n19281), .A(n17194), .B(n17193), .ZN(
        P3_U2648) );
  AOI21_X1 U20324 ( .B1(n17462), .B2(n17200), .A(n17468), .ZN(n17227) );
  NOR2_X1 U20325 ( .A1(n17474), .A2(n17200), .ZN(n17196) );
  NAND2_X1 U20326 ( .A1(n17196), .A2(n19277), .ZN(n17215) );
  AOI211_X1 U20327 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17213), .A(n17197), .B(
        n17481), .ZN(n17206) );
  AOI211_X1 U20328 ( .C1(n18112), .C2(n17199), .A(n17198), .B(n17431), .ZN(
        n17205) );
  NOR4_X1 U20329 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17474), .A3(n19277), 
        .A4(n17200), .ZN(n17204) );
  OAI22_X1 U20330 ( .A1(n17202), .A2(n17471), .B1(n17482), .B2(n17201), .ZN(
        n17203) );
  NOR4_X1 U20331 ( .A1(n17206), .A2(n17205), .A3(n17204), .A4(n17203), .ZN(
        n17207) );
  OAI221_X1 U20332 ( .B1(n19279), .B2(n17227), .C1(n19279), .C2(n17215), .A(
        n17207), .ZN(P3_U2649) );
  INV_X1 U20333 ( .A(n17227), .ZN(n17212) );
  AOI211_X1 U20334 ( .C1(n18124), .C2(n17209), .A(n17208), .B(n17431), .ZN(
        n17211) );
  INV_X1 U20335 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18128) );
  OAI22_X1 U20336 ( .A1(n18128), .A2(n17471), .B1(n17482), .B2(n17576), .ZN(
        n17210) );
  AOI211_X1 U20337 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n17212), .A(n17211), 
        .B(n17210), .ZN(n17216) );
  OAI211_X1 U20338 ( .C1(n17220), .C2(n17576), .A(n17470), .B(n17213), .ZN(
        n17214) );
  NAND3_X1 U20339 ( .A1(n17216), .A2(n17215), .A3(n17214), .ZN(P3_U2650) );
  INV_X1 U20340 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19275) );
  INV_X1 U20341 ( .A(n17217), .ZN(n17218) );
  AOI211_X1 U20342 ( .C1(n18139), .C2(n17219), .A(n17218), .B(n17431), .ZN(
        n17225) );
  AOI211_X1 U20343 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17236), .A(n17220), .B(
        n17481), .ZN(n17224) );
  INV_X1 U20344 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19273) );
  INV_X1 U20345 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19271) );
  NAND2_X1 U20346 ( .A1(n17462), .A2(n17228), .ZN(n17232) );
  NOR4_X1 U20347 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n19273), .A3(n19271), 
        .A4(n17232), .ZN(n17223) );
  OAI22_X1 U20348 ( .A1(n17221), .A2(n17471), .B1(n17482), .B2(n17590), .ZN(
        n17222) );
  NOR4_X1 U20349 ( .A1(n17225), .A2(n17224), .A3(n17223), .A4(n17222), .ZN(
        n17226) );
  OAI21_X1 U20350 ( .B1(n17227), .B2(n19275), .A(n17226), .ZN(P3_U2651) );
  INV_X1 U20351 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17240) );
  NOR2_X1 U20352 ( .A1(n17474), .A2(n17228), .ZN(n17252) );
  NOR2_X1 U20353 ( .A1(n17468), .A2(n17252), .ZN(n17259) );
  OAI21_X1 U20354 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n17474), .A(n17259), 
        .ZN(n17247) );
  AOI21_X1 U20355 ( .B1(n17240), .B2(n17241), .A(n17229), .ZN(n17230) );
  INV_X1 U20356 ( .A(n17230), .ZN(n18151) );
  INV_X1 U20357 ( .A(n17243), .ZN(n17231) );
  AOI221_X1 U20358 ( .B1(n17243), .B2(n18151), .C1(n17231), .C2(n17230), .A(
        n17431), .ZN(n17235) );
  INV_X1 U20359 ( .A(n17232), .ZN(n17248) );
  NAND3_X1 U20360 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n17248), .A3(n19273), 
        .ZN(n17233) );
  OAI211_X1 U20361 ( .C1(n17482), .C2(n17237), .A(n18701), .B(n17233), .ZN(
        n17234) );
  AOI211_X1 U20362 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n17247), .A(n17235), 
        .B(n17234), .ZN(n17239) );
  OAI211_X1 U20363 ( .C1(n17244), .C2(n17237), .A(n17470), .B(n17236), .ZN(
        n17238) );
  OAI211_X1 U20364 ( .C1(n17471), .C2(n17240), .A(n17239), .B(n17238), .ZN(
        P3_U2652) );
  AOI21_X1 U20365 ( .B1(n17408), .B2(P3_EBX_REG_18__SCAN_IN), .A(n18695), .ZN(
        n17251) );
  OAI21_X1 U20366 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18148), .A(
        n17241), .ZN(n18156) );
  NOR2_X1 U20367 ( .A1(n10321), .A2(n17431), .ZN(n17422) );
  INV_X1 U20368 ( .A(n17422), .ZN(n17457) );
  INV_X1 U20369 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18159) );
  OAI221_X1 U20370 ( .B1(n18156), .B2(n17275), .C1(n18156), .C2(n18159), .A(
        n19216), .ZN(n17242) );
  AOI22_X1 U20371 ( .A1(n17243), .A2(n18156), .B1(n17457), .B2(n17242), .ZN(
        n17246) );
  AOI211_X1 U20372 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17262), .A(n17244), .B(
        n17481), .ZN(n17245) );
  AOI211_X1 U20373 ( .C1(n17460), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17246), .B(n17245), .ZN(n17250) );
  OAI21_X1 U20374 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n17248), .A(n17247), 
        .ZN(n17249) );
  NAND3_X1 U20375 ( .A1(n17251), .A2(n17250), .A3(n17249), .ZN(P3_U2653) );
  INV_X1 U20376 ( .A(n17252), .ZN(n17253) );
  OAI22_X1 U20377 ( .A1(n17482), .A2(n17263), .B1(n17254), .B2(n17253), .ZN(
        n17261) );
  NAND2_X1 U20378 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9791), .ZN(
        n17255) );
  AOI21_X1 U20379 ( .B1(n10313), .B2(n17255), .A(n18148), .ZN(n18173) );
  INV_X1 U20380 ( .A(n17276), .ZN(n17256) );
  OAI21_X1 U20381 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17256), .A(
        n17255), .ZN(n18184) );
  AOI21_X1 U20382 ( .B1(n17275), .B2(n18184), .A(n17434), .ZN(n17257) );
  XNOR2_X1 U20383 ( .A(n18173), .B(n17257), .ZN(n17258) );
  OAI22_X1 U20384 ( .A1(n17259), .A2(n19270), .B1(n17431), .B2(n17258), .ZN(
        n17260) );
  NOR3_X1 U20385 ( .A1(n18695), .A2(n17261), .A3(n17260), .ZN(n17265) );
  OAI211_X1 U20386 ( .C1(n17267), .C2(n17263), .A(n17470), .B(n17262), .ZN(
        n17264) );
  OAI211_X1 U20387 ( .C1(n17471), .C2(n10313), .A(n17265), .B(n17264), .ZN(
        P3_U2654) );
  XOR2_X1 U20388 ( .A(n17266), .B(n18184), .Z(n17274) );
  AOI211_X1 U20389 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17278), .A(n17267), .B(
        n17481), .ZN(n17269) );
  OAI21_X1 U20390 ( .B1(n17482), .B2(n17618), .A(n18701), .ZN(n17268) );
  AOI211_X1 U20391 ( .C1(n17460), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n17269), .B(n17268), .ZN(n17273) );
  OAI21_X1 U20392 ( .B1(n17270), .B2(n17474), .A(n17485), .ZN(n17294) );
  NOR3_X1 U20393 ( .A1(n17474), .A2(n19263), .A3(n17293), .ZN(n17282) );
  INV_X1 U20394 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19265) );
  XNOR2_X1 U20395 ( .A(P3_REIP_REG_16__SCAN_IN), .B(n19265), .ZN(n17271) );
  AOI22_X1 U20396 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n17294), .B1(n17282), 
        .B2(n17271), .ZN(n17272) );
  OAI211_X1 U20397 ( .C1(n17431), .C2(n17274), .A(n17273), .B(n17272), .ZN(
        P3_U2655) );
  NOR2_X1 U20398 ( .A1(n17275), .A2(n17472), .ZN(n17277) );
  OAI21_X1 U20399 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18180), .A(
        n17276), .ZN(n18190) );
  AOI22_X1 U20400 ( .A1(n17408), .A2(P3_EBX_REG_15__SCAN_IN), .B1(n17277), 
        .B2(n18190), .ZN(n17286) );
  INV_X1 U20401 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18193) );
  OAI211_X1 U20402 ( .C1(n17288), .C2(n17279), .A(n17470), .B(n17278), .ZN(
        n17280) );
  OAI21_X1 U20403 ( .B1(n17471), .B2(n18193), .A(n17280), .ZN(n17281) );
  AOI221_X1 U20404 ( .B1(n17282), .B2(n19265), .C1(n17294), .C2(
        P3_REIP_REG_15__SCAN_IN), .A(n17281), .ZN(n17285) );
  INV_X1 U20405 ( .A(n18190), .ZN(n17283) );
  AOI21_X1 U20406 ( .B1(n10321), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n17431), .ZN(n17478) );
  OAI211_X1 U20407 ( .C1(n18180), .C2(n17422), .A(n17283), .B(n17478), .ZN(
        n17284) );
  NAND4_X1 U20408 ( .A1(n17286), .A2(n17285), .A3(n18701), .A4(n17284), .ZN(
        P3_U2656) );
  NAND2_X1 U20409 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17287), .ZN(
        n17299) );
  AOI21_X1 U20410 ( .B1(n10312), .B2(n17299), .A(n18180), .ZN(n18214) );
  NOR2_X1 U20411 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17299), .ZN(
        n17289) );
  NOR2_X1 U20412 ( .A1(n17289), .A2(n17472), .ZN(n17300) );
  INV_X1 U20413 ( .A(n17300), .ZN(n17298) );
  AOI211_X1 U20414 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17307), .A(n17288), .B(
        n17481), .ZN(n17292) );
  INV_X1 U20415 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17654) );
  OAI211_X1 U20416 ( .C1(n17289), .C2(n17434), .A(n19216), .B(n18214), .ZN(
        n17290) );
  OAI211_X1 U20417 ( .C1(n17482), .C2(n17654), .A(n18701), .B(n17290), .ZN(
        n17291) );
  AOI211_X1 U20418 ( .C1(n17460), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17292), .B(n17291), .ZN(n17297) );
  NOR2_X1 U20419 ( .A1(n17474), .A2(n17293), .ZN(n17295) );
  OAI21_X1 U20420 ( .B1(P3_REIP_REG_14__SCAN_IN), .B2(n17295), .A(n17294), 
        .ZN(n17296) );
  OAI211_X1 U20421 ( .C1(n18214), .C2(n17298), .A(n17297), .B(n17296), .ZN(
        P3_U2657) );
  INV_X1 U20422 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18242) );
  INV_X1 U20423 ( .A(n18314), .ZN(n18313) );
  NAND2_X1 U20424 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18313), .ZN(
        n17403) );
  NOR2_X1 U20425 ( .A1(n18318), .A2(n17403), .ZN(n17391) );
  NAND2_X1 U20426 ( .A1(n18252), .A2(n17391), .ZN(n18218) );
  NOR2_X1 U20427 ( .A1(n18242), .A2(n18218), .ZN(n17318) );
  OAI21_X1 U20428 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17318), .A(
        n17299), .ZN(n18225) );
  AOI22_X1 U20429 ( .A1(n17408), .A2(P3_EBX_REG_13__SCAN_IN), .B1(n17300), 
        .B2(n18225), .ZN(n17312) );
  INV_X1 U20430 ( .A(n17301), .ZN(n17317) );
  OAI21_X1 U20431 ( .B1(n17317), .B2(n17474), .A(n17485), .ZN(n17313) );
  NOR2_X1 U20432 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17474), .ZN(n17316) );
  INV_X1 U20433 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17304) );
  INV_X1 U20434 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n21260) );
  NAND3_X1 U20435 ( .A1(n17462), .A2(n17302), .A3(n21260), .ZN(n17303) );
  OAI211_X1 U20436 ( .C1(n17304), .C2(n17471), .A(n18701), .B(n17303), .ZN(
        n17305) );
  AOI221_X1 U20437 ( .B1(n17313), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n17316), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n17305), .ZN(n17311) );
  INV_X1 U20438 ( .A(n18225), .ZN(n17306) );
  OAI211_X1 U20439 ( .C1(n17318), .C2(n17434), .A(n17306), .B(n17478), .ZN(
        n17310) );
  OAI211_X1 U20440 ( .C1(n17314), .C2(n17308), .A(n17470), .B(n17307), .ZN(
        n17309) );
  NAND4_X1 U20441 ( .A1(n17312), .A2(n17311), .A3(n17310), .A4(n17309), .ZN(
        P3_U2658) );
  INV_X1 U20442 ( .A(n17313), .ZN(n17333) );
  AOI211_X1 U20443 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17336), .A(n17314), .B(
        n17481), .ZN(n17315) );
  AOI211_X1 U20444 ( .C1(n17317), .C2(n17316), .A(n18695), .B(n17315), .ZN(
        n17325) );
  AOI21_X1 U20445 ( .B1(n18242), .B2(n18218), .A(n17318), .ZN(n18237) );
  INV_X1 U20446 ( .A(n17391), .ZN(n17328) );
  NOR2_X1 U20447 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17328), .ZN(
        n17319) );
  AOI21_X1 U20448 ( .B1(n18252), .B2(n17319), .A(n17434), .ZN(n17320) );
  XOR2_X1 U20449 ( .A(n18237), .B(n17320), .Z(n17323) );
  OAI22_X1 U20450 ( .A1(n18242), .A2(n17471), .B1(n17482), .B2(n17321), .ZN(
        n17322) );
  AOI21_X1 U20451 ( .B1(n17323), .B2(n19216), .A(n17322), .ZN(n17324) );
  OAI211_X1 U20452 ( .C1(n19260), .C2(n17333), .A(n17325), .B(n17324), .ZN(
        P3_U2659) );
  INV_X1 U20453 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19257) );
  INV_X1 U20454 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19255) );
  NOR2_X1 U20455 ( .A1(n19257), .A2(n19255), .ZN(n17326) );
  INV_X1 U20456 ( .A(n17341), .ZN(n17371) );
  NOR2_X1 U20457 ( .A1(n17474), .A2(n17371), .ZN(n17364) );
  AOI21_X1 U20458 ( .B1(n17326), .B2(n17364), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n17334) );
  INV_X1 U20459 ( .A(n17327), .ZN(n17329) );
  NOR2_X1 U20460 ( .A1(n17329), .A2(n17328), .ZN(n17367) );
  AND3_X1 U20461 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(n17367), .ZN(n17347) );
  OAI21_X1 U20462 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17347), .A(
        n18218), .ZN(n18249) );
  INV_X1 U20463 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17473) );
  AOI21_X1 U20464 ( .B1(n17391), .B2(n17473), .A(n17434), .ZN(n17400) );
  AOI21_X1 U20465 ( .B1(n10321), .B2(n17330), .A(n17400), .ZN(n17331) );
  INV_X1 U20466 ( .A(n17331), .ZN(n17350) );
  XOR2_X1 U20467 ( .A(n18249), .B(n17350), .Z(n17332) );
  OAI22_X1 U20468 ( .A1(n17334), .A2(n17333), .B1(n17431), .B2(n17332), .ZN(
        n17335) );
  AOI211_X1 U20469 ( .C1(n17408), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18695), .B(
        n17335), .ZN(n17339) );
  OAI211_X1 U20470 ( .C1(n17342), .C2(n17337), .A(n17470), .B(n17336), .ZN(
        n17338) );
  OAI211_X1 U20471 ( .C1(n17471), .C2(n17340), .A(n17339), .B(n17338), .ZN(
        P3_U2660) );
  OAI21_X1 U20472 ( .B1(n17341), .B2(n17474), .A(n17485), .ZN(n17375) );
  AOI21_X1 U20473 ( .B1(n17364), .B2(n19255), .A(n17375), .ZN(n17353) );
  AOI211_X1 U20474 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17343), .A(n17342), .B(
        n17481), .ZN(n17346) );
  NAND3_X1 U20475 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n17364), .A3(n19257), 
        .ZN(n17344) );
  OAI211_X1 U20476 ( .C1(n17482), .C2(n17697), .A(n18701), .B(n17344), .ZN(
        n17345) );
  AOI211_X1 U20477 ( .C1(n17460), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n17346), .B(n17345), .ZN(n17352) );
  INV_X1 U20478 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17348) );
  NAND2_X1 U20479 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17367), .ZN(
        n17354) );
  AOI21_X1 U20480 ( .B1(n17348), .B2(n17354), .A(n17347), .ZN(n18260) );
  NAND3_X1 U20481 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17367), .A3(
        n17473), .ZN(n17355) );
  NAND3_X1 U20482 ( .A1(n18260), .A2(n10321), .A3(n17355), .ZN(n17349) );
  OAI211_X1 U20483 ( .C1(n18260), .C2(n17350), .A(n19216), .B(n17349), .ZN(
        n17351) );
  OAI211_X1 U20484 ( .C1(n17353), .C2(n19257), .A(n17352), .B(n17351), .ZN(
        P3_U2661) );
  OAI21_X1 U20485 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17367), .A(
        n17354), .ZN(n18277) );
  INV_X1 U20486 ( .A(n17355), .ZN(n17357) );
  AOI22_X1 U20487 ( .A1(n10321), .A2(n18277), .B1(n17367), .B2(n17473), .ZN(
        n17356) );
  NOR3_X1 U20488 ( .A1(n17357), .A2(n17356), .A3(n17431), .ZN(n17363) );
  AOI21_X1 U20489 ( .B1(n17470), .B2(n17358), .A(n17408), .ZN(n17360) );
  NOR2_X1 U20490 ( .A1(n17358), .A2(n17481), .ZN(n17370) );
  AOI22_X1 U20491 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17460), .B1(
        n17370), .B2(n17361), .ZN(n17359) );
  OAI211_X1 U20492 ( .C1(n17361), .C2(n17360), .A(n17359), .B(n18701), .ZN(
        n17362) );
  AOI211_X1 U20493 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(n17375), .A(n17363), .B(
        n17362), .ZN(n17366) );
  NAND2_X1 U20494 ( .A1(n17364), .A2(n19255), .ZN(n17365) );
  OAI211_X1 U20495 ( .C1(n17457), .C2(n18277), .A(n17366), .B(n17365), .ZN(
        P3_U2662) );
  NAND2_X1 U20496 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17391), .ZN(
        n17379) );
  AOI21_X1 U20497 ( .B1(n18288), .B2(n17379), .A(n17367), .ZN(n18291) );
  OAI21_X1 U20498 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17379), .A(
        n10321), .ZN(n17368) );
  XOR2_X1 U20499 ( .A(n18291), .B(n17368), .Z(n17378) );
  NAND2_X1 U20500 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17385), .ZN(n17369) );
  AOI22_X1 U20501 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17460), .B1(
        n17370), .B2(n17369), .ZN(n17377) );
  NAND2_X1 U20502 ( .A1(n17462), .A2(n17371), .ZN(n17372) );
  OAI22_X1 U20503 ( .A1(n17482), .A2(n17731), .B1(n17373), .B2(n17372), .ZN(
        n17374) );
  AOI211_X1 U20504 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n17375), .A(n18695), .B(
        n17374), .ZN(n17376) );
  OAI211_X1 U20505 ( .C1(n17431), .C2(n17378), .A(n17377), .B(n17376), .ZN(
        P3_U2663) );
  OAI21_X1 U20506 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17391), .A(
        n17379), .ZN(n18310) );
  XNOR2_X1 U20507 ( .A(n17400), .B(n18310), .ZN(n17381) );
  OAI22_X1 U20508 ( .A1(n18298), .A2(n17471), .B1(n17482), .B2(n17386), .ZN(
        n17380) );
  AOI211_X1 U20509 ( .C1(n19216), .C2(n17381), .A(n18695), .B(n17380), .ZN(
        n17390) );
  NOR3_X1 U20510 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17474), .A3(n17382), .ZN(
        n17398) );
  AOI21_X1 U20511 ( .B1(n17382), .B2(n17462), .A(n17468), .ZN(n17406) );
  INV_X1 U20512 ( .A(n17406), .ZN(n17383) );
  OAI21_X1 U20513 ( .B1(n17398), .B2(n17383), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n17389) );
  INV_X1 U20514 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19251) );
  NAND3_X1 U20515 ( .A1(n17462), .A2(n17384), .A3(n19251), .ZN(n17388) );
  OAI211_X1 U20516 ( .C1(n17392), .C2(n17386), .A(n17470), .B(n17385), .ZN(
        n17387) );
  NAND4_X1 U20517 ( .A1(n17390), .A2(n17389), .A3(n17388), .A4(n17387), .ZN(
        P3_U2664) );
  AOI21_X1 U20518 ( .B1(n18318), .B2(n17403), .A(n17391), .ZN(n18321) );
  NOR2_X1 U20519 ( .A1(n18321), .A2(n17431), .ZN(n17399) );
  AOI211_X1 U20520 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17409), .A(n17392), .B(
        n17481), .ZN(n17393) );
  AOI211_X1 U20521 ( .C1(n17408), .C2(P3_EBX_REG_6__SCAN_IN), .A(n18695), .B(
        n17393), .ZN(n17396) );
  INV_X1 U20522 ( .A(n17403), .ZN(n17394) );
  OAI211_X1 U20523 ( .C1(n17394), .C2(n17434), .A(n18321), .B(n17478), .ZN(
        n17395) );
  OAI211_X1 U20524 ( .C1(n17471), .C2(n18318), .A(n17396), .B(n17395), .ZN(
        n17397) );
  AOI211_X1 U20525 ( .C1(n17400), .C2(n17399), .A(n17398), .B(n17397), .ZN(
        n17401) );
  OAI21_X1 U20526 ( .B1(n17406), .B2(n19249), .A(n17401), .ZN(P3_U2665) );
  INV_X1 U20527 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17413) );
  NOR3_X1 U20528 ( .A1(n17474), .A2(n19244), .A3(n17461), .ZN(n17428) );
  AOI21_X1 U20529 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n17428), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17405) );
  INV_X1 U20530 ( .A(n18323), .ZN(n17402) );
  NOR2_X1 U20531 ( .A1(n17477), .A2(n17402), .ZN(n17415) );
  AOI21_X1 U20532 ( .B1(n17415), .B2(n17473), .A(n17434), .ZN(n17417) );
  OAI21_X1 U20533 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17415), .A(
        n17403), .ZN(n18329) );
  XOR2_X1 U20534 ( .A(n17417), .B(n18329), .Z(n17404) );
  OAI22_X1 U20535 ( .A1(n17406), .A2(n17405), .B1(n17431), .B2(n17404), .ZN(
        n17407) );
  AOI211_X1 U20536 ( .C1(n17408), .C2(P3_EBX_REG_5__SCAN_IN), .A(n18695), .B(
        n17407), .ZN(n17412) );
  OAI211_X1 U20537 ( .C1(n17419), .C2(n17410), .A(n17470), .B(n17409), .ZN(
        n17411) );
  OAI211_X1 U20538 ( .C1(n17471), .C2(n17413), .A(n17412), .B(n17411), .ZN(
        P3_U2666) );
  NOR2_X1 U20539 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17477), .ZN(
        n17454) );
  NOR2_X1 U20540 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18339), .ZN(
        n17418) );
  INV_X1 U20541 ( .A(n18339), .ZN(n17414) );
  NAND2_X1 U20542 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17414), .ZN(
        n17433) );
  AOI21_X1 U20543 ( .B1(n18347), .B2(n17433), .A(n17415), .ZN(n18344) );
  INV_X1 U20544 ( .A(n18344), .ZN(n17416) );
  AOI22_X1 U20545 ( .A1(n17454), .A2(n17418), .B1(n17417), .B2(n17416), .ZN(
        n17432) );
  NOR2_X1 U20546 ( .A1(n18347), .A2(n17471), .ZN(n17421) );
  AOI211_X1 U20547 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17443), .A(n17419), .B(
        n17481), .ZN(n17420) );
  AOI211_X1 U20548 ( .C1(n17422), .C2(n18344), .A(n17421), .B(n17420), .ZN(
        n17430) );
  OAI21_X1 U20549 ( .B1(n17423), .B2(n17474), .A(n17485), .ZN(n17442) );
  INV_X1 U20550 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19246) );
  NOR2_X1 U20551 ( .A1(n17424), .A2(n19372), .ZN(n17452) );
  OAI21_X1 U20552 ( .B1(n17738), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n17452), .ZN(n17425) );
  OAI211_X1 U20553 ( .C1(n17482), .C2(n17426), .A(n18701), .B(n17425), .ZN(
        n17427) );
  AOI221_X1 U20554 ( .B1(n17442), .B2(P3_REIP_REG_4__SCAN_IN), .C1(n17428), 
        .C2(n19246), .A(n17427), .ZN(n17429) );
  OAI211_X1 U20555 ( .C1(n17432), .C2(n17431), .A(n17430), .B(n17429), .ZN(
        P3_U2667) );
  INV_X1 U20556 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17447) );
  OAI21_X1 U20557 ( .B1(n17474), .B2(n17461), .A(n19244), .ZN(n17441) );
  INV_X1 U20558 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18367) );
  NOR2_X1 U20559 ( .A1(n17477), .A2(n18367), .ZN(n17449) );
  OAI21_X1 U20560 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17449), .A(
        n17433), .ZN(n18355) );
  AOI21_X1 U20561 ( .B1(n17473), .B2(n17449), .A(n17434), .ZN(n17453) );
  INV_X1 U20562 ( .A(n17453), .ZN(n17436) );
  OAI21_X1 U20563 ( .B1(n18355), .B2(n17436), .A(n19216), .ZN(n17435) );
  AOI21_X1 U20564 ( .B1(n18355), .B2(n17436), .A(n17435), .ZN(n17440) );
  INV_X1 U20565 ( .A(n17452), .ZN(n19374) );
  NOR2_X1 U20566 ( .A1(n19325), .A2(n12710), .ZN(n19172) );
  NAND2_X1 U20567 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19172), .ZN(
        n19165) );
  AOI21_X1 U20568 ( .B1(n17437), .B2(n19165), .A(n17738), .ZN(n19313) );
  INV_X1 U20569 ( .A(n19313), .ZN(n17438) );
  OAI22_X1 U20570 ( .A1(n17482), .A2(n17444), .B1(n19374), .B2(n17438), .ZN(
        n17439) );
  AOI211_X1 U20571 ( .C1(n17442), .C2(n17441), .A(n17440), .B(n17439), .ZN(
        n17446) );
  OAI211_X1 U20572 ( .C1(n17448), .C2(n17444), .A(n17470), .B(n17443), .ZN(
        n17445) );
  OAI211_X1 U20573 ( .C1(n17471), .C2(n17447), .A(n17446), .B(n17445), .ZN(
        P3_U2668) );
  INV_X1 U20574 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17465) );
  INV_X1 U20575 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17770) );
  INV_X1 U20576 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17777) );
  NAND2_X1 U20577 ( .A1(n17770), .A2(n17777), .ZN(n17467) );
  AOI211_X1 U20578 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17467), .A(n17448), .B(
        n17481), .ZN(n17459) );
  AOI21_X1 U20579 ( .B1(n17477), .B2(n18367), .A(n17449), .ZN(n17450) );
  INV_X1 U20580 ( .A(n17450), .ZN(n18365) );
  INV_X1 U20581 ( .A(n19165), .ZN(n17451) );
  AOI21_X1 U20582 ( .B1(n19325), .B2(n19179), .A(n17451), .ZN(n19323) );
  AOI22_X1 U20583 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n17468), .B1(n19323), 
        .B2(n17452), .ZN(n17456) );
  OAI211_X1 U20584 ( .C1(n17454), .C2(n18365), .A(n19216), .B(n17453), .ZN(
        n17455) );
  OAI211_X1 U20585 ( .C1(n17457), .C2(n18365), .A(n17456), .B(n17455), .ZN(
        n17458) );
  AOI211_X1 U20586 ( .C1(n17460), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n17459), .B(n17458), .ZN(n17464) );
  OAI211_X1 U20587 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17462), .B(n17461), .ZN(n17463) );
  OAI211_X1 U20588 ( .C1(n17465), .C2(n17482), .A(n17464), .B(n17463), .ZN(
        P3_U2669) );
  NAND2_X1 U20589 ( .A1(n17466), .A2(n19179), .ZN(n19326) );
  OAI21_X1 U20590 ( .B1(n17777), .B2(n17770), .A(n17467), .ZN(n17778) );
  INV_X1 U20591 ( .A(n17778), .ZN(n17469) );
  AOI22_X1 U20592 ( .A1(n17470), .A2(n17469), .B1(P3_REIP_REG_1__SCAN_IN), 
        .B2(n17468), .ZN(n17480) );
  OAI21_X1 U20593 ( .B1(n17473), .B2(n17472), .A(n17471), .ZN(n17476) );
  OAI22_X1 U20594 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17474), .B1(n17482), 
        .B2(n17777), .ZN(n17475) );
  AOI221_X1 U20595 ( .B1(n17478), .B2(n17477), .C1(n17476), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n17475), .ZN(n17479) );
  OAI211_X1 U20596 ( .C1(n19326), .C2(n19374), .A(n17480), .B(n17479), .ZN(
        P3_U2670) );
  NAND2_X1 U20597 ( .A1(n17482), .A2(n17481), .ZN(n17484) );
  AOI22_X1 U20598 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17484), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n17483), .ZN(n17487) );
  NAND3_X1 U20599 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19370), .A3(
        n17485), .ZN(n17486) );
  OAI211_X1 U20600 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n19374), .A(
        n17487), .B(n17486), .ZN(P3_U2671) );
  AOI22_X1 U20601 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9610), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17498) );
  AOI22_X1 U20602 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17738), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17497) );
  AOI22_X1 U20603 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n9590), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17720), .ZN(n17488) );
  OAI21_X1 U20604 ( .B1(n17489), .B2(n21273), .A(n17488), .ZN(n17495) );
  AOI22_X1 U20605 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n9597), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n17733), .ZN(n17493) );
  AOI22_X1 U20606 ( .A1(n17684), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12813), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17492) );
  AOI22_X1 U20607 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17734), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17491) );
  AOI22_X1 U20608 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n9628), .ZN(n17490) );
  NAND4_X1 U20609 ( .A1(n17493), .A2(n17492), .A3(n17491), .A4(n17490), .ZN(
        n17494) );
  AOI211_X1 U20610 ( .C1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .C2(n17719), .A(
        n17495), .B(n17494), .ZN(n17496) );
  NAND3_X1 U20611 ( .A1(n17498), .A2(n17497), .A3(n17496), .ZN(n17511) );
  AOI22_X1 U20612 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17734), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17503) );
  AOI22_X1 U20613 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17502) );
  AOI22_X1 U20614 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17684), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17501) );
  AOI22_X1 U20615 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17500) );
  NAND4_X1 U20616 ( .A1(n17503), .A2(n17502), .A3(n17501), .A4(n17500), .ZN(
        n17509) );
  AOI22_X1 U20617 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9611), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17507) );
  AOI22_X1 U20618 ( .A1(n17738), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12813), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17506) );
  AOI22_X1 U20619 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17737), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17505) );
  AOI22_X1 U20620 ( .A1(n17720), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17504) );
  NAND4_X1 U20621 ( .A1(n17507), .A2(n17506), .A3(n17505), .A4(n17504), .ZN(
        n17508) );
  NOR2_X1 U20622 ( .A1(n17509), .A2(n17508), .ZN(n17518) );
  INV_X1 U20623 ( .A(n17524), .ZN(n17517) );
  NOR3_X1 U20624 ( .A1(n17518), .A2(n17516), .A3(n17517), .ZN(n17510) );
  XNOR2_X1 U20625 ( .A(n17511), .B(n17510), .ZN(n17791) );
  NOR2_X1 U20626 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17512), .ZN(n17514) );
  OAI22_X1 U20627 ( .A1(n17791), .A2(n17766), .B1(n17514), .B2(n17513), .ZN(
        P3_U2673) );
  NAND2_X1 U20628 ( .A1(n17574), .A2(n17515), .ZN(n17522) );
  NOR2_X1 U20629 ( .A1(n17517), .A2(n17516), .ZN(n17519) );
  XNOR2_X1 U20630 ( .A(n17519), .B(n17518), .ZN(n17795) );
  AOI22_X1 U20631 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17520), .B1(n17760), 
        .B2(n17795), .ZN(n17521) );
  OAI21_X1 U20632 ( .B1(n17523), .B2(n17522), .A(n17521), .ZN(P3_U2674) );
  AOI21_X1 U20633 ( .B1(n17525), .B2(n17530), .A(n17524), .ZN(n17804) );
  NAND2_X1 U20634 ( .A1(n17760), .A2(n17804), .ZN(n17526) );
  OAI221_X1 U20635 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17529), .C1(n17528), 
        .C2(n17527), .A(n17526), .ZN(P3_U2676) );
  AOI21_X1 U20636 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17766), .A(n17538), .ZN(
        n17533) );
  OAI21_X1 U20637 ( .B1(n17532), .B2(n17531), .A(n17530), .ZN(n17810) );
  OAI22_X1 U20638 ( .A1(n17534), .A2(n17533), .B1(n17766), .B2(n17810), .ZN(
        P3_U2677) );
  NOR2_X1 U20639 ( .A1(n17535), .A2(n17539), .ZN(n17544) );
  AOI21_X1 U20640 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17766), .A(n17544), .ZN(
        n17537) );
  XNOR2_X1 U20641 ( .A(n17536), .B(n17540), .ZN(n17815) );
  OAI22_X1 U20642 ( .A1(n17538), .A2(n17537), .B1(n17766), .B2(n17815), .ZN(
        P3_U2678) );
  INV_X1 U20643 ( .A(n17539), .ZN(n17548) );
  AOI21_X1 U20644 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17766), .A(n17548), .ZN(
        n17543) );
  OAI21_X1 U20645 ( .B1(n17542), .B2(n17541), .A(n17540), .ZN(n17820) );
  OAI22_X1 U20646 ( .A1(n17544), .A2(n17543), .B1(n17766), .B2(n17820), .ZN(
        P3_U2679) );
  AOI21_X1 U20647 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17766), .A(n9753), .ZN(
        n17547) );
  XNOR2_X1 U20648 ( .A(n17546), .B(n17545), .ZN(n17825) );
  OAI22_X1 U20649 ( .A1(n17548), .A2(n17547), .B1(n17775), .B2(n17825), .ZN(
        P3_U2680) );
  AOI22_X1 U20650 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17738), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17552) );
  AOI22_X1 U20651 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12836), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17551) );
  AOI22_X1 U20652 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17550) );
  AOI22_X1 U20653 ( .A1(n9628), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17549) );
  NAND4_X1 U20654 ( .A1(n17552), .A2(n17551), .A3(n17550), .A4(n17549), .ZN(
        n17558) );
  AOI22_X1 U20655 ( .A1(n17684), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17556) );
  AOI22_X1 U20656 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12843), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17555) );
  AOI22_X1 U20657 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12813), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17554) );
  AOI22_X1 U20658 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17553) );
  NAND4_X1 U20659 ( .A1(n17556), .A2(n17555), .A3(n17554), .A4(n17553), .ZN(
        n17557) );
  NOR2_X1 U20660 ( .A1(n17558), .A2(n17557), .ZN(n17829) );
  NAND3_X1 U20661 ( .A1(n17560), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17775), 
        .ZN(n17559) );
  OAI221_X1 U20662 ( .B1(n17560), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17775), 
        .C2(n17829), .A(n17559), .ZN(P3_U2681) );
  NAND2_X1 U20663 ( .A1(n17775), .A2(n17561), .ZN(n17591) );
  AOI22_X1 U20664 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17573) );
  AOI22_X1 U20665 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17572) );
  AOI22_X1 U20666 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17734), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17562) );
  OAI21_X1 U20667 ( .B1(n17563), .B2(n21256), .A(n17562), .ZN(n17569) );
  AOI22_X1 U20668 ( .A1(n12813), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17567) );
  AOI22_X1 U20669 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17684), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17566) );
  AOI22_X1 U20670 ( .A1(n17714), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17565) );
  AOI22_X1 U20671 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17564) );
  NAND4_X1 U20672 ( .A1(n17567), .A2(n17566), .A3(n17565), .A4(n17564), .ZN(
        n17568) );
  AOI211_X1 U20673 ( .C1(n17570), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n17569), .B(n17568), .ZN(n17571) );
  NAND3_X1 U20674 ( .A1(n17573), .A2(n17572), .A3(n17571), .ZN(n17833) );
  AOI22_X1 U20675 ( .A1(n17760), .A2(n17833), .B1(n17574), .B2(n17576), .ZN(
        n17575) );
  OAI21_X1 U20676 ( .B1(n17576), .B2(n17591), .A(n17575), .ZN(P3_U2682) );
  AOI22_X1 U20677 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17684), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17587) );
  AOI22_X1 U20678 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17586) );
  AOI22_X1 U20679 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17577) );
  OAI21_X1 U20680 ( .B1(n17578), .B2(n17763), .A(n17577), .ZN(n17584) );
  AOI22_X1 U20681 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12843), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17582) );
  AOI22_X1 U20682 ( .A1(n12813), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17581) );
  AOI22_X1 U20683 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17580) );
  AOI22_X1 U20684 ( .A1(n12836), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17579) );
  NAND4_X1 U20685 ( .A1(n17582), .A2(n17581), .A3(n17580), .A4(n17579), .ZN(
        n17583) );
  AOI211_X1 U20686 ( .C1(n17738), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n17584), .B(n17583), .ZN(n17585) );
  NAND3_X1 U20687 ( .A1(n17587), .A2(n17586), .A3(n17585), .ZN(n17838) );
  NAND2_X1 U20688 ( .A1(n17760), .A2(n17838), .ZN(n17588) );
  OAI221_X1 U20689 ( .B1(n17591), .B2(n17590), .C1(n17591), .C2(n17589), .A(
        n17588), .ZN(P3_U2683) );
  INV_X1 U20690 ( .A(n17615), .ZN(n17592) );
  OAI21_X1 U20691 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17592), .A(n17775), .ZN(
        n17603) );
  AOI22_X1 U20692 ( .A1(n12813), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17596) );
  AOI22_X1 U20693 ( .A1(n17684), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17595) );
  AOI22_X1 U20694 ( .A1(n17734), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12843), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17594) );
  AOI22_X1 U20695 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17593) );
  NAND4_X1 U20696 ( .A1(n17596), .A2(n17595), .A3(n17594), .A4(n17593), .ZN(
        n17602) );
  AOI22_X1 U20697 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17600) );
  AOI22_X1 U20698 ( .A1(n17714), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12786), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17599) );
  AOI22_X1 U20699 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14270), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17598) );
  AOI22_X1 U20700 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17597) );
  NAND4_X1 U20701 ( .A1(n17600), .A2(n17599), .A3(n17598), .A4(n17597), .ZN(
        n17601) );
  NOR2_X1 U20702 ( .A1(n17602), .A2(n17601), .ZN(n17847) );
  OAI22_X1 U20703 ( .A1(n17604), .A2(n17603), .B1(n17847), .B2(n17766), .ZN(
        P3_U2684) );
  AOI22_X1 U20704 ( .A1(n17684), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12786), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17608) );
  AOI22_X1 U20705 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17738), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17607) );
  AOI22_X1 U20706 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17606) );
  AOI22_X1 U20707 ( .A1(n9628), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17605) );
  NAND4_X1 U20708 ( .A1(n17608), .A2(n17607), .A3(n17606), .A4(n17605), .ZN(
        n17614) );
  AOI22_X1 U20709 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17612) );
  AOI22_X1 U20710 ( .A1(n9611), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17734), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17611) );
  AOI22_X1 U20711 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17610) );
  AOI22_X1 U20712 ( .A1(n12813), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17609) );
  NAND4_X1 U20713 ( .A1(n17612), .A2(n17611), .A3(n17610), .A4(n17609), .ZN(
        n17613) );
  NOR2_X1 U20714 ( .A1(n17614), .A2(n17613), .ZN(n17852) );
  OAI21_X1 U20715 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n9739), .A(n17615), .ZN(
        n17616) );
  AOI22_X1 U20716 ( .A1(n17760), .A2(n17852), .B1(n17616), .B2(n17775), .ZN(
        P3_U2685) );
  NOR3_X1 U20717 ( .A1(n17826), .A2(n17657), .A3(n17617), .ZN(n17630) );
  INV_X1 U20718 ( .A(n17630), .ZN(n17655) );
  NOR2_X1 U20719 ( .A1(n17618), .A2(n17655), .ZN(n17642) );
  AOI21_X1 U20720 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17766), .A(n17642), .ZN(
        n17629) );
  AOI22_X1 U20721 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12836), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17622) );
  AOI22_X1 U20722 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17621) );
  AOI22_X1 U20723 ( .A1(n17720), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17620) );
  AOI22_X1 U20724 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17619) );
  NAND4_X1 U20725 ( .A1(n17622), .A2(n17621), .A3(n17620), .A4(n17619), .ZN(
        n17628) );
  AOI22_X1 U20726 ( .A1(n17684), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12813), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17626) );
  AOI22_X1 U20727 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17625) );
  AOI22_X1 U20728 ( .A1(n17738), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17624) );
  AOI22_X1 U20729 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17721), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17623) );
  NAND4_X1 U20730 ( .A1(n17626), .A2(n17625), .A3(n17624), .A4(n17623), .ZN(
        n17627) );
  NOR2_X1 U20731 ( .A1(n17628), .A2(n17627), .ZN(n17857) );
  OAI22_X1 U20732 ( .A1(n9739), .A2(n17629), .B1(n17857), .B2(n17766), .ZN(
        P3_U2686) );
  AOI21_X1 U20733 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17766), .A(n17630), .ZN(
        n17641) );
  AOI22_X1 U20734 ( .A1(n12813), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17634) );
  AOI22_X1 U20735 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17633) );
  AOI22_X1 U20736 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16791), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17632) );
  AOI22_X1 U20737 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17631) );
  NAND4_X1 U20738 ( .A1(n17634), .A2(n17633), .A3(n17632), .A4(n17631), .ZN(
        n17640) );
  AOI22_X1 U20739 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9610), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17638) );
  AOI22_X1 U20740 ( .A1(n17714), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17637) );
  AOI22_X1 U20741 ( .A1(n17684), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17734), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17636) );
  AOI22_X1 U20742 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17635) );
  NAND4_X1 U20743 ( .A1(n17638), .A2(n17637), .A3(n17636), .A4(n17635), .ZN(
        n17639) );
  NOR2_X1 U20744 ( .A1(n17640), .A2(n17639), .ZN(n17863) );
  OAI22_X1 U20745 ( .A1(n17642), .A2(n17641), .B1(n17863), .B2(n17766), .ZN(
        P3_U2687) );
  AOI22_X1 U20746 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17720), .ZN(n17647) );
  AOI22_X1 U20747 ( .A1(n17684), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17738), .ZN(n17646) );
  AOI22_X1 U20748 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n17643), .ZN(n17645) );
  AOI22_X1 U20749 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n9628), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17719), .ZN(n17644) );
  NAND4_X1 U20750 ( .A1(n17647), .A2(n17646), .A3(n17645), .A4(n17644), .ZN(
        n17653) );
  AOI22_X1 U20751 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17651) );
  AOI22_X1 U20752 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n9610), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17650) );
  AOI22_X1 U20753 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17734), .ZN(n17649) );
  AOI22_X1 U20754 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12813), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17733), .ZN(n17648) );
  NAND4_X1 U20755 ( .A1(n17651), .A2(n17650), .A3(n17649), .A4(n17648), .ZN(
        n17652) );
  NOR2_X1 U20756 ( .A1(n17653), .A2(n17652), .ZN(n17865) );
  NOR2_X1 U20757 ( .A1(n17654), .A2(n17657), .ZN(n17670) );
  OAI21_X1 U20758 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17670), .A(n17655), .ZN(
        n17656) );
  AOI22_X1 U20759 ( .A1(n17760), .A2(n17865), .B1(n17656), .B2(n17775), .ZN(
        P3_U2688) );
  INV_X1 U20760 ( .A(n17657), .ZN(n17658) );
  OAI21_X1 U20761 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17658), .A(n17775), .ZN(
        n17669) );
  AOI22_X1 U20762 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17662) );
  AOI22_X1 U20763 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17661) );
  AOI22_X1 U20764 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17660) );
  AOI22_X1 U20765 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17659) );
  NAND4_X1 U20766 ( .A1(n17662), .A2(n17661), .A3(n17660), .A4(n17659), .ZN(
        n17668) );
  AOI22_X1 U20767 ( .A1(n17714), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17666) );
  AOI22_X1 U20768 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12836), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17665) );
  AOI22_X1 U20769 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17664) );
  AOI22_X1 U20770 ( .A1(n17684), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12813), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17663) );
  NAND4_X1 U20771 ( .A1(n17666), .A2(n17665), .A3(n17664), .A4(n17663), .ZN(
        n17667) );
  NOR2_X1 U20772 ( .A1(n17668), .A2(n17667), .ZN(n17874) );
  OAI22_X1 U20773 ( .A1(n17670), .A2(n17669), .B1(n17874), .B2(n17766), .ZN(
        P3_U2689) );
  OR2_X1 U20774 ( .A1(n17826), .A2(n17671), .ZN(n17695) );
  AOI22_X1 U20775 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17675) );
  AOI22_X1 U20776 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17674) );
  AOI22_X1 U20777 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9611), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17673) );
  AOI22_X1 U20778 ( .A1(n9628), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17672) );
  NAND4_X1 U20779 ( .A1(n17675), .A2(n17674), .A3(n17673), .A4(n17672), .ZN(
        n17682) );
  AOI22_X1 U20780 ( .A1(n17714), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12813), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17680) );
  AOI22_X1 U20781 ( .A1(n17684), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12786), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17679) );
  AOI22_X1 U20782 ( .A1(n17734), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17678) );
  AOI22_X1 U20783 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17677) );
  NAND4_X1 U20784 ( .A1(n17680), .A2(n17679), .A3(n17678), .A4(n17677), .ZN(
        n17681) );
  NOR2_X1 U20785 ( .A1(n17682), .A2(n17681), .ZN(n17879) );
  NAND3_X1 U20786 ( .A1(n17695), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n17775), 
        .ZN(n17683) );
  OAI221_X1 U20787 ( .B1(n17695), .B2(P3_EBX_REG_12__SCAN_IN), .C1(n17775), 
        .C2(n17879), .A(n17683), .ZN(P3_U2691) );
  AOI22_X1 U20788 ( .A1(n17714), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17688) );
  AOI22_X1 U20789 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17687) );
  AOI22_X1 U20790 ( .A1(n17734), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17686) );
  AOI22_X1 U20791 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17684), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17685) );
  NAND4_X1 U20792 ( .A1(n17688), .A2(n17687), .A3(n17686), .A4(n17685), .ZN(
        n17694) );
  AOI22_X1 U20793 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17692) );
  AOI22_X1 U20794 ( .A1(n12813), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17643), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17691) );
  AOI22_X1 U20795 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17690) );
  AOI22_X1 U20796 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9597), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17689) );
  NAND4_X1 U20797 ( .A1(n17692), .A2(n17691), .A3(n17690), .A4(n17689), .ZN(
        n17693) );
  NOR2_X1 U20798 ( .A1(n17694), .A2(n17693), .ZN(n17884) );
  OAI211_X1 U20799 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n17713), .A(n17695), .B(
        n17766), .ZN(n17696) );
  OAI21_X1 U20800 ( .B1(n17884), .B2(n17775), .A(n17696), .ZN(P3_U2692) );
  AOI21_X1 U20801 ( .B1(n17697), .B2(n17728), .A(n17760), .ZN(n17698) );
  INV_X1 U20802 ( .A(n17698), .ZN(n17712) );
  AOI22_X1 U20803 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12813), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17710) );
  AOI22_X1 U20804 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17709) );
  AOI22_X1 U20805 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14270), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17699) );
  OAI21_X1 U20806 ( .B1(n17700), .B2(n17774), .A(n17699), .ZN(n17707) );
  AOI22_X1 U20807 ( .A1(n17714), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17705) );
  AOI22_X1 U20808 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9591), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17704) );
  AOI22_X1 U20809 ( .A1(n17684), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17701), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17703) );
  AOI22_X1 U20810 ( .A1(n17734), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17702) );
  NAND4_X1 U20811 ( .A1(n17705), .A2(n17704), .A3(n17703), .A4(n17702), .ZN(
        n17706) );
  AOI211_X1 U20812 ( .C1(n12842), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n17707), .B(n17706), .ZN(n17708) );
  NAND3_X1 U20813 ( .A1(n17710), .A2(n17709), .A3(n17708), .ZN(n17888) );
  INV_X1 U20814 ( .A(n17888), .ZN(n17711) );
  OAI22_X1 U20815 ( .A1(n17713), .A2(n17712), .B1(n17711), .B2(n17766), .ZN(
        P3_U2693) );
  AOI22_X1 U20816 ( .A1(n17734), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17733), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17718) );
  AOI22_X1 U20817 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12786), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17717) );
  AOI22_X1 U20818 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9611), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17716) );
  AOI22_X1 U20819 ( .A1(n17714), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17715) );
  NAND4_X1 U20820 ( .A1(n17718), .A2(n17717), .A3(n17716), .A4(n17715), .ZN(
        n17727) );
  AOI22_X1 U20821 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17725) );
  AOI22_X1 U20822 ( .A1(n14270), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12813), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17724) );
  AOI22_X1 U20823 ( .A1(n17684), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17723) );
  AOI22_X1 U20824 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17722) );
  NAND4_X1 U20825 ( .A1(n17725), .A2(n17724), .A3(n17723), .A4(n17722), .ZN(
        n17726) );
  NOR2_X1 U20826 ( .A1(n17727), .A2(n17726), .ZN(n17893) );
  OAI21_X1 U20827 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n9766), .A(n17728), .ZN(
        n17729) );
  AOI22_X1 U20828 ( .A1(n17760), .A2(n17893), .B1(n17729), .B2(n17775), .ZN(
        P3_U2694) );
  AOI21_X1 U20829 ( .B1(n17731), .B2(n17730), .A(n9766), .ZN(n17748) );
  AOI22_X1 U20830 ( .A1(n17701), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17747) );
  AOI22_X1 U20831 ( .A1(n17733), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17732), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17746) );
  AOI22_X1 U20832 ( .A1(n12813), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17734), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17735) );
  OAI21_X1 U20833 ( .B1(n17736), .B2(n21267), .A(n17735), .ZN(n17744) );
  AOI22_X1 U20834 ( .A1(n17737), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17742) );
  AOI22_X1 U20835 ( .A1(n12842), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14270), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17741) );
  AOI22_X1 U20836 ( .A1(n17570), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17738), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17740) );
  AOI22_X1 U20837 ( .A1(n9610), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17739) );
  NAND4_X1 U20838 ( .A1(n17742), .A2(n17741), .A3(n17740), .A4(n17739), .ZN(
        n17743) );
  AOI211_X1 U20839 ( .C1(n9597), .C2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n17744), .B(n17743), .ZN(n17745) );
  NAND3_X1 U20840 ( .A1(n17747), .A2(n17746), .A3(n17745), .ZN(n17897) );
  MUX2_X1 U20841 ( .A(n17748), .B(n17897), .S(n17760), .Z(P3_U2695) );
  NAND2_X1 U20842 ( .A1(n12696), .A2(n17749), .ZN(n17751) );
  NOR2_X1 U20843 ( .A1(n17760), .A2(n17749), .ZN(n17752) );
  AOI22_X1 U20844 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17760), .B1(
        P3_EBX_REG_7__SCAN_IN), .B2(n17752), .ZN(n17750) );
  OAI21_X1 U20845 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17751), .A(n17750), .ZN(
        P3_U2696) );
  OAI21_X1 U20846 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17753), .A(n17752), .ZN(
        n17754) );
  OAI21_X1 U20847 ( .B1(n17775), .B2(n17755), .A(n17754), .ZN(P3_U2697) );
  INV_X1 U20848 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17759) );
  OAI21_X1 U20849 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17757), .A(n17756), .ZN(
        n17758) );
  AOI22_X1 U20850 ( .A1(n17760), .A2(n17759), .B1(n17758), .B2(n17766), .ZN(
        P3_U2698) );
  NOR2_X1 U20851 ( .A1(n17761), .A2(n17782), .ZN(n17769) );
  INV_X1 U20852 ( .A(n17769), .ZN(n17764) );
  NAND3_X1 U20853 ( .A1(n17764), .A2(P3_EBX_REG_4__SCAN_IN), .A3(n17775), .ZN(
        n17762) );
  OAI221_X1 U20854 ( .B1(n17764), .B2(P3_EBX_REG_4__SCAN_IN), .C1(n17775), 
        .C2(n17763), .A(n17762), .ZN(P3_U2699) );
  NAND3_X1 U20855 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17765) );
  NOR2_X1 U20856 ( .A1(n17765), .A2(n17782), .ZN(n17772) );
  AOI21_X1 U20857 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17766), .A(n17772), .ZN(
        n17768) );
  INV_X1 U20858 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17767) );
  OAI22_X1 U20859 ( .A1(n17769), .A2(n17768), .B1(n17767), .B2(n17766), .ZN(
        P3_U2700) );
  NOR2_X1 U20860 ( .A1(n17770), .A2(n17777), .ZN(n17771) );
  AOI221_X1 U20861 ( .B1(n17771), .B2(n17779), .C1(n17826), .C2(n17779), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17773) );
  AOI211_X1 U20862 ( .C1(n17760), .C2(n17774), .A(n17773), .B(n17772), .ZN(
        P3_U2701) );
  INV_X1 U20863 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17776) );
  OAI222_X1 U20864 ( .A1(n17778), .A2(n17782), .B1(n17777), .B2(n17779), .C1(
        n17776), .C2(n17775), .ZN(P3_U2702) );
  AOI22_X1 U20865 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17760), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17780), .ZN(n17781) );
  OAI21_X1 U20866 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17782), .A(n17781), .ZN(
        P3_U2703) );
  INV_X1 U20867 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18003) );
  INV_X1 U20868 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17995) );
  INV_X1 U20869 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18042) );
  INV_X1 U20870 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n18037) );
  INV_X1 U20871 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18035) );
  INV_X1 U20872 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18033) );
  INV_X1 U20873 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18029) );
  INV_X1 U20874 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18027) );
  NOR4_X1 U20875 ( .A1(n18035), .A2(n18033), .A3(n18029), .A4(n18027), .ZN(
        n17783) );
  NAND3_X1 U20876 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(n17783), .ZN(n17869) );
  NOR2_X1 U20877 ( .A1(n18037), .A2(n17869), .ZN(n17864) );
  NAND2_X1 U20878 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .ZN(n17827) );
  NAND4_X1 U20879 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .A3(P3_EAX_REG_20__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17784)
         );
  NAND2_X1 U20880 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17822), .ZN(n17821) );
  NOR2_X1 U20881 ( .A1(n17826), .A2(n17821), .ZN(n17816) );
  NAND2_X1 U20882 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17816), .ZN(n17817) );
  INV_X1 U20883 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17999) );
  NAND2_X1 U20884 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17792), .ZN(n17788) );
  NAND2_X1 U20885 ( .A1(n17788), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n17787) );
  NOR2_X2 U20886 ( .A1(n17785), .A2(n17930), .ZN(n17858) );
  NAND2_X1 U20887 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17858), .ZN(n17786) );
  OAI221_X1 U20888 ( .B1(n17788), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n17787), 
        .C2(n17921), .A(n17786), .ZN(P3_U2704) );
  NOR2_X2 U20889 ( .A1(n18745), .A2(n17930), .ZN(n17859) );
  AOI22_X1 U20890 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17859), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17858), .ZN(n17790) );
  OAI211_X1 U20891 ( .C1(n17792), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17930), .B(
        n17788), .ZN(n17789) );
  OAI211_X1 U20892 ( .C1(n17791), .C2(n17917), .A(n17790), .B(n17789), .ZN(
        P3_U2705) );
  INV_X1 U20893 ( .A(n17792), .ZN(n17794) );
  OAI21_X1 U20894 ( .B1(n17921), .B2(n18003), .A(n17799), .ZN(n17793) );
  AOI22_X1 U20895 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n17858), .B1(n17794), .B2(
        n17793), .ZN(n17797) );
  AOI22_X1 U20896 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17859), .B1(n17795), .B2(
        n17927), .ZN(n17796) );
  NAND2_X1 U20897 ( .A1(n17797), .A2(n17796), .ZN(P3_U2706) );
  AOI22_X1 U20898 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17859), .B1(n17798), .B2(
        n17927), .ZN(n17801) );
  OAI211_X1 U20899 ( .C1(n17802), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17930), .B(
        n17799), .ZN(n17800) );
  OAI211_X1 U20900 ( .C1(n17842), .C2(n21246), .A(n17801), .B(n17800), .ZN(
        P3_U2707) );
  OAI21_X1 U20901 ( .B1(n17921), .B2(n17999), .A(n17807), .ZN(n17803) );
  AOI22_X1 U20902 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n17858), .B1(n10189), .B2(
        n17803), .ZN(n17806) );
  AOI22_X1 U20903 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17859), .B1(n17804), .B2(
        n17927), .ZN(n17805) );
  NAND2_X1 U20904 ( .A1(n17806), .A2(n17805), .ZN(P3_U2708) );
  AOI22_X1 U20905 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17859), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17858), .ZN(n17809) );
  OAI211_X1 U20906 ( .C1(n17811), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17930), .B(
        n17807), .ZN(n17808) );
  OAI211_X1 U20907 ( .C1(n17917), .C2(n17810), .A(n17809), .B(n17808), .ZN(
        P3_U2709) );
  AOI22_X1 U20908 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17859), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17858), .ZN(n17814) );
  AOI211_X1 U20909 ( .C1(n17995), .C2(n17817), .A(n17811), .B(n17921), .ZN(
        n17812) );
  INV_X1 U20910 ( .A(n17812), .ZN(n17813) );
  OAI211_X1 U20911 ( .C1(n17917), .C2(n17815), .A(n17814), .B(n17813), .ZN(
        P3_U2710) );
  AOI22_X1 U20912 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17859), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17858), .ZN(n17819) );
  OAI211_X1 U20913 ( .C1(n17816), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17930), .B(
        n17817), .ZN(n17818) );
  OAI211_X1 U20914 ( .C1(n17820), .C2(n17917), .A(n17819), .B(n17818), .ZN(
        P3_U2711) );
  AOI22_X1 U20915 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17859), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17858), .ZN(n17824) );
  OAI211_X1 U20916 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17822), .A(n17930), .B(
        n17821), .ZN(n17823) );
  OAI211_X1 U20917 ( .C1(n17825), .C2(n17917), .A(n17824), .B(n17823), .ZN(
        P3_U2712) );
  INV_X1 U20918 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17979) );
  INV_X1 U20919 ( .A(n17849), .ZN(n17853) );
  NAND2_X1 U20920 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17843), .ZN(n17839) );
  NAND2_X1 U20921 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17835), .ZN(n17834) );
  INV_X1 U20922 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17989) );
  INV_X1 U20923 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17987) );
  AOI22_X1 U20924 ( .A1(n17828), .A2(n17987), .B1(n17930), .B2(n17839), .ZN(
        n17832) );
  OAI22_X1 U20925 ( .A1(n17829), .A2(n17917), .B1(n19564), .B2(n17842), .ZN(
        n17830) );
  AOI21_X1 U20926 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n17859), .A(n17830), .ZN(
        n17831) );
  OAI221_X1 U20927 ( .B1(P3_EAX_REG_22__SCAN_IN), .B2(n17834), .C1(n17989), 
        .C2(n17832), .A(n17831), .ZN(P3_U2713) );
  AOI22_X1 U20928 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17859), .B1(n17927), .B2(
        n17833), .ZN(n17837) );
  OAI211_X1 U20929 ( .C1(n17835), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17930), .B(
        n17834), .ZN(n17836) );
  OAI211_X1 U20930 ( .C1(n17842), .C2(n19558), .A(n17837), .B(n17836), .ZN(
        P3_U2714) );
  AOI22_X1 U20931 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17859), .B1(n17927), .B2(
        n17838), .ZN(n17841) );
  OAI211_X1 U20932 ( .C1(n17843), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17930), .B(
        n17839), .ZN(n17840) );
  OAI211_X1 U20933 ( .C1(n17842), .C2(n19551), .A(n17841), .B(n17840), .ZN(
        P3_U2715) );
  AOI22_X1 U20934 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17859), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17858), .ZN(n17846) );
  INV_X1 U20935 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17983) );
  NAND2_X1 U20936 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17849), .ZN(n17848) );
  AOI211_X1 U20937 ( .C1(n17983), .C2(n17848), .A(n17843), .B(n17921), .ZN(
        n17844) );
  INV_X1 U20938 ( .A(n17844), .ZN(n17845) );
  OAI211_X1 U20939 ( .C1(n17847), .C2(n17917), .A(n17846), .B(n17845), .ZN(
        P3_U2716) );
  AOI22_X1 U20940 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17859), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17858), .ZN(n17851) );
  OAI211_X1 U20941 ( .C1(n17849), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17930), .B(
        n17848), .ZN(n17850) );
  OAI211_X1 U20942 ( .C1(n17852), .C2(n17917), .A(n17851), .B(n17850), .ZN(
        P3_U2717) );
  AOI22_X1 U20943 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17859), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17858), .ZN(n17856) );
  INV_X1 U20944 ( .A(n17860), .ZN(n17854) );
  OAI211_X1 U20945 ( .C1(n17854), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17930), .B(
        n17853), .ZN(n17855) );
  OAI211_X1 U20946 ( .C1(n17857), .C2(n17917), .A(n17856), .B(n17855), .ZN(
        P3_U2718) );
  AOI22_X1 U20947 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17859), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17858), .ZN(n17862) );
  OAI211_X1 U20948 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17867), .A(n17930), .B(
        n17860), .ZN(n17861) );
  OAI211_X1 U20949 ( .C1(n17863), .C2(n17917), .A(n17862), .B(n17861), .ZN(
        P3_U2719) );
  AND2_X1 U20950 ( .A1(n12696), .A2(n17899), .ZN(n17904) );
  AOI22_X1 U20951 ( .A1(n17904), .A2(n17864), .B1(P3_EAX_REG_15__SCAN_IN), 
        .B2(n17930), .ZN(n17866) );
  OAI222_X1 U20952 ( .A1(n17868), .A2(n17920), .B1(n17867), .B2(n17866), .C1(
        n17917), .C2(n17865), .ZN(P3_U2720) );
  NOR2_X1 U20953 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17869), .ZN(n17870) );
  AOI22_X1 U20954 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17928), .B1(n17904), .B2(
        n17870), .ZN(n17873) );
  NAND3_X1 U20955 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17930), .A3(n17871), 
        .ZN(n17872) );
  OAI211_X1 U20956 ( .C1(n17874), .C2(n17917), .A(n17873), .B(n17872), .ZN(
        P3_U2721) );
  INV_X1 U20957 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18025) );
  NAND2_X1 U20958 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17904), .ZN(n17898) );
  NAND2_X1 U20959 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17895), .ZN(n17889) );
  NAND2_X1 U20960 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17886), .ZN(n17878) );
  NAND2_X1 U20961 ( .A1(n17878), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n17877) );
  AOI22_X1 U20962 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17928), .B1(n17927), .B2(
        n17875), .ZN(n17876) );
  OAI221_X1 U20963 ( .B1(n17878), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n17877), 
        .C2(n17921), .A(n17876), .ZN(P3_U2722) );
  INV_X1 U20964 ( .A(n17878), .ZN(n17881) );
  AOI21_X1 U20965 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17930), .A(n17886), .ZN(
        n17880) );
  OAI222_X1 U20966 ( .A1(n17920), .A2(n17882), .B1(n17881), .B2(n17880), .C1(
        n17917), .C2(n17879), .ZN(P3_U2723) );
  INV_X1 U20967 ( .A(n17889), .ZN(n17883) );
  AOI21_X1 U20968 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17930), .A(n17883), .ZN(
        n17885) );
  OAI222_X1 U20969 ( .A1(n17920), .A2(n17887), .B1(n17886), .B2(n17885), .C1(
        n17917), .C2(n17884), .ZN(P3_U2724) );
  AOI22_X1 U20970 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17928), .B1(n17927), .B2(
        n17888), .ZN(n17891) );
  OAI211_X1 U20971 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17895), .A(n17930), .B(
        n17889), .ZN(n17890) );
  NAND2_X1 U20972 ( .A1(n17891), .A2(n17890), .ZN(P3_U2725) );
  INV_X1 U20973 ( .A(n17898), .ZN(n17892) );
  AOI21_X1 U20974 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17930), .A(n17892), .ZN(
        n17894) );
  OAI222_X1 U20975 ( .A1(n17920), .A2(n17896), .B1(n17895), .B2(n17894), .C1(
        n17917), .C2(n17893), .ZN(P3_U2726) );
  AOI22_X1 U20976 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17928), .B1(n17927), .B2(
        n17897), .ZN(n17901) );
  OAI211_X1 U20977 ( .C1(n17899), .C2(P3_EAX_REG_8__SCAN_IN), .A(n17930), .B(
        n17898), .ZN(n17900) );
  NAND2_X1 U20978 ( .A1(n17901), .A2(n17900), .ZN(P3_U2727) );
  INV_X1 U20979 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18019) );
  INV_X1 U20980 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18013) );
  INV_X1 U20981 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18011) );
  NAND3_X1 U20982 ( .A1(n12696), .A2(n9660), .A3(P3_EAX_REG_1__SCAN_IN), .ZN(
        n17929) );
  NOR2_X1 U20983 ( .A1(n18011), .A2(n17929), .ZN(n17915) );
  INV_X1 U20984 ( .A(n17915), .ZN(n17924) );
  NAND2_X1 U20985 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17914), .ZN(n17905) );
  NOR2_X1 U20986 ( .A1(n18019), .A2(n17905), .ZN(n17908) );
  AOI21_X1 U20987 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17930), .A(n17908), .ZN(
        n17903) );
  OAI222_X1 U20988 ( .A1(n17920), .A2(n21237), .B1(n17904), .B2(n17903), .C1(
        n17917), .C2(n17902), .ZN(P3_U2728) );
  INV_X1 U20989 ( .A(n17905), .ZN(n17911) );
  AOI21_X1 U20990 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17930), .A(n17911), .ZN(
        n17907) );
  OAI222_X1 U20991 ( .A1(n18751), .A2(n17920), .B1(n17908), .B2(n17907), .C1(
        n17917), .C2(n17906), .ZN(P3_U2729) );
  AOI21_X1 U20992 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17930), .A(n17914), .ZN(
        n17910) );
  OAI222_X1 U20993 ( .A1(n18746), .A2(n17920), .B1(n17911), .B2(n17910), .C1(
        n17917), .C2(n17909), .ZN(P3_U2730) );
  AOI21_X1 U20994 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17930), .A(n17919), .ZN(
        n17913) );
  OAI222_X1 U20995 ( .A1(n18741), .A2(n17920), .B1(n17914), .B2(n17913), .C1(
        n17917), .C2(n17912), .ZN(P3_U2731) );
  AOI21_X1 U20996 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17930), .A(n17915), .ZN(
        n17918) );
  OAI222_X1 U20997 ( .A1(n18737), .A2(n17920), .B1(n17919), .B2(n17918), .C1(
        n17917), .C2(n17916), .ZN(P3_U2732) );
  OAI21_X1 U20998 ( .B1(n18011), .B2(n17921), .A(n17929), .ZN(n17923) );
  AOI222_X1 U20999 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17928), .B1(n17924), .B2(
        n17923), .C1(n17927), .C2(n17922), .ZN(n17925) );
  INV_X1 U21000 ( .A(n17925), .ZN(P3_U2733) );
  AOI22_X1 U21001 ( .A1(n17928), .A2(BUF2_REG_1__SCAN_IN), .B1(n17927), .B2(
        n17926), .ZN(n17932) );
  OAI211_X1 U21002 ( .C1(n9660), .C2(P3_EAX_REG_1__SCAN_IN), .A(n17930), .B(
        n17929), .ZN(n17931) );
  NAND2_X1 U21003 ( .A1(n17932), .A2(n17931), .ZN(P3_U2734) );
  NOR2_X1 U21004 ( .A1(n17950), .A2(n17934), .ZN(P3_U2736) );
  INV_X1 U21005 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n21224) );
  NOR2_X1 U21006 ( .A1(n18721), .A2(n17970), .ZN(n17936) );
  INV_X2 U21007 ( .A(n19354), .ZN(n19217) );
  AOI22_X1 U21008 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17936), .B1(n19217), 
        .B2(P3_UWORD_REG_14__SCAN_IN), .ZN(n17935) );
  OAI21_X1 U21009 ( .B1(n21224), .B2(n17950), .A(n17935), .ZN(P3_U2737) );
  AOI22_X1 U21010 ( .A1(n19217), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17937) );
  OAI21_X1 U21011 ( .B1(n18003), .B2(n17952), .A(n17937), .ZN(P3_U2738) );
  INV_X1 U21012 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18001) );
  AOI22_X1 U21013 ( .A1(n19217), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17938) );
  OAI21_X1 U21014 ( .B1(n18001), .B2(n17952), .A(n17938), .ZN(P3_U2739) );
  AOI22_X1 U21015 ( .A1(n19217), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17939) );
  OAI21_X1 U21016 ( .B1(n17999), .B2(n17952), .A(n17939), .ZN(P3_U2740) );
  INV_X1 U21017 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17997) );
  AOI22_X1 U21018 ( .A1(n19217), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17940) );
  OAI21_X1 U21019 ( .B1(n17997), .B2(n17952), .A(n17940), .ZN(P3_U2741) );
  AOI22_X1 U21020 ( .A1(n19217), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17941) );
  OAI21_X1 U21021 ( .B1(n17995), .B2(n17952), .A(n17941), .ZN(P3_U2742) );
  INV_X1 U21022 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17993) );
  AOI22_X1 U21023 ( .A1(n19217), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17942) );
  OAI21_X1 U21024 ( .B1(n17993), .B2(n17952), .A(n17942), .ZN(P3_U2743) );
  INV_X1 U21025 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17991) );
  AOI22_X1 U21026 ( .A1(n19217), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17943) );
  OAI21_X1 U21027 ( .B1(n17991), .B2(n17952), .A(n17943), .ZN(P3_U2744) );
  AOI22_X1 U21028 ( .A1(n19217), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17944) );
  OAI21_X1 U21029 ( .B1(n17989), .B2(n17952), .A(n17944), .ZN(P3_U2745) );
  AOI22_X1 U21030 ( .A1(n19217), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17945) );
  OAI21_X1 U21031 ( .B1(n17987), .B2(n17952), .A(n17945), .ZN(P3_U2746) );
  INV_X1 U21032 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17985) );
  AOI22_X1 U21033 ( .A1(n19217), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17946) );
  OAI21_X1 U21034 ( .B1(n17985), .B2(n17952), .A(n17946), .ZN(P3_U2747) );
  AOI22_X1 U21035 ( .A1(n19217), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17947) );
  OAI21_X1 U21036 ( .B1(n17983), .B2(n17952), .A(n17947), .ZN(P3_U2748) );
  INV_X1 U21037 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17981) );
  AOI22_X1 U21038 ( .A1(n19217), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17948) );
  OAI21_X1 U21039 ( .B1(n17981), .B2(n17952), .A(n17948), .ZN(P3_U2749) );
  INV_X1 U21040 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n21293) );
  INV_X1 U21041 ( .A(P3_UWORD_REG_1__SCAN_IN), .ZN(n17949) );
  OAI222_X1 U21042 ( .A1(n17950), .A2(n21293), .B1(n17952), .B2(n17979), .C1(
        n19354), .C2(n17949), .ZN(P3_U2750) );
  INV_X1 U21043 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17977) );
  AOI22_X1 U21044 ( .A1(n19217), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17951) );
  OAI21_X1 U21045 ( .B1(n17977), .B2(n17952), .A(n17951), .ZN(P3_U2751) );
  AOI22_X1 U21046 ( .A1(n19217), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17953) );
  OAI21_X1 U21047 ( .B1(n18042), .B2(n17970), .A(n17953), .ZN(P3_U2752) );
  AOI22_X1 U21048 ( .A1(n19217), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17954) );
  OAI21_X1 U21049 ( .B1(n18037), .B2(n17970), .A(n17954), .ZN(P3_U2753) );
  AOI22_X1 U21050 ( .A1(n19217), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17955) );
  OAI21_X1 U21051 ( .B1(n18035), .B2(n17970), .A(n17955), .ZN(P3_U2754) );
  AOI22_X1 U21052 ( .A1(n19217), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17956) );
  OAI21_X1 U21053 ( .B1(n18033), .B2(n17970), .A(n17956), .ZN(P3_U2755) );
  AOI22_X1 U21054 ( .A1(n19217), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17957) );
  OAI21_X1 U21055 ( .B1(n18029), .B2(n17970), .A(n17957), .ZN(P3_U2756) );
  AOI22_X1 U21056 ( .A1(n19217), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17958) );
  OAI21_X1 U21057 ( .B1(n18027), .B2(n17970), .A(n17958), .ZN(P3_U2757) );
  AOI22_X1 U21058 ( .A1(n19217), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17959) );
  OAI21_X1 U21059 ( .B1(n18025), .B2(n17970), .A(n17959), .ZN(P3_U2758) );
  INV_X1 U21060 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18023) );
  AOI22_X1 U21061 ( .A1(n19217), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17960) );
  OAI21_X1 U21062 ( .B1(n18023), .B2(n17970), .A(n17960), .ZN(P3_U2759) );
  INV_X1 U21063 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18021) );
  AOI22_X1 U21064 ( .A1(n19217), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17961) );
  OAI21_X1 U21065 ( .B1(n18021), .B2(n17970), .A(n17961), .ZN(P3_U2760) );
  AOI22_X1 U21066 ( .A1(n19217), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17962) );
  OAI21_X1 U21067 ( .B1(n18019), .B2(n17970), .A(n17962), .ZN(P3_U2761) );
  INV_X1 U21068 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18017) );
  AOI22_X1 U21069 ( .A1(n19217), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17964) );
  OAI21_X1 U21070 ( .B1(n18017), .B2(n17970), .A(n17964), .ZN(P3_U2762) );
  INV_X1 U21071 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18015) );
  AOI22_X1 U21072 ( .A1(n19217), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17965) );
  OAI21_X1 U21073 ( .B1(n18015), .B2(n17970), .A(n17965), .ZN(P3_U2763) );
  AOI22_X1 U21074 ( .A1(n19217), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17966) );
  OAI21_X1 U21075 ( .B1(n18013), .B2(n17970), .A(n17966), .ZN(P3_U2764) );
  AOI22_X1 U21076 ( .A1(n19217), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17967) );
  OAI21_X1 U21077 ( .B1(n18011), .B2(n17970), .A(n17967), .ZN(P3_U2765) );
  INV_X1 U21078 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18009) );
  AOI22_X1 U21079 ( .A1(n19217), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17968) );
  OAI21_X1 U21080 ( .B1(n18009), .B2(n17970), .A(n17968), .ZN(P3_U2766) );
  INV_X1 U21081 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18007) );
  AOI22_X1 U21082 ( .A1(n19217), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17963), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17969) );
  OAI21_X1 U21083 ( .B1(n18007), .B2(n17970), .A(n17969), .ZN(P3_U2767) );
  NOR2_X1 U21084 ( .A1(n17972), .A2(n17973), .ZN(n19205) );
  NAND2_X2 U21085 ( .A1(n17974), .A2(n19205), .ZN(n18041) );
  INV_X1 U21086 ( .A(n17973), .ZN(n17975) );
  AOI22_X1 U21087 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18039), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18030), .ZN(n17976) );
  OAI21_X1 U21088 ( .B1(n17977), .B2(n18041), .A(n17976), .ZN(P3_U2768) );
  AOI22_X1 U21089 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18039), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18030), .ZN(n17978) );
  OAI21_X1 U21090 ( .B1(n17979), .B2(n18041), .A(n17978), .ZN(P3_U2769) );
  AOI22_X1 U21091 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18039), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18030), .ZN(n17980) );
  OAI21_X1 U21092 ( .B1(n17981), .B2(n18041), .A(n17980), .ZN(P3_U2770) );
  AOI22_X1 U21093 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18039), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18030), .ZN(n17982) );
  OAI21_X1 U21094 ( .B1(n17983), .B2(n18041), .A(n17982), .ZN(P3_U2771) );
  AOI22_X1 U21095 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18031), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18030), .ZN(n17984) );
  OAI21_X1 U21096 ( .B1(n17985), .B2(n18041), .A(n17984), .ZN(P3_U2772) );
  AOI22_X1 U21097 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18031), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18030), .ZN(n17986) );
  OAI21_X1 U21098 ( .B1(n17987), .B2(n18041), .A(n17986), .ZN(P3_U2773) );
  AOI22_X1 U21099 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18031), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18030), .ZN(n17988) );
  OAI21_X1 U21100 ( .B1(n17989), .B2(n18041), .A(n17988), .ZN(P3_U2774) );
  AOI22_X1 U21101 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18031), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18030), .ZN(n17990) );
  OAI21_X1 U21102 ( .B1(n17991), .B2(n18041), .A(n17990), .ZN(P3_U2775) );
  AOI22_X1 U21103 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18031), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18030), .ZN(n17992) );
  OAI21_X1 U21104 ( .B1(n17993), .B2(n18041), .A(n17992), .ZN(P3_U2776) );
  AOI22_X1 U21105 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18031), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18030), .ZN(n17994) );
  OAI21_X1 U21106 ( .B1(n17995), .B2(n18041), .A(n17994), .ZN(P3_U2777) );
  AOI22_X1 U21107 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18031), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18030), .ZN(n17996) );
  OAI21_X1 U21108 ( .B1(n17997), .B2(n18041), .A(n17996), .ZN(P3_U2778) );
  AOI22_X1 U21109 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18031), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18030), .ZN(n17998) );
  OAI21_X1 U21110 ( .B1(n17999), .B2(n18041), .A(n17998), .ZN(P3_U2779) );
  AOI22_X1 U21111 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18039), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18030), .ZN(n18000) );
  OAI21_X1 U21112 ( .B1(n18001), .B2(n18041), .A(n18000), .ZN(P3_U2780) );
  AOI22_X1 U21113 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18039), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18030), .ZN(n18002) );
  OAI21_X1 U21114 ( .B1(n18003), .B2(n18041), .A(n18002), .ZN(P3_U2781) );
  INV_X1 U21115 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18005) );
  AOI22_X1 U21116 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18039), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18030), .ZN(n18004) );
  OAI21_X1 U21117 ( .B1(n18005), .B2(n18041), .A(n18004), .ZN(P3_U2782) );
  AOI22_X1 U21118 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18039), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18030), .ZN(n18006) );
  OAI21_X1 U21119 ( .B1(n18007), .B2(n18041), .A(n18006), .ZN(P3_U2783) );
  AOI22_X1 U21120 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18039), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18030), .ZN(n18008) );
  OAI21_X1 U21121 ( .B1(n18009), .B2(n18041), .A(n18008), .ZN(P3_U2784) );
  AOI22_X1 U21122 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18039), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18030), .ZN(n18010) );
  OAI21_X1 U21123 ( .B1(n18011), .B2(n18041), .A(n18010), .ZN(P3_U2785) );
  AOI22_X1 U21124 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18039), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18030), .ZN(n18012) );
  OAI21_X1 U21125 ( .B1(n18013), .B2(n18041), .A(n18012), .ZN(P3_U2786) );
  AOI22_X1 U21126 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18039), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18038), .ZN(n18014) );
  OAI21_X1 U21127 ( .B1(n18015), .B2(n18041), .A(n18014), .ZN(P3_U2787) );
  AOI22_X1 U21128 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18039), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18038), .ZN(n18016) );
  OAI21_X1 U21129 ( .B1(n18017), .B2(n18041), .A(n18016), .ZN(P3_U2788) );
  AOI22_X1 U21130 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18039), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18038), .ZN(n18018) );
  OAI21_X1 U21131 ( .B1(n18019), .B2(n18041), .A(n18018), .ZN(P3_U2789) );
  AOI22_X1 U21132 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18039), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18038), .ZN(n18020) );
  OAI21_X1 U21133 ( .B1(n18021), .B2(n18041), .A(n18020), .ZN(P3_U2790) );
  AOI22_X1 U21134 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18039), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18038), .ZN(n18022) );
  OAI21_X1 U21135 ( .B1(n18023), .B2(n18041), .A(n18022), .ZN(P3_U2791) );
  AOI22_X1 U21136 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18031), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18038), .ZN(n18024) );
  OAI21_X1 U21137 ( .B1(n18025), .B2(n18041), .A(n18024), .ZN(P3_U2792) );
  AOI22_X1 U21138 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18031), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18030), .ZN(n18026) );
  OAI21_X1 U21139 ( .B1(n18027), .B2(n18041), .A(n18026), .ZN(P3_U2793) );
  AOI22_X1 U21140 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18039), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18038), .ZN(n18028) );
  OAI21_X1 U21141 ( .B1(n18029), .B2(n18041), .A(n18028), .ZN(P3_U2794) );
  AOI22_X1 U21142 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18031), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18030), .ZN(n18032) );
  OAI21_X1 U21143 ( .B1(n18033), .B2(n18041), .A(n18032), .ZN(P3_U2795) );
  AOI22_X1 U21144 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18039), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18038), .ZN(n18034) );
  OAI21_X1 U21145 ( .B1(n18035), .B2(n18041), .A(n18034), .ZN(P3_U2796) );
  AOI22_X1 U21146 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18039), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18038), .ZN(n18036) );
  OAI21_X1 U21147 ( .B1(n18037), .B2(n18041), .A(n18036), .ZN(P3_U2797) );
  AOI22_X1 U21148 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18039), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18038), .ZN(n18040) );
  OAI21_X1 U21149 ( .B1(n18042), .B2(n18041), .A(n18040), .ZN(P3_U2798) );
  AOI22_X1 U21150 ( .A1(n18140), .A2(n18044), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18043), .ZN(n18053) );
  NAND2_X1 U21151 ( .A1(n18045), .A2(n13037), .ZN(n18046) );
  XNOR2_X1 U21152 ( .A(n18046), .B(n10304), .ZN(n18399) );
  INV_X1 U21153 ( .A(n18408), .ZN(n18411) );
  NAND3_X1 U21154 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18411), .A3(
        n18407), .ZN(n18400) );
  INV_X1 U21155 ( .A(n18169), .ZN(n18058) );
  AOI21_X1 U21156 ( .B1(n18054), .B2(n19036), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18055) );
  NAND2_X1 U21157 ( .A1(n18695), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18405) );
  OAI21_X1 U21158 ( .B1(n18056), .B2(n18055), .A(n18405), .ZN(n18057) );
  AOI221_X1 U21159 ( .B1(n18140), .B2(n18059), .C1(n18058), .C2(n18059), .A(
        n18057), .ZN(n18064) );
  OAI21_X1 U21160 ( .B1(n18060), .B2(n18407), .A(n18061), .ZN(n18402) );
  AOI22_X1 U21161 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18062), .B1(
        n18293), .B2(n18402), .ZN(n18063) );
  OAI211_X1 U21162 ( .C1(n18103), .C2(n18400), .A(n18064), .B(n18063), .ZN(
        P3_U2804) );
  OAI21_X1 U21163 ( .B1(n18065), .B2(n18380), .A(n18381), .ZN(n18066) );
  AOI21_X1 U21164 ( .B1(n19036), .B2(n12597), .A(n18066), .ZN(n18093) );
  OAI21_X1 U21165 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18169), .A(
        n18093), .ZN(n18084) );
  AOI22_X1 U21166 ( .A1(n18140), .A2(n18067), .B1(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18084), .ZN(n18079) );
  XNOR2_X1 U21167 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n18068), .ZN(
        n18421) );
  XNOR2_X1 U21168 ( .A(n18069), .B(n18413), .ZN(n18423) );
  INV_X1 U21169 ( .A(n18070), .ZN(n18072) );
  OAI21_X1 U21170 ( .B1(n10304), .B2(n18072), .A(n18071), .ZN(n18073) );
  XNOR2_X1 U21171 ( .A(n18073), .B(n18413), .ZN(n18419) );
  OAI22_X1 U21172 ( .A1(n10295), .A2(n18423), .B1(n18248), .B2(n18419), .ZN(
        n18074) );
  AOI21_X1 U21173 ( .B1(n18371), .B2(n18421), .A(n18074), .ZN(n18078) );
  NAND2_X1 U21174 ( .A1(n18695), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18417) );
  INV_X1 U21175 ( .A(n18075), .ZN(n18221) );
  NOR2_X1 U21176 ( .A1(n18221), .A2(n12597), .ZN(n18086) );
  OAI211_X1 U21177 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n18086), .B(n18076), .ZN(n18077) );
  NAND4_X1 U21178 ( .A1(n18079), .A2(n18078), .A3(n18417), .A4(n18077), .ZN(
        P3_U2805) );
  INV_X1 U21179 ( .A(n18174), .ZN(n18188) );
  OR2_X1 U21180 ( .A1(n18080), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18439) );
  AOI22_X1 U21181 ( .A1(n18695), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18140), 
        .B2(n18081), .ZN(n18082) );
  INV_X1 U21182 ( .A(n18082), .ZN(n18083) );
  AOI221_X1 U21183 ( .B1(n18086), .B2(n18085), .C1(n18084), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18083), .ZN(n18089) );
  OAI22_X1 U21184 ( .A1(n18428), .A2(n10295), .B1(n18427), .B2(n18385), .ZN(
        n18100) );
  OAI21_X1 U21185 ( .B1(n18087), .B2(n18433), .A(n18070), .ZN(n18437) );
  AOI22_X1 U21186 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18100), .B1(
        n18293), .B2(n18437), .ZN(n18088) );
  OAI211_X1 U21187 ( .C1(n18188), .C2(n18439), .A(n18089), .B(n18088), .ZN(
        P3_U2806) );
  NOR2_X1 U21188 ( .A1(n18701), .A2(n19281), .ZN(n18443) );
  AOI21_X1 U21189 ( .B1(n12600), .B2(n19036), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18092) );
  OR2_X1 U21190 ( .A1(n18169), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18090) );
  OAI22_X1 U21191 ( .A1(n18093), .A2(n18092), .B1(n18091), .B2(n18090), .ZN(
        n18094) );
  AOI211_X1 U21192 ( .C1(n18095), .C2(n18140), .A(n18443), .B(n18094), .ZN(
        n18102) );
  OAI22_X1 U21193 ( .A1(n18096), .A2(n18104), .B1(n10304), .B2(n18117), .ZN(
        n18097) );
  NOR2_X1 U21194 ( .A1(n18097), .A2(n18133), .ZN(n18099) );
  XNOR2_X1 U21195 ( .A(n18099), .B(n18098), .ZN(n18444) );
  AOI22_X1 U21196 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18100), .B1(
        n18293), .B2(n18444), .ZN(n18101) );
  OAI211_X1 U21197 ( .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n18103), .A(
        n18102), .B(n18101), .ZN(P3_U2807) );
  INV_X1 U21198 ( .A(n18104), .ZN(n18105) );
  XNOR2_X1 U21199 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n18106), .ZN(
        n18460) );
  NOR2_X1 U21200 ( .A1(n18453), .A2(n18188), .ZN(n18118) );
  INV_X1 U21201 ( .A(n18453), .ZN(n18107) );
  AOI22_X1 U21202 ( .A1(n18294), .A2(n18514), .B1(n18371), .B2(n18523), .ZN(
        n18187) );
  OAI21_X1 U21203 ( .B1(n18107), .B2(n18142), .A(n18187), .ZN(n18130) );
  INV_X1 U21204 ( .A(n18381), .ZN(n18368) );
  AOI21_X1 U21205 ( .B1(n18108), .B2(n18334), .A(n18368), .ZN(n18109) );
  INV_X1 U21206 ( .A(n18109), .ZN(n18110) );
  AOI21_X1 U21207 ( .B1(n18219), .B2(n18111), .A(n18110), .ZN(n18137) );
  OAI21_X1 U21208 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18169), .A(
        n18137), .ZN(n18127) );
  AOI22_X1 U21209 ( .A1(n18140), .A2(n18112), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18127), .ZN(n18115) );
  NOR2_X1 U21210 ( .A1(n18221), .A2(n18108), .ZN(n18129) );
  OAI211_X1 U21211 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n18129), .B(n18113), .ZN(n18114) );
  OAI211_X1 U21212 ( .C1(n19279), .C2(n18701), .A(n18115), .B(n18114), .ZN(
        n18116) );
  AOI221_X1 U21213 ( .B1(n18118), .B2(n18117), .C1(n18130), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n18116), .ZN(n18119) );
  OAI21_X1 U21214 ( .B1(n18248), .B2(n18460), .A(n18119), .ZN(P3_U2808) );
  NAND3_X1 U21215 ( .A1(n10304), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n18120), .ZN(n18145) );
  INV_X1 U21216 ( .A(n18121), .ZN(n18146) );
  OAI22_X1 U21217 ( .A1(n18464), .A2(n18145), .B1(n18146), .B2(n18122), .ZN(
        n18123) );
  XNOR2_X1 U21218 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18123), .ZN(
        n18469) );
  AOI22_X1 U21219 ( .A1(n18695), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18140), 
        .B2(n18124), .ZN(n18125) );
  INV_X1 U21220 ( .A(n18125), .ZN(n18126) );
  AOI221_X1 U21221 ( .B1(n18129), .B2(n18128), .C1(n18127), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18126), .ZN(n18132) );
  NAND2_X1 U21222 ( .A1(n18161), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18461) );
  NOR3_X1 U21223 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18464), .A3(
        n18461), .ZN(n18468) );
  AOI22_X1 U21224 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18130), .B1(
        n18174), .B2(n18468), .ZN(n18131) );
  OAI211_X1 U21225 ( .C1(n18469), .C2(n18248), .A(n18132), .B(n18131), .ZN(
        P3_U2809) );
  INV_X1 U21226 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18141) );
  XNOR2_X1 U21227 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n18134), .ZN(
        n18477) );
  AOI21_X1 U21228 ( .B1(n18135), .B2(n19036), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18136) );
  OAI22_X1 U21229 ( .A1(n18137), .A2(n18136), .B1(n18701), .B2(n19275), .ZN(
        n18138) );
  AOI221_X1 U21230 ( .B1(n18140), .B2(n18139), .C1(n18058), .C2(n18139), .A(
        n18138), .ZN(n18144) );
  NOR2_X1 U21231 ( .A1(n18141), .A2(n18461), .ZN(n18448) );
  OAI21_X1 U21232 ( .B1(n18142), .B2(n18448), .A(n18187), .ZN(n18153) );
  INV_X1 U21233 ( .A(n18448), .ZN(n18472) );
  NOR2_X1 U21234 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18472), .ZN(
        n18470) );
  AOI22_X1 U21235 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18153), .B1(
        n18174), .B2(n18470), .ZN(n18143) );
  OAI211_X1 U21236 ( .C1(n18248), .C2(n18477), .A(n18144), .B(n18143), .ZN(
        P3_U2810) );
  OAI21_X1 U21237 ( .B1(n18162), .B2(n18146), .A(n18145), .ZN(n18147) );
  XNOR2_X1 U21238 ( .A(n18147), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18483) );
  OAI21_X1 U21239 ( .B1(n18368), .B2(n12602), .A(n18374), .ZN(n18170) );
  OAI21_X1 U21240 ( .B1(n18148), .B2(n18380), .A(n18170), .ZN(n18158) );
  NOR2_X1 U21241 ( .A1(n18221), .A2(n12602), .ZN(n18160) );
  OAI211_X1 U21242 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18160), .B(n18149), .ZN(n18150) );
  NAND2_X1 U21243 ( .A1(n18695), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18481) );
  OAI211_X1 U21244 ( .C1(n18239), .C2(n18151), .A(n18150), .B(n18481), .ZN(
        n18152) );
  AOI21_X1 U21245 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18158), .A(
        n18152), .ZN(n18155) );
  NOR2_X1 U21246 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18461), .ZN(
        n18478) );
  AOI22_X1 U21247 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18153), .B1(
        n18174), .B2(n18478), .ZN(n18154) );
  OAI211_X1 U21248 ( .C1(n18483), .C2(n18248), .A(n18155), .B(n18154), .ZN(
        P3_U2811) );
  NAND2_X1 U21249 ( .A1(n18161), .A2(n18163), .ZN(n18496) );
  OAI22_X1 U21250 ( .A1(n18701), .A2(n19271), .B1(n18239), .B2(n18156), .ZN(
        n18157) );
  AOI221_X1 U21251 ( .B1(n18160), .B2(n18159), .C1(n18158), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n18157), .ZN(n18166) );
  OAI21_X1 U21252 ( .B1(n18161), .B2(n18188), .A(n18187), .ZN(n18175) );
  OAI21_X1 U21253 ( .B1(n18228), .B2(n18163), .A(n18162), .ZN(n18164) );
  XNOR2_X1 U21254 ( .A(n18164), .B(n18121), .ZN(n18492) );
  AOI22_X1 U21255 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18175), .B1(
        n18293), .B2(n18492), .ZN(n18165) );
  OAI211_X1 U21256 ( .C1(n18188), .C2(n18496), .A(n18166), .B(n18165), .ZN(
        P3_U2812) );
  AOI21_X1 U21257 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18168), .A(
        n18167), .ZN(n18503) );
  AOI21_X1 U21258 ( .B1(n9791), .B2(n19036), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18171) );
  OAI22_X1 U21259 ( .A1(n18171), .A2(n18170), .B1(n18701), .B2(n19270), .ZN(
        n18172) );
  AOI21_X1 U21260 ( .B1(n18173), .B2(n18343), .A(n18172), .ZN(n18177) );
  NOR2_X1 U21261 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18512), .ZN(
        n18499) );
  AOI22_X1 U21262 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18175), .B1(
        n18174), .B2(n18499), .ZN(n18176) );
  OAI211_X1 U21263 ( .C1(n18503), .C2(n18248), .A(n18177), .B(n18176), .ZN(
        P3_U2813) );
  NOR2_X1 U21264 ( .A1(n18228), .A2(n12890), .ZN(n18266) );
  AOI22_X1 U21265 ( .A1(n18266), .A2(n10179), .B1(n18178), .B2(n18228), .ZN(
        n18179) );
  XNOR2_X1 U21266 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n18179), .ZN(
        n18509) );
  AOI21_X1 U21267 ( .B1(n18334), .B2(n12607), .A(n18368), .ZN(n18207) );
  OAI21_X1 U21268 ( .B1(n18180), .B2(n18380), .A(n18207), .ZN(n18192) );
  AOI22_X1 U21269 ( .A1(n18695), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18192), .ZN(n18183) );
  NOR2_X1 U21270 ( .A1(n18221), .A2(n12607), .ZN(n18194) );
  OAI211_X1 U21271 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18194), .B(n18181), .ZN(n18182) );
  OAI211_X1 U21272 ( .C1(n18239), .C2(n18184), .A(n18183), .B(n18182), .ZN(
        n18185) );
  AOI21_X1 U21273 ( .B1(n18293), .B2(n18509), .A(n18185), .ZN(n18186) );
  OAI221_X1 U21274 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18188), 
        .C1(n18512), .C2(n18187), .A(n18186), .ZN(P3_U2814) );
  NOR2_X1 U21275 ( .A1(n18189), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18519) );
  NAND2_X1 U21276 ( .A1(n18294), .A2(n18514), .ZN(n18203) );
  OAI22_X1 U21277 ( .A1(n18701), .A2(n19265), .B1(n18239), .B2(n18190), .ZN(
        n18191) );
  AOI221_X1 U21278 ( .B1(n18194), .B2(n18193), .C1(n18192), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18191), .ZN(n18202) );
  NAND2_X1 U21279 ( .A1(n12865), .A2(n18228), .ZN(n18274) );
  NOR3_X1 U21280 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18255), .A3(
        n18274), .ZN(n18234) );
  INV_X1 U21281 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18216) );
  NOR3_X1 U21282 ( .A1(n18562), .A2(n18196), .A3(n18195), .ZN(n18198) );
  AOI22_X1 U21283 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18228), .B1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18561), .ZN(n18197) );
  OAI221_X1 U21284 ( .B1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n18234), 
        .C1(n18216), .C2(n18198), .A(n18197), .ZN(n18199) );
  XNOR2_X1 U21285 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18199), .ZN(
        n18520) );
  AND2_X1 U21286 ( .A1(n18523), .A2(n18371), .ZN(n18200) );
  NAND4_X1 U21287 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18558), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(n18544), .ZN(n18211) );
  NAND2_X1 U21288 ( .A1(n9996), .A2(n18211), .ZN(n18522) );
  AOI22_X1 U21289 ( .A1(n18293), .A2(n18520), .B1(n18200), .B2(n18522), .ZN(
        n18201) );
  OAI211_X1 U21290 ( .C1(n18519), .C2(n18203), .A(n18202), .B(n18201), .ZN(
        P3_U2815) );
  AND2_X1 U21291 ( .A1(n18204), .A2(n18558), .ZN(n18550) );
  OAI221_X1 U21292 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18550), .A(n18205), .ZN(
        n18540) );
  AOI21_X1 U21293 ( .B1(n17287), .B2(n19036), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18206) );
  OAI22_X1 U21294 ( .A1(n18207), .A2(n18206), .B1(n18701), .B2(n19263), .ZN(
        n18213) );
  INV_X1 U21295 ( .A(n18266), .ZN(n18273) );
  NAND2_X1 U21296 ( .A1(n18208), .A2(n18561), .ZN(n18209) );
  OAI22_X1 U21297 ( .A1(n18528), .A2(n18273), .B1(n18274), .B2(n18209), .ZN(
        n18210) );
  XNOR2_X1 U21298 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18210), .ZN(
        n18536) );
  NAND2_X1 U21299 ( .A1(n18558), .A2(n18544), .ZN(n18552) );
  INV_X1 U21300 ( .A(n18552), .ZN(n18227) );
  OAI221_X1 U21301 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18227), .A(n18211), .ZN(
        n18535) );
  OAI22_X1 U21302 ( .A1(n18536), .A2(n18248), .B1(n18385), .B2(n18535), .ZN(
        n18212) );
  AOI211_X1 U21303 ( .C1(n18214), .C2(n18343), .A(n18213), .B(n18212), .ZN(
        n18215) );
  OAI21_X1 U21304 ( .B1(n10295), .B2(n18540), .A(n18215), .ZN(P3_U2816) );
  NAND2_X1 U21305 ( .A1(n18558), .A2(n18216), .ZN(n18557) );
  AOI22_X1 U21306 ( .A1(n18334), .A2(n18217), .B1(n18219), .B2(n18218), .ZN(
        n18220) );
  NAND2_X1 U21307 ( .A1(n18220), .A2(n18381), .ZN(n18241) );
  NOR2_X1 U21308 ( .A1(n18221), .A2(n18217), .ZN(n18243) );
  OAI211_X1 U21309 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18243), .B(n18222), .ZN(n18224) );
  NAND2_X1 U21310 ( .A1(n18695), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n18223) );
  OAI211_X1 U21311 ( .C1(n18239), .C2(n18225), .A(n18224), .B(n18223), .ZN(
        n18226) );
  AOI21_X1 U21312 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18241), .A(
        n18226), .ZN(n18233) );
  OAI22_X1 U21313 ( .A1(n18227), .A2(n18385), .B1(n18550), .B2(n10295), .ZN(
        n18244) );
  NOR2_X1 U21314 ( .A1(n18562), .A2(n18195), .ZN(n18230) );
  NOR2_X1 U21315 ( .A1(n18228), .A2(n18561), .ZN(n18229) );
  OAI22_X1 U21316 ( .A1(n18230), .A2(n18561), .B1(n18234), .B2(n18229), .ZN(
        n18231) );
  XNOR2_X1 U21317 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18231), .ZN(
        n18545) );
  AOI22_X1 U21318 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18244), .B1(
        n18293), .B2(n18545), .ZN(n18232) );
  OAI211_X1 U21319 ( .C1(n18283), .C2(n18557), .A(n18233), .B(n18232), .ZN(
        P3_U2817) );
  INV_X1 U21320 ( .A(n18562), .ZN(n18235) );
  AOI21_X1 U21321 ( .B1(n18266), .B2(n18235), .A(n18234), .ZN(n18236) );
  XNOR2_X1 U21322 ( .A(n18236), .B(n18561), .ZN(n18568) );
  INV_X1 U21323 ( .A(n18237), .ZN(n18238) );
  OAI22_X1 U21324 ( .A1(n18701), .A2(n19260), .B1(n18239), .B2(n18238), .ZN(
        n18240) );
  AOI221_X1 U21325 ( .B1(n18243), .B2(n18242), .C1(n18241), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n18240), .ZN(n18247) );
  OAI21_X1 U21326 ( .B1(n18562), .B2(n18283), .A(n18561), .ZN(n18245) );
  NAND2_X1 U21327 ( .A1(n18245), .A2(n18244), .ZN(n18246) );
  OAI211_X1 U21328 ( .C1(n18568), .C2(n18248), .A(n18247), .B(n18246), .ZN(
        P3_U2818) );
  INV_X1 U21329 ( .A(n18265), .ZN(n18577) );
  OR2_X1 U21330 ( .A1(n18577), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18582) );
  INV_X1 U21331 ( .A(n18249), .ZN(n18254) );
  INV_X1 U21332 ( .A(n18286), .ZN(n18287) );
  NOR2_X1 U21333 ( .A1(n18287), .A2(n19061), .ZN(n18299) );
  NAND3_X1 U21334 ( .A1(n18286), .A2(n17327), .A3(n19036), .ZN(n18259) );
  NOR2_X1 U21335 ( .A1(n18250), .A2(n18259), .ZN(n18272) );
  AOI21_X1 U21336 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18374), .A(
        n18272), .ZN(n18251) );
  AOI21_X1 U21337 ( .B1(n18299), .B2(n18252), .A(n18251), .ZN(n18253) );
  INV_X1 U21338 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19259) );
  NOR2_X1 U21339 ( .A1(n18701), .A2(n19259), .ZN(n18569) );
  AOI211_X1 U21340 ( .C1(n18254), .C2(n18343), .A(n18253), .B(n18569), .ZN(
        n18258) );
  INV_X1 U21341 ( .A(n18544), .ZN(n18572) );
  AOI22_X1 U21342 ( .A1(n18294), .A2(n12890), .B1(n18371), .B2(n18572), .ZN(
        n18282) );
  OAI21_X1 U21343 ( .B1(n18265), .B2(n18283), .A(n18282), .ZN(n18267) );
  OAI22_X1 U21344 ( .A1(n18577), .A2(n18273), .B1(n18255), .B2(n18274), .ZN(
        n18256) );
  XOR2_X1 U21345 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18256), .Z(
        n18570) );
  AOI22_X1 U21346 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18267), .B1(
        n18293), .B2(n18570), .ZN(n18257) );
  OAI211_X1 U21347 ( .C1(n18283), .C2(n18582), .A(n18258), .B(n18257), .ZN(
        P3_U2819) );
  INV_X1 U21348 ( .A(n18259), .ZN(n18276) );
  AND2_X1 U21349 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18276), .ZN(
        n18279) );
  AOI21_X1 U21350 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18374), .A(
        n18279), .ZN(n18271) );
  AOI22_X1 U21351 ( .A1(n18695), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18260), 
        .B2(n18343), .ZN(n18270) );
  NOR4_X1 U21352 ( .A1(n10304), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n18583), .A4(n18261), .ZN(n18264) );
  OAI221_X1 U21353 ( .B1(n18601), .B2(n18273), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18274), .A(n18583), .ZN(
        n18262) );
  INV_X1 U21354 ( .A(n18262), .ZN(n18263) );
  AOI211_X1 U21355 ( .C1(n18266), .C2(n18265), .A(n18264), .B(n18263), .ZN(
        n18584) );
  OAI21_X1 U21356 ( .B1(n18283), .B2(n18601), .A(n18583), .ZN(n18268) );
  AOI22_X1 U21357 ( .A1(n18293), .A2(n18584), .B1(n18268), .B2(n18267), .ZN(
        n18269) );
  OAI211_X1 U21358 ( .C1(n18272), .C2(n18271), .A(n18270), .B(n18269), .ZN(
        P3_U2820) );
  NAND2_X1 U21359 ( .A1(n18274), .A2(n18273), .ZN(n18275) );
  XNOR2_X1 U21360 ( .A(n18275), .B(n18601), .ZN(n18598) );
  NOR2_X1 U21361 ( .A1(n18701), .A2(n19255), .ZN(n18597) );
  AOI21_X1 U21362 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18374), .A(
        n18276), .ZN(n18278) );
  OAI22_X1 U21363 ( .A1(n18279), .A2(n18278), .B1(n18378), .B2(n18277), .ZN(
        n18280) );
  AOI211_X1 U21364 ( .C1(n18293), .C2(n18598), .A(n18597), .B(n18280), .ZN(
        n18281) );
  OAI221_X1 U21365 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18283), .C1(
        n18601), .C2(n18282), .A(n18281), .ZN(P3_U2821) );
  OAI21_X1 U21366 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18285), .A(
        n18284), .ZN(n18621) );
  NOR2_X1 U21367 ( .A1(n18701), .A2(n19254), .ZN(n18611) );
  OAI211_X1 U21368 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18286), .B(n19036), .ZN(n18289)
         );
  AOI21_X1 U21369 ( .B1(n18334), .B2(n18287), .A(n18368), .ZN(n18297) );
  OAI22_X1 U21370 ( .A1(n17327), .A2(n18289), .B1(n18288), .B2(n18297), .ZN(
        n18290) );
  AOI211_X1 U21371 ( .C1(n18291), .C2(n18343), .A(n18611), .B(n18290), .ZN(
        n18296) );
  OAI21_X1 U21372 ( .B1(n10304), .B2(n18618), .A(n18292), .ZN(n18615) );
  AOI22_X1 U21373 ( .A1(n18294), .A2(n18618), .B1(n18293), .B2(n18615), .ZN(
        n18295) );
  OAI211_X1 U21374 ( .C1(n18385), .C2(n18621), .A(n18296), .B(n18295), .ZN(
        P3_U2822) );
  INV_X1 U21375 ( .A(n18297), .ZN(n18300) );
  NOR2_X1 U21376 ( .A1(n18701), .A2(n19251), .ZN(n18625) );
  AOI221_X1 U21377 ( .B1(n18300), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n18299), .C2(n18298), .A(n18625), .ZN(n18309) );
  AOI21_X1 U21378 ( .B1(n18302), .B2(n18306), .A(n18301), .ZN(n18626) );
  AOI21_X1 U21379 ( .B1(n18305), .B2(n18304), .A(n18303), .ZN(n18307) );
  XNOR2_X1 U21380 ( .A(n18307), .B(n18306), .ZN(n18627) );
  AOI22_X1 U21381 ( .A1(n18375), .A2(n18626), .B1(n18371), .B2(n18627), .ZN(
        n18308) );
  OAI211_X1 U21382 ( .C1(n18378), .C2(n18310), .A(n18309), .B(n18308), .ZN(
        P3_U2823) );
  OAI21_X1 U21383 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18312), .A(
        n18311), .ZN(n18639) );
  NAND2_X1 U21384 ( .A1(n18313), .A2(n19036), .ZN(n18319) );
  OAI21_X1 U21385 ( .B1(n18314), .B2(n19061), .A(n18374), .ZN(n18332) );
  AOI21_X1 U21386 ( .B1(n9759), .B2(n18316), .A(n18315), .ZN(n18637) );
  AOI22_X1 U21387 ( .A1(n18375), .A2(n18637), .B1(n18695), .B2(
        P3_REIP_REG_6__SCAN_IN), .ZN(n18317) );
  OAI221_X1 U21388 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18319), .C1(
        n18318), .C2(n18332), .A(n18317), .ZN(n18320) );
  AOI21_X1 U21389 ( .B1(n18321), .B2(n18343), .A(n18320), .ZN(n18322) );
  OAI21_X1 U21390 ( .B1(n18385), .B2(n18639), .A(n18322), .ZN(P3_U2824) );
  AOI21_X1 U21391 ( .B1(n18323), .B2(n18381), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18333) );
  AOI21_X1 U21392 ( .B1(n18647), .B2(n18324), .A(n18325), .ZN(n18644) );
  INV_X1 U21393 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n21236) );
  NOR2_X1 U21394 ( .A1(n18701), .A2(n21236), .ZN(n18643) );
  OAI21_X1 U21395 ( .B1(n18328), .B2(n18327), .A(n18326), .ZN(n18641) );
  OAI22_X1 U21396 ( .A1(n18378), .A2(n18329), .B1(n18385), .B2(n18641), .ZN(
        n18330) );
  AOI211_X1 U21397 ( .C1(n18375), .C2(n18644), .A(n18643), .B(n18330), .ZN(
        n18331) );
  OAI21_X1 U21398 ( .B1(n18333), .B2(n18332), .A(n18331), .ZN(P3_U2825) );
  AOI21_X1 U21399 ( .B1(n18334), .B2(n18339), .A(n18368), .ZN(n18357) );
  AOI21_X1 U21400 ( .B1(n18337), .B2(n18336), .A(n18335), .ZN(n18338) );
  XNOR2_X1 U21401 ( .A(n18338), .B(n18658), .ZN(n18655) );
  NOR2_X1 U21402 ( .A1(n18701), .A2(n19246), .ZN(n18652) );
  NOR3_X1 U21403 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18339), .A3(
        n19061), .ZN(n18340) );
  AOI211_X1 U21404 ( .C1(n18371), .C2(n18655), .A(n18652), .B(n18340), .ZN(
        n18346) );
  AOI21_X1 U21405 ( .B1(n18342), .B2(n18341), .A(n9776), .ZN(n18653) );
  AOI22_X1 U21406 ( .A1(n18375), .A2(n18653), .B1(n18344), .B2(n18343), .ZN(
        n18345) );
  OAI211_X1 U21407 ( .C1(n18357), .C2(n18347), .A(n18346), .B(n18345), .ZN(
        P3_U2826) );
  OAI21_X1 U21408 ( .B1(n18350), .B2(n18349), .A(n18348), .ZN(n18661) );
  OAI21_X1 U21409 ( .B1(n18353), .B2(n18352), .A(n18351), .ZN(n18354) );
  XNOR2_X1 U21410 ( .A(n18354), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n18664) );
  AOI21_X1 U21411 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18381), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18356) );
  OAI22_X1 U21412 ( .A1(n18357), .A2(n18356), .B1(n18378), .B2(n18355), .ZN(
        n18358) );
  AOI21_X1 U21413 ( .B1(n18375), .B2(n18664), .A(n18358), .ZN(n18359) );
  NAND2_X1 U21414 ( .A1(n18695), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18660) );
  OAI211_X1 U21415 ( .C1(n18385), .C2(n18661), .A(n18359), .B(n18660), .ZN(
        P3_U2827) );
  OAI21_X1 U21416 ( .B1(n18362), .B2(n18361), .A(n18360), .ZN(n18676) );
  XNOR2_X1 U21417 ( .A(n18364), .B(n18363), .ZN(n18675) );
  OAI22_X1 U21418 ( .A1(n18378), .A2(n18365), .B1(n18384), .B2(n18675), .ZN(
        n18366) );
  AOI221_X1 U21419 ( .B1(n18368), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n19036), .C2(n18367), .A(n18366), .ZN(n18369) );
  NAND2_X1 U21420 ( .A1(n18695), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18680) );
  OAI211_X1 U21421 ( .C1(n18385), .C2(n18676), .A(n18369), .B(n18680), .ZN(
        P3_U2828) );
  NOR2_X1 U21422 ( .A1(n18379), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18370) );
  XNOR2_X1 U21423 ( .A(n18370), .B(n18373), .ZN(n18690) );
  AOI22_X1 U21424 ( .A1(n18371), .A2(n18690), .B1(n18695), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18377) );
  AOI22_X1 U21425 ( .A1(n18375), .A2(n18683), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18374), .ZN(n18376) );
  OAI211_X1 U21426 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n18378), .A(
        n18377), .B(n18376), .ZN(P3_U2829) );
  OAI21_X1 U21427 ( .B1(n18379), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18372), .ZN(n18697) );
  INV_X1 U21428 ( .A(n18697), .ZN(n18699) );
  NAND3_X1 U21429 ( .A1(n19214), .A2(n18381), .A3(n18380), .ZN(n18382) );
  AOI22_X1 U21430 ( .A1(n18695), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18382), .ZN(n18383) );
  OAI221_X1 U21431 ( .B1(n18699), .B2(n18385), .C1(n18697), .C2(n18384), .A(
        n18383), .ZN(P3_U2830) );
  NOR2_X1 U21432 ( .A1(n18386), .A2(n18453), .ZN(n18457) );
  NAND2_X1 U21433 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18457), .ZN(
        n18441) );
  NOR2_X1 U21434 ( .A1(n18387), .A2(n18441), .ZN(n18395) );
  OAI22_X1 U21435 ( .A1(n18389), .A2(n18549), .B1(n18388), .B2(n18450), .ZN(
        n18393) );
  NOR2_X1 U21436 ( .A1(n19182), .A2(n18703), .ZN(n18605) );
  INV_X1 U21437 ( .A(n18605), .ZN(n18606) );
  NOR2_X1 U21438 ( .A1(n19169), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18425) );
  AOI221_X1 U21439 ( .B1(n18424), .B2(n18606), .C1(n18408), .C2(n18606), .A(
        n18425), .ZN(n18414) );
  OAI211_X1 U21440 ( .C1(n18391), .C2(n18605), .A(n18390), .B(n18414), .ZN(
        n18392) );
  INV_X1 U21441 ( .A(n18401), .ZN(n18394) );
  MUX2_X1 U21442 ( .A(n18395), .B(n18394), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n18396) );
  AOI22_X1 U21443 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18650), .B1(
        n12963), .B2(n18396), .ZN(n18398) );
  NAND2_X1 U21444 ( .A1(n18695), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18397) );
  OAI211_X1 U21445 ( .C1(n18399), .C2(n18567), .A(n18398), .B(n18397), .ZN(
        P3_U2835) );
  OAI22_X1 U21446 ( .A1(n18401), .A2(n18407), .B1(n18441), .B2(n18400), .ZN(
        n18404) );
  OAI221_X1 U21447 ( .B1(n18404), .B2(n18403), .C1(n18404), .C2(n18402), .A(
        n12963), .ZN(n18406) );
  OAI211_X1 U21448 ( .C1(n18685), .C2(n18407), .A(n18406), .B(n18405), .ZN(
        P3_U2836) );
  INV_X1 U21449 ( .A(n18617), .ZN(n18541) );
  AOI211_X1 U21450 ( .C1(n10298), .C2(n18408), .A(n18413), .B(n18432), .ZN(
        n18415) );
  NAND3_X1 U21451 ( .A1(n18411), .A2(n18410), .A3(n18409), .ZN(n18412) );
  AOI22_X1 U21452 ( .A1(n18415), .A2(n18414), .B1(n18413), .B2(n18412), .ZN(
        n18416) );
  AOI22_X1 U21453 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18650), .B1(
        n12963), .B2(n18416), .ZN(n18418) );
  OAI211_X1 U21454 ( .C1(n18419), .C2(n18567), .A(n18418), .B(n18417), .ZN(
        n18420) );
  AOI21_X1 U21455 ( .B1(n18698), .B2(n18421), .A(n18420), .ZN(n18422) );
  OAI21_X1 U21456 ( .B1(n18541), .B2(n18423), .A(n18422), .ZN(P3_U2837) );
  INV_X1 U21457 ( .A(n18479), .ZN(n18440) );
  NOR2_X1 U21458 ( .A1(n18701), .A2(n19284), .ZN(n18436) );
  INV_X1 U21459 ( .A(n18424), .ZN(n18426) );
  INV_X1 U21460 ( .A(n18425), .ZN(n18604) );
  OAI21_X1 U21461 ( .B1(n18426), .B2(n18605), .A(n18604), .ZN(n18430) );
  OAI22_X1 U21462 ( .A1(n18428), .A2(n18549), .B1(n18427), .B2(n18450), .ZN(
        n18429) );
  NOR3_X1 U21463 ( .A1(n18650), .A2(n18430), .A3(n18429), .ZN(n18434) );
  NAND2_X1 U21464 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18434), .ZN(
        n18431) );
  OAI21_X1 U21465 ( .B1(n18432), .B2(n18431), .A(n18701), .ZN(n18446) );
  AOI211_X1 U21466 ( .C1(n18608), .C2(n18434), .A(n18433), .B(n18446), .ZN(
        n18435) );
  AOI211_X1 U21467 ( .C1(n18616), .C2(n18437), .A(n18436), .B(n18435), .ZN(
        n18438) );
  OAI21_X1 U21468 ( .B1(n18440), .B2(n18439), .A(n18438), .ZN(P3_U2838) );
  INV_X1 U21469 ( .A(n18441), .ZN(n18442) );
  AOI21_X1 U21470 ( .B1(n18442), .B2(n18685), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18447) );
  AOI21_X1 U21471 ( .B1(n18444), .B2(n18616), .A(n18443), .ZN(n18445) );
  OAI21_X1 U21472 ( .B1(n18447), .B2(n18446), .A(n18445), .ZN(P3_U2839) );
  AOI22_X1 U21473 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18650), .B1(
        n18695), .B2(P3_REIP_REG_22__SCAN_IN), .ZN(n18459) );
  AOI22_X1 U21474 ( .A1(n10298), .A2(n18464), .B1(n18465), .B2(n18547), .ZN(
        n18455) );
  NAND2_X1 U21475 ( .A1(n18450), .A2(n18549), .ZN(n18576) );
  AOI22_X1 U21476 ( .A1(n18703), .A2(n18451), .B1(n18453), .B2(n18576), .ZN(
        n18466) );
  INV_X1 U21477 ( .A(n18466), .ZN(n18452) );
  AOI221_X1 U21478 ( .B1(n18453), .B2(n19182), .C1(n18505), .C2(n19182), .A(
        n18452), .ZN(n18454) );
  NAND4_X1 U21479 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18463), .A3(
        n18455), .A4(n18454), .ZN(n18456) );
  OAI211_X1 U21480 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n18457), .A(
        n12963), .B(n18456), .ZN(n18458) );
  OAI211_X1 U21481 ( .C1(n18460), .C2(n18567), .A(n18459), .B(n18458), .ZN(
        P3_U2840) );
  NOR2_X1 U21482 ( .A1(n18701), .A2(n19277), .ZN(n18467) );
  OAI21_X1 U21483 ( .B1(n18505), .B2(n18461), .A(n19182), .ZN(n18462) );
  NAND3_X1 U21484 ( .A1(n18463), .A2(n12963), .A3(n18462), .ZN(n18471) );
  AOI22_X1 U21485 ( .A1(n18695), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18479), 
        .B2(n18470), .ZN(n18476) );
  AOI21_X1 U21486 ( .B1(n18576), .B2(n18472), .A(n18471), .ZN(n18473) );
  NOR2_X1 U21487 ( .A1(n18695), .A2(n18473), .ZN(n18480) );
  INV_X1 U21488 ( .A(n18684), .ZN(n18531) );
  NOR3_X1 U21489 ( .A1(n18531), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n18707), .ZN(n18474) );
  OAI21_X1 U21490 ( .B1(n18480), .B2(n18474), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18475) );
  OAI211_X1 U21491 ( .C1(n18567), .C2(n18477), .A(n18476), .B(n18475), .ZN(
        P3_U2842) );
  AOI22_X1 U21492 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18480), .B1(
        n18479), .B2(n18478), .ZN(n18482) );
  OAI211_X1 U21493 ( .C1(n18483), .C2(n18567), .A(n18482), .B(n18481), .ZN(
        P3_U2843) );
  NAND2_X1 U21494 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18485) );
  INV_X1 U21495 ( .A(n18671), .ZN(n18484) );
  OAI22_X1 U21496 ( .A1(n18603), .A2(n19177), .B1(n18485), .B2(n18484), .ZN(
        n18666) );
  NAND2_X1 U21497 ( .A1(n12963), .A2(n18666), .ZN(n18640) );
  NOR2_X1 U21498 ( .A1(n18515), .A2(n18640), .ZN(n18542) );
  AOI22_X1 U21499 ( .A1(n10179), .A2(n18542), .B1(n12963), .B2(n18486), .ZN(
        n18513) );
  NAND3_X1 U21500 ( .A1(n18487), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18604), .ZN(n18488) );
  AOI22_X1 U21501 ( .A1(n18489), .A2(n18576), .B1(n18606), .B2(n18488), .ZN(
        n18491) );
  AND4_X1 U21502 ( .A1(n12963), .A2(n18504), .A3(n18491), .A4(n18490), .ZN(
        n18497) );
  AOI221_X1 U21503 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18497), 
        .C1(n18605), .C2(n18497), .A(n18695), .ZN(n18493) );
  AOI22_X1 U21504 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18493), .B1(
        n18616), .B2(n18492), .ZN(n18495) );
  NAND2_X1 U21505 ( .A1(n18695), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18494) );
  OAI211_X1 U21506 ( .C1(n18513), .C2(n18496), .A(n18495), .B(n18494), .ZN(
        P3_U2844) );
  NOR2_X1 U21507 ( .A1(n18695), .A2(n18497), .ZN(n18500) );
  INV_X1 U21508 ( .A(n18513), .ZN(n18498) );
  AOI22_X1 U21509 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18500), .B1(
        n18499), .B2(n18498), .ZN(n18502) );
  NAND2_X1 U21510 ( .A1(n18695), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18501) );
  OAI211_X1 U21511 ( .C1(n18503), .C2(n18567), .A(n18502), .B(n18501), .ZN(
        P3_U2845) );
  NAND2_X1 U21512 ( .A1(n12963), .A2(n18504), .ZN(n18508) );
  INV_X1 U21513 ( .A(n18608), .ZN(n18610) );
  INV_X1 U21514 ( .A(n18547), .ZN(n18586) );
  AOI22_X1 U21515 ( .A1(n10298), .A2(n18548), .B1(n18703), .B2(n18546), .ZN(
        n18530) );
  OAI21_X1 U21516 ( .B1(n9996), .B2(n19182), .A(n18505), .ZN(n18506) );
  OAI211_X1 U21517 ( .C1(n18507), .C2(n18586), .A(n18530), .B(n18506), .ZN(
        n18516) );
  OAI221_X1 U21518 ( .B1(n18508), .B2(n18610), .C1(n18508), .C2(n18516), .A(
        n18701), .ZN(n18511) );
  AOI22_X1 U21519 ( .A1(n18695), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18616), 
        .B2(n18509), .ZN(n18510) );
  OAI221_X1 U21520 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18513), 
        .C1(n18512), .C2(n18511), .A(n18510), .ZN(P3_U2846) );
  AOI22_X1 U21521 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18650), .B1(
        n18695), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n18526) );
  NAND2_X1 U21522 ( .A1(n18571), .A2(n18514), .ZN(n18518) );
  INV_X1 U21523 ( .A(n18666), .ZN(n18623) );
  NOR3_X1 U21524 ( .A1(n18623), .A2(n18515), .A3(n18528), .ZN(n18533) );
  OAI221_X1 U21525 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18533), .A(n18516), .ZN(
        n18517) );
  OAI21_X1 U21526 ( .B1(n18519), .B2(n18518), .A(n18517), .ZN(n18521) );
  AOI22_X1 U21527 ( .A1(n12963), .A2(n18521), .B1(n18616), .B2(n18520), .ZN(
        n18525) );
  NAND3_X1 U21528 ( .A1(n18698), .A2(n18523), .A3(n18522), .ZN(n18524) );
  NAND3_X1 U21529 ( .A1(n18526), .A2(n18525), .A3(n18524), .ZN(P3_U2847) );
  AOI21_X1 U21530 ( .B1(n18558), .B2(n18593), .A(n19169), .ZN(n18554) );
  OAI21_X1 U21531 ( .B1(n18558), .B2(n19177), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18527) );
  AOI211_X1 U21532 ( .C1(n18703), .C2(n18528), .A(n18554), .B(n18527), .ZN(
        n18529) );
  OAI211_X1 U21533 ( .C1(n18531), .C2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n18530), .B(n18529), .ZN(n18532) );
  OAI211_X1 U21534 ( .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18533), .A(
        n12963), .B(n18532), .ZN(n18534) );
  OAI21_X1 U21535 ( .B1(n19263), .B2(n18701), .A(n18534), .ZN(n18538) );
  OAI22_X1 U21536 ( .A1(n18536), .A2(n18567), .B1(n18677), .B2(n18535), .ZN(
        n18537) );
  AOI211_X1 U21537 ( .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18650), .A(
        n18538), .B(n18537), .ZN(n18539) );
  OAI21_X1 U21538 ( .B1(n18541), .B2(n18540), .A(n18539), .ZN(P3_U2848) );
  NOR2_X1 U21539 ( .A1(n12890), .A2(n18541), .ZN(n18543) );
  AOI211_X1 U21540 ( .C1(n18698), .C2(n18544), .A(n18543), .B(n18542), .ZN(
        n18602) );
  AOI22_X1 U21541 ( .A1(n18695), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18616), 
        .B2(n18545), .ZN(n18556) );
  AND2_X1 U21542 ( .A1(n18703), .A2(n18546), .ZN(n18588) );
  OAI21_X1 U21543 ( .B1(n18588), .B2(n18562), .A(n18547), .ZN(n18578) );
  NAND2_X1 U21544 ( .A1(n10298), .A2(n18548), .ZN(n18573) );
  OAI211_X1 U21545 ( .C1(n18550), .C2(n18549), .A(n18578), .B(n18573), .ZN(
        n18551) );
  AOI21_X1 U21546 ( .B1(n19150), .B2(n18552), .A(n18551), .ZN(n18559) );
  OAI211_X1 U21547 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18586), .A(
        n12963), .B(n18559), .ZN(n18553) );
  OAI211_X1 U21548 ( .C1(n18554), .C2(n18553), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18701), .ZN(n18555) );
  OAI211_X1 U21549 ( .C1(n18602), .C2(n18557), .A(n18556), .B(n18555), .ZN(
        P3_U2849) );
  AND2_X1 U21550 ( .A1(n18558), .A2(n18593), .ZN(n18560) );
  OAI211_X1 U21551 ( .C1(n18560), .C2(n19169), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n18559), .ZN(n18564) );
  OAI22_X1 U21552 ( .A1(n18602), .A2(n18562), .B1(n18561), .B2(n18702), .ZN(
        n18563) );
  AOI22_X1 U21553 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18650), .B1(
        n18564), .B2(n18563), .ZN(n18566) );
  NAND2_X1 U21554 ( .A1(n18695), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18565) );
  OAI211_X1 U21555 ( .C1(n18568), .C2(n18567), .A(n18566), .B(n18565), .ZN(
        P3_U2850) );
  AOI21_X1 U21556 ( .B1(n18616), .B2(n18570), .A(n18569), .ZN(n18581) );
  AOI21_X1 U21557 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18593), .A(
        n19169), .ZN(n18575) );
  AOI22_X1 U21558 ( .A1(n19150), .A2(n18572), .B1(n18571), .B2(n12890), .ZN(
        n18574) );
  NAND3_X1 U21559 ( .A1(n12963), .A2(n18574), .A3(n18573), .ZN(n18596) );
  AOI211_X1 U21560 ( .C1(n18577), .C2(n18576), .A(n18575), .B(n18596), .ZN(
        n18585) );
  OAI211_X1 U21561 ( .C1(n19169), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18585), .B(n18578), .ZN(n18579) );
  NAND3_X1 U21562 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18701), .A3(
        n18579), .ZN(n18580) );
  OAI211_X1 U21563 ( .C1(n18602), .C2(n18582), .A(n18581), .B(n18580), .ZN(
        P3_U2851) );
  NAND2_X1 U21564 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18583), .ZN(
        n18591) );
  AOI22_X1 U21565 ( .A1(n18695), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18616), 
        .B2(n18584), .ZN(n18590) );
  OAI21_X1 U21566 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18586), .A(
        n18585), .ZN(n18587) );
  OAI211_X1 U21567 ( .C1(n18588), .C2(n18587), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18701), .ZN(n18589) );
  OAI211_X1 U21568 ( .C1(n18602), .C2(n18591), .A(n18590), .B(n18589), .ZN(
        P3_U2852) );
  AOI21_X1 U21569 ( .B1(n18703), .B2(n18613), .A(n19182), .ZN(n18592) );
  OAI22_X1 U21570 ( .A1(n19184), .A2(n18594), .B1(n18593), .B2(n18592), .ZN(
        n18595) );
  OAI21_X1 U21571 ( .B1(n18596), .B2(n18595), .A(n18701), .ZN(n18600) );
  AOI21_X1 U21572 ( .B1(n18616), .B2(n18598), .A(n18597), .ZN(n18599) );
  OAI221_X1 U21573 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18602), .C1(
        n18601), .C2(n18600), .A(n18599), .ZN(P3_U2853) );
  NAND3_X1 U21574 ( .A1(n18607), .A2(n12963), .A3(n18666), .ZN(n18635) );
  NOR2_X1 U21575 ( .A1(n18609), .A2(n18635), .ZN(n18614) );
  NAND2_X1 U21576 ( .A1(n10298), .A2(n18603), .ZN(n18673) );
  OAI211_X1 U21577 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n18605), .A(
        n18673), .B(n18604), .ZN(n18669) );
  AOI21_X1 U21578 ( .B1(n18682), .B2(n18606), .A(n18669), .ZN(n18649) );
  OAI21_X1 U21579 ( .B1(n18608), .B2(n18607), .A(n18649), .ZN(n18632) );
  AOI21_X1 U21580 ( .B1(n18610), .B2(n18609), .A(n18632), .ZN(n18631) );
  OAI21_X1 U21581 ( .B1(n18631), .B2(n18686), .A(n18685), .ZN(n18612) );
  AOI221_X1 U21582 ( .B1(n18614), .B2(n18613), .C1(n18612), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18611), .ZN(n18620) );
  AOI22_X1 U21583 ( .A1(n18618), .A2(n18617), .B1(n18616), .B2(n18615), .ZN(
        n18619) );
  OAI211_X1 U21584 ( .C1(n18677), .C2(n18621), .A(n18620), .B(n18619), .ZN(
        P3_U2854) );
  NOR2_X1 U21585 ( .A1(n18623), .A2(n18622), .ZN(n18624) );
  OAI221_X1 U21586 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18624), .A(n12963), .ZN(
        n18630) );
  AOI21_X1 U21587 ( .B1(n18650), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18625), .ZN(n18629) );
  AOI22_X1 U21588 ( .A1(n18698), .A2(n18627), .B1(n18700), .B2(n18626), .ZN(
        n18628) );
  OAI211_X1 U21589 ( .C1(n18631), .C2(n18630), .A(n18629), .B(n18628), .ZN(
        P3_U2855) );
  INV_X1 U21590 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18634) );
  AOI21_X1 U21591 ( .B1(n12963), .B2(n18632), .A(n18650), .ZN(n18646) );
  NAND2_X1 U21592 ( .A1(n18695), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n18633) );
  OAI221_X1 U21593 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18635), .C1(
        n18634), .C2(n18646), .A(n18633), .ZN(n18636) );
  AOI21_X1 U21594 ( .B1(n18700), .B2(n18637), .A(n18636), .ZN(n18638) );
  OAI21_X1 U21595 ( .B1(n18677), .B2(n18639), .A(n18638), .ZN(P3_U2856) );
  NOR2_X1 U21596 ( .A1(n12853), .A2(n18640), .ZN(n18654) );
  NAND2_X1 U21597 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18654), .ZN(
        n18648) );
  NOR2_X1 U21598 ( .A1(n18677), .A2(n18641), .ZN(n18642) );
  AOI211_X1 U21599 ( .C1(n18700), .C2(n18644), .A(n18643), .B(n18642), .ZN(
        n18645) );
  OAI221_X1 U21600 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18648), .C1(
        n18647), .C2(n18646), .A(n18645), .ZN(P3_U2857) );
  NAND2_X1 U21601 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18649), .ZN(
        n18665) );
  AOI21_X1 U21602 ( .B1(n18651), .B2(n18665), .A(n18650), .ZN(n18659) );
  AOI21_X1 U21603 ( .B1(n18653), .B2(n18700), .A(n18652), .ZN(n18657) );
  AOI22_X1 U21604 ( .A1(n18655), .A2(n18698), .B1(n18654), .B2(n18658), .ZN(
        n18656) );
  OAI211_X1 U21605 ( .C1(n18659), .C2(n18658), .A(n18657), .B(n18656), .ZN(
        P3_U2858) );
  INV_X1 U21606 ( .A(n18660), .ZN(n18663) );
  OAI22_X1 U21607 ( .A1(n12853), .A2(n18685), .B1(n18677), .B2(n18661), .ZN(
        n18662) );
  AOI211_X1 U21608 ( .C1(n18664), .C2(n18700), .A(n18663), .B(n18662), .ZN(
        n18668) );
  OAI211_X1 U21609 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18666), .A(
        n12963), .B(n18665), .ZN(n18667) );
  NAND2_X1 U21610 ( .A1(n18668), .A2(n18667), .ZN(P3_U2859) );
  NOR2_X1 U21611 ( .A1(n19320), .A2(n18687), .ZN(n18670) );
  AOI21_X1 U21612 ( .B1(n10298), .B2(n18670), .A(n18669), .ZN(n18674) );
  NAND3_X1 U21613 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18671), .A3(
        n18682), .ZN(n18672) );
  OAI211_X1 U21614 ( .C1(n18674), .C2(n18682), .A(n18673), .B(n18672), .ZN(
        n18679) );
  OAI22_X1 U21615 ( .A1(n18677), .A2(n18676), .B1(n18693), .B2(n18675), .ZN(
        n18678) );
  AOI21_X1 U21616 ( .B1(n12963), .B2(n18679), .A(n18678), .ZN(n18681) );
  OAI211_X1 U21617 ( .C1(n18685), .C2(n18682), .A(n18681), .B(n18680), .ZN(
        P3_U2860) );
  INV_X1 U21618 ( .A(n18683), .ZN(n18694) );
  NAND3_X1 U21619 ( .A1(n12963), .A2(n18684), .A3(n18687), .ZN(n18705) );
  AOI21_X1 U21620 ( .B1(n18685), .B2(n18705), .A(n19320), .ZN(n18689) );
  AOI211_X1 U21621 ( .C1(n19184), .C2(n18687), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18686), .ZN(n18688) );
  AOI211_X1 U21622 ( .C1(n18698), .C2(n18690), .A(n18689), .B(n18688), .ZN(
        n18692) );
  NAND2_X1 U21623 ( .A1(n18695), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18691) );
  OAI211_X1 U21624 ( .C1(n18694), .C2(n18693), .A(n18692), .B(n18691), .ZN(
        P3_U2861) );
  AND2_X1 U21625 ( .A1(n18695), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18696) );
  AOI221_X1 U21626 ( .B1(n18700), .B2(n18699), .C1(n18698), .C2(n18697), .A(
        n18696), .ZN(n18706) );
  OAI211_X1 U21627 ( .C1(n18703), .C2(n18702), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18701), .ZN(n18704) );
  NAND3_X1 U21628 ( .A1(n18706), .A2(n18705), .A3(n18704), .ZN(P3_U2862) );
  AOI211_X1 U21629 ( .C1(n21320), .C2(n18708), .A(n18707), .B(n19214), .ZN(
        n19209) );
  INV_X1 U21630 ( .A(n18760), .ZN(n18709) );
  OAI21_X1 U21631 ( .B1(n19209), .B2(n18709), .A(n18718), .ZN(n18710) );
  OAI221_X1 U21632 ( .B1(n19188), .B2(n19352), .C1(n19188), .C2(n18718), .A(
        n18710), .ZN(P3_U2863) );
  NAND2_X1 U21633 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18870) );
  AOI221_X1 U21634 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18870), .C1(n18712), 
        .C2(n18870), .A(n18711), .ZN(n18717) );
  INV_X1 U21635 ( .A(n18713), .ZN(n18714) );
  AOI22_X1 U21636 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18714), .B1(
        n18781), .B2(n18718), .ZN(n18716) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18717), .B1(
        n18716), .B2(n19193), .ZN(P3_U2865) );
  NAND2_X1 U21638 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19196), .ZN(
        n18848) );
  INV_X1 U21639 ( .A(n18848), .ZN(n18894) );
  NOR2_X1 U21640 ( .A1(n18985), .A2(n18894), .ZN(n18715) );
  OAI22_X1 U21641 ( .A1(n18717), .A2(n19196), .B1(n18716), .B2(n18715), .ZN(
        P3_U2866) );
  NOR2_X1 U21642 ( .A1(n19197), .A2(n18718), .ZN(P3_U2867) );
  NOR2_X1 U21643 ( .A1(n18720), .A2(n18719), .ZN(n18750) );
  INV_X1 U21644 ( .A(n18750), .ZN(n18756) );
  NOR2_X1 U21645 ( .A1(n18721), .A2(n18756), .ZN(n19096) );
  NAND2_X1 U21646 ( .A1(n19189), .A2(n19188), .ZN(n19190) );
  INV_X1 U21647 ( .A(n19190), .ZN(n19006) );
  NOR2_X1 U21648 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18804) );
  NAND2_X1 U21649 ( .A1(n19006), .A2(n18804), .ZN(n18824) );
  NAND2_X1 U21650 ( .A1(n19036), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19099) );
  INV_X1 U21651 ( .A(n19099), .ZN(n19033) );
  INV_X1 U21652 ( .A(n18870), .ZN(n18722) );
  NAND2_X1 U21653 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18722), .ZN(
        n19090) );
  NOR2_X2 U21654 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19090), .ZN(
        n19085) );
  NOR2_X2 U21655 ( .A1(n19063), .A2(n18723), .ZN(n19093) );
  NOR2_X2 U21656 ( .A1(n19188), .A2(n19090), .ZN(n19143) );
  NOR2_X1 U21657 ( .A1(n19143), .A2(n18817), .ZN(n18782) );
  NOR2_X1 U21658 ( .A1(n19091), .A2(n18782), .ZN(n18755) );
  AOI22_X1 U21659 ( .A1(n19033), .A2(n19085), .B1(n19093), .B2(n18755), .ZN(
        n18729) );
  NAND2_X1 U21660 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19189), .ZN(
        n18849) );
  INV_X1 U21661 ( .A(n18849), .ZN(n18937) );
  NOR2_X1 U21662 ( .A1(n19193), .A2(n19196), .ZN(n19095) );
  NAND2_X1 U21663 ( .A1(n18937), .A2(n19095), .ZN(n19105) );
  NAND2_X1 U21664 ( .A1(n19105), .A2(n19083), .ZN(n19060) );
  NOR2_X1 U21665 ( .A1(n18782), .A2(n19063), .ZN(n18726) );
  INV_X1 U21666 ( .A(n18724), .ZN(n18725) );
  AOI22_X1 U21667 ( .A1(n19036), .A2(n19060), .B1(n18726), .B2(n18725), .ZN(
        n18757) );
  NOR2_X2 U21668 ( .A1(n18727), .A2(n19061), .ZN(n19092) );
  INV_X1 U21669 ( .A(n19105), .ZN(n19141) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18757), .B1(
        n19092), .B2(n19141), .ZN(n18728) );
  OAI211_X1 U21671 ( .C1(n19039), .C2(n18824), .A(n18729), .B(n18728), .ZN(
        P3_U2868) );
  NAND2_X1 U21672 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19036), .ZN(n19043) );
  NAND2_X1 U21673 ( .A1(n19036), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19106) );
  INV_X1 U21674 ( .A(n19106), .ZN(n19040) );
  AND2_X1 U21675 ( .A1(n19010), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19100) );
  AOI22_X1 U21676 ( .A1(n19040), .A2(n19085), .B1(n19100), .B2(n18755), .ZN(
        n18731) );
  NOR2_X2 U21677 ( .A1(n19360), .A2(n18756), .ZN(n19102) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18757), .B1(
        n19102), .B2(n18817), .ZN(n18730) );
  OAI211_X1 U21679 ( .C1(n19043), .C2(n19105), .A(n18731), .B(n18730), .ZN(
        P3_U2869) );
  NAND2_X1 U21680 ( .A1(n18750), .A2(n18732), .ZN(n19112) );
  AND2_X1 U21681 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19036), .ZN(n19109) );
  NOR2_X2 U21682 ( .A1(n19063), .A2(n18733), .ZN(n19107) );
  AOI22_X1 U21683 ( .A1(n19109), .A2(n19141), .B1(n19107), .B2(n18755), .ZN(
        n18735) );
  AND2_X1 U21684 ( .A1(n19036), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19108) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18757), .B1(
        n19108), .B2(n19085), .ZN(n18734) );
  OAI211_X1 U21686 ( .C1(n19112), .C2(n18824), .A(n18735), .B(n18734), .ZN(
        P3_U2870) );
  NAND2_X1 U21687 ( .A1(n18750), .A2(n18736), .ZN(n19118) );
  AND2_X1 U21688 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19036), .ZN(n19115) );
  NOR2_X2 U21689 ( .A1(n19063), .A2(n18737), .ZN(n19113) );
  AOI22_X1 U21690 ( .A1(n19115), .A2(n19141), .B1(n19113), .B2(n18755), .ZN(
        n18740) );
  NOR2_X2 U21691 ( .A1(n19061), .A2(n18738), .ZN(n19114) );
  AOI22_X1 U21692 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18757), .B1(
        n19114), .B2(n19085), .ZN(n18739) );
  OAI211_X1 U21693 ( .C1(n19118), .C2(n18824), .A(n18740), .B(n18739), .ZN(
        P3_U2871) );
  NOR2_X1 U21694 ( .A1(n21246), .A2(n19061), .ZN(n19074) );
  NAND2_X1 U21695 ( .A1(n19036), .A2(BUF2_REG_20__SCAN_IN), .ZN(n19077) );
  INV_X1 U21696 ( .A(n19077), .ZN(n19120) );
  NOR2_X2 U21697 ( .A1(n19063), .A2(n18741), .ZN(n19119) );
  AOI22_X1 U21698 ( .A1(n19120), .A2(n19085), .B1(n19119), .B2(n18755), .ZN(
        n18744) );
  NOR2_X2 U21699 ( .A1(n18742), .A2(n18756), .ZN(n19121) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18757), .B1(
        n19121), .B2(n18817), .ZN(n18743) );
  OAI211_X1 U21701 ( .C1(n19124), .C2(n19105), .A(n18744), .B(n18743), .ZN(
        P3_U2872) );
  NAND2_X1 U21702 ( .A1(n18750), .A2(n18745), .ZN(n19130) );
  NOR2_X2 U21703 ( .A1(n19061), .A2(n19558), .ZN(n19127) );
  NOR2_X2 U21704 ( .A1(n19063), .A2(n18746), .ZN(n19125) );
  AOI22_X1 U21705 ( .A1(n19127), .A2(n19085), .B1(n19125), .B2(n18755), .ZN(
        n18748) );
  AND2_X1 U21706 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19036), .ZN(n19126) );
  AOI22_X1 U21707 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18757), .B1(
        n19126), .B2(n19141), .ZN(n18747) );
  OAI211_X1 U21708 ( .C1(n19130), .C2(n18824), .A(n18748), .B(n18747), .ZN(
        P3_U2873) );
  NAND2_X1 U21709 ( .A1(n18750), .A2(n18749), .ZN(n19138) );
  NOR2_X2 U21710 ( .A1(n19063), .A2(n18751), .ZN(n19131) );
  AOI22_X1 U21711 ( .A1(n19134), .A2(n19141), .B1(n19131), .B2(n18755), .ZN(
        n18753) );
  NOR2_X2 U21712 ( .A1(n19061), .A2(n19564), .ZN(n19132) );
  AOI22_X1 U21713 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18757), .B1(
        n19132), .B2(n19085), .ZN(n18752) );
  OAI211_X1 U21714 ( .C1(n19138), .C2(n18824), .A(n18753), .B(n18752), .ZN(
        P3_U2874) );
  NOR2_X1 U21715 ( .A1(n19061), .A2(n18754), .ZN(n18978) );
  NAND2_X1 U21716 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19036), .ZN(n18983) );
  INV_X1 U21717 ( .A(n18983), .ZN(n19142) );
  NOR2_X2 U21718 ( .A1(n21237), .A2(n19063), .ZN(n19140) );
  AOI22_X1 U21719 ( .A1(n19142), .A2(n19085), .B1(n19140), .B2(n18755), .ZN(
        n18759) );
  NOR2_X2 U21720 ( .A1(n12696), .A2(n18756), .ZN(n19144) );
  AOI22_X1 U21721 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18757), .B1(
        n19144), .B2(n18817), .ZN(n18758) );
  OAI211_X1 U21722 ( .C1(n19149), .C2(n19105), .A(n18759), .B(n18758), .ZN(
        P3_U2875) );
  NAND2_X1 U21723 ( .A1(n18937), .A2(n18804), .ZN(n18846) );
  INV_X1 U21724 ( .A(n18804), .ZN(n18780) );
  OR2_X1 U21725 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19091), .ZN(
        n19031) );
  NOR2_X1 U21726 ( .A1(n18780), .A2(n19031), .ZN(n18776) );
  AOI22_X1 U21727 ( .A1(n19033), .A2(n19143), .B1(n19093), .B2(n18776), .ZN(
        n18763) );
  INV_X1 U21728 ( .A(n19090), .ZN(n18761) );
  NAND2_X1 U21729 ( .A1(n19010), .A2(n18760), .ZN(n18803) );
  NOR2_X1 U21730 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18803), .ZN(
        n19034) );
  AOI22_X1 U21731 ( .A1(n19036), .A2(n18761), .B1(n18804), .B2(n19034), .ZN(
        n18777) );
  AOI22_X1 U21732 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18777), .B1(
        n19092), .B2(n19085), .ZN(n18762) );
  OAI211_X1 U21733 ( .C1(n19039), .C2(n18846), .A(n18763), .B(n18762), .ZN(
        P3_U2876) );
  AOI22_X1 U21734 ( .A1(n19040), .A2(n19143), .B1(n19100), .B2(n18776), .ZN(
        n18765) );
  AOI22_X1 U21735 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18777), .B1(
        n19102), .B2(n18839), .ZN(n18764) );
  OAI211_X1 U21736 ( .C1(n19043), .C2(n19083), .A(n18765), .B(n18764), .ZN(
        P3_U2877) );
  AOI22_X1 U21737 ( .A1(n19108), .A2(n19143), .B1(n19107), .B2(n18776), .ZN(
        n18767) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18777), .B1(
        n19109), .B2(n19085), .ZN(n18766) );
  OAI211_X1 U21739 ( .C1(n19112), .C2(n18846), .A(n18767), .B(n18766), .ZN(
        P3_U2878) );
  AOI22_X1 U21740 ( .A1(n19114), .A2(n19143), .B1(n19113), .B2(n18776), .ZN(
        n18769) );
  AOI22_X1 U21741 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18777), .B1(
        n19115), .B2(n19085), .ZN(n18768) );
  OAI211_X1 U21742 ( .C1(n19118), .C2(n18846), .A(n18769), .B(n18768), .ZN(
        P3_U2879) );
  AOI22_X1 U21743 ( .A1(n19120), .A2(n19143), .B1(n19119), .B2(n18776), .ZN(
        n18771) );
  AOI22_X1 U21744 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18777), .B1(
        n19121), .B2(n18839), .ZN(n18770) );
  OAI211_X1 U21745 ( .C1(n19124), .C2(n19083), .A(n18771), .B(n18770), .ZN(
        P3_U2880) );
  AOI22_X1 U21746 ( .A1(n19127), .A2(n19143), .B1(n19125), .B2(n18776), .ZN(
        n18773) );
  AOI22_X1 U21747 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18777), .B1(
        n19126), .B2(n19085), .ZN(n18772) );
  OAI211_X1 U21748 ( .C1(n19130), .C2(n18846), .A(n18773), .B(n18772), .ZN(
        P3_U2881) );
  AOI22_X1 U21749 ( .A1(n19134), .A2(n19085), .B1(n19131), .B2(n18776), .ZN(
        n18775) );
  AOI22_X1 U21750 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18777), .B1(
        n19132), .B2(n19143), .ZN(n18774) );
  OAI211_X1 U21751 ( .C1(n19138), .C2(n18846), .A(n18775), .B(n18774), .ZN(
        P3_U2882) );
  AOI22_X1 U21752 ( .A1(n19142), .A2(n19143), .B1(n19140), .B2(n18776), .ZN(
        n18779) );
  AOI22_X1 U21753 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18777), .B1(
        n19144), .B2(n18839), .ZN(n18778) );
  OAI211_X1 U21754 ( .C1(n19149), .C2(n19083), .A(n18779), .B(n18778), .ZN(
        P3_U2883) );
  NOR2_X1 U21755 ( .A1(n19189), .A2(n18780), .ZN(n18847) );
  NAND2_X1 U21756 ( .A1(n18847), .A2(n19188), .ZN(n18860) );
  NOR2_X1 U21757 ( .A1(n18839), .A2(n18865), .ZN(n18825) );
  NOR2_X1 U21758 ( .A1(n19091), .A2(n18825), .ZN(n18798) );
  AOI22_X1 U21759 ( .A1(n19033), .A2(n18817), .B1(n19093), .B2(n18798), .ZN(
        n18785) );
  INV_X1 U21760 ( .A(n18781), .ZN(n19007) );
  OAI21_X1 U21761 ( .B1(n18782), .B2(n19007), .A(n18825), .ZN(n18783) );
  OAI211_X1 U21762 ( .C1(n18865), .C2(n19335), .A(n19010), .B(n18783), .ZN(
        n18799) );
  AOI22_X1 U21763 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18799), .B1(
        n19092), .B2(n19143), .ZN(n18784) );
  OAI211_X1 U21764 ( .C1(n19039), .C2(n18860), .A(n18785), .B(n18784), .ZN(
        P3_U2884) );
  INV_X1 U21765 ( .A(n19043), .ZN(n19101) );
  AOI22_X1 U21766 ( .A1(n19101), .A2(n19143), .B1(n19100), .B2(n18798), .ZN(
        n18787) );
  AOI22_X1 U21767 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18799), .B1(
        n19102), .B2(n18865), .ZN(n18786) );
  OAI211_X1 U21768 ( .C1(n19106), .C2(n18824), .A(n18787), .B(n18786), .ZN(
        P3_U2885) );
  AOI22_X1 U21769 ( .A1(n19108), .A2(n18817), .B1(n19107), .B2(n18798), .ZN(
        n18789) );
  AOI22_X1 U21770 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18799), .B1(
        n19109), .B2(n19143), .ZN(n18788) );
  OAI211_X1 U21771 ( .C1(n19112), .C2(n18860), .A(n18789), .B(n18788), .ZN(
        P3_U2886) );
  AOI22_X1 U21772 ( .A1(n19114), .A2(n18817), .B1(n19113), .B2(n18798), .ZN(
        n18791) );
  AOI22_X1 U21773 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18799), .B1(
        n19115), .B2(n19143), .ZN(n18790) );
  OAI211_X1 U21774 ( .C1(n19118), .C2(n18860), .A(n18791), .B(n18790), .ZN(
        P3_U2887) );
  AOI22_X1 U21775 ( .A1(n19074), .A2(n19143), .B1(n19119), .B2(n18798), .ZN(
        n18793) );
  AOI22_X1 U21776 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18799), .B1(
        n19121), .B2(n18865), .ZN(n18792) );
  OAI211_X1 U21777 ( .C1(n19077), .C2(n18824), .A(n18793), .B(n18792), .ZN(
        P3_U2888) );
  AOI22_X1 U21778 ( .A1(n19127), .A2(n18817), .B1(n19125), .B2(n18798), .ZN(
        n18795) );
  AOI22_X1 U21779 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18799), .B1(
        n19126), .B2(n19143), .ZN(n18794) );
  OAI211_X1 U21780 ( .C1(n19130), .C2(n18860), .A(n18795), .B(n18794), .ZN(
        P3_U2889) );
  AOI22_X1 U21781 ( .A1(n19132), .A2(n18817), .B1(n19131), .B2(n18798), .ZN(
        n18797) );
  AOI22_X1 U21782 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18799), .B1(
        n19134), .B2(n19143), .ZN(n18796) );
  OAI211_X1 U21783 ( .C1(n19138), .C2(n18860), .A(n18797), .B(n18796), .ZN(
        P3_U2890) );
  INV_X1 U21784 ( .A(n19143), .ZN(n19137) );
  AOI22_X1 U21785 ( .A1(n19142), .A2(n18817), .B1(n19140), .B2(n18798), .ZN(
        n18801) );
  AOI22_X1 U21786 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18799), .B1(
        n19144), .B2(n18865), .ZN(n18800) );
  OAI211_X1 U21787 ( .C1(n19149), .C2(n19137), .A(n18801), .B(n18800), .ZN(
        P3_U2891) );
  NAND2_X1 U21788 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18847), .ZN(
        n18892) );
  INV_X1 U21789 ( .A(n18847), .ZN(n18802) );
  NOR2_X1 U21790 ( .A1(n19091), .A2(n18802), .ZN(n18820) );
  AOI22_X1 U21791 ( .A1(n19093), .A2(n18820), .B1(n19092), .B2(n18817), .ZN(
        n18806) );
  OAI21_X1 U21792 ( .B1(n19189), .B2(n18803), .A(n19061), .ZN(n19094) );
  NAND2_X1 U21793 ( .A1(n18804), .A2(n19094), .ZN(n18821) );
  AOI22_X1 U21794 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18821), .B1(
        n19033), .B2(n18839), .ZN(n18805) );
  OAI211_X1 U21795 ( .C1(n19039), .C2(n18892), .A(n18806), .B(n18805), .ZN(
        P3_U2892) );
  AOI22_X1 U21796 ( .A1(n19040), .A2(n18839), .B1(n19100), .B2(n18820), .ZN(
        n18808) );
  AOI22_X1 U21797 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18821), .B1(
        n19102), .B2(n18885), .ZN(n18807) );
  OAI211_X1 U21798 ( .C1(n19043), .C2(n18824), .A(n18808), .B(n18807), .ZN(
        P3_U2893) );
  AOI22_X1 U21799 ( .A1(n19109), .A2(n18817), .B1(n19107), .B2(n18820), .ZN(
        n18810) );
  AOI22_X1 U21800 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18821), .B1(
        n19108), .B2(n18839), .ZN(n18809) );
  OAI211_X1 U21801 ( .C1(n19112), .C2(n18892), .A(n18810), .B(n18809), .ZN(
        P3_U2894) );
  AOI22_X1 U21802 ( .A1(n19115), .A2(n18817), .B1(n19113), .B2(n18820), .ZN(
        n18812) );
  AOI22_X1 U21803 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18821), .B1(
        n19114), .B2(n18839), .ZN(n18811) );
  OAI211_X1 U21804 ( .C1(n19118), .C2(n18892), .A(n18812), .B(n18811), .ZN(
        P3_U2895) );
  AOI22_X1 U21805 ( .A1(n19120), .A2(n18839), .B1(n19119), .B2(n18820), .ZN(
        n18814) );
  AOI22_X1 U21806 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18821), .B1(
        n19121), .B2(n18885), .ZN(n18813) );
  OAI211_X1 U21807 ( .C1(n19124), .C2(n18824), .A(n18814), .B(n18813), .ZN(
        P3_U2896) );
  AOI22_X1 U21808 ( .A1(n19127), .A2(n18839), .B1(n19125), .B2(n18820), .ZN(
        n18816) );
  AOI22_X1 U21809 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18821), .B1(
        n19126), .B2(n18817), .ZN(n18815) );
  OAI211_X1 U21810 ( .C1(n19130), .C2(n18892), .A(n18816), .B(n18815), .ZN(
        P3_U2897) );
  AOI22_X1 U21811 ( .A1(n19132), .A2(n18839), .B1(n19131), .B2(n18820), .ZN(
        n18819) );
  AOI22_X1 U21812 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18821), .B1(
        n19134), .B2(n18817), .ZN(n18818) );
  OAI211_X1 U21813 ( .C1(n19138), .C2(n18892), .A(n18819), .B(n18818), .ZN(
        P3_U2898) );
  AOI22_X1 U21814 ( .A1(n19142), .A2(n18839), .B1(n19140), .B2(n18820), .ZN(
        n18823) );
  AOI22_X1 U21815 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18821), .B1(
        n19144), .B2(n18885), .ZN(n18822) );
  OAI211_X1 U21816 ( .C1(n19149), .C2(n18824), .A(n18823), .B(n18822), .ZN(
        P3_U2899) );
  NOR2_X2 U21817 ( .A1(n19190), .A2(n18848), .ZN(n18903) );
  NOR2_X1 U21818 ( .A1(n18885), .A2(n18903), .ZN(n18871) );
  NOR2_X1 U21819 ( .A1(n19091), .A2(n18871), .ZN(n18842) );
  AOI22_X1 U21820 ( .A1(n19093), .A2(n18842), .B1(n19092), .B2(n18839), .ZN(
        n18828) );
  OAI21_X1 U21821 ( .B1(n18825), .B2(n19007), .A(n18871), .ZN(n18826) );
  OAI211_X1 U21822 ( .C1(n18903), .C2(n19335), .A(n19010), .B(n18826), .ZN(
        n18843) );
  AOI22_X1 U21823 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18843), .B1(
        n19096), .B2(n18903), .ZN(n18827) );
  OAI211_X1 U21824 ( .C1(n19099), .C2(n18860), .A(n18828), .B(n18827), .ZN(
        P3_U2900) );
  AOI22_X1 U21825 ( .A1(n19040), .A2(n18865), .B1(n19100), .B2(n18842), .ZN(
        n18830) );
  AOI22_X1 U21826 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18843), .B1(
        n19102), .B2(n18903), .ZN(n18829) );
  OAI211_X1 U21827 ( .C1(n19043), .C2(n18846), .A(n18830), .B(n18829), .ZN(
        P3_U2901) );
  INV_X1 U21828 ( .A(n18903), .ZN(n18915) );
  AOI22_X1 U21829 ( .A1(n19108), .A2(n18865), .B1(n19107), .B2(n18842), .ZN(
        n18832) );
  AOI22_X1 U21830 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18843), .B1(
        n19109), .B2(n18839), .ZN(n18831) );
  OAI211_X1 U21831 ( .C1(n19112), .C2(n18915), .A(n18832), .B(n18831), .ZN(
        P3_U2902) );
  AOI22_X1 U21832 ( .A1(n19114), .A2(n18865), .B1(n19113), .B2(n18842), .ZN(
        n18834) );
  AOI22_X1 U21833 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18843), .B1(
        n19115), .B2(n18839), .ZN(n18833) );
  OAI211_X1 U21834 ( .C1(n19118), .C2(n18915), .A(n18834), .B(n18833), .ZN(
        P3_U2903) );
  AOI22_X1 U21835 ( .A1(n19074), .A2(n18839), .B1(n19119), .B2(n18842), .ZN(
        n18836) );
  AOI22_X1 U21836 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18843), .B1(
        n19121), .B2(n18903), .ZN(n18835) );
  OAI211_X1 U21837 ( .C1(n19077), .C2(n18860), .A(n18836), .B(n18835), .ZN(
        P3_U2904) );
  AOI22_X1 U21838 ( .A1(n19126), .A2(n18839), .B1(n19125), .B2(n18842), .ZN(
        n18838) );
  AOI22_X1 U21839 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18843), .B1(
        n19127), .B2(n18865), .ZN(n18837) );
  OAI211_X1 U21840 ( .C1(n19130), .C2(n18915), .A(n18838), .B(n18837), .ZN(
        P3_U2905) );
  AOI22_X1 U21841 ( .A1(n19134), .A2(n18839), .B1(n19131), .B2(n18842), .ZN(
        n18841) );
  AOI22_X1 U21842 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18843), .B1(
        n19132), .B2(n18865), .ZN(n18840) );
  OAI211_X1 U21843 ( .C1(n19138), .C2(n18915), .A(n18841), .B(n18840), .ZN(
        P3_U2906) );
  AOI22_X1 U21844 ( .A1(n19142), .A2(n18865), .B1(n19140), .B2(n18842), .ZN(
        n18845) );
  AOI22_X1 U21845 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18843), .B1(
        n19144), .B2(n18903), .ZN(n18844) );
  OAI211_X1 U21846 ( .C1(n19149), .C2(n18846), .A(n18845), .B(n18844), .ZN(
        P3_U2907) );
  NOR2_X1 U21847 ( .A1(n18848), .A2(n19031), .ZN(n18866) );
  AOI22_X1 U21848 ( .A1(n19093), .A2(n18866), .B1(n19092), .B2(n18865), .ZN(
        n18851) );
  AOI22_X1 U21849 ( .A1(n19036), .A2(n18847), .B1(n18894), .B2(n19034), .ZN(
        n18867) );
  NOR2_X2 U21850 ( .A1(n18849), .A2(n18848), .ZN(n18933) );
  AOI22_X1 U21851 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18867), .B1(
        n18933), .B2(n19096), .ZN(n18850) );
  OAI211_X1 U21852 ( .C1(n19099), .C2(n18892), .A(n18851), .B(n18850), .ZN(
        P3_U2908) );
  AOI22_X1 U21853 ( .A1(n19101), .A2(n18865), .B1(n19100), .B2(n18866), .ZN(
        n18853) );
  AOI22_X1 U21854 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18867), .B1(
        n18933), .B2(n19102), .ZN(n18852) );
  OAI211_X1 U21855 ( .C1(n19106), .C2(n18892), .A(n18853), .B(n18852), .ZN(
        P3_U2909) );
  INV_X1 U21856 ( .A(n18933), .ZN(n18906) );
  AOI22_X1 U21857 ( .A1(n19108), .A2(n18885), .B1(n19107), .B2(n18866), .ZN(
        n18855) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18867), .B1(
        n19109), .B2(n18865), .ZN(n18854) );
  OAI211_X1 U21859 ( .C1(n18906), .C2(n19112), .A(n18855), .B(n18854), .ZN(
        P3_U2910) );
  AOI22_X1 U21860 ( .A1(n19114), .A2(n18885), .B1(n19113), .B2(n18866), .ZN(
        n18857) );
  AOI22_X1 U21861 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18867), .B1(
        n19115), .B2(n18865), .ZN(n18856) );
  OAI211_X1 U21862 ( .C1(n18906), .C2(n19118), .A(n18857), .B(n18856), .ZN(
        P3_U2911) );
  AOI22_X1 U21863 ( .A1(n19120), .A2(n18885), .B1(n19119), .B2(n18866), .ZN(
        n18859) );
  AOI22_X1 U21864 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18867), .B1(
        n18933), .B2(n19121), .ZN(n18858) );
  OAI211_X1 U21865 ( .C1(n19124), .C2(n18860), .A(n18859), .B(n18858), .ZN(
        P3_U2912) );
  AOI22_X1 U21866 ( .A1(n19126), .A2(n18865), .B1(n19125), .B2(n18866), .ZN(
        n18862) );
  AOI22_X1 U21867 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18867), .B1(
        n19127), .B2(n18885), .ZN(n18861) );
  OAI211_X1 U21868 ( .C1(n18906), .C2(n19130), .A(n18862), .B(n18861), .ZN(
        P3_U2913) );
  AOI22_X1 U21869 ( .A1(n19134), .A2(n18865), .B1(n19131), .B2(n18866), .ZN(
        n18864) );
  AOI22_X1 U21870 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18867), .B1(
        n19132), .B2(n18885), .ZN(n18863) );
  OAI211_X1 U21871 ( .C1(n18906), .C2(n19138), .A(n18864), .B(n18863), .ZN(
        P3_U2914) );
  AOI22_X1 U21872 ( .A1(n19140), .A2(n18866), .B1(n18978), .B2(n18865), .ZN(
        n18869) );
  AOI22_X1 U21873 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18867), .B1(
        n18933), .B2(n19144), .ZN(n18868) );
  OAI211_X1 U21874 ( .C1(n18983), .C2(n18892), .A(n18869), .B(n18868), .ZN(
        P3_U2915) );
  NOR2_X1 U21875 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18870), .ZN(
        n18939) );
  NAND2_X1 U21876 ( .A1(n18939), .A2(n19188), .ZN(n18950) );
  INV_X1 U21877 ( .A(n18950), .ZN(n18956) );
  NOR2_X1 U21878 ( .A1(n18956), .A2(n18933), .ZN(n18916) );
  NOR2_X1 U21879 ( .A1(n19091), .A2(n18916), .ZN(n18888) );
  AOI22_X1 U21880 ( .A1(n19033), .A2(n18903), .B1(n19093), .B2(n18888), .ZN(
        n18874) );
  OAI21_X1 U21881 ( .B1(n18871), .B2(n19007), .A(n18916), .ZN(n18872) );
  OAI211_X1 U21882 ( .C1(n18956), .C2(n19335), .A(n19010), .B(n18872), .ZN(
        n18889) );
  AOI22_X1 U21883 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18889), .B1(
        n19092), .B2(n18885), .ZN(n18873) );
  OAI211_X1 U21884 ( .C1(n18950), .C2(n19039), .A(n18874), .B(n18873), .ZN(
        P3_U2916) );
  AOI22_X1 U21885 ( .A1(n19101), .A2(n18885), .B1(n19100), .B2(n18888), .ZN(
        n18876) );
  AOI22_X1 U21886 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18889), .B1(
        n18956), .B2(n19102), .ZN(n18875) );
  OAI211_X1 U21887 ( .C1(n19106), .C2(n18915), .A(n18876), .B(n18875), .ZN(
        P3_U2917) );
  AOI22_X1 U21888 ( .A1(n19108), .A2(n18903), .B1(n19107), .B2(n18888), .ZN(
        n18878) );
  AOI22_X1 U21889 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18889), .B1(
        n19109), .B2(n18885), .ZN(n18877) );
  OAI211_X1 U21890 ( .C1(n18950), .C2(n19112), .A(n18878), .B(n18877), .ZN(
        P3_U2918) );
  AOI22_X1 U21891 ( .A1(n19115), .A2(n18885), .B1(n19113), .B2(n18888), .ZN(
        n18880) );
  AOI22_X1 U21892 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18889), .B1(
        n19114), .B2(n18903), .ZN(n18879) );
  OAI211_X1 U21893 ( .C1(n18950), .C2(n19118), .A(n18880), .B(n18879), .ZN(
        P3_U2919) );
  AOI22_X1 U21894 ( .A1(n19120), .A2(n18903), .B1(n19119), .B2(n18888), .ZN(
        n18882) );
  AOI22_X1 U21895 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18889), .B1(
        n18956), .B2(n19121), .ZN(n18881) );
  OAI211_X1 U21896 ( .C1(n19124), .C2(n18892), .A(n18882), .B(n18881), .ZN(
        P3_U2920) );
  AOI22_X1 U21897 ( .A1(n19126), .A2(n18885), .B1(n19125), .B2(n18888), .ZN(
        n18884) );
  AOI22_X1 U21898 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18889), .B1(
        n19127), .B2(n18903), .ZN(n18883) );
  OAI211_X1 U21899 ( .C1(n18950), .C2(n19130), .A(n18884), .B(n18883), .ZN(
        P3_U2921) );
  AOI22_X1 U21900 ( .A1(n19134), .A2(n18885), .B1(n19131), .B2(n18888), .ZN(
        n18887) );
  AOI22_X1 U21901 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18889), .B1(
        n19132), .B2(n18903), .ZN(n18886) );
  OAI211_X1 U21902 ( .C1(n18950), .C2(n19138), .A(n18887), .B(n18886), .ZN(
        P3_U2922) );
  AOI22_X1 U21903 ( .A1(n19142), .A2(n18903), .B1(n19140), .B2(n18888), .ZN(
        n18891) );
  AOI22_X1 U21904 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18889), .B1(
        n18956), .B2(n19144), .ZN(n18890) );
  OAI211_X1 U21905 ( .C1(n19149), .C2(n18892), .A(n18891), .B(n18890), .ZN(
        P3_U2923) );
  NAND2_X1 U21906 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18939), .ZN(
        n18972) );
  INV_X1 U21907 ( .A(n18939), .ZN(n18893) );
  NOR2_X1 U21908 ( .A1(n19091), .A2(n18893), .ZN(n18911) );
  AOI22_X1 U21909 ( .A1(n19033), .A2(n18933), .B1(n19093), .B2(n18911), .ZN(
        n18896) );
  NAND2_X1 U21910 ( .A1(n18894), .A2(n19094), .ZN(n18912) );
  AOI22_X1 U21911 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18912), .B1(
        n19092), .B2(n18903), .ZN(n18895) );
  OAI211_X1 U21912 ( .C1(n18972), .C2(n19039), .A(n18896), .B(n18895), .ZN(
        P3_U2924) );
  AOI22_X1 U21913 ( .A1(n19101), .A2(n18903), .B1(n19100), .B2(n18911), .ZN(
        n18898) );
  AOI22_X1 U21914 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18912), .B1(
        n18979), .B2(n19102), .ZN(n18897) );
  OAI211_X1 U21915 ( .C1(n18906), .C2(n19106), .A(n18898), .B(n18897), .ZN(
        P3_U2925) );
  AOI22_X1 U21916 ( .A1(n18933), .A2(n19108), .B1(n19107), .B2(n18911), .ZN(
        n18900) );
  AOI22_X1 U21917 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18912), .B1(
        n19109), .B2(n18903), .ZN(n18899) );
  OAI211_X1 U21918 ( .C1(n18972), .C2(n19112), .A(n18900), .B(n18899), .ZN(
        P3_U2926) );
  AOI22_X1 U21919 ( .A1(n19115), .A2(n18903), .B1(n19113), .B2(n18911), .ZN(
        n18902) );
  AOI22_X1 U21920 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18912), .B1(
        n18933), .B2(n19114), .ZN(n18901) );
  OAI211_X1 U21921 ( .C1(n18972), .C2(n19118), .A(n18902), .B(n18901), .ZN(
        P3_U2927) );
  AOI22_X1 U21922 ( .A1(n19074), .A2(n18903), .B1(n19119), .B2(n18911), .ZN(
        n18905) );
  AOI22_X1 U21923 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18912), .B1(
        n18979), .B2(n19121), .ZN(n18904) );
  OAI211_X1 U21924 ( .C1(n18906), .C2(n19077), .A(n18905), .B(n18904), .ZN(
        P3_U2928) );
  AOI22_X1 U21925 ( .A1(n19126), .A2(n18903), .B1(n19125), .B2(n18911), .ZN(
        n18908) );
  AOI22_X1 U21926 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18912), .B1(
        n18933), .B2(n19127), .ZN(n18907) );
  OAI211_X1 U21927 ( .C1(n18972), .C2(n19130), .A(n18908), .B(n18907), .ZN(
        P3_U2929) );
  AOI22_X1 U21928 ( .A1(n18933), .A2(n19132), .B1(n19131), .B2(n18911), .ZN(
        n18910) );
  AOI22_X1 U21929 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18912), .B1(
        n19134), .B2(n18903), .ZN(n18909) );
  OAI211_X1 U21930 ( .C1(n18972), .C2(n19138), .A(n18910), .B(n18909), .ZN(
        P3_U2930) );
  AOI22_X1 U21931 ( .A1(n18933), .A2(n19142), .B1(n19140), .B2(n18911), .ZN(
        n18914) );
  AOI22_X1 U21932 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18912), .B1(
        n18979), .B2(n19144), .ZN(n18913) );
  OAI211_X1 U21933 ( .C1(n19149), .C2(n18915), .A(n18914), .B(n18913), .ZN(
        P3_U2931) );
  NAND2_X1 U21934 ( .A1(n19006), .A2(n18985), .ZN(n19005) );
  AOI21_X1 U21935 ( .B1(n19005), .B2(n18972), .A(n19091), .ZN(n18932) );
  AOI22_X1 U21936 ( .A1(n18933), .A2(n19092), .B1(n19093), .B2(n18932), .ZN(
        n18919) );
  AOI221_X1 U21937 ( .B1(n18916), .B2(n18972), .C1(n19007), .C2(n18972), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18917) );
  OAI21_X1 U21938 ( .B1(n18998), .B2(n18917), .A(n19010), .ZN(n18934) );
  AOI22_X1 U21939 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18934), .B1(
        n18998), .B2(n19096), .ZN(n18918) );
  OAI211_X1 U21940 ( .C1(n19099), .C2(n18950), .A(n18919), .B(n18918), .ZN(
        P3_U2932) );
  AOI22_X1 U21941 ( .A1(n18933), .A2(n19101), .B1(n18932), .B2(n19100), .ZN(
        n18921) );
  AOI22_X1 U21942 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18934), .B1(
        n18998), .B2(n19102), .ZN(n18920) );
  OAI211_X1 U21943 ( .C1(n18950), .C2(n19106), .A(n18921), .B(n18920), .ZN(
        P3_U2933) );
  AOI22_X1 U21944 ( .A1(n18956), .A2(n19108), .B1(n18932), .B2(n19107), .ZN(
        n18923) );
  AOI22_X1 U21945 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18934), .B1(
        n18933), .B2(n19109), .ZN(n18922) );
  OAI211_X1 U21946 ( .C1(n19005), .C2(n19112), .A(n18923), .B(n18922), .ZN(
        P3_U2934) );
  AOI22_X1 U21947 ( .A1(n18956), .A2(n19114), .B1(n18932), .B2(n19113), .ZN(
        n18925) );
  AOI22_X1 U21948 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18934), .B1(
        n18933), .B2(n19115), .ZN(n18924) );
  OAI211_X1 U21949 ( .C1(n19005), .C2(n19118), .A(n18925), .B(n18924), .ZN(
        P3_U2935) );
  AOI22_X1 U21950 ( .A1(n18933), .A2(n19074), .B1(n18932), .B2(n19119), .ZN(
        n18927) );
  AOI22_X1 U21951 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18934), .B1(
        n18998), .B2(n19121), .ZN(n18926) );
  OAI211_X1 U21952 ( .C1(n18950), .C2(n19077), .A(n18927), .B(n18926), .ZN(
        P3_U2936) );
  AOI22_X1 U21953 ( .A1(n18956), .A2(n19127), .B1(n18932), .B2(n19125), .ZN(
        n18929) );
  AOI22_X1 U21954 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18934), .B1(
        n18933), .B2(n19126), .ZN(n18928) );
  OAI211_X1 U21955 ( .C1(n19005), .C2(n19130), .A(n18929), .B(n18928), .ZN(
        P3_U2937) );
  AOI22_X1 U21956 ( .A1(n18956), .A2(n19132), .B1(n18932), .B2(n19131), .ZN(
        n18931) );
  AOI22_X1 U21957 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18934), .B1(
        n18933), .B2(n19134), .ZN(n18930) );
  OAI211_X1 U21958 ( .C1(n19005), .C2(n19138), .A(n18931), .B(n18930), .ZN(
        P3_U2938) );
  AOI22_X1 U21959 ( .A1(n18933), .A2(n18978), .B1(n18932), .B2(n19140), .ZN(
        n18936) );
  AOI22_X1 U21960 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18934), .B1(
        n18998), .B2(n19144), .ZN(n18935) );
  OAI211_X1 U21961 ( .C1(n18950), .C2(n18983), .A(n18936), .B(n18935), .ZN(
        P3_U2939) );
  NAND2_X1 U21962 ( .A1(n18985), .A2(n18937), .ZN(n19030) );
  INV_X1 U21963 ( .A(n18985), .ZN(n18938) );
  NOR2_X1 U21964 ( .A1(n18938), .A2(n19031), .ZN(n18955) );
  AOI22_X1 U21965 ( .A1(n18956), .A2(n19092), .B1(n19093), .B2(n18955), .ZN(
        n18941) );
  AOI22_X1 U21966 ( .A1(n19036), .A2(n18939), .B1(n18985), .B2(n19034), .ZN(
        n18957) );
  AOI22_X1 U21967 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18957), .B1(
        n19033), .B2(n18979), .ZN(n18940) );
  OAI211_X1 U21968 ( .C1(n19039), .C2(n19030), .A(n18941), .B(n18940), .ZN(
        P3_U2940) );
  AOI22_X1 U21969 ( .A1(n18979), .A2(n19040), .B1(n19100), .B2(n18955), .ZN(
        n18943) );
  INV_X1 U21970 ( .A(n19030), .ZN(n19023) );
  AOI22_X1 U21971 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18957), .B1(
        n19102), .B2(n19023), .ZN(n18942) );
  OAI211_X1 U21972 ( .C1(n18950), .C2(n19043), .A(n18943), .B(n18942), .ZN(
        P3_U2941) );
  AOI22_X1 U21973 ( .A1(n18979), .A2(n19108), .B1(n19107), .B2(n18955), .ZN(
        n18945) );
  AOI22_X1 U21974 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18957), .B1(
        n18956), .B2(n19109), .ZN(n18944) );
  OAI211_X1 U21975 ( .C1(n19112), .C2(n19030), .A(n18945), .B(n18944), .ZN(
        P3_U2942) );
  AOI22_X1 U21976 ( .A1(n18979), .A2(n19114), .B1(n19113), .B2(n18955), .ZN(
        n18947) );
  AOI22_X1 U21977 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18957), .B1(
        n18956), .B2(n19115), .ZN(n18946) );
  OAI211_X1 U21978 ( .C1(n19118), .C2(n19030), .A(n18947), .B(n18946), .ZN(
        P3_U2943) );
  AOI22_X1 U21979 ( .A1(n18979), .A2(n19120), .B1(n19119), .B2(n18955), .ZN(
        n18949) );
  AOI22_X1 U21980 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18957), .B1(
        n19121), .B2(n19023), .ZN(n18948) );
  OAI211_X1 U21981 ( .C1(n18950), .C2(n19124), .A(n18949), .B(n18948), .ZN(
        P3_U2944) );
  AOI22_X1 U21982 ( .A1(n18956), .A2(n19126), .B1(n19125), .B2(n18955), .ZN(
        n18952) );
  AOI22_X1 U21983 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18957), .B1(
        n18979), .B2(n19127), .ZN(n18951) );
  OAI211_X1 U21984 ( .C1(n19130), .C2(n19030), .A(n18952), .B(n18951), .ZN(
        P3_U2945) );
  AOI22_X1 U21985 ( .A1(n18956), .A2(n19134), .B1(n19131), .B2(n18955), .ZN(
        n18954) );
  AOI22_X1 U21986 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18957), .B1(
        n18979), .B2(n19132), .ZN(n18953) );
  OAI211_X1 U21987 ( .C1(n19138), .C2(n19030), .A(n18954), .B(n18953), .ZN(
        P3_U2946) );
  AOI22_X1 U21988 ( .A1(n18956), .A2(n18978), .B1(n19140), .B2(n18955), .ZN(
        n18959) );
  AOI22_X1 U21989 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18957), .B1(
        n19144), .B2(n19023), .ZN(n18958) );
  OAI211_X1 U21990 ( .C1(n18972), .C2(n18983), .A(n18959), .B(n18958), .ZN(
        P3_U2947) );
  NAND2_X1 U21991 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18985), .ZN(
        n18984) );
  NOR2_X2 U21992 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18984), .ZN(
        n19052) );
  NOR2_X1 U21993 ( .A1(n19023), .A2(n19052), .ZN(n19008) );
  NOR2_X1 U21994 ( .A1(n19091), .A2(n19008), .ZN(n18977) );
  AOI22_X1 U21995 ( .A1(n18979), .A2(n19092), .B1(n19093), .B2(n18977), .ZN(
        n18963) );
  NOR2_X1 U21996 ( .A1(n18998), .A2(n18979), .ZN(n18960) );
  OAI21_X1 U21997 ( .B1(n18960), .B2(n19007), .A(n19008), .ZN(n18961) );
  OAI211_X1 U21998 ( .C1(n19052), .C2(n19335), .A(n19010), .B(n18961), .ZN(
        n18980) );
  AOI22_X1 U21999 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18980), .B1(
        n19096), .B2(n19052), .ZN(n18962) );
  OAI211_X1 U22000 ( .C1(n19099), .C2(n19005), .A(n18963), .B(n18962), .ZN(
        P3_U2948) );
  AOI22_X1 U22001 ( .A1(n18979), .A2(n19101), .B1(n19100), .B2(n18977), .ZN(
        n18965) );
  AOI22_X1 U22002 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18980), .B1(
        n19102), .B2(n19052), .ZN(n18964) );
  OAI211_X1 U22003 ( .C1(n19005), .C2(n19106), .A(n18965), .B(n18964), .ZN(
        P3_U2949) );
  INV_X1 U22004 ( .A(n19052), .ZN(n19059) );
  AOI22_X1 U22005 ( .A1(n18998), .A2(n19108), .B1(n19107), .B2(n18977), .ZN(
        n18967) );
  AOI22_X1 U22006 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18980), .B1(
        n18979), .B2(n19109), .ZN(n18966) );
  OAI211_X1 U22007 ( .C1(n19112), .C2(n19059), .A(n18967), .B(n18966), .ZN(
        P3_U2950) );
  AOI22_X1 U22008 ( .A1(n18998), .A2(n19114), .B1(n19113), .B2(n18977), .ZN(
        n18969) );
  AOI22_X1 U22009 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18980), .B1(
        n18979), .B2(n19115), .ZN(n18968) );
  OAI211_X1 U22010 ( .C1(n19118), .C2(n19059), .A(n18969), .B(n18968), .ZN(
        P3_U2951) );
  AOI22_X1 U22011 ( .A1(n18998), .A2(n19120), .B1(n19119), .B2(n18977), .ZN(
        n18971) );
  AOI22_X1 U22012 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18980), .B1(
        n19121), .B2(n19052), .ZN(n18970) );
  OAI211_X1 U22013 ( .C1(n18972), .C2(n19124), .A(n18971), .B(n18970), .ZN(
        P3_U2952) );
  AOI22_X1 U22014 ( .A1(n18979), .A2(n19126), .B1(n19125), .B2(n18977), .ZN(
        n18974) );
  AOI22_X1 U22015 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18980), .B1(
        n18998), .B2(n19127), .ZN(n18973) );
  OAI211_X1 U22016 ( .C1(n19130), .C2(n19059), .A(n18974), .B(n18973), .ZN(
        P3_U2953) );
  AOI22_X1 U22017 ( .A1(n18998), .A2(n19132), .B1(n19131), .B2(n18977), .ZN(
        n18976) );
  AOI22_X1 U22018 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18980), .B1(
        n18979), .B2(n19134), .ZN(n18975) );
  OAI211_X1 U22019 ( .C1(n19138), .C2(n19059), .A(n18976), .B(n18975), .ZN(
        P3_U2954) );
  AOI22_X1 U22020 ( .A1(n18979), .A2(n18978), .B1(n19140), .B2(n18977), .ZN(
        n18982) );
  AOI22_X1 U22021 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18980), .B1(
        n19144), .B2(n19052), .ZN(n18981) );
  OAI211_X1 U22022 ( .C1(n19005), .C2(n18983), .A(n18982), .B(n18981), .ZN(
        P3_U2955) );
  INV_X1 U22023 ( .A(n18984), .ZN(n19035) );
  NAND2_X1 U22024 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19035), .ZN(
        n19089) );
  NOR2_X1 U22025 ( .A1(n19091), .A2(n18984), .ZN(n19001) );
  AOI22_X1 U22026 ( .A1(n19033), .A2(n19023), .B1(n19093), .B2(n19001), .ZN(
        n18987) );
  NAND2_X1 U22027 ( .A1(n18985), .A2(n19094), .ZN(n19002) );
  AOI22_X1 U22028 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19002), .B1(
        n18998), .B2(n19092), .ZN(n18986) );
  OAI211_X1 U22029 ( .C1(n19039), .C2(n19089), .A(n18987), .B(n18986), .ZN(
        P3_U2956) );
  AOI22_X1 U22030 ( .A1(n18998), .A2(n19101), .B1(n19100), .B2(n19001), .ZN(
        n18989) );
  AOI22_X1 U22031 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19002), .B1(
        n19102), .B2(n19080), .ZN(n18988) );
  OAI211_X1 U22032 ( .C1(n19106), .C2(n19030), .A(n18989), .B(n18988), .ZN(
        P3_U2957) );
  AOI22_X1 U22033 ( .A1(n18998), .A2(n19109), .B1(n19107), .B2(n19001), .ZN(
        n18991) );
  AOI22_X1 U22034 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19002), .B1(
        n19108), .B2(n19023), .ZN(n18990) );
  OAI211_X1 U22035 ( .C1(n19112), .C2(n19089), .A(n18991), .B(n18990), .ZN(
        P3_U2958) );
  AOI22_X1 U22036 ( .A1(n19114), .A2(n19023), .B1(n19113), .B2(n19001), .ZN(
        n18993) );
  AOI22_X1 U22037 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19002), .B1(
        n18998), .B2(n19115), .ZN(n18992) );
  OAI211_X1 U22038 ( .C1(n19118), .C2(n19089), .A(n18993), .B(n18992), .ZN(
        P3_U2959) );
  AOI22_X1 U22039 ( .A1(n18998), .A2(n19074), .B1(n19119), .B2(n19001), .ZN(
        n18995) );
  AOI22_X1 U22040 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19002), .B1(
        n19121), .B2(n19080), .ZN(n18994) );
  OAI211_X1 U22041 ( .C1(n19077), .C2(n19030), .A(n18995), .B(n18994), .ZN(
        P3_U2960) );
  AOI22_X1 U22042 ( .A1(n19127), .A2(n19023), .B1(n19125), .B2(n19001), .ZN(
        n18997) );
  AOI22_X1 U22043 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19002), .B1(
        n18998), .B2(n19126), .ZN(n18996) );
  OAI211_X1 U22044 ( .C1(n19130), .C2(n19089), .A(n18997), .B(n18996), .ZN(
        P3_U2961) );
  AOI22_X1 U22045 ( .A1(n19132), .A2(n19023), .B1(n19131), .B2(n19001), .ZN(
        n19000) );
  AOI22_X1 U22046 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19002), .B1(
        n18998), .B2(n19134), .ZN(n18999) );
  OAI211_X1 U22047 ( .C1(n19138), .C2(n19089), .A(n19000), .B(n18999), .ZN(
        P3_U2962) );
  AOI22_X1 U22048 ( .A1(n19142), .A2(n19023), .B1(n19140), .B2(n19001), .ZN(
        n19004) );
  AOI22_X1 U22049 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19002), .B1(
        n19144), .B2(n19080), .ZN(n19003) );
  OAI211_X1 U22050 ( .C1(n19005), .C2(n19149), .A(n19004), .B(n19003), .ZN(
        P3_U2963) );
  NAND2_X1 U22051 ( .A1(n19006), .A2(n19095), .ZN(n19148) );
  INV_X1 U22052 ( .A(n19148), .ZN(n19133) );
  NOR2_X1 U22053 ( .A1(n19080), .A2(n19133), .ZN(n19062) );
  NOR2_X1 U22054 ( .A1(n19091), .A2(n19062), .ZN(n19026) );
  AOI22_X1 U22055 ( .A1(n19093), .A2(n19026), .B1(n19092), .B2(n19023), .ZN(
        n19012) );
  OAI21_X1 U22056 ( .B1(n19008), .B2(n19007), .A(n19062), .ZN(n19009) );
  OAI211_X1 U22057 ( .C1(n19133), .C2(n19335), .A(n19010), .B(n19009), .ZN(
        n19027) );
  AOI22_X1 U22058 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19027), .B1(
        n19033), .B2(n19052), .ZN(n19011) );
  OAI211_X1 U22059 ( .C1(n19039), .C2(n19148), .A(n19012), .B(n19011), .ZN(
        P3_U2964) );
  AOI22_X1 U22060 ( .A1(n19040), .A2(n19052), .B1(n19100), .B2(n19026), .ZN(
        n19014) );
  AOI22_X1 U22061 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19027), .B1(
        n19102), .B2(n19133), .ZN(n19013) );
  OAI211_X1 U22062 ( .C1(n19043), .C2(n19030), .A(n19014), .B(n19013), .ZN(
        P3_U2965) );
  AOI22_X1 U22063 ( .A1(n19108), .A2(n19052), .B1(n19107), .B2(n19026), .ZN(
        n19016) );
  AOI22_X1 U22064 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19027), .B1(
        n19109), .B2(n19023), .ZN(n19015) );
  OAI211_X1 U22065 ( .C1(n19112), .C2(n19148), .A(n19016), .B(n19015), .ZN(
        P3_U2966) );
  AOI22_X1 U22066 ( .A1(n19115), .A2(n19023), .B1(n19113), .B2(n19026), .ZN(
        n19018) );
  AOI22_X1 U22067 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19027), .B1(
        n19114), .B2(n19052), .ZN(n19017) );
  OAI211_X1 U22068 ( .C1(n19118), .C2(n19148), .A(n19018), .B(n19017), .ZN(
        P3_U2967) );
  AOI22_X1 U22069 ( .A1(n19074), .A2(n19023), .B1(n19119), .B2(n19026), .ZN(
        n19020) );
  AOI22_X1 U22070 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19027), .B1(
        n19121), .B2(n19133), .ZN(n19019) );
  OAI211_X1 U22071 ( .C1(n19077), .C2(n19059), .A(n19020), .B(n19019), .ZN(
        P3_U2968) );
  AOI22_X1 U22072 ( .A1(n19126), .A2(n19023), .B1(n19125), .B2(n19026), .ZN(
        n19022) );
  AOI22_X1 U22073 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19027), .B1(
        n19127), .B2(n19052), .ZN(n19021) );
  OAI211_X1 U22074 ( .C1(n19130), .C2(n19148), .A(n19022), .B(n19021), .ZN(
        P3_U2969) );
  AOI22_X1 U22075 ( .A1(n19132), .A2(n19052), .B1(n19131), .B2(n19026), .ZN(
        n19025) );
  AOI22_X1 U22076 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19027), .B1(
        n19134), .B2(n19023), .ZN(n19024) );
  OAI211_X1 U22077 ( .C1(n19138), .C2(n19148), .A(n19025), .B(n19024), .ZN(
        P3_U2970) );
  AOI22_X1 U22078 ( .A1(n19142), .A2(n19052), .B1(n19140), .B2(n19026), .ZN(
        n19029) );
  AOI22_X1 U22079 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19027), .B1(
        n19144), .B2(n19133), .ZN(n19028) );
  OAI211_X1 U22080 ( .C1(n19149), .C2(n19030), .A(n19029), .B(n19028), .ZN(
        P3_U2971) );
  INV_X1 U22081 ( .A(n19095), .ZN(n19032) );
  NOR2_X1 U22082 ( .A1(n19032), .A2(n19031), .ZN(n19055) );
  AOI22_X1 U22083 ( .A1(n19033), .A2(n19080), .B1(n19093), .B2(n19055), .ZN(
        n19038) );
  AOI22_X1 U22084 ( .A1(n19036), .A2(n19035), .B1(n19095), .B2(n19034), .ZN(
        n19056) );
  AOI22_X1 U22085 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19056), .B1(
        n19092), .B2(n19052), .ZN(n19037) );
  OAI211_X1 U22086 ( .C1(n19039), .C2(n19105), .A(n19038), .B(n19037), .ZN(
        P3_U2972) );
  AOI22_X1 U22087 ( .A1(n19040), .A2(n19080), .B1(n19100), .B2(n19055), .ZN(
        n19042) );
  AOI22_X1 U22088 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19056), .B1(
        n19102), .B2(n19141), .ZN(n19041) );
  OAI211_X1 U22089 ( .C1(n19043), .C2(n19059), .A(n19042), .B(n19041), .ZN(
        P3_U2973) );
  AOI22_X1 U22090 ( .A1(n19109), .A2(n19052), .B1(n19107), .B2(n19055), .ZN(
        n19045) );
  AOI22_X1 U22091 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19056), .B1(
        n19108), .B2(n19080), .ZN(n19044) );
  OAI211_X1 U22092 ( .C1(n19112), .C2(n19105), .A(n19045), .B(n19044), .ZN(
        P3_U2974) );
  AOI22_X1 U22093 ( .A1(n19114), .A2(n19080), .B1(n19113), .B2(n19055), .ZN(
        n19047) );
  AOI22_X1 U22094 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19056), .B1(
        n19115), .B2(n19052), .ZN(n19046) );
  OAI211_X1 U22095 ( .C1(n19118), .C2(n19105), .A(n19047), .B(n19046), .ZN(
        P3_U2975) );
  AOI22_X1 U22096 ( .A1(n19120), .A2(n19080), .B1(n19119), .B2(n19055), .ZN(
        n19049) );
  AOI22_X1 U22097 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19056), .B1(
        n19121), .B2(n19141), .ZN(n19048) );
  OAI211_X1 U22098 ( .C1(n19124), .C2(n19059), .A(n19049), .B(n19048), .ZN(
        P3_U2976) );
  AOI22_X1 U22099 ( .A1(n19126), .A2(n19052), .B1(n19125), .B2(n19055), .ZN(
        n19051) );
  AOI22_X1 U22100 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19056), .B1(
        n19127), .B2(n19080), .ZN(n19050) );
  OAI211_X1 U22101 ( .C1(n19130), .C2(n19105), .A(n19051), .B(n19050), .ZN(
        P3_U2977) );
  AOI22_X1 U22102 ( .A1(n19134), .A2(n19052), .B1(n19131), .B2(n19055), .ZN(
        n19054) );
  AOI22_X1 U22103 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19056), .B1(
        n19132), .B2(n19080), .ZN(n19053) );
  OAI211_X1 U22104 ( .C1(n19138), .C2(n19105), .A(n19054), .B(n19053), .ZN(
        P3_U2978) );
  AOI22_X1 U22105 ( .A1(n19142), .A2(n19080), .B1(n19140), .B2(n19055), .ZN(
        n19058) );
  AOI22_X1 U22106 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19056), .B1(
        n19144), .B2(n19141), .ZN(n19057) );
  OAI211_X1 U22107 ( .C1(n19149), .C2(n19059), .A(n19058), .B(n19057), .ZN(
        P3_U2979) );
  INV_X1 U22108 ( .A(n19060), .ZN(n19064) );
  NOR2_X1 U22109 ( .A1(n19091), .A2(n19064), .ZN(n19084) );
  AOI22_X1 U22110 ( .A1(n19093), .A2(n19084), .B1(n19092), .B2(n19080), .ZN(
        n19067) );
  OAI22_X1 U22111 ( .A1(n19064), .A2(n19063), .B1(n19062), .B2(n19061), .ZN(
        n19065) );
  OAI21_X1 U22112 ( .B1(n19085), .B2(n19335), .A(n19065), .ZN(n19086) );
  AOI22_X1 U22113 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19086), .B1(
        n19096), .B2(n19085), .ZN(n19066) );
  OAI211_X1 U22114 ( .C1(n19099), .C2(n19148), .A(n19067), .B(n19066), .ZN(
        P3_U2980) );
  AOI22_X1 U22115 ( .A1(n19101), .A2(n19080), .B1(n19100), .B2(n19084), .ZN(
        n19069) );
  AOI22_X1 U22116 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19086), .B1(
        n19102), .B2(n19085), .ZN(n19068) );
  OAI211_X1 U22117 ( .C1(n19106), .C2(n19148), .A(n19069), .B(n19068), .ZN(
        P3_U2981) );
  AOI22_X1 U22118 ( .A1(n19109), .A2(n19080), .B1(n19107), .B2(n19084), .ZN(
        n19071) );
  AOI22_X1 U22119 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19086), .B1(
        n19108), .B2(n19133), .ZN(n19070) );
  OAI211_X1 U22120 ( .C1(n19112), .C2(n19083), .A(n19071), .B(n19070), .ZN(
        P3_U2982) );
  AOI22_X1 U22121 ( .A1(n19115), .A2(n19080), .B1(n19113), .B2(n19084), .ZN(
        n19073) );
  AOI22_X1 U22122 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19086), .B1(
        n19114), .B2(n19133), .ZN(n19072) );
  OAI211_X1 U22123 ( .C1(n19118), .C2(n19083), .A(n19073), .B(n19072), .ZN(
        P3_U2983) );
  AOI22_X1 U22124 ( .A1(n19074), .A2(n19080), .B1(n19119), .B2(n19084), .ZN(
        n19076) );
  AOI22_X1 U22125 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19086), .B1(
        n19121), .B2(n19085), .ZN(n19075) );
  OAI211_X1 U22126 ( .C1(n19077), .C2(n19148), .A(n19076), .B(n19075), .ZN(
        P3_U2984) );
  AOI22_X1 U22127 ( .A1(n19126), .A2(n19080), .B1(n19125), .B2(n19084), .ZN(
        n19079) );
  AOI22_X1 U22128 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19086), .B1(
        n19127), .B2(n19133), .ZN(n19078) );
  OAI211_X1 U22129 ( .C1(n19130), .C2(n19083), .A(n19079), .B(n19078), .ZN(
        P3_U2985) );
  AOI22_X1 U22130 ( .A1(n19132), .A2(n19133), .B1(n19131), .B2(n19084), .ZN(
        n19082) );
  AOI22_X1 U22131 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19086), .B1(
        n19134), .B2(n19080), .ZN(n19081) );
  OAI211_X1 U22132 ( .C1(n19138), .C2(n19083), .A(n19082), .B(n19081), .ZN(
        P3_U2986) );
  AOI22_X1 U22133 ( .A1(n19142), .A2(n19133), .B1(n19140), .B2(n19084), .ZN(
        n19088) );
  AOI22_X1 U22134 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19086), .B1(
        n19144), .B2(n19085), .ZN(n19087) );
  OAI211_X1 U22135 ( .C1(n19149), .C2(n19089), .A(n19088), .B(n19087), .ZN(
        P3_U2987) );
  NOR2_X1 U22136 ( .A1(n19091), .A2(n19090), .ZN(n19139) );
  AOI22_X1 U22137 ( .A1(n19093), .A2(n19139), .B1(n19092), .B2(n19133), .ZN(
        n19098) );
  NAND2_X1 U22138 ( .A1(n19095), .A2(n19094), .ZN(n19145) );
  AOI22_X1 U22139 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19145), .B1(
        n19096), .B2(n19143), .ZN(n19097) );
  OAI211_X1 U22140 ( .C1(n19099), .C2(n19105), .A(n19098), .B(n19097), .ZN(
        P3_U2988) );
  AOI22_X1 U22141 ( .A1(n19101), .A2(n19133), .B1(n19100), .B2(n19139), .ZN(
        n19104) );
  AOI22_X1 U22142 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19145), .B1(
        n19102), .B2(n19143), .ZN(n19103) );
  OAI211_X1 U22143 ( .C1(n19106), .C2(n19105), .A(n19104), .B(n19103), .ZN(
        P3_U2989) );
  AOI22_X1 U22144 ( .A1(n19108), .A2(n19141), .B1(n19107), .B2(n19139), .ZN(
        n19111) );
  AOI22_X1 U22145 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19145), .B1(
        n19109), .B2(n19133), .ZN(n19110) );
  OAI211_X1 U22146 ( .C1(n19112), .C2(n19137), .A(n19111), .B(n19110), .ZN(
        P3_U2990) );
  AOI22_X1 U22147 ( .A1(n19114), .A2(n19141), .B1(n19113), .B2(n19139), .ZN(
        n19117) );
  AOI22_X1 U22148 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19145), .B1(
        n19115), .B2(n19133), .ZN(n19116) );
  OAI211_X1 U22149 ( .C1(n19118), .C2(n19137), .A(n19117), .B(n19116), .ZN(
        P3_U2991) );
  AOI22_X1 U22150 ( .A1(n19120), .A2(n19141), .B1(n19119), .B2(n19139), .ZN(
        n19123) );
  AOI22_X1 U22151 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19145), .B1(
        n19121), .B2(n19143), .ZN(n19122) );
  OAI211_X1 U22152 ( .C1(n19124), .C2(n19148), .A(n19123), .B(n19122), .ZN(
        P3_U2992) );
  AOI22_X1 U22153 ( .A1(n19126), .A2(n19133), .B1(n19125), .B2(n19139), .ZN(
        n19129) );
  AOI22_X1 U22154 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19145), .B1(
        n19127), .B2(n19141), .ZN(n19128) );
  OAI211_X1 U22155 ( .C1(n19130), .C2(n19137), .A(n19129), .B(n19128), .ZN(
        P3_U2993) );
  AOI22_X1 U22156 ( .A1(n19132), .A2(n19141), .B1(n19131), .B2(n19139), .ZN(
        n19136) );
  AOI22_X1 U22157 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19145), .B1(
        n19134), .B2(n19133), .ZN(n19135) );
  OAI211_X1 U22158 ( .C1(n19138), .C2(n19137), .A(n19136), .B(n19135), .ZN(
        P3_U2994) );
  AOI22_X1 U22159 ( .A1(n19142), .A2(n19141), .B1(n19140), .B2(n19139), .ZN(
        n19147) );
  AOI22_X1 U22160 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19145), .B1(
        n19144), .B2(n19143), .ZN(n19146) );
  OAI211_X1 U22161 ( .C1(n19149), .C2(n19148), .A(n19147), .B(n19146), .ZN(
        P3_U2995) );
  NOR2_X1 U22162 ( .A1(n10298), .A2(n19150), .ZN(n19151) );
  OAI222_X1 U22163 ( .A1(n19155), .A2(n19154), .B1(n19153), .B2(n19152), .C1(
        n19151), .C2(n9744), .ZN(n19351) );
  OAI21_X1 U22164 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n19156), .ZN(n19157) );
  OAI211_X1 U22165 ( .C1(n19181), .C2(n19203), .A(n19158), .B(n19157), .ZN(
        n19201) );
  NAND2_X1 U22166 ( .A1(n19325), .A2(n19179), .ZN(n19159) );
  NAND2_X1 U22167 ( .A1(n19184), .A2(n12709), .ZN(n19185) );
  AOI22_X1 U22168 ( .A1(n10298), .A2(n19159), .B1(n19172), .B2(n19185), .ZN(
        n19160) );
  NOR2_X1 U22169 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19160), .ZN(
        n19314) );
  AOI21_X1 U22170 ( .B1(n19163), .B2(n19162), .A(n19161), .ZN(n19168) );
  OAI21_X1 U22171 ( .B1(n19184), .B2(n19172), .A(n19168), .ZN(n19164) );
  AOI22_X1 U22172 ( .A1(n19325), .A2(n19179), .B1(n19165), .B2(n19164), .ZN(
        n19315) );
  NAND2_X1 U22173 ( .A1(n19181), .A2(n19315), .ZN(n19166) );
  AOI22_X1 U22174 ( .A1(n19181), .A2(n19314), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19166), .ZN(n19200) );
  AOI221_X1 U22175 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19168), 
        .C1(n19167), .C2(n19168), .A(n19325), .ZN(n19180) );
  NOR2_X1 U22176 ( .A1(n19169), .A2(n12709), .ZN(n19171) );
  OAI211_X1 U22177 ( .C1(n19171), .C2(n19170), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n19325), .ZN(n19176) );
  AOI211_X1 U22178 ( .C1(n19325), .C2(n12710), .A(n19173), .B(n19172), .ZN(
        n19174) );
  INV_X1 U22179 ( .A(n19174), .ZN(n19175) );
  OAI211_X1 U22180 ( .C1(n19323), .C2(n19177), .A(n19176), .B(n19175), .ZN(
        n19178) );
  AOI21_X1 U22181 ( .B1(n19180), .B2(n19179), .A(n19178), .ZN(n19321) );
  AOI22_X1 U22182 ( .A1(n19191), .A2(n19325), .B1(n19321), .B2(n19181), .ZN(
        n19195) );
  NOR2_X1 U22183 ( .A1(n19183), .A2(n19182), .ZN(n19187) );
  AOI22_X1 U22184 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19184), .B1(
        n19187), .B2(n12709), .ZN(n19336) );
  INV_X1 U22185 ( .A(n19185), .ZN(n19186) );
  OAI22_X1 U22186 ( .A1(n19187), .A2(n19326), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19186), .ZN(n19331) );
  OAI221_X1 U22187 ( .B1(n19195), .B2(n19194), .C1(n19193), .C2(n19192), .A(
        n19197), .ZN(n19199) );
  AOI21_X1 U22188 ( .B1(n19197), .B2(n19196), .A(n19195), .ZN(n19198) );
  INV_X1 U22189 ( .A(n19361), .ZN(n19355) );
  AOI22_X1 U22190 ( .A1(n19217), .A2(n19355), .B1(n19204), .B2(n19203), .ZN(
        n19210) );
  NOR2_X1 U22191 ( .A1(n19207), .A2(n19215), .ZN(n19312) );
  OAI211_X1 U22192 ( .C1(P3_STATE2_REG_2__SCAN_IN), .C2(n19361), .A(n19312), 
        .B(n19208), .ZN(n19219) );
  OAI22_X1 U22193 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19210), .B1(n19209), 
        .B2(n19219), .ZN(n19211) );
  OAI21_X1 U22194 ( .B1(n19213), .B2(n19212), .A(n19211), .ZN(P3_U2996) );
  NOR4_X1 U22195 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19215), .A3(n19214), 
        .A4(n19361), .ZN(n19221) );
  AOI211_X1 U22196 ( .C1(n19355), .C2(n19217), .A(n19216), .B(n19221), .ZN(
        n19218) );
  OAI21_X1 U22197 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n19219), .A(n19218), 
        .ZN(P3_U2997) );
  NOR2_X1 U22198 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19363) );
  NOR4_X1 U22199 ( .A1(n19363), .A2(n19222), .A3(n19221), .A4(n19220), .ZN(
        P3_U2998) );
  AND2_X1 U22200 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19223), .ZN(
        P3_U2999) );
  INV_X1 U22201 ( .A(P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n21333) );
  NOR2_X1 U22202 ( .A1(n21333), .A2(n19310), .ZN(P3_U3000) );
  AND2_X1 U22203 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19223), .ZN(
        P3_U3001) );
  AND2_X1 U22204 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19223), .ZN(
        P3_U3002) );
  AND2_X1 U22205 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19223), .ZN(
        P3_U3003) );
  AND2_X1 U22206 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19223), .ZN(
        P3_U3004) );
  AND2_X1 U22207 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19223), .ZN(
        P3_U3005) );
  AND2_X1 U22208 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19223), .ZN(
        P3_U3006) );
  AND2_X1 U22209 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19223), .ZN(
        P3_U3007) );
  AND2_X1 U22210 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19223), .ZN(
        P3_U3008) );
  AND2_X1 U22211 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19223), .ZN(
        P3_U3009) );
  AND2_X1 U22212 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19223), .ZN(
        P3_U3010) );
  AND2_X1 U22213 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19223), .ZN(
        P3_U3011) );
  AND2_X1 U22214 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19223), .ZN(
        P3_U3012) );
  AND2_X1 U22215 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19223), .ZN(
        P3_U3013) );
  AND2_X1 U22216 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19223), .ZN(
        P3_U3014) );
  AND2_X1 U22217 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19223), .ZN(
        P3_U3015) );
  AND2_X1 U22218 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19223), .ZN(
        P3_U3016) );
  AND2_X1 U22219 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19223), .ZN(
        P3_U3017) );
  AND2_X1 U22220 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19223), .ZN(
        P3_U3018) );
  AND2_X1 U22221 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19223), .ZN(
        P3_U3019) );
  AND2_X1 U22222 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19223), .ZN(
        P3_U3020) );
  AND2_X1 U22223 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19223), .ZN(P3_U3021) );
  AND2_X1 U22224 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19223), .ZN(P3_U3022) );
  AND2_X1 U22225 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19223), .ZN(P3_U3023) );
  AND2_X1 U22226 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19223), .ZN(P3_U3024) );
  AND2_X1 U22227 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19223), .ZN(P3_U3025) );
  AND2_X1 U22228 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19223), .ZN(P3_U3026) );
  AND2_X1 U22229 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19223), .ZN(P3_U3027) );
  AND2_X1 U22230 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19223), .ZN(P3_U3028) );
  OAI21_X1 U22231 ( .B1(n19224), .B2(n21090), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19225) );
  AOI22_X1 U22232 ( .A1(n19237), .A2(n19240), .B1(n19368), .B2(n19225), .ZN(
        n19226) );
  INV_X1 U22233 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n21318) );
  NAND3_X1 U22234 ( .A1(NA), .A2(n19237), .A3(n21318), .ZN(n19231) );
  OAI211_X1 U22235 ( .C1(n19361), .C2(n19230), .A(n19226), .B(n19231), .ZN(
        P3_U3029) );
  NOR2_X1 U22236 ( .A1(n19240), .A2(n21090), .ZN(n19235) );
  NOR2_X1 U22237 ( .A1(n19237), .A2(n19235), .ZN(n19227) );
  NOR2_X1 U22238 ( .A1(n19361), .A2(n21318), .ZN(n19232) );
  AOI21_X1 U22239 ( .B1(n19227), .B2(P3_REQUESTPENDING_REG_SCAN_IN), .A(n19232), .ZN(n19229) );
  INV_X1 U22240 ( .A(n19228), .ZN(n19358) );
  OAI211_X1 U22241 ( .C1(n21090), .C2(n19230), .A(n19229), .B(n19358), .ZN(
        P3_U3030) );
  AOI21_X1 U22242 ( .B1(n19237), .B2(n19231), .A(n19232), .ZN(n19238) );
  INV_X1 U22243 ( .A(n19232), .ZN(n19233) );
  OAI22_X1 U22244 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19233), .ZN(n19234) );
  OAI22_X1 U22245 ( .A1(n19235), .A2(n19234), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19236) );
  OAI22_X1 U22246 ( .A1(n19238), .A2(n19240), .B1(n19237), .B2(n19236), .ZN(
        P3_U3031) );
  INV_X2 U22247 ( .A(n19239), .ZN(n19300) );
  INV_X1 U22248 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19242) );
  NAND2_X1 U22249 ( .A1(n19349), .A2(n19240), .ZN(n19295) );
  CLKBUF_X1 U22250 ( .A(n19295), .Z(n19296) );
  OAI222_X1 U22251 ( .A1(n19342), .A2(n19300), .B1(n19241), .B2(n19349), .C1(
        n19242), .C2(n19296), .ZN(P3_U3032) );
  OAI222_X1 U22252 ( .A1(n19296), .A2(n19244), .B1(n19243), .B2(n19349), .C1(
        n19242), .C2(n19300), .ZN(P3_U3033) );
  OAI222_X1 U22253 ( .A1(n19296), .A2(n19246), .B1(n19245), .B2(n19349), .C1(
        n19244), .C2(n19300), .ZN(P3_U3034) );
  OAI222_X1 U22254 ( .A1(n19296), .A2(n21236), .B1(n19247), .B2(n19349), .C1(
        n19246), .C2(n19300), .ZN(P3_U3035) );
  OAI222_X1 U22255 ( .A1(n19296), .A2(n19249), .B1(n19248), .B2(n19349), .C1(
        n21236), .C2(n19300), .ZN(P3_U3036) );
  OAI222_X1 U22256 ( .A1(n19296), .A2(n19251), .B1(n19250), .B2(n19349), .C1(
        n19249), .C2(n19300), .ZN(P3_U3037) );
  OAI222_X1 U22257 ( .A1(n19295), .A2(n19254), .B1(n19252), .B2(n19349), .C1(
        n19251), .C2(n19300), .ZN(P3_U3038) );
  OAI222_X1 U22258 ( .A1(n19254), .A2(n19300), .B1(n19253), .B2(n19349), .C1(
        n19255), .C2(n19296), .ZN(P3_U3039) );
  OAI222_X1 U22259 ( .A1(n19296), .A2(n19257), .B1(n19256), .B2(n19349), .C1(
        n19255), .C2(n19300), .ZN(P3_U3040) );
  OAI222_X1 U22260 ( .A1(n19296), .A2(n19259), .B1(n19258), .B2(n19349), .C1(
        n19257), .C2(n19300), .ZN(P3_U3041) );
  OAI222_X1 U22261 ( .A1(n19296), .A2(n19260), .B1(n21291), .B2(n19349), .C1(
        n19259), .C2(n19300), .ZN(P3_U3042) );
  OAI222_X1 U22262 ( .A1(n19296), .A2(n21260), .B1(n19261), .B2(n19349), .C1(
        n19260), .C2(n19300), .ZN(P3_U3043) );
  OAI222_X1 U22263 ( .A1(n19296), .A2(n19263), .B1(n19262), .B2(n19349), .C1(
        n21260), .C2(n19300), .ZN(P3_U3044) );
  OAI222_X1 U22264 ( .A1(n19295), .A2(n19265), .B1(n19264), .B2(n19349), .C1(
        n19263), .C2(n19300), .ZN(P3_U3045) );
  INV_X1 U22265 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19267) );
  OAI222_X1 U22266 ( .A1(n19295), .A2(n19267), .B1(n19266), .B2(n19349), .C1(
        n19265), .C2(n19300), .ZN(P3_U3046) );
  OAI222_X1 U22267 ( .A1(n19295), .A2(n19270), .B1(n19268), .B2(n19349), .C1(
        n19267), .C2(n19300), .ZN(P3_U3047) );
  OAI222_X1 U22268 ( .A1(n19270), .A2(n19300), .B1(n19269), .B2(n19349), .C1(
        n19271), .C2(n19296), .ZN(P3_U3048) );
  OAI222_X1 U22269 ( .A1(n19295), .A2(n19273), .B1(n19272), .B2(n19349), .C1(
        n19271), .C2(n19300), .ZN(P3_U3049) );
  OAI222_X1 U22270 ( .A1(n19295), .A2(n19275), .B1(n19274), .B2(n19349), .C1(
        n19273), .C2(n19300), .ZN(P3_U3050) );
  OAI222_X1 U22271 ( .A1(n19295), .A2(n19277), .B1(n19276), .B2(n19349), .C1(
        n19275), .C2(n19300), .ZN(P3_U3051) );
  OAI222_X1 U22272 ( .A1(n19295), .A2(n19279), .B1(n19278), .B2(n19349), .C1(
        n19277), .C2(n19300), .ZN(P3_U3052) );
  OAI222_X1 U22273 ( .A1(n19296), .A2(n19281), .B1(n19280), .B2(n19349), .C1(
        n19279), .C2(n19300), .ZN(P3_U3053) );
  OAI222_X1 U22274 ( .A1(n19296), .A2(n19284), .B1(n19282), .B2(n19349), .C1(
        n19281), .C2(n19300), .ZN(P3_U3054) );
  OAI222_X1 U22275 ( .A1(n19284), .A2(n19300), .B1(n19283), .B2(n19349), .C1(
        n19285), .C2(n19296), .ZN(P3_U3055) );
  OAI222_X1 U22276 ( .A1(n19296), .A2(n19287), .B1(n19286), .B2(n19349), .C1(
        n19285), .C2(n19300), .ZN(P3_U3056) );
  OAI222_X1 U22277 ( .A1(n19296), .A2(n19289), .B1(n19288), .B2(n19349), .C1(
        n19287), .C2(n19300), .ZN(P3_U3057) );
  OAI222_X1 U22278 ( .A1(n19296), .A2(n19291), .B1(n19290), .B2(n19349), .C1(
        n19289), .C2(n19300), .ZN(P3_U3058) );
  OAI222_X1 U22279 ( .A1(n19296), .A2(n19293), .B1(n19292), .B2(n19349), .C1(
        n19291), .C2(n19300), .ZN(P3_U3059) );
  OAI222_X1 U22280 ( .A1(n19295), .A2(n19299), .B1(n19294), .B2(n19349), .C1(
        n19293), .C2(n19300), .ZN(P3_U3060) );
  OAI222_X1 U22281 ( .A1(n19300), .A2(n19299), .B1(n19298), .B2(n19349), .C1(
        n19297), .C2(n19296), .ZN(P3_U3061) );
  INV_X1 U22282 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n19301) );
  AOI22_X1 U22283 ( .A1(n19349), .A2(n19302), .B1(n19301), .B2(n19368), .ZN(
        P3_U3274) );
  INV_X1 U22284 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19343) );
  INV_X1 U22285 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n19303) );
  AOI22_X1 U22286 ( .A1(n19349), .A2(n19343), .B1(n19303), .B2(n19368), .ZN(
        P3_U3275) );
  INV_X1 U22287 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n19304) );
  AOI22_X1 U22288 ( .A1(n19349), .A2(n19305), .B1(n19304), .B2(n19368), .ZN(
        P3_U3276) );
  INV_X1 U22289 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21294) );
  INV_X1 U22290 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n19306) );
  AOI22_X1 U22291 ( .A1(n19349), .A2(n21294), .B1(n19306), .B2(n19368), .ZN(
        P3_U3277) );
  OAI21_X1 U22292 ( .B1(n19310), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19308), 
        .ZN(n19307) );
  INV_X1 U22293 ( .A(n19307), .ZN(P3_U3280) );
  OAI21_X1 U22294 ( .B1(n19310), .B2(n19309), .A(n19308), .ZN(P3_U3281) );
  OAI21_X1 U22295 ( .B1(n19312), .B2(n19335), .A(n19311), .ZN(P3_U3282) );
  AOI22_X1 U22296 ( .A1(n19330), .A2(n19314), .B1(n19337), .B2(n19313), .ZN(
        n19318) );
  INV_X1 U22297 ( .A(n19315), .ZN(n19316) );
  AOI21_X1 U22298 ( .B1(n19330), .B2(n19316), .A(n19340), .ZN(n19317) );
  OAI22_X1 U22299 ( .A1(n19340), .A2(n19318), .B1(n19317), .B2(n17437), .ZN(
        P3_U3285) );
  NAND2_X1 U22300 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19334) );
  AOI22_X1 U22301 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n19320), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n19319), .ZN(n19328) );
  OAI22_X1 U22302 ( .A1(n19321), .A2(n19370), .B1(n19334), .B2(n19328), .ZN(
        n19322) );
  AOI21_X1 U22303 ( .B1(n19337), .B2(n19323), .A(n19322), .ZN(n19324) );
  AOI22_X1 U22304 ( .A1(n19340), .A2(n19325), .B1(n19324), .B2(n19332), .ZN(
        P3_U3288) );
  INV_X1 U22305 ( .A(n19326), .ZN(n19329) );
  INV_X1 U22306 ( .A(n19334), .ZN(n19327) );
  AOI222_X1 U22307 ( .A1(n19331), .A2(n19330), .B1(n19337), .B2(n19329), .C1(
        n19328), .C2(n19327), .ZN(n19333) );
  AOI22_X1 U22308 ( .A1(n19340), .A2(n12710), .B1(n19333), .B2(n19332), .ZN(
        P3_U3289) );
  OAI221_X1 U22309 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n19336), .C1(
        P3_STATE2_REG_1__SCAN_IN), .C2(n19335), .A(n19334), .ZN(n19339) );
  AOI21_X1 U22310 ( .B1(n12709), .B2(n19337), .A(n19340), .ZN(n19338) );
  AOI22_X1 U22311 ( .A1(n12709), .A2(n19340), .B1(n19339), .B2(n19338), .ZN(
        P3_U3290) );
  AOI21_X1 U22312 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19341) );
  OAI22_X1 U22313 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n19342), .B1(
        P3_REIP_REG_1__SCAN_IN), .B2(n19341), .ZN(n19344) );
  AOI22_X1 U22314 ( .A1(n19347), .A2(n19344), .B1(n19343), .B2(n19345), .ZN(
        P3_U3292) );
  NOR2_X1 U22315 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n19346) );
  AOI22_X1 U22316 ( .A1(n19347), .A2(n19346), .B1(n21294), .B2(n19345), .ZN(
        P3_U3293) );
  INV_X1 U22317 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19348) );
  AOI22_X1 U22318 ( .A1(n19349), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19348), 
        .B2(n19368), .ZN(P3_U3294) );
  MUX2_X1 U22319 ( .A(P3_MORE_REG_SCAN_IN), .B(n19351), .S(n19350), .Z(
        P3_U3295) );
  OAI22_X1 U22320 ( .A1(n19355), .A2(n19354), .B1(n19353), .B2(n19352), .ZN(
        n19356) );
  NOR2_X1 U22321 ( .A1(n19357), .A2(n19356), .ZN(n19367) );
  AOI21_X1 U22322 ( .B1(n19360), .B2(n19359), .A(n19358), .ZN(n19362) );
  OAI211_X1 U22323 ( .C1(n19371), .C2(n19362), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19361), .ZN(n19364) );
  AOI21_X1 U22324 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19364), .A(n19363), 
        .ZN(n19366) );
  NAND2_X1 U22325 ( .A1(n19367), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19365) );
  OAI21_X1 U22326 ( .B1(n19367), .B2(n19366), .A(n19365), .ZN(P3_U3296) );
  OAI22_X1 U22327 ( .A1(n19368), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n19349), .ZN(n19369) );
  INV_X1 U22328 ( .A(n19369), .ZN(P3_U3297) );
  OAI21_X1 U22329 ( .B1(n19370), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n19372), 
        .ZN(n19375) );
  OAI22_X1 U22330 ( .A1(n19375), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19372), 
        .B2(n19371), .ZN(n19373) );
  INV_X1 U22331 ( .A(n19373), .ZN(P3_U3298) );
  OAI21_X1 U22332 ( .B1(n19375), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n19374), 
        .ZN(n19376) );
  INV_X1 U22333 ( .A(n19376), .ZN(P3_U3299) );
  INV_X1 U22334 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19378) );
  NAND2_X1 U22335 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n21286), .ZN(n20175) );
  NOR2_X1 U22336 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n20171) );
  INV_X1 U22337 ( .A(n20171), .ZN(n19377) );
  OAI21_X1 U22338 ( .B1(n20167), .B2(n20175), .A(n19377), .ZN(n20250) );
  OAI21_X1 U22339 ( .B1(n20167), .B2(n19378), .A(n20165), .ZN(P2_U2815) );
  AOI221_X1 U22340 ( .B1(P2_STATE_REG_1__SCAN_IN), .B2(n20167), .C1(n21286), 
        .C2(n20167), .A(P2_D_C_N_REG_SCAN_IN), .ZN(n19379) );
  AOI21_X1 U22341 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n20287), .A(n19379), 
        .ZN(P2_U2817) );
  OAI21_X1 U22342 ( .B1(n19380), .B2(BS16), .A(n20250), .ZN(n20248) );
  OAI21_X1 U22343 ( .B1(n20250), .B2(n20036), .A(n20248), .ZN(P2_U2818) );
  NOR2_X1 U22344 ( .A1(n19382), .A2(n19381), .ZN(n20282) );
  OAI21_X1 U22345 ( .B1(n20282), .B2(n11751), .A(n19383), .ZN(P2_U2819) );
  NOR4_X1 U22346 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19387) );
  NOR4_X1 U22347 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19386) );
  NOR4_X1 U22348 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19385) );
  NOR4_X1 U22349 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19384) );
  NAND4_X1 U22350 ( .A1(n19387), .A2(n19386), .A3(n19385), .A4(n19384), .ZN(
        n19393) );
  NOR4_X1 U22351 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19391) );
  AOI211_X1 U22352 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_13__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19390) );
  NOR4_X1 U22353 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19389) );
  NOR4_X1 U22354 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19388) );
  NAND4_X1 U22355 ( .A1(n19391), .A2(n19390), .A3(n19389), .A4(n19388), .ZN(
        n19392) );
  NOR2_X1 U22356 ( .A1(n19393), .A2(n19392), .ZN(n19401) );
  INV_X1 U22357 ( .A(n19401), .ZN(n19400) );
  NOR2_X1 U22358 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19400), .ZN(n19394) );
  INV_X1 U22359 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20246) );
  AOI22_X1 U22360 ( .A1(n19394), .A2(n19395), .B1(n19400), .B2(n20246), .ZN(
        P2_U2820) );
  OR3_X1 U22361 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19399) );
  INV_X1 U22362 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20244) );
  AOI22_X1 U22363 ( .A1(n19394), .A2(n19399), .B1(n19400), .B2(n20244), .ZN(
        P2_U2821) );
  INV_X1 U22364 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20249) );
  NAND2_X1 U22365 ( .A1(n19394), .A2(n20249), .ZN(n19398) );
  OAI21_X1 U22366 ( .B1(n20184), .B2(n19395), .A(n19401), .ZN(n19396) );
  OAI21_X1 U22367 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19401), .A(n19396), 
        .ZN(n19397) );
  OAI221_X1 U22368 ( .B1(n19398), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19398), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19397), .ZN(P2_U2822) );
  INV_X1 U22369 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20242) );
  OAI221_X1 U22370 ( .B1(n19401), .B2(n20242), .C1(n19400), .C2(n19399), .A(
        n19398), .ZN(P2_U2823) );
  AOI21_X1 U22371 ( .B1(n19402), .B2(P2_REIP_REG_6__SCAN_IN), .A(n16434), .ZN(
        n19403) );
  OAI21_X1 U22372 ( .B1(n19404), .B2(n21330), .A(n19403), .ZN(n19405) );
  AOI21_X1 U22373 ( .B1(n19407), .B2(n19406), .A(n19405), .ZN(n19423) );
  NAND2_X1 U22374 ( .A1(n19408), .A2(n19411), .ZN(n19410) );
  MUX2_X1 U22375 ( .A(n19411), .B(n19410), .S(n19409), .Z(n19421) );
  AND2_X1 U22376 ( .A1(n19413), .A2(n19412), .ZN(n19420) );
  NAND2_X1 U22377 ( .A1(n19415), .A2(n19414), .ZN(n19418) );
  NAND2_X1 U22378 ( .A1(n19416), .A2(n13130), .ZN(n19417) );
  NAND2_X1 U22379 ( .A1(n19418), .A2(n19417), .ZN(n19419) );
  AOI21_X1 U22380 ( .B1(n19421), .B2(n19420), .A(n19419), .ZN(n19422) );
  OAI211_X1 U22381 ( .C1(n16437), .C2(n19424), .A(n19423), .B(n19422), .ZN(
        P2_U2849) );
  AOI22_X1 U22382 ( .A1(n20259), .A2(n19433), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19431), .ZN(n19430) );
  OAI21_X1 U22383 ( .B1(n19427), .B2(n19426), .A(n19425), .ZN(n19428) );
  NAND2_X1 U22384 ( .A1(n19428), .A2(n19437), .ZN(n19429) );
  OAI211_X1 U22385 ( .C1(n19547), .C2(n19441), .A(n19430), .B(n19429), .ZN(
        P2_U2916) );
  AOI22_X1 U22386 ( .A1(n19433), .A2(n19432), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19431), .ZN(n19440) );
  OAI21_X1 U22387 ( .B1(n19436), .B2(n19435), .A(n19434), .ZN(n19438) );
  NAND2_X1 U22388 ( .A1(n19438), .A2(n19437), .ZN(n19439) );
  OAI211_X1 U22389 ( .C1(n19497), .C2(n19441), .A(n19440), .B(n19439), .ZN(
        P2_U2918) );
  NOR2_X1 U22390 ( .A1(n19445), .A2(n19442), .ZN(P2_U2920) );
  AOI22_X1 U22391 ( .A1(n19443), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n19476), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n19444) );
  OAI21_X1 U22392 ( .B1(n21339), .B2(n19445), .A(n19444), .ZN(P2_U2927) );
  AOI22_X1 U22393 ( .A1(n19477), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n19476), 
        .B2(P2_LWORD_REG_15__SCAN_IN), .ZN(n19446) );
  OAI21_X1 U22394 ( .B1(n19447), .B2(n19479), .A(n19446), .ZN(P2_U2936) );
  AOI22_X1 U22395 ( .A1(n19477), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n19476), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19448) );
  OAI21_X1 U22396 ( .B1(n19449), .B2(n19479), .A(n19448), .ZN(P2_U2937) );
  AOI22_X1 U22397 ( .A1(n19477), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n19476), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n19450) );
  OAI21_X1 U22398 ( .B1(n19451), .B2(n19479), .A(n19450), .ZN(P2_U2938) );
  AOI22_X1 U22399 ( .A1(n19477), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n19476), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n19452) );
  OAI21_X1 U22400 ( .B1(n19453), .B2(n19479), .A(n19452), .ZN(P2_U2939) );
  AOI22_X1 U22401 ( .A1(n19477), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n19476), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n19454) );
  OAI21_X1 U22402 ( .B1(n19455), .B2(n19479), .A(n19454), .ZN(P2_U2940) );
  AOI22_X1 U22403 ( .A1(n19477), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n19476), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n19456) );
  OAI21_X1 U22404 ( .B1(n19457), .B2(n19479), .A(n19456), .ZN(P2_U2941) );
  AOI22_X1 U22405 ( .A1(n19477), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n19476), 
        .B2(P2_LWORD_REG_9__SCAN_IN), .ZN(n19458) );
  OAI21_X1 U22406 ( .B1(n19459), .B2(n19479), .A(n19458), .ZN(P2_U2942) );
  INV_X1 U22407 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19461) );
  AOI22_X1 U22408 ( .A1(n19477), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n19476), 
        .B2(P2_LWORD_REG_8__SCAN_IN), .ZN(n19460) );
  OAI21_X1 U22409 ( .B1(n19461), .B2(n19479), .A(n19460), .ZN(P2_U2943) );
  AOI22_X1 U22410 ( .A1(n19477), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n19476), 
        .B2(P2_LWORD_REG_7__SCAN_IN), .ZN(n19462) );
  OAI21_X1 U22411 ( .B1(n19463), .B2(n19479), .A(n19462), .ZN(P2_U2944) );
  AOI22_X1 U22412 ( .A1(n19477), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n19476), 
        .B2(P2_LWORD_REG_6__SCAN_IN), .ZN(n19464) );
  OAI21_X1 U22413 ( .B1(n19465), .B2(n19479), .A(n19464), .ZN(P2_U2945) );
  INV_X1 U22414 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19467) );
  AOI22_X1 U22415 ( .A1(n19477), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n19476), 
        .B2(P2_LWORD_REG_5__SCAN_IN), .ZN(n19466) );
  OAI21_X1 U22416 ( .B1(n19467), .B2(n19479), .A(n19466), .ZN(P2_U2946) );
  INV_X1 U22417 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19469) );
  AOI22_X1 U22418 ( .A1(n19477), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n19476), 
        .B2(P2_LWORD_REG_4__SCAN_IN), .ZN(n19468) );
  OAI21_X1 U22419 ( .B1(n19469), .B2(n19479), .A(n19468), .ZN(P2_U2947) );
  INV_X1 U22420 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19471) );
  AOI22_X1 U22421 ( .A1(n19477), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n19476), 
        .B2(P2_LWORD_REG_3__SCAN_IN), .ZN(n19470) );
  OAI21_X1 U22422 ( .B1(n19471), .B2(n19479), .A(n19470), .ZN(P2_U2948) );
  AOI22_X1 U22423 ( .A1(n19477), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n19476), 
        .B2(P2_LWORD_REG_2__SCAN_IN), .ZN(n19472) );
  OAI21_X1 U22424 ( .B1(n19473), .B2(n19479), .A(n19472), .ZN(P2_U2949) );
  INV_X1 U22425 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19475) );
  AOI22_X1 U22426 ( .A1(n19477), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n19476), 
        .B2(P2_LWORD_REG_1__SCAN_IN), .ZN(n19474) );
  OAI21_X1 U22427 ( .B1(n19475), .B2(n19479), .A(n19474), .ZN(P2_U2950) );
  INV_X1 U22428 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19480) );
  AOI22_X1 U22429 ( .A1(n19477), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(n19476), 
        .B2(P2_LWORD_REG_0__SCAN_IN), .ZN(n19478) );
  OAI21_X1 U22430 ( .B1(n19480), .B2(n19479), .A(n19478), .ZN(P2_U2951) );
  AOI22_X1 U22431 ( .A1(n19518), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n19517), .ZN(n19481) );
  OAI21_X1 U22432 ( .B1(n19497), .B2(n19520), .A(n19481), .ZN(P2_U2953) );
  AOI22_X1 U22433 ( .A1(n19518), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n19517), .ZN(n19482) );
  OAI21_X1 U22434 ( .B1(n19499), .B2(n19520), .A(n19482), .ZN(P2_U2954) );
  AOI22_X1 U22435 ( .A1(n19518), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_19__SCAN_IN), .B2(n19517), .ZN(n19483) );
  OAI21_X1 U22436 ( .B1(n19547), .B2(n19520), .A(n19483), .ZN(P2_U2955) );
  AOI22_X1 U22437 ( .A1(n19518), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n19517), .ZN(n19484) );
  OAI21_X1 U22438 ( .B1(n19502), .B2(n19520), .A(n19484), .ZN(P2_U2956) );
  AOI22_X1 U22439 ( .A1(n19518), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_21__SCAN_IN), .B2(n19517), .ZN(n19485) );
  OAI21_X1 U22440 ( .B1(n19504), .B2(n19520), .A(n19485), .ZN(P2_U2957) );
  AOI22_X1 U22441 ( .A1(n19518), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n19517), .ZN(n19486) );
  OAI21_X1 U22442 ( .B1(n19506), .B2(n19520), .A(n19486), .ZN(P2_U2958) );
  AOI22_X1 U22443 ( .A1(n19518), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_23__SCAN_IN), .B2(n19517), .ZN(n19487) );
  OAI21_X1 U22444 ( .B1(n19508), .B2(n19520), .A(n19487), .ZN(P2_U2959) );
  AOI22_X1 U22445 ( .A1(n19518), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n19517), .ZN(n19490) );
  NAND2_X1 U22446 ( .A1(n19489), .A2(n19488), .ZN(n19509) );
  NAND2_X1 U22447 ( .A1(n19490), .A2(n19509), .ZN(P2_U2960) );
  AOI22_X1 U22448 ( .A1(n19518), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n19517), .ZN(n19491) );
  OAI21_X1 U22449 ( .B1(n19512), .B2(n19520), .A(n19491), .ZN(P2_U2963) );
  AOI22_X1 U22450 ( .A1(n19518), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n19517), .ZN(n19492) );
  OAI21_X1 U22451 ( .B1(n19514), .B2(n19520), .A(n19492), .ZN(P2_U2964) );
  AOI22_X1 U22452 ( .A1(n19518), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19517), .ZN(n19493) );
  OAI21_X1 U22453 ( .B1(n19516), .B2(n19520), .A(n19493), .ZN(P2_U2965) );
  AOI22_X1 U22454 ( .A1(n19518), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n19517), .ZN(n19494) );
  OAI21_X1 U22455 ( .B1(n19495), .B2(n19520), .A(n19494), .ZN(P2_U2967) );
  AOI22_X1 U22456 ( .A1(n19518), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_1__SCAN_IN), .B2(n19517), .ZN(n19496) );
  OAI21_X1 U22457 ( .B1(n19497), .B2(n19520), .A(n19496), .ZN(P2_U2968) );
  AOI22_X1 U22458 ( .A1(n19518), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n19517), .ZN(n19498) );
  OAI21_X1 U22459 ( .B1(n19499), .B2(n19520), .A(n19498), .ZN(P2_U2969) );
  AOI22_X1 U22460 ( .A1(n19518), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n19517), .ZN(n19500) );
  OAI21_X1 U22461 ( .B1(n19547), .B2(n19520), .A(n19500), .ZN(P2_U2970) );
  AOI22_X1 U22462 ( .A1(n19518), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n19517), .ZN(n19501) );
  OAI21_X1 U22463 ( .B1(n19502), .B2(n19520), .A(n19501), .ZN(P2_U2971) );
  AOI22_X1 U22464 ( .A1(n19518), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n19517), .ZN(n19503) );
  OAI21_X1 U22465 ( .B1(n19504), .B2(n19520), .A(n19503), .ZN(P2_U2972) );
  AOI22_X1 U22466 ( .A1(n19518), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_6__SCAN_IN), .B2(n19517), .ZN(n19505) );
  OAI21_X1 U22467 ( .B1(n19506), .B2(n19520), .A(n19505), .ZN(P2_U2973) );
  AOI22_X1 U22468 ( .A1(n19518), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_7__SCAN_IN), .B2(n19517), .ZN(n19507) );
  OAI21_X1 U22469 ( .B1(n19508), .B2(n19520), .A(n19507), .ZN(P2_U2974) );
  AOI22_X1 U22470 ( .A1(n19518), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_8__SCAN_IN), .B2(n19517), .ZN(n19510) );
  NAND2_X1 U22471 ( .A1(n19510), .A2(n19509), .ZN(P2_U2975) );
  AOI22_X1 U22472 ( .A1(n19518), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n19517), .ZN(n19511) );
  OAI21_X1 U22473 ( .B1(n19512), .B2(n19520), .A(n19511), .ZN(P2_U2978) );
  AOI22_X1 U22474 ( .A1(n19518), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n19517), .ZN(n19513) );
  OAI21_X1 U22475 ( .B1(n19514), .B2(n19520), .A(n19513), .ZN(P2_U2979) );
  AOI22_X1 U22476 ( .A1(n19518), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n19517), .ZN(n19515) );
  OAI21_X1 U22477 ( .B1(n19516), .B2(n19520), .A(n19515), .ZN(P2_U2980) );
  AOI22_X1 U22478 ( .A1(n19518), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(
        P2_EAX_REG_15__SCAN_IN), .B2(n19517), .ZN(n19519) );
  OAI21_X1 U22479 ( .B1(n19521), .B2(n19520), .A(n19519), .ZN(P2_U2982) );
  INV_X1 U22480 ( .A(n20098), .ZN(n20030) );
  NAND2_X1 U22481 ( .A1(n20262), .A2(n20271), .ZN(n19626) );
  OR2_X1 U22482 ( .A1(n19626), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19593) );
  NOR2_X1 U22483 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19593), .ZN(
        n19529) );
  INV_X1 U22484 ( .A(n19529), .ZN(n19579) );
  OAI22_X1 U22485 ( .A1(n20152), .A2(n20051), .B1(n20094), .B2(n19579), .ZN(
        n19524) );
  INV_X1 U22486 ( .A(n19524), .ZN(n19534) );
  AOI21_X1 U22487 ( .B1(n20152), .B2(n19625), .A(n20036), .ZN(n19525) );
  NOR2_X1 U22488 ( .A1(n19525), .A2(n20037), .ZN(n19528) );
  OAI21_X1 U22489 ( .B1(n19530), .B2(n20258), .A(n20104), .ZN(n19526) );
  AOI21_X1 U22490 ( .B1(n19528), .B2(n20155), .A(n19526), .ZN(n19527) );
  OAI21_X1 U22491 ( .B1(n19527), .B2(n19529), .A(n20102), .ZN(n19583) );
  OAI21_X1 U22492 ( .B1(n20105), .B2(n19529), .A(n19528), .ZN(n19532) );
  OAI21_X1 U22493 ( .B1(n19530), .B2(n19529), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19531) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19583), .B1(
        n20048), .B2(n19582), .ZN(n19533) );
  OAI211_X1 U22495 ( .C1(n20109), .C2(n19625), .A(n19534), .B(n19533), .ZN(
        P2_U3048) );
  AOI22_X1 U22496 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19576), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19575), .ZN(n20116) );
  OAI22_X1 U22497 ( .A1(n20152), .A2(n20116), .B1(n19579), .B2(n20110), .ZN(
        n19537) );
  INV_X1 U22498 ( .A(n19537), .ZN(n19540) );
  AOI22_X1 U22499 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19583), .B1(
        n20053), .B2(n19582), .ZN(n19539) );
  OAI211_X1 U22500 ( .C1(n20006), .C2(n19625), .A(n19540), .B(n19539), .ZN(
        P2_U3049) );
  AOI22_X1 U22501 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19576), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19575), .ZN(n20123) );
  AOI22_X1 U22502 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19576), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19575), .ZN(n20060) );
  OAI22_X1 U22503 ( .A1(n20152), .A2(n20060), .B1(n19579), .B2(n20117), .ZN(
        n19541) );
  INV_X1 U22504 ( .A(n19541), .ZN(n19544) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19583), .B1(
        n20057), .B2(n19582), .ZN(n19543) );
  OAI211_X1 U22506 ( .C1(n20123), .C2(n19625), .A(n19544), .B(n19543), .ZN(
        P2_U3050) );
  AOI22_X2 U22507 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19576), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19575), .ZN(n20130) );
  AOI22_X1 U22508 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19576), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19575), .ZN(n20066) );
  NAND2_X1 U22509 ( .A1(n19578), .A2(n19545), .ZN(n20124) );
  OAI22_X1 U22510 ( .A1(n20152), .A2(n20066), .B1(n19579), .B2(n20124), .ZN(
        n19546) );
  INV_X1 U22511 ( .A(n19546), .ZN(n19550) );
  INV_X1 U22512 ( .A(n19547), .ZN(n19548) );
  AOI22_X1 U22513 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19583), .B1(
        n20063), .B2(n19582), .ZN(n19549) );
  OAI211_X1 U22514 ( .C1(n20130), .C2(n19625), .A(n19550), .B(n19549), .ZN(
        P2_U3051) );
  AOI22_X1 U22515 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19575), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19576), .ZN(n20067) );
  OAI22_X1 U22516 ( .A1(n20152), .A2(n20067), .B1(n20131), .B2(n19579), .ZN(
        n19554) );
  INV_X1 U22517 ( .A(n19554), .ZN(n19557) );
  AOI22_X1 U22518 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19583), .B1(
        n20069), .B2(n19582), .ZN(n19556) );
  OAI211_X1 U22519 ( .C1(n20137), .C2(n19625), .A(n19557), .B(n19556), .ZN(
        P2_U3052) );
  AOI22_X1 U22520 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19575), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19576), .ZN(n20077) );
  OAI22_X1 U22521 ( .A1(n20152), .A2(n20077), .B1(n19579), .B2(n20138), .ZN(
        n19560) );
  INV_X1 U22522 ( .A(n19560), .ZN(n19563) );
  AOI22_X1 U22523 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19583), .B1(
        n20074), .B2(n19582), .ZN(n19562) );
  OAI211_X1 U22524 ( .C1(n20144), .C2(n19625), .A(n19563), .B(n19562), .ZN(
        P2_U3053) );
  AOI22_X1 U22525 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19576), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19575), .ZN(n20079) );
  AND2_X1 U22526 ( .A1(n19578), .A2(n19566), .ZN(n19976) );
  OAI22_X1 U22527 ( .A1(n20152), .A2(n20079), .B1(n20145), .B2(n19579), .ZN(
        n19567) );
  INV_X1 U22528 ( .A(n19567), .ZN(n19570) );
  AOI22_X1 U22529 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19583), .B1(
        n20081), .B2(n19582), .ZN(n19569) );
  OAI211_X1 U22530 ( .C1(n20153), .C2(n19625), .A(n19570), .B(n19569), .ZN(
        P2_U3054) );
  AOI22_X1 U22531 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19576), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19575), .ZN(n20164) );
  OAI22_X1 U22532 ( .A1(n20152), .A2(n20164), .B1(n19579), .B2(n20154), .ZN(
        n19580) );
  INV_X1 U22533 ( .A(n19580), .ZN(n19585) );
  AOI22_X1 U22534 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19583), .B1(
        n20087), .B2(n19582), .ZN(n19584) );
  OAI211_X1 U22535 ( .C1(n20029), .C2(n19625), .A(n19585), .B(n19584), .ZN(
        P2_U3055) );
  OR2_X1 U22536 ( .A1(n19855), .A2(n19626), .ZN(n19619) );
  NAND2_X1 U22537 ( .A1(n19619), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19586) );
  NOR2_X1 U22538 ( .A1(n19587), .A2(n19586), .ZN(n19592) );
  INV_X1 U22539 ( .A(n19593), .ZN(n19588) );
  OAI21_X1 U22540 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19588), .A(n19785), 
        .ZN(n19589) );
  INV_X1 U22541 ( .A(n20048), .ZN(n20095) );
  OAI22_X1 U22542 ( .A1(n19620), .A2(n20095), .B1(n20094), .B2(n19619), .ZN(
        n19590) );
  INV_X1 U22543 ( .A(n19590), .ZN(n19600) );
  INV_X1 U22544 ( .A(n19619), .ZN(n19596) );
  NAND2_X1 U22545 ( .A1(n19598), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19788) );
  INV_X1 U22546 ( .A(n19788), .ZN(n19591) );
  NAND2_X1 U22547 ( .A1(n19591), .A2(n19820), .ZN(n19594) );
  AOI21_X1 U22548 ( .B1(n19594), .B2(n19593), .A(n19592), .ZN(n19595) );
  OAI211_X1 U22549 ( .C1(n19596), .C2(n20104), .A(n19595), .B(n20102), .ZN(
        n19622) );
  NAND2_X1 U22550 ( .A1(n19820), .A2(n19792), .ZN(n19631) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19622), .B1(
        n19652), .B2(n19928), .ZN(n19599) );
  OAI211_X1 U22552 ( .C1(n20051), .C2(n19625), .A(n19600), .B(n19599), .ZN(
        P2_U3056) );
  INV_X1 U22553 ( .A(n20053), .ZN(n20111) );
  OAI22_X1 U22554 ( .A1(n19620), .A2(n20111), .B1(n20110), .B2(n19619), .ZN(
        n19601) );
  INV_X1 U22555 ( .A(n19601), .ZN(n19603) );
  AOI22_X1 U22556 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19622), .B1(
        n19652), .B2(n20113), .ZN(n19602) );
  OAI211_X1 U22557 ( .C1(n20116), .C2(n19625), .A(n19603), .B(n19602), .ZN(
        P2_U3057) );
  INV_X1 U22558 ( .A(n20057), .ZN(n20118) );
  OAI22_X1 U22559 ( .A1(n19620), .A2(n20118), .B1(n20117), .B2(n19619), .ZN(
        n19604) );
  INV_X1 U22560 ( .A(n19604), .ZN(n19606) );
  INV_X1 U22561 ( .A(n20123), .ZN(n19959) );
  AOI22_X1 U22562 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19622), .B1(
        n19652), .B2(n19959), .ZN(n19605) );
  OAI211_X1 U22563 ( .C1(n20060), .C2(n19625), .A(n19606), .B(n19605), .ZN(
        P2_U3058) );
  INV_X1 U22564 ( .A(n20063), .ZN(n20125) );
  OAI22_X1 U22565 ( .A1(n19620), .A2(n20125), .B1(n20124), .B2(n19619), .ZN(
        n19607) );
  INV_X1 U22566 ( .A(n19607), .ZN(n19609) );
  INV_X1 U22567 ( .A(n20130), .ZN(n19964) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19622), .B1(
        n19652), .B2(n19964), .ZN(n19608) );
  OAI211_X1 U22569 ( .C1(n20066), .C2(n19625), .A(n19609), .B(n19608), .ZN(
        P2_U3059) );
  INV_X1 U22570 ( .A(n20069), .ZN(n20132) );
  OAI22_X1 U22571 ( .A1(n19620), .A2(n20132), .B1(n20131), .B2(n19619), .ZN(
        n19610) );
  INV_X1 U22572 ( .A(n19610), .ZN(n19612) );
  AOI22_X1 U22573 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19622), .B1(
        n19652), .B2(n19969), .ZN(n19611) );
  OAI211_X1 U22574 ( .C1(n20067), .C2(n19625), .A(n19612), .B(n19611), .ZN(
        P2_U3060) );
  INV_X1 U22575 ( .A(n20074), .ZN(n20139) );
  OAI22_X1 U22576 ( .A1(n19620), .A2(n20139), .B1(n20138), .B2(n19619), .ZN(
        n19613) );
  INV_X1 U22577 ( .A(n19613), .ZN(n19615) );
  AOI22_X1 U22578 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19622), .B1(
        n19652), .B2(n20073), .ZN(n19614) );
  OAI211_X1 U22579 ( .C1(n20077), .C2(n19625), .A(n19615), .B(n19614), .ZN(
        P2_U3061) );
  INV_X1 U22580 ( .A(n20081), .ZN(n20146) );
  OAI22_X1 U22581 ( .A1(n19620), .A2(n20146), .B1(n20145), .B2(n19619), .ZN(
        n19616) );
  INV_X1 U22582 ( .A(n19616), .ZN(n19618) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19622), .B1(
        n19652), .B2(n19977), .ZN(n19617) );
  OAI211_X1 U22584 ( .C1(n20079), .C2(n19625), .A(n19618), .B(n19617), .ZN(
        P2_U3062) );
  INV_X1 U22585 ( .A(n20087), .ZN(n20156) );
  OAI22_X1 U22586 ( .A1(n19620), .A2(n20156), .B1(n20154), .B2(n19619), .ZN(
        n19621) );
  INV_X1 U22587 ( .A(n19621), .ZN(n19624) );
  AOI22_X1 U22588 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19622), .B1(
        n19652), .B2(n20159), .ZN(n19623) );
  OAI211_X1 U22589 ( .C1(n20164), .C2(n19625), .A(n19624), .B(n19623), .ZN(
        P2_U3063) );
  INV_X1 U22590 ( .A(n19626), .ZN(n19628) );
  AND2_X1 U22591 ( .A1(n19660), .A2(n20034), .ZN(n19650) );
  OAI21_X1 U22592 ( .B1(n19627), .B2(n19650), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19629) );
  NAND2_X1 U22593 ( .A1(n19889), .A2(n19628), .ZN(n19632) );
  NAND2_X1 U22594 ( .A1(n19629), .A2(n19632), .ZN(n19651) );
  AOI22_X1 U22595 ( .A1(n19651), .A2(n20048), .B1(n19894), .B2(n19650), .ZN(
        n19637) );
  AOI21_X1 U22596 ( .B1(n19630), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19635) );
  AND2_X1 U22597 ( .A1(n19683), .A2(n19631), .ZN(n19633) );
  OAI211_X1 U22598 ( .C1(n19633), .C2(n20036), .A(n20258), .B(n19632), .ZN(
        n19634) );
  OAI211_X1 U22599 ( .C1(n19650), .C2(n19635), .A(n19634), .B(n20102), .ZN(
        n19653) );
  AOI22_X1 U22600 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19653), .B1(
        n19652), .B2(n20106), .ZN(n19636) );
  OAI211_X1 U22601 ( .C1(n20109), .C2(n19683), .A(n19637), .B(n19636), .ZN(
        P2_U3064) );
  AOI22_X1 U22602 ( .A1(n19651), .A2(n20053), .B1(n19650), .B2(n20052), .ZN(
        n19639) );
  INV_X1 U22603 ( .A(n20116), .ZN(n20003) );
  AOI22_X1 U22604 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19653), .B1(
        n19652), .B2(n20003), .ZN(n19638) );
  OAI211_X1 U22605 ( .C1(n20006), .C2(n19683), .A(n19639), .B(n19638), .ZN(
        P2_U3065) );
  AOI22_X1 U22606 ( .A1(n19651), .A2(n20057), .B1(n19650), .B2(n19958), .ZN(
        n19641) );
  INV_X1 U22607 ( .A(n20060), .ZN(n20120) );
  AOI22_X1 U22608 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19653), .B1(
        n19652), .B2(n20120), .ZN(n19640) );
  OAI211_X1 U22609 ( .C1(n20123), .C2(n19683), .A(n19641), .B(n19640), .ZN(
        P2_U3066) );
  AOI22_X1 U22610 ( .A1(n19651), .A2(n20063), .B1(n19650), .B2(n19963), .ZN(
        n19643) );
  INV_X1 U22611 ( .A(n20066), .ZN(n20127) );
  AOI22_X1 U22612 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19653), .B1(
        n19652), .B2(n20127), .ZN(n19642) );
  OAI211_X1 U22613 ( .C1(n20130), .C2(n19683), .A(n19643), .B(n19642), .ZN(
        P2_U3067) );
  AOI22_X1 U22614 ( .A1(n19651), .A2(n20069), .B1(n19650), .B2(n19968), .ZN(
        n19645) );
  INV_X1 U22615 ( .A(n20067), .ZN(n20134) );
  AOI22_X1 U22616 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19653), .B1(
        n19652), .B2(n20134), .ZN(n19644) );
  OAI211_X1 U22617 ( .C1(n20137), .C2(n19683), .A(n19645), .B(n19644), .ZN(
        P2_U3068) );
  AOI22_X1 U22618 ( .A1(n19651), .A2(n20074), .B1(n19650), .B2(n20072), .ZN(
        n19647) );
  INV_X1 U22619 ( .A(n20077), .ZN(n20141) );
  AOI22_X1 U22620 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19653), .B1(
        n19652), .B2(n20141), .ZN(n19646) );
  OAI211_X1 U22621 ( .C1(n20144), .C2(n19683), .A(n19647), .B(n19646), .ZN(
        P2_U3069) );
  AOI22_X1 U22622 ( .A1(n19651), .A2(n20081), .B1(n19650), .B2(n19976), .ZN(
        n19649) );
  INV_X1 U22623 ( .A(n20079), .ZN(n20148) );
  AOI22_X1 U22624 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19653), .B1(
        n19652), .B2(n20148), .ZN(n19648) );
  OAI211_X1 U22625 ( .C1(n20153), .C2(n19683), .A(n19649), .B(n19648), .ZN(
        P2_U3070) );
  AOI22_X1 U22626 ( .A1(n19651), .A2(n20087), .B1(n19650), .B2(n20084), .ZN(
        n19655) );
  INV_X1 U22627 ( .A(n20164), .ZN(n20024) );
  AOI22_X1 U22628 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19653), .B1(
        n19652), .B2(n20024), .ZN(n19654) );
  OAI211_X1 U22629 ( .C1(n20029), .C2(n19683), .A(n19655), .B(n19654), .ZN(
        P2_U3071) );
  INV_X1 U22630 ( .A(n19719), .ZN(n19689) );
  AND2_X1 U22631 ( .A1(n19660), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19679) );
  INV_X1 U22632 ( .A(n19679), .ZN(n19682) );
  OAI22_X1 U22633 ( .A1(n19683), .A2(n20051), .B1(n20094), .B2(n19682), .ZN(
        n19656) );
  INV_X1 U22634 ( .A(n19656), .ZN(n19666) );
  OAI21_X1 U22635 ( .B1(n19788), .B2(n19657), .A(n20258), .ZN(n19664) );
  INV_X1 U22636 ( .A(n19661), .ZN(n19658) );
  OAI211_X1 U22637 ( .C1(n19658), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20037), 
        .B(n19682), .ZN(n19659) );
  OAI211_X1 U22638 ( .C1(n19664), .C2(n19660), .A(n20102), .B(n19659), .ZN(
        n19686) );
  INV_X1 U22639 ( .A(n19660), .ZN(n19663) );
  OAI21_X1 U22640 ( .B1(n19661), .B2(n19679), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19662) );
  AOI22_X1 U22641 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19686), .B1(
        n20048), .B2(n19685), .ZN(n19665) );
  OAI211_X1 U22642 ( .C1(n20109), .C2(n19689), .A(n19666), .B(n19665), .ZN(
        P2_U3072) );
  OAI22_X1 U22643 ( .A1(n19683), .A2(n20116), .B1(n19682), .B2(n20110), .ZN(
        n19667) );
  INV_X1 U22644 ( .A(n19667), .ZN(n19669) );
  AOI22_X1 U22645 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19686), .B1(
        n20053), .B2(n19685), .ZN(n19668) );
  OAI211_X1 U22646 ( .C1(n20006), .C2(n19689), .A(n19669), .B(n19668), .ZN(
        P2_U3073) );
  AOI22_X1 U22647 ( .A1(n19719), .A2(n19959), .B1(n19679), .B2(n19958), .ZN(
        n19671) );
  AOI22_X1 U22648 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19686), .B1(
        n20057), .B2(n19685), .ZN(n19670) );
  OAI211_X1 U22649 ( .C1(n20060), .C2(n19683), .A(n19671), .B(n19670), .ZN(
        P2_U3074) );
  AOI22_X1 U22650 ( .A1(n19719), .A2(n19964), .B1(n19679), .B2(n19963), .ZN(
        n19673) );
  AOI22_X1 U22651 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19686), .B1(
        n20063), .B2(n19685), .ZN(n19672) );
  OAI211_X1 U22652 ( .C1(n20066), .C2(n19683), .A(n19673), .B(n19672), .ZN(
        P2_U3075) );
  AOI22_X1 U22653 ( .A1(n19969), .A2(n19719), .B1(n19679), .B2(n19968), .ZN(
        n19675) );
  AOI22_X1 U22654 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19686), .B1(
        n20069), .B2(n19685), .ZN(n19674) );
  OAI211_X1 U22655 ( .C1(n20067), .C2(n19683), .A(n19675), .B(n19674), .ZN(
        P2_U3076) );
  OAI22_X1 U22656 ( .A1(n19683), .A2(n20077), .B1(n19682), .B2(n20138), .ZN(
        n19676) );
  INV_X1 U22657 ( .A(n19676), .ZN(n19678) );
  AOI22_X1 U22658 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19686), .B1(
        n20074), .B2(n19685), .ZN(n19677) );
  OAI211_X1 U22659 ( .C1(n20144), .C2(n19689), .A(n19678), .B(n19677), .ZN(
        P2_U3077) );
  AOI22_X1 U22660 ( .A1(n19977), .A2(n19719), .B1(n19679), .B2(n19976), .ZN(
        n19681) );
  AOI22_X1 U22661 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19686), .B1(
        n20081), .B2(n19685), .ZN(n19680) );
  OAI211_X1 U22662 ( .C1(n20079), .C2(n19683), .A(n19681), .B(n19680), .ZN(
        P2_U3078) );
  OAI22_X1 U22663 ( .A1(n19683), .A2(n20164), .B1(n19682), .B2(n20154), .ZN(
        n19684) );
  INV_X1 U22664 ( .A(n19684), .ZN(n19688) );
  AOI22_X1 U22665 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19686), .B1(
        n20087), .B2(n19685), .ZN(n19687) );
  OAI211_X1 U22666 ( .C1(n20029), .C2(n19689), .A(n19688), .B(n19687), .ZN(
        P2_U3079) );
  INV_X1 U22667 ( .A(n19690), .ZN(n19691) );
  NAND2_X1 U22668 ( .A1(n19691), .A2(n20262), .ZN(n19699) );
  NOR2_X1 U22669 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19692) );
  AND2_X1 U22670 ( .A1(n19726), .A2(n20034), .ZN(n19717) );
  OAI21_X1 U22671 ( .B1(n19693), .B2(n19717), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19694) );
  AOI22_X1 U22672 ( .A1(n19718), .A2(n20048), .B1(n19894), .B2(n19717), .ZN(
        n19704) );
  AOI21_X1 U22673 ( .B1(n19696), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19702) );
  INV_X1 U22674 ( .A(n19697), .ZN(n19700) );
  OAI21_X1 U22675 ( .B1(n19719), .B2(n19747), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19698) );
  OAI21_X1 U22676 ( .B1(n19700), .B2(n19699), .A(n19698), .ZN(n19701) );
  OAI211_X1 U22677 ( .C1(n19702), .C2(n19717), .A(n20102), .B(n19701), .ZN(
        n19720) );
  AOI22_X1 U22678 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19720), .B1(
        n19719), .B2(n20106), .ZN(n19703) );
  OAI211_X1 U22679 ( .C1(n20109), .C2(n19745), .A(n19704), .B(n19703), .ZN(
        P2_U3080) );
  AOI22_X1 U22680 ( .A1(n19718), .A2(n20053), .B1(n20052), .B2(n19717), .ZN(
        n19706) );
  AOI22_X1 U22681 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19720), .B1(
        n19719), .B2(n20003), .ZN(n19705) );
  OAI211_X1 U22682 ( .C1(n20006), .C2(n19745), .A(n19706), .B(n19705), .ZN(
        P2_U3081) );
  AOI22_X1 U22683 ( .A1(n19718), .A2(n20057), .B1(n19958), .B2(n19717), .ZN(
        n19708) );
  AOI22_X1 U22684 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19720), .B1(
        n19719), .B2(n20120), .ZN(n19707) );
  OAI211_X1 U22685 ( .C1(n20123), .C2(n19745), .A(n19708), .B(n19707), .ZN(
        P2_U3082) );
  AOI22_X1 U22686 ( .A1(n19718), .A2(n20063), .B1(n19963), .B2(n19717), .ZN(
        n19710) );
  AOI22_X1 U22687 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19720), .B1(
        n19719), .B2(n20127), .ZN(n19709) );
  OAI211_X1 U22688 ( .C1(n20130), .C2(n19745), .A(n19710), .B(n19709), .ZN(
        P2_U3083) );
  AOI22_X1 U22689 ( .A1(n19718), .A2(n20069), .B1(n19968), .B2(n19717), .ZN(
        n19712) );
  AOI22_X1 U22690 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19720), .B1(
        n19719), .B2(n20134), .ZN(n19711) );
  OAI211_X1 U22691 ( .C1(n20137), .C2(n19745), .A(n19712), .B(n19711), .ZN(
        P2_U3084) );
  AOI22_X1 U22692 ( .A1(n19718), .A2(n20074), .B1(n20072), .B2(n19717), .ZN(
        n19714) );
  AOI22_X1 U22693 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19720), .B1(
        n19719), .B2(n20141), .ZN(n19713) );
  OAI211_X1 U22694 ( .C1(n20144), .C2(n19745), .A(n19714), .B(n19713), .ZN(
        P2_U3085) );
  AOI22_X1 U22695 ( .A1(n19718), .A2(n20081), .B1(n19976), .B2(n19717), .ZN(
        n19716) );
  AOI22_X1 U22696 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19720), .B1(
        n19719), .B2(n20148), .ZN(n19715) );
  OAI211_X1 U22697 ( .C1(n20153), .C2(n19745), .A(n19716), .B(n19715), .ZN(
        P2_U3086) );
  AOI22_X1 U22698 ( .A1(n19718), .A2(n20087), .B1(n20084), .B2(n19717), .ZN(
        n19722) );
  AOI22_X1 U22699 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19720), .B1(
        n19719), .B2(n20024), .ZN(n19721) );
  OAI211_X1 U22700 ( .C1(n20029), .C2(n19745), .A(n19722), .B(n19721), .ZN(
        P2_U3087) );
  INV_X1 U22701 ( .A(n19780), .ZN(n19752) );
  AOI22_X1 U22702 ( .A1(n19747), .A2(n20106), .B1(n19894), .B2(n19746), .ZN(
        n19732) );
  OAI21_X1 U22703 ( .B1(n19788), .B2(n19993), .A(n20258), .ZN(n19730) );
  OAI21_X1 U22704 ( .B1(n19727), .B2(n20044), .A(n20104), .ZN(n19724) );
  INV_X1 U22705 ( .A(n19746), .ZN(n19761) );
  AOI21_X1 U22706 ( .B1(n19724), .B2(n19761), .A(n19996), .ZN(n19725) );
  INV_X1 U22707 ( .A(n19726), .ZN(n19729) );
  OAI21_X1 U22708 ( .B1(n19727), .B2(n19746), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19728) );
  AOI22_X1 U22709 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19749), .B1(
        n20048), .B2(n19748), .ZN(n19731) );
  OAI211_X1 U22710 ( .C1(n20109), .C2(n19752), .A(n19732), .B(n19731), .ZN(
        P2_U3088) );
  AOI22_X1 U22711 ( .A1(n19747), .A2(n20003), .B1(n19746), .B2(n20052), .ZN(
        n19734) );
  AOI22_X1 U22712 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19749), .B1(
        n20053), .B2(n19748), .ZN(n19733) );
  OAI211_X1 U22713 ( .C1(n20006), .C2(n19752), .A(n19734), .B(n19733), .ZN(
        P2_U3089) );
  AOI22_X1 U22714 ( .A1(n19780), .A2(n19959), .B1(n19746), .B2(n19958), .ZN(
        n19736) );
  AOI22_X1 U22715 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19749), .B1(
        n20057), .B2(n19748), .ZN(n19735) );
  OAI211_X1 U22716 ( .C1(n20060), .C2(n19745), .A(n19736), .B(n19735), .ZN(
        P2_U3090) );
  AOI22_X1 U22717 ( .A1(n19747), .A2(n20127), .B1(n19746), .B2(n19963), .ZN(
        n19738) );
  AOI22_X1 U22718 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19749), .B1(
        n20063), .B2(n19748), .ZN(n19737) );
  OAI211_X1 U22719 ( .C1(n20130), .C2(n19752), .A(n19738), .B(n19737), .ZN(
        P2_U3091) );
  AOI22_X1 U22720 ( .A1(n19969), .A2(n19780), .B1(n19746), .B2(n19968), .ZN(
        n19740) );
  AOI22_X1 U22721 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19749), .B1(
        n20069), .B2(n19748), .ZN(n19739) );
  OAI211_X1 U22722 ( .C1(n20067), .C2(n19745), .A(n19740), .B(n19739), .ZN(
        P2_U3092) );
  AOI22_X1 U22723 ( .A1(n19747), .A2(n20141), .B1(n19746), .B2(n20072), .ZN(
        n19742) );
  AOI22_X1 U22724 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19749), .B1(
        n20074), .B2(n19748), .ZN(n19741) );
  OAI211_X1 U22725 ( .C1(n20144), .C2(n19752), .A(n19742), .B(n19741), .ZN(
        P2_U3093) );
  AOI22_X1 U22726 ( .A1(n19977), .A2(n19780), .B1(n19746), .B2(n19976), .ZN(
        n19744) );
  AOI22_X1 U22727 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19749), .B1(
        n20081), .B2(n19748), .ZN(n19743) );
  OAI211_X1 U22728 ( .C1(n20079), .C2(n19745), .A(n19744), .B(n19743), .ZN(
        P2_U3094) );
  AOI22_X1 U22729 ( .A1(n19747), .A2(n20024), .B1(n19746), .B2(n20084), .ZN(
        n19751) );
  AOI22_X1 U22730 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19749), .B1(
        n20087), .B2(n19748), .ZN(n19750) );
  OAI211_X1 U22731 ( .C1(n20029), .C2(n19752), .A(n19751), .B(n19750), .ZN(
        P2_U3095) );
  AND2_X1 U22732 ( .A1(n19754), .A2(n20262), .ZN(n19791) );
  NAND2_X1 U22733 ( .A1(n19791), .A2(n20034), .ZN(n19757) );
  NOR2_X1 U22734 ( .A1(n20258), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19756) );
  OAI222_X1 U22735 ( .A1(n19761), .A2(n20037), .B1(n19757), .B2(n19756), .C1(
        n20044), .C2(n19755), .ZN(n19779) );
  INV_X1 U22736 ( .A(n19757), .ZN(n19778) );
  AOI22_X1 U22737 ( .A1(n19779), .A2(n20048), .B1(n19894), .B2(n19778), .ZN(
        n19765) );
  INV_X1 U22738 ( .A(n19819), .ZN(n19758) );
  OAI21_X1 U22739 ( .B1(n19780), .B2(n19758), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19762) );
  NOR2_X1 U22740 ( .A1(n19759), .A2(n20258), .ZN(n19760) );
  AOI211_X1 U22741 ( .C1(n19762), .C2(n19761), .A(P2_STATE2_REG_3__SCAN_IN), 
        .B(n19760), .ZN(n19763) );
  OAI21_X1 U22742 ( .B1(n19763), .B2(n19778), .A(n20102), .ZN(n19781) );
  AOI22_X1 U22743 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19781), .B1(
        n19780), .B2(n20106), .ZN(n19764) );
  OAI211_X1 U22744 ( .C1(n20109), .C2(n19819), .A(n19765), .B(n19764), .ZN(
        P2_U3096) );
  AOI22_X1 U22745 ( .A1(n19779), .A2(n20053), .B1(n20052), .B2(n19778), .ZN(
        n19767) );
  AOI22_X1 U22746 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19781), .B1(
        n19780), .B2(n20003), .ZN(n19766) );
  OAI211_X1 U22747 ( .C1(n20006), .C2(n19819), .A(n19767), .B(n19766), .ZN(
        P2_U3097) );
  AOI22_X1 U22748 ( .A1(n19779), .A2(n20057), .B1(n19958), .B2(n19778), .ZN(
        n19769) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19781), .B1(
        n19780), .B2(n20120), .ZN(n19768) );
  OAI211_X1 U22750 ( .C1(n20123), .C2(n19819), .A(n19769), .B(n19768), .ZN(
        P2_U3098) );
  AOI22_X1 U22751 ( .A1(n19779), .A2(n20063), .B1(n19963), .B2(n19778), .ZN(
        n19771) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19781), .B1(
        n19780), .B2(n20127), .ZN(n19770) );
  OAI211_X1 U22753 ( .C1(n20130), .C2(n19819), .A(n19771), .B(n19770), .ZN(
        P2_U3099) );
  AOI22_X1 U22754 ( .A1(n19779), .A2(n20069), .B1(n19968), .B2(n19778), .ZN(
        n19773) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19781), .B1(
        n19780), .B2(n20134), .ZN(n19772) );
  OAI211_X1 U22756 ( .C1(n20137), .C2(n19819), .A(n19773), .B(n19772), .ZN(
        P2_U3100) );
  AOI22_X1 U22757 ( .A1(n19779), .A2(n20074), .B1(n20072), .B2(n19778), .ZN(
        n19775) );
  AOI22_X1 U22758 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19781), .B1(
        n19780), .B2(n20141), .ZN(n19774) );
  OAI211_X1 U22759 ( .C1(n20144), .C2(n19819), .A(n19775), .B(n19774), .ZN(
        P2_U3101) );
  AOI22_X1 U22760 ( .A1(n19779), .A2(n20081), .B1(n19976), .B2(n19778), .ZN(
        n19777) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19781), .B1(
        n19780), .B2(n20148), .ZN(n19776) );
  OAI211_X1 U22762 ( .C1(n20153), .C2(n19819), .A(n19777), .B(n19776), .ZN(
        P2_U3102) );
  AOI22_X1 U22763 ( .A1(n19779), .A2(n20087), .B1(n20084), .B2(n19778), .ZN(
        n19783) );
  AOI22_X1 U22764 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19781), .B1(
        n19780), .B2(n20024), .ZN(n19782) );
  OAI211_X1 U22765 ( .C1(n20029), .C2(n19819), .A(n19783), .B(n19782), .ZN(
        P2_U3103) );
  NAND2_X1 U22766 ( .A1(n19791), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19825) );
  NAND2_X1 U22767 ( .A1(n19825), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19784) );
  NOR2_X1 U22768 ( .A1(n11956), .A2(n19784), .ZN(n19789) );
  OAI21_X1 U22769 ( .B1(n19791), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n19785), 
        .ZN(n19786) );
  OAI22_X1 U22770 ( .A1(n19813), .A2(n20095), .B1(n20094), .B2(n19825), .ZN(
        n19787) );
  INV_X1 U22771 ( .A(n19787), .ZN(n19794) );
  NOR2_X1 U22772 ( .A1(n20030), .A2(n19788), .ZN(n20257) );
  AOI211_X1 U22773 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19825), .A(n19996), 
        .B(n19789), .ZN(n19790) );
  AOI22_X1 U22774 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n19928), .ZN(n19793) );
  OAI211_X1 U22775 ( .C1(n20051), .C2(n19819), .A(n19794), .B(n19793), .ZN(
        P2_U3104) );
  OAI22_X1 U22776 ( .A1(n19813), .A2(n20111), .B1(n19825), .B2(n20110), .ZN(
        n19795) );
  INV_X1 U22777 ( .A(n19795), .ZN(n19797) );
  AOI22_X1 U22778 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n20113), .ZN(n19796) );
  OAI211_X1 U22779 ( .C1(n20116), .C2(n19819), .A(n19797), .B(n19796), .ZN(
        P2_U3105) );
  OAI22_X1 U22780 ( .A1(n19813), .A2(n20118), .B1(n19825), .B2(n20117), .ZN(
        n19798) );
  INV_X1 U22781 ( .A(n19798), .ZN(n19800) );
  AOI22_X1 U22782 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n19959), .ZN(n19799) );
  OAI211_X1 U22783 ( .C1(n20060), .C2(n19819), .A(n19800), .B(n19799), .ZN(
        P2_U3106) );
  OAI22_X1 U22784 ( .A1(n19813), .A2(n20125), .B1(n19825), .B2(n20124), .ZN(
        n19801) );
  INV_X1 U22785 ( .A(n19801), .ZN(n19803) );
  AOI22_X1 U22786 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n19964), .ZN(n19802) );
  OAI211_X1 U22787 ( .C1(n20066), .C2(n19819), .A(n19803), .B(n19802), .ZN(
        P2_U3107) );
  OAI22_X1 U22788 ( .A1(n19813), .A2(n20132), .B1(n19825), .B2(n20131), .ZN(
        n19804) );
  INV_X1 U22789 ( .A(n19804), .ZN(n19806) );
  AOI22_X1 U22790 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n19969), .ZN(n19805) );
  OAI211_X1 U22791 ( .C1(n20067), .C2(n19819), .A(n19806), .B(n19805), .ZN(
        P2_U3108) );
  OAI22_X1 U22792 ( .A1(n19813), .A2(n20139), .B1(n19825), .B2(n20138), .ZN(
        n19807) );
  INV_X1 U22793 ( .A(n19807), .ZN(n19809) );
  AOI22_X1 U22794 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n20073), .ZN(n19808) );
  OAI211_X1 U22795 ( .C1(n20077), .C2(n19819), .A(n19809), .B(n19808), .ZN(
        P2_U3109) );
  OAI22_X1 U22796 ( .A1(n19813), .A2(n20146), .B1(n19825), .B2(n20145), .ZN(
        n19810) );
  INV_X1 U22797 ( .A(n19810), .ZN(n19812) );
  AOI22_X1 U22798 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n19977), .ZN(n19811) );
  OAI211_X1 U22799 ( .C1(n20079), .C2(n19819), .A(n19812), .B(n19811), .ZN(
        P2_U3110) );
  OAI22_X1 U22800 ( .A1(n19813), .A2(n20156), .B1(n19825), .B2(n20154), .ZN(
        n19814) );
  INV_X1 U22801 ( .A(n19814), .ZN(n19818) );
  AOI22_X1 U22802 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n20159), .ZN(n19817) );
  OAI211_X1 U22803 ( .C1(n20164), .C2(n19819), .A(n19818), .B(n19817), .ZN(
        P2_U3111) );
  NAND2_X1 U22804 ( .A1(n20271), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19893) );
  NOR2_X1 U22805 ( .A1(n19893), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19859) );
  INV_X1 U22806 ( .A(n19859), .ZN(n19862) );
  NOR2_X1 U22807 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19862), .ZN(
        n19848) );
  INV_X1 U22808 ( .A(n19848), .ZN(n19838) );
  OAI22_X1 U22809 ( .A1(n19854), .A2(n20051), .B1(n20094), .B2(n19838), .ZN(
        n19821) );
  INV_X1 U22810 ( .A(n19821), .ZN(n19832) );
  AOI21_X1 U22811 ( .B1(n19854), .B2(n19883), .A(n20036), .ZN(n19822) );
  NOR2_X1 U22812 ( .A1(n19822), .A2(n20037), .ZN(n19826) );
  OAI21_X1 U22813 ( .B1(n19828), .B2(n20044), .A(n20104), .ZN(n19823) );
  AOI21_X1 U22814 ( .B1(n19826), .B2(n19825), .A(n19823), .ZN(n19824) );
  OAI21_X1 U22815 ( .B1(n19824), .B2(n19848), .A(n20102), .ZN(n19851) );
  INV_X1 U22816 ( .A(n19825), .ZN(n19827) );
  OAI21_X1 U22817 ( .B1(n19848), .B2(n19827), .A(n19826), .ZN(n19830) );
  OAI21_X1 U22818 ( .B1(n19828), .B2(n19848), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19829) );
  AOI22_X1 U22819 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19851), .B1(
        n20048), .B2(n19850), .ZN(n19831) );
  OAI211_X1 U22820 ( .C1(n20109), .C2(n19883), .A(n19832), .B(n19831), .ZN(
        P2_U3112) );
  AOI22_X1 U22821 ( .A1(n20113), .A2(n19849), .B1(n20052), .B2(n19848), .ZN(
        n19834) );
  AOI22_X1 U22822 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n20053), .ZN(n19833) );
  OAI211_X1 U22823 ( .C1(n20116), .C2(n19854), .A(n19834), .B(n19833), .ZN(
        P2_U3113) );
  OAI22_X1 U22824 ( .A1(n19854), .A2(n20060), .B1(n20117), .B2(n19838), .ZN(
        n19835) );
  INV_X1 U22825 ( .A(n19835), .ZN(n19837) );
  AOI22_X1 U22826 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n20057), .ZN(n19836) );
  OAI211_X1 U22827 ( .C1(n20123), .C2(n19883), .A(n19837), .B(n19836), .ZN(
        P2_U3114) );
  OAI22_X1 U22828 ( .A1(n19883), .A2(n20130), .B1(n20124), .B2(n19838), .ZN(
        n19839) );
  INV_X1 U22829 ( .A(n19839), .ZN(n19841) );
  AOI22_X1 U22830 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n20063), .ZN(n19840) );
  OAI211_X1 U22831 ( .C1(n20066), .C2(n19854), .A(n19841), .B(n19840), .ZN(
        P2_U3115) );
  AOI22_X1 U22832 ( .A1(n19969), .A2(n19849), .B1(n19968), .B2(n19848), .ZN(
        n19843) );
  AOI22_X1 U22833 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n20069), .ZN(n19842) );
  OAI211_X1 U22834 ( .C1(n20067), .C2(n19854), .A(n19843), .B(n19842), .ZN(
        P2_U3116) );
  AOI22_X1 U22835 ( .A1(n20073), .A2(n19849), .B1(n20072), .B2(n19848), .ZN(
        n19845) );
  AOI22_X1 U22836 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n20074), .ZN(n19844) );
  OAI211_X1 U22837 ( .C1(n20077), .C2(n19854), .A(n19845), .B(n19844), .ZN(
        P2_U3117) );
  AOI22_X1 U22838 ( .A1(n19977), .A2(n19849), .B1(n19976), .B2(n19848), .ZN(
        n19847) );
  AOI22_X1 U22839 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n20081), .ZN(n19846) );
  OAI211_X1 U22840 ( .C1(n20079), .C2(n19854), .A(n19847), .B(n19846), .ZN(
        P2_U3118) );
  AOI22_X1 U22841 ( .A1(n20159), .A2(n19849), .B1(n20084), .B2(n19848), .ZN(
        n19853) );
  AOI22_X1 U22842 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n20087), .ZN(n19852) );
  OAI211_X1 U22843 ( .C1(n20164), .C2(n19854), .A(n19853), .B(n19852), .ZN(
        P2_U3119) );
  OR2_X1 U22844 ( .A1(n19855), .A2(n19893), .ZN(n19882) );
  OAI22_X1 U22845 ( .A1(n19883), .A2(n20051), .B1(n20094), .B2(n19882), .ZN(
        n19856) );
  INV_X1 U22846 ( .A(n19856), .ZN(n19865) );
  NAND2_X1 U22847 ( .A1(n10027), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19994) );
  OAI21_X1 U22848 ( .B1(n19994), .B2(n19857), .A(n20258), .ZN(n19863) );
  OAI211_X1 U22849 ( .C1(n10015), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20037), 
        .B(n19882), .ZN(n19858) );
  OAI211_X1 U22850 ( .C1(n19863), .C2(n19859), .A(n20102), .B(n19858), .ZN(
        n19886) );
  INV_X1 U22851 ( .A(n19882), .ZN(n19896) );
  OAI21_X1 U22852 ( .B1(n19860), .B2(n19896), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19861) );
  AOI22_X1 U22853 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19886), .B1(
        n20048), .B2(n19885), .ZN(n19864) );
  OAI211_X1 U22854 ( .C1(n20109), .C2(n19895), .A(n19865), .B(n19864), .ZN(
        P2_U3120) );
  OAI22_X1 U22855 ( .A1(n19883), .A2(n20116), .B1(n19882), .B2(n20110), .ZN(
        n19866) );
  INV_X1 U22856 ( .A(n19866), .ZN(n19868) );
  AOI22_X1 U22857 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19886), .B1(
        n20053), .B2(n19885), .ZN(n19867) );
  OAI211_X1 U22858 ( .C1(n20006), .C2(n19895), .A(n19868), .B(n19867), .ZN(
        P2_U3121) );
  OAI22_X1 U22859 ( .A1(n19895), .A2(n20123), .B1(n19882), .B2(n20117), .ZN(
        n19869) );
  INV_X1 U22860 ( .A(n19869), .ZN(n19871) );
  AOI22_X1 U22861 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19886), .B1(
        n20057), .B2(n19885), .ZN(n19870) );
  OAI211_X1 U22862 ( .C1(n20060), .C2(n19883), .A(n19871), .B(n19870), .ZN(
        P2_U3122) );
  OAI22_X1 U22863 ( .A1(n19895), .A2(n20130), .B1(n19882), .B2(n20124), .ZN(
        n19872) );
  INV_X1 U22864 ( .A(n19872), .ZN(n19874) );
  AOI22_X1 U22865 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19886), .B1(
        n20063), .B2(n19885), .ZN(n19873) );
  OAI211_X1 U22866 ( .C1(n20066), .C2(n19883), .A(n19874), .B(n19873), .ZN(
        P2_U3123) );
  OAI22_X1 U22867 ( .A1(n19883), .A2(n20067), .B1(n19882), .B2(n20131), .ZN(
        n19875) );
  INV_X1 U22868 ( .A(n19875), .ZN(n19877) );
  AOI22_X1 U22869 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19886), .B1(
        n20069), .B2(n19885), .ZN(n19876) );
  OAI211_X1 U22870 ( .C1(n20137), .C2(n19895), .A(n19877), .B(n19876), .ZN(
        P2_U3124) );
  AOI22_X1 U22871 ( .A1(n20073), .A2(n19914), .B1(n19896), .B2(n20072), .ZN(
        n19879) );
  AOI22_X1 U22872 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19886), .B1(
        n20074), .B2(n19885), .ZN(n19878) );
  OAI211_X1 U22873 ( .C1(n20077), .C2(n19883), .A(n19879), .B(n19878), .ZN(
        P2_U3125) );
  AOI22_X1 U22874 ( .A1(n19977), .A2(n19914), .B1(n19896), .B2(n19976), .ZN(
        n19881) );
  AOI22_X1 U22875 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19886), .B1(
        n20081), .B2(n19885), .ZN(n19880) );
  OAI211_X1 U22876 ( .C1(n20079), .C2(n19883), .A(n19881), .B(n19880), .ZN(
        P2_U3126) );
  OAI22_X1 U22877 ( .A1(n19883), .A2(n20164), .B1(n19882), .B2(n20154), .ZN(
        n19884) );
  INV_X1 U22878 ( .A(n19884), .ZN(n19888) );
  AOI22_X1 U22879 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19886), .B1(
        n20087), .B2(n19885), .ZN(n19887) );
  OAI211_X1 U22880 ( .C1(n20029), .C2(n19895), .A(n19888), .B(n19887), .ZN(
        P2_U3127) );
  INV_X1 U22881 ( .A(n19889), .ZN(n19892) );
  INV_X1 U22882 ( .A(n19893), .ZN(n19890) );
  NAND2_X1 U22883 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19890), .ZN(
        n19924) );
  NOR2_X1 U22884 ( .A1(n19924), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19912) );
  OAI21_X1 U22885 ( .B1(n9621), .B2(n19912), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19891) );
  AOI22_X1 U22886 ( .A1(n19913), .A2(n20048), .B1(n19894), .B2(n19912), .ZN(
        n19899) );
  AOI21_X1 U22887 ( .B1(n19895), .B2(n19955), .A(n20036), .ZN(n19897) );
  AOI22_X1 U22888 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19915), .B1(
        n19914), .B2(n20106), .ZN(n19898) );
  OAI211_X1 U22889 ( .C1(n20109), .C2(n19955), .A(n19899), .B(n19898), .ZN(
        P2_U3128) );
  AOI22_X1 U22890 ( .A1(n19913), .A2(n20053), .B1(n19912), .B2(n20052), .ZN(
        n19901) );
  AOI22_X1 U22891 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19915), .B1(
        n19914), .B2(n20003), .ZN(n19900) );
  OAI211_X1 U22892 ( .C1(n20006), .C2(n19955), .A(n19901), .B(n19900), .ZN(
        P2_U3129) );
  AOI22_X1 U22893 ( .A1(n19913), .A2(n20057), .B1(n19912), .B2(n19958), .ZN(
        n19903) );
  AOI22_X1 U22894 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19915), .B1(
        n19914), .B2(n20120), .ZN(n19902) );
  OAI211_X1 U22895 ( .C1(n20123), .C2(n19955), .A(n19903), .B(n19902), .ZN(
        P2_U3130) );
  AOI22_X1 U22896 ( .A1(n19913), .A2(n20063), .B1(n19912), .B2(n19963), .ZN(
        n19905) );
  AOI22_X1 U22897 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19915), .B1(
        n19914), .B2(n20127), .ZN(n19904) );
  OAI211_X1 U22898 ( .C1(n20130), .C2(n19955), .A(n19905), .B(n19904), .ZN(
        P2_U3131) );
  AOI22_X1 U22899 ( .A1(n19913), .A2(n20069), .B1(n19912), .B2(n19968), .ZN(
        n19907) );
  AOI22_X1 U22900 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19915), .B1(
        n19914), .B2(n20134), .ZN(n19906) );
  OAI211_X1 U22901 ( .C1(n20137), .C2(n19955), .A(n19907), .B(n19906), .ZN(
        P2_U3132) );
  AOI22_X1 U22902 ( .A1(n19913), .A2(n20074), .B1(n19912), .B2(n20072), .ZN(
        n19909) );
  AOI22_X1 U22903 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19915), .B1(
        n19914), .B2(n20141), .ZN(n19908) );
  OAI211_X1 U22904 ( .C1(n20144), .C2(n19955), .A(n19909), .B(n19908), .ZN(
        P2_U3133) );
  AOI22_X1 U22905 ( .A1(n19913), .A2(n20081), .B1(n19912), .B2(n19976), .ZN(
        n19911) );
  AOI22_X1 U22906 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19915), .B1(
        n19914), .B2(n20148), .ZN(n19910) );
  OAI211_X1 U22907 ( .C1(n20153), .C2(n19955), .A(n19911), .B(n19910), .ZN(
        P2_U3134) );
  AOI22_X1 U22908 ( .A1(n19913), .A2(n20087), .B1(n19912), .B2(n20084), .ZN(
        n19917) );
  AOI22_X1 U22909 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19915), .B1(
        n19914), .B2(n20024), .ZN(n19916) );
  OAI211_X1 U22910 ( .C1(n20029), .C2(n19955), .A(n19917), .B(n19916), .ZN(
        P2_U3135) );
  NOR2_X1 U22911 ( .A1(n19924), .A2(n20034), .ZN(n19927) );
  OR2_X1 U22912 ( .A1(n19927), .A2(n20044), .ZN(n19918) );
  NOR2_X1 U22913 ( .A1(n19919), .A2(n19918), .ZN(n19923) );
  OAI21_X1 U22914 ( .B1(n19924), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20044), 
        .ZN(n19920) );
  INV_X1 U22915 ( .A(n19920), .ZN(n19921) );
  INV_X1 U22916 ( .A(n19927), .ZN(n19949) );
  OAI22_X1 U22917 ( .A1(n19950), .A2(n20095), .B1(n20094), .B2(n19949), .ZN(
        n19922) );
  INV_X1 U22918 ( .A(n19922), .ZN(n19930) );
  INV_X1 U22919 ( .A(n19994), .ZN(n20099) );
  NAND2_X1 U22920 ( .A1(n20099), .A2(n20252), .ZN(n19925) );
  AOI21_X1 U22921 ( .B1(n19925), .B2(n19924), .A(n19923), .ZN(n19926) );
  OAI211_X1 U22922 ( .C1(n19927), .C2(n20104), .A(n19926), .B(n20102), .ZN(
        n19952) );
  AOI22_X1 U22923 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19952), .B1(
        n19983), .B2(n19928), .ZN(n19929) );
  OAI211_X1 U22924 ( .C1(n20051), .C2(n19955), .A(n19930), .B(n19929), .ZN(
        P2_U3136) );
  OAI22_X1 U22925 ( .A1(n19950), .A2(n20111), .B1(n20110), .B2(n19949), .ZN(
        n19931) );
  INV_X1 U22926 ( .A(n19931), .ZN(n19933) );
  AOI22_X1 U22927 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19952), .B1(
        n19983), .B2(n20113), .ZN(n19932) );
  OAI211_X1 U22928 ( .C1(n20116), .C2(n19955), .A(n19933), .B(n19932), .ZN(
        P2_U3137) );
  OAI22_X1 U22929 ( .A1(n19950), .A2(n20118), .B1(n20117), .B2(n19949), .ZN(
        n19934) );
  INV_X1 U22930 ( .A(n19934), .ZN(n19936) );
  AOI22_X1 U22931 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19952), .B1(
        n19983), .B2(n19959), .ZN(n19935) );
  OAI211_X1 U22932 ( .C1(n20060), .C2(n19955), .A(n19936), .B(n19935), .ZN(
        P2_U3138) );
  OAI22_X1 U22933 ( .A1(n19950), .A2(n20125), .B1(n20124), .B2(n19949), .ZN(
        n19937) );
  INV_X1 U22934 ( .A(n19937), .ZN(n19939) );
  AOI22_X1 U22935 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19952), .B1(
        n19983), .B2(n19964), .ZN(n19938) );
  OAI211_X1 U22936 ( .C1(n20066), .C2(n19955), .A(n19939), .B(n19938), .ZN(
        P2_U3139) );
  OAI22_X1 U22937 ( .A1(n19950), .A2(n20132), .B1(n20131), .B2(n19949), .ZN(
        n19940) );
  INV_X1 U22938 ( .A(n19940), .ZN(n19942) );
  AOI22_X1 U22939 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19952), .B1(
        n19983), .B2(n19969), .ZN(n19941) );
  OAI211_X1 U22940 ( .C1(n20067), .C2(n19955), .A(n19942), .B(n19941), .ZN(
        P2_U3140) );
  OAI22_X1 U22941 ( .A1(n19950), .A2(n20139), .B1(n20138), .B2(n19949), .ZN(
        n19943) );
  INV_X1 U22942 ( .A(n19943), .ZN(n19945) );
  AOI22_X1 U22943 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19952), .B1(
        n19983), .B2(n20073), .ZN(n19944) );
  OAI211_X1 U22944 ( .C1(n20077), .C2(n19955), .A(n19945), .B(n19944), .ZN(
        P2_U3141) );
  OAI22_X1 U22945 ( .A1(n19950), .A2(n20146), .B1(n20145), .B2(n19949), .ZN(
        n19946) );
  INV_X1 U22946 ( .A(n19946), .ZN(n19948) );
  AOI22_X1 U22947 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19952), .B1(
        n19983), .B2(n19977), .ZN(n19947) );
  OAI211_X1 U22948 ( .C1(n20079), .C2(n19955), .A(n19948), .B(n19947), .ZN(
        P2_U3142) );
  OAI22_X1 U22949 ( .A1(n19950), .A2(n20156), .B1(n20154), .B2(n19949), .ZN(
        n19951) );
  INV_X1 U22950 ( .A(n19951), .ZN(n19954) );
  AOI22_X1 U22951 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19952), .B1(
        n19983), .B2(n20159), .ZN(n19953) );
  OAI211_X1 U22952 ( .C1(n20164), .C2(n19955), .A(n19954), .B(n19953), .ZN(
        P2_U3143) );
  AOI22_X1 U22953 ( .A1(n19982), .A2(n20053), .B1(n19981), .B2(n20052), .ZN(
        n19957) );
  AOI22_X1 U22954 ( .A1(n20025), .A2(n20113), .B1(n19983), .B2(n20003), .ZN(
        n19956) );
  OAI211_X1 U22955 ( .C1(n19987), .C2(n11855), .A(n19957), .B(n19956), .ZN(
        P2_U3145) );
  INV_X1 U22956 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n19962) );
  AOI22_X1 U22957 ( .A1(n19982), .A2(n20057), .B1(n19981), .B2(n19958), .ZN(
        n19961) );
  AOI22_X1 U22958 ( .A1(n19983), .A2(n20120), .B1(n20025), .B2(n19959), .ZN(
        n19960) );
  OAI211_X1 U22959 ( .C1(n19987), .C2(n19962), .A(n19961), .B(n19960), .ZN(
        P2_U3146) );
  INV_X1 U22960 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n19967) );
  AOI22_X1 U22961 ( .A1(n19982), .A2(n20063), .B1(n19981), .B2(n19963), .ZN(
        n19966) );
  AOI22_X1 U22962 ( .A1(n20025), .A2(n19964), .B1(n19983), .B2(n20127), .ZN(
        n19965) );
  OAI211_X1 U22963 ( .C1(n19987), .C2(n19967), .A(n19966), .B(n19965), .ZN(
        P2_U3147) );
  INV_X1 U22964 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n19972) );
  AOI22_X1 U22965 ( .A1(n19982), .A2(n20069), .B1(n19981), .B2(n19968), .ZN(
        n19971) );
  AOI22_X1 U22966 ( .A1(n20025), .A2(n19969), .B1(n19983), .B2(n20134), .ZN(
        n19970) );
  OAI211_X1 U22967 ( .C1(n19987), .C2(n19972), .A(n19971), .B(n19970), .ZN(
        P2_U3148) );
  INV_X1 U22968 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n19975) );
  AOI22_X1 U22969 ( .A1(n19982), .A2(n20074), .B1(n19981), .B2(n20072), .ZN(
        n19974) );
  AOI22_X1 U22970 ( .A1(n20025), .A2(n20073), .B1(n19983), .B2(n20141), .ZN(
        n19973) );
  OAI211_X1 U22971 ( .C1(n19987), .C2(n19975), .A(n19974), .B(n19973), .ZN(
        P2_U3149) );
  INV_X1 U22972 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n19980) );
  AOI22_X1 U22973 ( .A1(n19982), .A2(n20081), .B1(n19981), .B2(n19976), .ZN(
        n19979) );
  AOI22_X1 U22974 ( .A1(n20025), .A2(n19977), .B1(n19983), .B2(n20148), .ZN(
        n19978) );
  OAI211_X1 U22975 ( .C1(n19987), .C2(n19980), .A(n19979), .B(n19978), .ZN(
        P2_U3150) );
  INV_X1 U22976 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n19986) );
  AOI22_X1 U22977 ( .A1(n19982), .A2(n20087), .B1(n19981), .B2(n20084), .ZN(
        n19985) );
  AOI22_X1 U22978 ( .A1(n20025), .A2(n20159), .B1(n19983), .B2(n20024), .ZN(
        n19984) );
  OAI211_X1 U22979 ( .C1(n19987), .C2(n19986), .A(n19985), .B(n19984), .ZN(
        P2_U3151) );
  OR2_X2 U22980 ( .A1(n19988), .A2(n19993), .ZN(n20091) );
  NAND2_X1 U22981 ( .A1(n19998), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20046) );
  NAND2_X1 U22982 ( .A1(n20046), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19989) );
  NOR2_X1 U22983 ( .A1(n19990), .A2(n19989), .ZN(n19995) );
  AOI21_X1 U22984 ( .B1(n19998), .B2(n20104), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19991) );
  OAI22_X1 U22985 ( .A1(n20022), .A2(n20095), .B1(n20094), .B2(n20046), .ZN(
        n19992) );
  INV_X1 U22986 ( .A(n19992), .ZN(n20001) );
  NOR2_X1 U22987 ( .A1(n19994), .A2(n19993), .ZN(n19999) );
  AOI211_X1 U22988 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20046), .A(n19996), 
        .B(n19995), .ZN(n19997) );
  AOI22_X1 U22989 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20026), .B1(
        n20025), .B2(n20106), .ZN(n20000) );
  OAI211_X1 U22990 ( .C1(n20109), .C2(n20091), .A(n20001), .B(n20000), .ZN(
        P2_U3152) );
  OAI22_X1 U22991 ( .A1(n20022), .A2(n20111), .B1(n20046), .B2(n20110), .ZN(
        n20002) );
  INV_X1 U22992 ( .A(n20002), .ZN(n20005) );
  AOI22_X1 U22993 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20026), .B1(
        n20025), .B2(n20003), .ZN(n20004) );
  OAI211_X1 U22994 ( .C1(n20006), .C2(n20091), .A(n20005), .B(n20004), .ZN(
        P2_U3153) );
  OAI22_X1 U22995 ( .A1(n20022), .A2(n20118), .B1(n20046), .B2(n20117), .ZN(
        n20007) );
  INV_X1 U22996 ( .A(n20007), .ZN(n20009) );
  AOI22_X1 U22997 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20026), .B1(
        n20025), .B2(n20120), .ZN(n20008) );
  OAI211_X1 U22998 ( .C1(n20123), .C2(n20091), .A(n20009), .B(n20008), .ZN(
        P2_U3154) );
  OAI22_X1 U22999 ( .A1(n20022), .A2(n20125), .B1(n20046), .B2(n20124), .ZN(
        n20010) );
  INV_X1 U23000 ( .A(n20010), .ZN(n20012) );
  AOI22_X1 U23001 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20026), .B1(
        n20025), .B2(n20127), .ZN(n20011) );
  OAI211_X1 U23002 ( .C1(n20130), .C2(n20091), .A(n20012), .B(n20011), .ZN(
        P2_U3155) );
  OAI22_X1 U23003 ( .A1(n20022), .A2(n20132), .B1(n20046), .B2(n20131), .ZN(
        n20013) );
  INV_X1 U23004 ( .A(n20013), .ZN(n20015) );
  AOI22_X1 U23005 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20026), .B1(
        n20025), .B2(n20134), .ZN(n20014) );
  OAI211_X1 U23006 ( .C1(n20137), .C2(n20091), .A(n20015), .B(n20014), .ZN(
        P2_U3156) );
  OAI22_X1 U23007 ( .A1(n20022), .A2(n20139), .B1(n20046), .B2(n20138), .ZN(
        n20016) );
  INV_X1 U23008 ( .A(n20016), .ZN(n20018) );
  AOI22_X1 U23009 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20026), .B1(
        n20025), .B2(n20141), .ZN(n20017) );
  OAI211_X1 U23010 ( .C1(n20144), .C2(n20091), .A(n20018), .B(n20017), .ZN(
        P2_U3157) );
  OAI22_X1 U23011 ( .A1(n20022), .A2(n20146), .B1(n20046), .B2(n20145), .ZN(
        n20019) );
  INV_X1 U23012 ( .A(n20019), .ZN(n20021) );
  AOI22_X1 U23013 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20026), .B1(
        n20025), .B2(n20148), .ZN(n20020) );
  OAI211_X1 U23014 ( .C1(n20153), .C2(n20091), .A(n20021), .B(n20020), .ZN(
        P2_U3158) );
  OAI22_X1 U23015 ( .A1(n20022), .A2(n20156), .B1(n20046), .B2(n20154), .ZN(
        n20023) );
  INV_X1 U23016 ( .A(n20023), .ZN(n20028) );
  AOI22_X1 U23017 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20026), .B1(
        n20025), .B2(n20024), .ZN(n20027) );
  OAI211_X1 U23018 ( .C1(n20029), .C2(n20091), .A(n20028), .B(n20027), .ZN(
        P2_U3159) );
  NOR2_X1 U23019 ( .A1(n20033), .A2(n20032), .ZN(n20097) );
  AND2_X1 U23020 ( .A1(n20097), .A2(n20034), .ZN(n20085) );
  INV_X1 U23021 ( .A(n20085), .ZN(n20078) );
  OAI22_X1 U23022 ( .A1(n20061), .A2(n20109), .B1(n20094), .B2(n20078), .ZN(
        n20035) );
  INV_X1 U23023 ( .A(n20035), .ZN(n20050) );
  AOI21_X1 U23024 ( .B1(n20061), .B2(n20091), .A(n20036), .ZN(n20038) );
  OAI21_X1 U23025 ( .B1(n20039), .B2(n20258), .A(n20104), .ZN(n20040) );
  AOI21_X1 U23026 ( .B1(n20042), .B2(n20046), .A(n20040), .ZN(n20041) );
  OAI21_X1 U23027 ( .B1(n20041), .B2(n20085), .A(n20102), .ZN(n20088) );
  INV_X1 U23028 ( .A(n20042), .ZN(n20047) );
  NOR2_X1 U23029 ( .A1(n20042), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20045) );
  AOI22_X1 U23030 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20088), .B1(
        n20048), .B2(n20086), .ZN(n20049) );
  OAI211_X1 U23031 ( .C1(n20051), .C2(n20091), .A(n20050), .B(n20049), .ZN(
        P2_U3160) );
  AOI22_X1 U23032 ( .A1(n20113), .A2(n20149), .B1(n20085), .B2(n20052), .ZN(
        n20055) );
  AOI22_X1 U23033 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20088), .B1(
        n20053), .B2(n20086), .ZN(n20054) );
  OAI211_X1 U23034 ( .C1(n20116), .C2(n20091), .A(n20055), .B(n20054), .ZN(
        P2_U3161) );
  OAI22_X1 U23035 ( .A1(n20061), .A2(n20123), .B1(n20078), .B2(n20117), .ZN(
        n20056) );
  INV_X1 U23036 ( .A(n20056), .ZN(n20059) );
  AOI22_X1 U23037 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20088), .B1(
        n20057), .B2(n20086), .ZN(n20058) );
  OAI211_X1 U23038 ( .C1(n20060), .C2(n20091), .A(n20059), .B(n20058), .ZN(
        P2_U3162) );
  OAI22_X1 U23039 ( .A1(n20061), .A2(n20130), .B1(n20078), .B2(n20124), .ZN(
        n20062) );
  INV_X1 U23040 ( .A(n20062), .ZN(n20065) );
  AOI22_X1 U23041 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20088), .B1(
        n20063), .B2(n20086), .ZN(n20064) );
  OAI211_X1 U23042 ( .C1(n20066), .C2(n20091), .A(n20065), .B(n20064), .ZN(
        P2_U3163) );
  OAI22_X1 U23043 ( .A1(n20091), .A2(n20067), .B1(n20078), .B2(n20131), .ZN(
        n20068) );
  INV_X1 U23044 ( .A(n20068), .ZN(n20071) );
  AOI22_X1 U23045 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20088), .B1(
        n20069), .B2(n20086), .ZN(n20070) );
  OAI211_X1 U23046 ( .C1(n20137), .C2(n20061), .A(n20071), .B(n20070), .ZN(
        P2_U3164) );
  AOI22_X1 U23047 ( .A1(n20073), .A2(n20149), .B1(n20085), .B2(n20072), .ZN(
        n20076) );
  AOI22_X1 U23048 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20088), .B1(
        n20074), .B2(n20086), .ZN(n20075) );
  OAI211_X1 U23049 ( .C1(n20077), .C2(n20091), .A(n20076), .B(n20075), .ZN(
        P2_U3165) );
  OAI22_X1 U23050 ( .A1(n20091), .A2(n20079), .B1(n20078), .B2(n20145), .ZN(
        n20080) );
  INV_X1 U23051 ( .A(n20080), .ZN(n20083) );
  AOI22_X1 U23052 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20088), .B1(
        n20081), .B2(n20086), .ZN(n20082) );
  OAI211_X1 U23053 ( .C1(n20153), .C2(n20061), .A(n20083), .B(n20082), .ZN(
        P2_U3166) );
  AOI22_X1 U23054 ( .A1(n20159), .A2(n20149), .B1(n20085), .B2(n20084), .ZN(
        n20090) );
  AOI22_X1 U23055 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20088), .B1(
        n20087), .B2(n20086), .ZN(n20089) );
  OAI211_X1 U23056 ( .C1(n20164), .C2(n20091), .A(n20090), .B(n20089), .ZN(
        P2_U3167) );
  NAND2_X1 U23057 ( .A1(n20155), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20092) );
  NOR2_X1 U23058 ( .A1(n9662), .A2(n20092), .ZN(n20100) );
  AOI21_X1 U23059 ( .B1(n20097), .B2(n20104), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20093) );
  OAI22_X1 U23060 ( .A1(n20157), .A2(n20095), .B1(n20155), .B2(n20094), .ZN(
        n20096) );
  INV_X1 U23061 ( .A(n20096), .ZN(n20108) );
  AOI21_X1 U23062 ( .B1(n20099), .B2(n20098), .A(n20097), .ZN(n20101) );
  NOR2_X1 U23063 ( .A1(n20101), .A2(n20100), .ZN(n20103) );
  OAI211_X1 U23064 ( .C1(n20105), .C2(n20104), .A(n20103), .B(n20102), .ZN(
        n20161) );
  AOI22_X1 U23065 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20161), .B1(
        n20149), .B2(n20106), .ZN(n20107) );
  OAI211_X1 U23066 ( .C1(n20109), .C2(n20152), .A(n20108), .B(n20107), .ZN(
        P2_U3168) );
  OAI22_X1 U23067 ( .A1(n20157), .A2(n20111), .B1(n20155), .B2(n20110), .ZN(
        n20112) );
  INV_X1 U23068 ( .A(n20112), .ZN(n20115) );
  INV_X1 U23069 ( .A(n20152), .ZN(n20160) );
  AOI22_X1 U23070 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20161), .B1(
        n20160), .B2(n20113), .ZN(n20114) );
  OAI211_X1 U23071 ( .C1(n20116), .C2(n20061), .A(n20115), .B(n20114), .ZN(
        P2_U3169) );
  OAI22_X1 U23072 ( .A1(n20157), .A2(n20118), .B1(n20155), .B2(n20117), .ZN(
        n20119) );
  INV_X1 U23073 ( .A(n20119), .ZN(n20122) );
  AOI22_X1 U23074 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20161), .B1(
        n20149), .B2(n20120), .ZN(n20121) );
  OAI211_X1 U23075 ( .C1(n20123), .C2(n20152), .A(n20122), .B(n20121), .ZN(
        P2_U3170) );
  OAI22_X1 U23076 ( .A1(n20157), .A2(n20125), .B1(n20155), .B2(n20124), .ZN(
        n20126) );
  INV_X1 U23077 ( .A(n20126), .ZN(n20129) );
  AOI22_X1 U23078 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20161), .B1(
        n20149), .B2(n20127), .ZN(n20128) );
  OAI211_X1 U23079 ( .C1(n20130), .C2(n20152), .A(n20129), .B(n20128), .ZN(
        P2_U3171) );
  OAI22_X1 U23080 ( .A1(n20157), .A2(n20132), .B1(n20155), .B2(n20131), .ZN(
        n20133) );
  INV_X1 U23081 ( .A(n20133), .ZN(n20136) );
  AOI22_X1 U23082 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20161), .B1(
        n20149), .B2(n20134), .ZN(n20135) );
  OAI211_X1 U23083 ( .C1(n20137), .C2(n20152), .A(n20136), .B(n20135), .ZN(
        P2_U3172) );
  OAI22_X1 U23084 ( .A1(n20157), .A2(n20139), .B1(n20155), .B2(n20138), .ZN(
        n20140) );
  INV_X1 U23085 ( .A(n20140), .ZN(n20143) );
  AOI22_X1 U23086 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20161), .B1(
        n20149), .B2(n20141), .ZN(n20142) );
  OAI211_X1 U23087 ( .C1(n20144), .C2(n20152), .A(n20143), .B(n20142), .ZN(
        P2_U3173) );
  OAI22_X1 U23088 ( .A1(n20157), .A2(n20146), .B1(n20155), .B2(n20145), .ZN(
        n20147) );
  INV_X1 U23089 ( .A(n20147), .ZN(n20151) );
  AOI22_X1 U23090 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20161), .B1(
        n20149), .B2(n20148), .ZN(n20150) );
  OAI211_X1 U23091 ( .C1(n20153), .C2(n20152), .A(n20151), .B(n20150), .ZN(
        P2_U3174) );
  OAI22_X1 U23092 ( .A1(n20157), .A2(n20156), .B1(n20155), .B2(n20154), .ZN(
        n20158) );
  INV_X1 U23093 ( .A(n20158), .ZN(n20163) );
  AOI22_X1 U23094 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20161), .B1(
        n20160), .B2(n20159), .ZN(n20162) );
  OAI211_X1 U23095 ( .C1(n20164), .C2(n20061), .A(n20163), .B(n20162), .ZN(
        P2_U3175) );
  AND2_X1 U23096 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20165), .ZN(
        P2_U3179) );
  AND2_X1 U23097 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20165), .ZN(
        P2_U3180) );
  AND2_X1 U23098 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20165), .ZN(
        P2_U3181) );
  AND2_X1 U23099 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20165), .ZN(
        P2_U3182) );
  AND2_X1 U23100 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20165), .ZN(
        P2_U3183) );
  AND2_X1 U23101 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20165), .ZN(
        P2_U3184) );
  AND2_X1 U23102 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20165), .ZN(
        P2_U3185) );
  AND2_X1 U23103 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20165), .ZN(
        P2_U3186) );
  AND2_X1 U23104 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20165), .ZN(
        P2_U3187) );
  AND2_X1 U23105 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20165), .ZN(
        P2_U3188) );
  AND2_X1 U23106 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20165), .ZN(
        P2_U3189) );
  AND2_X1 U23107 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20165), .ZN(
        P2_U3190) );
  AND2_X1 U23108 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20165), .ZN(
        P2_U3191) );
  AND2_X1 U23109 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20165), .ZN(
        P2_U3192) );
  AND2_X1 U23110 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20165), .ZN(
        P2_U3193) );
  AND2_X1 U23111 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20165), .ZN(
        P2_U3194) );
  AND2_X1 U23112 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20165), .ZN(
        P2_U3195) );
  AND2_X1 U23113 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20165), .ZN(
        P2_U3196) );
  INV_X1 U23114 ( .A(P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n21323) );
  NOR2_X1 U23115 ( .A1(n21323), .A2(n20250), .ZN(P2_U3197) );
  AND2_X1 U23116 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20165), .ZN(
        P2_U3198) );
  AND2_X1 U23117 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20165), .ZN(
        P2_U3199) );
  AND2_X1 U23118 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20165), .ZN(
        P2_U3200) );
  AND2_X1 U23119 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20165), .ZN(P2_U3201) );
  AND2_X1 U23120 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20165), .ZN(P2_U3202) );
  AND2_X1 U23121 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20165), .ZN(P2_U3203) );
  AND2_X1 U23122 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20165), .ZN(P2_U3204) );
  AND2_X1 U23123 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20165), .ZN(P2_U3205) );
  AND2_X1 U23124 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20165), .ZN(P2_U3206) );
  AND2_X1 U23125 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20165), .ZN(P2_U3207) );
  AND2_X1 U23126 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20165), .ZN(P2_U3208) );
  NAND2_X1 U23127 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20166), .ZN(n20176) );
  INV_X1 U23128 ( .A(n20176), .ZN(n20181) );
  INV_X1 U23129 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20168) );
  NOR3_X1 U23130 ( .A1(n20181), .A2(n20168), .A3(n20167), .ZN(n20170) );
  OAI211_X1 U23131 ( .C1(HOLD), .C2(n20168), .A(n20284), .B(n20177), .ZN(
        n20169) );
  NAND2_X1 U23132 ( .A1(NA), .A2(n20171), .ZN(n20179) );
  OAI211_X1 U23133 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n20170), .A(n20169), 
        .B(n20179), .ZN(P2_U3209) );
  NAND2_X1 U23134 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n21090), .ZN(n20180) );
  OAI21_X1 U23135 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n20171), .A(n20180), 
        .ZN(n20172) );
  AOI21_X1 U23136 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(n20172), .A(n20181), .ZN(n20174) );
  OAI211_X1 U23137 ( .C1(n21090), .C2(n20175), .A(n20174), .B(n20173), .ZN(
        P2_U3210) );
  OAI22_X1 U23138 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20177), .B1(NA), 
        .B2(n20176), .ZN(n20178) );
  OAI211_X1 U23139 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20178), .ZN(n20183) );
  OAI211_X1 U23140 ( .C1(n20181), .C2(n20180), .A(P2_STATE_REG_2__SCAN_IN), 
        .B(n20179), .ZN(n20182) );
  NAND2_X1 U23141 ( .A1(n20183), .A2(n20182), .ZN(P2_U3211) );
  NAND2_X2 U23142 ( .A1(n20287), .A2(n21286), .ZN(n20240) );
  INV_X1 U23143 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20186) );
  OAI222_X1 U23144 ( .A1(n20240), .A2(n20186), .B1(n20185), .B2(n20287), .C1(
        n20184), .C2(n20237), .ZN(P2_U3212) );
  OAI222_X1 U23145 ( .A1(n20240), .A2(n20188), .B1(n20187), .B2(n20287), .C1(
        n20186), .C2(n20237), .ZN(P2_U3213) );
  OAI222_X1 U23146 ( .A1(n20240), .A2(n20190), .B1(n20189), .B2(n20287), .C1(
        n20188), .C2(n20237), .ZN(P2_U3214) );
  OAI222_X1 U23147 ( .A1(n20240), .A2(n12040), .B1(n20191), .B2(n20287), .C1(
        n20190), .C2(n20237), .ZN(P2_U3215) );
  OAI222_X1 U23148 ( .A1(n20240), .A2(n20193), .B1(n20192), .B2(n20287), .C1(
        n12040), .C2(n20237), .ZN(P2_U3216) );
  OAI222_X1 U23149 ( .A1(n20240), .A2(n20195), .B1(n20194), .B2(n20287), .C1(
        n20193), .C2(n20237), .ZN(P2_U3217) );
  OAI222_X1 U23150 ( .A1(n20240), .A2(n20197), .B1(n20196), .B2(n20287), .C1(
        n20195), .C2(n20237), .ZN(P2_U3218) );
  OAI222_X1 U23151 ( .A1(n20240), .A2(n20199), .B1(n20198), .B2(n20287), .C1(
        n20197), .C2(n20237), .ZN(P2_U3219) );
  INV_X1 U23152 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20201) );
  OAI222_X1 U23153 ( .A1(n20240), .A2(n20201), .B1(n20200), .B2(n20287), .C1(
        n20199), .C2(n20237), .ZN(P2_U3220) );
  INV_X1 U23154 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n20203) );
  OAI222_X1 U23155 ( .A1(n20240), .A2(n20203), .B1(n20202), .B2(n20287), .C1(
        n20201), .C2(n20237), .ZN(P2_U3221) );
  OAI222_X1 U23156 ( .A1(n20240), .A2(n20205), .B1(n20204), .B2(n20287), .C1(
        n20203), .C2(n20237), .ZN(P2_U3222) );
  OAI222_X1 U23157 ( .A1(n20240), .A2(n20207), .B1(n20206), .B2(n20287), .C1(
        n20205), .C2(n20237), .ZN(P2_U3223) );
  OAI222_X1 U23158 ( .A1(n20240), .A2(n21272), .B1(n20208), .B2(n20287), .C1(
        n20207), .C2(n20237), .ZN(P2_U3224) );
  OAI222_X1 U23159 ( .A1(n20240), .A2(n20210), .B1(n20209), .B2(n20287), .C1(
        n21272), .C2(n20237), .ZN(P2_U3225) );
  OAI222_X1 U23160 ( .A1(n20240), .A2(n12163), .B1(n20211), .B2(n20287), .C1(
        n20210), .C2(n20237), .ZN(P2_U3226) );
  INV_X1 U23161 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20213) );
  OAI222_X1 U23162 ( .A1(n20240), .A2(n20213), .B1(n20212), .B2(n20287), .C1(
        n12163), .C2(n20237), .ZN(P2_U3227) );
  OAI222_X1 U23163 ( .A1(n20240), .A2(n20215), .B1(n20214), .B2(n20287), .C1(
        n20213), .C2(n20237), .ZN(P2_U3228) );
  OAI222_X1 U23164 ( .A1(n20240), .A2(n20217), .B1(n20216), .B2(n20287), .C1(
        n20215), .C2(n20237), .ZN(P2_U3229) );
  OAI222_X1 U23165 ( .A1(n20240), .A2(n20219), .B1(n20218), .B2(n20287), .C1(
        n20217), .C2(n20237), .ZN(P2_U3230) );
  INV_X1 U23166 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20221) );
  NOR2_X1 U23167 ( .A1(n20219), .A2(n21286), .ZN(n21206) );
  AOI22_X1 U23168 ( .A1(n20287), .A2(n21206), .B1(P2_ADDRESS_REG_19__SCAN_IN), 
        .B2(n20284), .ZN(n20220) );
  OAI21_X1 U23169 ( .B1(n20221), .B2(n20240), .A(n20220), .ZN(P2_U3231) );
  INV_X1 U23170 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20223) );
  OAI222_X1 U23171 ( .A1(n20240), .A2(n20223), .B1(n20222), .B2(n20287), .C1(
        n20221), .C2(n20237), .ZN(P2_U3232) );
  OAI222_X1 U23172 ( .A1(n20240), .A2(n20225), .B1(n20224), .B2(n20287), .C1(
        n20223), .C2(n20237), .ZN(P2_U3233) );
  INV_X1 U23173 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20227) );
  OAI222_X1 U23174 ( .A1(n20240), .A2(n20227), .B1(n20226), .B2(n20287), .C1(
        n20225), .C2(n20237), .ZN(P2_U3234) );
  INV_X1 U23175 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20229) );
  OAI222_X1 U23176 ( .A1(n20240), .A2(n20229), .B1(n20228), .B2(n20287), .C1(
        n20227), .C2(n20237), .ZN(P2_U3235) );
  OAI222_X1 U23177 ( .A1(n20240), .A2(n20230), .B1(n21239), .B2(n20287), .C1(
        n20229), .C2(n20237), .ZN(P2_U3236) );
  OAI222_X1 U23178 ( .A1(n20240), .A2(n20233), .B1(n20231), .B2(n20287), .C1(
        n20230), .C2(n20237), .ZN(P2_U3237) );
  OAI222_X1 U23179 ( .A1(n20237), .A2(n20233), .B1(n20232), .B2(n20287), .C1(
        n20234), .C2(n20240), .ZN(P2_U3238) );
  INV_X1 U23180 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20235) );
  OAI222_X1 U23181 ( .A1(n20240), .A2(n20235), .B1(n21252), .B2(n20287), .C1(
        n20234), .C2(n20237), .ZN(P2_U3239) );
  INV_X1 U23182 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20238) );
  OAI222_X1 U23183 ( .A1(n20240), .A2(n20238), .B1(n20236), .B2(n20287), .C1(
        n20235), .C2(n20237), .ZN(P2_U3240) );
  OAI222_X1 U23184 ( .A1(n20240), .A2(n14359), .B1(n20239), .B2(n20287), .C1(
        n20238), .C2(n20237), .ZN(P2_U3241) );
  INV_X1 U23185 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20241) );
  AOI22_X1 U23186 ( .A1(n20287), .A2(n20242), .B1(n20241), .B2(n20284), .ZN(
        P2_U3585) );
  MUX2_X1 U23187 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20287), .Z(P2_U3586) );
  INV_X1 U23188 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20243) );
  AOI22_X1 U23189 ( .A1(n20287), .A2(n20244), .B1(n20243), .B2(n20284), .ZN(
        P2_U3587) );
  INV_X1 U23190 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20245) );
  AOI22_X1 U23191 ( .A1(n20287), .A2(n20246), .B1(n20245), .B2(n20284), .ZN(
        P2_U3588) );
  OAI21_X1 U23192 ( .B1(n20250), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20248), 
        .ZN(n20247) );
  INV_X1 U23193 ( .A(n20247), .ZN(P2_U3591) );
  OAI21_X1 U23194 ( .B1(n20250), .B2(n20249), .A(n20248), .ZN(P2_U3592) );
  NAND2_X1 U23195 ( .A1(n20252), .A2(n20251), .ZN(n20265) );
  NAND3_X1 U23196 ( .A1(n20254), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20253), 
        .ZN(n20256) );
  NAND2_X1 U23197 ( .A1(n20256), .A2(n20255), .ZN(n20263) );
  NAND2_X1 U23198 ( .A1(n20265), .A2(n20263), .ZN(n20260) );
  AOI222_X1 U23199 ( .A1(n20260), .A2(n10027), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20259), .C1(n20258), .C2(n20257), .ZN(n20261) );
  AOI22_X1 U23200 ( .A1(n20272), .A2(n20262), .B1(n20261), .B2(n20269), .ZN(
        P2_U3602) );
  NOR2_X1 U23201 ( .A1(n20264), .A2(n20263), .ZN(n20267) );
  INV_X1 U23202 ( .A(n20265), .ZN(n20266) );
  AOI211_X1 U23203 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20268), .A(n20267), 
        .B(n20266), .ZN(n20270) );
  AOI22_X1 U23204 ( .A1(n20272), .A2(n20271), .B1(n20270), .B2(n20269), .ZN(
        P2_U3603) );
  INV_X1 U23205 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20273) );
  AOI22_X1 U23206 ( .A1(n20287), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20273), 
        .B2(n20284), .ZN(P2_U3608) );
  INV_X1 U23207 ( .A(n20274), .ZN(n20281) );
  INV_X1 U23208 ( .A(n20275), .ZN(n20277) );
  AOI22_X1 U23209 ( .A1(n20279), .A2(n20278), .B1(n20277), .B2(n20276), .ZN(
        n20280) );
  NAND2_X1 U23210 ( .A1(n20281), .A2(n20280), .ZN(n20283) );
  MUX2_X1 U23211 ( .A(P2_MORE_REG_SCAN_IN), .B(n20283), .S(n20282), .Z(
        P2_U3609) );
  INV_X1 U23212 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n20285) );
  AOI22_X1 U23213 ( .A1(n20287), .A2(n20286), .B1(n20285), .B2(n20284), .ZN(
        P2_U3611) );
  AOI21_X1 U23214 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21092), .A(n21080), 
        .ZN(n21082) );
  INV_X1 U23215 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n21243) );
  INV_X2 U23216 ( .A(n21170), .ZN(n21172) );
  AOI21_X1 U23217 ( .B1(n21082), .B2(n21243), .A(n21172), .ZN(P1_U2802) );
  OAI21_X1 U23218 ( .B1(n20289), .B2(n20288), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20290) );
  OAI21_X1 U23219 ( .B1(n20291), .B2(n10144), .A(n20290), .ZN(P1_U2803) );
  NOR2_X1 U23220 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n21084) );
  OAI21_X1 U23221 ( .B1(n21084), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21170), .ZN(
        n20292) );
  OAI21_X1 U23222 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21170), .A(n20292), 
        .ZN(P1_U2804) );
  OAI21_X1 U23223 ( .B1(BS16), .B2(n21084), .A(n21157), .ZN(n21155) );
  OAI21_X1 U23224 ( .B1(n21157), .B2(n20979), .A(n21155), .ZN(P1_U2805) );
  OAI21_X1 U23225 ( .B1(n20294), .B2(n15541), .A(n20293), .ZN(P1_U2806) );
  NOR4_X1 U23226 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20298) );
  NOR4_X1 U23227 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20297) );
  NOR4_X1 U23228 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20296) );
  NOR4_X1 U23229 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20295) );
  NAND4_X1 U23230 ( .A1(n20298), .A2(n20297), .A3(n20296), .A4(n20295), .ZN(
        n20304) );
  NOR4_X1 U23231 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20302) );
  AOI211_X1 U23232 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_16__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20301) );
  NOR4_X1 U23233 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20300) );
  NOR4_X1 U23234 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20299) );
  NAND4_X1 U23235 ( .A1(n20302), .A2(n20301), .A3(n20300), .A4(n20299), .ZN(
        n20303) );
  NOR2_X1 U23236 ( .A1(n20304), .A2(n20303), .ZN(n21169) );
  INV_X1 U23237 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21150) );
  NOR3_X1 U23238 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20306) );
  OAI21_X1 U23239 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20306), .A(n21169), .ZN(
        n20305) );
  OAI21_X1 U23240 ( .B1(n21169), .B2(n21150), .A(n20305), .ZN(P1_U2807) );
  INV_X1 U23241 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21156) );
  AOI21_X1 U23242 ( .B1(n21162), .B2(n21156), .A(n20306), .ZN(n20307) );
  INV_X1 U23243 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21147) );
  INV_X1 U23244 ( .A(n21169), .ZN(n21164) );
  AOI22_X1 U23245 ( .A1(n21169), .A2(n20307), .B1(n21147), .B2(n21164), .ZN(
        P1_U2808) );
  AOI22_X1 U23246 ( .A1(n20308), .A2(n15238), .B1(n20350), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n20314) );
  AOI22_X1 U23247 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n20369), .B1(
        n20367), .B2(n20383), .ZN(n20313) );
  AOI21_X1 U23248 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n20309), .A(n16962), .ZN(
        n20312) );
  AOI22_X1 U23249 ( .A1(n20384), .A2(n20333), .B1(n20375), .B2(n20310), .ZN(
        n20311) );
  NAND4_X1 U23250 ( .A1(n20314), .A2(n20313), .A3(n20312), .A4(n20311), .ZN(
        P1_U2831) );
  AOI221_X1 U23251 ( .B1(n20351), .B2(n20327), .C1(n20315), .C2(n20327), .A(
        n20326), .ZN(n20329) );
  NOR4_X1 U23252 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20354), .A3(n20351), .A4(
        n20315), .ZN(n20316) );
  AOI211_X1 U23253 ( .C1(n20369), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n16962), .B(n20316), .ZN(n20318) );
  AOI22_X1 U23254 ( .A1(n20367), .A2(n9646), .B1(n20350), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n20317) );
  OAI211_X1 U23255 ( .C1(n20319), .C2(n20358), .A(n20318), .B(n20317), .ZN(
        n20320) );
  AOI21_X1 U23256 ( .B1(n20333), .B2(n20387), .A(n20320), .ZN(n20321) );
  OAI21_X1 U23257 ( .B1(n20329), .B2(n21225), .A(n20321), .ZN(P1_U2833) );
  AOI21_X1 U23258 ( .B1(n20369), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16962), .ZN(n20323) );
  NAND2_X1 U23259 ( .A1(n20350), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n20322) );
  OAI211_X1 U23260 ( .C1(n20325), .C2(n20324), .A(n20323), .B(n20322), .ZN(
        n20331) );
  INV_X1 U23261 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21102) );
  AOI21_X1 U23262 ( .B1(n20327), .B2(n20351), .A(n20326), .ZN(n20328) );
  NAND2_X1 U23263 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n20328), .ZN(n20341) );
  AOI21_X1 U23264 ( .B1(n21102), .B2(n20341), .A(n20329), .ZN(n20330) );
  AOI211_X1 U23265 ( .C1(n20333), .C2(n20332), .A(n20331), .B(n20330), .ZN(
        n20334) );
  OAI21_X1 U23266 ( .B1(n20335), .B2(n20358), .A(n20334), .ZN(P1_U2834) );
  OAI22_X1 U23267 ( .A1(n20338), .A2(n20395), .B1(n20337), .B2(n20336), .ZN(
        n20339) );
  AOI211_X1 U23268 ( .C1(n20367), .C2(n20390), .A(n16962), .B(n20339), .ZN(
        n20343) );
  INV_X1 U23269 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21100) );
  OAI21_X1 U23270 ( .B1(n20354), .B2(n20351), .A(n21100), .ZN(n20340) );
  AOI22_X1 U23271 ( .A1(n20393), .A2(n20377), .B1(n20341), .B2(n20340), .ZN(
        n20342) );
  OAI211_X1 U23272 ( .C1(n20344), .C2(n20358), .A(n20343), .B(n20342), .ZN(
        P1_U2835) );
  NAND4_X1 U23273 ( .A1(n20345), .A2(P1_REIP_REG_3__SCAN_IN), .A3(
        P1_REIP_REG_2__SCAN_IN), .A4(P1_REIP_REG_1__SCAN_IN), .ZN(n20352) );
  NAND2_X1 U23274 ( .A1(n20346), .A2(n20352), .ZN(n20381) );
  NAND2_X1 U23275 ( .A1(n20369), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20347) );
  OAI211_X1 U23276 ( .C1(n20381), .C2(n21097), .A(n20348), .B(n20347), .ZN(
        n20349) );
  AOI21_X1 U23277 ( .B1(n20350), .B2(P1_EBX_REG_4__SCAN_IN), .A(n20349), .ZN(
        n20365) );
  INV_X1 U23278 ( .A(n20351), .ZN(n20353) );
  NOR3_X1 U23279 ( .A1(n20354), .A2(n20353), .A3(n20352), .ZN(n20355) );
  AOI21_X1 U23280 ( .B1(n20368), .B2(n20356), .A(n20355), .ZN(n20357) );
  INV_X1 U23281 ( .A(n20357), .ZN(n20363) );
  OAI22_X1 U23282 ( .A1(n20361), .A2(n20360), .B1(n20359), .B2(n20358), .ZN(
        n20362) );
  AOI211_X1 U23283 ( .C1(n20367), .C2(n20465), .A(n20363), .B(n20362), .ZN(
        n20364) );
  NAND2_X1 U23284 ( .A1(n20365), .A2(n20364), .ZN(P1_U2836) );
  AOI21_X1 U23285 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(n20366), .A(
        P1_REIP_REG_3__SCAN_IN), .ZN(n20382) );
  NAND2_X1 U23286 ( .A1(n20367), .A2(n20472), .ZN(n20373) );
  NAND2_X1 U23287 ( .A1(n20350), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n20372) );
  NAND2_X1 U23288 ( .A1(n20774), .A2(n20368), .ZN(n20371) );
  NAND2_X1 U23289 ( .A1(n20369), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n20370) );
  AND4_X1 U23290 ( .A1(n20373), .A2(n20372), .A3(n20371), .A4(n20370), .ZN(
        n20380) );
  INV_X1 U23291 ( .A(n20374), .ZN(n20376) );
  AOI22_X1 U23292 ( .A1(n20378), .A2(n20377), .B1(n20376), .B2(n20375), .ZN(
        n20379) );
  OAI211_X1 U23293 ( .C1(n20382), .C2(n20381), .A(n20380), .B(n20379), .ZN(
        P1_U2837) );
  AOI22_X1 U23294 ( .A1(n20384), .A2(n20392), .B1(n20391), .B2(n20383), .ZN(
        n20385) );
  OAI21_X1 U23295 ( .B1(n20396), .B2(n20386), .A(n20385), .ZN(P1_U2863) );
  AOI22_X1 U23296 ( .A1(n20387), .A2(n20392), .B1(n20391), .B2(n9646), .ZN(
        n20388) );
  OAI21_X1 U23297 ( .B1(n20396), .B2(n20389), .A(n20388), .ZN(P1_U2865) );
  AOI22_X1 U23298 ( .A1(n20393), .A2(n20392), .B1(n20391), .B2(n20390), .ZN(
        n20394) );
  OAI21_X1 U23299 ( .B1(n20396), .B2(n20395), .A(n20394), .ZN(P1_U2867) );
  INV_X1 U23300 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n21337) );
  INV_X1 U23301 ( .A(n20397), .ZN(n20400) );
  AOI22_X1 U23302 ( .A1(n20400), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n21176), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20398) );
  OAI21_X1 U23303 ( .B1(n21337), .B2(n20399), .A(n20398), .ZN(P1_U2910) );
  INV_X1 U23304 ( .A(P1_UWORD_REG_4__SCAN_IN), .ZN(n21242) );
  AOI22_X1 U23305 ( .A1(n20426), .A2(P1_DATAO_REG_20__SCAN_IN), .B1(n20400), 
        .B2(P1_EAX_REG_20__SCAN_IN), .ZN(n20401) );
  OAI21_X1 U23306 ( .B1(n21242), .B2(n20410), .A(n20401), .ZN(P1_U2916) );
  AOI22_X1 U23307 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20408), .B1(n20426), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20402) );
  OAI21_X1 U23308 ( .B1(n20403), .B2(n20410), .A(n20402), .ZN(P1_U2921) );
  AOI22_X1 U23309 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20404) );
  OAI21_X1 U23310 ( .B1(n15025), .B2(n20428), .A(n20404), .ZN(P1_U2922) );
  INV_X1 U23311 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20406) );
  AOI22_X1 U23312 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20405) );
  OAI21_X1 U23313 ( .B1(n20406), .B2(n20428), .A(n20405), .ZN(P1_U2923) );
  INV_X1 U23314 ( .A(P1_LWORD_REG_12__SCAN_IN), .ZN(n21266) );
  AOI22_X1 U23315 ( .A1(P1_EAX_REG_12__SCAN_IN), .A2(n20408), .B1(n20426), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20407) );
  OAI21_X1 U23316 ( .B1(n21266), .B2(n20410), .A(n20407), .ZN(P1_U2924) );
  INV_X1 U23317 ( .A(P1_LWORD_REG_11__SCAN_IN), .ZN(n21321) );
  AOI22_X1 U23318 ( .A1(P1_EAX_REG_11__SCAN_IN), .A2(n20408), .B1(n20426), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20409) );
  OAI21_X1 U23319 ( .B1(n21321), .B2(n20410), .A(n20409), .ZN(P1_U2925) );
  INV_X1 U23320 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20412) );
  AOI22_X1 U23321 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20411) );
  OAI21_X1 U23322 ( .B1(n20412), .B2(n20428), .A(n20411), .ZN(P1_U2926) );
  INV_X1 U23323 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20414) );
  AOI22_X1 U23324 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20413) );
  OAI21_X1 U23325 ( .B1(n20414), .B2(n20428), .A(n20413), .ZN(P1_U2927) );
  AOI22_X1 U23326 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20415) );
  OAI21_X1 U23327 ( .B1(n14165), .B2(n20428), .A(n20415), .ZN(P1_U2928) );
  AOI22_X1 U23328 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20416) );
  OAI21_X1 U23329 ( .B1(n11088), .B2(n20428), .A(n20416), .ZN(P1_U2929) );
  AOI22_X1 U23330 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20417) );
  OAI21_X1 U23331 ( .B1(n20418), .B2(n20428), .A(n20417), .ZN(P1_U2930) );
  AOI22_X1 U23332 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20419) );
  OAI21_X1 U23333 ( .B1(n20420), .B2(n20428), .A(n20419), .ZN(P1_U2931) );
  AOI22_X1 U23334 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20421) );
  OAI21_X1 U23335 ( .B1(n20422), .B2(n20428), .A(n20421), .ZN(P1_U2932) );
  AOI22_X1 U23336 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20423) );
  OAI21_X1 U23337 ( .B1(n11002), .B2(n20428), .A(n20423), .ZN(P1_U2933) );
  AOI22_X1 U23338 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20424) );
  OAI21_X1 U23339 ( .B1(n10970), .B2(n20428), .A(n20424), .ZN(P1_U2934) );
  AOI22_X1 U23340 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20425) );
  OAI21_X1 U23341 ( .B1(n10977), .B2(n20428), .A(n20425), .ZN(P1_U2935) );
  AOI22_X1 U23342 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n21176), .B1(n20426), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20427) );
  OAI21_X1 U23343 ( .B1(n20429), .B2(n20428), .A(n20427), .ZN(P1_U2936) );
  AOI22_X1 U23344 ( .A1(n20454), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20453), .ZN(n20431) );
  NAND2_X1 U23345 ( .A1(n20439), .A2(n20430), .ZN(n20441) );
  NAND2_X1 U23346 ( .A1(n20431), .A2(n20441), .ZN(P1_U2945) );
  AOI22_X1 U23347 ( .A1(n20454), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20453), .ZN(n20433) );
  NAND2_X1 U23348 ( .A1(n20439), .A2(n20432), .ZN(n20445) );
  NAND2_X1 U23349 ( .A1(n20433), .A2(n20445), .ZN(P1_U2947) );
  AOI22_X1 U23350 ( .A1(n20454), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20453), .ZN(n20435) );
  NAND2_X1 U23351 ( .A1(n20439), .A2(n20434), .ZN(n20447) );
  NAND2_X1 U23352 ( .A1(n20435), .A2(n20447), .ZN(P1_U2948) );
  AOI22_X1 U23353 ( .A1(n20454), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20453), .ZN(n20437) );
  NAND2_X1 U23354 ( .A1(n20439), .A2(n20436), .ZN(n20449) );
  NAND2_X1 U23355 ( .A1(n20437), .A2(n20449), .ZN(P1_U2949) );
  AOI22_X1 U23356 ( .A1(n20454), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20453), .ZN(n20440) );
  NAND2_X1 U23357 ( .A1(n20439), .A2(n20438), .ZN(n20455) );
  NAND2_X1 U23358 ( .A1(n20440), .A2(n20455), .ZN(P1_U2951) );
  AOI22_X1 U23359 ( .A1(n20454), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20453), .ZN(n20442) );
  NAND2_X1 U23360 ( .A1(n20442), .A2(n20441), .ZN(P1_U2960) );
  AOI22_X1 U23361 ( .A1(n20454), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20453), .ZN(n20444) );
  NAND2_X1 U23362 ( .A1(n20444), .A2(n20443), .ZN(P1_U2961) );
  AOI22_X1 U23363 ( .A1(n20454), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20453), .ZN(n20446) );
  NAND2_X1 U23364 ( .A1(n20446), .A2(n20445), .ZN(P1_U2962) );
  AOI22_X1 U23365 ( .A1(n20454), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20453), .ZN(n20448) );
  NAND2_X1 U23366 ( .A1(n20448), .A2(n20447), .ZN(P1_U2963) );
  AOI22_X1 U23367 ( .A1(n20454), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20453), .ZN(n20450) );
  NAND2_X1 U23368 ( .A1(n20450), .A2(n20449), .ZN(P1_U2964) );
  AOI22_X1 U23369 ( .A1(n20454), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20453), .ZN(n20452) );
  NAND2_X1 U23370 ( .A1(n20452), .A2(n20451), .ZN(P1_U2965) );
  AOI22_X1 U23371 ( .A1(n20454), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20453), .ZN(n20456) );
  NAND2_X1 U23372 ( .A1(n20456), .A2(n20455), .ZN(P1_U2966) );
  OAI21_X1 U23373 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20457), .ZN(n20467) );
  AOI21_X1 U23374 ( .B1(n20460), .B2(n20459), .A(n20458), .ZN(n20475) );
  OAI22_X1 U23375 ( .A1(n20462), .A2(n20481), .B1(n20475), .B2(n20461), .ZN(
        n20463) );
  AOI211_X1 U23376 ( .C1(n20473), .C2(n20465), .A(n20464), .B(n20463), .ZN(
        n20466) );
  OAI21_X1 U23377 ( .B1(n20468), .B2(n20467), .A(n20466), .ZN(P1_U3027) );
  INV_X1 U23378 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21096) );
  NOR2_X1 U23379 ( .A1(n20348), .A2(n21096), .ZN(n20471) );
  OAI22_X1 U23380 ( .A1(n20469), .A2(n20481), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20468), .ZN(n20470) );
  AOI211_X1 U23381 ( .C1(n20473), .C2(n20472), .A(n20471), .B(n20470), .ZN(
        n20474) );
  OAI21_X1 U23382 ( .B1(n20475), .B2(n13206), .A(n20474), .ZN(P1_U3028) );
  INV_X1 U23383 ( .A(n20476), .ZN(n20480) );
  OAI21_X1 U23384 ( .B1(n20478), .B2(n20477), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20479) );
  OAI211_X1 U23385 ( .C1(n20482), .C2(n20481), .A(n20480), .B(n20479), .ZN(
        n20483) );
  INV_X1 U23386 ( .A(n20483), .ZN(n20485) );
  OAI211_X1 U23387 ( .C1(n20487), .C2(n20486), .A(n20485), .B(n20484), .ZN(
        P1_U3031) );
  NOR2_X1 U23388 ( .A1(n20489), .A2(n20488), .ZN(P1_U3032) );
  INV_X1 U23389 ( .A(n20492), .ZN(n20490) );
  AOI22_X1 U23390 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20531), .B1(DATAI_16_), 
        .B2(n20493), .ZN(n20942) );
  INV_X1 U23391 ( .A(n21023), .ZN(n20939) );
  NAND2_X1 U23392 ( .A1(n20533), .A2(n10837), .ZN(n20698) );
  NAND3_X1 U23393 ( .A1(n20873), .A2(n20836), .A3(n20901), .ZN(n20545) );
  NOR2_X1 U23394 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20545), .ZN(
        n20534) );
  AOI22_X1 U23395 ( .A1(n21065), .A2(n20939), .B1(n21014), .B2(n20534), .ZN(
        n20507) );
  NAND2_X1 U23396 ( .A1(n20503), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20976) );
  NAND2_X1 U23397 ( .A1(n20563), .A2(n20934), .ZN(n20498) );
  NAND2_X1 U23398 ( .A1(n20934), .A2(n20979), .ZN(n20902) );
  OAI21_X1 U23399 ( .B1(n21065), .B2(n20498), .A(n20902), .ZN(n20502) );
  OR2_X1 U23400 ( .A1(n20774), .A2(n20499), .ZN(n20540) );
  OR2_X1 U23401 ( .A1(n20540), .A2(n20981), .ZN(n20504) );
  NAND2_X1 U23402 ( .A1(n20833), .A2(n20775), .ZN(n20646) );
  AOI22_X1 U23403 ( .A1(n20502), .A2(n20504), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20646), .ZN(n20500) );
  NOR2_X2 U23404 ( .A1(n20649), .A2(n20501), .ZN(n21013) );
  INV_X1 U23405 ( .A(n20502), .ZN(n20505) );
  NOR2_X1 U23406 ( .A1(n20503), .A2(n21074), .ZN(n20834) );
  INV_X1 U23407 ( .A(n20834), .ZN(n20777) );
  AOI22_X1 U23408 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20537), .B1(
        n21013), .B2(n20536), .ZN(n20506) );
  OAI211_X1 U23409 ( .C1(n20942), .C2(n20563), .A(n20507), .B(n20506), .ZN(
        P1_U3033) );
  AOI22_X1 U23410 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20531), .B1(DATAI_17_), 
        .B2(n20493), .ZN(n20946) );
  AOI22_X1 U23411 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20531), .B1(DATAI_25_), 
        .B2(n20493), .ZN(n21029) );
  INV_X1 U23412 ( .A(n21029), .ZN(n20943) );
  NAND2_X1 U23413 ( .A1(n20533), .A2(n20508), .ZN(n20709) );
  AOI22_X1 U23414 ( .A1(n21065), .A2(n20943), .B1(n20534), .B2(n21025), .ZN(
        n20511) );
  NOR2_X2 U23415 ( .A1(n20649), .A2(n20509), .ZN(n21024) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20537), .B1(
        n21024), .B2(n20536), .ZN(n20510) );
  OAI211_X1 U23417 ( .C1(n20946), .C2(n20563), .A(n20511), .B(n20510), .ZN(
        P1_U3034) );
  AOI22_X1 U23418 ( .A1(DATAI_18_), .A2(n20493), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20531), .ZN(n20950) );
  AOI22_X1 U23419 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20531), .B1(DATAI_26_), 
        .B2(n20493), .ZN(n21035) );
  INV_X1 U23420 ( .A(n21035), .ZN(n20947) );
  NAND2_X1 U23421 ( .A1(n20533), .A2(n20512), .ZN(n20713) );
  AOI22_X1 U23422 ( .A1(n21065), .A2(n20947), .B1(n21031), .B2(n20534), .ZN(
        n20515) );
  NOR2_X2 U23423 ( .A1(n20649), .A2(n20513), .ZN(n21030) );
  AOI22_X1 U23424 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20537), .B1(
        n21030), .B2(n20536), .ZN(n20514) );
  OAI211_X1 U23425 ( .C1(n20950), .C2(n20563), .A(n20515), .B(n20514), .ZN(
        P1_U3035) );
  AOI22_X1 U23426 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20531), .B1(DATAI_19_), 
        .B2(n20493), .ZN(n20954) );
  AOI22_X1 U23427 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20531), .B1(DATAI_27_), 
        .B2(n20493), .ZN(n21041) );
  INV_X1 U23428 ( .A(n21041), .ZN(n20951) );
  NAND2_X1 U23429 ( .A1(n20533), .A2(n20516), .ZN(n20717) );
  AOI22_X1 U23430 ( .A1(n21065), .A2(n20951), .B1(n21037), .B2(n20534), .ZN(
        n20519) );
  NOR2_X2 U23431 ( .A1(n20649), .A2(n20517), .ZN(n21036) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20537), .B1(
        n21036), .B2(n20536), .ZN(n20518) );
  OAI211_X1 U23433 ( .C1(n20954), .C2(n20563), .A(n20519), .B(n20518), .ZN(
        P1_U3036) );
  AOI22_X1 U23434 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20531), .B1(DATAI_20_), 
        .B2(n20493), .ZN(n20958) );
  AOI22_X1 U23435 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20531), .B1(DATAI_28_), 
        .B2(n20493), .ZN(n21047) );
  INV_X1 U23436 ( .A(n21047), .ZN(n20955) );
  NAND2_X1 U23437 ( .A1(n20533), .A2(n20520), .ZN(n20721) );
  AOI22_X1 U23438 ( .A1(n21065), .A2(n20955), .B1(n20534), .B2(n21043), .ZN(
        n20523) );
  NOR2_X2 U23439 ( .A1(n20649), .A2(n20521), .ZN(n21042) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20537), .B1(
        n21042), .B2(n20536), .ZN(n20522) );
  OAI211_X1 U23441 ( .C1(n20958), .C2(n20563), .A(n20523), .B(n20522), .ZN(
        P1_U3037) );
  AOI22_X1 U23442 ( .A1(DATAI_21_), .A2(n20493), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20531), .ZN(n20962) );
  INV_X1 U23443 ( .A(n21053), .ZN(n20959) );
  NAND2_X1 U23444 ( .A1(n20533), .A2(n20524), .ZN(n20725) );
  AOI22_X1 U23445 ( .A1(n21065), .A2(n20959), .B1(n20534), .B2(n21049), .ZN(
        n20527) );
  NOR2_X2 U23446 ( .A1(n20649), .A2(n20525), .ZN(n21048) );
  AOI22_X1 U23447 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20537), .B1(
        n21048), .B2(n20536), .ZN(n20526) );
  OAI211_X1 U23448 ( .C1(n20962), .C2(n20563), .A(n20527), .B(n20526), .ZN(
        P1_U3038) );
  AOI22_X1 U23449 ( .A1(DATAI_22_), .A2(n20493), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20531), .ZN(n20966) );
  AOI22_X1 U23450 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20531), .B1(DATAI_30_), 
        .B2(n20493), .ZN(n21059) );
  INV_X1 U23451 ( .A(n21059), .ZN(n20963) );
  AOI22_X1 U23452 ( .A1(n21065), .A2(n20963), .B1(n21055), .B2(n20534), .ZN(
        n20530) );
  NOR2_X2 U23453 ( .A1(n20649), .A2(n20528), .ZN(n21054) );
  AOI22_X1 U23454 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20537), .B1(
        n21054), .B2(n20536), .ZN(n20529) );
  OAI211_X1 U23455 ( .C1(n20966), .C2(n20563), .A(n20530), .B(n20529), .ZN(
        P1_U3039) );
  AOI22_X1 U23456 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20531), .B1(DATAI_23_), 
        .B2(n20493), .ZN(n20974) );
  AOI22_X1 U23457 ( .A1(DATAI_31_), .A2(n20493), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20531), .ZN(n21070) );
  INV_X1 U23458 ( .A(n21070), .ZN(n20969) );
  NAND2_X1 U23459 ( .A1(n20533), .A2(n20532), .ZN(n20733) );
  AOI22_X1 U23460 ( .A1(n21065), .A2(n20969), .B1(n20534), .B2(n21063), .ZN(
        n20539) );
  NOR2_X2 U23461 ( .A1(n20649), .A2(n20535), .ZN(n21061) );
  AOI22_X1 U23462 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20537), .B1(
        n21061), .B2(n20536), .ZN(n20538) );
  OAI211_X1 U23463 ( .C1(n20974), .C2(n20563), .A(n20539), .B(n20538), .ZN(
        P1_U3040) );
  NOR2_X1 U23464 ( .A1(n20933), .A2(n20545), .ZN(n20565) );
  INV_X1 U23465 ( .A(n20541), .ZN(n20803) );
  AOI21_X1 U23466 ( .B1(n20609), .B2(n20803), .A(n20565), .ZN(n20542) );
  OAI22_X1 U23467 ( .A1(n20542), .A2(n21010), .B1(n20545), .B2(n21074), .ZN(
        n20564) );
  AOI22_X1 U23468 ( .A1(n21014), .A2(n20565), .B1(n21013), .B2(n20564), .ZN(
        n20549) );
  INV_X1 U23469 ( .A(n20543), .ZN(n20544) );
  NOR2_X1 U23470 ( .A1(n20610), .A2(n20544), .ZN(n20547) );
  INV_X1 U23471 ( .A(n20545), .ZN(n20546) );
  INV_X1 U23472 ( .A(n20599), .ZN(n20560) );
  INV_X1 U23473 ( .A(n20942), .ZN(n21020) );
  AOI22_X1 U23474 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20567), .B1(
        n20560), .B2(n21020), .ZN(n20548) );
  OAI211_X1 U23475 ( .C1(n21023), .C2(n20563), .A(n20549), .B(n20548), .ZN(
        P1_U3041) );
  AOI22_X1 U23476 ( .A1(n21025), .A2(n20565), .B1(n21024), .B2(n20564), .ZN(
        n20551) );
  INV_X1 U23477 ( .A(n20946), .ZN(n21026) );
  AOI22_X1 U23478 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20567), .B1(
        n20560), .B2(n21026), .ZN(n20550) );
  OAI211_X1 U23479 ( .C1(n21029), .C2(n20563), .A(n20551), .B(n20550), .ZN(
        P1_U3042) );
  AOI22_X1 U23480 ( .A1(n21031), .A2(n20565), .B1(n21030), .B2(n20564), .ZN(
        n20553) );
  INV_X1 U23481 ( .A(n20563), .ZN(n20566) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20567), .B1(
        n20566), .B2(n20947), .ZN(n20552) );
  OAI211_X1 U23483 ( .C1(n20950), .C2(n20599), .A(n20553), .B(n20552), .ZN(
        P1_U3043) );
  AOI22_X1 U23484 ( .A1(n21037), .A2(n20565), .B1(n21036), .B2(n20564), .ZN(
        n20555) );
  INV_X1 U23485 ( .A(n20954), .ZN(n21038) );
  AOI22_X1 U23486 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20567), .B1(
        n20560), .B2(n21038), .ZN(n20554) );
  OAI211_X1 U23487 ( .C1(n21041), .C2(n20563), .A(n20555), .B(n20554), .ZN(
        P1_U3044) );
  AOI22_X1 U23488 ( .A1(n21043), .A2(n20565), .B1(n21042), .B2(n20564), .ZN(
        n20557) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20567), .B1(
        n20566), .B2(n20955), .ZN(n20556) );
  OAI211_X1 U23490 ( .C1(n20958), .C2(n20599), .A(n20557), .B(n20556), .ZN(
        P1_U3045) );
  AOI22_X1 U23491 ( .A1(n21049), .A2(n20565), .B1(n21048), .B2(n20564), .ZN(
        n20559) );
  INV_X1 U23492 ( .A(n20962), .ZN(n21050) );
  AOI22_X1 U23493 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20567), .B1(
        n20560), .B2(n21050), .ZN(n20558) );
  OAI211_X1 U23494 ( .C1(n21053), .C2(n20563), .A(n20559), .B(n20558), .ZN(
        P1_U3046) );
  AOI22_X1 U23495 ( .A1(n21055), .A2(n20565), .B1(n21054), .B2(n20564), .ZN(
        n20562) );
  INV_X1 U23496 ( .A(n20966), .ZN(n21056) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20567), .B1(
        n20560), .B2(n21056), .ZN(n20561) );
  OAI211_X1 U23498 ( .C1(n21059), .C2(n20563), .A(n20562), .B(n20561), .ZN(
        P1_U3047) );
  AOI22_X1 U23499 ( .A1(n21063), .A2(n20565), .B1(n21061), .B2(n20564), .ZN(
        n20569) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20567), .B1(
        n20566), .B2(n20969), .ZN(n20568) );
  OAI211_X1 U23501 ( .C1(n20974), .C2(n20599), .A(n20569), .B(n20568), .ZN(
        P1_U3048) );
  NAND2_X1 U23502 ( .A1(n15553), .A2(n20570), .ZN(n20831) );
  NAND3_X1 U23503 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20873), .A3(
        n20836), .ZN(n20614) );
  OR2_X1 U23504 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20614), .ZN(
        n20598) );
  OAI22_X1 U23505 ( .A1(n20643), .A2(n20942), .B1(n20698), .B2(n20598), .ZN(
        n20571) );
  INV_X1 U23506 ( .A(n20571), .ZN(n20579) );
  NAND2_X1 U23507 ( .A1(n20643), .A2(n20599), .ZN(n20572) );
  AOI21_X1 U23508 ( .B1(n20572), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21010), 
        .ZN(n20574) );
  NAND2_X1 U23509 ( .A1(n20609), .A2(n20981), .ZN(n20576) );
  AOI22_X1 U23510 ( .A1(n20574), .A2(n20576), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20598), .ZN(n20573) );
  OAI21_X1 U23511 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20833), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20701) );
  NAND3_X1 U23512 ( .A1(n20842), .A2(n20573), .A3(n20701), .ZN(n20602) );
  INV_X1 U23513 ( .A(n20574), .ZN(n20577) );
  INV_X1 U23514 ( .A(n20833), .ZN(n20575) );
  NAND2_X1 U23515 ( .A1(n20575), .A2(n20873), .ZN(n20704) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20602), .B1(
        n21013), .B2(n20601), .ZN(n20578) );
  OAI211_X1 U23517 ( .C1(n21023), .C2(n20599), .A(n20579), .B(n20578), .ZN(
        P1_U3049) );
  OAI22_X1 U23518 ( .A1(n20599), .A2(n21029), .B1(n20709), .B2(n20598), .ZN(
        n20580) );
  INV_X1 U23519 ( .A(n20580), .ZN(n20582) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20602), .B1(
        n21024), .B2(n20601), .ZN(n20581) );
  OAI211_X1 U23521 ( .C1(n20946), .C2(n20643), .A(n20582), .B(n20581), .ZN(
        P1_U3050) );
  OAI22_X1 U23522 ( .A1(n20599), .A2(n21035), .B1(n20713), .B2(n20598), .ZN(
        n20583) );
  INV_X1 U23523 ( .A(n20583), .ZN(n20585) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20602), .B1(
        n21030), .B2(n20601), .ZN(n20584) );
  OAI211_X1 U23525 ( .C1(n20950), .C2(n20643), .A(n20585), .B(n20584), .ZN(
        P1_U3051) );
  OAI22_X1 U23526 ( .A1(n20599), .A2(n21041), .B1(n20717), .B2(n20598), .ZN(
        n20586) );
  INV_X1 U23527 ( .A(n20586), .ZN(n20588) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20602), .B1(
        n21036), .B2(n20601), .ZN(n20587) );
  OAI211_X1 U23529 ( .C1(n20954), .C2(n20643), .A(n20588), .B(n20587), .ZN(
        P1_U3052) );
  OAI22_X1 U23530 ( .A1(n20643), .A2(n20958), .B1(n20721), .B2(n20598), .ZN(
        n20589) );
  INV_X1 U23531 ( .A(n20589), .ZN(n20591) );
  AOI22_X1 U23532 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20602), .B1(
        n21042), .B2(n20601), .ZN(n20590) );
  OAI211_X1 U23533 ( .C1(n21047), .C2(n20599), .A(n20591), .B(n20590), .ZN(
        P1_U3053) );
  OAI22_X1 U23534 ( .A1(n20643), .A2(n20962), .B1(n20725), .B2(n20598), .ZN(
        n20592) );
  INV_X1 U23535 ( .A(n20592), .ZN(n20594) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20602), .B1(
        n21048), .B2(n20601), .ZN(n20593) );
  OAI211_X1 U23537 ( .C1(n21053), .C2(n20599), .A(n20594), .B(n20593), .ZN(
        P1_U3054) );
  OAI22_X1 U23538 ( .A1(n20599), .A2(n21059), .B1(n20729), .B2(n20598), .ZN(
        n20595) );
  INV_X1 U23539 ( .A(n20595), .ZN(n20597) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20602), .B1(
        n21054), .B2(n20601), .ZN(n20596) );
  OAI211_X1 U23541 ( .C1(n20966), .C2(n20643), .A(n20597), .B(n20596), .ZN(
        P1_U3055) );
  OAI22_X1 U23542 ( .A1(n20599), .A2(n21070), .B1(n20733), .B2(n20598), .ZN(
        n20600) );
  INV_X1 U23543 ( .A(n20600), .ZN(n20604) );
  AOI22_X1 U23544 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20602), .B1(
        n21061), .B2(n20601), .ZN(n20603) );
  OAI211_X1 U23545 ( .C1(n20974), .C2(n20643), .A(n20604), .B(n20603), .ZN(
        P1_U3056) );
  OR2_X1 U23546 ( .A1(n20874), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20637) );
  OAI22_X1 U23547 ( .A1(n20643), .A2(n21023), .B1(n20698), .B2(n20637), .ZN(
        n20605) );
  INV_X1 U23548 ( .A(n20605), .ZN(n20618) );
  AND2_X1 U23549 ( .A1(n20607), .A2(n20606), .ZN(n21008) );
  INV_X1 U23550 ( .A(n20637), .ZN(n20608) );
  AOI21_X1 U23551 ( .B1(n20609), .B2(n21008), .A(n20608), .ZN(n20616) );
  OR2_X1 U23552 ( .A1(n20610), .A2(n20877), .ZN(n20611) );
  AOI22_X1 U23553 ( .A1(n20616), .A2(n20613), .B1(n21010), .B2(n20614), .ZN(
        n20612) );
  NAND2_X1 U23554 ( .A1(n21018), .A2(n20612), .ZN(n20640) );
  INV_X1 U23555 ( .A(n20613), .ZN(n20615) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20640), .B1(
        n21013), .B2(n20639), .ZN(n20617) );
  OAI211_X1 U23557 ( .C1(n20942), .C2(n20663), .A(n20618), .B(n20617), .ZN(
        P1_U3057) );
  OAI22_X1 U23558 ( .A1(n20663), .A2(n20946), .B1(n20709), .B2(n20637), .ZN(
        n20619) );
  INV_X1 U23559 ( .A(n20619), .ZN(n20621) );
  AOI22_X1 U23560 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20640), .B1(
        n21024), .B2(n20639), .ZN(n20620) );
  OAI211_X1 U23561 ( .C1(n21029), .C2(n20643), .A(n20621), .B(n20620), .ZN(
        P1_U3058) );
  OAI22_X1 U23562 ( .A1(n20663), .A2(n20950), .B1(n20713), .B2(n20637), .ZN(
        n20622) );
  INV_X1 U23563 ( .A(n20622), .ZN(n20624) );
  AOI22_X1 U23564 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20640), .B1(
        n21030), .B2(n20639), .ZN(n20623) );
  OAI211_X1 U23565 ( .C1(n21035), .C2(n20643), .A(n20624), .B(n20623), .ZN(
        P1_U3059) );
  OAI22_X1 U23566 ( .A1(n20663), .A2(n20954), .B1(n20717), .B2(n20637), .ZN(
        n20625) );
  INV_X1 U23567 ( .A(n20625), .ZN(n20627) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20640), .B1(
        n21036), .B2(n20639), .ZN(n20626) );
  OAI211_X1 U23569 ( .C1(n21041), .C2(n20643), .A(n20627), .B(n20626), .ZN(
        P1_U3060) );
  OAI22_X1 U23570 ( .A1(n20643), .A2(n21047), .B1(n20721), .B2(n20637), .ZN(
        n20628) );
  INV_X1 U23571 ( .A(n20628), .ZN(n20630) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20640), .B1(
        n21042), .B2(n20639), .ZN(n20629) );
  OAI211_X1 U23573 ( .C1(n20958), .C2(n20663), .A(n20630), .B(n20629), .ZN(
        P1_U3061) );
  OAI22_X1 U23574 ( .A1(n20663), .A2(n20962), .B1(n20725), .B2(n20637), .ZN(
        n20631) );
  INV_X1 U23575 ( .A(n20631), .ZN(n20633) );
  AOI22_X1 U23576 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20640), .B1(
        n21048), .B2(n20639), .ZN(n20632) );
  OAI211_X1 U23577 ( .C1(n21053), .C2(n20643), .A(n20633), .B(n20632), .ZN(
        P1_U3062) );
  OAI22_X1 U23578 ( .A1(n20663), .A2(n20966), .B1(n20729), .B2(n20637), .ZN(
        n20634) );
  INV_X1 U23579 ( .A(n20634), .ZN(n20636) );
  AOI22_X1 U23580 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20640), .B1(
        n21054), .B2(n20639), .ZN(n20635) );
  OAI211_X1 U23581 ( .C1(n21059), .C2(n20643), .A(n20636), .B(n20635), .ZN(
        P1_U3063) );
  OAI22_X1 U23582 ( .A1(n20663), .A2(n20974), .B1(n20733), .B2(n20637), .ZN(
        n20638) );
  INV_X1 U23583 ( .A(n20638), .ZN(n20642) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20640), .B1(
        n21061), .B2(n20639), .ZN(n20641) );
  OAI211_X1 U23585 ( .C1(n21070), .C2(n20643), .A(n20642), .B(n20641), .ZN(
        P1_U3064) );
  NAND3_X1 U23586 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20873), .A3(
        n20901), .ZN(n20672) );
  NOR2_X1 U23587 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20672), .ZN(
        n20667) );
  OR2_X1 U23588 ( .A1(n13452), .A2(n20644), .ZN(n20648) );
  NAND3_X1 U23589 ( .A1(n20742), .A2(n20934), .A3(n13484), .ZN(n20645) );
  AOI22_X1 U23590 ( .A1(n21014), .A2(n20667), .B1(n21013), .B2(n20666), .ZN(
        n20652) );
  OAI21_X1 U23591 ( .B1(n20668), .B2(n20688), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20647) );
  OAI21_X1 U23592 ( .B1(n20981), .B2(n20648), .A(n20647), .ZN(n20650) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20669), .B1(
        n20688), .B2(n21020), .ZN(n20651) );
  OAI211_X1 U23594 ( .C1(n21023), .C2(n20663), .A(n20652), .B(n20651), .ZN(
        P1_U3065) );
  AOI22_X1 U23595 ( .A1(n21025), .A2(n20667), .B1(n21024), .B2(n20666), .ZN(
        n20654) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20943), .ZN(n20653) );
  OAI211_X1 U23597 ( .C1(n20946), .C2(n20697), .A(n20654), .B(n20653), .ZN(
        P1_U3066) );
  AOI22_X1 U23598 ( .A1(n21031), .A2(n20667), .B1(n21030), .B2(n20666), .ZN(
        n20656) );
  AOI22_X1 U23599 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20947), .ZN(n20655) );
  OAI211_X1 U23600 ( .C1(n20950), .C2(n20697), .A(n20656), .B(n20655), .ZN(
        P1_U3067) );
  AOI22_X1 U23601 ( .A1(n21037), .A2(n20667), .B1(n21036), .B2(n20666), .ZN(
        n20658) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20951), .ZN(n20657) );
  OAI211_X1 U23603 ( .C1(n20954), .C2(n20697), .A(n20658), .B(n20657), .ZN(
        P1_U3068) );
  AOI22_X1 U23604 ( .A1(n21043), .A2(n20667), .B1(n21042), .B2(n20666), .ZN(
        n20660) );
  INV_X1 U23605 ( .A(n20958), .ZN(n21044) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20669), .B1(
        n20688), .B2(n21044), .ZN(n20659) );
  OAI211_X1 U23607 ( .C1(n21047), .C2(n20663), .A(n20660), .B(n20659), .ZN(
        P1_U3069) );
  AOI22_X1 U23608 ( .A1(n21049), .A2(n20667), .B1(n21048), .B2(n20666), .ZN(
        n20662) );
  AOI22_X1 U23609 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20669), .B1(
        n20688), .B2(n21050), .ZN(n20661) );
  OAI211_X1 U23610 ( .C1(n21053), .C2(n20663), .A(n20662), .B(n20661), .ZN(
        P1_U3070) );
  AOI22_X1 U23611 ( .A1(n21055), .A2(n20667), .B1(n21054), .B2(n20666), .ZN(
        n20665) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20963), .ZN(n20664) );
  OAI211_X1 U23613 ( .C1(n20966), .C2(n20697), .A(n20665), .B(n20664), .ZN(
        P1_U3071) );
  AOI22_X1 U23614 ( .A1(n21063), .A2(n20667), .B1(n21061), .B2(n20666), .ZN(
        n20671) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20969), .ZN(n20670) );
  OAI211_X1 U23616 ( .C1(n20974), .C2(n20697), .A(n20671), .B(n20670), .ZN(
        P1_U3072) );
  NOR2_X1 U23617 ( .A1(n20933), .A2(n20672), .ZN(n20692) );
  AOI21_X1 U23618 ( .B1(n20742), .B2(n20803), .A(n20692), .ZN(n20673) );
  OAI22_X1 U23619 ( .A1(n20673), .A2(n21010), .B1(n20672), .B2(n21074), .ZN(
        n20691) );
  AOI22_X1 U23620 ( .A1(n21014), .A2(n20692), .B1(n21013), .B2(n20691), .ZN(
        n20677) );
  INV_X1 U23621 ( .A(n20672), .ZN(n20675) );
  OAI21_X1 U23622 ( .B1(n20750), .B2(n20806), .A(n20673), .ZN(n20674) );
  OAI221_X1 U23623 ( .B1(n20934), .B2(n20675), .C1(n21010), .C2(n20674), .A(
        n21018), .ZN(n20694) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20694), .B1(
        n20693), .B2(n21020), .ZN(n20676) );
  OAI211_X1 U23625 ( .C1(n21023), .C2(n20697), .A(n20677), .B(n20676), .ZN(
        P1_U3073) );
  AOI22_X1 U23626 ( .A1(n21025), .A2(n20692), .B1(n21024), .B2(n20691), .ZN(
        n20679) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20694), .B1(
        n20688), .B2(n20943), .ZN(n20678) );
  OAI211_X1 U23628 ( .C1(n20946), .C2(n20735), .A(n20679), .B(n20678), .ZN(
        P1_U3074) );
  AOI22_X1 U23629 ( .A1(n21031), .A2(n20692), .B1(n21030), .B2(n20691), .ZN(
        n20681) );
  INV_X1 U23630 ( .A(n20950), .ZN(n21032) );
  AOI22_X1 U23631 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20694), .B1(
        n20693), .B2(n21032), .ZN(n20680) );
  OAI211_X1 U23632 ( .C1(n21035), .C2(n20697), .A(n20681), .B(n20680), .ZN(
        P1_U3075) );
  AOI22_X1 U23633 ( .A1(n21037), .A2(n20692), .B1(n21036), .B2(n20691), .ZN(
        n20683) );
  AOI22_X1 U23634 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20694), .B1(
        n20693), .B2(n21038), .ZN(n20682) );
  OAI211_X1 U23635 ( .C1(n21041), .C2(n20697), .A(n20683), .B(n20682), .ZN(
        P1_U3076) );
  AOI22_X1 U23636 ( .A1(n21043), .A2(n20692), .B1(n21042), .B2(n20691), .ZN(
        n20685) );
  AOI22_X1 U23637 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20694), .B1(
        n20688), .B2(n20955), .ZN(n20684) );
  OAI211_X1 U23638 ( .C1(n20958), .C2(n20735), .A(n20685), .B(n20684), .ZN(
        P1_U3077) );
  AOI22_X1 U23639 ( .A1(n21049), .A2(n20692), .B1(n21048), .B2(n20691), .ZN(
        n20687) );
  AOI22_X1 U23640 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20694), .B1(
        n20693), .B2(n21050), .ZN(n20686) );
  OAI211_X1 U23641 ( .C1(n21053), .C2(n20697), .A(n20687), .B(n20686), .ZN(
        P1_U3078) );
  AOI22_X1 U23642 ( .A1(n21055), .A2(n20692), .B1(n21054), .B2(n20691), .ZN(
        n20690) );
  AOI22_X1 U23643 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20694), .B1(
        n20688), .B2(n20963), .ZN(n20689) );
  OAI211_X1 U23644 ( .C1(n20966), .C2(n20735), .A(n20690), .B(n20689), .ZN(
        P1_U3079) );
  AOI22_X1 U23645 ( .A1(n21063), .A2(n20692), .B1(n21061), .B2(n20691), .ZN(
        n20696) );
  INV_X1 U23646 ( .A(n20974), .ZN(n21064) );
  AOI22_X1 U23647 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20694), .B1(
        n20693), .B2(n21064), .ZN(n20695) );
  OAI211_X1 U23648 ( .C1(n21070), .C2(n20697), .A(n20696), .B(n20695), .ZN(
        P1_U3080) );
  INV_X1 U23649 ( .A(n20748), .ZN(n20743) );
  OAI22_X1 U23650 ( .A1(n20765), .A2(n20942), .B1(n20698), .B2(n20734), .ZN(
        n20699) );
  INV_X1 U23651 ( .A(n20699), .ZN(n20708) );
  NAND3_X1 U23652 ( .A1(n20765), .A2(n20735), .A3(n20934), .ZN(n20700) );
  NAND2_X1 U23653 ( .A1(n20700), .A2(n20902), .ZN(n20703) );
  NAND2_X1 U23654 ( .A1(n20742), .A2(n20981), .ZN(n20705) );
  AOI22_X1 U23655 ( .A1(n20703), .A2(n20705), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20734), .ZN(n20702) );
  NAND3_X1 U23656 ( .A1(n20985), .A2(n20702), .A3(n20701), .ZN(n20738) );
  INV_X1 U23657 ( .A(n20703), .ZN(n20706) );
  AOI22_X1 U23658 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20738), .B1(
        n21013), .B2(n20737), .ZN(n20707) );
  OAI211_X1 U23659 ( .C1(n21023), .C2(n20735), .A(n20708), .B(n20707), .ZN(
        P1_U3081) );
  OAI22_X1 U23660 ( .A1(n20735), .A2(n21029), .B1(n20734), .B2(n20709), .ZN(
        n20710) );
  INV_X1 U23661 ( .A(n20710), .ZN(n20712) );
  AOI22_X1 U23662 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20738), .B1(
        n21024), .B2(n20737), .ZN(n20711) );
  OAI211_X1 U23663 ( .C1(n20946), .C2(n20765), .A(n20712), .B(n20711), .ZN(
        P1_U3082) );
  OAI22_X1 U23664 ( .A1(n20765), .A2(n20950), .B1(n20734), .B2(n20713), .ZN(
        n20714) );
  INV_X1 U23665 ( .A(n20714), .ZN(n20716) );
  AOI22_X1 U23666 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20738), .B1(
        n21030), .B2(n20737), .ZN(n20715) );
  OAI211_X1 U23667 ( .C1(n21035), .C2(n20735), .A(n20716), .B(n20715), .ZN(
        P1_U3083) );
  OAI22_X1 U23668 ( .A1(n20765), .A2(n20954), .B1(n20734), .B2(n20717), .ZN(
        n20718) );
  INV_X1 U23669 ( .A(n20718), .ZN(n20720) );
  AOI22_X1 U23670 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20738), .B1(
        n21036), .B2(n20737), .ZN(n20719) );
  OAI211_X1 U23671 ( .C1(n21041), .C2(n20735), .A(n20720), .B(n20719), .ZN(
        P1_U3084) );
  OAI22_X1 U23672 ( .A1(n20735), .A2(n21047), .B1(n20734), .B2(n20721), .ZN(
        n20722) );
  INV_X1 U23673 ( .A(n20722), .ZN(n20724) );
  AOI22_X1 U23674 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20738), .B1(
        n21042), .B2(n20737), .ZN(n20723) );
  OAI211_X1 U23675 ( .C1(n20958), .C2(n20765), .A(n20724), .B(n20723), .ZN(
        P1_U3085) );
  OAI22_X1 U23676 ( .A1(n20735), .A2(n21053), .B1(n20734), .B2(n20725), .ZN(
        n20726) );
  INV_X1 U23677 ( .A(n20726), .ZN(n20728) );
  AOI22_X1 U23678 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20738), .B1(
        n21048), .B2(n20737), .ZN(n20727) );
  OAI211_X1 U23679 ( .C1(n20962), .C2(n20765), .A(n20728), .B(n20727), .ZN(
        P1_U3086) );
  OAI22_X1 U23680 ( .A1(n20765), .A2(n20966), .B1(n20734), .B2(n20729), .ZN(
        n20730) );
  INV_X1 U23681 ( .A(n20730), .ZN(n20732) );
  AOI22_X1 U23682 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20738), .B1(
        n21054), .B2(n20737), .ZN(n20731) );
  OAI211_X1 U23683 ( .C1(n21059), .C2(n20735), .A(n20732), .B(n20731), .ZN(
        P1_U3087) );
  OAI22_X1 U23684 ( .A1(n20735), .A2(n21070), .B1(n20734), .B2(n20733), .ZN(
        n20736) );
  INV_X1 U23685 ( .A(n20736), .ZN(n20740) );
  AOI22_X1 U23686 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20738), .B1(
        n21061), .B2(n20737), .ZN(n20739) );
  OAI211_X1 U23687 ( .C1(n20974), .C2(n20765), .A(n20740), .B(n20739), .ZN(
        P1_U3088) );
  INV_X1 U23688 ( .A(n20741), .ZN(n20767) );
  AOI21_X1 U23689 ( .B1(n20742), .B2(n21008), .A(n20767), .ZN(n20745) );
  OAI22_X1 U23690 ( .A1(n20745), .A2(n21010), .B1(n21074), .B2(n20743), .ZN(
        n20766) );
  AOI22_X1 U23691 ( .A1(n21014), .A2(n20767), .B1(n21013), .B2(n20766), .ZN(
        n20752) );
  INV_X1 U23692 ( .A(n20744), .ZN(n20746) );
  NAND2_X1 U23693 ( .A1(n20746), .A2(n20745), .ZN(n20747) );
  OAI221_X1 U23694 ( .B1(n20934), .B2(n20748), .C1(n21010), .C2(n20747), .A(
        n21018), .ZN(n20769) );
  AOI22_X1 U23695 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20769), .B1(
        n20799), .B2(n21020), .ZN(n20751) );
  OAI211_X1 U23696 ( .C1(n21023), .C2(n20765), .A(n20752), .B(n20751), .ZN(
        P1_U3089) );
  AOI22_X1 U23697 ( .A1(n21025), .A2(n20767), .B1(n21024), .B2(n20766), .ZN(
        n20754) );
  INV_X1 U23698 ( .A(n20765), .ZN(n20768) );
  AOI22_X1 U23699 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20769), .B1(
        n20768), .B2(n20943), .ZN(n20753) );
  OAI211_X1 U23700 ( .C1(n20946), .C2(n20772), .A(n20754), .B(n20753), .ZN(
        P1_U3090) );
  AOI22_X1 U23701 ( .A1(n21031), .A2(n20767), .B1(n21030), .B2(n20766), .ZN(
        n20756) );
  AOI22_X1 U23702 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20769), .B1(
        n20799), .B2(n21032), .ZN(n20755) );
  OAI211_X1 U23703 ( .C1(n21035), .C2(n20765), .A(n20756), .B(n20755), .ZN(
        P1_U3091) );
  AOI22_X1 U23704 ( .A1(n21037), .A2(n20767), .B1(n21036), .B2(n20766), .ZN(
        n20758) );
  AOI22_X1 U23705 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20769), .B1(
        n20799), .B2(n21038), .ZN(n20757) );
  OAI211_X1 U23706 ( .C1(n21041), .C2(n20765), .A(n20758), .B(n20757), .ZN(
        P1_U3092) );
  AOI22_X1 U23707 ( .A1(n21043), .A2(n20767), .B1(n21042), .B2(n20766), .ZN(
        n20760) );
  AOI22_X1 U23708 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20769), .B1(
        n20799), .B2(n21044), .ZN(n20759) );
  OAI211_X1 U23709 ( .C1(n21047), .C2(n20765), .A(n20760), .B(n20759), .ZN(
        P1_U3093) );
  AOI22_X1 U23710 ( .A1(n21049), .A2(n20767), .B1(n21048), .B2(n20766), .ZN(
        n20762) );
  AOI22_X1 U23711 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20769), .B1(
        n20799), .B2(n21050), .ZN(n20761) );
  OAI211_X1 U23712 ( .C1(n21053), .C2(n20765), .A(n20762), .B(n20761), .ZN(
        P1_U3094) );
  AOI22_X1 U23713 ( .A1(n21055), .A2(n20767), .B1(n21054), .B2(n20766), .ZN(
        n20764) );
  AOI22_X1 U23714 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20769), .B1(
        n20799), .B2(n21056), .ZN(n20763) );
  OAI211_X1 U23715 ( .C1(n21059), .C2(n20765), .A(n20764), .B(n20763), .ZN(
        P1_U3095) );
  AOI22_X1 U23716 ( .A1(n21063), .A2(n20767), .B1(n21061), .B2(n20766), .ZN(
        n20771) );
  AOI22_X1 U23717 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20769), .B1(
        n20768), .B2(n20969), .ZN(n20770) );
  OAI211_X1 U23718 ( .C1(n20974), .C2(n20772), .A(n20771), .B(n20770), .ZN(
        P1_U3096) );
  INV_X1 U23719 ( .A(n20900), .ZN(n20773) );
  NAND3_X1 U23720 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20836), .A3(
        n20901), .ZN(n20804) );
  NOR2_X1 U23721 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20804), .ZN(
        n20798) );
  AND2_X1 U23722 ( .A1(n20774), .A2(n13452), .ZN(n20875) );
  AOI21_X1 U23723 ( .B1(n20875), .B2(n13484), .A(n20798), .ZN(n20779) );
  INV_X1 U23724 ( .A(n20775), .ZN(n20776) );
  NAND2_X1 U23725 ( .A1(n20776), .A2(n20833), .ZN(n20909) );
  OAI22_X1 U23726 ( .A1(n20779), .A2(n21010), .B1(n20909), .B2(n20777), .ZN(
        n20797) );
  AOI22_X1 U23727 ( .A1(n21014), .A2(n20798), .B1(n20797), .B2(n21013), .ZN(
        n20784) );
  INV_X1 U23728 ( .A(n20829), .ZN(n20778) );
  OAI21_X1 U23729 ( .B1(n20778), .B2(n20799), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20780) );
  NAND2_X1 U23730 ( .A1(n20780), .A2(n20779), .ZN(n20781) );
  AOI22_X1 U23731 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20800), .B1(
        n20799), .B2(n20939), .ZN(n20783) );
  OAI211_X1 U23732 ( .C1(n20942), .C2(n20829), .A(n20784), .B(n20783), .ZN(
        P1_U3097) );
  AOI22_X1 U23733 ( .A1(n21025), .A2(n20798), .B1(n20797), .B2(n21024), .ZN(
        n20786) );
  AOI22_X1 U23734 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20800), .B1(
        n20799), .B2(n20943), .ZN(n20785) );
  OAI211_X1 U23735 ( .C1(n20946), .C2(n20829), .A(n20786), .B(n20785), .ZN(
        P1_U3098) );
  AOI22_X1 U23736 ( .A1(n21031), .A2(n20798), .B1(n20797), .B2(n21030), .ZN(
        n20788) );
  AOI22_X1 U23737 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20800), .B1(
        n20799), .B2(n20947), .ZN(n20787) );
  OAI211_X1 U23738 ( .C1(n20950), .C2(n20829), .A(n20788), .B(n20787), .ZN(
        P1_U3099) );
  AOI22_X1 U23739 ( .A1(n21037), .A2(n20798), .B1(n20797), .B2(n21036), .ZN(
        n20790) );
  AOI22_X1 U23740 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20800), .B1(
        n20799), .B2(n20951), .ZN(n20789) );
  OAI211_X1 U23741 ( .C1(n20954), .C2(n20829), .A(n20790), .B(n20789), .ZN(
        P1_U3100) );
  AOI22_X1 U23742 ( .A1(n21043), .A2(n20798), .B1(n20797), .B2(n21042), .ZN(
        n20792) );
  AOI22_X1 U23743 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20800), .B1(
        n20799), .B2(n20955), .ZN(n20791) );
  OAI211_X1 U23744 ( .C1(n20958), .C2(n20829), .A(n20792), .B(n20791), .ZN(
        P1_U3101) );
  AOI22_X1 U23745 ( .A1(n21049), .A2(n20798), .B1(n20797), .B2(n21048), .ZN(
        n20794) );
  AOI22_X1 U23746 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20800), .B1(
        n20799), .B2(n20959), .ZN(n20793) );
  OAI211_X1 U23747 ( .C1(n20962), .C2(n20829), .A(n20794), .B(n20793), .ZN(
        P1_U3102) );
  AOI22_X1 U23748 ( .A1(n21055), .A2(n20798), .B1(n20797), .B2(n21054), .ZN(
        n20796) );
  AOI22_X1 U23749 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20800), .B1(
        n20799), .B2(n20963), .ZN(n20795) );
  OAI211_X1 U23750 ( .C1(n20966), .C2(n20829), .A(n20796), .B(n20795), .ZN(
        P1_U3103) );
  AOI22_X1 U23751 ( .A1(n21063), .A2(n20798), .B1(n20797), .B2(n21061), .ZN(
        n20802) );
  AOI22_X1 U23752 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20800), .B1(
        n20799), .B2(n20969), .ZN(n20801) );
  OAI211_X1 U23753 ( .C1(n20974), .C2(n20829), .A(n20802), .B(n20801), .ZN(
        P1_U3104) );
  NOR2_X1 U23754 ( .A1(n20933), .A2(n20804), .ZN(n20825) );
  AOI21_X1 U23755 ( .B1(n20875), .B2(n20803), .A(n20825), .ZN(n20805) );
  OAI22_X1 U23756 ( .A1(n20805), .A2(n21010), .B1(n20804), .B2(n21074), .ZN(
        n20824) );
  AOI22_X1 U23757 ( .A1(n21014), .A2(n20825), .B1(n20824), .B2(n21013), .ZN(
        n20811) );
  INV_X1 U23758 ( .A(n20804), .ZN(n20808) );
  INV_X1 U23759 ( .A(n20872), .ZN(n20879) );
  OAI21_X1 U23760 ( .B1(n20879), .B2(n20806), .A(n20805), .ZN(n20807) );
  OAI221_X1 U23761 ( .B1(n20934), .B2(n20808), .C1(n21010), .C2(n20807), .A(
        n21018), .ZN(n20826) );
  AOI22_X1 U23762 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20826), .B1(
        n20865), .B2(n21020), .ZN(n20810) );
  OAI211_X1 U23763 ( .C1(n21023), .C2(n20829), .A(n20811), .B(n20810), .ZN(
        P1_U3105) );
  AOI22_X1 U23764 ( .A1(n21025), .A2(n20825), .B1(n20824), .B2(n21024), .ZN(
        n20813) );
  AOI22_X1 U23765 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20826), .B1(
        n20865), .B2(n21026), .ZN(n20812) );
  OAI211_X1 U23766 ( .C1(n21029), .C2(n20829), .A(n20813), .B(n20812), .ZN(
        P1_U3106) );
  AOI22_X1 U23767 ( .A1(n21031), .A2(n20825), .B1(n20824), .B2(n21030), .ZN(
        n20815) );
  AOI22_X1 U23768 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20826), .B1(
        n20865), .B2(n21032), .ZN(n20814) );
  OAI211_X1 U23769 ( .C1(n21035), .C2(n20829), .A(n20815), .B(n20814), .ZN(
        P1_U3107) );
  AOI22_X1 U23770 ( .A1(n21037), .A2(n20825), .B1(n20824), .B2(n21036), .ZN(
        n20817) );
  AOI22_X1 U23771 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20826), .B1(
        n20865), .B2(n21038), .ZN(n20816) );
  OAI211_X1 U23772 ( .C1(n21041), .C2(n20829), .A(n20817), .B(n20816), .ZN(
        P1_U3108) );
  AOI22_X1 U23773 ( .A1(n21043), .A2(n20825), .B1(n20824), .B2(n21042), .ZN(
        n20819) );
  AOI22_X1 U23774 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20826), .B1(
        n20865), .B2(n21044), .ZN(n20818) );
  OAI211_X1 U23775 ( .C1(n21047), .C2(n20829), .A(n20819), .B(n20818), .ZN(
        P1_U3109) );
  AOI22_X1 U23776 ( .A1(n21049), .A2(n20825), .B1(n20824), .B2(n21048), .ZN(
        n20821) );
  AOI22_X1 U23777 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20826), .B1(
        n20865), .B2(n21050), .ZN(n20820) );
  OAI211_X1 U23778 ( .C1(n21053), .C2(n20829), .A(n20821), .B(n20820), .ZN(
        P1_U3110) );
  AOI22_X1 U23779 ( .A1(n21055), .A2(n20825), .B1(n20824), .B2(n21054), .ZN(
        n20823) );
  AOI22_X1 U23780 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20826), .B1(
        n20865), .B2(n21056), .ZN(n20822) );
  OAI211_X1 U23781 ( .C1(n21059), .C2(n20829), .A(n20823), .B(n20822), .ZN(
        P1_U3111) );
  AOI22_X1 U23782 ( .A1(n21063), .A2(n20825), .B1(n20824), .B2(n21061), .ZN(
        n20828) );
  AOI22_X1 U23783 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20826), .B1(
        n20865), .B2(n21064), .ZN(n20827) );
  OAI211_X1 U23784 ( .C1(n21070), .C2(n20829), .A(n20828), .B(n20827), .ZN(
        P1_U3112) );
  INV_X1 U23785 ( .A(n20865), .ZN(n20830) );
  NAND2_X1 U23786 ( .A1(n20830), .A2(n20934), .ZN(n20832) );
  INV_X1 U23787 ( .A(n20831), .ZN(n20977) );
  OAI21_X1 U23788 ( .B1(n20832), .B2(n20896), .A(n20902), .ZN(n20840) );
  OR2_X1 U23789 ( .A1(n20833), .A2(n20873), .ZN(n20975) );
  INV_X1 U23790 ( .A(n20975), .ZN(n20835) );
  INV_X1 U23791 ( .A(n21013), .ZN(n20845) );
  NAND3_X1 U23792 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20836), .ZN(n20878) );
  NOR2_X1 U23793 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20878), .ZN(
        n20864) );
  AOI22_X1 U23794 ( .A1(n20865), .A2(n20939), .B1(n21014), .B2(n20864), .ZN(
        n20844) );
  INV_X1 U23795 ( .A(n20837), .ZN(n20839) );
  INV_X1 U23796 ( .A(n20864), .ZN(n20838) );
  AOI22_X1 U23797 ( .A1(n20840), .A2(n20839), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20838), .ZN(n20841) );
  NAND2_X1 U23798 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20975), .ZN(n20984) );
  NAND3_X1 U23799 ( .A1(n20842), .A2(n20841), .A3(n20984), .ZN(n20866) );
  AOI22_X1 U23800 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20866), .B1(
        n20896), .B2(n21020), .ZN(n20843) );
  OAI211_X1 U23801 ( .C1(n20870), .C2(n20845), .A(n20844), .B(n20843), .ZN(
        P1_U3113) );
  INV_X1 U23802 ( .A(n21024), .ZN(n20848) );
  AOI22_X1 U23803 ( .A1(n20896), .A2(n21026), .B1(n21025), .B2(n20864), .ZN(
        n20847) );
  AOI22_X1 U23804 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20866), .B1(
        n20865), .B2(n20943), .ZN(n20846) );
  OAI211_X1 U23805 ( .C1(n20870), .C2(n20848), .A(n20847), .B(n20846), .ZN(
        P1_U3114) );
  INV_X1 U23806 ( .A(n21030), .ZN(n20851) );
  AOI22_X1 U23807 ( .A1(n20896), .A2(n21032), .B1(n21031), .B2(n20864), .ZN(
        n20850) );
  AOI22_X1 U23808 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20866), .B1(
        n20865), .B2(n20947), .ZN(n20849) );
  OAI211_X1 U23809 ( .C1(n20870), .C2(n20851), .A(n20850), .B(n20849), .ZN(
        P1_U3115) );
  INV_X1 U23810 ( .A(n21036), .ZN(n20854) );
  AOI22_X1 U23811 ( .A1(n20865), .A2(n20951), .B1(n21037), .B2(n20864), .ZN(
        n20853) );
  AOI22_X1 U23812 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20866), .B1(
        n20896), .B2(n21038), .ZN(n20852) );
  OAI211_X1 U23813 ( .C1(n20870), .C2(n20854), .A(n20853), .B(n20852), .ZN(
        P1_U3116) );
  INV_X1 U23814 ( .A(n21042), .ZN(n20857) );
  AOI22_X1 U23815 ( .A1(n20865), .A2(n20955), .B1(n21043), .B2(n20864), .ZN(
        n20856) );
  AOI22_X1 U23816 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20866), .B1(
        n20896), .B2(n21044), .ZN(n20855) );
  OAI211_X1 U23817 ( .C1(n20870), .C2(n20857), .A(n20856), .B(n20855), .ZN(
        P1_U3117) );
  INV_X1 U23818 ( .A(n21048), .ZN(n20860) );
  AOI22_X1 U23819 ( .A1(n20896), .A2(n21050), .B1(n21049), .B2(n20864), .ZN(
        n20859) );
  AOI22_X1 U23820 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20866), .B1(
        n20865), .B2(n20959), .ZN(n20858) );
  OAI211_X1 U23821 ( .C1(n20870), .C2(n20860), .A(n20859), .B(n20858), .ZN(
        P1_U3118) );
  INV_X1 U23822 ( .A(n21054), .ZN(n20863) );
  AOI22_X1 U23823 ( .A1(n20865), .A2(n20963), .B1(n21055), .B2(n20864), .ZN(
        n20862) );
  AOI22_X1 U23824 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20866), .B1(
        n20896), .B2(n21056), .ZN(n20861) );
  OAI211_X1 U23825 ( .C1(n20870), .C2(n20863), .A(n20862), .B(n20861), .ZN(
        P1_U3119) );
  INV_X1 U23826 ( .A(n21061), .ZN(n20869) );
  AOI22_X1 U23827 ( .A1(n20865), .A2(n20969), .B1(n21063), .B2(n20864), .ZN(
        n20868) );
  AOI22_X1 U23828 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20866), .B1(
        n20896), .B2(n21064), .ZN(n20867) );
  OAI211_X1 U23829 ( .C1(n20870), .C2(n20869), .A(n20868), .B(n20867), .ZN(
        P1_U3120) );
  AOI21_X1 U23830 ( .B1(n20875), .B2(n21008), .A(n10553), .ZN(n20876) );
  OAI22_X1 U23831 ( .A1(n20876), .A2(n21010), .B1(n20878), .B2(n21074), .ZN(
        n20895) );
  AOI22_X1 U23832 ( .A1(n21014), .A2(n10553), .B1(n21013), .B2(n20895), .ZN(
        n20882) );
  OR2_X1 U23833 ( .A1(n20877), .A2(n21010), .ZN(n21016) );
  OAI21_X1 U23834 ( .B1(n20879), .B2(n21016), .A(n20878), .ZN(n20880) );
  NAND2_X1 U23835 ( .A1(n20880), .A2(n21018), .ZN(n20897) );
  AOI22_X1 U23836 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20897), .B1(
        n20896), .B2(n20939), .ZN(n20881) );
  OAI211_X1 U23837 ( .C1(n20942), .C2(n20931), .A(n20882), .B(n20881), .ZN(
        P1_U3121) );
  AOI22_X1 U23838 ( .A1(n21025), .A2(n10553), .B1(n21024), .B2(n20895), .ZN(
        n20884) );
  AOI22_X1 U23839 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20897), .B1(
        n20896), .B2(n20943), .ZN(n20883) );
  OAI211_X1 U23840 ( .C1(n20946), .C2(n20931), .A(n20884), .B(n20883), .ZN(
        P1_U3122) );
  AOI22_X1 U23841 ( .A1(n21031), .A2(n10553), .B1(n21030), .B2(n20895), .ZN(
        n20886) );
  AOI22_X1 U23842 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20897), .B1(
        n20896), .B2(n20947), .ZN(n20885) );
  OAI211_X1 U23843 ( .C1(n20950), .C2(n20931), .A(n20886), .B(n20885), .ZN(
        P1_U3123) );
  AOI22_X1 U23844 ( .A1(n21037), .A2(n10553), .B1(n21036), .B2(n20895), .ZN(
        n20888) );
  AOI22_X1 U23845 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20897), .B1(
        n20896), .B2(n20951), .ZN(n20887) );
  OAI211_X1 U23846 ( .C1(n20954), .C2(n20931), .A(n20888), .B(n20887), .ZN(
        P1_U3124) );
  AOI22_X1 U23847 ( .A1(n21043), .A2(n10553), .B1(n21042), .B2(n20895), .ZN(
        n20890) );
  AOI22_X1 U23848 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20897), .B1(
        n20896), .B2(n20955), .ZN(n20889) );
  OAI211_X1 U23849 ( .C1(n20958), .C2(n20931), .A(n20890), .B(n20889), .ZN(
        P1_U3125) );
  AOI22_X1 U23850 ( .A1(n21049), .A2(n10553), .B1(n21048), .B2(n20895), .ZN(
        n20892) );
  AOI22_X1 U23851 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20897), .B1(
        n20896), .B2(n20959), .ZN(n20891) );
  OAI211_X1 U23852 ( .C1(n20962), .C2(n20931), .A(n20892), .B(n20891), .ZN(
        P1_U3126) );
  AOI22_X1 U23853 ( .A1(n21055), .A2(n10553), .B1(n21054), .B2(n20895), .ZN(
        n20894) );
  AOI22_X1 U23854 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20897), .B1(
        n20896), .B2(n20963), .ZN(n20893) );
  OAI211_X1 U23855 ( .C1(n20966), .C2(n20931), .A(n20894), .B(n20893), .ZN(
        P1_U3127) );
  AOI22_X1 U23856 ( .A1(n21063), .A2(n10553), .B1(n21061), .B2(n20895), .ZN(
        n20899) );
  AOI22_X1 U23857 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20897), .B1(
        n20896), .B2(n20969), .ZN(n20898) );
  OAI211_X1 U23858 ( .C1(n20974), .C2(n20931), .A(n20899), .B(n20898), .ZN(
        P1_U3128) );
  NAND3_X1 U23859 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20901), .ZN(n20936) );
  NOR2_X1 U23860 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20936), .ZN(
        n20926) );
  AOI22_X1 U23861 ( .A1(n20970), .A2(n21020), .B1(n21014), .B2(n20926), .ZN(
        n20913) );
  INV_X1 U23862 ( .A(n20909), .ZN(n20907) );
  NAND2_X1 U23863 ( .A1(n20931), .A2(n20934), .ZN(n20903) );
  OAI21_X1 U23864 ( .B1(n20970), .B2(n20903), .A(n20902), .ZN(n20908) );
  NOR2_X1 U23865 ( .A1(n13452), .A2(n20904), .ZN(n20982) );
  NAND2_X1 U23866 ( .A1(n20982), .A2(n13484), .ZN(n20910) );
  INV_X1 U23867 ( .A(n20926), .ZN(n20905) );
  AOI22_X1 U23868 ( .A1(n20908), .A2(n20910), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20905), .ZN(n20906) );
  INV_X1 U23869 ( .A(n20908), .ZN(n20911) );
  AOI22_X1 U23870 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20928), .B1(
        n21013), .B2(n20927), .ZN(n20912) );
  OAI211_X1 U23871 ( .C1(n21023), .C2(n20931), .A(n20913), .B(n20912), .ZN(
        P1_U3129) );
  AOI22_X1 U23872 ( .A1(n20970), .A2(n21026), .B1(n21025), .B2(n20926), .ZN(
        n20915) );
  AOI22_X1 U23873 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20928), .B1(
        n21024), .B2(n20927), .ZN(n20914) );
  OAI211_X1 U23874 ( .C1(n21029), .C2(n20931), .A(n20915), .B(n20914), .ZN(
        P1_U3130) );
  AOI22_X1 U23875 ( .A1(n20970), .A2(n21032), .B1(n21031), .B2(n20926), .ZN(
        n20917) );
  AOI22_X1 U23876 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20928), .B1(
        n21030), .B2(n20927), .ZN(n20916) );
  OAI211_X1 U23877 ( .C1(n21035), .C2(n20931), .A(n20917), .B(n20916), .ZN(
        P1_U3131) );
  AOI22_X1 U23878 ( .A1(n20970), .A2(n21038), .B1(n21037), .B2(n20926), .ZN(
        n20919) );
  AOI22_X1 U23879 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20928), .B1(
        n21036), .B2(n20927), .ZN(n20918) );
  OAI211_X1 U23880 ( .C1(n21041), .C2(n20931), .A(n20919), .B(n20918), .ZN(
        P1_U3132) );
  AOI22_X1 U23881 ( .A1(n20970), .A2(n21044), .B1(n21043), .B2(n20926), .ZN(
        n20921) );
  AOI22_X1 U23882 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20928), .B1(
        n21042), .B2(n20927), .ZN(n20920) );
  OAI211_X1 U23883 ( .C1(n21047), .C2(n20931), .A(n20921), .B(n20920), .ZN(
        P1_U3133) );
  AOI22_X1 U23884 ( .A1(n20970), .A2(n21050), .B1(n21049), .B2(n20926), .ZN(
        n20923) );
  AOI22_X1 U23885 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20928), .B1(
        n21048), .B2(n20927), .ZN(n20922) );
  OAI211_X1 U23886 ( .C1(n21053), .C2(n20931), .A(n20923), .B(n20922), .ZN(
        P1_U3134) );
  AOI22_X1 U23887 ( .A1(n20970), .A2(n21056), .B1(n21055), .B2(n20926), .ZN(
        n20925) );
  AOI22_X1 U23888 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20928), .B1(
        n21054), .B2(n20927), .ZN(n20924) );
  OAI211_X1 U23889 ( .C1(n21059), .C2(n20931), .A(n20925), .B(n20924), .ZN(
        P1_U3135) );
  AOI22_X1 U23890 ( .A1(n20970), .A2(n21064), .B1(n21063), .B2(n20926), .ZN(
        n20930) );
  AOI22_X1 U23891 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20928), .B1(
        n21061), .B2(n20927), .ZN(n20929) );
  OAI211_X1 U23892 ( .C1(n21070), .C2(n20931), .A(n20930), .B(n20929), .ZN(
        P1_U3136) );
  NOR2_X1 U23893 ( .A1(n20933), .A2(n20936), .ZN(n20968) );
  NAND2_X1 U23894 ( .A1(n20982), .A2(n20934), .ZN(n21012) );
  INV_X1 U23895 ( .A(n20968), .ZN(n20935) );
  OAI222_X1 U23896 ( .A1(n21012), .A2(n20541), .B1(n21074), .B2(n20936), .C1(
        n21010), .C2(n20935), .ZN(n20967) );
  AOI22_X1 U23897 ( .A1(n21014), .A2(n20968), .B1(n21013), .B2(n20967), .ZN(
        n20941) );
  INV_X1 U23898 ( .A(n20936), .ZN(n20938) );
  AOI22_X1 U23899 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20971), .B1(
        n20970), .B2(n20939), .ZN(n20940) );
  OAI211_X1 U23900 ( .C1(n20942), .C2(n21007), .A(n20941), .B(n20940), .ZN(
        P1_U3137) );
  AOI22_X1 U23901 ( .A1(n21025), .A2(n20968), .B1(n21024), .B2(n20967), .ZN(
        n20945) );
  AOI22_X1 U23902 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20971), .B1(
        n20970), .B2(n20943), .ZN(n20944) );
  OAI211_X1 U23903 ( .C1(n20946), .C2(n21007), .A(n20945), .B(n20944), .ZN(
        P1_U3138) );
  AOI22_X1 U23904 ( .A1(n21031), .A2(n20968), .B1(n21030), .B2(n20967), .ZN(
        n20949) );
  AOI22_X1 U23905 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20971), .B1(
        n20970), .B2(n20947), .ZN(n20948) );
  OAI211_X1 U23906 ( .C1(n20950), .C2(n21007), .A(n20949), .B(n20948), .ZN(
        P1_U3139) );
  AOI22_X1 U23907 ( .A1(n21037), .A2(n20968), .B1(n21036), .B2(n20967), .ZN(
        n20953) );
  AOI22_X1 U23908 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20971), .B1(
        n20970), .B2(n20951), .ZN(n20952) );
  OAI211_X1 U23909 ( .C1(n20954), .C2(n21007), .A(n20953), .B(n20952), .ZN(
        P1_U3140) );
  AOI22_X1 U23910 ( .A1(n21043), .A2(n20968), .B1(n21042), .B2(n20967), .ZN(
        n20957) );
  AOI22_X1 U23911 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20971), .B1(
        n20970), .B2(n20955), .ZN(n20956) );
  OAI211_X1 U23912 ( .C1(n20958), .C2(n21007), .A(n20957), .B(n20956), .ZN(
        P1_U3141) );
  AOI22_X1 U23913 ( .A1(n21049), .A2(n20968), .B1(n21048), .B2(n20967), .ZN(
        n20961) );
  AOI22_X1 U23914 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20971), .B1(
        n20970), .B2(n20959), .ZN(n20960) );
  OAI211_X1 U23915 ( .C1(n20962), .C2(n21007), .A(n20961), .B(n20960), .ZN(
        P1_U3142) );
  AOI22_X1 U23916 ( .A1(n21055), .A2(n20968), .B1(n21054), .B2(n20967), .ZN(
        n20965) );
  AOI22_X1 U23917 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20971), .B1(
        n20970), .B2(n20963), .ZN(n20964) );
  OAI211_X1 U23918 ( .C1(n20966), .C2(n21007), .A(n20965), .B(n20964), .ZN(
        P1_U3143) );
  AOI22_X1 U23919 ( .A1(n21063), .A2(n20968), .B1(n21061), .B2(n20967), .ZN(
        n20973) );
  AOI22_X1 U23920 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20971), .B1(
        n20970), .B2(n20969), .ZN(n20972) );
  OAI211_X1 U23921 ( .C1(n20974), .C2(n21007), .A(n20973), .B(n20972), .ZN(
        P1_U3144) );
  NOR2_X1 U23922 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21015), .ZN(
        n21002) );
  OAI22_X1 U23923 ( .A1(n21012), .A2(n13484), .B1(n20976), .B2(n20975), .ZN(
        n21001) );
  AOI22_X1 U23924 ( .A1(n21014), .A2(n21002), .B1(n21013), .B2(n21001), .ZN(
        n20988) );
  AOI21_X1 U23925 ( .B1(n21069), .B2(n21007), .A(n20979), .ZN(n20980) );
  AOI21_X1 U23926 ( .B1(n20982), .B2(n20981), .A(n20980), .ZN(n20983) );
  NOR2_X1 U23927 ( .A1(n20983), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20986) );
  AOI22_X1 U23928 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n21004), .B1(
        n21003), .B2(n21020), .ZN(n20987) );
  OAI211_X1 U23929 ( .C1(n21023), .C2(n21007), .A(n20988), .B(n20987), .ZN(
        P1_U3145) );
  AOI22_X1 U23930 ( .A1(n21025), .A2(n21002), .B1(n21024), .B2(n21001), .ZN(
        n20990) );
  AOI22_X1 U23931 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21004), .B1(
        n21003), .B2(n21026), .ZN(n20989) );
  OAI211_X1 U23932 ( .C1(n21029), .C2(n21007), .A(n20990), .B(n20989), .ZN(
        P1_U3146) );
  AOI22_X1 U23933 ( .A1(n21031), .A2(n21002), .B1(n21030), .B2(n21001), .ZN(
        n20992) );
  AOI22_X1 U23934 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n21004), .B1(
        n21003), .B2(n21032), .ZN(n20991) );
  OAI211_X1 U23935 ( .C1(n21035), .C2(n21007), .A(n20992), .B(n20991), .ZN(
        P1_U3147) );
  AOI22_X1 U23936 ( .A1(n21037), .A2(n21002), .B1(n21036), .B2(n21001), .ZN(
        n20994) );
  AOI22_X1 U23937 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n21004), .B1(
        n21003), .B2(n21038), .ZN(n20993) );
  OAI211_X1 U23938 ( .C1(n21041), .C2(n21007), .A(n20994), .B(n20993), .ZN(
        P1_U3148) );
  AOI22_X1 U23939 ( .A1(n21043), .A2(n21002), .B1(n21042), .B2(n21001), .ZN(
        n20996) );
  AOI22_X1 U23940 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n21004), .B1(
        n21003), .B2(n21044), .ZN(n20995) );
  OAI211_X1 U23941 ( .C1(n21047), .C2(n21007), .A(n20996), .B(n20995), .ZN(
        P1_U3149) );
  AOI22_X1 U23942 ( .A1(n21049), .A2(n21002), .B1(n21048), .B2(n21001), .ZN(
        n20998) );
  AOI22_X1 U23943 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n21004), .B1(
        n21003), .B2(n21050), .ZN(n20997) );
  OAI211_X1 U23944 ( .C1(n21053), .C2(n21007), .A(n20998), .B(n20997), .ZN(
        P1_U3150) );
  AOI22_X1 U23945 ( .A1(n21055), .A2(n21002), .B1(n21054), .B2(n21001), .ZN(
        n21000) );
  AOI22_X1 U23946 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n21004), .B1(
        n21003), .B2(n21056), .ZN(n20999) );
  OAI211_X1 U23947 ( .C1(n21059), .C2(n21007), .A(n21000), .B(n20999), .ZN(
        P1_U3151) );
  AOI22_X1 U23948 ( .A1(n21063), .A2(n21002), .B1(n21061), .B2(n21001), .ZN(
        n21006) );
  AOI22_X1 U23949 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n21004), .B1(
        n21003), .B2(n21064), .ZN(n21005) );
  OAI211_X1 U23950 ( .C1(n21070), .C2(n21007), .A(n21006), .B(n21005), .ZN(
        P1_U3152) );
  INV_X1 U23951 ( .A(n21009), .ZN(n21062) );
  INV_X1 U23952 ( .A(n21008), .ZN(n21011) );
  OAI222_X1 U23953 ( .A1(n21012), .A2(n21011), .B1(n21074), .B2(n21015), .C1(
        n21010), .C2(n21009), .ZN(n21060) );
  AOI22_X1 U23954 ( .A1(n21014), .A2(n21062), .B1(n21013), .B2(n21060), .ZN(
        n21022) );
  OAI21_X1 U23955 ( .B1(n21017), .B2(n21016), .A(n21015), .ZN(n21019) );
  NAND2_X1 U23956 ( .A1(n21019), .A2(n21018), .ZN(n21066) );
  AOI22_X1 U23957 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21066), .B1(
        n21065), .B2(n21020), .ZN(n21021) );
  OAI211_X1 U23958 ( .C1(n21023), .C2(n21069), .A(n21022), .B(n21021), .ZN(
        P1_U3153) );
  AOI22_X1 U23959 ( .A1(n21025), .A2(n21062), .B1(n21024), .B2(n21060), .ZN(
        n21028) );
  AOI22_X1 U23960 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21066), .B1(
        n21065), .B2(n21026), .ZN(n21027) );
  OAI211_X1 U23961 ( .C1(n21029), .C2(n21069), .A(n21028), .B(n21027), .ZN(
        P1_U3154) );
  AOI22_X1 U23962 ( .A1(n21031), .A2(n21062), .B1(n21030), .B2(n21060), .ZN(
        n21034) );
  AOI22_X1 U23963 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21066), .B1(
        n21065), .B2(n21032), .ZN(n21033) );
  OAI211_X1 U23964 ( .C1(n21035), .C2(n21069), .A(n21034), .B(n21033), .ZN(
        P1_U3155) );
  AOI22_X1 U23965 ( .A1(n21037), .A2(n21062), .B1(n21036), .B2(n21060), .ZN(
        n21040) );
  AOI22_X1 U23966 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21066), .B1(
        n21065), .B2(n21038), .ZN(n21039) );
  OAI211_X1 U23967 ( .C1(n21041), .C2(n21069), .A(n21040), .B(n21039), .ZN(
        P1_U3156) );
  AOI22_X1 U23968 ( .A1(n21043), .A2(n21062), .B1(n21042), .B2(n21060), .ZN(
        n21046) );
  AOI22_X1 U23969 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21066), .B1(
        n21065), .B2(n21044), .ZN(n21045) );
  OAI211_X1 U23970 ( .C1(n21047), .C2(n21069), .A(n21046), .B(n21045), .ZN(
        P1_U3157) );
  AOI22_X1 U23971 ( .A1(n21049), .A2(n21062), .B1(n21048), .B2(n21060), .ZN(
        n21052) );
  AOI22_X1 U23972 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21066), .B1(
        n21065), .B2(n21050), .ZN(n21051) );
  OAI211_X1 U23973 ( .C1(n21053), .C2(n21069), .A(n21052), .B(n21051), .ZN(
        P1_U3158) );
  AOI22_X1 U23974 ( .A1(n21055), .A2(n21062), .B1(n21054), .B2(n21060), .ZN(
        n21058) );
  AOI22_X1 U23975 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21066), .B1(
        n21065), .B2(n21056), .ZN(n21057) );
  OAI211_X1 U23976 ( .C1(n21059), .C2(n21069), .A(n21058), .B(n21057), .ZN(
        P1_U3159) );
  AOI22_X1 U23977 ( .A1(n21063), .A2(n21062), .B1(n21061), .B2(n21060), .ZN(
        n21068) );
  AOI22_X1 U23978 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21066), .B1(
        n21065), .B2(n21064), .ZN(n21067) );
  OAI211_X1 U23979 ( .C1(n21070), .C2(n21069), .A(n21068), .B(n21067), .ZN(
        P1_U3160) );
  NOR2_X1 U23980 ( .A1(n10144), .A2(n21185), .ZN(n21073) );
  INV_X1 U23981 ( .A(n21071), .ZN(n21072) );
  OAI21_X1 U23982 ( .B1(n21074), .B2(n21073), .A(n21072), .ZN(P1_U3163) );
  AND2_X1 U23983 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21153), .ZN(
        P1_U3164) );
  AND2_X1 U23984 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21153), .ZN(
        P1_U3165) );
  AND2_X1 U23985 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21153), .ZN(
        P1_U3166) );
  AND2_X1 U23986 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21153), .ZN(
        P1_U3167) );
  AND2_X1 U23987 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21153), .ZN(
        P1_U3168) );
  AND2_X1 U23988 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21153), .ZN(
        P1_U3169) );
  AND2_X1 U23989 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21153), .ZN(
        P1_U3170) );
  AND2_X1 U23990 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21153), .ZN(
        P1_U3171) );
  AND2_X1 U23991 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21153), .ZN(
        P1_U3172) );
  AND2_X1 U23992 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21153), .ZN(
        P1_U3173) );
  AND2_X1 U23993 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21153), .ZN(
        P1_U3174) );
  AND2_X1 U23994 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21153), .ZN(
        P1_U3175) );
  AND2_X1 U23995 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21153), .ZN(
        P1_U3176) );
  AND2_X1 U23996 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21153), .ZN(
        P1_U3177) );
  AND2_X1 U23997 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21153), .ZN(
        P1_U3178) );
  INV_X1 U23998 ( .A(P1_DATAWIDTH_REG_16__SCAN_IN), .ZN(n21221) );
  NOR2_X1 U23999 ( .A1(n21157), .A2(n21221), .ZN(P1_U3179) );
  AND2_X1 U24000 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21153), .ZN(
        P1_U3180) );
  AND2_X1 U24001 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21153), .ZN(
        P1_U3181) );
  AND2_X1 U24002 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21153), .ZN(
        P1_U3182) );
  AND2_X1 U24003 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21153), .ZN(
        P1_U3183) );
  AND2_X1 U24004 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21153), .ZN(
        P1_U3184) );
  AND2_X1 U24005 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21153), .ZN(
        P1_U3185) );
  AND2_X1 U24006 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21153), .ZN(P1_U3186) );
  AND2_X1 U24007 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21153), .ZN(P1_U3187) );
  AND2_X1 U24008 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21153), .ZN(P1_U3188) );
  AND2_X1 U24009 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21153), .ZN(P1_U3189) );
  AND2_X1 U24010 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21153), .ZN(P1_U3190) );
  AND2_X1 U24011 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21153), .ZN(P1_U3191) );
  AND2_X1 U24012 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21153), .ZN(P1_U3192) );
  AND2_X1 U24013 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21153), .ZN(P1_U3193) );
  AOI21_X1 U24014 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21075), .A(n21080), 
        .ZN(n21085) );
  NOR2_X1 U24015 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n21077) );
  NAND2_X1 U24016 ( .A1(n21080), .A2(NA), .ZN(n21076) );
  OAI211_X1 U24017 ( .C1(n21090), .C2(n21077), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .B(n21076), .ZN(n21078) );
  INV_X1 U24018 ( .A(n21078), .ZN(n21079) );
  OAI22_X1 U24019 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21085), .B1(n21172), 
        .B2(n21079), .ZN(P1_U3194) );
  NOR3_X1 U24020 ( .A1(NA), .A2(n21080), .A3(n21175), .ZN(n21081) );
  OAI22_X1 U24021 ( .A1(n21082), .A2(n21081), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n21083), .ZN(n21091) );
  NOR2_X1 U24022 ( .A1(NA), .A2(n21083), .ZN(n21088) );
  AOI211_X1 U24023 ( .C1(NA), .C2(n21086), .A(n21085), .B(n21084), .ZN(n21087)
         );
  OAI21_X1 U24024 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n21088), .A(n21087), 
        .ZN(n21089) );
  OAI21_X1 U24025 ( .B1(n21091), .B2(n21090), .A(n21089), .ZN(P1_U3196) );
  NAND2_X1 U24026 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21172), .ZN(n21141) );
  NAND2_X1 U24027 ( .A1(n21172), .A2(n21092), .ZN(n21137) );
  INV_X1 U24028 ( .A(n21137), .ZN(n21143) );
  AOI222_X1 U24029 ( .A1(n21144), .A2(P1_REIP_REG_1__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n21170), .C1(P1_REIP_REG_2__SCAN_IN), 
        .C2(n21143), .ZN(n21093) );
  INV_X1 U24030 ( .A(n21093), .ZN(P1_U3197) );
  AOI222_X1 U24031 ( .A1(n21143), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n21170), .C1(P1_REIP_REG_2__SCAN_IN), 
        .C2(n21144), .ZN(n21094) );
  INV_X1 U24032 ( .A(n21094), .ZN(P1_U3198) );
  OAI222_X1 U24033 ( .A1(n21141), .A2(n21096), .B1(n21095), .B2(n21172), .C1(
        n21097), .C2(n21137), .ZN(P1_U3199) );
  INV_X1 U24034 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n21098) );
  OAI222_X1 U24035 ( .A1(n21137), .A2(n21100), .B1(n21098), .B2(n21172), .C1(
        n21097), .C2(n21141), .ZN(P1_U3200) );
  INV_X1 U24036 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n21099) );
  OAI222_X1 U24037 ( .A1(n21141), .A2(n21100), .B1(n21099), .B2(n21172), .C1(
        n21102), .C2(n21137), .ZN(P1_U3201) );
  INV_X1 U24038 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n21101) );
  OAI222_X1 U24039 ( .A1(n21141), .A2(n21102), .B1(n21101), .B2(n21172), .C1(
        n21225), .C2(n21137), .ZN(P1_U3202) );
  INV_X1 U24040 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n21300) );
  OAI222_X1 U24041 ( .A1(n21141), .A2(n21225), .B1(n21300), .B2(n21172), .C1(
        n21103), .C2(n21137), .ZN(P1_U3203) );
  INV_X1 U24042 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n21104) );
  OAI222_X1 U24043 ( .A1(n21137), .A2(n15238), .B1(n21104), .B2(n21172), .C1(
        n21103), .C2(n21141), .ZN(P1_U3204) );
  INV_X1 U24044 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n21228) );
  OAI222_X1 U24045 ( .A1(n21141), .A2(n15238), .B1(n21228), .B2(n21172), .C1(
        n21106), .C2(n21137), .ZN(P1_U3205) );
  INV_X1 U24046 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n21105) );
  OAI222_X1 U24047 ( .A1(n21141), .A2(n21106), .B1(n21105), .B2(n21172), .C1(
        n21108), .C2(n21137), .ZN(P1_U3206) );
  AOI22_X1 U24048 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n21170), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n21143), .ZN(n21107) );
  OAI21_X1 U24049 ( .B1(n21108), .B2(n21141), .A(n21107), .ZN(P1_U3207) );
  AOI22_X1 U24050 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n21170), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n21144), .ZN(n21109) );
  OAI21_X1 U24051 ( .B1(n21111), .B2(n21137), .A(n21109), .ZN(P1_U3208) );
  INV_X1 U24052 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n21110) );
  OAI222_X1 U24053 ( .A1(n21141), .A2(n21111), .B1(n21110), .B2(n21172), .C1(
        n21112), .C2(n21137), .ZN(P1_U3209) );
  INV_X1 U24054 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n21113) );
  OAI222_X1 U24055 ( .A1(n21137), .A2(n21115), .B1(n21113), .B2(n21172), .C1(
        n21112), .C2(n21141), .ZN(P1_U3210) );
  INV_X1 U24056 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n21114) );
  OAI222_X1 U24057 ( .A1(n21141), .A2(n21115), .B1(n21114), .B2(n21172), .C1(
        n21117), .C2(n21137), .ZN(P1_U3211) );
  AOI22_X1 U24058 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n21170), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n21143), .ZN(n21116) );
  OAI21_X1 U24059 ( .B1(n21117), .B2(n21141), .A(n21116), .ZN(P1_U3212) );
  AOI22_X1 U24060 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n21170), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n21144), .ZN(n21118) );
  OAI21_X1 U24061 ( .B1(n21120), .B2(n21137), .A(n21118), .ZN(P1_U3213) );
  INV_X1 U24062 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n21119) );
  OAI222_X1 U24063 ( .A1(n21141), .A2(n21120), .B1(n21119), .B2(n21172), .C1(
        n21121), .C2(n21137), .ZN(P1_U3214) );
  INV_X1 U24064 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n21122) );
  OAI222_X1 U24065 ( .A1(n21137), .A2(n21124), .B1(n21122), .B2(n21172), .C1(
        n21121), .C2(n21141), .ZN(P1_U3215) );
  INV_X1 U24066 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n21123) );
  OAI222_X1 U24067 ( .A1(n21141), .A2(n21124), .B1(n21123), .B2(n21172), .C1(
        n21126), .C2(n21137), .ZN(P1_U3216) );
  INV_X1 U24068 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n21125) );
  OAI222_X1 U24069 ( .A1(n21141), .A2(n21126), .B1(n21125), .B2(n21172), .C1(
        n21128), .C2(n21137), .ZN(P1_U3217) );
  AOI22_X1 U24070 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n21170), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21143), .ZN(n21127) );
  OAI21_X1 U24071 ( .B1(n21128), .B2(n21141), .A(n21127), .ZN(P1_U3218) );
  AOI22_X1 U24072 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n21170), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21144), .ZN(n21129) );
  OAI21_X1 U24073 ( .B1(n21131), .B2(n21137), .A(n21129), .ZN(P1_U3219) );
  INV_X1 U24074 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n21130) );
  OAI222_X1 U24075 ( .A1(n21141), .A2(n21131), .B1(n21130), .B2(n21172), .C1(
        n21133), .C2(n21137), .ZN(P1_U3220) );
  INV_X1 U24076 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n21132) );
  OAI222_X1 U24077 ( .A1(n21141), .A2(n21133), .B1(n21132), .B2(n21172), .C1(
        n21135), .C2(n21137), .ZN(P1_U3221) );
  AOI22_X1 U24078 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n21143), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21170), .ZN(n21134) );
  OAI21_X1 U24079 ( .B1(n21135), .B2(n21141), .A(n21134), .ZN(P1_U3222) );
  AOI22_X1 U24080 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n21144), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21170), .ZN(n21136) );
  OAI21_X1 U24081 ( .B1(n21140), .B2(n21137), .A(n21136), .ZN(P1_U3223) );
  INV_X1 U24082 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n21139) );
  OAI222_X1 U24083 ( .A1(n21141), .A2(n21140), .B1(n21139), .B2(n21172), .C1(
        n21138), .C2(n21137), .ZN(P1_U3224) );
  AOI222_X1 U24084 ( .A1(n21143), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21170), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n21144), .ZN(n21142) );
  INV_X1 U24085 ( .A(n21142), .ZN(P1_U3225) );
  AOI222_X1 U24086 ( .A1(n21144), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21170), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n21143), .ZN(n21145) );
  INV_X1 U24087 ( .A(n21145), .ZN(P1_U3226) );
  INV_X1 U24088 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n21146) );
  AOI22_X1 U24089 ( .A1(n21172), .A2(n21147), .B1(n21146), .B2(n21170), .ZN(
        P1_U3458) );
  INV_X1 U24090 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21165) );
  INV_X1 U24091 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n21148) );
  AOI22_X1 U24092 ( .A1(n21172), .A2(n21165), .B1(n21148), .B2(n21170), .ZN(
        P1_U3459) );
  INV_X1 U24093 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n21149) );
  AOI22_X1 U24094 ( .A1(n21172), .A2(n21150), .B1(n21149), .B2(n21170), .ZN(
        P1_U3460) );
  INV_X1 U24095 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21168) );
  INV_X1 U24096 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n21151) );
  AOI22_X1 U24097 ( .A1(n21172), .A2(n21168), .B1(n21151), .B2(n21170), .ZN(
        P1_U3461) );
  INV_X1 U24098 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21154) );
  INV_X1 U24099 ( .A(n21155), .ZN(n21152) );
  AOI21_X1 U24100 ( .B1(n21154), .B2(n21153), .A(n21152), .ZN(P1_U3464) );
  OAI21_X1 U24101 ( .B1(n21157), .B2(n21156), .A(n21155), .ZN(P1_U3465) );
  INV_X1 U24102 ( .A(n21158), .ZN(n21160) );
  OAI22_X1 U24103 ( .A1(n21160), .A2(n21189), .B1(n21159), .B2(n21186), .ZN(
        n21161) );
  MUX2_X1 U24104 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n21161), .S(
        n21192), .Z(P1_U3469) );
  AOI21_X1 U24105 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21163) );
  AOI22_X1 U24106 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21163), .B2(n21162), .ZN(n21166) );
  AOI22_X1 U24107 ( .A1(n21169), .A2(n21166), .B1(n21165), .B2(n21164), .ZN(
        P1_U3481) );
  OAI21_X1 U24108 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n21169), .ZN(n21167) );
  OAI21_X1 U24109 ( .B1(n21169), .B2(n21168), .A(n21167), .ZN(P1_U3482) );
  AOI22_X1 U24110 ( .A1(n21172), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21171), 
        .B2(n21170), .ZN(P1_U3483) );
  AOI211_X1 U24111 ( .C1(n21176), .C2(n21175), .A(n21174), .B(n21173), .ZN(
        n21183) );
  INV_X1 U24112 ( .A(n10847), .ZN(n21178) );
  OAI211_X1 U24113 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21178), .A(n21177), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21180) );
  AOI21_X1 U24114 ( .B1(n21180), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n21179), 
        .ZN(n21182) );
  NAND2_X1 U24115 ( .A1(n21183), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21181) );
  OAI21_X1 U24116 ( .B1(n21183), .B2(n21182), .A(n21181), .ZN(P1_U3485) );
  MUX2_X1 U24117 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n21172), .Z(P1_U3486) );
  OAI21_X1 U24118 ( .B1(n21184), .B2(n21189), .A(n21192), .ZN(n21193) );
  OAI22_X1 U24119 ( .A1(n21186), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21185), .ZN(n21187) );
  INV_X1 U24120 ( .A(n21187), .ZN(n21188) );
  OAI21_X1 U24121 ( .B1(n21190), .B2(n21189), .A(n21188), .ZN(n21191) );
  AOI22_X1 U24122 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21193), .B1(
        n21192), .B2(n21191), .ZN(n21354) );
  NAND4_X1 U24123 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n21303), .A3(n21272), 
        .A4(n21267), .ZN(n21205) );
  NOR4_X1 U24124 ( .A1(BUF1_REG_13__SCAN_IN), .A2(P3_DATAO_REG_17__SCAN_IN), 
        .A3(P3_ADDRESS_REG_10__SCAN_IN), .A4(n21294), .ZN(n21198) );
  INV_X1 U24125 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n21301) );
  NOR3_X1 U24126 ( .A1(P2_EAX_REG_28__SCAN_IN), .A2(P2_EAX_REG_31__SCAN_IN), 
        .A3(n21301), .ZN(n21197) );
  INV_X1 U24127 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n21195) );
  NOR4_X1 U24128 ( .A1(n21195), .A2(n21300), .A3(n21194), .A4(
        P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n21196) );
  NAND4_X1 U24129 ( .A1(n21198), .A2(n21197), .A3(n21196), .A4(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n21204) );
  NAND4_X1 U24130 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_LWORD_REG_11__SCAN_IN), .A4(
        n21320), .ZN(n21203) );
  NOR4_X1 U24131 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(
        P2_EBX_REG_6__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_UWORD_REG_3__SCAN_IN), .ZN(n21201) );
  NOR3_X1 U24132 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(P2_DATAO_REG_24__SCAN_IN), 
        .ZN(n21200) );
  NOR4_X1 U24133 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_15__3__SCAN_IN), .A3(n21315), .A4(n21318), .ZN(n21199) );
  NAND4_X1 U24134 ( .A1(n21201), .A2(P1_DATAO_REG_26__SCAN_IN), .A3(n21200), 
        .A4(n21199), .ZN(n21202) );
  NOR4_X1 U24135 ( .A1(n21205), .A2(n21204), .A3(n21203), .A4(n21202), .ZN(
        n21352) );
  INV_X1 U24136 ( .A(n21206), .ZN(n21219) );
  INV_X1 U24137 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n21227) );
  INV_X1 U24138 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n21207) );
  NOR4_X1 U24139 ( .A1(n21227), .A2(n21285), .A3(n21207), .A4(
        P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n21211) );
  NAND2_X1 U24140 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n21209) );
  NOR4_X1 U24141 ( .A1(n21209), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        P1_ADDRESS_REG_8__SCAN_IN), .A4(n21208), .ZN(n21210) );
  NAND3_X1 U24142 ( .A1(n21211), .A2(n21210), .A3(
        P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n21218) );
  INV_X1 U24143 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n21240) );
  NOR4_X1 U24144 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(n21237), .A4(n21240), .ZN(n21215)
         );
  NOR4_X1 U24145 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_UWORD_REG_4__SCAN_IN), 
        .A3(n21246), .A4(n21239), .ZN(n21214) );
  NOR4_X1 U24146 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A4(
        n15706), .ZN(n21213) );
  INV_X1 U24147 ( .A(DATAI_17_), .ZN(n21269) );
  NOR4_X1 U24148 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .A3(P3_REIP_REG_13__SCAN_IN), .A4(
        n21269), .ZN(n21212) );
  NAND4_X1 U24149 ( .A1(n21215), .A2(n21214), .A3(n21213), .A4(n21212), .ZN(
        n21217) );
  NAND4_X1 U24150 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(
        P3_DATAO_REG_30__SCAN_IN), .A3(n21304), .A4(n21225), .ZN(n21216) );
  NOR4_X1 U24151 ( .A1(n21219), .A2(n21218), .A3(n21217), .A4(n21216), .ZN(
        n21351) );
  AOI22_X1 U24152 ( .A1(n21222), .A2(keyinput43), .B1(keyinput44), .B2(n21221), 
        .ZN(n21220) );
  OAI221_X1 U24153 ( .B1(n21222), .B2(keyinput43), .C1(n21221), .C2(keyinput44), .A(n21220), .ZN(n21234) );
  AOI22_X1 U24154 ( .A1(n21225), .A2(keyinput46), .B1(keyinput42), .B2(n21224), 
        .ZN(n21223) );
  OAI221_X1 U24155 ( .B1(n21225), .B2(keyinput46), .C1(n21224), .C2(keyinput42), .A(n21223), .ZN(n21233) );
  AOI22_X1 U24156 ( .A1(n21228), .A2(keyinput45), .B1(n21227), .B2(keyinput59), 
        .ZN(n21226) );
  OAI221_X1 U24157 ( .B1(n21228), .B2(keyinput45), .C1(n21227), .C2(keyinput59), .A(n21226), .ZN(n21232) );
  XNOR2_X1 U24158 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B(keyinput49), .ZN(
        n21230) );
  XNOR2_X1 U24159 ( .A(keyinput10), .B(P1_EBX_REG_1__SCAN_IN), .ZN(n21229) );
  NAND2_X1 U24160 ( .A1(n21230), .A2(n21229), .ZN(n21231) );
  NOR4_X1 U24161 ( .A1(n21234), .A2(n21233), .A3(n21232), .A4(n21231), .ZN(
        n21283) );
  AOI22_X1 U24162 ( .A1(n21237), .A2(keyinput37), .B1(keyinput22), .B2(n21236), 
        .ZN(n21235) );
  OAI221_X1 U24163 ( .B1(n21237), .B2(keyinput37), .C1(n21236), .C2(keyinput22), .A(n21235), .ZN(n21250) );
  AOI22_X1 U24164 ( .A1(n21240), .A2(keyinput53), .B1(keyinput3), .B2(n21239), 
        .ZN(n21238) );
  OAI221_X1 U24165 ( .B1(n21240), .B2(keyinput53), .C1(n21239), .C2(keyinput3), 
        .A(n21238), .ZN(n21249) );
  AOI22_X1 U24166 ( .A1(n21243), .A2(keyinput23), .B1(keyinput57), .B2(n21242), 
        .ZN(n21241) );
  OAI221_X1 U24167 ( .B1(n21243), .B2(keyinput23), .C1(n21242), .C2(keyinput57), .A(n21241), .ZN(n21248) );
  AOI22_X1 U24168 ( .A1(n21246), .A2(keyinput5), .B1(keyinput26), .B2(n21245), 
        .ZN(n21244) );
  OAI221_X1 U24169 ( .B1(n21246), .B2(keyinput5), .C1(n21245), .C2(keyinput26), 
        .A(n21244), .ZN(n21247) );
  NOR4_X1 U24170 ( .A1(n21250), .A2(n21249), .A3(n21248), .A4(n21247), .ZN(
        n21282) );
  INV_X1 U24171 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n21253) );
  AOI22_X1 U24172 ( .A1(n21253), .A2(keyinput60), .B1(n21252), .B2(keyinput38), 
        .ZN(n21251) );
  OAI221_X1 U24173 ( .B1(n21253), .B2(keyinput60), .C1(n21252), .C2(keyinput38), .A(n21251), .ZN(n21264) );
  INV_X1 U24174 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n21255) );
  AOI22_X1 U24175 ( .A1(n21256), .A2(keyinput14), .B1(n21255), .B2(keyinput21), 
        .ZN(n21254) );
  OAI221_X1 U24176 ( .B1(n21256), .B2(keyinput14), .C1(n21255), .C2(keyinput21), .A(n21254), .ZN(n21263) );
  XOR2_X1 U24177 ( .A(n15706), .B(keyinput33), .Z(n21259) );
  XNOR2_X1 U24178 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B(keyinput7), .ZN(
        n21258) );
  XNOR2_X1 U24179 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B(keyinput41), .ZN(
        n21257) );
  NAND3_X1 U24180 ( .A1(n21259), .A2(n21258), .A3(n21257), .ZN(n21262) );
  XNOR2_X1 U24181 ( .A(n21260), .B(keyinput58), .ZN(n21261) );
  NOR4_X1 U24182 ( .A1(n21264), .A2(n21263), .A3(n21262), .A4(n21261), .ZN(
        n21281) );
  AOI22_X1 U24183 ( .A1(n21267), .A2(keyinput62), .B1(keyinput18), .B2(n21266), 
        .ZN(n21265) );
  OAI221_X1 U24184 ( .B1(n21267), .B2(keyinput62), .C1(n21266), .C2(keyinput18), .A(n21265), .ZN(n21279) );
  AOI22_X1 U24185 ( .A1(n21270), .A2(keyinput16), .B1(keyinput2), .B2(n21269), 
        .ZN(n21268) );
  OAI221_X1 U24186 ( .B1(n21270), .B2(keyinput16), .C1(n21269), .C2(keyinput2), 
        .A(n21268), .ZN(n21278) );
  AOI22_X1 U24187 ( .A1(n21273), .A2(keyinput34), .B1(n21272), .B2(keyinput8), 
        .ZN(n21271) );
  OAI221_X1 U24188 ( .B1(n21273), .B2(keyinput34), .C1(n21272), .C2(keyinput8), 
        .A(n21271), .ZN(n21277) );
  XNOR2_X1 U24189 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B(keyinput24), .ZN(
        n21275) );
  XNOR2_X1 U24190 ( .A(P2_REIP_REG_20__SCAN_IN), .B(keyinput35), .ZN(n21274)
         );
  NAND2_X1 U24191 ( .A1(n21275), .A2(n21274), .ZN(n21276) );
  NOR4_X1 U24192 ( .A1(n21279), .A2(n21278), .A3(n21277), .A4(n21276), .ZN(
        n21280) );
  NAND4_X1 U24193 ( .A1(n21283), .A2(n21282), .A3(n21281), .A4(n21280), .ZN(
        n21350) );
  AOI22_X1 U24194 ( .A1(n21286), .A2(keyinput11), .B1(keyinput55), .B2(n21285), 
        .ZN(n21284) );
  OAI221_X1 U24195 ( .B1(n21286), .B2(keyinput11), .C1(n21285), .C2(keyinput55), .A(n21284), .ZN(n21298) );
  INV_X1 U24196 ( .A(P2_EAX_REG_31__SCAN_IN), .ZN(n21289) );
  AOI22_X1 U24197 ( .A1(n21289), .A2(keyinput36), .B1(n21288), .B2(keyinput56), 
        .ZN(n21287) );
  OAI221_X1 U24198 ( .B1(n21289), .B2(keyinput36), .C1(n21288), .C2(keyinput56), .A(n21287), .ZN(n21297) );
  AOI22_X1 U24199 ( .A1(n21291), .A2(keyinput51), .B1(n13849), .B2(keyinput6), 
        .ZN(n21290) );
  OAI221_X1 U24200 ( .B1(n21291), .B2(keyinput51), .C1(n13849), .C2(keyinput6), 
        .A(n21290), .ZN(n21296) );
  AOI22_X1 U24201 ( .A1(n21294), .A2(keyinput61), .B1(keyinput30), .B2(n21293), 
        .ZN(n21292) );
  OAI221_X1 U24202 ( .B1(n21294), .B2(keyinput61), .C1(n21293), .C2(keyinput30), .A(n21292), .ZN(n21295) );
  NOR4_X1 U24203 ( .A1(n21298), .A2(n21297), .A3(n21296), .A4(n21295), .ZN(
        n21348) );
  AOI22_X1 U24204 ( .A1(n21301), .A2(keyinput1), .B1(keyinput12), .B2(n21300), 
        .ZN(n21299) );
  OAI221_X1 U24205 ( .B1(n21301), .B2(keyinput1), .C1(n21300), .C2(keyinput12), 
        .A(n21299), .ZN(n21312) );
  AOI22_X1 U24206 ( .A1(n21304), .A2(keyinput17), .B1(n21303), .B2(keyinput47), 
        .ZN(n21302) );
  OAI221_X1 U24207 ( .B1(n21304), .B2(keyinput17), .C1(n21303), .C2(keyinput47), .A(n21302), .ZN(n21311) );
  XNOR2_X1 U24208 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B(keyinput50), .ZN(
        n21307) );
  XNOR2_X1 U24209 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B(keyinput28), .ZN(
        n21306) );
  XNOR2_X1 U24210 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B(keyinput19), .ZN(
        n21305) );
  NAND3_X1 U24211 ( .A1(n21307), .A2(n21306), .A3(n21305), .ZN(n21310) );
  XNOR2_X1 U24212 ( .A(n21308), .B(keyinput48), .ZN(n21309) );
  NOR4_X1 U24213 ( .A1(n21312), .A2(n21311), .A3(n21310), .A4(n21309), .ZN(
        n21347) );
  INV_X1 U24214 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n21314) );
  AOI22_X1 U24215 ( .A1(n21315), .A2(keyinput15), .B1(n21314), .B2(keyinput27), 
        .ZN(n21313) );
  OAI221_X1 U24216 ( .B1(n21315), .B2(keyinput15), .C1(n21314), .C2(keyinput27), .A(n21313), .ZN(n21328) );
  INV_X1 U24217 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n21317) );
  AOI22_X1 U24218 ( .A1(n21318), .A2(keyinput0), .B1(n21317), .B2(keyinput32), 
        .ZN(n21316) );
  OAI221_X1 U24219 ( .B1(n21318), .B2(keyinput0), .C1(n21317), .C2(keyinput32), 
        .A(n21316), .ZN(n21327) );
  AOI22_X1 U24220 ( .A1(n21321), .A2(keyinput54), .B1(n21320), .B2(keyinput29), 
        .ZN(n21319) );
  OAI221_X1 U24221 ( .B1(n21321), .B2(keyinput54), .C1(n21320), .C2(keyinput29), .A(n21319), .ZN(n21326) );
  INV_X1 U24222 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n21324) );
  AOI22_X1 U24223 ( .A1(n21324), .A2(keyinput4), .B1(keyinput9), .B2(n21323), 
        .ZN(n21322) );
  OAI221_X1 U24224 ( .B1(n21324), .B2(keyinput4), .C1(n21323), .C2(keyinput9), 
        .A(n21322), .ZN(n21325) );
  NOR4_X1 U24225 ( .A1(n21328), .A2(n21327), .A3(n21326), .A4(n21325), .ZN(
        n21346) );
  AOI22_X1 U24226 ( .A1(n21331), .A2(keyinput52), .B1(n21330), .B2(keyinput40), 
        .ZN(n21329) );
  OAI221_X1 U24227 ( .B1(n21331), .B2(keyinput52), .C1(n21330), .C2(keyinput40), .A(n21329), .ZN(n21344) );
  INV_X1 U24228 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n21334) );
  AOI22_X1 U24229 ( .A1(n21334), .A2(keyinput25), .B1(keyinput39), .B2(n21333), 
        .ZN(n21332) );
  OAI221_X1 U24230 ( .B1(n21334), .B2(keyinput25), .C1(n21333), .C2(keyinput39), .A(n21332), .ZN(n21343) );
  AOI22_X1 U24231 ( .A1(n21337), .A2(keyinput63), .B1(n21336), .B2(keyinput31), 
        .ZN(n21335) );
  OAI221_X1 U24232 ( .B1(n21337), .B2(keyinput63), .C1(n21336), .C2(keyinput31), .A(n21335), .ZN(n21342) );
  INV_X1 U24233 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n21340) );
  AOI22_X1 U24234 ( .A1(n21340), .A2(keyinput20), .B1(keyinput13), .B2(n21339), 
        .ZN(n21338) );
  OAI221_X1 U24235 ( .B1(n21340), .B2(keyinput20), .C1(n21339), .C2(keyinput13), .A(n21338), .ZN(n21341) );
  NOR4_X1 U24236 ( .A1(n21344), .A2(n21343), .A3(n21342), .A4(n21341), .ZN(
        n21345) );
  NAND4_X1 U24237 ( .A1(n21348), .A2(n21347), .A3(n21346), .A4(n21345), .ZN(
        n21349) );
  AOI211_X1 U24238 ( .C1(n21352), .C2(n21351), .A(n21350), .B(n21349), .ZN(
        n21353) );
  XNOR2_X1 U24239 ( .A(n21354), .B(n21353), .ZN(P1_U3474) );
  AND2_X1 U13098 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17327) );
  NOR2_X2 U12983 ( .A1(n18108), .A2(n18113), .ZN(n12600) );
  NOR2_X2 U13408 ( .A1(n17199), .A2(n18112), .ZN(n17198) );
  OR2_X2 U13415 ( .A1(n17137), .A2(n17138), .ZN(n10326) );
  INV_X2 U13410 ( .A(n18217), .ZN(n10309) );
  AND2_X2 U13920 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13457) );
  INV_X1 U13242 ( .A(n17563), .ZN(n14305) );
  BUF_X2 U11036 ( .A(n11890), .Z(n14461) );
  CLKBUF_X2 U11059 ( .A(n10705), .Z(n11268) );
  CLKBUF_X1 U11066 ( .A(n10791), .Z(n11303) );
  CLKBUF_X2 U11076 ( .A(n10732), .Z(n11280) );
  CLKBUF_X1 U11108 ( .A(n11436), .Z(n13712) );
  NAND2_X2 U11182 ( .A1(n10778), .A2(n9659), .ZN(n11438) );
  CLKBUF_X1 U11347 ( .A(n12230), .Z(n12563) );
  NOR2_X1 U11366 ( .A1(n18059), .A2(n17156), .ZN(n17155) );
  CLKBUF_X1 U11440 ( .A(n14109), .Z(n14110) );
  CLKBUF_X2 U11546 ( .A(n10319), .Z(n17434) );
  AOI211_X1 U11618 ( .C1(n17142), .C2(n17141), .A(n17140), .B(n17139), .ZN(
        n17143) );
  CLKBUF_X1 U11680 ( .A(n17085), .Z(n17090) );
  NOR2_X2 U12349 ( .A1(n14013), .A2(n14010), .ZN(n21355) );
  CLKBUF_X1 U12631 ( .A(n18031), .Z(n18039) );
endmodule

