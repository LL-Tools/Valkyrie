

module b14_C_gen_AntiSAT_k_256_10 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085;

  OR2_X1 U2462 ( .A1(n3148), .A2(n2424), .ZN(n2423) );
  AND2_X1 U2464 ( .A1(n2841), .A2(n2840), .ZN(n4404) );
  XNOR2_X2 U2465 ( .A(n2788), .B(n2787), .ZN(n3831) );
  AND2_X2 U2466 ( .A1(n2417), .A2(n2416), .ZN(n3132) );
  NOR2_X1 U2467 ( .A1(n4454), .A2(n3916), .ZN(n4466) );
  NAND2_X1 U2468 ( .A1(n2542), .A2(n2478), .ZN(n3853) );
  AND2_X2 U2469 ( .A1(n2932), .A2(n4694), .ZN(n3513) );
  NOR2_X1 U2470 ( .A1(n4445), .A2(n4444), .ZN(n4443) );
  NAND3_X1 U2471 ( .A1(n4404), .A2(n4405), .A3(n2323), .ZN(n3034) );
  AND2_X2 U2472 ( .A1(n2508), .A2(n2509), .ZN(n3706) );
  AND3_X1 U2473 ( .A1(n2467), .A2(n2243), .A3(n2316), .ZN(n2495) );
  XNOR2_X1 U2474 ( .A(n2785), .B(n2784), .ZN(n3940) );
  NAND2_X1 U2475 ( .A1(n2316), .A2(n2344), .ZN(n2727) );
  NOR2_X1 U2476 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2475)
         );
  NOR2_X1 U2477 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2480)
         );
  NOR2_X1 U2478 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2481)
         );
  NOR2_X1 U2479 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2482)
         );
  INV_X1 U2480 ( .A(n2976), .ZN(n3008) );
  NOR2_X1 U2481 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2494)
         );
  NAND2_X1 U2482 ( .A1(n2882), .A2(IR_REG_28__SCAN_IN), .ZN(n2398) );
  INV_X1 U2483 ( .A(n2468), .ZN(n2467) );
  AND2_X1 U2484 ( .A1(n2317), .A2(n2456), .ZN(n2316) );
  AND2_X1 U2485 ( .A1(n2396), .A2(n2488), .ZN(n2317) );
  INV_X1 U2486 ( .A(IR_REG_18__SCAN_IN), .ZN(n2488) );
  NOR2_X1 U2487 ( .A1(n4091), .A2(n2459), .ZN(n2458) );
  INV_X1 U2488 ( .A(n2719), .ZN(n2459) );
  NAND2_X1 U2489 ( .A1(n3757), .A2(n3831), .ZN(n2976) );
  INV_X1 U2490 ( .A(n4471), .ZN(n2265) );
  NOR2_X1 U2491 ( .A1(n2295), .A2(n2245), .ZN(n2292) );
  OR2_X1 U2492 ( .A1(n3222), .A2(n3220), .ZN(n2800) );
  INV_X1 U2493 ( .A(n3327), .ZN(n3314) );
  NAND2_X1 U2494 ( .A1(n3755), .A2(n3758), .ZN(n4620) );
  NOR2_X1 U2495 ( .A1(n2907), .A2(n2858), .ZN(n2938) );
  INV_X1 U2496 ( .A(n2550), .ZN(n2397) );
  NAND2_X1 U2497 ( .A1(n2469), .A2(n2789), .ZN(n2468) );
  INV_X1 U2498 ( .A(n2470), .ZN(n2469) );
  INV_X1 U2499 ( .A(n2483), .ZN(n2456) );
  AND4_X1 U2500 ( .A1(n2693), .A2(n2484), .A3(n2485), .A4(n2669), .ZN(n2486)
         );
  INV_X1 U2501 ( .A(IR_REG_16__SCAN_IN), .ZN(n2484) );
  INV_X1 U2502 ( .A(IR_REG_14__SCAN_IN), .ZN(n2485) );
  AOI21_X1 U2503 ( .B1(n2331), .B2(n2329), .A(n2225), .ZN(n2328) );
  INV_X1 U2504 ( .A(n3513), .ZN(n3548) );
  AOI22_X1 U2505 ( .A1(n4614), .A2(n3479), .B1(n2933), .B2(n2932), .ZN(n2981)
         );
  NAND2_X1 U2506 ( .A1(n2931), .A2(n2930), .ZN(n2936) );
  INV_X1 U2507 ( .A(n2929), .ZN(n2930) );
  OAI22_X1 U2508 ( .A1(n3551), .A2(n4629), .B1(n3034), .B2(n2928), .ZN(n2929)
         );
  NAND2_X1 U2509 ( .A1(n4406), .A2(n3940), .ZN(n2447) );
  INV_X1 U2510 ( .A(n3706), .ZN(n2772) );
  XNOR2_X1 U2511 ( .A(n3891), .B(n2386), .ZN(n4476) );
  XNOR2_X1 U2512 ( .A(n3894), .B(n2385), .ZN(n4497) );
  XNOR2_X1 U2513 ( .A(n3897), .B(n2384), .ZN(n4518) );
  AOI21_X1 U2514 ( .B1(n4072), .B2(n2745), .A(n2744), .ZN(n4061) );
  INV_X2 U2515 ( .A(n2553), .ZN(n2544) );
  NAND2_X1 U2516 ( .A1(n3852), .A2(n3763), .ZN(n2285) );
  INV_X1 U2517 ( .A(n2543), .ZN(n2287) );
  AND2_X1 U2518 ( .A1(n2486), .A2(n2397), .ZN(n2344) );
  XNOR2_X1 U2519 ( .A(n2342), .B(n2473), .ZN(n2509) );
  NAND2_X1 U2520 ( .A1(n2507), .A2(IR_REG_31__SCAN_IN), .ZN(n2342) );
  NAND2_X1 U2521 ( .A1(n2394), .A2(n2705), .ZN(n2393) );
  INV_X1 U2522 ( .A(n3482), .ZN(n2442) );
  NAND2_X1 U2523 ( .A1(n3482), .A2(n2441), .ZN(n2440) );
  INV_X1 U2524 ( .A(n2443), .ZN(n2441) );
  AND2_X1 U2525 ( .A1(n4425), .A2(n3606), .ZN(n2320) );
  INV_X1 U2526 ( .A(n4450), .ZN(n2268) );
  NAND2_X1 U2527 ( .A1(n3671), .A2(n4011), .ZN(n2453) );
  INV_X1 U2528 ( .A(n4000), .ZN(n2454) );
  INV_X1 U2529 ( .A(n2449), .ZN(n2311) );
  INV_X1 U2530 ( .A(n3729), .ZN(n2448) );
  NAND2_X1 U2531 ( .A1(n2369), .A2(n2464), .ZN(n2367) );
  AOI21_X1 U2532 ( .B1(n3794), .B2(n3793), .A(n2358), .ZN(n2357) );
  INV_X1 U2533 ( .A(n3797), .ZN(n2358) );
  NOR2_X1 U2534 ( .A1(n2245), .A2(n2294), .ZN(n2293) );
  INV_X1 U2535 ( .A(n3775), .ZN(n2380) );
  INV_X1 U2536 ( .A(n3781), .ZN(n2377) );
  NOR2_X1 U2537 ( .A1(n2410), .A2(n4029), .ZN(n2408) );
  NAND2_X1 U2538 ( .A1(n4118), .A2(n2807), .ZN(n2406) );
  NAND2_X1 U2539 ( .A1(n4187), .A2(n2682), .ZN(n2465) );
  AND2_X1 U2540 ( .A1(n2401), .A2(n3401), .ZN(n2400) );
  AND2_X1 U2541 ( .A1(n3314), .A2(n4604), .ZN(n2401) );
  OR2_X1 U2542 ( .A1(n3193), .A2(n3265), .ZN(n3225) );
  NAND2_X1 U2543 ( .A1(n2471), .A2(n2782), .ZN(n2470) );
  INV_X1 U2544 ( .A(n2489), .ZN(n2471) );
  INV_X1 U2545 ( .A(IR_REG_20__SCAN_IN), .ZN(n2787) );
  INV_X1 U2546 ( .A(IR_REG_15__SCAN_IN), .ZN(n2693) );
  NAND2_X1 U2547 ( .A1(n2421), .A2(n3208), .ZN(n2420) );
  INV_X1 U2548 ( .A(n3205), .ZN(n2421) );
  OR2_X1 U2549 ( .A1(n2767), .A2(n3515), .ZN(n2774) );
  INV_X1 U2550 ( .A(n4614), .ZN(n2990) );
  XNOR2_X1 U2551 ( .A(n3137), .B(n3399), .ZN(n3138) );
  NAND2_X1 U2552 ( .A1(n3454), .A2(n3453), .ZN(n3455) );
  INV_X1 U2553 ( .A(n3452), .ZN(n3454) );
  INV_X1 U2554 ( .A(n3336), .ZN(n2336) );
  NOR2_X1 U2555 ( .A1(n3581), .A2(n2434), .ZN(n2433) );
  INV_X1 U2556 ( .A(n2436), .ZN(n2434) );
  INV_X1 U2557 ( .A(n2335), .ZN(n2334) );
  OAI21_X1 U2558 ( .B1(n2230), .B2(n2336), .A(n2432), .ZN(n2335) );
  AND2_X1 U2559 ( .A1(n2437), .A2(n3582), .ZN(n2432) );
  AOI22_X1 U2560 ( .A1(n3853), .A2(n3479), .B1(n2932), .B2(n3048), .ZN(n3015)
         );
  AND2_X1 U2561 ( .A1(n2537), .A2(REG3_REG_0__SCAN_IN), .ZN(n2522) );
  AOI21_X1 U2562 ( .B1(n2962), .B2(REG2_REG_3__SCAN_IN), .A(n2269), .ZN(n3886)
         );
  AND2_X1 U2563 ( .A1(n2270), .A2(n4409), .ZN(n2269) );
  AND2_X1 U2564 ( .A1(n3910), .A2(n2339), .ZN(n4445) );
  NAND2_X1 U2565 ( .A1(n3911), .A2(n4408), .ZN(n2339) );
  OAI21_X1 U2566 ( .B1(n4459), .B2(n2265), .A(n2263), .ZN(n3891) );
  INV_X1 U2567 ( .A(n2264), .ZN(n2263) );
  OAI21_X1 U2568 ( .B1(n3889), .B2(n2265), .A(n3890), .ZN(n2264) );
  NAND2_X1 U2569 ( .A1(n4485), .A2(n4486), .ZN(n4484) );
  NAND2_X1 U2570 ( .A1(n4487), .A2(n3893), .ZN(n3894) );
  NAND2_X1 U2571 ( .A1(n4497), .A2(REG2_REG_10__SCAN_IN), .ZN(n4496) );
  NAND2_X1 U2572 ( .A1(n4506), .A2(n4507), .ZN(n4505) );
  NAND2_X1 U2573 ( .A1(n4508), .A2(n3896), .ZN(n3897) );
  NAND2_X1 U2574 ( .A1(n4518), .A2(REG2_REG_12__SCAN_IN), .ZN(n4517) );
  OAI22_X1 U2575 ( .A1(n4530), .A2(n4526), .B1(REG2_REG_13__SCAN_IN), .B2(
        n3907), .ZN(n3899) );
  NAND2_X1 U2576 ( .A1(n4569), .A2(n2392), .ZN(n2391) );
  NAND2_X1 U2577 ( .A1(n4645), .A2(n4155), .ZN(n2392) );
  NAND2_X1 U2578 ( .A1(n4005), .A2(n3992), .ZN(n2452) );
  AND2_X1 U2579 ( .A1(n2251), .A2(n2766), .ZN(n2304) );
  NAND2_X1 U2580 ( .A1(n4061), .A2(n4060), .ZN(n2450) );
  AND2_X1 U2581 ( .A1(n2457), .A2(n2277), .ZN(n2276) );
  NAND2_X1 U2582 ( .A1(n2280), .A2(n2709), .ZN(n4129) );
  NAND2_X1 U2583 ( .A1(n4150), .A2(n2708), .ZN(n2280) );
  NAND2_X1 U2584 ( .A1(n2802), .A2(n3792), .ZN(n3366) );
  NAND2_X1 U2585 ( .A1(n2347), .A2(n2345), .ZN(n2802) );
  AOI21_X1 U2586 ( .B1(n2348), .B2(n2351), .A(n2346), .ZN(n2345) );
  NAND2_X1 U2587 ( .A1(n2256), .A2(n2224), .ZN(n2295) );
  NAND2_X1 U2588 ( .A1(n2246), .A2(n2634), .ZN(n2296) );
  NAND2_X1 U2589 ( .A1(n2634), .A2(n2224), .ZN(n2294) );
  OAI21_X1 U2590 ( .B1(n3224), .B2(n2624), .A(n2623), .ZN(n3297) );
  OAI21_X1 U2591 ( .B1(n3093), .B2(n3092), .A(n3778), .ZN(n3118) );
  OAI21_X1 U2592 ( .B1(n3100), .B2(n2574), .A(n2575), .ZN(n3117) );
  AND2_X1 U2593 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2564) );
  AND2_X1 U2594 ( .A1(n2794), .A2(n2536), .ZN(n2451) );
  NAND2_X1 U2595 ( .A1(n2791), .A2(n3940), .ZN(n4621) );
  AND2_X1 U2596 ( .A1(n3970), .A2(n3559), .ZN(n2888) );
  AND2_X1 U2597 ( .A1(n3990), .A2(n3976), .ZN(n3970) );
  AND2_X1 U2598 ( .A1(n2780), .A2(n2779), .ZN(n4240) );
  NOR2_X1 U2599 ( .A1(n4010), .A2(n3500), .ZN(n3990) );
  INV_X1 U2600 ( .A(n3474), .ZN(n4064) );
  AND2_X1 U2601 ( .A1(n4077), .A2(n4064), .ZN(n4066) );
  NOR2_X1 U2602 ( .A1(n4095), .A2(n4266), .ZN(n4077) );
  NOR2_X1 U2603 ( .A1(n4210), .A2(n4316), .ZN(n4211) );
  OR2_X1 U2604 ( .A1(n2996), .A2(n3831), .ZN(n4328) );
  INV_X1 U2605 ( .A(n3853), .ZN(n4617) );
  NAND2_X1 U2606 ( .A1(n2997), .A2(n2829), .ZN(n4695) );
  OR2_X1 U2607 ( .A1(n2996), .A2(n4407), .ZN(n4694) );
  NAND2_X1 U2608 ( .A1(n2842), .A2(n4404), .ZN(n2907) );
  INV_X1 U2609 ( .A(n2495), .ZN(n2838) );
  NAND2_X1 U2610 ( .A1(n2495), .A2(n2492), .ZN(n2840) );
  INV_X1 U2611 ( .A(IR_REG_26__SCAN_IN), .ZN(n2492) );
  OAI21_X1 U2612 ( .B1(n2727), .B2(n2468), .A(IR_REG_31__SCAN_IN), .ZN(n2846)
         );
  INV_X1 U2613 ( .A(IR_REG_31__SCAN_IN), .ZN(n2705) );
  NOR2_X2 U2614 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2534)
         );
  NOR2_X1 U2615 ( .A1(n2226), .A2(n3678), .ZN(n2325) );
  NAND2_X1 U2616 ( .A1(n2328), .A2(n2330), .ZN(n2327) );
  INV_X1 U2617 ( .A(n2331), .ZN(n2330) );
  NAND2_X1 U2618 ( .A1(n3408), .A2(n2318), .ZN(n3523) );
  NAND2_X1 U2619 ( .A1(n3635), .A2(n3637), .ZN(n2318) );
  OAI21_X1 U2620 ( .B1(n3593), .B2(n2329), .A(n2425), .ZN(n3558) );
  AND2_X1 U2621 ( .A1(n2429), .A2(n2426), .ZN(n2425) );
  NAND2_X1 U2622 ( .A1(n2428), .A2(n2427), .ZN(n2426) );
  NOR2_X1 U2623 ( .A1(n2430), .A2(n3666), .ZN(n2429) );
  OR2_X1 U2624 ( .A1(n2982), .A2(n3399), .ZN(n2983) );
  NAND2_X1 U2625 ( .A1(n2515), .A2(n2514), .ZN(n4026) );
  NAND4_X1 U2626 ( .A1(n2549), .A2(n2548), .A3(n2547), .A4(n2546), .ZN(n3852)
         );
  NAND2_X1 U2627 ( .A1(n2231), .A2(n2533), .ZN(n2979) );
  NAND2_X1 U2628 ( .A1(n2381), .A2(n2916), .ZN(n3871) );
  NAND2_X1 U2629 ( .A1(n2382), .A2(n2262), .ZN(n2381) );
  NAND2_X1 U2630 ( .A1(n4459), .A2(n3889), .ZN(n4470) );
  NAND2_X1 U2631 ( .A1(n4488), .A2(n4489), .ZN(n4487) );
  NAND2_X1 U2632 ( .A1(n4509), .A2(n4510), .ZN(n4508) );
  NAND2_X1 U2633 ( .A1(n4568), .A2(n4570), .ZN(n4569) );
  AND2_X1 U2634 ( .A1(n2918), .A2(n2906), .ZN(n4583) );
  INV_X1 U2635 ( .A(n2390), .ZN(n2389) );
  AOI21_X1 U2636 ( .B1(n2391), .B2(n4581), .A(n4579), .ZN(n2390) );
  NOR2_X1 U2637 ( .A1(n2391), .A2(n4581), .ZN(n4580) );
  AND2_X1 U2638 ( .A1(n4439), .A2(n2958), .ZN(n4585) );
  AOI21_X1 U2639 ( .B1(n3983), .B2(n2361), .A(n2359), .ZN(n2877) );
  NOR2_X1 U2640 ( .A1(n2822), .A2(n2362), .ZN(n2361) );
  INV_X1 U2641 ( .A(n3940), .ZN(n4143) );
  NAND2_X1 U2642 ( .A1(n4717), .A2(n4133), .ZN(n4339) );
  INV_X1 U2643 ( .A(n4404), .ZN(n2912) );
  AND2_X1 U2644 ( .A1(n2472), .A2(n2315), .ZN(n2313) );
  AND2_X1 U2645 ( .A1(n2474), .A2(n2473), .ZN(n2472) );
  AND2_X1 U2646 ( .A1(n2452), .A2(n2233), .ZN(n2306) );
  NOR2_X1 U2647 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2619)
         );
  NOR2_X1 U2648 ( .A1(n3648), .A2(n2444), .ZN(n2443) );
  INV_X1 U2649 ( .A(n3471), .ZN(n2444) );
  OAI21_X1 U2650 ( .B1(n3523), .B2(n3519), .A(n3520), .ZN(n3419) );
  NOR2_X1 U2651 ( .A1(n2303), .A2(n2299), .ZN(n2298) );
  INV_X1 U2652 ( .A(n2453), .ZN(n2299) );
  INV_X1 U2653 ( .A(n2306), .ZN(n2303) );
  NAND2_X1 U2654 ( .A1(n2306), .A2(n2302), .ZN(n2301) );
  INV_X1 U2655 ( .A(n2304), .ZN(n2302) );
  NOR2_X1 U2656 ( .A1(n2279), .A2(n2275), .ZN(n2274) );
  INV_X1 U2657 ( .A(n2708), .ZN(n2275) );
  INV_X1 U2658 ( .A(n2458), .ZN(n2279) );
  AOI21_X1 U2659 ( .B1(n4136), .B2(n2458), .A(n2222), .ZN(n2457) );
  NAND2_X1 U2660 ( .A1(n2458), .A2(n2278), .ZN(n2277) );
  INV_X1 U2661 ( .A(n2709), .ZN(n2278) );
  INV_X1 U2662 ( .A(n3791), .ZN(n2346) );
  AOI21_X1 U2663 ( .B1(n2350), .B2(n3790), .A(n2349), .ZN(n2348) );
  INV_X1 U2664 ( .A(n3776), .ZN(n2350) );
  INV_X1 U2665 ( .A(n3790), .ZN(n2351) );
  NAND2_X1 U2666 ( .A1(n2272), .A2(n2597), .ZN(n3235) );
  NAND2_X1 U2667 ( .A1(n3201), .A2(n3722), .ZN(n2272) );
  NAND2_X1 U2668 ( .A1(n2950), .A2(n4612), .ZN(n3758) );
  NAND2_X1 U2669 ( .A1(n2979), .A2(n4630), .ZN(n3755) );
  NOR2_X1 U2670 ( .A1(n2697), .A2(n2516), .ZN(n3474) );
  INV_X1 U2671 ( .A(IR_REG_27__SCAN_IN), .ZN(n2496) );
  AND2_X1 U2672 ( .A1(n2840), .A2(n2493), .ZN(n2882) );
  AND2_X1 U2673 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2493)
         );
  AND2_X1 U2674 ( .A1(n2475), .A2(n2487), .ZN(n2396) );
  OR2_X1 U2675 ( .A1(n2642), .A2(IR_REG_10__SCAN_IN), .ZN(n2643) );
  OR2_X1 U2676 ( .A1(n2632), .A2(IR_REG_9__SCAN_IN), .ZN(n2642) );
  INV_X1 U2677 ( .A(IR_REG_1__SCAN_IN), .ZN(n2394) );
  NOR2_X1 U2678 ( .A1(n3547), .A2(n3666), .ZN(n2331) );
  NAND2_X1 U2679 ( .A1(n3529), .A2(n3482), .ZN(n3532) );
  INV_X1 U2680 ( .A(n3547), .ZN(n2430) );
  INV_X1 U2681 ( .A(n3594), .ZN(n2427) );
  NAND2_X1 U2682 ( .A1(n2439), .A2(n2438), .ZN(n2437) );
  INV_X1 U2683 ( .A(n3395), .ZN(n2438) );
  INV_X1 U2684 ( .A(n3394), .ZN(n2439) );
  NAND2_X1 U2685 ( .A1(n3394), .A2(n3395), .ZN(n2436) );
  OAI21_X1 U2686 ( .B1(n3575), .B2(n2221), .A(n2237), .ZN(n3614) );
  AND2_X1 U2687 ( .A1(n3489), .A2(n3490), .ZN(n3486) );
  OR2_X1 U2688 ( .A1(n2728), .A2(n4976), .ZN(n2736) );
  NAND2_X1 U2689 ( .A1(n3623), .A2(n2337), .ZN(n2445) );
  AND2_X1 U2690 ( .A1(n2446), .A2(n3627), .ZN(n2337) );
  NAND2_X1 U2691 ( .A1(n2414), .A2(n2230), .ZN(n3337) );
  NAND2_X1 U2692 ( .A1(n3429), .A2(n3606), .ZN(n2322) );
  NAND2_X1 U2693 ( .A1(n3419), .A2(n3418), .ZN(n4423) );
  OR2_X1 U2694 ( .A1(n2655), .A2(n5058), .ZN(n2671) );
  NAND2_X1 U2695 ( .A1(n3871), .A2(n2235), .ZN(n2270) );
  NAND2_X1 U2696 ( .A1(n2966), .A2(REG1_REG_4__SCAN_IN), .ZN(n3910) );
  OAI21_X1 U2697 ( .B1(n3884), .B2(n2268), .A(n2266), .ZN(n3888) );
  INV_X1 U2698 ( .A(n2267), .ZN(n2266) );
  OAI21_X1 U2699 ( .B1(n2228), .B2(n2268), .A(n3887), .ZN(n2267) );
  AOI21_X1 U2700 ( .B1(REG1_REG_5__SCAN_IN), .B2(n3913), .A(n4443), .ZN(n3915)
         );
  AND2_X1 U2701 ( .A1(n2338), .A2(n2261), .ZN(n3918) );
  NAND2_X1 U2702 ( .A1(n4466), .A2(n4463), .ZN(n2338) );
  NAND2_X1 U2703 ( .A1(n4484), .A2(n3920), .ZN(n3921) );
  NAND2_X1 U2704 ( .A1(n4505), .A2(n2253), .ZN(n3923) );
  NAND2_X1 U2705 ( .A1(n4534), .A2(n3925), .ZN(n3927) );
  NAND2_X1 U2706 ( .A1(n4553), .A2(n3929), .ZN(n3931) );
  NAND2_X1 U2707 ( .A1(n3702), .A2(n3818), .ZN(n2362) );
  NOR2_X1 U2708 ( .A1(n2363), .A2(n2360), .ZN(n2359) );
  INV_X1 U2709 ( .A(n3702), .ZN(n2360) );
  INV_X1 U2710 ( .A(n2364), .ZN(n2363) );
  OAI21_X1 U2711 ( .B1(n2220), .B2(n2822), .A(n3704), .ZN(n2364) );
  NAND2_X1 U2712 ( .A1(n2297), .A2(n2300), .ZN(n2874) );
  AND2_X1 U2713 ( .A1(n2301), .A2(n2307), .ZN(n2300) );
  NAND2_X1 U2714 ( .A1(n2454), .A2(n2298), .ZN(n2297) );
  NAND2_X1 U2715 ( .A1(n3844), .A2(n4236), .ZN(n2307) );
  NOR2_X1 U2716 ( .A1(n3967), .A2(n2822), .ZN(n2876) );
  AND2_X1 U2717 ( .A1(n2365), .A2(n2220), .ZN(n3967) );
  NAND2_X1 U2718 ( .A1(n2310), .A2(n2309), .ZN(n4018) );
  NAND2_X1 U2719 ( .A1(n2227), .A2(n2448), .ZN(n2309) );
  NAND2_X1 U2720 ( .A1(n4267), .A2(n3474), .ZN(n2449) );
  INV_X1 U2721 ( .A(n2369), .ZN(n2368) );
  AND2_X1 U2722 ( .A1(n2814), .A2(n2367), .ZN(n2366) );
  AND2_X1 U2723 ( .A1(n2370), .A2(n3803), .ZN(n2369) );
  INV_X1 U2724 ( .A(n3805), .ZN(n2370) );
  NAND2_X1 U2725 ( .A1(n4163), .A2(n4173), .ZN(n2371) );
  NAND2_X1 U2726 ( .A1(n4127), .A2(n2719), .ZN(n4116) );
  OR2_X1 U2727 ( .A1(n4129), .A2(n4136), .ZN(n4127) );
  NAND2_X1 U2728 ( .A1(n2371), .A2(n3803), .ZN(n4147) );
  AOI21_X1 U2729 ( .B1(n2461), .B2(n2462), .A(n2249), .ZN(n2460) );
  INV_X1 U2730 ( .A(n2682), .ZN(n2461) );
  NAND2_X1 U2731 ( .A1(n3366), .A2(n3793), .ZN(n2353) );
  OAI21_X1 U2732 ( .B1(n3366), .B2(n2356), .A(n2354), .ZN(n4206) );
  INV_X1 U2733 ( .A(n2357), .ZN(n2356) );
  AOI21_X1 U2734 ( .B1(n2357), .B2(n2355), .A(n4208), .ZN(n2354) );
  INV_X1 U2735 ( .A(n3793), .ZN(n2355) );
  NOR2_X1 U2736 ( .A1(n2292), .A2(n2247), .ZN(n2289) );
  AND2_X1 U2737 ( .A1(n2635), .A2(REG3_REG_11__SCAN_IN), .ZN(n2645) );
  OAI21_X1 U2738 ( .B1(n2800), .B2(n2351), .A(n2348), .ZN(n4591) );
  NAND2_X1 U2739 ( .A1(n2800), .A2(n3776), .ZN(n3298) );
  AOI21_X1 U2740 ( .B1(n2379), .B2(n2377), .A(n2376), .ZN(n2375) );
  INV_X1 U2741 ( .A(n2379), .ZN(n2378) );
  INV_X1 U2742 ( .A(n3780), .ZN(n2376) );
  OAI21_X1 U2743 ( .B1(n2797), .B2(n2374), .A(n2372), .ZN(n3093) );
  NAND2_X1 U2744 ( .A1(n3766), .A2(n3765), .ZN(n2374) );
  INV_X1 U2745 ( .A(n2282), .ZN(n2281) );
  AND2_X1 U2746 ( .A1(n3768), .A2(n3778), .ZN(n3741) );
  NAND2_X1 U2747 ( .A1(n3068), .A2(n3765), .ZN(n3082) );
  NAND2_X1 U2748 ( .A1(n4617), .A2(n3048), .ZN(n3759) );
  NAND2_X1 U2749 ( .A1(n2796), .A2(n2795), .ZN(n3066) );
  NAND2_X1 U2750 ( .A1(n4609), .A2(n3758), .ZN(n2796) );
  NAND2_X1 U2751 ( .A1(n2797), .A2(n3065), .ZN(n3068) );
  NOR2_X1 U2752 ( .A1(n4695), .A2(n3757), .ZN(n2953) );
  NAND3_X1 U2753 ( .A1(n2352), .A2(n3755), .A3(n3758), .ZN(n4609) );
  NOR2_X1 U2754 ( .A1(n2697), .A2(n4746), .ZN(n4233) );
  INV_X1 U2755 ( .A(n3500), .ZN(n3992) );
  NAND2_X1 U2756 ( .A1(n4077), .A2(n2259), .ZN(n4010) );
  INV_X1 U2757 ( .A(n4023), .ZN(n4029) );
  NAND2_X1 U2758 ( .A1(n4077), .A2(n2408), .ZN(n4031) );
  NAND2_X1 U2759 ( .A1(n4077), .A2(n2409), .ZN(n4046) );
  INV_X1 U2760 ( .A(n3534), .ZN(n4047) );
  NAND2_X1 U2761 ( .A1(n2405), .A2(n2404), .ZN(n2403) );
  NOR2_X1 U2762 ( .A1(n4138), .A2(n3629), .ZN(n2404) );
  INV_X1 U2763 ( .A(n2406), .ZN(n2405) );
  NOR2_X1 U2764 ( .A1(n2697), .A2(n2743), .ZN(n4266) );
  INV_X1 U2765 ( .A(n3541), .ZN(n4118) );
  NOR3_X1 U2766 ( .A1(n4170), .A2(n4138), .A3(n4292), .ZN(n4132) );
  NOR2_X1 U2767 ( .A1(n4170), .A2(n4292), .ZN(n4151) );
  OR2_X1 U2768 ( .A1(n4192), .A2(n4168), .ZN(n4170) );
  NAND2_X1 U2769 ( .A1(n2465), .A2(n2462), .ZN(n4176) );
  NAND2_X1 U2770 ( .A1(n2465), .A2(n2684), .ZN(n4174) );
  NAND2_X1 U2771 ( .A1(n3305), .A2(n2254), .ZN(n4210) );
  INV_X1 U2772 ( .A(n4320), .ZN(n4613) );
  INV_X1 U2773 ( .A(n4317), .ZN(n4616) );
  NAND2_X1 U2774 ( .A1(n3305), .A2(n2400), .ZN(n3360) );
  NAND2_X1 U2775 ( .A1(n3305), .A2(n2401), .ZN(n4603) );
  OAI21_X1 U2776 ( .B1(n3297), .B2(n2246), .A(n2634), .ZN(n4596) );
  AND2_X1 U2777 ( .A1(n3305), .A2(n3314), .ZN(n4685) );
  AND2_X1 U2778 ( .A1(n3119), .A2(n3170), .ZN(n3192) );
  INV_X1 U2779 ( .A(n4333), .ZN(n4625) );
  OR2_X1 U2780 ( .A1(n3078), .A2(n3385), .ZN(n3095) );
  NOR2_X1 U2781 ( .A1(n3095), .A2(n3157), .ZN(n3119) );
  NOR2_X1 U2782 ( .A1(n4628), .A2(n3048), .ZN(n3072) );
  NAND2_X1 U2783 ( .A1(n3072), .A2(n3108), .ZN(n3078) );
  INV_X1 U2784 ( .A(n4328), .ZN(n4611) );
  AND2_X1 U2785 ( .A1(n4413), .A2(n2904), .ZN(n4317) );
  OR2_X1 U2786 ( .A1(n4413), .A2(n2941), .ZN(n4320) );
  OAI21_X1 U2787 ( .B1(n2907), .B2(D_REG_0__SCAN_IN), .A(n2862), .ZN(n3004) );
  AND2_X1 U2788 ( .A1(n2861), .A2(n2860), .ZN(n2868) );
  NAND2_X1 U2789 ( .A1(n2467), .A2(n2466), .ZN(n2314) );
  NOR2_X1 U2790 ( .A1(n2491), .A2(IR_REG_25__SCAN_IN), .ZN(n2315) );
  AND2_X1 U2791 ( .A1(n2792), .A2(n2494), .ZN(n2474) );
  XNOR2_X1 U2792 ( .A(n2846), .B(n2845), .ZN(n3033) );
  XNOR2_X1 U2793 ( .A(n2790), .B(n2789), .ZN(n2829) );
  NAND2_X1 U2794 ( .A1(n2236), .A2(IR_REG_31__SCAN_IN), .ZN(n2790) );
  XNOR2_X1 U2795 ( .A(n2783), .B(n2782), .ZN(n3751) );
  NAND2_X1 U2796 ( .A1(n2232), .A2(IR_REG_31__SCAN_IN), .ZN(n2783) );
  NAND2_X1 U2797 ( .A1(n2786), .A2(IR_REG_31__SCAN_IN), .ZN(n2788) );
  NAND2_X1 U2798 ( .A1(n2727), .A2(IR_REG_31__SCAN_IN), .ZN(n2785) );
  AND3_X1 U2799 ( .A1(n2455), .A2(n2456), .A3(n2486), .ZN(n2706) );
  INV_X1 U2800 ( .A(n2572), .ZN(n2455) );
  OR2_X1 U2801 ( .A1(n2679), .A2(IR_REG_14__SCAN_IN), .ZN(n2680) );
  AOI22_X1 U2802 ( .A1(n2422), .A2(n3205), .B1(n3206), .B2(n2423), .ZN(n2418)
         );
  OR2_X1 U2803 ( .A1(n2423), .A2(n3206), .ZN(n2422) );
  NAND2_X1 U2804 ( .A1(n3028), .A2(n3029), .ZN(n2416) );
  AND2_X1 U2805 ( .A1(n3951), .A2(n2775), .ZN(n3959) );
  INV_X1 U2806 ( .A(n3558), .ZN(n3564) );
  NAND2_X1 U2807 ( .A1(n3623), .A2(n3627), .ZN(n3575) );
  NAND2_X1 U2808 ( .A1(n2435), .A2(n2436), .ZN(n3584) );
  NAND2_X1 U2809 ( .A1(n3396), .A2(n2437), .ZN(n2435) );
  INV_X1 U2810 ( .A(n3672), .ZN(n4421) );
  XOR2_X1 U2811 ( .A(n3139), .B(n3138), .Z(n3382) );
  AOI21_X1 U2812 ( .B1(n2334), .B2(n2336), .A(n2238), .ZN(n2333) );
  INV_X1 U2813 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3650) );
  NAND2_X1 U2814 ( .A1(n2445), .A2(n3471), .ZN(n3647) );
  OR2_X1 U2815 ( .A1(n3149), .A2(n2423), .ZN(n3207) );
  INV_X1 U2816 ( .A(n2447), .ZN(n2975) );
  NAND4_X1 U2817 ( .A1(n2571), .A2(n2570), .A3(n2569), .A4(n2568), .ZN(n3850)
         );
  NAND4_X1 U2818 ( .A1(n2558), .A2(n2557), .A3(n2556), .A4(n2555), .ZN(n3851)
         );
  NAND2_X1 U2819 ( .A1(n2527), .A2(n2526), .ZN(n4614) );
  NOR2_X1 U2820 ( .A1(n2479), .A2(n2522), .ZN(n2527) );
  AND2_X1 U2821 ( .A1(n2525), .A2(n2524), .ZN(n2526) );
  NAND2_X1 U2822 ( .A1(REG2_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2383) );
  XNOR2_X1 U2823 ( .A(n2270), .B(n2923), .ZN(n2962) );
  NAND2_X1 U2824 ( .A1(n3884), .A2(n2228), .ZN(n4449) );
  XNOR2_X1 U2825 ( .A(n3888), .B(n4656), .ZN(n4460) );
  XNOR2_X1 U2826 ( .A(n3918), .B(n2386), .ZN(n4481) );
  NAND2_X1 U2827 ( .A1(n4481), .A2(REG1_REG_8__SCAN_IN), .ZN(n4480) );
  NAND2_X1 U2828 ( .A1(n4475), .A2(n3892), .ZN(n4488) );
  XNOR2_X1 U2829 ( .A(n3921), .B(n2385), .ZN(n4502) );
  NAND2_X1 U2830 ( .A1(n4502), .A2(REG1_REG_10__SCAN_IN), .ZN(n4501) );
  NAND2_X1 U2831 ( .A1(n4496), .A2(n3895), .ZN(n4509) );
  XNOR2_X1 U2832 ( .A(n3923), .B(n2384), .ZN(n4523) );
  NAND2_X1 U2833 ( .A1(n4523), .A2(REG1_REG_12__SCAN_IN), .ZN(n4522) );
  NAND2_X1 U2834 ( .A1(n4517), .A2(n3898), .ZN(n4530) );
  NAND2_X1 U2835 ( .A1(n4535), .A2(n4536), .ZN(n4534) );
  XNOR2_X1 U2836 ( .A(n3927), .B(n4650), .ZN(n4545) );
  NAND2_X1 U2837 ( .A1(n4545), .A2(REG1_REG_14__SCAN_IN), .ZN(n4544) );
  NAND2_X1 U2838 ( .A1(n4554), .A2(n4555), .ZN(n4553) );
  XNOR2_X1 U2839 ( .A(n3931), .B(n3930), .ZN(n4564) );
  NOR2_X1 U2840 ( .A1(n4564), .A2(REG1_REG_16__SCAN_IN), .ZN(n4565) );
  NAND2_X1 U2841 ( .A1(n4560), .A2(n3903), .ZN(n4568) );
  AOI21_X1 U2842 ( .B1(n4583), .B2(ADDR_REG_18__SCAN_IN), .A(n4582), .ZN(n2388) );
  INV_X1 U2843 ( .A(n4528), .ZN(n4579) );
  NAND2_X1 U2844 ( .A1(n2305), .A2(n2304), .ZN(n2308) );
  AND2_X1 U2845 ( .A1(n2305), .A2(n2251), .ZN(n3981) );
  INV_X1 U2846 ( .A(n2450), .ZN(n4063) );
  INV_X1 U2847 ( .A(n4307), .ZN(n4198) );
  OR2_X1 U2848 ( .A1(n3366), .A2(n3794), .ZN(n3346) );
  NAND2_X1 U2849 ( .A1(n2290), .A2(n2295), .ZN(n3358) );
  NAND2_X1 U2850 ( .A1(n3297), .A2(n2291), .ZN(n2290) );
  INV_X1 U2851 ( .A(n2294), .ZN(n2291) );
  NAND2_X1 U2852 ( .A1(n2286), .A2(n2285), .ZN(n3080) );
  NAND2_X1 U2853 ( .A1(n3045), .A2(n2543), .ZN(n3063) );
  AND3_X1 U2854 ( .A1(n2541), .A2(n2540), .A3(n2539), .ZN(n2478) );
  NAND2_X1 U2855 ( .A1(n4618), .A2(n2536), .ZN(n3046) );
  NAND2_X1 U2856 ( .A1(n4172), .A2(n3050), .ZN(n4160) );
  INV_X1 U2857 ( .A(n4171), .ZN(n4627) );
  INV_X1 U2858 ( .A(n4717), .ZN(n4714) );
  OR2_X1 U2859 ( .A1(n4066), .A2(n4065), .ZN(n4369) );
  AND2_X2 U2860 ( .A1(n2868), .A2(n3004), .ZN(n4701) );
  OR2_X1 U2861 ( .A1(n3391), .A2(n2705), .ZN(n2343) );
  INV_X1 U2862 ( .A(n2509), .ZN(n2899) );
  MUX2_X1 U2863 ( .A(IR_REG_31__SCAN_IN), .B(n2839), .S(IR_REG_26__SCAN_IN), 
        .Z(n2841) );
  XNOR2_X1 U2864 ( .A(n2836), .B(IR_REG_24__SCAN_IN), .ZN(n4405) );
  NAND2_X1 U2865 ( .A1(n2835), .A2(IR_REG_31__SCAN_IN), .ZN(n2836) );
  AND2_X1 U2866 ( .A1(n3033), .A2(STATE_REG_SCAN_IN), .ZN(n4643) );
  INV_X1 U2867 ( .A(n2829), .ZN(n4406) );
  INV_X1 U2868 ( .A(n3751), .ZN(n3757) );
  XNOR2_X1 U2869 ( .A(n2694), .B(IR_REG_15__SCAN_IN), .ZN(n4648) );
  NOR2_X1 U2870 ( .A1(n2534), .A2(n2705), .ZN(n2341) );
  INV_X2 U2871 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U2872 ( .A1(n2327), .A2(n4427), .ZN(n2326) );
  NAND2_X1 U2873 ( .A1(n3019), .A2(n3018), .ZN(n3020) );
  NAND2_X1 U2874 ( .A1(n4449), .A2(n4450), .ZN(n4448) );
  NAND2_X1 U2875 ( .A1(n4470), .A2(n4471), .ZN(n4469) );
  INV_X1 U2876 ( .A(n2387), .ZN(n4589) );
  OAI21_X1 U2877 ( .B1(n4580), .B2(n2389), .A(n2388), .ZN(n2387) );
  NAND2_X1 U2878 ( .A1(n2413), .A2(n2411), .ZN(U3354) );
  AOI21_X1 U2879 ( .B1(n3957), .B2(n4191), .A(n2412), .ZN(n2411) );
  OAI21_X1 U2880 ( .B1(n3953), .B2(n3954), .A(n4172), .ZN(n2413) );
  NAND2_X1 U2881 ( .A1(n3955), .A2(n2258), .ZN(n2412) );
  OR2_X1 U2882 ( .A1(n3952), .A2(n4339), .ZN(n2889) );
  OR2_X1 U2883 ( .A1(n3961), .A2(n4339), .ZN(n2866) );
  OR2_X1 U2884 ( .A1(n3952), .A2(n4402), .ZN(n2893) );
  OR2_X1 U2885 ( .A1(n3961), .A2(n4402), .ZN(n2871) );
  INV_X1 U2886 ( .A(n3399), .ZN(n3277) );
  INV_X1 U2887 ( .A(n2932), .ZN(n3550) );
  AND2_X2 U2888 ( .A1(n3034), .A2(n2976), .ZN(n2932) );
  NAND2_X1 U2889 ( .A1(n2845), .A2(n2490), .ZN(n2491) );
  NAND2_X1 U2890 ( .A1(n2454), .A2(n2453), .ZN(n2305) );
  AND2_X1 U2891 ( .A1(n3969), .A2(n3822), .ZN(n2220) );
  OR2_X1 U2892 ( .A1(n2442), .A2(n3472), .ZN(n2221) );
  NAND2_X1 U2893 ( .A1(n4092), .A2(n3730), .ZN(n2222) );
  AND2_X1 U2894 ( .A1(n2431), .A2(n2248), .ZN(n2223) );
  INV_X1 U2895 ( .A(n2697), .ZN(n3709) );
  OR2_X1 U2896 ( .A1(n3845), .A2(n4592), .ZN(n2224) );
  AND2_X1 U2897 ( .A1(n3666), .A2(n3547), .ZN(n2225) );
  AND2_X1 U2898 ( .A1(n2328), .A2(n2255), .ZN(n2226) );
  OR2_X1 U2899 ( .A1(n2250), .A2(n2311), .ZN(n2227) );
  AND2_X1 U2900 ( .A1(n3806), .A2(n3803), .ZN(n4173) );
  INV_X1 U2901 ( .A(n4173), .ZN(n2464) );
  INV_X1 U2902 ( .A(n3678), .ZN(n4427) );
  INV_X1 U2903 ( .A(IR_REG_0__SCAN_IN), .ZN(n2928) );
  NOR2_X1 U2904 ( .A1(n2271), .A2(n2383), .ZN(n3873) );
  OR2_X1 U2905 ( .A1(n3886), .A2(n3885), .ZN(n2228) );
  NAND2_X1 U2906 ( .A1(n2510), .A2(n2509), .ZN(n2553) );
  AND2_X1 U2907 ( .A1(n2353), .A2(n2357), .ZN(n2229) );
  AND2_X1 U2908 ( .A1(n3323), .A2(n3321), .ZN(n2230) );
  AND3_X1 U2909 ( .A1(n2532), .A2(n2530), .A3(n2531), .ZN(n2231) );
  XNOR2_X1 U2910 ( .A(n2343), .B(IR_REG_30__SCAN_IN), .ZN(n2508) );
  OR2_X1 U2911 ( .A1(n2727), .A2(n2489), .ZN(n2232) );
  INV_X1 U2912 ( .A(n4630), .ZN(n4612) );
  OR2_X1 U2913 ( .A1(n3844), .A2(n4236), .ZN(n2233) );
  NOR2_X1 U2914 ( .A1(n2551), .A2(n2287), .ZN(n2234) );
  INV_X1 U2915 ( .A(IR_REG_2__SCAN_IN), .ZN(n2340) );
  OR2_X1 U2916 ( .A1(n3867), .A2(n3869), .ZN(n2235) );
  OR2_X1 U2917 ( .A1(n2727), .A2(n2470), .ZN(n2236) );
  INV_X1 U2918 ( .A(n2491), .ZN(n2466) );
  INV_X1 U2919 ( .A(IR_REG_25__SCAN_IN), .ZN(n2832) );
  AND2_X1 U2920 ( .A1(n2440), .A2(n3486), .ZN(n2237) );
  NOR2_X1 U2921 ( .A1(n2433), .A2(n3405), .ZN(n2238) );
  INV_X1 U2922 ( .A(IR_REG_23__SCAN_IN), .ZN(n2845) );
  AND2_X1 U2923 ( .A1(n2450), .A2(n2449), .ZN(n2239) );
  AND2_X1 U2924 ( .A1(n2308), .A2(n2452), .ZN(n2240) );
  AND2_X1 U2925 ( .A1(n2448), .A2(n4060), .ZN(n2241) );
  AND2_X1 U2926 ( .A1(n2365), .A2(n3822), .ZN(n2242) );
  AND2_X1 U2927 ( .A1(n2344), .A2(n2315), .ZN(n2243) );
  OR2_X1 U2928 ( .A1(n2314), .A2(n2727), .ZN(n2244) );
  INV_X1 U2929 ( .A(IR_REG_28__SCAN_IN), .ZN(n2792) );
  AND2_X1 U2930 ( .A1(n4595), .A2(n3401), .ZN(n2245) );
  AND2_X1 U2931 ( .A1(n4593), .A2(n3327), .ZN(n2246) );
  NAND2_X1 U2932 ( .A1(n2321), .A2(n3430), .ZN(n3607) );
  NAND2_X1 U2933 ( .A1(n3337), .A2(n3336), .ZN(n3396) );
  AND2_X1 U2934 ( .A1(n4331), .A2(n3586), .ZN(n2247) );
  INV_X1 U2935 ( .A(n3639), .ZN(n4327) );
  OR2_X1 U2936 ( .A1(n3499), .A2(n3498), .ZN(n2248) );
  AND2_X1 U2937 ( .A1(n4308), .A2(n4168), .ZN(n2249) );
  INV_X1 U2938 ( .A(IR_REG_29__SCAN_IN), .ZN(n2473) );
  AND2_X1 U2939 ( .A1(n4055), .A2(n3534), .ZN(n2250) );
  NAND2_X1 U2940 ( .A1(n2414), .A2(n3321), .ZN(n3322) );
  NAND2_X1 U2941 ( .A1(n4026), .A2(n3596), .ZN(n2251) );
  AND2_X1 U2942 ( .A1(n2371), .A2(n2369), .ZN(n2252) );
  INV_X1 U2943 ( .A(n3420), .ZN(n4422) );
  INV_X1 U2944 ( .A(n2402), .ZN(n4120) );
  NOR3_X1 U2945 ( .A1(n4170), .A2(n2406), .A3(n4138), .ZN(n2402) );
  NOR2_X1 U2946 ( .A1(n4170), .A2(n2403), .ZN(n2407) );
  OR2_X1 U2947 ( .A1(n4653), .A2(n4715), .ZN(n2253) );
  AND2_X1 U2948 ( .A1(n2400), .A2(n4327), .ZN(n2254) );
  NAND2_X1 U2949 ( .A1(n3547), .A2(n2428), .ZN(n2255) );
  NAND2_X1 U2950 ( .A1(n2296), .A2(n4597), .ZN(n2256) );
  AND2_X1 U2951 ( .A1(n3667), .A2(n2248), .ZN(n2428) );
  INV_X1 U2952 ( .A(n2428), .ZN(n2329) );
  AND2_X1 U2953 ( .A1(n2322), .A2(n3605), .ZN(n2257) );
  INV_X1 U2954 ( .A(n2463), .ZN(n2462) );
  NAND2_X1 U2955 ( .A1(n2464), .A2(n2684), .ZN(n2463) );
  NAND2_X2 U2956 ( .A1(n3007), .A2(n4171), .ZN(n4172) );
  INV_X1 U2957 ( .A(n4138), .ZN(n4135) );
  AND2_X1 U2958 ( .A1(n2508), .A2(n2899), .ZN(n2537) );
  OAI22_X1 U2959 ( .A1(n3235), .A2(n2608), .B1(n3265), .B2(n3847), .ZN(n3224)
         );
  OAI21_X1 U2960 ( .B1(n3117), .B2(n2585), .A(n2584), .ZN(n3201) );
  NOR2_X1 U2961 ( .A1(n2697), .A2(n2499), .ZN(n3596) );
  INV_X1 U2962 ( .A(n3786), .ZN(n2349) );
  OR2_X1 U2963 ( .A1(n4221), .A2(n3956), .ZN(n2258) );
  NAND2_X1 U2964 ( .A1(n2451), .A2(n4618), .ZN(n3045) );
  AND2_X1 U2965 ( .A1(n2408), .A2(n4011), .ZN(n2259) );
  NOR2_X1 U2966 ( .A1(n3149), .A2(n3148), .ZN(n2260) );
  INV_X1 U2967 ( .A(n2410), .ZN(n2409) );
  NAND2_X1 U2968 ( .A1(n4047), .A2(n4064), .ZN(n2410) );
  NAND2_X1 U2969 ( .A1(n2397), .A2(n2475), .ZN(n2572) );
  INV_X1 U2970 ( .A(n3721), .ZN(n2284) );
  INV_X1 U2971 ( .A(n4236), .ZN(n3976) );
  NOR2_X1 U2972 ( .A1(n2697), .A2(n2773), .ZN(n4236) );
  NAND2_X1 U2973 ( .A1(n2986), .A2(n2985), .ZN(n3019) );
  INV_X1 U2974 ( .A(n4495), .ZN(n2385) );
  INV_X1 U2975 ( .A(n4516), .ZN(n2384) );
  INV_X1 U2976 ( .A(n4474), .ZN(n2386) );
  INV_X1 U2977 ( .A(IR_REG_3__SCAN_IN), .ZN(n2559) );
  INV_X1 U2978 ( .A(DATAI_1_), .ZN(n2399) );
  INV_X1 U2979 ( .A(IR_REG_22__SCAN_IN), .ZN(n2789) );
  INV_X1 U2980 ( .A(IR_REG_19__SCAN_IN), .ZN(n2784) );
  OR2_X1 U2981 ( .A1(n3917), .A2(REG1_REG_7__SCAN_IN), .ZN(n2261) );
  OR2_X1 U2982 ( .A1(n3859), .A2(n2915), .ZN(n2262) );
  INV_X1 U2983 ( .A(n2312), .ZN(n3391) );
  MUX2_X1 U2984 ( .A(REG2_REG_1__SCAN_IN), .B(n2915), .S(n3859), .Z(n2271) );
  NAND3_X1 U2985 ( .A1(n2395), .A2(n2393), .A3(n2535), .ZN(n3859) );
  INV_X1 U2986 ( .A(n2979), .ZN(n2950) );
  NAND2_X1 U2987 ( .A1(n4150), .A2(n2274), .ZN(n2273) );
  NAND2_X1 U2988 ( .A1(n2273), .A2(n2276), .ZN(n2734) );
  NAND2_X1 U2989 ( .A1(n2283), .A2(n2281), .ZN(n3100) );
  OAI21_X1 U2990 ( .B1(n2285), .B2(n2284), .A(n2563), .ZN(n2282) );
  NAND3_X1 U2991 ( .A1(n2234), .A2(n3045), .A3(n3721), .ZN(n2283) );
  NAND2_X1 U2992 ( .A1(n2234), .A2(n3045), .ZN(n2286) );
  NAND2_X1 U2993 ( .A1(n3297), .A2(n2293), .ZN(n2288) );
  NAND2_X1 U2994 ( .A1(n2288), .A2(n2289), .ZN(n3349) );
  NAND2_X1 U2995 ( .A1(n4061), .A2(n2241), .ZN(n2310) );
  NAND4_X1 U2996 ( .A1(n2467), .A2(n2316), .A3(n2344), .A4(n2313), .ZN(n2312)
         );
  NAND2_X1 U2997 ( .A1(n2319), .A2(n2257), .ZN(n3656) );
  NAND3_X1 U2998 ( .A1(n3428), .A2(n2320), .A3(n4422), .ZN(n2319) );
  NAND3_X1 U2999 ( .A1(n3428), .A2(n4422), .A3(n4425), .ZN(n2321) );
  INV_X1 U3000 ( .A(n4405), .ZN(n2908) );
  NAND2_X4 U3001 ( .A1(n3008), .A2(n3034), .ZN(n3551) );
  INV_X1 U3002 ( .A(n2911), .ZN(n2323) );
  NAND2_X1 U3003 ( .A1(n2431), .A2(n2325), .ZN(n2324) );
  OAI211_X1 U3004 ( .C1(n2431), .C2(n2326), .A(n3518), .B(n2324), .ZN(U3211)
         );
  NAND2_X1 U3005 ( .A1(n2414), .A2(n2334), .ZN(n2332) );
  NAND2_X1 U3006 ( .A1(n2332), .A2(n2333), .ZN(n3635) );
  NAND2_X1 U3007 ( .A1(n2445), .A2(n2443), .ZN(n3529) );
  XNOR2_X2 U3008 ( .A(n2341), .B(n2340), .ZN(n4410) );
  NAND3_X1 U3009 ( .A1(n2344), .A2(n2456), .A3(n2396), .ZN(n2716) );
  NAND2_X1 U3010 ( .A1(n2800), .A2(n2348), .ZN(n2347) );
  INV_X1 U3011 ( .A(n3754), .ZN(n2352) );
  NAND2_X1 U3012 ( .A1(n3983), .A2(n3818), .ZN(n2365) );
  OAI21_X1 U3013 ( .B1(n4163), .B2(n2368), .A(n2366), .ZN(n2815) );
  INV_X1 U3014 ( .A(n2373), .ZN(n2372) );
  OAI21_X1 U3015 ( .B1(n2374), .B2(n3065), .A(n3769), .ZN(n2373) );
  OAI21_X1 U3016 ( .B1(n3196), .B2(n2378), .A(n2375), .ZN(n3222) );
  OAI21_X1 U3017 ( .B1(n3196), .B2(n2799), .A(n3781), .ZN(n3236) );
  AOI21_X1 U3018 ( .B1(n2799), .B2(n3781), .A(n2380), .ZN(n2379) );
  AOI211_X1 U3019 ( .C1(n3957), .C2(n4678), .A(n3954), .B(n2886), .ZN(n2891)
         );
  NAND2_X1 U3020 ( .A1(n2815), .A2(n3809), .ZN(n4074) );
  NAND2_X4 U3021 ( .A1(n2498), .A2(n2398), .ZN(n2697) );
  NAND2_X1 U3022 ( .A1(n3317), .A2(n3316), .ZN(n2414) );
  NAND2_X1 U3024 ( .A1(n3254), .A2(n3253), .ZN(n3274) );
  NAND2_X1 U3025 ( .A1(n2419), .A2(n2418), .ZN(n3250) );
  INV_X1 U3026 ( .A(n3873), .ZN(n2382) );
  NAND3_X1 U3027 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .A3(
        IR_REG_31__SCAN_IN), .ZN(n2395) );
  MUX2_X1 U3028 ( .A(n2399), .B(n3859), .S(n2697), .Z(n4630) );
  INV_X1 U3029 ( .A(n2407), .ZN(n4095) );
  INV_X1 U3030 ( .A(n3021), .ZN(n2415) );
  NAND3_X1 U3031 ( .A1(n3019), .A2(n3018), .A3(n2415), .ZN(n2417) );
  INV_X1 U3032 ( .A(n2417), .ZN(n3027) );
  NAND2_X1 U3033 ( .A1(n3149), .A2(n2420), .ZN(n2419) );
  NOR2_X1 U3034 ( .A1(n3167), .A2(n3168), .ZN(n2424) );
  NAND2_X1 U3035 ( .A1(n3593), .A2(n3594), .ZN(n2431) );
  INV_X1 U3036 ( .A(n3472), .ZN(n2446) );
  NAND2_X2 U3037 ( .A1(n2447), .A2(n2976), .ZN(n3399) );
  NOR2_X1 U3038 ( .A1(n2572), .A2(n2483), .ZN(n2661) );
  OAI21_X1 U3039 ( .B1(n4187), .B2(n2463), .A(n2460), .ZN(n4150) );
  NAND2_X1 U3040 ( .A1(n2495), .A2(n2474), .ZN(n2507) );
  NAND2_X1 U3041 ( .A1(n2495), .A2(n2494), .ZN(n2506) );
  XNOR2_X1 U3042 ( .A(n3017), .B(n2980), .ZN(n2986) );
  XNOR2_X1 U3043 ( .A(n2977), .B(n3399), .ZN(n3017) );
  AOI21_X1 U3044 ( .B1(n2979), .B2(n3479), .A(n2974), .ZN(n2977) );
  INV_X2 U3045 ( .A(n4172), .ZN(n4626) );
  INV_X1 U3046 ( .A(DATAI_25_), .ZN(n2499) );
  AND2_X1 U3047 ( .A1(n3565), .A2(n4427), .ZN(n2476) );
  AND2_X1 U3048 ( .A1(n3557), .A2(n2476), .ZN(n2477) );
  INV_X1 U3049 ( .A(DATAI_27_), .ZN(n2773) );
  INV_X1 U3050 ( .A(DATAI_21_), .ZN(n2743) );
  AND2_X1 U3051 ( .A1(n3706), .A2(REG2_REG_0__SCAN_IN), .ZN(n2479) );
  INV_X1 U3052 ( .A(n3581), .ZN(n3406) );
  AND2_X1 U3053 ( .A1(n4186), .A2(n2683), .ZN(n2681) );
  AND2_X1 U3054 ( .A1(n4208), .A2(n2681), .ZN(n2682) );
  INV_X1 U3055 ( .A(IR_REG_24__SCAN_IN), .ZN(n2490) );
  INV_X1 U3056 ( .A(IR_REG_17__SCAN_IN), .ZN(n2487) );
  INV_X1 U3057 ( .A(n3582), .ZN(n3405) );
  INV_X1 U3058 ( .A(n3325), .ZN(n3323) );
  INV_X1 U3059 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4976) );
  INV_X1 U3060 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4839) );
  INV_X1 U3061 ( .A(DATAI_22_), .ZN(n2516) );
  INV_X1 U3062 ( .A(IR_REG_13__SCAN_IN), .ZN(n2669) );
  OAI21_X1 U3063 ( .B1(n3635), .B2(n3637), .A(n3636), .ZN(n3408) );
  INV_X1 U3064 ( .A(REG3_REG_10__SCAN_IN), .ZN(n5045) );
  OR2_X1 U3065 ( .A1(n3252), .A2(n3251), .ZN(n3253) );
  NAND2_X1 U3066 ( .A1(n3144), .A2(n3150), .ZN(n3145) );
  NOR2_X1 U3067 ( .A1(n2907), .A2(D_REG_1__SCAN_IN), .ZN(n3003) );
  OR2_X1 U3068 ( .A1(n2738), .A2(n3650), .ZN(n2747) );
  OR2_X1 U3069 ( .A1(n2754), .A2(n4839), .ZN(n2760) );
  OR2_X1 U3070 ( .A1(n2710), .A2(n4578), .ZN(n2721) );
  OR2_X1 U3071 ( .A1(n2612), .A2(n2500), .ZN(n2626) );
  INV_X1 U3072 ( .A(n3179), .ZN(n3170) );
  NAND2_X1 U3073 ( .A1(n3759), .A2(n3761), .ZN(n2794) );
  INV_X1 U3074 ( .A(DATAI_20_), .ZN(n4978) );
  INV_X1 U3075 ( .A(n4592), .ZN(n4604) );
  INV_X1 U3076 ( .A(IR_REG_21__SCAN_IN), .ZN(n2782) );
  INV_X1 U3077 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3515) );
  INV_X1 U3078 ( .A(DATAI_23_), .ZN(n2753) );
  INV_X1 U3079 ( .A(n3168), .ZN(n3143) );
  AND2_X1 U3080 ( .A1(n2954), .A2(n4171), .ZN(n4416) );
  NOR2_X1 U3081 ( .A1(n3551), .A2(n2948), .ZN(n3836) );
  INV_X1 U3082 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3172) );
  INV_X1 U3083 ( .A(REG3_REG_13__SCAN_IN), .ZN(n5058) );
  INV_X1 U3084 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4578) );
  AND2_X1 U3085 ( .A1(n3701), .A2(n3821), .ZN(n3969) );
  AND2_X1 U3086 ( .A1(n4107), .A2(n4106), .ZN(n4149) );
  NAND2_X1 U3087 ( .A1(n3001), .A2(n2953), .ZN(n4171) );
  NOR2_X1 U3088 ( .A1(n2697), .A2(n4879), .ZN(n3500) );
  NOR2_X1 U3089 ( .A1(n2697), .A2(n4978), .ZN(n3629) );
  AND2_X1 U3090 ( .A1(n2824), .A2(n2823), .ZN(n4333) );
  NAND2_X1 U3091 ( .A1(n2834), .A2(n2838), .ZN(n2911) );
  NOR2_X1 U3092 ( .A1(n2697), .A2(n2753), .ZN(n3534) );
  INV_X1 U3093 ( .A(n4416), .ZN(n3682) );
  INV_X1 U3094 ( .A(n4417), .ZN(n3681) );
  OR2_X1 U3095 ( .A1(n2774), .A2(n3560), .ZN(n3951) );
  AND2_X1 U3096 ( .A1(n2918), .A2(n2917), .ZN(n4439) );
  AND2_X1 U3097 ( .A1(n4439), .A2(n3835), .ZN(n4528) );
  AND2_X1 U3098 ( .A1(n4109), .A2(n4110), .ZN(n4136) );
  INV_X1 U3099 ( .A(n4208), .ZN(n4205) );
  AND2_X1 U3100 ( .A1(n3797), .A2(n3347), .ZN(n3738) );
  AND2_X1 U3101 ( .A1(n4172), .A2(n3102), .ZN(n4191) );
  INV_X1 U3102 ( .A(n4160), .ZN(n4632) );
  INV_X1 U3103 ( .A(n4694), .ZN(n4133) );
  NAND2_X1 U3104 ( .A1(n4621), .A2(n4695), .ZN(n4678) );
  INV_X1 U3105 ( .A(n4695), .ZN(n4689) );
  AND2_X1 U3106 ( .A1(n3034), .A2(n4643), .ZN(n3001) );
  INV_X1 U3107 ( .A(n4643), .ZN(n2895) );
  NAND2_X1 U3108 ( .A1(n3558), .A2(n2477), .ZN(n3571) );
  AND2_X1 U3109 ( .A1(n3038), .A2(n3037), .ZN(n4432) );
  OR2_X1 U3110 ( .A1(n2989), .A2(n2944), .ZN(n3678) );
  INV_X1 U3111 ( .A(n4240), .ZN(n3972) );
  OR2_X1 U3112 ( .A1(n2758), .A2(n2757), .ZN(n4007) );
  INV_X2 U3113 ( .A(U4043), .ZN(n3854) );
  NAND2_X1 U3114 ( .A1(n4439), .A2(n4413), .ZN(n4590) );
  INV_X1 U3115 ( .A(n4191), .ZN(n4177) );
  INV_X1 U3116 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4715) );
  AND2_X2 U3117 ( .A1(n2868), .A2(n2863), .ZN(n4717) );
  NAND2_X1 U3118 ( .A1(n4701), .A2(n4133), .ZN(n4402) );
  INV_X1 U3119 ( .A(n4701), .ZN(n4699) );
  INV_X1 U3120 ( .A(D_REG_23__SCAN_IN), .ZN(n5034) );
  INV_X1 U3121 ( .A(D_REG_7__SCAN_IN), .ZN(n5017) );
  INV_X1 U3122 ( .A(DATAI_30_), .ZN(n4746) );
  INV_X1 U3123 ( .A(n3908), .ZN(n4653) );
  NOR2_X1 U3124 ( .A1(n3034), .A2(n2895), .ZN(U4043) );
  INV_X1 U3125 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2864) );
  NAND2_X1 U3126 ( .A1(n2534), .A2(n2340), .ZN(n2550) );
  NAND4_X1 U3127 ( .A1(n2619), .A2(n2482), .A3(n2481), .A4(n2480), .ZN(n2483)
         );
  NAND2_X1 U3128 ( .A1(n2787), .A2(n2784), .ZN(n2489) );
  NAND2_X1 U3129 ( .A1(n2705), .A2(n2496), .ZN(n2497) );
  NAND2_X1 U3130 ( .A1(n2506), .A2(n2497), .ZN(n2883) );
  NAND2_X1 U3131 ( .A1(n2883), .A2(n2792), .ZN(n2498) );
  NAND2_X1 U3132 ( .A1(n2564), .A2(REG3_REG_5__SCAN_IN), .ZN(n2577) );
  NOR2_X1 U3133 ( .A1(n2577), .A2(n3172), .ZN(n2588) );
  NAND2_X1 U3134 ( .A1(n2588), .A2(REG3_REG_7__SCAN_IN), .ZN(n2612) );
  NAND2_X1 U3135 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2500) );
  NOR2_X1 U3136 ( .A1(n2626), .A2(n5045), .ZN(n2635) );
  NAND2_X1 U3137 ( .A1(n2645), .A2(REG3_REG_12__SCAN_IN), .ZN(n2655) );
  NAND2_X1 U3138 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2501) );
  NOR2_X1 U3139 ( .A1(n2671), .A2(n2501), .ZN(n2685) );
  NAND2_X1 U3140 ( .A1(n2685), .A2(REG3_REG_16__SCAN_IN), .ZN(n2699) );
  INV_X1 U3141 ( .A(n2699), .ZN(n2502) );
  NAND2_X1 U3142 ( .A1(n2502), .A2(REG3_REG_17__SCAN_IN), .ZN(n2710) );
  INV_X1 U3143 ( .A(n2721), .ZN(n2503) );
  NAND2_X1 U3144 ( .A1(n2503), .A2(REG3_REG_19__SCAN_IN), .ZN(n2728) );
  INV_X1 U3145 ( .A(n2736), .ZN(n2504) );
  NAND2_X1 U3146 ( .A1(n2504), .A2(REG3_REG_21__SCAN_IN), .ZN(n2738) );
  INV_X1 U3147 ( .A(n2747), .ZN(n2505) );
  NAND2_X1 U31480 ( .A1(n2505), .A2(REG3_REG_23__SCAN_IN), .ZN(n2754) );
  XNOR2_X1 U31490 ( .A(n2760), .B(REG3_REG_25__SCAN_IN), .ZN(n4013) );
  NAND2_X1 U3150 ( .A1(n4013), .A2(n2537), .ZN(n2515) );
  INV_X1 U3151 ( .A(n2508), .ZN(n2510) );
  AND2_X2 U3152 ( .A1(n2510), .A2(n2899), .ZN(n2538) );
  INV_X1 U3153 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4251) );
  NAND2_X1 U3154 ( .A1(n3706), .A2(REG2_REG_25__SCAN_IN), .ZN(n2512) );
  NAND2_X1 U3155 ( .A1(n2544), .A2(REG0_REG_25__SCAN_IN), .ZN(n2511) );
  OAI211_X1 U3156 ( .C1(n2566), .C2(n4251), .A(n2512), .B(n2511), .ZN(n2513)
         );
  INV_X1 U3157 ( .A(n2513), .ZN(n2514) );
  INV_X1 U3158 ( .A(n4026), .ZN(n3671) );
  INV_X1 U3159 ( .A(n3596), .ZN(n4011) );
  NAND2_X1 U3160 ( .A1(n2544), .A2(REG0_REG_22__SCAN_IN), .ZN(n2521) );
  NAND2_X1 U3161 ( .A1(n2738), .A2(n3650), .ZN(n2517) );
  NAND2_X1 U3162 ( .A1(n2747), .A2(n2517), .ZN(n3649) );
  OR2_X1 U3163 ( .A1(n2828), .A2(n3649), .ZN(n2520) );
  NAND2_X1 U3164 ( .A1(n2538), .A2(REG1_REG_22__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U3165 ( .A1(n3706), .A2(REG2_REG_22__SCAN_IN), .ZN(n2518) );
  NAND4_X1 U3166 ( .A1(n2521), .A2(n2520), .A3(n2519), .A4(n2518), .ZN(n4267)
         );
  INV_X1 U3167 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2523) );
  OR2_X1 U3168 ( .A1(n2553), .A2(n2523), .ZN(n2525) );
  NAND2_X1 U3169 ( .A1(n2538), .A2(REG1_REG_0__SCAN_IN), .ZN(n2524) );
  INV_X1 U3170 ( .A(DATAI_0_), .ZN(n2528) );
  MUX2_X1 U3171 ( .A(n2528), .B(n2928), .S(n2697), .Z(n4629) );
  NOR2_X1 U3172 ( .A1(n2990), .A2(n4629), .ZN(n4619) );
  NAND2_X1 U3173 ( .A1(n2537), .A2(REG3_REG_1__SCAN_IN), .ZN(n2533) );
  INV_X1 U3174 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2529) );
  OR2_X1 U3175 ( .A1(n2553), .A2(n2529), .ZN(n2532) );
  NAND2_X1 U3176 ( .A1(n2538), .A2(REG1_REG_1__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U3177 ( .A1(n3706), .A2(REG2_REG_1__SCAN_IN), .ZN(n2530) );
  INV_X1 U3178 ( .A(n2534), .ZN(n2535) );
  INV_X1 U3179 ( .A(n3859), .ZN(n4411) );
  NAND2_X1 U3180 ( .A1(n4619), .A2(n4620), .ZN(n4618) );
  NAND2_X1 U3181 ( .A1(n2979), .A2(n4612), .ZN(n2536) );
  INV_X1 U3182 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3051) );
  OR2_X1 U3183 ( .A1(n2828), .A2(n3051), .ZN(n2542) );
  NAND2_X1 U3184 ( .A1(n2544), .A2(REG0_REG_2__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U3185 ( .A1(n3706), .A2(REG2_REG_2__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U3186 ( .A1(n2538), .A2(REG1_REG_2__SCAN_IN), .ZN(n2539) );
  MUX2_X1 U3187 ( .A(DATAI_2_), .B(n4410), .S(n2697), .Z(n3048) );
  INV_X1 U3188 ( .A(n3048), .ZN(n3055) );
  NAND2_X1 U3189 ( .A1(n3853), .A2(n3055), .ZN(n3761) );
  NAND2_X1 U3190 ( .A1(n4617), .A2(n3055), .ZN(n2543) );
  OR2_X1 U3191 ( .A1(n2828), .A2(REG3_REG_3__SCAN_IN), .ZN(n2549) );
  INV_X1 U3192 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2545) );
  OR2_X1 U3193 ( .A1(n2553), .A2(n2545), .ZN(n2548) );
  NAND2_X1 U3194 ( .A1(n2538), .A2(REG1_REG_3__SCAN_IN), .ZN(n2547) );
  NAND2_X1 U3195 ( .A1(n3706), .A2(REG2_REG_3__SCAN_IN), .ZN(n2546) );
  NAND2_X1 U3196 ( .A1(n2550), .A2(IR_REG_31__SCAN_IN), .ZN(n2560) );
  XNOR2_X1 U3197 ( .A(n2560), .B(IR_REG_3__SCAN_IN), .ZN(n4409) );
  MUX2_X1 U3198 ( .A(DATAI_3_), .B(n4409), .S(n2697), .Z(n3763) );
  NOR2_X1 U3199 ( .A1(n3852), .A2(n3763), .ZN(n2551) );
  INV_X1 U3200 ( .A(n3852), .ZN(n3764) );
  INV_X1 U3201 ( .A(n3763), .ZN(n3108) );
  INV_X1 U3202 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2552) );
  OR2_X1 U3203 ( .A1(n2553), .A2(n2552), .ZN(n2558) );
  NAND2_X1 U3204 ( .A1(n2538), .A2(REG1_REG_4__SCAN_IN), .ZN(n2557) );
  NOR2_X1 U3205 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2554) );
  NOR2_X1 U3206 ( .A1(n2564), .A2(n2554), .ZN(n3383) );
  NAND2_X1 U3207 ( .A1(n2537), .A2(n3383), .ZN(n2556) );
  NAND2_X1 U3208 ( .A1(n3706), .A2(REG2_REG_4__SCAN_IN), .ZN(n2555) );
  INV_X1 U3209 ( .A(n3851), .ZN(n3160) );
  NAND2_X1 U32100 ( .A1(n2560), .A2(n2559), .ZN(n2561) );
  NAND2_X1 U32110 ( .A1(n2561), .A2(IR_REG_31__SCAN_IN), .ZN(n2562) );
  XNOR2_X1 U32120 ( .A(n2562), .B(IR_REG_4__SCAN_IN), .ZN(n4408) );
  MUX2_X1 U32130 ( .A(DATAI_4_), .B(n4408), .S(n2697), .Z(n3385) );
  NAND2_X1 U32140 ( .A1(n3160), .A2(n3385), .ZN(n3766) );
  INV_X1 U32150 ( .A(n3385), .ZN(n3133) );
  NAND2_X1 U32160 ( .A1(n3851), .A2(n3133), .ZN(n3769) );
  NAND2_X1 U32170 ( .A1(n3766), .A2(n3769), .ZN(n3721) );
  NAND2_X1 U32180 ( .A1(n3851), .A2(n3385), .ZN(n2563) );
  OAI21_X1 U32190 ( .B1(n2564), .B2(REG3_REG_5__SCAN_IN), .A(n2577), .ZN(n3156) );
  OR2_X1 U32200 ( .A1(n2828), .A2(n3156), .ZN(n2571) );
  INV_X2 U32210 ( .A(n2538), .ZN(n2566) );
  INV_X1 U32220 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2565) );
  OR2_X1 U32230 ( .A1(n2566), .A2(n2565), .ZN(n2570) );
  INV_X1 U32240 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2567) );
  OR2_X1 U32250 ( .A1(n2772), .A2(n2567), .ZN(n2569) );
  NAND2_X1 U32260 ( .A1(n2544), .A2(REG0_REG_5__SCAN_IN), .ZN(n2568) );
  NAND2_X1 U32270 ( .A1(n2572), .A2(IR_REG_31__SCAN_IN), .ZN(n2573) );
  XNOR2_X1 U32280 ( .A(n2573), .B(IR_REG_5__SCAN_IN), .ZN(n3913) );
  MUX2_X1 U32290 ( .A(DATAI_5_), .B(n3913), .S(n2697), .Z(n3157) );
  AND2_X1 U32300 ( .A1(n3850), .A2(n3157), .ZN(n2574) );
  INV_X1 U32310 ( .A(n3850), .ZN(n3181) );
  INV_X1 U32320 ( .A(n3157), .ZN(n3152) );
  NAND2_X1 U32330 ( .A1(n3181), .A2(n3152), .ZN(n2575) );
  INV_X1 U32340 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2576) );
  OR2_X1 U32350 ( .A1(n2553), .A2(n2576), .ZN(n2582) );
  INV_X2 U32360 ( .A(n2537), .ZN(n2828) );
  AND2_X1 U32370 ( .A1(n2577), .A2(n3172), .ZN(n2578) );
  OR2_X1 U32380 ( .A1(n2578), .A2(n2588), .ZN(n3175) );
  OR2_X1 U32390 ( .A1(n2828), .A2(n3175), .ZN(n2581) );
  NAND2_X1 U32400 ( .A1(n2538), .A2(REG1_REG_6__SCAN_IN), .ZN(n2580) );
  NAND2_X1 U32410 ( .A1(n3706), .A2(REG2_REG_6__SCAN_IN), .ZN(n2579) );
  NAND4_X1 U32420 ( .A1(n2582), .A2(n2581), .A3(n2580), .A4(n2579), .ZN(n3849)
         );
  NOR2_X1 U32430 ( .A1(n2572), .A2(IR_REG_5__SCAN_IN), .ZN(n2621) );
  OR2_X1 U32440 ( .A1(n2621), .A2(n2705), .ZN(n2583) );
  XNOR2_X1 U32450 ( .A(n2583), .B(IR_REG_6__SCAN_IN), .ZN(n3914) );
  MUX2_X1 U32460 ( .A(DATAI_6_), .B(n3914), .S(n2697), .Z(n3179) );
  NOR2_X1 U32470 ( .A1(n3849), .A2(n3179), .ZN(n2585) );
  NAND2_X1 U32480 ( .A1(n3849), .A2(n3179), .ZN(n2584) );
  INV_X1 U32490 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2586) );
  OR2_X1 U32500 ( .A1(n2553), .A2(n2586), .ZN(n2594) );
  INV_X1 U32510 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2587) );
  OR2_X1 U32520 ( .A1(n2566), .A2(n2587), .ZN(n2593) );
  OR2_X1 U32530 ( .A1(n2588), .A2(REG3_REG_7__SCAN_IN), .ZN(n2589) );
  NAND2_X1 U32540 ( .A1(n2612), .A2(n2589), .ZN(n3216) );
  OR2_X1 U32550 ( .A1(n2828), .A2(n3216), .ZN(n2592) );
  INV_X1 U32560 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2590) );
  OR2_X1 U32570 ( .A1(n2772), .A2(n2590), .ZN(n2591) );
  NAND4_X1 U32580 ( .A1(n2594), .A2(n2593), .A3(n2592), .A4(n2591), .ZN(n3848)
         );
  INV_X1 U32590 ( .A(n3848), .ZN(n3238) );
  INV_X1 U32600 ( .A(IR_REG_6__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U32610 ( .A1(n2621), .A2(n2595), .ZN(n2596) );
  NAND2_X1 U32620 ( .A1(n2596), .A2(IR_REG_31__SCAN_IN), .ZN(n2605) );
  XNOR2_X1 U32630 ( .A(n2605), .B(IR_REG_7__SCAN_IN), .ZN(n3917) );
  MUX2_X1 U32640 ( .A(DATAI_7_), .B(n3917), .S(n2697), .Z(n3213) );
  NAND2_X1 U32650 ( .A1(n3238), .A2(n3213), .ZN(n3772) );
  INV_X1 U32660 ( .A(n3213), .ZN(n3210) );
  NAND2_X1 U32670 ( .A1(n3848), .A2(n3210), .ZN(n3781) );
  NAND2_X1 U32680 ( .A1(n3772), .A2(n3781), .ZN(n3722) );
  NAND2_X1 U32690 ( .A1(n3848), .A2(n3213), .ZN(n2597) );
  INV_X1 U32700 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2598) );
  OR2_X1 U32710 ( .A1(n2553), .A2(n2598), .ZN(n2603) );
  INV_X1 U32720 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2599) );
  OR2_X1 U32730 ( .A1(n2566), .A2(n2599), .ZN(n2602) );
  INV_X1 U32740 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2611) );
  XNOR2_X1 U32750 ( .A(n2612), .B(n2611), .ZN(n3268) );
  OR2_X1 U32760 ( .A1(n2828), .A2(n3268), .ZN(n2601) );
  INV_X1 U32770 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3244) );
  OR2_X1 U32780 ( .A1(n2772), .A2(n3244), .ZN(n2600) );
  NAND4_X1 U32790 ( .A1(n2603), .A2(n2602), .A3(n2601), .A4(n2600), .ZN(n3847)
         );
  INV_X1 U32800 ( .A(IR_REG_7__SCAN_IN), .ZN(n2604) );
  NAND2_X1 U32810 ( .A1(n2605), .A2(n2604), .ZN(n2606) );
  NAND2_X1 U32820 ( .A1(n2606), .A2(IR_REG_31__SCAN_IN), .ZN(n2607) );
  XNOR2_X1 U32830 ( .A(n2607), .B(IR_REG_8__SCAN_IN), .ZN(n4474) );
  MUX2_X1 U32840 ( .A(DATAI_8_), .B(n4474), .S(n2697), .Z(n3265) );
  AND2_X1 U32850 ( .A1(n3847), .A2(n3265), .ZN(n2608) );
  INV_X1 U32860 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3294) );
  OR2_X1 U32870 ( .A1(n2566), .A2(n3294), .ZN(n2617) );
  INV_X1 U32880 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2609) );
  OR2_X1 U32890 ( .A1(n2772), .A2(n2609), .ZN(n2616) );
  INV_X1 U32900 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2610) );
  OAI21_X1 U32910 ( .B1(n2612), .B2(n2611), .A(n2610), .ZN(n2613) );
  NAND2_X1 U32920 ( .A1(n2613), .A2(n2626), .ZN(n3281) );
  OR2_X1 U32930 ( .A1(n2828), .A2(n3281), .ZN(n2615) );
  NAND2_X1 U32940 ( .A1(n2544), .A2(REG0_REG_9__SCAN_IN), .ZN(n2614) );
  NAND4_X1 U32950 ( .A1(n2617), .A2(n2616), .A3(n2615), .A4(n2614), .ZN(n3846)
         );
  INV_X1 U32960 ( .A(IR_REG_8__SCAN_IN), .ZN(n2618) );
  AND2_X1 U32970 ( .A1(n2619), .A2(n2618), .ZN(n2620) );
  NAND2_X1 U32980 ( .A1(n2621), .A2(n2620), .ZN(n2632) );
  NAND2_X1 U32990 ( .A1(n2632), .A2(IR_REG_31__SCAN_IN), .ZN(n2622) );
  XNOR2_X1 U33000 ( .A(n2622), .B(IR_REG_9__SCAN_IN), .ZN(n3909) );
  MUX2_X1 U33010 ( .A(DATAI_9_), .B(n3909), .S(n2697), .Z(n3285) );
  NOR2_X1 U33020 ( .A1(n3846), .A2(n3285), .ZN(n2624) );
  NAND2_X1 U33030 ( .A1(n3846), .A2(n3285), .ZN(n2623) );
  INV_X1 U33040 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2625) );
  OR2_X1 U33050 ( .A1(n2566), .A2(n2625), .ZN(n2631) );
  AND2_X1 U33060 ( .A1(n2626), .A2(n5045), .ZN(n2627) );
  OR2_X1 U33070 ( .A1(n2627), .A2(n2635), .ZN(n3330) );
  OR2_X1 U33080 ( .A1(n2828), .A2(n3330), .ZN(n2630) );
  INV_X1 U33090 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3306) );
  OR2_X1 U33100 ( .A1(n2772), .A2(n3306), .ZN(n2629) );
  NAND2_X1 U33110 ( .A1(n2544), .A2(REG0_REG_10__SCAN_IN), .ZN(n2628) );
  NAND4_X1 U33120 ( .A1(n2631), .A2(n2630), .A3(n2629), .A4(n2628), .ZN(n4593)
         );
  NAND2_X1 U33130 ( .A1(n2642), .A2(IR_REG_31__SCAN_IN), .ZN(n2633) );
  XNOR2_X1 U33140 ( .A(n2633), .B(IR_REG_10__SCAN_IN), .ZN(n4495) );
  MUX2_X1 U33150 ( .A(DATAI_10_), .B(n4495), .S(n2697), .Z(n3327) );
  INV_X1 U33160 ( .A(n4593), .ZN(n2801) );
  NAND2_X1 U33170 ( .A1(n2801), .A2(n3314), .ZN(n2634) );
  NOR2_X1 U33180 ( .A1(n2635), .A2(REG3_REG_11__SCAN_IN), .ZN(n2636) );
  OR2_X1 U33190 ( .A1(n2645), .A2(n2636), .ZN(n4601) );
  OR2_X1 U33200 ( .A1(n2828), .A2(n4601), .ZN(n2641) );
  INV_X1 U33210 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2637) );
  OR2_X1 U33220 ( .A1(n2772), .A2(n2637), .ZN(n2640) );
  NAND2_X1 U33230 ( .A1(n2538), .A2(REG1_REG_11__SCAN_IN), .ZN(n2639) );
  NAND2_X1 U33240 ( .A1(n2544), .A2(REG0_REG_11__SCAN_IN), .ZN(n2638) );
  NAND4_X1 U33250 ( .A1(n2641), .A2(n2640), .A3(n2639), .A4(n2638), .ZN(n3845)
         );
  INV_X1 U33260 ( .A(n3845), .ZN(n3373) );
  NAND2_X1 U33270 ( .A1(n2643), .A2(IR_REG_31__SCAN_IN), .ZN(n2652) );
  XNOR2_X1 U33280 ( .A(n2652), .B(IR_REG_11__SCAN_IN), .ZN(n3908) );
  MUX2_X1 U33290 ( .A(DATAI_11_), .B(n3908), .S(n2697), .Z(n4592) );
  NAND2_X1 U33300 ( .A1(n3373), .A2(n4592), .ZN(n3792) );
  NAND2_X1 U33310 ( .A1(n3845), .A2(n4604), .ZN(n3791) );
  NAND2_X1 U33320 ( .A1(n3792), .A2(n3791), .ZN(n4597) );
  INV_X1 U33330 ( .A(REG1_REG_12__SCAN_IN), .ZN(n2644) );
  OR2_X1 U33340 ( .A1(n2566), .A2(n2644), .ZN(n2650) );
  OR2_X1 U33350 ( .A1(n2645), .A2(REG3_REG_12__SCAN_IN), .ZN(n2646) );
  NAND2_X1 U33360 ( .A1(n2655), .A2(n2646), .ZN(n3589) );
  OR2_X1 U33370 ( .A1(n2828), .A2(n3589), .ZN(n2649) );
  INV_X1 U33380 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3361) );
  OR2_X1 U33390 ( .A1(n2772), .A2(n3361), .ZN(n2648) );
  NAND2_X1 U33400 ( .A1(n2544), .A2(REG0_REG_12__SCAN_IN), .ZN(n2647) );
  NAND4_X1 U33410 ( .A1(n2650), .A2(n2649), .A3(n2648), .A4(n2647), .ZN(n4331)
         );
  INV_X1 U33420 ( .A(n4331), .ZN(n4595) );
  INV_X1 U33430 ( .A(IR_REG_11__SCAN_IN), .ZN(n2651) );
  NAND2_X1 U33440 ( .A1(n2652), .A2(n2651), .ZN(n2653) );
  NAND2_X1 U33450 ( .A1(n2653), .A2(IR_REG_31__SCAN_IN), .ZN(n2654) );
  XNOR2_X1 U33460 ( .A(n2654), .B(IR_REG_12__SCAN_IN), .ZN(n4516) );
  MUX2_X1 U33470 ( .A(DATAI_12_), .B(n4516), .S(n2697), .Z(n3586) );
  INV_X1 U33480 ( .A(n3586), .ZN(n3401) );
  INV_X1 U33490 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4337) );
  OR2_X1 U33500 ( .A1(n2566), .A2(n4337), .ZN(n2660) );
  NAND2_X1 U33510 ( .A1(n2655), .A2(n5058), .ZN(n2656) );
  NAND2_X1 U33520 ( .A1(n2671), .A2(n2656), .ZN(n3642) );
  OR2_X1 U3353 ( .A1(n2828), .A2(n3642), .ZN(n2659) );
  NAND2_X1 U33540 ( .A1(n2544), .A2(REG0_REG_13__SCAN_IN), .ZN(n2658) );
  NAND2_X1 U3355 ( .A1(n3706), .A2(REG2_REG_13__SCAN_IN), .ZN(n2657) );
  NAND4_X1 U3356 ( .A1(n2660), .A2(n2659), .A3(n2658), .A4(n2657), .ZN(n4215)
         );
  INV_X1 U3357 ( .A(n4215), .ZN(n4321) );
  OR2_X1 U3358 ( .A1(n2661), .A2(n2705), .ZN(n2662) );
  XNOR2_X1 U3359 ( .A(n2662), .B(IR_REG_13__SCAN_IN), .ZN(n3907) );
  MUX2_X1 U3360 ( .A(DATAI_13_), .B(n3907), .S(n2697), .Z(n3639) );
  NAND2_X1 U3361 ( .A1(n4321), .A2(n4327), .ZN(n2663) );
  NAND2_X1 U3362 ( .A1(n3349), .A2(n2663), .ZN(n4187) );
  INV_X1 U3363 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4325) );
  OR2_X1 U3364 ( .A1(n2566), .A2(n4325), .ZN(n2668) );
  INV_X1 U3365 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2664) );
  XNOR2_X1 U3366 ( .A(n2671), .B(n2664), .ZN(n4217) );
  OR2_X1 U3367 ( .A1(n2828), .A2(n4217), .ZN(n2667) );
  NAND2_X1 U3368 ( .A1(n2544), .A2(REG0_REG_14__SCAN_IN), .ZN(n2666) );
  NAND2_X1 U3369 ( .A1(n3706), .A2(REG2_REG_14__SCAN_IN), .ZN(n2665) );
  NAND4_X1 U3370 ( .A1(n2668), .A2(n2667), .A3(n2666), .A4(n2665), .ZN(n4193)
         );
  INV_X1 U3371 ( .A(n4193), .ZN(n4329) );
  NAND2_X1 U3372 ( .A1(n2661), .A2(n2669), .ZN(n2679) );
  NAND2_X1 U3373 ( .A1(n2679), .A2(IR_REG_31__SCAN_IN), .ZN(n2670) );
  XNOR2_X1 U3374 ( .A(n2670), .B(IR_REG_14__SCAN_IN), .ZN(n3926) );
  MUX2_X1 U3375 ( .A(DATAI_14_), .B(n3926), .S(n2697), .Z(n4316) );
  NAND2_X1 U3376 ( .A1(n4329), .A2(n4316), .ZN(n4182) );
  INV_X1 U3377 ( .A(n4316), .ZN(n4222) );
  NAND2_X1 U3378 ( .A1(n4193), .A2(n4222), .ZN(n3688) );
  NAND2_X1 U3379 ( .A1(n4182), .A2(n3688), .ZN(n4208) );
  NAND2_X1 U3380 ( .A1(n4215), .A2(n3639), .ZN(n4186) );
  INV_X1 U3381 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4313) );
  OR2_X1 U3382 ( .A1(n2566), .A2(n4313), .ZN(n2678) );
  INV_X1 U3383 ( .A(n2671), .ZN(n2672) );
  AOI21_X1 U3384 ( .B1(n2672), .B2(REG3_REG_14__SCAN_IN), .A(
        REG3_REG_15__SCAN_IN), .ZN(n2673) );
  OR2_X1 U3385 ( .A1(n2673), .A2(n2685), .ZN(n4194) );
  OR2_X1 U3386 ( .A1(n2828), .A2(n4194), .ZN(n2677) );
  INV_X1 U3387 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2674) );
  OR2_X1 U3388 ( .A1(n2772), .A2(n2674), .ZN(n2676) );
  NAND2_X1 U3389 ( .A1(n2544), .A2(REG0_REG_15__SCAN_IN), .ZN(n2675) );
  NAND4_X1 U3390 ( .A1(n2678), .A2(n2677), .A3(n2676), .A4(n2675), .ZN(n4318)
         );
  NAND2_X1 U3391 ( .A1(n2680), .A2(IR_REG_31__SCAN_IN), .ZN(n2694) );
  MUX2_X1 U3392 ( .A(DATAI_15_), .B(n4648), .S(n2697), .Z(n4307) );
  NAND2_X1 U3393 ( .A1(n4318), .A2(n4307), .ZN(n2683) );
  NOR2_X1 U3394 ( .A1(n4193), .A2(n4316), .ZN(n4188) );
  INV_X1 U3395 ( .A(n4318), .ZN(n4418) );
  AOI22_X1 U3396 ( .A1(n4188), .A2(n2683), .B1(n4418), .B2(n4198), .ZN(n2684)
         );
  INV_X1 U3397 ( .A(n2685), .ZN(n2686) );
  INV_X1 U3398 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4414) );
  NAND2_X1 U3399 ( .A1(n2686), .A2(n4414), .ZN(n2687) );
  NAND2_X1 U3400 ( .A1(n2699), .A2(n2687), .ZN(n4431) );
  OR2_X1 U3401 ( .A1(n2828), .A2(n4431), .ZN(n2692) );
  INV_X1 U3402 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2688) );
  OR2_X1 U3403 ( .A1(n2566), .A2(n2688), .ZN(n2691) );
  NAND2_X1 U3404 ( .A1(n3706), .A2(REG2_REG_16__SCAN_IN), .ZN(n2690) );
  NAND2_X1 U3405 ( .A1(n2544), .A2(REG0_REG_16__SCAN_IN), .ZN(n2689) );
  NAND4_X1 U3406 ( .A1(n2692), .A2(n2691), .A3(n2690), .A4(n2689), .ZN(n4308)
         );
  INV_X1 U3407 ( .A(n4308), .ZN(n4296) );
  NAND2_X1 U3408 ( .A1(n2694), .A2(n2693), .ZN(n2695) );
  NAND2_X1 U3409 ( .A1(n2695), .A2(IR_REG_31__SCAN_IN), .ZN(n2696) );
  XNOR2_X1 U3410 ( .A(n2696), .B(IR_REG_16__SCAN_IN), .ZN(n3930) );
  MUX2_X1 U3411 ( .A(DATAI_16_), .B(n3930), .S(n2697), .Z(n4168) );
  NAND2_X1 U3412 ( .A1(n4296), .A2(n4168), .ZN(n3806) );
  INV_X1 U3413 ( .A(n4168), .ZN(n4415) );
  NAND2_X1 U3414 ( .A1(n4308), .A2(n4415), .ZN(n3803) );
  INV_X1 U3415 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2698) );
  NAND2_X1 U3416 ( .A1(n2699), .A2(n2698), .ZN(n2700) );
  NAND2_X1 U3417 ( .A1(n2710), .A2(n2700), .ZN(n4154) );
  OR2_X1 U3418 ( .A1(n2828), .A2(n4154), .ZN(n2704) );
  INV_X1 U3419 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4299) );
  OR2_X1 U3420 ( .A1(n2566), .A2(n4299), .ZN(n2703) );
  INV_X1 U3421 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4155) );
  OR2_X1 U3422 ( .A1(n2772), .A2(n4155), .ZN(n2702) );
  NAND2_X1 U3423 ( .A1(n2544), .A2(REG0_REG_17__SCAN_IN), .ZN(n2701) );
  NAND4_X1 U3424 ( .A1(n2704), .A2(n2703), .A3(n2702), .A4(n2701), .ZN(n4420)
         );
  INV_X1 U3425 ( .A(n4420), .ZN(n4140) );
  OR2_X1 U3426 ( .A1(n2706), .A2(n2705), .ZN(n2707) );
  XNOR2_X1 U3427 ( .A(n2707), .B(IR_REG_17__SCAN_IN), .ZN(n3933) );
  MUX2_X1 U3428 ( .A(DATAI_17_), .B(n3933), .S(n2697), .Z(n4292) );
  INV_X1 U3429 ( .A(n4292), .ZN(n2807) );
  NAND2_X1 U3430 ( .A1(n4140), .A2(n2807), .ZN(n2708) );
  NAND2_X1 U3431 ( .A1(n4420), .A2(n4292), .ZN(n2709) );
  INV_X1 U3432 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3935) );
  OR2_X1 U3433 ( .A1(n2566), .A2(n3935), .ZN(n2715) );
  NAND2_X1 U3434 ( .A1(n2710), .A2(n4578), .ZN(n2711) );
  NAND2_X1 U3435 ( .A1(n2721), .A2(n2711), .ZN(n4130) );
  OR2_X1 U3436 ( .A1(n2828), .A2(n4130), .ZN(n2714) );
  NAND2_X1 U3437 ( .A1(n2544), .A2(REG0_REG_18__SCAN_IN), .ZN(n2713) );
  NAND2_X1 U3438 ( .A1(n3706), .A2(REG2_REG_18__SCAN_IN), .ZN(n2712) );
  NAND4_X1 U3439 ( .A1(n2715), .A2(n2714), .A3(n2713), .A4(n2712), .ZN(n4293)
         );
  INV_X1 U3440 ( .A(n4293), .ZN(n2718) );
  NAND2_X1 U3441 ( .A1(n2716), .A2(IR_REG_31__SCAN_IN), .ZN(n2717) );
  XNOR2_X1 U3442 ( .A(n2717), .B(IR_REG_18__SCAN_IN), .ZN(n3906) );
  MUX2_X1 U3443 ( .A(DATAI_18_), .B(n3906), .S(n2697), .Z(n4138) );
  NAND2_X1 U3444 ( .A1(n2718), .A2(n4138), .ZN(n4109) );
  NAND2_X1 U3445 ( .A1(n4293), .A2(n4135), .ZN(n4110) );
  NAND2_X1 U3446 ( .A1(n2718), .A2(n4135), .ZN(n2719) );
  INV_X1 U3447 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4287) );
  OR2_X1 U3448 ( .A1(n2566), .A2(n4287), .ZN(n2726) );
  INV_X1 U3449 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2720) );
  NAND2_X1 U3450 ( .A1(n2721), .A2(n2720), .ZN(n2722) );
  NAND2_X1 U3451 ( .A1(n2728), .A2(n2722), .ZN(n4121) );
  OR2_X1 U3452 ( .A1(n2828), .A2(n4121), .ZN(n2725) );
  INV_X1 U3453 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4122) );
  OR2_X1 U3454 ( .A1(n2772), .A2(n4122), .ZN(n2724) );
  NAND2_X1 U3455 ( .A1(n2544), .A2(REG0_REG_19__SCAN_IN), .ZN(n2723) );
  NAND4_X1 U3456 ( .A1(n2726), .A2(n2725), .A3(n2724), .A4(n2723), .ZN(n4278)
         );
  MUX2_X1 U3457 ( .A(DATAI_19_), .B(n4143), .S(n2697), .Z(n3541) );
  NOR2_X1 U34580 ( .A1(n4278), .A2(n3541), .ZN(n4091) );
  NAND2_X1 U34590 ( .A1(n2544), .A2(REG0_REG_20__SCAN_IN), .ZN(n2733) );
  NAND2_X1 U3460 ( .A1(n2728), .A2(n4976), .ZN(n2729) );
  NAND2_X1 U3461 ( .A1(n2736), .A2(n2729), .ZN(n4097) );
  OR2_X1 U3462 ( .A1(n2828), .A2(n4097), .ZN(n2732) );
  NAND2_X1 U3463 ( .A1(n2538), .A2(REG1_REG_20__SCAN_IN), .ZN(n2731) );
  NAND2_X1 U3464 ( .A1(n3706), .A2(REG2_REG_20__SCAN_IN), .ZN(n2730) );
  NAND4_X1 U3465 ( .A1(n2733), .A2(n2732), .A3(n2731), .A4(n2730), .ZN(n4079)
         );
  NAND2_X1 U3466 ( .A1(n4079), .A2(n3629), .ZN(n3730) );
  NAND2_X1 U34670 ( .A1(n4278), .A2(n3541), .ZN(n4092) );
  INV_X1 U3468 ( .A(n4079), .ZN(n4269) );
  INV_X1 U34690 ( .A(n3629), .ZN(n4275) );
  NAND2_X1 U3470 ( .A1(n4269), .A2(n4275), .ZN(n3731) );
  NAND2_X1 U34710 ( .A1(n2734), .A2(n3731), .ZN(n4072) );
  NAND2_X1 U3472 ( .A1(n2544), .A2(REG0_REG_21__SCAN_IN), .ZN(n2742) );
  INV_X1 U34730 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2735) );
  NAND2_X1 U3474 ( .A1(n2736), .A2(n2735), .ZN(n2737) );
  NAND2_X1 U34750 ( .A1(n2738), .A2(n2737), .ZN(n4080) );
  OR2_X1 U3476 ( .A1(n2828), .A2(n4080), .ZN(n2741) );
  NAND2_X1 U34770 ( .A1(n2538), .A2(REG1_REG_21__SCAN_IN), .ZN(n2740) );
  NAND2_X1 U3478 ( .A1(n3706), .A2(REG2_REG_21__SCAN_IN), .ZN(n2739) );
  NAND4_X1 U34790 ( .A1(n2742), .A2(n2741), .A3(n2740), .A4(n2739), .ZN(n4096)
         );
  NAND2_X1 U3480 ( .A1(n4096), .A2(n4266), .ZN(n2745) );
  NOR2_X1 U34810 ( .A1(n4096), .A2(n4266), .ZN(n2744) );
  INV_X1 U3482 ( .A(n4267), .ZN(n2746) );
  NAND2_X1 U34830 ( .A1(n2746), .A2(n3474), .ZN(n4039) );
  NAND2_X1 U3484 ( .A1(n4267), .A2(n4064), .ZN(n2817) );
  NAND2_X1 U34850 ( .A1(n4039), .A2(n2817), .ZN(n4060) );
  NAND2_X1 U3486 ( .A1(n2544), .A2(REG0_REG_23__SCAN_IN), .ZN(n2752) );
  INV_X1 U34870 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4826) );
  NAND2_X1 U3488 ( .A1(n2747), .A2(n4826), .ZN(n2748) );
  NAND2_X1 U34890 ( .A1(n2754), .A2(n2748), .ZN(n4048) );
  OR2_X1 U3490 ( .A1(n2828), .A2(n4048), .ZN(n2751) );
  NAND2_X1 U34910 ( .A1(n2538), .A2(REG1_REG_23__SCAN_IN), .ZN(n2750) );
  NAND2_X1 U3492 ( .A1(n3706), .A2(REG2_REG_23__SCAN_IN), .ZN(n2749) );
  NAND4_X1 U34930 ( .A1(n2752), .A2(n2751), .A3(n2750), .A4(n2749), .ZN(n4055)
         );
  NOR2_X1 U3494 ( .A1(n4055), .A2(n3534), .ZN(n3729) );
  NAND2_X1 U34950 ( .A1(n2754), .A2(n4839), .ZN(n2755) );
  NAND2_X1 U3496 ( .A1(n2760), .A2(n2755), .ZN(n4032) );
  INV_X1 U34970 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4033) );
  OAI22_X1 U3498 ( .A1(n4032), .A2(n2828), .B1(n2772), .B2(n4033), .ZN(n2758)
         );
  INV_X1 U34990 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4255) );
  NAND2_X1 U3500 ( .A1(n2544), .A2(REG0_REG_24__SCAN_IN), .ZN(n2756) );
  OAI21_X1 U35010 ( .B1(n2566), .B2(n4255), .A(n2756), .ZN(n2757) );
  INV_X1 U3502 ( .A(n4007), .ZN(n4042) );
  NAND2_X1 U35030 ( .A1(n3709), .A2(DATAI_24_), .ZN(n4023) );
  NOR2_X1 U3504 ( .A1(n4042), .A2(n4023), .ZN(n2759) );
  OAI22_X1 U35050 ( .A1(n4018), .A2(n2759), .B1(n4029), .B2(n4007), .ZN(n4000)
         );
  INV_X1 U35060 ( .A(REG2_REG_26__SCAN_IN), .ZN(n3994) );
  INV_X1 U35070 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3597) );
  INV_X1 U35080 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3670) );
  OAI21_X1 U35090 ( .B1(n2760), .B2(n3597), .A(n3670), .ZN(n2763) );
  INV_X1 U35100 ( .A(n2760), .ZN(n2762) );
  AND2_X1 U35110 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2761) );
  NAND2_X1 U35120 ( .A1(n2762), .A2(n2761), .ZN(n2767) );
  NAND2_X1 U35130 ( .A1(n2763), .A2(n2767), .ZN(n3995) );
  OR2_X1 U35140 ( .A1(n3995), .A2(n2828), .ZN(n2765) );
  AOI22_X1 U35150 ( .A1(n2538), .A2(REG1_REG_26__SCAN_IN), .B1(n2544), .B2(
        REG0_REG_26__SCAN_IN), .ZN(n2764) );
  OAI211_X1 U35160 ( .C1(n2772), .C2(n3994), .A(n2765), .B(n2764), .ZN(n4237)
         );
  INV_X1 U35170 ( .A(DATAI_26_), .ZN(n4879) );
  NAND2_X1 U35180 ( .A1(n4237), .A2(n3500), .ZN(n2766) );
  INV_X1 U35190 ( .A(n4237), .ZN(n4005) );
  INV_X1 U35200 ( .A(REG2_REG_27__SCAN_IN), .ZN(n2771) );
  NAND2_X1 U35210 ( .A1(n2767), .A2(n3515), .ZN(n2768) );
  NAND2_X1 U35220 ( .A1(n2774), .A2(n2768), .ZN(n3514) );
  OR2_X1 U35230 ( .A1(n3514), .A2(n2828), .ZN(n2770) );
  AOI22_X1 U35240 ( .A1(n2538), .A2(REG1_REG_27__SCAN_IN), .B1(n2544), .B2(
        REG0_REG_27__SCAN_IN), .ZN(n2769) );
  OAI211_X1 U35250 ( .C1(n2772), .C2(n2771), .A(n2770), .B(n2769), .ZN(n3844)
         );
  INV_X1 U35260 ( .A(n3844), .ZN(n3986) );
  INV_X1 U35270 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3560) );
  NAND2_X1 U35280 ( .A1(n2774), .A2(n3560), .ZN(n2775) );
  NAND2_X1 U35290 ( .A1(n3959), .A2(n2537), .ZN(n2780) );
  NAND2_X1 U35300 ( .A1(n2544), .A2(REG0_REG_28__SCAN_IN), .ZN(n2777) );
  NAND2_X1 U35310 ( .A1(n3706), .A2(REG2_REG_28__SCAN_IN), .ZN(n2776) );
  OAI211_X1 U35320 ( .C1(n2566), .C2(n2864), .A(n2777), .B(n2776), .ZN(n2778)
         );
  INV_X1 U35330 ( .A(n2778), .ZN(n2779) );
  NAND2_X1 U35340 ( .A1(n3709), .A2(DATAI_28_), .ZN(n3559) );
  NAND2_X1 U35350 ( .A1(n3972), .A2(n3559), .ZN(n3704) );
  INV_X1 U35360 ( .A(n3559), .ZN(n2873) );
  NAND2_X1 U35370 ( .A1(n4240), .A2(n2873), .ZN(n3702) );
  NAND2_X1 U35380 ( .A1(n3704), .A2(n3702), .ZN(n3718) );
  INV_X1 U35390 ( .A(n3718), .ZN(n2781) );
  XNOR2_X1 U35400 ( .A(n2874), .B(n2781), .ZN(n3958) );
  NAND2_X1 U35410 ( .A1(n2785), .A2(n2784), .ZN(n2786) );
  XNOR2_X1 U35420 ( .A(n3008), .B(n2829), .ZN(n2791) );
  AND2_X1 U35430 ( .A1(n3831), .A2(n4143), .ZN(n2997) );
  NAND2_X1 U35440 ( .A1(n2506), .A2(IR_REG_31__SCAN_IN), .ZN(n2793) );
  XNOR2_X1 U35450 ( .A(n2793), .B(n2792), .ZN(n4413) );
  NAND2_X1 U35460 ( .A1(n4406), .A2(n3757), .ZN(n2941) );
  INV_X1 U35470 ( .A(n4629), .ZN(n2933) );
  NAND2_X1 U35480 ( .A1(n2990), .A2(n2933), .ZN(n3754) );
  INV_X1 U35490 ( .A(n2794), .ZN(n2795) );
  NAND2_X1 U35500 ( .A1(n3066), .A2(n3759), .ZN(n2797) );
  XNOR2_X1 U35510 ( .A(n3852), .B(n3763), .ZN(n3065) );
  NAND2_X1 U35520 ( .A1(n3764), .A2(n3763), .ZN(n3765) );
  AND2_X1 U35530 ( .A1(n3850), .A2(n3152), .ZN(n3092) );
  NAND2_X1 U35540 ( .A1(n3181), .A2(n3157), .ZN(n3778) );
  NAND2_X1 U35550 ( .A1(n3849), .A2(n3170), .ZN(n3779) );
  NAND2_X1 U35560 ( .A1(n3118), .A2(n3779), .ZN(n2798) );
  INV_X1 U35570 ( .A(n3849), .ZN(n3200) );
  NAND2_X1 U35580 ( .A1(n3200), .A2(n3179), .ZN(n3771) );
  NAND2_X1 U35590 ( .A1(n2798), .A2(n3771), .ZN(n3196) );
  INV_X1 U35600 ( .A(n3772), .ZN(n2799) );
  INV_X1 U35610 ( .A(n3847), .ZN(n3288) );
  NAND2_X1 U35620 ( .A1(n3288), .A2(n3265), .ZN(n3775) );
  INV_X1 U35630 ( .A(n3265), .ZN(n3258) );
  NAND2_X1 U35640 ( .A1(n3847), .A2(n3258), .ZN(n3780) );
  INV_X1 U35650 ( .A(n3285), .ZN(n3227) );
  AND2_X1 U35660 ( .A1(n3846), .A2(n3227), .ZN(n3220) );
  INV_X1 U35670 ( .A(n3846), .ZN(n3300) );
  NAND2_X1 U35680 ( .A1(n3300), .A2(n3285), .ZN(n3776) );
  NAND2_X1 U35690 ( .A1(n4593), .A2(n3314), .ZN(n3790) );
  NAND2_X1 U35700 ( .A1(n2801), .A2(n3327), .ZN(n3786) );
  NOR2_X1 U35710 ( .A1(n4331), .A2(n3401), .ZN(n3794) );
  NAND2_X1 U35720 ( .A1(n4215), .A2(n4327), .ZN(n3347) );
  NAND2_X1 U35730 ( .A1(n4331), .A2(n3401), .ZN(n3345) );
  AND2_X1 U35740 ( .A1(n3347), .A2(n3345), .ZN(n3793) );
  NAND2_X1 U35750 ( .A1(n4321), .A2(n3639), .ZN(n3797) );
  NAND2_X1 U35760 ( .A1(n4418), .A2(n4307), .ZN(n3796) );
  NAND2_X1 U35770 ( .A1(n4318), .A2(n4198), .ZN(n3689) );
  NAND2_X1 U35780 ( .A1(n3796), .A2(n3689), .ZN(n4190) );
  INV_X1 U35790 ( .A(n4182), .ZN(n2803) );
  NOR2_X1 U35800 ( .A1(n4190), .A2(n2803), .ZN(n2804) );
  NAND2_X1 U35810 ( .A1(n4206), .A2(n2804), .ZN(n2805) );
  NAND2_X1 U3582 ( .A1(n2805), .A2(n3689), .ZN(n4163) );
  NAND2_X1 U3583 ( .A1(n4278), .A2(n4118), .ZN(n2806) );
  AND2_X1 U3584 ( .A1(n4110), .A2(n2806), .ZN(n2808) );
  NAND2_X1 U3585 ( .A1(n4420), .A2(n2807), .ZN(n4106) );
  NAND2_X1 U3586 ( .A1(n2808), .A2(n4106), .ZN(n3805) );
  NAND2_X1 U3587 ( .A1(n4140), .A2(n4292), .ZN(n4107) );
  NAND2_X1 U3588 ( .A1(n4109), .A2(n4107), .ZN(n2809) );
  NAND2_X1 U3589 ( .A1(n2809), .A2(n2808), .ZN(n2812) );
  INV_X1 U3590 ( .A(n4278), .ZN(n2810) );
  NAND2_X1 U3591 ( .A1(n2810), .A2(n3541), .ZN(n2811) );
  NAND2_X1 U3592 ( .A1(n2812), .A2(n2811), .ZN(n4089) );
  NOR2_X1 U3593 ( .A1(n4079), .A2(n4275), .ZN(n2813) );
  OR2_X1 U3594 ( .A1(n4089), .A2(n2813), .ZN(n3810) );
  INV_X1 U3595 ( .A(n3810), .ZN(n2814) );
  NAND2_X1 U3596 ( .A1(n4079), .A2(n4275), .ZN(n3809) );
  INV_X1 U3597 ( .A(n4096), .ZN(n4276) );
  NAND2_X1 U3598 ( .A1(n4276), .A2(n4266), .ZN(n4038) );
  AND2_X1 U3599 ( .A1(n4039), .A2(n4038), .ZN(n3814) );
  NAND2_X1 U3600 ( .A1(n4074), .A2(n3814), .ZN(n2821) );
  NAND2_X1 U3601 ( .A1(n4055), .A2(n4047), .ZN(n2816) );
  NAND2_X1 U3602 ( .A1(n2817), .A2(n2816), .ZN(n3812) );
  INV_X1 U3603 ( .A(n3812), .ZN(n2820) );
  INV_X1 U3604 ( .A(n4266), .ZN(n4084) );
  NAND2_X1 U3605 ( .A1(n4096), .A2(n4084), .ZN(n3808) );
  INV_X1 U3606 ( .A(n3808), .ZN(n2818) );
  NAND2_X1 U3607 ( .A1(n2818), .A2(n4039), .ZN(n2819) );
  AND2_X1 U3608 ( .A1(n2820), .A2(n2819), .ZN(n3697) );
  NAND2_X1 U3609 ( .A1(n2821), .A2(n3697), .ZN(n4020) );
  NAND2_X1 U3610 ( .A1(n4042), .A2(n4029), .ZN(n3736) );
  INV_X1 U3611 ( .A(n4055), .ZN(n4024) );
  NAND2_X1 U3612 ( .A1(n4024), .A2(n3534), .ZN(n4019) );
  AND2_X1 U3613 ( .A1(n3736), .A2(n4019), .ZN(n3695) );
  NAND2_X1 U3614 ( .A1(n4020), .A2(n3695), .ZN(n4002) );
  NAND2_X1 U3615 ( .A1(n4026), .A2(n4011), .ZN(n3732) );
  NAND2_X1 U3616 ( .A1(n4007), .A2(n4023), .ZN(n4001) );
  AND2_X1 U3617 ( .A1(n3732), .A2(n4001), .ZN(n3815) );
  NAND2_X1 U3618 ( .A1(n4002), .A2(n3815), .ZN(n3983) );
  OR2_X1 U3619 ( .A1(n4237), .A2(n3992), .ZN(n3717) );
  OR2_X1 U3620 ( .A1(n4026), .A2(n4011), .ZN(n3982) );
  AND2_X1 U3621 ( .A1(n3717), .A2(n3982), .ZN(n3818) );
  NAND2_X1 U3622 ( .A1(n4237), .A2(n3992), .ZN(n3822) );
  NAND2_X1 U3623 ( .A1(n3986), .A2(n4236), .ZN(n3701) );
  NAND2_X1 U3624 ( .A1(n3844), .A2(n3976), .ZN(n3821) );
  INV_X1 U3625 ( .A(n3701), .ZN(n2822) );
  XNOR2_X1 U3626 ( .A(n2876), .B(n3718), .ZN(n2825) );
  OR2_X1 U3627 ( .A1(n2829), .A2(n3940), .ZN(n2824) );
  OR2_X1 U3628 ( .A1(n3751), .A2(n3831), .ZN(n2823) );
  NAND2_X1 U3629 ( .A1(n2825), .A2(n4625), .ZN(n2831) );
  AOI22_X1 U3630 ( .A1(n2544), .A2(REG0_REG_29__SCAN_IN), .B1(n2538), .B2(
        REG1_REG_29__SCAN_IN), .ZN(n2827) );
  NAND2_X1 U3631 ( .A1(n3706), .A2(REG2_REG_29__SCAN_IN), .ZN(n2826) );
  OAI211_X1 U3632 ( .C1(n3951), .C2(n2828), .A(n2827), .B(n2826), .ZN(n3843)
         );
  INV_X1 U3633 ( .A(n2941), .ZN(n2904) );
  NAND2_X1 U3634 ( .A1(n2829), .A2(n3751), .ZN(n2996) );
  AOI22_X1 U3635 ( .A1(n3843), .A2(n4317), .B1(n4611), .B2(n2873), .ZN(n2830)
         );
  OAI211_X1 U3636 ( .C1(n3986), .C2(n4320), .A(n2831), .B(n2830), .ZN(n3963)
         );
  AOI21_X1 U3637 ( .B1(n3958), .B2(n4678), .A(n3963), .ZN(n2869) );
  NAND2_X1 U3638 ( .A1(n2244), .A2(IR_REG_31__SCAN_IN), .ZN(n2833) );
  MUX2_X1 U3639 ( .A(n2833), .B(IR_REG_31__SCAN_IN), .S(n2832), .Z(n2834) );
  NAND2_X1 U3640 ( .A1(n2911), .A2(B_REG_SCAN_IN), .ZN(n2837) );
  NAND2_X1 U3641 ( .A1(n2846), .A2(n2845), .ZN(n2835) );
  MUX2_X1 U3642 ( .A(n2837), .B(B_REG_SCAN_IN), .S(n4405), .Z(n2842) );
  NAND2_X1 U3643 ( .A1(n2838), .A2(IR_REG_31__SCAN_IN), .ZN(n2839) );
  INV_X1 U3644 ( .A(n3003), .ZN(n2844) );
  AND2_X1 U3645 ( .A1(n2912), .A2(n2911), .ZN(n2937) );
  INV_X1 U3646 ( .A(n2937), .ZN(n2843) );
  NAND2_X1 U3647 ( .A1(n2844), .A2(n2843), .ZN(n2861) );
  AND2_X1 U3648 ( .A1(n3831), .A2(n3940), .ZN(n2940) );
  OR2_X1 U3649 ( .A1(n2941), .A2(n2940), .ZN(n3000) );
  INV_X1 U3650 ( .A(n2953), .ZN(n2847) );
  NAND3_X1 U3651 ( .A1(n3001), .A2(n3000), .A3(n2847), .ZN(n2859) );
  NOR4_X1 U3652 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2851) );
  NOR4_X1 U3653 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2850) );
  NOR4_X1 U3654 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n2849) );
  NOR4_X1 U3655 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2848) );
  NAND4_X1 U3656 ( .A1(n2851), .A2(n2850), .A3(n2849), .A4(n2848), .ZN(n2857)
         );
  NOR2_X1 U3657 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_14__SCAN_IN), .ZN(n2855)
         );
  NOR4_X1 U3658 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2854) );
  NOR4_X1 U3659 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_29__SCAN_IN), .ZN(n2853) );
  NOR4_X1 U3660 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2852) );
  NAND4_X1 U3661 ( .A1(n2855), .A2(n2854), .A3(n2853), .A4(n2852), .ZN(n2856)
         );
  NOR2_X1 U3662 ( .A1(n2857), .A2(n2856), .ZN(n2858) );
  NOR2_X1 U3663 ( .A1(n2859), .A2(n2938), .ZN(n2860) );
  NAND2_X1 U3664 ( .A1(n2912), .A2(n2908), .ZN(n2862) );
  INV_X1 U3665 ( .A(n3004), .ZN(n2863) );
  MUX2_X1 U3666 ( .A(n2864), .B(n2869), .S(n4717), .Z(n2867) );
  NAND2_X1 U3667 ( .A1(n4630), .A2(n4629), .ZN(n4628) );
  NAND2_X1 U3668 ( .A1(n3192), .A2(n3210), .ZN(n3193) );
  NOR2_X1 U3669 ( .A1(n3225), .A2(n3285), .ZN(n3305) );
  NAND2_X1 U3670 ( .A1(n4211), .A2(n4198), .ZN(n4192) );
  INV_X1 U3671 ( .A(n2888), .ZN(n2865) );
  OAI21_X1 U3672 ( .B1(n3970), .B2(n3559), .A(n2865), .ZN(n3961) );
  INV_X1 U3673 ( .A(n3831), .ZN(n4407) );
  NAND2_X1 U3674 ( .A1(n2867), .A2(n2866), .ZN(U3546) );
  INV_X1 U3675 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2870) );
  MUX2_X1 U3676 ( .A(n2870), .B(n2869), .S(n4701), .Z(n2872) );
  NAND2_X1 U3677 ( .A1(n2872), .A2(n2871), .ZN(U3514) );
  INV_X1 U3678 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2887) );
  AOI22_X1 U3679 ( .A1(n2874), .A2(n3718), .B1(n2873), .B2(n3972), .ZN(n2875)
         );
  NAND2_X1 U3680 ( .A1(n3709), .A2(DATAI_29_), .ZN(n3956) );
  XNOR2_X1 U3681 ( .A(n3843), .B(n3956), .ZN(n3749) );
  XNOR2_X1 U3682 ( .A(n2875), .B(n3749), .ZN(n3957) );
  XNOR2_X1 U3683 ( .A(n2877), .B(n3749), .ZN(n2885) );
  NAND2_X1 U3684 ( .A1(n2538), .A2(REG1_REG_30__SCAN_IN), .ZN(n2881) );
  NAND2_X1 U3685 ( .A1(n3706), .A2(REG2_REG_30__SCAN_IN), .ZN(n2880) );
  INV_X1 U3686 ( .A(REG0_REG_30__SCAN_IN), .ZN(n2878) );
  OR2_X1 U3687 ( .A1(n2553), .A2(n2878), .ZN(n2879) );
  AND3_X1 U3688 ( .A1(n2881), .A2(n2880), .A3(n2879), .ZN(n3712) );
  INV_X1 U3689 ( .A(B_REG_SCAN_IN), .ZN(n2884) );
  OR2_X1 U3690 ( .A1(n2883), .A2(n2882), .ZN(n2958) );
  OAI21_X1 U3691 ( .B1(n2884), .B2(n2958), .A(n4317), .ZN(n3946) );
  OAI22_X1 U3692 ( .A1(n2885), .A2(n4333), .B1(n3712), .B2(n3946), .ZN(n3954)
         );
  OAI22_X1 U3693 ( .A1(n4240), .A2(n4320), .B1(n4328), .B2(n3956), .ZN(n2886)
         );
  MUX2_X1 U3694 ( .A(n2887), .B(n2891), .S(n4717), .Z(n2890) );
  NAND2_X1 U3695 ( .A1(n2888), .A2(n3956), .ZN(n4231) );
  OAI21_X1 U3696 ( .B1(n2888), .B2(n3956), .A(n4231), .ZN(n3952) );
  NAND2_X1 U3697 ( .A1(n2890), .A2(n2889), .ZN(U3547) );
  INV_X1 U3698 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2892) );
  MUX2_X1 U3699 ( .A(n2892), .B(n2891), .S(n4701), .Z(n2894) );
  NAND2_X1 U3700 ( .A1(n2894), .A2(n2893), .ZN(U3515) );
  INV_X1 U3701 ( .A(DATAI_19_), .ZN(n4852) );
  MUX2_X1 U3702 ( .A(n3940), .B(n4852), .S(U3149), .Z(n2896) );
  INV_X1 U3703 ( .A(n2896), .ZN(U3333) );
  NAND2_X1 U3704 ( .A1(n3757), .A2(STATE_REG_SCAN_IN), .ZN(n2897) );
  OAI21_X1 U3705 ( .B1(STATE_REG_SCAN_IN), .B2(n2743), .A(n2897), .ZN(U3331)
         );
  NAND2_X1 U3706 ( .A1(n2323), .A2(STATE_REG_SCAN_IN), .ZN(n2898) );
  OAI21_X1 U3707 ( .B1(STATE_REG_SCAN_IN), .B2(n2499), .A(n2898), .ZN(U3327)
         );
  INV_X1 U3708 ( .A(DATAI_29_), .ZN(n4979) );
  NAND2_X1 U3709 ( .A1(n2899), .A2(STATE_REG_SCAN_IN), .ZN(n2900) );
  OAI21_X1 U3710 ( .B1(STATE_REG_SCAN_IN), .B2(n4979), .A(n2900), .ZN(U3323)
         );
  INV_X1 U3711 ( .A(n2958), .ZN(n4437) );
  NAND2_X1 U3712 ( .A1(n4437), .A2(STATE_REG_SCAN_IN), .ZN(n2901) );
  OAI21_X1 U3713 ( .B1(STATE_REG_SCAN_IN), .B2(n2773), .A(n2901), .ZN(U3325)
         );
  NAND2_X1 U3714 ( .A1(n2508), .A2(STATE_REG_SCAN_IN), .ZN(n2902) );
  OAI21_X1 U3715 ( .B1(STATE_REG_SCAN_IN), .B2(n4746), .A(n2902), .ZN(U3322)
         );
  INV_X1 U3716 ( .A(n3001), .ZN(n2903) );
  OR2_X1 U3717 ( .A1(n3033), .A2(U3149), .ZN(n3839) );
  NAND2_X1 U3718 ( .A1(n2903), .A2(n3839), .ZN(n2918) );
  AND2_X1 U3719 ( .A1(n2904), .A2(n3033), .ZN(n2905) );
  NOR2_X1 U3720 ( .A1(n2697), .A2(n2905), .ZN(n2917) );
  INV_X1 U3721 ( .A(n2917), .ZN(n2906) );
  NOR2_X1 U3722 ( .A1(n4583), .A2(U4043), .ZN(U3148) );
  AND2_X2 U3723 ( .A1(n2907), .A2(n3001), .ZN(n4642) );
  NAND3_X1 U3724 ( .A1(n2912), .A2(n4643), .A3(n2908), .ZN(n2909) );
  OAI21_X1 U3725 ( .B1(n4642), .B2(D_REG_0__SCAN_IN), .A(n2909), .ZN(n2910) );
  INV_X1 U3726 ( .A(n2910), .ZN(U3458) );
  NAND3_X1 U3727 ( .A1(n2912), .A2(n4643), .A3(n2911), .ZN(n2913) );
  OAI21_X1 U3728 ( .B1(n4642), .B2(D_REG_1__SCAN_IN), .A(n2913), .ZN(n2914) );
  INV_X1 U3729 ( .A(n2914), .ZN(U3459) );
  INV_X1 U3730 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3869) );
  INV_X1 U3731 ( .A(n4410), .ZN(n3867) );
  INV_X1 U3732 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2915) );
  INV_X1 U3733 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3011) );
  MUX2_X1 U3734 ( .A(REG2_REG_2__SCAN_IN), .B(n3869), .S(n4410), .Z(n2916) );
  XNOR2_X1 U3735 ( .A(n2962), .B(REG2_REG_3__SCAN_IN), .ZN(n2927) );
  NOR2_X1 U3736 ( .A1(n4413), .A2(n2958), .ZN(n3835) );
  INV_X1 U3737 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3106) );
  NOR2_X1 U3738 ( .A1(STATE_REG_SCAN_IN), .A2(n3106), .ZN(n3039) );
  INV_X1 U3739 ( .A(n4409), .ZN(n2923) );
  NOR2_X1 U3740 ( .A1(n4590), .A2(n2923), .ZN(n2919) );
  AOI211_X1 U3741 ( .C1(n4583), .C2(ADDR_REG_3__SCAN_IN), .A(n3039), .B(n2919), 
        .ZN(n2926) );
  XNOR2_X1 U3742 ( .A(n3859), .B(REG1_REG_1__SCAN_IN), .ZN(n3858) );
  AND2_X1 U3743 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3857)
         );
  NAND2_X1 U3744 ( .A1(n3858), .A2(n3857), .ZN(n3856) );
  NAND2_X1 U3745 ( .A1(n4411), .A2(REG1_REG_1__SCAN_IN), .ZN(n2920) );
  NAND2_X1 U3746 ( .A1(n3856), .A2(n2920), .ZN(n3875) );
  INV_X1 U3747 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2921) );
  MUX2_X1 U3748 ( .A(REG1_REG_2__SCAN_IN), .B(n2921), .S(n4410), .Z(n3876) );
  NAND2_X1 U3749 ( .A1(n3875), .A2(n3876), .ZN(n3874) );
  NAND2_X1 U3750 ( .A1(n4410), .A2(REG1_REG_2__SCAN_IN), .ZN(n2922) );
  NAND2_X1 U3751 ( .A1(n3874), .A2(n2922), .ZN(n2963) );
  XNOR2_X1 U3752 ( .A(n2963), .B(n2923), .ZN(n2924) );
  NAND2_X1 U3753 ( .A1(n2924), .A2(REG1_REG_3__SCAN_IN), .ZN(n2965) );
  OAI211_X1 U3754 ( .C1(REG1_REG_3__SCAN_IN), .C2(n2924), .A(n4585), .B(n2965), 
        .ZN(n2925) );
  OAI211_X1 U3755 ( .C1(n2927), .C2(n4579), .A(n2926), .B(n2925), .ZN(U3243)
         );
  NAND2_X1 U3756 ( .A1(n3513), .A2(n4614), .ZN(n2931) );
  INV_X1 U3757 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2934) );
  OAI21_X1 U3759 ( .B1(n3034), .B2(n2934), .A(n2981), .ZN(n2935) );
  NAND2_X1 U3760 ( .A1(n2936), .A2(n2935), .ZN(n2984) );
  OAI21_X1 U3761 ( .B1(n2936), .B2(n2935), .A(n2984), .ZN(n2959) );
  NOR2_X1 U3762 ( .A1(n2938), .A2(n2937), .ZN(n3006) );
  NOR2_X1 U3763 ( .A1(n3004), .A2(n3003), .ZN(n2939) );
  NAND2_X1 U3764 ( .A1(n3006), .A2(n2939), .ZN(n2989) );
  OR2_X1 U3765 ( .A1(n2996), .A2(n2940), .ZN(n2942) );
  NAND2_X1 U3766 ( .A1(n2942), .A2(n2941), .ZN(n2945) );
  INV_X1 U3767 ( .A(n2945), .ZN(n2943) );
  NAND2_X1 U3768 ( .A1(n3001), .A2(n2943), .ZN(n2944) );
  NAND2_X1 U3769 ( .A1(n2945), .A2(n4328), .ZN(n2946) );
  NAND2_X1 U3770 ( .A1(n2989), .A2(n2946), .ZN(n2947) );
  NAND2_X1 U3771 ( .A1(n2947), .A2(n3000), .ZN(n3036) );
  INV_X1 U3772 ( .A(n3036), .ZN(n2949) );
  NAND2_X1 U3773 ( .A1(n4643), .A2(n2975), .ZN(n2948) );
  NAND2_X1 U3774 ( .A1(n2989), .A2(n3836), .ZN(n3037) );
  NAND3_X1 U3775 ( .A1(n2949), .A2(n3001), .A3(n3037), .ZN(n3024) );
  NAND2_X1 U3776 ( .A1(n3836), .A2(n4413), .ZN(n2951) );
  OR2_X1 U3777 ( .A1(n2989), .A2(n2951), .ZN(n3672) );
  NAND2_X1 U3778 ( .A1(n3001), .A2(n4611), .ZN(n2952) );
  OR2_X1 U3779 ( .A1(n2989), .A2(n2952), .ZN(n2954) );
  OAI22_X1 U3780 ( .A1(n2950), .A2(n3672), .B1(n4416), .B2(n4629), .ZN(n2955)
         );
  AOI21_X1 U3781 ( .B1(REG3_REG_0__SCAN_IN), .B2(n3024), .A(n2955), .ZN(n2956)
         );
  OAI21_X1 U3782 ( .B1(n2959), .B2(n3678), .A(n2956), .ZN(U3229) );
  INV_X1 U3783 ( .A(n4413), .ZN(n2987) );
  NAND2_X1 U3784 ( .A1(n4437), .A2(n3011), .ZN(n2957) );
  NAND2_X1 U3785 ( .A1(n2987), .A2(n2957), .ZN(n4438) );
  INV_X1 U3786 ( .A(n4438), .ZN(n4436) );
  NAND3_X1 U3787 ( .A1(n2959), .A2(n2987), .A3(n2958), .ZN(n2961) );
  AND2_X1 U3788 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3861)
         );
  AOI21_X1 U3789 ( .B1(n3835), .B2(n3861), .A(n3854), .ZN(n2960) );
  OAI211_X1 U3790 ( .C1(n4436), .C2(IR_REG_0__SCAN_IN), .A(n2961), .B(n2960), 
        .ZN(n3880) );
  XNOR2_X1 U3791 ( .A(n3886), .B(n4408), .ZN(n3883) );
  XOR2_X1 U3792 ( .A(REG2_REG_4__SCAN_IN), .B(n3883), .Z(n2972) );
  INV_X1 U3793 ( .A(n4408), .ZN(n3885) );
  NAND2_X1 U3794 ( .A1(n2963), .A2(n4409), .ZN(n2964) );
  NAND2_X1 U3795 ( .A1(n2965), .A2(n2964), .ZN(n3911) );
  XNOR2_X1 U3796 ( .A(n3911), .B(n3885), .ZN(n2966) );
  INV_X1 U3797 ( .A(n2966), .ZN(n2967) );
  INV_X1 U3798 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4709) );
  NAND2_X1 U3799 ( .A1(n2967), .A2(n4709), .ZN(n2968) );
  NAND3_X1 U3800 ( .A1(n4585), .A2(n3910), .A3(n2968), .ZN(n2970) );
  INV_X1 U3801 ( .A(REG3_REG_4__SCAN_IN), .ZN(n4988) );
  NOR2_X1 U3802 ( .A1(STATE_REG_SCAN_IN), .A2(n4988), .ZN(n3384) );
  AOI21_X1 U3803 ( .B1(n4583), .B2(ADDR_REG_4__SCAN_IN), .A(n3384), .ZN(n2969)
         );
  OAI211_X1 U3804 ( .C1(n4590), .C2(n3885), .A(n2970), .B(n2969), .ZN(n2971)
         );
  AOI21_X1 U3805 ( .B1(n4528), .B2(n2972), .A(n2971), .ZN(n2973) );
  NAND2_X1 U3806 ( .A1(n3880), .A2(n2973), .ZN(U3244) );
  INV_X1 U3807 ( .A(n3024), .ZN(n2995) );
  INV_X1 U3808 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2994) );
  NOR2_X1 U3809 ( .A1(n3550), .A2(n4630), .ZN(n2974) );
  NOR2_X1 U3810 ( .A1(n4630), .A2(n3551), .ZN(n2978) );
  AOI21_X1 U3811 ( .B1(n2979), .B2(n3513), .A(n2978), .ZN(n3016) );
  INV_X1 U3812 ( .A(n3016), .ZN(n2980) );
  INV_X1 U3813 ( .A(n2981), .ZN(n2982) );
  NAND2_X1 U3814 ( .A1(n2984), .A2(n2983), .ZN(n2985) );
  OAI211_X1 U3815 ( .C1(n2986), .C2(n2985), .A(n3019), .B(n4427), .ZN(n2993)
         );
  NAND2_X1 U3816 ( .A1(n3836), .A2(n2987), .ZN(n2988) );
  OR2_X1 U3817 ( .A1(n2989), .A2(n2988), .ZN(n4417) );
  OAI22_X1 U3818 ( .A1(n4617), .A2(n3672), .B1(n2990), .B2(n4417), .ZN(n2991)
         );
  AOI21_X1 U3819 ( .B1(n4612), .B2(n3682), .A(n2991), .ZN(n2992) );
  OAI211_X1 U3820 ( .C1(n2995), .C2(n2994), .A(n2993), .B(n2992), .ZN(U3219)
         );
  NOR2_X1 U3821 ( .A1(n4629), .A2(n2996), .ZN(n4659) );
  INV_X1 U3822 ( .A(n2997), .ZN(n2999) );
  INV_X1 U3823 ( .A(n4621), .ZN(n3081) );
  NAND2_X1 U3824 ( .A1(n4614), .A2(n4629), .ZN(n3756) );
  NAND2_X1 U3825 ( .A1(n3756), .A2(n3754), .ZN(n4660) );
  OAI21_X1 U3826 ( .B1(n3081), .B2(n4625), .A(n4660), .ZN(n2998) );
  OAI21_X1 U3827 ( .B1(n2950), .B2(n4616), .A(n2998), .ZN(n4658) );
  AOI21_X1 U3828 ( .B1(n4659), .B2(n2999), .A(n4658), .ZN(n3014) );
  NAND2_X1 U3829 ( .A1(n3001), .A2(n3000), .ZN(n3002) );
  NOR2_X1 U3830 ( .A1(n3003), .A2(n3002), .ZN(n3005) );
  NAND3_X1 U3831 ( .A1(n3006), .A2(n3005), .A3(n3004), .ZN(n3007) );
  NAND2_X1 U3832 ( .A1(n3008), .A2(n4143), .ZN(n3101) );
  INV_X1 U3833 ( .A(n3101), .ZN(n3009) );
  NAND2_X1 U3834 ( .A1(n4172), .A2(n3009), .ZN(n4227) );
  INV_X1 U3835 ( .A(n4227), .ZN(n4633) );
  INV_X1 U3836 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3010) );
  OAI22_X1 U3837 ( .A1(n4172), .A2(n3011), .B1(n3010), .B2(n4171), .ZN(n3012)
         );
  AOI21_X1 U3838 ( .B1(n4660), .B2(n4633), .A(n3012), .ZN(n3013) );
  OAI21_X1 U3839 ( .B1(n3014), .B2(n4626), .A(n3013), .ZN(U3290) );
  XNOR2_X1 U3840 ( .A(n3015), .B(n3399), .ZN(n3028) );
  AOI22_X1 U3841 ( .A1(n3853), .A2(n3513), .B1(n3479), .B2(n3048), .ZN(n3029)
         );
  XNOR2_X1 U3842 ( .A(n3028), .B(n3029), .ZN(n3021) );
  OR2_X1 U3843 ( .A1(n3017), .A2(n3016), .ZN(n3018) );
  AOI21_X1 U3844 ( .B1(n3021), .B2(n3020), .A(n3027), .ZN(n3026) );
  AOI22_X1 U3845 ( .A1(n4421), .A2(n3852), .B1(n3681), .B2(n2979), .ZN(n3022)
         );
  OAI21_X1 U3846 ( .B1(n4416), .B2(n3055), .A(n3022), .ZN(n3023) );
  AOI21_X1 U3847 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3024), .A(n3023), .ZN(n3025)
         );
  OAI21_X1 U3848 ( .B1(n3026), .B2(n3678), .A(n3025), .ZN(U3234) );
  AOI22_X1 U3849 ( .A1(n3852), .A2(n3513), .B1(n3479), .B2(n3763), .ZN(n3128)
         );
  NAND2_X1 U3850 ( .A1(n3852), .A2(n3479), .ZN(n3031) );
  NAND2_X1 U3851 ( .A1(n3763), .A2(n2932), .ZN(n3030) );
  NAND2_X1 U3852 ( .A1(n3031), .A2(n3030), .ZN(n3032) );
  XNOR2_X1 U3853 ( .A(n3032), .B(n3399), .ZN(n3130) );
  XOR2_X1 U3854 ( .A(n3128), .B(n3130), .Z(n3131) );
  XNOR2_X1 U3855 ( .A(n3132), .B(n3131), .ZN(n3043) );
  NAND2_X1 U3856 ( .A1(n3034), .A2(n3033), .ZN(n3035) );
  OAI21_X1 U3857 ( .B1(n3036), .B2(n3035), .A(STATE_REG_SCAN_IN), .ZN(n3038)
         );
  AOI21_X1 U3858 ( .B1(n4421), .B2(n3851), .A(n3039), .ZN(n3041) );
  AOI22_X1 U3859 ( .A1(n3682), .A2(n3763), .B1(n3681), .B2(n3853), .ZN(n3040)
         );
  OAI211_X1 U3860 ( .C1(n4432), .C2(REG3_REG_3__SCAN_IN), .A(n3041), .B(n3040), 
        .ZN(n3042) );
  AOI21_X1 U3861 ( .B1(n3043), .B2(n4427), .A(n3042), .ZN(n3044) );
  INV_X1 U3862 ( .A(n3044), .ZN(U3215) );
  NAND2_X1 U3863 ( .A1(n3046), .A2(n2795), .ZN(n3047) );
  NAND2_X1 U3864 ( .A1(n3045), .A2(n3047), .ZN(n4667) );
  AND2_X1 U3865 ( .A1(n4628), .A2(n3048), .ZN(n3049) );
  OR2_X1 U3866 ( .A1(n3049), .A2(n3072), .ZN(n4668) );
  NOR2_X1 U3867 ( .A1(n4694), .A2(n4143), .ZN(n3050) );
  OAI22_X1 U3868 ( .A1(n4668), .A2(n4160), .B1(n3051), .B2(n4171), .ZN(n3061)
         );
  NAND3_X1 U3869 ( .A1(n2794), .A2(n3758), .A3(n4609), .ZN(n3052) );
  NAND2_X1 U3870 ( .A1(n3066), .A2(n3052), .ZN(n3057) );
  NAND2_X1 U3871 ( .A1(n2979), .A2(n4613), .ZN(n3054) );
  NAND2_X1 U3872 ( .A1(n3852), .A2(n4317), .ZN(n3053) );
  OAI211_X1 U3873 ( .C1(n4328), .C2(n3055), .A(n3054), .B(n3053), .ZN(n3056)
         );
  AOI21_X1 U3874 ( .B1(n3057), .B2(n4625), .A(n3056), .ZN(n3059) );
  NAND2_X1 U3875 ( .A1(n4667), .A2(n3081), .ZN(n3058) );
  NAND2_X1 U3876 ( .A1(n3059), .A2(n3058), .ZN(n4666) );
  MUX2_X1 U3877 ( .A(n4666), .B(REG2_REG_2__SCAN_IN), .S(n4626), .Z(n3060) );
  AOI211_X1 U3878 ( .C1(n4633), .C2(n4667), .A(n3061), .B(n3060), .ZN(n3062)
         );
  INV_X1 U3879 ( .A(n3062), .ZN(U3288) );
  XNOR2_X1 U3880 ( .A(n3063), .B(n3065), .ZN(n3116) );
  INV_X1 U3881 ( .A(n3116), .ZN(n3071) );
  AOI22_X1 U3882 ( .A1(n3851), .A2(n4317), .B1(n4611), .B2(n3763), .ZN(n3064)
         );
  OAI21_X1 U3883 ( .B1(n4617), .B2(n4320), .A(n3064), .ZN(n3070) );
  INV_X1 U3884 ( .A(n3065), .ZN(n3748) );
  NAND3_X1 U3885 ( .A1(n3066), .A2(n3759), .A3(n3748), .ZN(n3067) );
  AND2_X1 U3886 ( .A1(n3068), .A2(n3067), .ZN(n3069) );
  OAI22_X1 U3887 ( .A1(n3116), .A2(n4621), .B1(n3069), .B2(n4333), .ZN(n3105)
         );
  AOI211_X1 U3888 ( .C1(n4689), .C2(n3071), .A(n3070), .B(n3105), .ZN(n3077)
         );
  INV_X1 U3889 ( .A(n3072), .ZN(n3074) );
  INV_X1 U3890 ( .A(n3078), .ZN(n3073) );
  AOI21_X1 U3891 ( .B1(n3763), .B2(n3074), .A(n3073), .ZN(n3109) );
  INV_X1 U3892 ( .A(n4402), .ZN(n4669) );
  AOI22_X1 U3893 ( .A1(n3109), .A2(n4669), .B1(REG0_REG_3__SCAN_IN), .B2(n4699), .ZN(n3075) );
  OAI21_X1 U3894 ( .B1(n3077), .B2(n4699), .A(n3075), .ZN(U3473) );
  INV_X1 U3895 ( .A(n4339), .ZN(n4705) );
  AOI22_X1 U3896 ( .A1(n3109), .A2(n4705), .B1(REG1_REG_3__SCAN_IN), .B2(n4714), .ZN(n3076) );
  OAI21_X1 U3897 ( .B1(n3077), .B2(n4714), .A(n3076), .ZN(U3521) );
  AOI21_X1 U3898 ( .B1(n3078), .B2(n3385), .A(n4694), .ZN(n3079) );
  NAND2_X1 U3899 ( .A1(n3079), .A2(n3095), .ZN(n4672) );
  NOR2_X1 U3900 ( .A1(n4672), .A2(n4143), .ZN(n3089) );
  XNOR2_X1 U3901 ( .A(n3080), .B(n2284), .ZN(n4671) );
  NAND2_X1 U3902 ( .A1(n4671), .A2(n3081), .ZN(n3088) );
  XNOR2_X1 U3903 ( .A(n3082), .B(n2284), .ZN(n3086) );
  NAND2_X1 U3904 ( .A1(n3852), .A2(n4613), .ZN(n3084) );
  NAND2_X1 U3905 ( .A1(n3850), .A2(n4317), .ZN(n3083) );
  OAI211_X1 U3906 ( .C1(n4328), .C2(n3133), .A(n3084), .B(n3083), .ZN(n3085)
         );
  AOI21_X1 U3907 ( .B1(n3086), .B2(n4625), .A(n3085), .ZN(n3087) );
  NAND2_X1 U3908 ( .A1(n3088), .A2(n3087), .ZN(n4675) );
  AOI211_X1 U3909 ( .C1(n4627), .C2(n3383), .A(n3089), .B(n4675), .ZN(n3091)
         );
  AOI22_X1 U3910 ( .A1(n4671), .A2(n4633), .B1(REG2_REG_4__SCAN_IN), .B2(n4626), .ZN(n3090) );
  OAI21_X1 U3911 ( .B1(n3091), .B2(n4626), .A(n3090), .ZN(U3286) );
  INV_X1 U3912 ( .A(n3092), .ZN(n3768) );
  XOR2_X1 U3913 ( .A(n3741), .B(n3093), .Z(n3094) );
  NAND2_X1 U3914 ( .A1(n3094), .A2(n4625), .ZN(n3159) );
  AND2_X1 U3915 ( .A1(n3095), .A2(n3157), .ZN(n3096) );
  NOR2_X1 U3916 ( .A1(n3119), .A2(n3096), .ZN(n3164) );
  AND2_X1 U3917 ( .A1(n4172), .A2(n4613), .ZN(n4216) );
  INV_X1 U3918 ( .A(n4216), .ZN(n3229) );
  NAND2_X1 U3919 ( .A1(n4172), .A2(n4611), .ZN(n4221) );
  INV_X1 U3920 ( .A(n4221), .ZN(n4157) );
  AND2_X1 U3921 ( .A1(n4172), .A2(n4317), .ZN(n4214) );
  AOI22_X1 U3922 ( .A1(n4157), .A2(n3157), .B1(n4214), .B2(n3849), .ZN(n3097)
         );
  OAI21_X1 U3923 ( .B1(n3160), .B2(n3229), .A(n3097), .ZN(n3099) );
  OAI22_X1 U3924 ( .A1(n3156), .A2(n4171), .B1(n2567), .B2(n4172), .ZN(n3098)
         );
  AOI211_X1 U3925 ( .C1(n3164), .C2(n4632), .A(n3099), .B(n3098), .ZN(n3104)
         );
  XNOR2_X1 U3926 ( .A(n3100), .B(n3741), .ZN(n3162) );
  NAND2_X1 U3927 ( .A1(n4621), .A2(n3101), .ZN(n3102) );
  NAND2_X1 U3928 ( .A1(n3162), .A2(n4191), .ZN(n3103) );
  OAI211_X1 U3929 ( .C1(n3159), .C2(n4626), .A(n3104), .B(n3103), .ZN(U3285)
         );
  NAND2_X1 U3930 ( .A1(n3105), .A2(n4172), .ZN(n3115) );
  AOI22_X1 U3931 ( .A1(n4626), .A2(REG2_REG_3__SCAN_IN), .B1(n4627), .B2(n3106), .ZN(n3107) );
  OAI21_X1 U3932 ( .B1(n3108), .B2(n4221), .A(n3107), .ZN(n3113) );
  INV_X1 U3933 ( .A(n3109), .ZN(n3111) );
  INV_X1 U3934 ( .A(n4214), .ZN(n3110) );
  OAI22_X1 U3935 ( .A1(n3111), .A2(n4160), .B1(n3160), .B2(n3110), .ZN(n3112)
         );
  AOI211_X1 U3936 ( .C1(n4216), .C2(n3853), .A(n3113), .B(n3112), .ZN(n3114)
         );
  OAI211_X1 U3937 ( .C1(n3116), .C2(n4227), .A(n3115), .B(n3114), .ZN(U3287)
         );
  NAND2_X1 U3938 ( .A1(n3771), .A2(n3779), .ZN(n3720) );
  XOR2_X1 U3939 ( .A(n3720), .B(n3117), .Z(n3185) );
  XOR2_X1 U3940 ( .A(n3720), .B(n3118), .Z(n3183) );
  NAND2_X1 U3941 ( .A1(n4172), .A2(n4625), .ZN(n4105) );
  INV_X1 U3942 ( .A(n4105), .ZN(n3126) );
  NOR2_X1 U3943 ( .A1(n3119), .A2(n3170), .ZN(n3120) );
  OR2_X1 U3944 ( .A1(n3192), .A2(n3120), .ZN(n3188) );
  INV_X1 U3945 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3121) );
  OAI22_X1 U3946 ( .A1(n4172), .A2(n3121), .B1(n3175), .B2(n4171), .ZN(n3122)
         );
  AOI21_X1 U3947 ( .B1(n3179), .B2(n4157), .A(n3122), .ZN(n3124) );
  AOI22_X1 U3948 ( .A1(n4214), .A2(n3848), .B1(n4216), .B2(n3850), .ZN(n3123)
         );
  OAI211_X1 U3949 ( .C1(n3188), .C2(n4160), .A(n3124), .B(n3123), .ZN(n3125)
         );
  AOI21_X1 U3950 ( .B1(n3183), .B2(n3126), .A(n3125), .ZN(n3127) );
  OAI21_X1 U3951 ( .B1(n4177), .B2(n3185), .A(n3127), .ZN(U3284) );
  INV_X1 U3952 ( .A(n3128), .ZN(n3129) );
  OAI22_X1 U3953 ( .A1(n3132), .A2(n3131), .B1(n3130), .B2(n3129), .ZN(n3146)
         );
  NOR2_X1 U3954 ( .A1(n3133), .A2(n3551), .ZN(n3134) );
  AOI21_X1 U3955 ( .B1(n3851), .B2(n3513), .A(n3134), .ZN(n3139) );
  NAND2_X1 U3956 ( .A1(n3851), .A2(n3479), .ZN(n3136) );
  NAND2_X1 U3957 ( .A1(n3385), .A2(n2932), .ZN(n3135) );
  NAND2_X1 U3958 ( .A1(n3136), .A2(n3135), .ZN(n3137) );
  NOR2_X1 U3959 ( .A1(n3146), .A2(n3382), .ZN(n3381) );
  INV_X1 U3960 ( .A(n3138), .ZN(n3140) );
  NOR2_X1 U3961 ( .A1(n3140), .A2(n3139), .ZN(n3147) );
  OR2_X1 U3962 ( .A1(n3381), .A2(n3147), .ZN(n3151) );
  AOI22_X1 U3963 ( .A1(n3850), .A2(n3479), .B1(n2932), .B2(n3157), .ZN(n3141)
         );
  XNOR2_X1 U3964 ( .A(n3141), .B(n3399), .ZN(n3167) );
  NOR2_X1 U3965 ( .A1(n3152), .A2(n3551), .ZN(n3142) );
  AOI21_X1 U3966 ( .B1(n3850), .B2(n3513), .A(n3142), .ZN(n3168) );
  XNOR2_X1 U3967 ( .A(n3167), .B(n3143), .ZN(n3150) );
  INV_X1 U3968 ( .A(n3382), .ZN(n3144) );
  NOR2_X1 U3969 ( .A1(n3146), .A2(n3145), .ZN(n3149) );
  AND2_X1 U3970 ( .A1(n3150), .A2(n3147), .ZN(n3148) );
  OAI211_X1 U3971 ( .C1(n3151), .C2(n3150), .A(n2260), .B(n4427), .ZN(n3155)
         );
  INV_X1 U3972 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4867) );
  NOR2_X1 U3973 ( .A1(STATE_REG_SCAN_IN), .A2(n4867), .ZN(n4446) );
  OAI22_X1 U3974 ( .A1(n3200), .A2(n3672), .B1(n4416), .B2(n3152), .ZN(n3153)
         );
  AOI211_X1 U3975 ( .C1(n3681), .C2(n3851), .A(n4446), .B(n3153), .ZN(n3154)
         );
  OAI211_X1 U3976 ( .C1(n4432), .C2(n3156), .A(n3155), .B(n3154), .ZN(U3224)
         );
  AOI22_X1 U3977 ( .A1(n3849), .A2(n4317), .B1(n4611), .B2(n3157), .ZN(n3158)
         );
  OAI211_X1 U3978 ( .C1(n3160), .C2(n4320), .A(n3159), .B(n3158), .ZN(n3161)
         );
  AOI21_X1 U3979 ( .B1(n3162), .B2(n4678), .A(n3161), .ZN(n3166) );
  AOI22_X1 U3980 ( .A1(n3164), .A2(n4705), .B1(REG1_REG_5__SCAN_IN), .B2(n4714), .ZN(n3163) );
  OAI21_X1 U3981 ( .B1(n3166), .B2(n4714), .A(n3163), .ZN(U3523) );
  AOI22_X1 U3982 ( .A1(n3164), .A2(n4669), .B1(REG0_REG_5__SCAN_IN), .B2(n4699), .ZN(n3165) );
  OAI21_X1 U3983 ( .B1(n3166), .B2(n4699), .A(n3165), .ZN(U3477) );
  AOI22_X1 U3984 ( .A1(n3849), .A2(n3479), .B1(n2932), .B2(n3179), .ZN(n3169)
         );
  XOR2_X1 U3985 ( .A(n3399), .B(n3169), .Z(n3205) );
  OAI22_X1 U3986 ( .A1(n3200), .A2(n3548), .B1(n3551), .B2(n3170), .ZN(n3206)
         );
  XNOR2_X1 U3987 ( .A(n3205), .B(n3206), .ZN(n3171) );
  XNOR2_X1 U3988 ( .A(n3207), .B(n3171), .ZN(n3177) );
  NOR2_X1 U3989 ( .A1(STATE_REG_SCAN_IN), .A2(n3172), .ZN(n4457) );
  AOI21_X1 U3990 ( .B1(n3681), .B2(n3850), .A(n4457), .ZN(n3174) );
  AOI22_X1 U3991 ( .A1(n3682), .A2(n3179), .B1(n4421), .B2(n3848), .ZN(n3173)
         );
  OAI211_X1 U3992 ( .C1(n4432), .C2(n3175), .A(n3174), .B(n3173), .ZN(n3176)
         );
  AOI21_X1 U3993 ( .B1(n3177), .B2(n4427), .A(n3176), .ZN(n3178) );
  INV_X1 U3994 ( .A(n3178), .ZN(U3236) );
  INV_X1 U3995 ( .A(n4678), .ZN(n4301) );
  AOI22_X1 U3996 ( .A1(n3848), .A2(n4317), .B1(n3179), .B2(n4611), .ZN(n3180)
         );
  OAI21_X1 U3997 ( .B1(n3181), .B2(n4320), .A(n3180), .ZN(n3182) );
  AOI21_X1 U3998 ( .B1(n3183), .B2(n4625), .A(n3182), .ZN(n3184) );
  OAI21_X1 U3999 ( .B1(n3185), .B2(n4301), .A(n3184), .ZN(n3190) );
  INV_X1 U4000 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4456) );
  OAI22_X1 U4001 ( .A1(n3188), .A2(n4339), .B1(n4717), .B2(n4456), .ZN(n3186)
         );
  AOI21_X1 U4002 ( .B1(n3190), .B2(n4717), .A(n3186), .ZN(n3187) );
  INV_X1 U4003 ( .A(n3187), .ZN(U3524) );
  OAI22_X1 U4004 ( .A1(n3188), .A2(n4402), .B1(n4701), .B2(n2576), .ZN(n3189)
         );
  AOI21_X1 U4005 ( .B1(n3190), .B2(n4701), .A(n3189), .ZN(n3191) );
  INV_X1 U4006 ( .A(n3191), .ZN(U3479) );
  INV_X1 U4007 ( .A(n3192), .ZN(n3194) );
  INV_X1 U4008 ( .A(n3193), .ZN(n3243) );
  AOI211_X1 U4009 ( .C1(n3213), .C2(n3194), .A(n4694), .B(n3243), .ZN(n4677)
         );
  INV_X1 U4010 ( .A(n3722), .ZN(n3195) );
  XNOR2_X1 U4011 ( .A(n3196), .B(n3195), .ZN(n3197) );
  NAND2_X1 U4012 ( .A1(n3197), .A2(n4625), .ZN(n3199) );
  AOI22_X1 U4013 ( .A1(n3847), .A2(n4317), .B1(n4611), .B2(n3213), .ZN(n3198)
         );
  OAI211_X1 U4014 ( .C1(n3200), .C2(n4320), .A(n3199), .B(n3198), .ZN(n4676)
         );
  AOI21_X1 U4015 ( .B1(n4677), .B2(n3940), .A(n4676), .ZN(n3204) );
  XOR2_X1 U4016 ( .A(n3201), .B(n3722), .Z(n4679) );
  OAI22_X1 U4017 ( .A1(n4172), .A2(n2590), .B1(n3216), .B2(n4171), .ZN(n3202)
         );
  AOI21_X1 U4018 ( .B1(n4679), .B2(n4191), .A(n3202), .ZN(n3203) );
  OAI21_X1 U4019 ( .B1(n3204), .B2(n4626), .A(n3203), .ZN(U3283) );
  INV_X1 U4020 ( .A(n3206), .ZN(n3208) );
  AOI22_X1 U4021 ( .A1(n3848), .A2(n3479), .B1(n2932), .B2(n3213), .ZN(n3209)
         );
  XNOR2_X1 U4022 ( .A(n3209), .B(n3399), .ZN(n3252) );
  NOR2_X1 U4023 ( .A1(n3210), .A2(n3551), .ZN(n3211) );
  AOI21_X1 U4024 ( .B1(n3848), .B2(n3513), .A(n3211), .ZN(n3251) );
  XOR2_X1 U4025 ( .A(n3252), .B(n3251), .Z(n3249) );
  XOR2_X1 U4026 ( .A(n3250), .B(n3249), .Z(n3218) );
  INV_X1 U4027 ( .A(REG3_REG_7__SCAN_IN), .ZN(n3212) );
  NOR2_X1 U4028 ( .A1(STATE_REG_SCAN_IN), .A2(n3212), .ZN(n4467) );
  AOI21_X1 U4029 ( .B1(n4421), .B2(n3847), .A(n4467), .ZN(n3215) );
  AOI22_X1 U4030 ( .A1(n3682), .A2(n3213), .B1(n3681), .B2(n3849), .ZN(n3214)
         );
  OAI211_X1 U4031 ( .C1(n4432), .C2(n3216), .A(n3215), .B(n3214), .ZN(n3217)
         );
  AOI21_X1 U4032 ( .B1(n3218), .B2(n4427), .A(n3217), .ZN(n3219) );
  INV_X1 U4033 ( .A(n3219), .ZN(U3210) );
  INV_X1 U4034 ( .A(n3220), .ZN(n3788) );
  AND2_X1 U4035 ( .A1(n3788), .A2(n3776), .ZN(n3742) );
  INV_X1 U4036 ( .A(n3742), .ZN(n3221) );
  XNOR2_X1 U4037 ( .A(n3222), .B(n3221), .ZN(n3223) );
  NAND2_X1 U4038 ( .A1(n3223), .A2(n4625), .ZN(n3287) );
  XOR2_X1 U4039 ( .A(n3742), .B(n3224), .Z(n3290) );
  NAND2_X1 U4040 ( .A1(n3290), .A2(n4191), .ZN(n3234) );
  INV_X1 U4041 ( .A(n3305), .ZN(n3226) );
  OAI21_X1 U4042 ( .B1(n4680), .B2(n3227), .A(n3226), .ZN(n3296) );
  INV_X1 U40430 ( .A(n3296), .ZN(n3232) );
  OAI22_X1 U4044 ( .A1(n3281), .A2(n4171), .B1(n2609), .B2(n4172), .ZN(n3231)
         );
  AOI22_X1 U4045 ( .A1(n4157), .A2(n3285), .B1(n4214), .B2(n4593), .ZN(n3228)
         );
  OAI21_X1 U4046 ( .B1(n3288), .B2(n3229), .A(n3228), .ZN(n3230) );
  AOI211_X1 U4047 ( .C1(n3232), .C2(n4632), .A(n3231), .B(n3230), .ZN(n3233)
         );
  OAI211_X1 U4048 ( .C1(n4626), .C2(n3287), .A(n3234), .B(n3233), .ZN(U3281)
         );
  NAND2_X1 U4049 ( .A1(n3775), .A2(n3780), .ZN(n3719) );
  XNOR2_X1 U4050 ( .A(n3235), .B(n3719), .ZN(n3242) );
  XNOR2_X1 U4051 ( .A(n3236), .B(n3719), .ZN(n3240) );
  AOI22_X1 U4052 ( .A1(n3846), .A2(n4317), .B1(n3265), .B2(n4611), .ZN(n3237)
         );
  OAI21_X1 U4053 ( .B1(n3238), .B2(n4320), .A(n3237), .ZN(n3239) );
  AOI21_X1 U4054 ( .B1(n3240), .B2(n4625), .A(n3239), .ZN(n3241) );
  OAI21_X1 U4055 ( .B1(n3242), .B2(n4621), .A(n3241), .ZN(n4682) );
  INV_X1 U4056 ( .A(n4682), .ZN(n3248) );
  INV_X1 U4057 ( .A(n3242), .ZN(n4684) );
  NOR2_X1 U4058 ( .A1(n3243), .A2(n3258), .ZN(n4681) );
  NOR3_X1 U4059 ( .A1(n4681), .A2(n4680), .A3(n4160), .ZN(n3246) );
  OAI22_X1 U4060 ( .A1(n4172), .A2(n3244), .B1(n3268), .B2(n4171), .ZN(n3245)
         );
  AOI211_X1 U4061 ( .C1(n4684), .C2(n4633), .A(n3246), .B(n3245), .ZN(n3247)
         );
  OAI21_X1 U4062 ( .B1(n3248), .B2(n4626), .A(n3247), .ZN(U3282) );
  NAND2_X1 U4063 ( .A1(n3250), .A2(n3249), .ZN(n3254) );
  NAND2_X1 U4064 ( .A1(n3847), .A2(n3479), .ZN(n3256) );
  NAND2_X1 U4065 ( .A1(n3265), .A2(n2932), .ZN(n3255) );
  NAND2_X1 U4066 ( .A1(n3256), .A2(n3255), .ZN(n3257) );
  XNOR2_X1 U4067 ( .A(n3257), .B(n3277), .ZN(n3261) );
  NOR2_X1 U4068 ( .A1(n3258), .A2(n3551), .ZN(n3259) );
  AOI21_X1 U4069 ( .B1(n3847), .B2(n3513), .A(n3259), .ZN(n3260) );
  NOR2_X1 U4070 ( .A1(n3261), .A2(n3260), .ZN(n3273) );
  INV_X1 U4071 ( .A(n3273), .ZN(n3262) );
  NAND2_X1 U4072 ( .A1(n3261), .A2(n3260), .ZN(n3272) );
  NAND2_X1 U4073 ( .A1(n3262), .A2(n3272), .ZN(n3263) );
  XNOR2_X1 U4074 ( .A(n3274), .B(n3263), .ZN(n3270) );
  NAND2_X1 U4075 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4477) );
  INV_X1 U4076 ( .A(n4477), .ZN(n3264) );
  AOI21_X1 U4077 ( .B1(n4421), .B2(n3846), .A(n3264), .ZN(n3267) );
  AOI22_X1 U4078 ( .A1(n3682), .A2(n3265), .B1(n3681), .B2(n3848), .ZN(n3266)
         );
  OAI211_X1 U4079 ( .C1(n4432), .C2(n3268), .A(n3267), .B(n3266), .ZN(n3269)
         );
  AOI21_X1 U4080 ( .B1(n3270), .B2(n4427), .A(n3269), .ZN(n3271) );
  INV_X1 U4081 ( .A(n3271), .ZN(U3218) );
  OAI21_X2 U4082 ( .B1(n3274), .B2(n3273), .A(n3272), .ZN(n3317) );
  NAND2_X1 U4083 ( .A1(n3846), .A2(n3479), .ZN(n3276) );
  NAND2_X1 U4084 ( .A1(n3285), .A2(n2932), .ZN(n3275) );
  NAND2_X1 U4085 ( .A1(n3276), .A2(n3275), .ZN(n3278) );
  XNOR2_X1 U4086 ( .A(n3278), .B(n3399), .ZN(n3318) );
  AOI22_X1 U4087 ( .A1(n3846), .A2(n3513), .B1(n3479), .B2(n3285), .ZN(n3319)
         );
  XNOR2_X1 U4088 ( .A(n3318), .B(n3319), .ZN(n3316) );
  XNOR2_X1 U4089 ( .A(n3317), .B(n3316), .ZN(n3283) );
  NOR2_X1 U4090 ( .A1(STATE_REG_SCAN_IN), .A2(n2610), .ZN(n4493) );
  AOI21_X1 U4091 ( .B1(n4421), .B2(n4593), .A(n4493), .ZN(n3280) );
  AOI22_X1 U4092 ( .A1(n3682), .A2(n3285), .B1(n3681), .B2(n3847), .ZN(n3279)
         );
  OAI211_X1 U4093 ( .C1(n4432), .C2(n3281), .A(n3280), .B(n3279), .ZN(n3282)
         );
  AOI21_X1 U4094 ( .B1(n3283), .B2(n4427), .A(n3282), .ZN(n3284) );
  INV_X1 U4095 ( .A(n3284), .ZN(U3228) );
  INV_X1 U4096 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4097 ( .A1(n4593), .A2(n4317), .B1(n4611), .B2(n3285), .ZN(n3286)
         );
  OAI211_X1 U4098 ( .C1(n3288), .C2(n4320), .A(n3287), .B(n3286), .ZN(n3289)
         );
  AOI21_X1 U4099 ( .B1(n3290), .B2(n4678), .A(n3289), .ZN(n3293) );
  MUX2_X1 U4100 ( .A(n3291), .B(n3293), .S(n4701), .Z(n3292) );
  OAI21_X1 U4101 ( .B1(n3296), .B2(n4402), .A(n3292), .ZN(U3485) );
  MUX2_X1 U4102 ( .A(n3294), .B(n3293), .S(n4717), .Z(n3295) );
  OAI21_X1 U4103 ( .B1(n4339), .B2(n3296), .A(n3295), .ZN(U3527) );
  AND2_X1 U4104 ( .A1(n3786), .A2(n3790), .ZN(n3740) );
  XOR2_X1 U4105 ( .A(n3740), .B(n3297), .Z(n3304) );
  XNOR2_X1 U4106 ( .A(n3298), .B(n3740), .ZN(n3302) );
  AOI22_X1 U4107 ( .A1(n3845), .A2(n4317), .B1(n4611), .B2(n3327), .ZN(n3299)
         );
  OAI21_X1 U4108 ( .B1(n3300), .B2(n4320), .A(n3299), .ZN(n3301) );
  AOI21_X1 U4109 ( .B1(n3302), .B2(n4625), .A(n3301), .ZN(n3303) );
  OAI21_X1 U4110 ( .B1(n3304), .B2(n4621), .A(n3303), .ZN(n4687) );
  INV_X1 U4111 ( .A(n4687), .ZN(n3310) );
  INV_X1 U4112 ( .A(n3304), .ZN(n4690) );
  NOR2_X1 U4113 ( .A1(n3305), .A2(n3314), .ZN(n4686) );
  NOR3_X1 U4114 ( .A1(n4686), .A2(n4685), .A3(n4160), .ZN(n3308) );
  OAI22_X1 U4115 ( .A1(n4172), .A2(n3306), .B1(n3330), .B2(n4171), .ZN(n3307)
         );
  AOI211_X1 U4116 ( .C1(n4690), .C2(n4633), .A(n3308), .B(n3307), .ZN(n3309)
         );
  OAI21_X1 U4117 ( .B1(n3310), .B2(n4626), .A(n3309), .ZN(U3280) );
  NAND2_X1 U4118 ( .A1(n4593), .A2(n3479), .ZN(n3312) );
  NAND2_X1 U4119 ( .A1(n3327), .A2(n2932), .ZN(n3311) );
  NAND2_X1 U4120 ( .A1(n3312), .A2(n3311), .ZN(n3313) );
  XNOR2_X1 U4121 ( .A(n3313), .B(n3399), .ZN(n3335) );
  NOR2_X1 U4122 ( .A1(n3314), .A2(n3551), .ZN(n3315) );
  AOI21_X1 U4123 ( .B1(n4593), .B2(n3513), .A(n3315), .ZN(n3333) );
  XOR2_X1 U4124 ( .A(n3335), .B(n3333), .Z(n3325) );
  INV_X1 U4125 ( .A(n3318), .ZN(n3320) );
  NAND2_X1 U4126 ( .A1(n3320), .A2(n3319), .ZN(n3321) );
  INV_X1 U4127 ( .A(n3337), .ZN(n3324) );
  AOI211_X1 U4128 ( .C1(n3325), .C2(n3322), .A(n3678), .B(n3324), .ZN(n3332)
         );
  NAND2_X1 U4129 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4498) );
  INV_X1 U4130 ( .A(n4498), .ZN(n3326) );
  AOI21_X1 U4131 ( .B1(n3681), .B2(n3846), .A(n3326), .ZN(n3329) );
  AOI22_X1 U4132 ( .A1(n3682), .A2(n3327), .B1(n4421), .B2(n3845), .ZN(n3328)
         );
  OAI211_X1 U4133 ( .C1(n4432), .C2(n3330), .A(n3329), .B(n3328), .ZN(n3331)
         );
  OR2_X1 U4134 ( .A1(n3332), .A2(n3331), .ZN(U3214) );
  INV_X1 U4135 ( .A(n3333), .ZN(n3334) );
  NAND2_X1 U4136 ( .A1(n3335), .A2(n3334), .ZN(n3336) );
  AOI22_X1 U4137 ( .A1(n3845), .A2(n3479), .B1(n2932), .B2(n4592), .ZN(n3338)
         );
  XOR2_X1 U4138 ( .A(n3399), .B(n3338), .Z(n3394) );
  OAI22_X1 U4139 ( .A1(n3373), .A2(n3548), .B1(n3551), .B2(n4604), .ZN(n3395)
         );
  XNOR2_X1 U4140 ( .A(n3394), .B(n3395), .ZN(n3339) );
  XNOR2_X1 U4141 ( .A(n3396), .B(n3339), .ZN(n3343) );
  AND2_X1 U4142 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4514) );
  AOI21_X1 U4143 ( .B1(n4421), .B2(n4331), .A(n4514), .ZN(n3341) );
  AOI22_X1 U4144 ( .A1(n3682), .A2(n4592), .B1(n3681), .B2(n4593), .ZN(n3340)
         );
  OAI211_X1 U4145 ( .C1(n4432), .C2(n4601), .A(n3341), .B(n3340), .ZN(n3342)
         );
  AOI21_X1 U4146 ( .B1(n3343), .B2(n4427), .A(n3342), .ZN(n3344) );
  INV_X1 U4147 ( .A(n3344), .ZN(U3233) );
  NAND2_X1 U4148 ( .A1(n3346), .A2(n3345), .ZN(n3348) );
  XNOR2_X1 U4149 ( .A(n3348), .B(n3738), .ZN(n4334) );
  XNOR2_X1 U4150 ( .A(n3349), .B(n3738), .ZN(n4336) );
  NAND2_X1 U4151 ( .A1(n4336), .A2(n4191), .ZN(n3357) );
  INV_X1 U4152 ( .A(n3360), .ZN(n3350) );
  OAI21_X1 U4153 ( .B1(n3350), .B2(n4327), .A(n4210), .ZN(n4403) );
  INV_X1 U4154 ( .A(n4403), .ZN(n3355) );
  AOI22_X1 U4155 ( .A1(n4216), .A2(n4331), .B1(n4214), .B2(n4193), .ZN(n3353)
         );
  INV_X1 U4156 ( .A(n3642), .ZN(n3351) );
  AOI22_X1 U4157 ( .A1(n4626), .A2(REG2_REG_13__SCAN_IN), .B1(n3351), .B2(
        n4627), .ZN(n3352) );
  OAI211_X1 U4158 ( .C1(n4327), .C2(n4221), .A(n3353), .B(n3352), .ZN(n3354)
         );
  AOI21_X1 U4159 ( .B1(n3355), .B2(n4632), .A(n3354), .ZN(n3356) );
  OAI211_X1 U4160 ( .C1(n4334), .C2(n4105), .A(n3357), .B(n3356), .ZN(U3277)
         );
  XNOR2_X1 U4161 ( .A(n4331), .B(n3401), .ZN(n3747) );
  XOR2_X1 U4162 ( .A(n3747), .B(n3358), .Z(n3375) );
  NAND2_X1 U4163 ( .A1(n4603), .A2(n3586), .ZN(n3359) );
  NAND2_X1 U4164 ( .A1(n3360), .A2(n3359), .ZN(n3380) );
  OAI22_X1 U4165 ( .A1(n4172), .A2(n3361), .B1(n3589), .B2(n4171), .ZN(n3362)
         );
  AOI21_X1 U4166 ( .B1(n3586), .B2(n4157), .A(n3362), .ZN(n3364) );
  AOI22_X1 U4167 ( .A1(n4216), .A2(n3845), .B1(n4214), .B2(n4215), .ZN(n3363)
         );
  OAI211_X1 U4168 ( .C1(n3380), .C2(n4160), .A(n3364), .B(n3363), .ZN(n3369)
         );
  INV_X1 U4169 ( .A(n3747), .ZN(n3365) );
  XNOR2_X1 U4170 ( .A(n3366), .B(n3365), .ZN(n3367) );
  NAND2_X1 U4171 ( .A1(n3367), .A2(n4625), .ZN(n3372) );
  NOR2_X1 U4172 ( .A1(n3372), .A2(n4626), .ZN(n3368) );
  AOI211_X1 U4173 ( .C1(n3375), .C2(n4191), .A(n3369), .B(n3368), .ZN(n3370)
         );
  INV_X1 U4174 ( .A(n3370), .ZN(U3278) );
  AOI22_X1 U4175 ( .A1(n4215), .A2(n4317), .B1(n4611), .B2(n3586), .ZN(n3371)
         );
  OAI211_X1 U4176 ( .C1(n3373), .C2(n4320), .A(n3372), .B(n3371), .ZN(n3374)
         );
  AOI21_X1 U4177 ( .B1(n3375), .B2(n4678), .A(n3374), .ZN(n3377) );
  MUX2_X1 U4178 ( .A(n2644), .B(n3377), .S(n4717), .Z(n3376) );
  OAI21_X1 U4179 ( .B1(n3380), .B2(n4339), .A(n3376), .ZN(U3530) );
  INV_X1 U4180 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3378) );
  MUX2_X1 U4181 ( .A(n3378), .B(n3377), .S(n4701), .Z(n3379) );
  OAI21_X1 U4182 ( .B1(n3380), .B2(n4402), .A(n3379), .ZN(U3491) );
  AOI211_X1 U4183 ( .C1(n3382), .C2(n3146), .A(n3678), .B(n3381), .ZN(n3390)
         );
  INV_X1 U4184 ( .A(n3383), .ZN(n3388) );
  AOI21_X1 U4185 ( .B1(n4421), .B2(n3850), .A(n3384), .ZN(n3387) );
  AOI22_X1 U4186 ( .A1(n3682), .A2(n3385), .B1(n3681), .B2(n3852), .ZN(n3386)
         );
  OAI211_X1 U4187 ( .C1(n4432), .C2(n3388), .A(n3387), .B(n3386), .ZN(n3389)
         );
  OR2_X1 U4188 ( .A1(n3390), .A2(n3389), .ZN(U3227) );
  INV_X1 U4189 ( .A(IR_REG_30__SCAN_IN), .ZN(n3392) );
  NAND3_X1 U4190 ( .A1(n3392), .A2(STATE_REG_SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n3393) );
  INV_X1 U4191 ( .A(DATAI_31_), .ZN(n4975) );
  OAI22_X1 U4192 ( .A1(n2312), .A2(n3393), .B1(STATE_REG_SCAN_IN), .B2(n4975), 
        .ZN(U3321) );
  NAND2_X1 U4193 ( .A1(n4331), .A2(n3479), .ZN(n3398) );
  NAND2_X1 U4194 ( .A1(n3586), .A2(n2932), .ZN(n3397) );
  NAND2_X1 U4195 ( .A1(n3398), .A2(n3397), .ZN(n3400) );
  XNOR2_X1 U4196 ( .A(n3400), .B(n3277), .ZN(n3404) );
  NOR2_X1 U4197 ( .A1(n3401), .A2(n3551), .ZN(n3402) );
  AOI21_X1 U4198 ( .B1(n4331), .B2(n3513), .A(n3402), .ZN(n3403) );
  NOR2_X1 U4199 ( .A1(n3404), .A2(n3403), .ZN(n3581) );
  NAND2_X1 U4200 ( .A1(n3404), .A2(n3403), .ZN(n3582) );
  AOI22_X1 U4201 ( .A1(n4215), .A2(n3479), .B1(n2932), .B2(n3639), .ZN(n3407)
         );
  XOR2_X1 U4202 ( .A(n3399), .B(n3407), .Z(n3637) );
  OAI22_X1 U4203 ( .A1(n4321), .A2(n3548), .B1(n3551), .B2(n4327), .ZN(n3636)
         );
  NAND2_X1 U4204 ( .A1(n4193), .A2(n3479), .ZN(n3410) );
  NAND2_X1 U4205 ( .A1(n4316), .A2(n2932), .ZN(n3409) );
  NAND2_X1 U4206 ( .A1(n3410), .A2(n3409), .ZN(n3411) );
  XNOR2_X1 U4207 ( .A(n3411), .B(n3277), .ZN(n3414) );
  NOR2_X1 U4208 ( .A1(n4222), .A2(n3551), .ZN(n3412) );
  AOI21_X1 U4209 ( .B1(n4193), .B2(n3513), .A(n3412), .ZN(n3413) );
  NOR2_X1 U4210 ( .A1(n3414), .A2(n3413), .ZN(n3519) );
  NAND2_X1 U4211 ( .A1(n3414), .A2(n3413), .ZN(n3520) );
  AOI22_X1 U4212 ( .A1(n4318), .A2(n3479), .B1(n2932), .B2(n4307), .ZN(n3415)
         );
  XNOR2_X1 U4213 ( .A(n3415), .B(n3399), .ZN(n3418) );
  NAND2_X1 U4214 ( .A1(n4318), .A2(n3513), .ZN(n3417) );
  NAND2_X1 U4215 ( .A1(n4307), .A2(n3479), .ZN(n3416) );
  NAND2_X1 U4216 ( .A1(n3417), .A2(n3416), .ZN(n4424) );
  NAND2_X1 U4217 ( .A1(n4423), .A2(n4424), .ZN(n3428) );
  NOR2_X1 U4218 ( .A1(n3419), .A2(n3418), .ZN(n3420) );
  NAND2_X1 U4219 ( .A1(n4308), .A2(n3479), .ZN(n3422) );
  NAND2_X1 U4220 ( .A1(n4168), .A2(n2932), .ZN(n3421) );
  NAND2_X1 U4221 ( .A1(n3422), .A2(n3421), .ZN(n3423) );
  XNOR2_X1 U4222 ( .A(n3423), .B(n3399), .ZN(n3427) );
  NAND2_X1 U4223 ( .A1(n4308), .A2(n3513), .ZN(n3425) );
  NAND2_X1 U4224 ( .A1(n4168), .A2(n3479), .ZN(n3424) );
  NAND2_X1 U4225 ( .A1(n3425), .A2(n3424), .ZN(n3426) );
  NOR2_X1 U4226 ( .A1(n3427), .A2(n3426), .ZN(n3429) );
  AOI21_X1 U4227 ( .B1(n3427), .B2(n3426), .A(n3429), .ZN(n4425) );
  INV_X1 U4228 ( .A(n3429), .ZN(n3430) );
  NAND2_X1 U4229 ( .A1(n4420), .A2(n3479), .ZN(n3432) );
  NAND2_X1 U4230 ( .A1(n4292), .A2(n2932), .ZN(n3431) );
  NAND2_X1 U4231 ( .A1(n3432), .A2(n3431), .ZN(n3433) );
  XNOR2_X1 U4232 ( .A(n3433), .B(n3399), .ZN(n3436) );
  NAND2_X1 U4233 ( .A1(n4420), .A2(n3513), .ZN(n3435) );
  NAND2_X1 U4234 ( .A1(n4292), .A2(n3479), .ZN(n3434) );
  NAND2_X1 U4235 ( .A1(n3435), .A2(n3434), .ZN(n3437) );
  NAND2_X1 U4236 ( .A1(n3436), .A2(n3437), .ZN(n3606) );
  INV_X1 U4237 ( .A(n3436), .ZN(n3439) );
  INV_X1 U4238 ( .A(n3437), .ZN(n3438) );
  NAND2_X1 U4239 ( .A1(n3439), .A2(n3438), .ZN(n3605) );
  NAND2_X1 U4240 ( .A1(n4293), .A2(n3479), .ZN(n3441) );
  NAND2_X1 U4241 ( .A1(n4138), .A2(n2932), .ZN(n3440) );
  NAND2_X1 U4242 ( .A1(n3441), .A2(n3440), .ZN(n3442) );
  XNOR2_X1 U4243 ( .A(n3442), .B(n3399), .ZN(n3445) );
  NAND2_X1 U4244 ( .A1(n4293), .A2(n3513), .ZN(n3444) );
  NAND2_X1 U4245 ( .A1(n4138), .A2(n3479), .ZN(n3443) );
  NAND2_X1 U4246 ( .A1(n3444), .A2(n3443), .ZN(n3446) );
  NAND2_X1 U4247 ( .A1(n3445), .A2(n3446), .ZN(n3657) );
  NAND2_X1 U4248 ( .A1(n3656), .A2(n3657), .ZN(n3655) );
  INV_X1 U4249 ( .A(n3445), .ZN(n3448) );
  INV_X1 U4250 ( .A(n3446), .ZN(n3447) );
  NAND2_X1 U4251 ( .A1(n3448), .A2(n3447), .ZN(n3659) );
  NAND2_X1 U4252 ( .A1(n3655), .A2(n3659), .ZN(n3540) );
  NAND2_X1 U4253 ( .A1(n4278), .A2(n3479), .ZN(n3450) );
  NAND2_X1 U4254 ( .A1(n3541), .A2(n2932), .ZN(n3449) );
  NAND2_X1 U4255 ( .A1(n3450), .A2(n3449), .ZN(n3451) );
  XNOR2_X1 U4256 ( .A(n3451), .B(n3399), .ZN(n3452) );
  AOI22_X1 U4257 ( .A1(n4278), .A2(n3513), .B1(n3479), .B2(n3541), .ZN(n3453)
         );
  XNOR2_X1 U4258 ( .A(n3452), .B(n3453), .ZN(n3539) );
  NAND2_X1 U4259 ( .A1(n3540), .A2(n3539), .ZN(n3456) );
  NAND2_X1 U4260 ( .A1(n3456), .A2(n3455), .ZN(n3624) );
  NAND2_X1 U4261 ( .A1(n4079), .A2(n3479), .ZN(n3458) );
  NAND2_X1 U4262 ( .A1(n3629), .A2(n2932), .ZN(n3457) );
  NAND2_X1 U4263 ( .A1(n3458), .A2(n3457), .ZN(n3459) );
  XNOR2_X1 U4264 ( .A(n3459), .B(n3399), .ZN(n3462) );
  NAND2_X1 U4265 ( .A1(n4079), .A2(n3513), .ZN(n3461) );
  NAND2_X1 U4266 ( .A1(n3629), .A2(n3479), .ZN(n3460) );
  NAND2_X1 U4267 ( .A1(n3461), .A2(n3460), .ZN(n3463) );
  NAND2_X1 U4268 ( .A1(n3462), .A2(n3463), .ZN(n3625) );
  NAND2_X1 U4269 ( .A1(n3624), .A2(n3625), .ZN(n3623) );
  INV_X1 U4270 ( .A(n3462), .ZN(n3465) );
  INV_X1 U4271 ( .A(n3463), .ZN(n3464) );
  NAND2_X1 U4272 ( .A1(n3465), .A2(n3464), .ZN(n3627) );
  NAND2_X1 U4273 ( .A1(n4096), .A2(n3479), .ZN(n3467) );
  NAND2_X1 U4274 ( .A1(n4266), .A2(n2932), .ZN(n3466) );
  NAND2_X1 U4275 ( .A1(n3467), .A2(n3466), .ZN(n3468) );
  XNOR2_X1 U4276 ( .A(n3468), .B(n3399), .ZN(n3572) );
  NAND2_X1 U4277 ( .A1(n4096), .A2(n3513), .ZN(n3470) );
  NAND2_X1 U4278 ( .A1(n4266), .A2(n3479), .ZN(n3469) );
  NAND2_X1 U4279 ( .A1(n3470), .A2(n3469), .ZN(n3573) );
  NOR2_X1 U4280 ( .A1(n3572), .A2(n3573), .ZN(n3472) );
  NAND2_X1 U4281 ( .A1(n3572), .A2(n3573), .ZN(n3471) );
  AOI22_X1 U4282 ( .A1(n4267), .A2(n3479), .B1(n2932), .B2(n3474), .ZN(n3473)
         );
  XNOR2_X1 U4283 ( .A(n3473), .B(n3399), .ZN(n3475) );
  AOI22_X1 U4284 ( .A1(n4267), .A2(n3513), .B1(n3479), .B2(n3474), .ZN(n3476)
         );
  XNOR2_X1 U4285 ( .A(n3475), .B(n3476), .ZN(n3648) );
  INV_X1 U4286 ( .A(n3475), .ZN(n3478) );
  INV_X1 U4287 ( .A(n3476), .ZN(n3477) );
  NOR2_X1 U4288 ( .A1(n3478), .A2(n3477), .ZN(n3531) );
  AOI22_X1 U4289 ( .A1(n4055), .A2(n3479), .B1(n2932), .B2(n3534), .ZN(n3480)
         );
  XNOR2_X1 U4290 ( .A(n3480), .B(n3399), .ZN(n3484) );
  NOR2_X1 U4291 ( .A1(n4047), .A2(n3551), .ZN(n3481) );
  AOI21_X1 U4292 ( .B1(n4055), .B2(n3513), .A(n3481), .ZN(n3483) );
  XNOR2_X1 U4293 ( .A(n3484), .B(n3483), .ZN(n3530) );
  NOR2_X1 U4294 ( .A1(n3531), .A2(n3530), .ZN(n3482) );
  OR2_X1 U4295 ( .A1(n3484), .A2(n3483), .ZN(n3489) );
  NOR2_X1 U4296 ( .A1(n4023), .A2(n3551), .ZN(n3485) );
  AOI21_X1 U4297 ( .B1(n4007), .B2(n3513), .A(n3485), .ZN(n3490) );
  AOI22_X1 U4298 ( .A1(n4007), .A2(n3479), .B1(n2932), .B2(n4029), .ZN(n3488)
         );
  XOR2_X1 U4299 ( .A(n3399), .B(n3488), .Z(n3616) );
  NAND2_X1 U4300 ( .A1(n3614), .A2(n3616), .ZN(n3493) );
  NAND2_X1 U4301 ( .A1(n3532), .A2(n3489), .ZN(n3492) );
  INV_X1 U4302 ( .A(n3490), .ZN(n3491) );
  NAND2_X1 U4303 ( .A1(n3492), .A2(n3491), .ZN(n3615) );
  NAND2_X1 U4304 ( .A1(n3493), .A2(n3615), .ZN(n3593) );
  NAND2_X1 U4305 ( .A1(n4026), .A2(n3479), .ZN(n3495) );
  NAND2_X1 U4306 ( .A1(n3596), .A2(n2932), .ZN(n3494) );
  NAND2_X1 U4307 ( .A1(n3495), .A2(n3494), .ZN(n3496) );
  XNOR2_X1 U4308 ( .A(n3496), .B(n3277), .ZN(n3499) );
  NOR2_X1 U4309 ( .A1(n4011), .A2(n3551), .ZN(n3497) );
  AOI21_X1 U4310 ( .B1(n4026), .B2(n3513), .A(n3497), .ZN(n3498) );
  NAND2_X1 U4311 ( .A1(n3499), .A2(n3498), .ZN(n3594) );
  NAND2_X1 U4312 ( .A1(n4237), .A2(n3479), .ZN(n3502) );
  NAND2_X1 U4313 ( .A1(n3500), .A2(n2932), .ZN(n3501) );
  NAND2_X1 U4314 ( .A1(n3502), .A2(n3501), .ZN(n3503) );
  XNOR2_X1 U4315 ( .A(n3503), .B(n3277), .ZN(n3508) );
  INV_X1 U4316 ( .A(n3508), .ZN(n3506) );
  NOR2_X1 U4317 ( .A1(n3992), .A2(n3551), .ZN(n3504) );
  AOI21_X1 U4318 ( .B1(n4237), .B2(n3513), .A(n3504), .ZN(n3507) );
  INV_X1 U4319 ( .A(n3507), .ZN(n3505) );
  NAND2_X1 U4320 ( .A1(n3506), .A2(n3505), .ZN(n3667) );
  AND2_X1 U4321 ( .A1(n3508), .A2(n3507), .ZN(n3666) );
  NAND2_X1 U4322 ( .A1(n3844), .A2(n3479), .ZN(n3510) );
  NAND2_X1 U4323 ( .A1(n4236), .A2(n2932), .ZN(n3509) );
  NAND2_X1 U4324 ( .A1(n3510), .A2(n3509), .ZN(n3511) );
  XNOR2_X1 U4325 ( .A(n3511), .B(n3399), .ZN(n3556) );
  NOR2_X1 U4326 ( .A1(n3976), .A2(n3551), .ZN(n3512) );
  AOI21_X1 U4327 ( .B1(n3844), .B2(n3513), .A(n3512), .ZN(n3554) );
  XNOR2_X1 U4328 ( .A(n3556), .B(n3554), .ZN(n3547) );
  INV_X1 U4329 ( .A(n3514), .ZN(n3973) );
  INV_X1 U4330 ( .A(n4432), .ZN(n3675) );
  OAI22_X1 U4331 ( .A1(n4005), .A2(n4417), .B1(n4416), .B2(n3976), .ZN(n3517)
         );
  OAI22_X1 U4332 ( .A1(n4240), .A2(n3672), .B1(STATE_REG_SCAN_IN), .B2(n3515), 
        .ZN(n3516) );
  AOI211_X1 U4333 ( .C1(n3973), .C2(n3675), .A(n3517), .B(n3516), .ZN(n3518)
         );
  INV_X1 U4334 ( .A(n3519), .ZN(n3521) );
  NAND2_X1 U4335 ( .A1(n3521), .A2(n3520), .ZN(n3522) );
  XNOR2_X1 U4336 ( .A(n3523), .B(n3522), .ZN(n3527) );
  AND2_X1 U4337 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4543) );
  AOI21_X1 U4338 ( .B1(n4421), .B2(n4318), .A(n4543), .ZN(n3525) );
  AOI22_X1 U4339 ( .A1(n3682), .A2(n4316), .B1(n3681), .B2(n4215), .ZN(n3524)
         );
  OAI211_X1 U4340 ( .C1(n4432), .C2(n4217), .A(n3525), .B(n3524), .ZN(n3526)
         );
  AOI21_X1 U4341 ( .B1(n3527), .B2(n4427), .A(n3526), .ZN(n3528) );
  INV_X1 U4342 ( .A(n3528), .ZN(U3212) );
  INV_X1 U4343 ( .A(n3529), .ZN(n3646) );
  OAI21_X1 U4344 ( .B1(n3646), .B2(n3531), .A(n3530), .ZN(n3533) );
  NAND3_X1 U4345 ( .A1(n3533), .A2(n4427), .A3(n3532), .ZN(n3538) );
  AOI22_X1 U4346 ( .A1(n4007), .A2(n4421), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3537) );
  AOI22_X1 U4347 ( .A1(n3682), .A2(n3534), .B1(n3681), .B2(n4267), .ZN(n3536)
         );
  OR2_X1 U4348 ( .A1(n4432), .A2(n4048), .ZN(n3535) );
  NAND4_X1 U4349 ( .A1(n3538), .A2(n3537), .A3(n3536), .A4(n3535), .ZN(U3213)
         );
  XNOR2_X1 U4350 ( .A(n3540), .B(n3539), .ZN(n3545) );
  AND2_X1 U4351 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3938) );
  AOI21_X1 U4352 ( .B1(n3681), .B2(n4293), .A(n3938), .ZN(n3543) );
  AOI22_X1 U4353 ( .A1(n3682), .A2(n3541), .B1(n4421), .B2(n4079), .ZN(n3542)
         );
  OAI211_X1 U4354 ( .C1(n4432), .C2(n4121), .A(n3543), .B(n3542), .ZN(n3544)
         );
  AOI21_X1 U4355 ( .B1(n3545), .B2(n4427), .A(n3544), .ZN(n3546) );
  INV_X1 U4356 ( .A(n3546), .ZN(U3216) );
  OAI22_X1 U4357 ( .A1(n4240), .A2(n3548), .B1(n3551), .B2(n3559), .ZN(n3549)
         );
  XNOR2_X1 U4358 ( .A(n3549), .B(n3399), .ZN(n3553) );
  OAI22_X1 U4359 ( .A1(n4240), .A2(n3551), .B1(n3550), .B2(n3559), .ZN(n3552)
         );
  XNOR2_X1 U4360 ( .A(n3553), .B(n3552), .ZN(n3567) );
  INV_X1 U4361 ( .A(n3567), .ZN(n3557) );
  INV_X1 U4362 ( .A(n3554), .ZN(n3555) );
  NAND2_X1 U4363 ( .A1(n3556), .A2(n3555), .ZN(n3565) );
  OAI22_X1 U4364 ( .A1(n3986), .A2(n4417), .B1(n4416), .B2(n3559), .ZN(n3563)
         );
  INV_X1 U4365 ( .A(n3843), .ZN(n3561) );
  OAI22_X1 U4366 ( .A1(n3561), .A2(n3672), .B1(STATE_REG_SCAN_IN), .B2(n3560), 
        .ZN(n3562) );
  AOI211_X1 U4367 ( .C1(n3959), .C2(n3675), .A(n3563), .B(n3562), .ZN(n3570)
         );
  NAND3_X1 U4368 ( .A1(n3564), .A2(n4427), .A3(n3567), .ZN(n3569) );
  INV_X1 U4369 ( .A(n3565), .ZN(n3566) );
  NAND3_X1 U4370 ( .A1(n3567), .A2(n4427), .A3(n3566), .ZN(n3568) );
  NAND4_X1 U4371 ( .A1(n3571), .A2(n3570), .A3(n3569), .A4(n3568), .ZN(U3217)
         );
  XOR2_X1 U4372 ( .A(n3573), .B(n3572), .Z(n3574) );
  XNOR2_X1 U4373 ( .A(n3575), .B(n3574), .ZN(n3579) );
  AOI22_X1 U4374 ( .A1(n3681), .A2(n4079), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3577) );
  AOI22_X1 U4375 ( .A1(n3682), .A2(n4266), .B1(n4421), .B2(n4267), .ZN(n3576)
         );
  OAI211_X1 U4376 ( .C1(n4432), .C2(n4080), .A(n3577), .B(n3576), .ZN(n3578)
         );
  AOI21_X1 U4377 ( .B1(n3579), .B2(n4427), .A(n3578), .ZN(n3580) );
  INV_X1 U4378 ( .A(n3580), .ZN(U3220) );
  NAND2_X1 U4379 ( .A1(n3406), .A2(n3582), .ZN(n3583) );
  XNOR2_X1 U4380 ( .A(n3584), .B(n3583), .ZN(n3591) );
  NAND2_X1 U4381 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4519) );
  INV_X1 U4382 ( .A(n4519), .ZN(n3585) );
  AOI21_X1 U4383 ( .B1(n3681), .B2(n3845), .A(n3585), .ZN(n3588) );
  AOI22_X1 U4384 ( .A1(n3682), .A2(n3586), .B1(n4421), .B2(n4215), .ZN(n3587)
         );
  OAI211_X1 U4385 ( .C1(n4432), .C2(n3589), .A(n3588), .B(n3587), .ZN(n3590)
         );
  AOI21_X1 U4386 ( .B1(n3591), .B2(n4427), .A(n3590), .ZN(n3592) );
  INV_X1 U4387 ( .A(n3592), .ZN(U3221) );
  NAND2_X1 U4388 ( .A1(n2248), .A2(n3594), .ZN(n3595) );
  XNOR2_X1 U4389 ( .A(n3593), .B(n3595), .ZN(n3603) );
  INV_X1 U4390 ( .A(n4013), .ZN(n3601) );
  AOI22_X1 U4391 ( .A1(n4237), .A2(n4421), .B1(n3682), .B2(n3596), .ZN(n3600)
         );
  NOR2_X1 U4392 ( .A1(n3597), .A2(STATE_REG_SCAN_IN), .ZN(n3598) );
  AOI21_X1 U4393 ( .B1(n4007), .B2(n3681), .A(n3598), .ZN(n3599) );
  OAI211_X1 U4394 ( .C1(n4432), .C2(n3601), .A(n3600), .B(n3599), .ZN(n3602)
         );
  AOI21_X1 U4395 ( .B1(n3603), .B2(n4427), .A(n3602), .ZN(n3604) );
  INV_X1 U4396 ( .A(n3604), .ZN(U3222) );
  NAND2_X1 U4397 ( .A1(n3606), .A2(n3605), .ZN(n3608) );
  XOR2_X1 U4398 ( .A(n3608), .B(n3607), .Z(n3612) );
  NOR2_X1 U4399 ( .A1(STATE_REG_SCAN_IN), .A2(n2698), .ZN(n4572) );
  AOI21_X1 U4400 ( .B1(n3681), .B2(n4308), .A(n4572), .ZN(n3610) );
  AOI22_X1 U4401 ( .A1(n3682), .A2(n4292), .B1(n4421), .B2(n4293), .ZN(n3609)
         );
  OAI211_X1 U4402 ( .C1(n4432), .C2(n4154), .A(n3610), .B(n3609), .ZN(n3611)
         );
  AOI21_X1 U4403 ( .B1(n3612), .B2(n4427), .A(n3611), .ZN(n3613) );
  INV_X1 U4404 ( .A(n3613), .ZN(U3225) );
  NAND2_X1 U4405 ( .A1(n3615), .A2(n3614), .ZN(n3617) );
  XNOR2_X1 U4406 ( .A(n3617), .B(n3616), .ZN(n3621) );
  AOI22_X1 U4407 ( .A1(n3682), .A2(n4029), .B1(n4026), .B2(n4421), .ZN(n3619)
         );
  AOI22_X1 U4408 ( .A1(n3681), .A2(n4055), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3618) );
  OAI211_X1 U4409 ( .C1(n4432), .C2(n4032), .A(n3619), .B(n3618), .ZN(n3620)
         );
  AOI21_X1 U4410 ( .B1(n3621), .B2(n4427), .A(n3620), .ZN(n3622) );
  INV_X1 U4411 ( .A(n3622), .ZN(U3226) );
  INV_X1 U4412 ( .A(n3623), .ZN(n3628) );
  AOI21_X1 U4413 ( .B1(n3627), .B2(n3625), .A(n3624), .ZN(n3626) );
  AOI21_X1 U4414 ( .B1(n3628), .B2(n3627), .A(n3626), .ZN(n3634) );
  AOI22_X1 U4415 ( .A1(n3681), .A2(n4278), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3631) );
  AOI22_X1 U4416 ( .A1(n3682), .A2(n3629), .B1(n4421), .B2(n4096), .ZN(n3630)
         );
  OAI211_X1 U4417 ( .C1(n4432), .C2(n4097), .A(n3631), .B(n3630), .ZN(n3632)
         );
  INV_X1 U4418 ( .A(n3632), .ZN(n3633) );
  OAI21_X1 U4419 ( .B1(n3634), .B2(n3678), .A(n3633), .ZN(U3230) );
  XNOR2_X1 U4420 ( .A(n3637), .B(n3636), .ZN(n3638) );
  XNOR2_X1 U4421 ( .A(n3635), .B(n3638), .ZN(n3644) );
  NOR2_X1 U4422 ( .A1(STATE_REG_SCAN_IN), .A2(n5058), .ZN(n4533) );
  AOI21_X1 U4423 ( .B1(n3681), .B2(n4331), .A(n4533), .ZN(n3641) );
  AOI22_X1 U4424 ( .A1(n3682), .A2(n3639), .B1(n4421), .B2(n4193), .ZN(n3640)
         );
  OAI211_X1 U4425 ( .C1(n4432), .C2(n3642), .A(n3641), .B(n3640), .ZN(n3643)
         );
  AOI21_X1 U4426 ( .B1(n3644), .B2(n4427), .A(n3643), .ZN(n3645) );
  INV_X1 U4427 ( .A(n3645), .ZN(U3231) );
  AOI21_X1 U4428 ( .B1(n3648), .B2(n3647), .A(n3646), .ZN(n3654) );
  INV_X1 U4429 ( .A(n3649), .ZN(n4067) );
  OAI22_X1 U4430 ( .A1(n4276), .A2(n4417), .B1(STATE_REG_SCAN_IN), .B2(n3650), 
        .ZN(n3652) );
  OAI22_X1 U4431 ( .A1(n4024), .A2(n3672), .B1(n4416), .B2(n4064), .ZN(n3651)
         );
  AOI211_X1 U4432 ( .C1(n4067), .C2(n3675), .A(n3652), .B(n3651), .ZN(n3653)
         );
  OAI21_X1 U4433 ( .B1(n3654), .B2(n3678), .A(n3653), .ZN(U3232) );
  INV_X1 U4434 ( .A(n3655), .ZN(n3660) );
  AOI21_X1 U4435 ( .B1(n3657), .B2(n3659), .A(n3656), .ZN(n3658) );
  AOI21_X1 U4436 ( .B1(n3660), .B2(n3659), .A(n3658), .ZN(n3665) );
  AOI22_X1 U4437 ( .A1(n4421), .A2(n4278), .B1(REG3_REG_18__SCAN_IN), .B2(
        U3149), .ZN(n3662) );
  AOI22_X1 U4438 ( .A1(n3682), .A2(n4138), .B1(n3681), .B2(n4420), .ZN(n3661)
         );
  OAI211_X1 U4439 ( .C1(n4432), .C2(n4130), .A(n3662), .B(n3661), .ZN(n3663)
         );
  INV_X1 U4440 ( .A(n3663), .ZN(n3664) );
  OAI21_X1 U4441 ( .B1(n3665), .B2(n3678), .A(n3664), .ZN(U3235) );
  INV_X1 U4442 ( .A(n3666), .ZN(n3668) );
  NAND2_X1 U4443 ( .A1(n3668), .A2(n3667), .ZN(n3669) );
  XNOR2_X1 U4444 ( .A(n2223), .B(n3669), .ZN(n3679) );
  INV_X1 U4445 ( .A(n3995), .ZN(n3676) );
  OAI22_X1 U4446 ( .A1(n3671), .A2(n4417), .B1(STATE_REG_SCAN_IN), .B2(n3670), 
        .ZN(n3674) );
  OAI22_X1 U4447 ( .A1(n3986), .A2(n3672), .B1(n4416), .B2(n3992), .ZN(n3673)
         );
  AOI211_X1 U4448 ( .C1(n3676), .C2(n3675), .A(n3674), .B(n3673), .ZN(n3677)
         );
  OAI21_X1 U4449 ( .B1(n3679), .B2(n3678), .A(n3677), .ZN(U3237) );
  NAND2_X1 U4450 ( .A1(n4422), .A2(n4423), .ZN(n3680) );
  XNOR2_X1 U4451 ( .A(n3680), .B(n4424), .ZN(n3686) );
  AND2_X1 U4452 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4552) );
  AOI21_X1 U4453 ( .B1(n4421), .B2(n4308), .A(n4552), .ZN(n3684) );
  AOI22_X1 U4454 ( .A1(n3682), .A2(n4307), .B1(n3681), .B2(n4193), .ZN(n3683)
         );
  OAI211_X1 U4455 ( .C1(n4432), .C2(n4194), .A(n3684), .B(n3683), .ZN(n3685)
         );
  AOI21_X1 U4456 ( .B1(n3686), .B2(n4427), .A(n3685), .ZN(n3687) );
  INV_X1 U4457 ( .A(n3687), .ZN(U3238) );
  NAND3_X1 U4458 ( .A1(n2229), .A2(n4182), .A3(n3796), .ZN(n3690) );
  NAND2_X1 U4459 ( .A1(n3689), .A2(n3688), .ZN(n3784) );
  NAND2_X1 U4460 ( .A1(n3784), .A2(n3796), .ZN(n3787) );
  NAND2_X1 U4461 ( .A1(n3690), .A2(n3787), .ZN(n3692) );
  INV_X1 U4462 ( .A(n3803), .ZN(n3691) );
  AOI211_X1 U4463 ( .C1(n3692), .C2(n3806), .A(n3691), .B(n3805), .ZN(n3693)
         );
  OAI21_X1 U4464 ( .B1(n3693), .B2(n3810), .A(n3809), .ZN(n3694) );
  NAND2_X1 U4465 ( .A1(n3694), .A2(n3814), .ZN(n3696) );
  INV_X1 U4466 ( .A(n3695), .ZN(n3817) );
  AOI21_X1 U4467 ( .B1(n3697), .B2(n3696), .A(n3817), .ZN(n3699) );
  INV_X1 U4468 ( .A(n3815), .ZN(n3698) );
  OAI21_X1 U4469 ( .B1(n3699), .B2(n3698), .A(n3818), .ZN(n3700) );
  AND3_X1 U4470 ( .A1(n3700), .A2(n3969), .A3(n3822), .ZN(n3705) );
  NAND2_X1 U4471 ( .A1(n3702), .A2(n3701), .ZN(n3824) );
  NAND2_X1 U4472 ( .A1(n3843), .A2(n3956), .ZN(n3703) );
  AND2_X1 U4473 ( .A1(n3704), .A2(n3703), .ZN(n3825) );
  OAI21_X1 U4474 ( .B1(n3705), .B2(n3824), .A(n3825), .ZN(n3716) );
  INV_X1 U4475 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4341) );
  NAND2_X1 U4476 ( .A1(n3706), .A2(REG2_REG_31__SCAN_IN), .ZN(n3708) );
  NAND2_X1 U4477 ( .A1(n2538), .A2(REG1_REG_31__SCAN_IN), .ZN(n3707) );
  OAI211_X1 U4478 ( .C1(n2553), .C2(n4341), .A(n3708), .B(n3707), .ZN(n3841)
         );
  INV_X1 U4479 ( .A(n3841), .ZN(n3947) );
  OR2_X1 U4480 ( .A1(n3843), .A2(n3956), .ZN(n3711) );
  NAND2_X1 U4481 ( .A1(n3712), .A2(n4233), .ZN(n3710) );
  NAND2_X1 U4482 ( .A1(n3709), .A2(DATAI_31_), .ZN(n3945) );
  NAND2_X1 U4483 ( .A1(n3841), .A2(n3945), .ZN(n3827) );
  AND2_X1 U4484 ( .A1(n3710), .A2(n3827), .ZN(n3735) );
  NAND2_X1 U4485 ( .A1(n3711), .A2(n3735), .ZN(n3823) );
  AOI21_X1 U4486 ( .B1(n4233), .B2(n3947), .A(n3823), .ZN(n3715) );
  INV_X1 U4487 ( .A(n3945), .ZN(n3948) );
  INV_X1 U4488 ( .A(n3712), .ZN(n3842) );
  INV_X1 U4489 ( .A(n4233), .ZN(n3713) );
  NAND2_X1 U4490 ( .A1(n3842), .A2(n3713), .ZN(n3728) );
  NAND2_X1 U4491 ( .A1(n3728), .A2(n3841), .ZN(n3714) );
  AOI22_X1 U4492 ( .A1(n3716), .A2(n3715), .B1(n3948), .B2(n3714), .ZN(n3753)
         );
  NAND2_X1 U4493 ( .A1(n3717), .A2(n3822), .ZN(n3984) );
  NAND2_X1 U4494 ( .A1(n4038), .A2(n3808), .ZN(n4073) );
  NOR3_X1 U4495 ( .A1(n3718), .A2(n3984), .A3(n4073), .ZN(n3726) );
  NOR4_X1 U4496 ( .A1(n4597), .A2(n3721), .A3(n3720), .A4(n3719), .ZN(n3725)
         );
  NOR4_X1 U4497 ( .A1(n2794), .A2(n2464), .A3(n4060), .A4(n3722), .ZN(n3724)
         );
  NOR4_X1 U4498 ( .A1(n4620), .A2(n4660), .A3(n4208), .A4(n4190), .ZN(n3723)
         );
  NAND4_X1 U4499 ( .A1(n3726), .A2(n3725), .A3(n3724), .A4(n3723), .ZN(n3746)
         );
  OR2_X1 U4500 ( .A1(n3841), .A2(n3945), .ZN(n3727) );
  AND2_X1 U4501 ( .A1(n3728), .A2(n3727), .ZN(n3826) );
  OR2_X1 U4502 ( .A1(n2250), .A2(n3729), .ZN(n4041) );
  NAND2_X1 U4503 ( .A1(n3731), .A2(n3730), .ZN(n4093) );
  NAND2_X1 U4504 ( .A1(n4041), .A2(n4093), .ZN(n3733) );
  NAND2_X1 U4505 ( .A1(n3982), .A2(n3732), .ZN(n4004) );
  NOR2_X1 U4506 ( .A1(n3733), .A2(n4004), .ZN(n3734) );
  NAND4_X1 U4507 ( .A1(n3969), .A2(n3826), .A3(n3735), .A4(n3734), .ZN(n3745)
         );
  NAND2_X1 U4508 ( .A1(n3736), .A2(n4001), .ZN(n4021) );
  INV_X1 U4509 ( .A(n4021), .ZN(n3739) );
  INV_X1 U4510 ( .A(n4092), .ZN(n3737) );
  OR2_X1 U4511 ( .A1(n3737), .A2(n4091), .ZN(n4117) );
  NAND4_X1 U4512 ( .A1(n3739), .A2(n4149), .A3(n3738), .A4(n4117), .ZN(n3744)
         );
  NAND4_X1 U4513 ( .A1(n3742), .A2(n3741), .A3(n4136), .A4(n3740), .ZN(n3743)
         );
  OR4_X1 U4514 ( .A1(n3746), .A2(n3745), .A3(n3744), .A4(n3743), .ZN(n3750) );
  NOR4_X1 U4515 ( .A1(n3750), .A2(n3749), .A3(n3748), .A4(n3747), .ZN(n3752)
         );
  MUX2_X1 U4516 ( .A(n3753), .B(n3752), .S(n3751), .Z(n3833) );
  OAI211_X1 U4517 ( .C1(n2352), .C2(n3757), .A(n3756), .B(n3755), .ZN(n3760)
         );
  NAND3_X1 U4518 ( .A1(n3760), .A2(n3759), .A3(n3758), .ZN(n3762) );
  OAI211_X1 U4519 ( .C1(n3764), .C2(n3763), .A(n3762), .B(n3761), .ZN(n3767)
         );
  NAND3_X1 U4520 ( .A1(n3767), .A2(n3766), .A3(n3765), .ZN(n3770) );
  NAND4_X1 U4521 ( .A1(n3770), .A2(n3769), .A3(n3779), .A4(n3768), .ZN(n3773)
         );
  NAND3_X1 U4522 ( .A1(n3773), .A2(n3772), .A3(n3771), .ZN(n3774) );
  NAND3_X1 U4523 ( .A1(n3774), .A2(n3781), .A3(n3780), .ZN(n3777) );
  AND3_X1 U4524 ( .A1(n3777), .A2(n3776), .A3(n3775), .ZN(n3785) );
  INV_X1 U4525 ( .A(n3787), .ZN(n3800) );
  INV_X1 U4526 ( .A(n3778), .ZN(n3782) );
  NAND4_X1 U4527 ( .A1(n3782), .A2(n3781), .A3(n3780), .A4(n3779), .ZN(n3783)
         );
  OAI22_X1 U4528 ( .A1(n3785), .A2(n3784), .B1(n3800), .B2(n3783), .ZN(n3789)
         );
  AOI22_X1 U4529 ( .A1(n3789), .A2(n3788), .B1(n2349), .B2(n3787), .ZN(n3802)
         );
  NAND3_X1 U4530 ( .A1(n3793), .A2(n3791), .A3(n3790), .ZN(n3801) );
  INV_X1 U4531 ( .A(n3792), .ZN(n3795) );
  OAI21_X1 U4532 ( .B1(n3795), .B2(n3794), .A(n3793), .ZN(n3798) );
  AND4_X1 U4533 ( .A1(n3798), .A2(n4182), .A3(n3797), .A4(n3796), .ZN(n3799)
         );
  OAI22_X1 U4534 ( .A1(n3802), .A2(n3801), .B1(n3800), .B2(n3799), .ZN(n3804)
         );
  NAND2_X1 U4535 ( .A1(n3804), .A2(n3803), .ZN(n3807) );
  AOI21_X1 U4536 ( .B1(n3807), .B2(n3806), .A(n3805), .ZN(n3811) );
  OAI211_X1 U4537 ( .C1(n3811), .C2(n3810), .A(n3809), .B(n3808), .ZN(n3813)
         );
  AOI21_X1 U4538 ( .B1(n3814), .B2(n3813), .A(n3812), .ZN(n3816) );
  OAI21_X1 U4539 ( .B1(n3817), .B2(n3816), .A(n3815), .ZN(n3819) );
  NAND2_X1 U4540 ( .A1(n3819), .A2(n3818), .ZN(n3820) );
  NAND4_X1 U4541 ( .A1(n3825), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3830)
         );
  AOI21_X1 U4542 ( .B1(n3825), .B2(n3824), .A(n3823), .ZN(n3829) );
  INV_X1 U4543 ( .A(n3826), .ZN(n3828) );
  AOI22_X1 U4544 ( .A1(n3830), .A2(n3829), .B1(n3828), .B2(n3827), .ZN(n3832)
         );
  MUX2_X1 U4545 ( .A(n3833), .B(n3832), .S(n3831), .Z(n3834) );
  XNOR2_X1 U4546 ( .A(n3834), .B(n4143), .ZN(n3840) );
  NAND2_X1 U4547 ( .A1(n3836), .A2(n3835), .ZN(n3837) );
  OAI211_X1 U4548 ( .C1(n4406), .C2(n3839), .A(n3837), .B(B_REG_SCAN_IN), .ZN(
        n3838) );
  OAI21_X1 U4549 ( .B1(n3840), .B2(n3839), .A(n3838), .ZN(U3239) );
  MUX2_X1 U4550 ( .A(DATAO_REG_31__SCAN_IN), .B(n3841), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4551 ( .A(n3842), .B(DATAO_REG_30__SCAN_IN), .S(n3854), .Z(U3580)
         );
  MUX2_X1 U4552 ( .A(DATAO_REG_29__SCAN_IN), .B(n3843), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4553 ( .A(n3972), .B(DATAO_REG_28__SCAN_IN), .S(n3854), .Z(U3578)
         );
  MUX2_X1 U4554 ( .A(n3844), .B(DATAO_REG_27__SCAN_IN), .S(n3854), .Z(U3577)
         );
  MUX2_X1 U4555 ( .A(n4237), .B(DATAO_REG_26__SCAN_IN), .S(n3854), .Z(U3576)
         );
  MUX2_X1 U4556 ( .A(n4026), .B(DATAO_REG_25__SCAN_IN), .S(n3854), .Z(U3575)
         );
  MUX2_X1 U4557 ( .A(n4007), .B(DATAO_REG_24__SCAN_IN), .S(n3854), .Z(U3574)
         );
  MUX2_X1 U4558 ( .A(n4055), .B(DATAO_REG_23__SCAN_IN), .S(n3854), .Z(U3573)
         );
  MUX2_X1 U4559 ( .A(n4267), .B(DATAO_REG_22__SCAN_IN), .S(n3854), .Z(U3572)
         );
  MUX2_X1 U4560 ( .A(n4096), .B(DATAO_REG_21__SCAN_IN), .S(n3854), .Z(U3571)
         );
  MUX2_X1 U4561 ( .A(n4079), .B(DATAO_REG_20__SCAN_IN), .S(n3854), .Z(U3570)
         );
  MUX2_X1 U4562 ( .A(n4278), .B(DATAO_REG_19__SCAN_IN), .S(n3854), .Z(U3569)
         );
  MUX2_X1 U4563 ( .A(n4293), .B(DATAO_REG_18__SCAN_IN), .S(n3854), .Z(U3568)
         );
  MUX2_X1 U4564 ( .A(n4420), .B(DATAO_REG_17__SCAN_IN), .S(n3854), .Z(U3567)
         );
  MUX2_X1 U4565 ( .A(n4308), .B(DATAO_REG_16__SCAN_IN), .S(n3854), .Z(U3566)
         );
  MUX2_X1 U4566 ( .A(n4318), .B(DATAO_REG_15__SCAN_IN), .S(n3854), .Z(U3565)
         );
  MUX2_X1 U4567 ( .A(n4193), .B(DATAO_REG_14__SCAN_IN), .S(n3854), .Z(U3564)
         );
  MUX2_X1 U4568 ( .A(n4215), .B(DATAO_REG_13__SCAN_IN), .S(n3854), .Z(U3563)
         );
  MUX2_X1 U4569 ( .A(n4331), .B(DATAO_REG_12__SCAN_IN), .S(n3854), .Z(U3562)
         );
  MUX2_X1 U4570 ( .A(n3845), .B(DATAO_REG_11__SCAN_IN), .S(n3854), .Z(U3561)
         );
  MUX2_X1 U4571 ( .A(n4593), .B(DATAO_REG_10__SCAN_IN), .S(n3854), .Z(U3560)
         );
  MUX2_X1 U4572 ( .A(n3846), .B(DATAO_REG_9__SCAN_IN), .S(n3854), .Z(U3559) );
  MUX2_X1 U4573 ( .A(n3847), .B(DATAO_REG_8__SCAN_IN), .S(n3854), .Z(U3558) );
  MUX2_X1 U4574 ( .A(n3848), .B(DATAO_REG_7__SCAN_IN), .S(n3854), .Z(U3557) );
  MUX2_X1 U4575 ( .A(n3849), .B(DATAO_REG_6__SCAN_IN), .S(n3854), .Z(U3556) );
  MUX2_X1 U4576 ( .A(n3850), .B(DATAO_REG_5__SCAN_IN), .S(n3854), .Z(U3555) );
  MUX2_X1 U4577 ( .A(n3851), .B(DATAO_REG_4__SCAN_IN), .S(n3854), .Z(U3554) );
  MUX2_X1 U4578 ( .A(n3852), .B(DATAO_REG_3__SCAN_IN), .S(n3854), .Z(U3553) );
  MUX2_X1 U4579 ( .A(n3853), .B(DATAO_REG_2__SCAN_IN), .S(n3854), .Z(U3552) );
  MUX2_X1 U4580 ( .A(n2979), .B(DATAO_REG_1__SCAN_IN), .S(n3854), .Z(U3551) );
  MUX2_X1 U4581 ( .A(DATAO_REG_0__SCAN_IN), .B(n4614), .S(U4043), .Z(U3550) );
  INV_X1 U4582 ( .A(n4590), .ZN(n3855) );
  NAND2_X1 U4583 ( .A1(n3855), .A2(n4411), .ZN(n3865) );
  OAI211_X1 U4584 ( .C1(n3858), .C2(n3857), .A(n4585), .B(n3856), .ZN(n3864)
         );
  MUX2_X1 U4585 ( .A(n2915), .B(REG2_REG_1__SCAN_IN), .S(n3859), .Z(n3860) );
  OAI211_X1 U4586 ( .C1(n3861), .C2(n3860), .A(n4528), .B(n2382), .ZN(n3863)
         );
  AOI22_X1 U4587 ( .A1(n4583), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3862) );
  NAND4_X1 U4588 ( .A1(n3865), .A2(n3864), .A3(n3863), .A4(n3862), .ZN(U3241)
         );
  AOI22_X1 U4589 ( .A1(n4583), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3866) );
  OAI21_X1 U4590 ( .B1(n4590), .B2(n3867), .A(n3866), .ZN(n3868) );
  INV_X1 U4591 ( .A(n3868), .ZN(n3879) );
  MUX2_X1 U4592 ( .A(n3869), .B(REG2_REG_2__SCAN_IN), .S(n4410), .Z(n3870) );
  NAND2_X1 U4593 ( .A1(n3870), .A2(n2262), .ZN(n3872) );
  OAI211_X1 U4594 ( .C1(n3873), .C2(n3872), .A(n4528), .B(n3871), .ZN(n3878)
         );
  OAI211_X1 U4595 ( .C1(n3876), .C2(n3875), .A(n4585), .B(n3874), .ZN(n3877)
         );
  NAND4_X1 U4596 ( .A1(n3880), .A2(n3879), .A3(n3878), .A4(n3877), .ZN(U3242)
         );
  MUX2_X1 U4597 ( .A(n4122), .B(REG2_REG_19__SCAN_IN), .S(n3940), .Z(n3905) );
  INV_X1 U4598 ( .A(n3906), .ZN(n4644) );
  INV_X1 U4599 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4600 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4644), .B1(n3906), .B2(
        n3881), .ZN(n4581) );
  NOR2_X1 U4601 ( .A1(n3933), .A2(REG2_REG_17__SCAN_IN), .ZN(n3882) );
  AOI21_X1 U4602 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3933), .A(n3882), .ZN(n4570) );
  INV_X1 U4603 ( .A(n3926), .ZN(n4650) );
  INV_X1 U4604 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4527) );
  INV_X1 U4605 ( .A(n3907), .ZN(n4651) );
  NOR2_X1 U4606 ( .A1(n4527), .A2(n4651), .ZN(n4526) );
  NAND2_X1 U4607 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3908), .ZN(n3896) );
  AOI22_X1 U4608 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3908), .B1(n4653), .B2(
        n2637), .ZN(n4510) );
  NAND2_X1 U4609 ( .A1(n3909), .A2(REG2_REG_9__SCAN_IN), .ZN(n3893) );
  INV_X1 U4610 ( .A(n3909), .ZN(n4654) );
  AOI22_X1 U4611 ( .A1(n3909), .A2(REG2_REG_9__SCAN_IN), .B1(n2609), .B2(n4654), .ZN(n4489) );
  NAND2_X1 U4612 ( .A1(n3917), .A2(REG2_REG_7__SCAN_IN), .ZN(n3890) );
  INV_X1 U4613 ( .A(n3917), .ZN(n4655) );
  AOI22_X1 U4614 ( .A1(n3917), .A2(REG2_REG_7__SCAN_IN), .B1(n2590), .B2(n4655), .ZN(n4471) );
  NAND2_X1 U4615 ( .A1(n3913), .A2(REG2_REG_5__SCAN_IN), .ZN(n3887) );
  INV_X1 U4616 ( .A(n3913), .ZN(n4657) );
  AOI22_X1 U4617 ( .A1(n3913), .A2(REG2_REG_5__SCAN_IN), .B1(n2567), .B2(n4657), .ZN(n4450) );
  NAND2_X1 U4618 ( .A1(n3883), .A2(REG2_REG_4__SCAN_IN), .ZN(n3884) );
  NAND2_X1 U4619 ( .A1(n3914), .A2(n3888), .ZN(n3889) );
  NAND2_X1 U4620 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4460), .ZN(n4459) );
  NAND2_X1 U4621 ( .A1(n4474), .A2(n3891), .ZN(n3892) );
  NAND2_X1 U4622 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4476), .ZN(n4475) );
  NAND2_X1 U4623 ( .A1(n4495), .A2(n3894), .ZN(n3895) );
  NAND2_X1 U4624 ( .A1(n4516), .A2(n3897), .ZN(n3898) );
  NOR2_X1 U4625 ( .A1(n4650), .A2(n3899), .ZN(n3900) );
  INV_X1 U4626 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4541) );
  XNOR2_X1 U4627 ( .A(n4650), .B(n3899), .ZN(n4540) );
  NOR2_X1 U4628 ( .A1(n4541), .A2(n4540), .ZN(n4539) );
  NOR2_X1 U4629 ( .A1(n3900), .A2(n4539), .ZN(n4550) );
  NAND2_X1 U4630 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4648), .ZN(n3901) );
  OAI21_X1 U4631 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4648), .A(n3901), .ZN(n4549) );
  NOR2_X1 U4632 ( .A1(n4550), .A2(n4549), .ZN(n4548) );
  AOI21_X1 U4633 ( .B1(n4648), .B2(REG2_REG_15__SCAN_IN), .A(n4548), .ZN(n3902) );
  INV_X1 U4634 ( .A(n3930), .ZN(n4647) );
  NAND2_X1 U4635 ( .A1(n3902), .A2(n4647), .ZN(n3903) );
  XOR2_X1 U4636 ( .A(n3902), .B(n4647), .Z(n4561) );
  INV_X1 U4637 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4559) );
  NAND2_X1 U4638 ( .A1(n4561), .A2(n4559), .ZN(n4560) );
  AOI21_X1 U4639 ( .B1(REG2_REG_18__SCAN_IN), .B2(n3906), .A(n4580), .ZN(n3904) );
  XOR2_X1 U4640 ( .A(n3905), .B(n3904), .Z(n3944) );
  AOI22_X1 U4641 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3906), .B1(n4644), .B2(
        n3935), .ZN(n4587) );
  NOR2_X1 U4642 ( .A1(n3933), .A2(REG1_REG_17__SCAN_IN), .ZN(n3934) );
  NAND2_X1 U4643 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4648), .ZN(n3929) );
  INV_X1 U4644 ( .A(n4648), .ZN(n4558) );
  AOI22_X1 U4645 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4648), .B1(n4558), .B2(
        n4313), .ZN(n4555) );
  NAND2_X1 U4646 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3907), .ZN(n3925) );
  AOI22_X1 U4647 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3907), .B1(n4651), .B2(
        n4337), .ZN(n4536) );
  AOI22_X1 U4648 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3908), .B1(n4653), .B2(
        n4715), .ZN(n4507) );
  NAND2_X1 U4649 ( .A1(n3909), .A2(REG1_REG_9__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4650 ( .A1(n3909), .A2(REG1_REG_9__SCAN_IN), .B1(n3294), .B2(n4654), .ZN(n4486) );
  NAND2_X1 U4651 ( .A1(n3913), .A2(REG1_REG_5__SCAN_IN), .ZN(n3912) );
  OAI21_X1 U4652 ( .B1(n3913), .B2(REG1_REG_5__SCAN_IN), .A(n3912), .ZN(n4444)
         );
  INV_X1 U4653 ( .A(n3914), .ZN(n4656) );
  NOR2_X1 U4654 ( .A1(n3915), .A2(n4656), .ZN(n3916) );
  XNOR2_X1 U4655 ( .A(n3915), .B(n4656), .ZN(n4455) );
  NOR2_X1 U4656 ( .A1(n4456), .A2(n4455), .ZN(n4454) );
  NAND2_X1 U4657 ( .A1(n3917), .A2(REG1_REG_7__SCAN_IN), .ZN(n4463) );
  NAND2_X1 U4658 ( .A1(n4474), .A2(n3918), .ZN(n3919) );
  NAND2_X1 U4659 ( .A1(n3919), .A2(n4480), .ZN(n4485) );
  NAND2_X1 U4660 ( .A1(n4495), .A2(n3921), .ZN(n3922) );
  NAND2_X1 U4661 ( .A1(n3922), .A2(n4501), .ZN(n4506) );
  NAND2_X1 U4662 ( .A1(n4516), .A2(n3923), .ZN(n3924) );
  NAND2_X1 U4663 ( .A1(n3924), .A2(n4522), .ZN(n4535) );
  NAND2_X1 U4664 ( .A1(n3926), .A2(n3927), .ZN(n3928) );
  NAND2_X1 U4665 ( .A1(n3928), .A2(n4544), .ZN(n4554) );
  NOR2_X1 U4666 ( .A1(n3930), .A2(n3931), .ZN(n3932) );
  NOR2_X1 U4667 ( .A1(n3932), .A2(n4565), .ZN(n4574) );
  INV_X1 U4668 ( .A(n3933), .ZN(n4645) );
  AOI22_X1 U4669 ( .A1(n3933), .A2(n4299), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4645), .ZN(n4573) );
  NOR2_X1 U4670 ( .A1(n4574), .A2(n4573), .ZN(n4575) );
  NOR2_X1 U4671 ( .A1(n3934), .A2(n4575), .ZN(n4586) );
  NAND2_X1 U4672 ( .A1(n4587), .A2(n4586), .ZN(n4584) );
  OAI21_X1 U4673 ( .B1(n4644), .B2(n3935), .A(n4584), .ZN(n3937) );
  MUX2_X1 U4674 ( .A(REG1_REG_19__SCAN_IN), .B(n4287), .S(n3940), .Z(n3936) );
  XNOR2_X1 U4675 ( .A(n3937), .B(n3936), .ZN(n3942) );
  AOI21_X1 U4676 ( .B1(n4583), .B2(ADDR_REG_19__SCAN_IN), .A(n3938), .ZN(n3939) );
  OAI21_X1 U4677 ( .B1(n4590), .B2(n3940), .A(n3939), .ZN(n3941) );
  AOI21_X1 U4678 ( .B1(n3942), .B2(n4585), .A(n3941), .ZN(n3943) );
  OAI21_X1 U4679 ( .B1(n3944), .B2(n4579), .A(n3943), .ZN(U3259) );
  NOR2_X1 U4680 ( .A1(n4231), .A2(n4233), .ZN(n4230) );
  XNOR2_X1 U4681 ( .A(n4230), .B(n3945), .ZN(n4343) );
  NOR2_X1 U4682 ( .A1(n3947), .A2(n3946), .ZN(n4232) );
  AOI21_X1 U4683 ( .B1(n3948), .B2(n4611), .A(n4232), .ZN(n4340) );
  NOR2_X1 U4684 ( .A1(n4340), .A2(n4626), .ZN(n3949) );
  AOI21_X1 U4685 ( .B1(REG2_REG_31__SCAN_IN), .B2(n4626), .A(n3949), .ZN(n3950) );
  OAI21_X1 U4686 ( .B1(n4343), .B2(n4160), .A(n3950), .ZN(U3260) );
  OAI22_X1 U4687 ( .A1(n3952), .A2(n4160), .B1(n3951), .B2(n4171), .ZN(n3953)
         );
  AOI22_X1 U4688 ( .A1(n3972), .A2(n4216), .B1(n4626), .B2(
        REG2_REG_29__SCAN_IN), .ZN(n3955) );
  INV_X1 U4689 ( .A(n3958), .ZN(n3965) );
  AOI22_X1 U4690 ( .A1(n3959), .A2(n4627), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4626), .ZN(n3960) );
  OAI21_X1 U4691 ( .B1(n3961), .B2(n4160), .A(n3960), .ZN(n3962) );
  AOI21_X1 U4692 ( .B1(n3963), .B2(n4172), .A(n3962), .ZN(n3964) );
  OAI21_X1 U4693 ( .B1(n3965), .B2(n4177), .A(n3964), .ZN(U3262) );
  NOR2_X1 U4694 ( .A1(n2242), .A2(n3969), .ZN(n3966) );
  OR2_X1 U4695 ( .A1(n3967), .A2(n3966), .ZN(n3968) );
  NAND2_X1 U4696 ( .A1(n3968), .A2(n4625), .ZN(n4239) );
  XNOR2_X1 U4697 ( .A(n2240), .B(n3969), .ZN(n4242) );
  NAND2_X1 U4698 ( .A1(n4242), .A2(n4191), .ZN(n3980) );
  INV_X1 U4699 ( .A(n3970), .ZN(n3971) );
  OAI21_X1 U4700 ( .B1(n3990), .B2(n3976), .A(n3971), .ZN(n4349) );
  INV_X1 U4701 ( .A(n4349), .ZN(n3978) );
  AOI22_X1 U4702 ( .A1(n3972), .A2(n4214), .B1(n4216), .B2(n4237), .ZN(n3975)
         );
  AOI22_X1 U4703 ( .A1(n3973), .A2(n4627), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4626), .ZN(n3974) );
  OAI211_X1 U4704 ( .C1(n3976), .C2(n4221), .A(n3975), .B(n3974), .ZN(n3977)
         );
  AOI21_X1 U4705 ( .B1(n3978), .B2(n4632), .A(n3977), .ZN(n3979) );
  OAI211_X1 U4706 ( .C1(n4626), .C2(n4239), .A(n3980), .B(n3979), .ZN(U3263)
         );
  XNOR2_X1 U4707 ( .A(n3981), .B(n3984), .ZN(n4246) );
  INV_X1 U4708 ( .A(n4246), .ZN(n3999) );
  NAND2_X1 U4709 ( .A1(n3983), .A2(n3982), .ZN(n3985) );
  XNOR2_X1 U4710 ( .A(n3985), .B(n3984), .ZN(n3989) );
  OAI22_X1 U4711 ( .A1(n3986), .A2(n4616), .B1(n4328), .B2(n3992), .ZN(n3987)
         );
  AOI21_X1 U4712 ( .B1(n4613), .B2(n4026), .A(n3987), .ZN(n3988) );
  OAI21_X1 U4713 ( .B1(n3989), .B2(n4333), .A(n3988), .ZN(n4245) );
  INV_X1 U4714 ( .A(n4010), .ZN(n3993) );
  INV_X1 U4715 ( .A(n3990), .ZN(n3991) );
  OAI21_X1 U4716 ( .B1(n3993), .B2(n3992), .A(n3991), .ZN(n4353) );
  NOR2_X1 U4717 ( .A1(n4353), .A2(n4160), .ZN(n3997) );
  OAI22_X1 U4718 ( .A1(n3995), .A2(n4171), .B1(n4172), .B2(n3994), .ZN(n3996)
         );
  AOI211_X1 U4719 ( .C1(n4245), .C2(n4172), .A(n3997), .B(n3996), .ZN(n3998)
         );
  OAI21_X1 U4720 ( .B1(n3999), .B2(n4177), .A(n3998), .ZN(U3264) );
  XNOR2_X1 U4721 ( .A(n4000), .B(n4004), .ZN(n4250) );
  INV_X1 U4722 ( .A(n4250), .ZN(n4017) );
  NAND2_X1 U4723 ( .A1(n4002), .A2(n4001), .ZN(n4003) );
  XOR2_X1 U4724 ( .A(n4004), .B(n4003), .Z(n4009) );
  OAI22_X1 U4725 ( .A1(n4005), .A2(n4616), .B1(n4328), .B2(n4011), .ZN(n4006)
         );
  AOI21_X1 U4726 ( .B1(n4613), .B2(n4007), .A(n4006), .ZN(n4008) );
  OAI21_X1 U4727 ( .B1(n4009), .B2(n4333), .A(n4008), .ZN(n4249) );
  INV_X1 U4728 ( .A(n4031), .ZN(n4012) );
  OAI21_X1 U4729 ( .B1(n4012), .B2(n4011), .A(n4010), .ZN(n4357) );
  AOI22_X1 U4730 ( .A1(n4626), .A2(REG2_REG_25__SCAN_IN), .B1(n4013), .B2(
        n4627), .ZN(n4014) );
  OAI21_X1 U4731 ( .B1(n4357), .B2(n4160), .A(n4014), .ZN(n4015) );
  AOI21_X1 U4732 ( .B1(n4249), .B2(n4172), .A(n4015), .ZN(n4016) );
  OAI21_X1 U4733 ( .B1(n4017), .B2(n4177), .A(n4016), .ZN(U3265) );
  XOR2_X1 U4734 ( .A(n4021), .B(n4018), .Z(n4254) );
  INV_X1 U4735 ( .A(n4254), .ZN(n4037) );
  NAND2_X1 U4736 ( .A1(n4020), .A2(n4019), .ZN(n4022) );
  XNOR2_X1 U4737 ( .A(n4022), .B(n4021), .ZN(n4028) );
  OAI22_X1 U4738 ( .A1(n4024), .A2(n4320), .B1(n4328), .B2(n4023), .ZN(n4025)
         );
  AOI21_X1 U4739 ( .B1(n4317), .B2(n4026), .A(n4025), .ZN(n4027) );
  OAI21_X1 U4740 ( .B1(n4028), .B2(n4333), .A(n4027), .ZN(n4253) );
  NAND2_X1 U4741 ( .A1(n4046), .A2(n4029), .ZN(n4030) );
  NAND2_X1 U4742 ( .A1(n4031), .A2(n4030), .ZN(n4361) );
  NOR2_X1 U4743 ( .A1(n4361), .A2(n4160), .ZN(n4035) );
  OAI22_X1 U4744 ( .A1(n4172), .A2(n4033), .B1(n4032), .B2(n4171), .ZN(n4034)
         );
  AOI211_X1 U4745 ( .C1(n4253), .C2(n4172), .A(n4035), .B(n4034), .ZN(n4036)
         );
  OAI21_X1 U4746 ( .B1(n4037), .B2(n4177), .A(n4036), .ZN(U3266) );
  XOR2_X1 U4747 ( .A(n4041), .B(n2239), .Z(n4258) );
  INV_X1 U4748 ( .A(n4258), .ZN(n4053) );
  OR2_X1 U4749 ( .A1(n4074), .A2(n4073), .ZN(n4076) );
  AND2_X1 U4750 ( .A1(n4076), .A2(n4038), .ZN(n4054) );
  OAI21_X1 U4751 ( .B1(n4054), .B2(n4060), .A(n4039), .ZN(n4040) );
  XOR2_X1 U4752 ( .A(n4041), .B(n4040), .Z(n4045) );
  OAI22_X1 U4753 ( .A1(n4042), .A2(n4616), .B1(n4047), .B2(n4328), .ZN(n4043)
         );
  AOI21_X1 U4754 ( .B1(n4613), .B2(n4267), .A(n4043), .ZN(n4044) );
  OAI21_X1 U4755 ( .B1(n4045), .B2(n4333), .A(n4044), .ZN(n4257) );
  OAI21_X1 U4756 ( .B1(n4066), .B2(n4047), .A(n4046), .ZN(n4365) );
  NOR2_X1 U4757 ( .A1(n4365), .A2(n4160), .ZN(n4051) );
  INV_X1 U4758 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4049) );
  OAI22_X1 U4759 ( .A1(n4172), .A2(n4049), .B1(n4048), .B2(n4171), .ZN(n4050)
         );
  AOI211_X1 U4760 ( .C1(n4257), .C2(n4172), .A(n4051), .B(n4050), .ZN(n4052)
         );
  OAI21_X1 U4761 ( .B1(n4053), .B2(n4177), .A(n4052), .ZN(U3267) );
  XNOR2_X1 U4762 ( .A(n4054), .B(n4060), .ZN(n4059) );
  NAND2_X1 U4763 ( .A1(n4096), .A2(n4613), .ZN(n4057) );
  NAND2_X1 U4764 ( .A1(n4055), .A2(n4317), .ZN(n4056) );
  OAI211_X1 U4765 ( .C1(n4328), .C2(n4064), .A(n4057), .B(n4056), .ZN(n4058)
         );
  AOI21_X1 U4766 ( .B1(n4059), .B2(n4625), .A(n4058), .ZN(n4262) );
  NOR2_X1 U4767 ( .A1(n4061), .A2(n4060), .ZN(n4062) );
  OR2_X1 U4768 ( .A1(n4063), .A2(n4062), .ZN(n4261) );
  INV_X1 U4769 ( .A(n4261), .ZN(n4070) );
  NOR2_X1 U4770 ( .A1(n4077), .A2(n4064), .ZN(n4065) );
  AOI22_X1 U4771 ( .A1(n4626), .A2(REG2_REG_22__SCAN_IN), .B1(n4067), .B2(
        n4627), .ZN(n4068) );
  OAI21_X1 U4772 ( .B1(n4369), .B2(n4160), .A(n4068), .ZN(n4069) );
  AOI21_X1 U4773 ( .B1(n4070), .B2(n4191), .A(n4069), .ZN(n4071) );
  OAI21_X1 U4774 ( .B1(n4626), .B2(n4262), .A(n4071), .ZN(U3268) );
  XNOR2_X1 U4775 ( .A(n4072), .B(n4073), .ZN(n4272) );
  INV_X1 U4776 ( .A(n4272), .ZN(n4088) );
  NAND2_X1 U4777 ( .A1(n4074), .A2(n4073), .ZN(n4075) );
  AOI21_X1 U4778 ( .B1(n4076), .B2(n4075), .A(n4333), .ZN(n4271) );
  INV_X1 U4779 ( .A(n4077), .ZN(n4078) );
  OAI21_X1 U4780 ( .B1(n2407), .B2(n4084), .A(n4078), .ZN(n4373) );
  NOR2_X1 U4781 ( .A1(n4373), .A2(n4160), .ZN(n4086) );
  AOI22_X1 U4782 ( .A1(n4216), .A2(n4079), .B1(n4214), .B2(n4267), .ZN(n4083)
         );
  INV_X1 U4783 ( .A(n4080), .ZN(n4081) );
  AOI22_X1 U4784 ( .A1(n4626), .A2(REG2_REG_21__SCAN_IN), .B1(n4081), .B2(
        n4627), .ZN(n4082) );
  OAI211_X1 U4785 ( .C1(n4084), .C2(n4221), .A(n4083), .B(n4082), .ZN(n4085)
         );
  AOI211_X1 U4786 ( .C1(n4271), .C2(n4172), .A(n4086), .B(n4085), .ZN(n4087)
         );
  OAI21_X1 U4787 ( .B1(n4088), .B2(n4177), .A(n4087), .ZN(U3269) );
  NOR2_X1 U4788 ( .A1(n2252), .A2(n4089), .ZN(n4090) );
  XNOR2_X1 U4789 ( .A(n4090), .B(n4093), .ZN(n4280) );
  AOI21_X1 U4790 ( .B1(n4116), .B2(n4092), .A(n4091), .ZN(n4094) );
  XNOR2_X1 U4791 ( .A(n4094), .B(n4093), .ZN(n4282) );
  NAND2_X1 U4792 ( .A1(n4282), .A2(n4191), .ZN(n4104) );
  OAI21_X1 U4793 ( .B1(n2402), .B2(n4275), .A(n4095), .ZN(n4377) );
  INV_X1 U4794 ( .A(n4377), .ZN(n4102) );
  AOI22_X1 U4795 ( .A1(n4216), .A2(n4278), .B1(n4214), .B2(n4096), .ZN(n4100)
         );
  INV_X1 U4796 ( .A(n4097), .ZN(n4098) );
  AOI22_X1 U4797 ( .A1(n4626), .A2(REG2_REG_20__SCAN_IN), .B1(n4098), .B2(
        n4627), .ZN(n4099) );
  OAI211_X1 U4798 ( .C1(n4275), .C2(n4221), .A(n4100), .B(n4099), .ZN(n4101)
         );
  AOI21_X1 U4799 ( .B1(n4102), .B2(n4632), .A(n4101), .ZN(n4103) );
  OAI211_X1 U4800 ( .C1(n4280), .C2(n4105), .A(n4104), .B(n4103), .ZN(U3270)
         );
  INV_X1 U4801 ( .A(n4106), .ZN(n4108) );
  OAI21_X1 U4802 ( .B1(n4147), .B2(n4108), .A(n4107), .ZN(n4137) );
  INV_X1 U4803 ( .A(n4109), .ZN(n4111) );
  OAI21_X1 U4804 ( .B1(n4137), .B2(n4111), .A(n4110), .ZN(n4112) );
  XNOR2_X1 U4805 ( .A(n4112), .B(n4117), .ZN(n4115) );
  OAI22_X1 U4806 ( .A1(n4269), .A2(n4616), .B1(n4328), .B2(n4118), .ZN(n4113)
         );
  AOI21_X1 U4807 ( .B1(n4613), .B2(n4293), .A(n4113), .ZN(n4114) );
  OAI21_X1 U4808 ( .B1(n4115), .B2(n4333), .A(n4114), .ZN(n4285) );
  INV_X1 U4809 ( .A(n4285), .ZN(n4126) );
  XOR2_X1 U4810 ( .A(n4117), .B(n4116), .Z(n4286) );
  OR2_X1 U4811 ( .A1(n4132), .A2(n4118), .ZN(n4119) );
  NAND2_X1 U4812 ( .A1(n4120), .A2(n4119), .ZN(n4381) );
  NOR2_X1 U4813 ( .A1(n4381), .A2(n4160), .ZN(n4124) );
  OAI22_X1 U4814 ( .A1(n4172), .A2(n4122), .B1(n4121), .B2(n4171), .ZN(n4123)
         );
  AOI211_X1 U4815 ( .C1(n4286), .C2(n4191), .A(n4124), .B(n4123), .ZN(n4125)
         );
  OAI21_X1 U4816 ( .B1(n4626), .B2(n4126), .A(n4125), .ZN(U3271) );
  INV_X1 U4817 ( .A(n4127), .ZN(n4128) );
  AOI21_X1 U4818 ( .B1(n4136), .B2(n4129), .A(n4128), .ZN(n4291) );
  INV_X1 U4819 ( .A(n4130), .ZN(n4131) );
  AOI22_X1 U4820 ( .A1(n4626), .A2(REG2_REG_18__SCAN_IN), .B1(n4131), .B2(
        n4627), .ZN(n4146) );
  INV_X1 U4821 ( .A(n4132), .ZN(n4134) );
  OAI211_X1 U4822 ( .C1(n4151), .C2(n4135), .A(n4134), .B(n4133), .ZN(n4289)
         );
  XNOR2_X1 U4823 ( .A(n4137), .B(n4136), .ZN(n4142) );
  AOI22_X1 U4824 ( .A1(n4278), .A2(n4317), .B1(n4138), .B2(n4611), .ZN(n4139)
         );
  OAI21_X1 U4825 ( .B1(n4140), .B2(n4320), .A(n4139), .ZN(n4141) );
  AOI21_X1 U4826 ( .B1(n4142), .B2(n4625), .A(n4141), .ZN(n4290) );
  OAI21_X1 U4827 ( .B1(n4143), .B2(n4289), .A(n4290), .ZN(n4144) );
  NAND2_X1 U4828 ( .A1(n4144), .A2(n4172), .ZN(n4145) );
  OAI211_X1 U4829 ( .C1(n4291), .C2(n4177), .A(n4146), .B(n4145), .ZN(U3272)
         );
  XOR2_X1 U4830 ( .A(n4149), .B(n4147), .Z(n4148) );
  NAND2_X1 U4831 ( .A1(n4148), .A2(n4625), .ZN(n4295) );
  XNOR2_X1 U4832 ( .A(n4150), .B(n4149), .ZN(n4298) );
  INV_X1 U4833 ( .A(n4151), .ZN(n4153) );
  NAND2_X1 U4834 ( .A1(n4170), .A2(n4292), .ZN(n4152) );
  NAND2_X1 U4835 ( .A1(n4153), .A2(n4152), .ZN(n4386) );
  OAI22_X1 U4836 ( .A1(n4172), .A2(n4155), .B1(n4154), .B2(n4171), .ZN(n4156)
         );
  AOI21_X1 U4837 ( .B1(n4292), .B2(n4157), .A(n4156), .ZN(n4159) );
  AOI22_X1 U4838 ( .A1(n4216), .A2(n4308), .B1(n4214), .B2(n4293), .ZN(n4158)
         );
  OAI211_X1 U4839 ( .C1(n4386), .C2(n4160), .A(n4159), .B(n4158), .ZN(n4161)
         );
  AOI21_X1 U4840 ( .B1(n4298), .B2(n4191), .A(n4161), .ZN(n4162) );
  OAI21_X1 U4841 ( .B1(n4626), .B2(n4295), .A(n4162), .ZN(U3273) );
  XNOR2_X1 U4842 ( .A(n4163), .B(n2464), .ZN(n4167) );
  NAND2_X1 U4843 ( .A1(n4318), .A2(n4613), .ZN(n4165) );
  NAND2_X1 U4844 ( .A1(n4420), .A2(n4317), .ZN(n4164) );
  OAI211_X1 U4845 ( .C1(n4328), .C2(n4415), .A(n4165), .B(n4164), .ZN(n4166)
         );
  AOI21_X1 U4846 ( .B1(n4167), .B2(n4625), .A(n4166), .ZN(n4304) );
  NAND2_X1 U4847 ( .A1(n4192), .A2(n4168), .ZN(n4169) );
  NAND2_X1 U4848 ( .A1(n4170), .A2(n4169), .ZN(n4390) );
  INV_X1 U4849 ( .A(n4390), .ZN(n4180) );
  OAI22_X1 U4850 ( .A1(n4172), .A2(n4559), .B1(n4431), .B2(n4171), .ZN(n4179)
         );
  NAND2_X1 U4851 ( .A1(n4174), .A2(n4173), .ZN(n4175) );
  NAND2_X1 U4852 ( .A1(n4176), .A2(n4175), .ZN(n4302) );
  NOR2_X1 U4853 ( .A1(n4302), .A2(n4177), .ZN(n4178) );
  AOI211_X1 U4854 ( .C1(n4180), .C2(n4632), .A(n4179), .B(n4178), .ZN(n4181)
         );
  OAI21_X1 U4855 ( .B1(n4626), .B2(n4304), .A(n4181), .ZN(U3274) );
  NAND2_X1 U4856 ( .A1(n4206), .A2(n4182), .ZN(n4184) );
  INV_X1 U4857 ( .A(n4190), .ZN(n4183) );
  XNOR2_X1 U4858 ( .A(n4184), .B(n4183), .ZN(n4185) );
  NAND2_X1 U4859 ( .A1(n4185), .A2(n4625), .ZN(n4310) );
  NAND2_X1 U4860 ( .A1(n4187), .A2(n4186), .ZN(n4204) );
  NOR2_X1 U4861 ( .A1(n4204), .A2(n4205), .ZN(n4203) );
  NOR2_X1 U4862 ( .A1(n4203), .A2(n4188), .ZN(n4189) );
  XOR2_X1 U4863 ( .A(n4190), .B(n4189), .Z(n4312) );
  NAND2_X1 U4864 ( .A1(n4312), .A2(n4191), .ZN(n4202) );
  OAI21_X1 U4865 ( .B1(n4211), .B2(n4198), .A(n4192), .ZN(n4394) );
  INV_X1 U4866 ( .A(n4394), .ZN(n4200) );
  AOI22_X1 U4867 ( .A1(n4216), .A2(n4193), .B1(n4214), .B2(n4308), .ZN(n4197)
         );
  INV_X1 U4868 ( .A(n4194), .ZN(n4195) );
  AOI22_X1 U4869 ( .A1(n4626), .A2(REG2_REG_15__SCAN_IN), .B1(n4195), .B2(
        n4627), .ZN(n4196) );
  OAI211_X1 U4870 ( .C1(n4198), .C2(n4221), .A(n4197), .B(n4196), .ZN(n4199)
         );
  AOI21_X1 U4871 ( .B1(n4200), .B2(n4632), .A(n4199), .ZN(n4201) );
  OAI211_X1 U4872 ( .C1(n4626), .C2(n4310), .A(n4202), .B(n4201), .ZN(U3275)
         );
  AOI21_X1 U4873 ( .B1(n4205), .B2(n4204), .A(n4203), .ZN(n4315) );
  INV_X1 U4874 ( .A(n4206), .ZN(n4207) );
  AOI21_X1 U4875 ( .B1(n2229), .B2(n4208), .A(n4207), .ZN(n4209) );
  OAI22_X1 U4876 ( .A1(n4315), .A2(n4621), .B1(n4333), .B2(n4209), .ZN(n4322)
         );
  NAND2_X1 U4877 ( .A1(n4322), .A2(n4172), .ZN(n4226) );
  INV_X1 U4878 ( .A(n4210), .ZN(n4213) );
  INV_X1 U4879 ( .A(n4211), .ZN(n4212) );
  OAI21_X1 U4880 ( .B1(n4213), .B2(n4222), .A(n4212), .ZN(n4398) );
  INV_X1 U4881 ( .A(n4398), .ZN(n4224) );
  AOI22_X1 U4882 ( .A1(n4216), .A2(n4215), .B1(n4214), .B2(n4318), .ZN(n4220)
         );
  INV_X1 U4883 ( .A(n4217), .ZN(n4218) );
  AOI22_X1 U4884 ( .A1(n4626), .A2(REG2_REG_14__SCAN_IN), .B1(n4218), .B2(
        n4627), .ZN(n4219) );
  OAI211_X1 U4885 ( .C1(n4222), .C2(n4221), .A(n4220), .B(n4219), .ZN(n4223)
         );
  AOI21_X1 U4886 ( .B1(n4224), .B2(n4632), .A(n4223), .ZN(n4225) );
  OAI211_X1 U4887 ( .C1(n4315), .C2(n4227), .A(n4226), .B(n4225), .ZN(U3276)
         );
  NOR2_X1 U4888 ( .A1(n4340), .A2(n4714), .ZN(n4228) );
  AOI21_X1 U4889 ( .B1(REG1_REG_31__SCAN_IN), .B2(n4714), .A(n4228), .ZN(n4229) );
  OAI21_X1 U4890 ( .B1(n4343), .B2(n4339), .A(n4229), .ZN(U3549) );
  AOI21_X1 U4891 ( .B1(n4233), .B2(n4231), .A(n4230), .ZN(n4433) );
  INV_X1 U4892 ( .A(n4433), .ZN(n4345) );
  INV_X1 U4893 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4234) );
  AOI21_X1 U4894 ( .B1(n4233), .B2(n4611), .A(n4232), .ZN(n4435) );
  MUX2_X1 U4895 ( .A(n4234), .B(n4435), .S(n4717), .Z(n4235) );
  OAI21_X1 U4896 ( .B1(n4345), .B2(n4339), .A(n4235), .ZN(U3548) );
  INV_X1 U4897 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4243) );
  AOI22_X1 U4898 ( .A1(n4237), .A2(n4613), .B1(n4236), .B2(n4611), .ZN(n4238)
         );
  OAI211_X1 U4899 ( .C1(n4240), .C2(n4616), .A(n4239), .B(n4238), .ZN(n4241)
         );
  AOI21_X1 U4900 ( .B1(n4242), .B2(n4678), .A(n4241), .ZN(n4346) );
  MUX2_X1 U4901 ( .A(n4243), .B(n4346), .S(n4717), .Z(n4244) );
  OAI21_X1 U4902 ( .B1(n4339), .B2(n4349), .A(n4244), .ZN(U3545) );
  INV_X1 U4903 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4247) );
  AOI21_X1 U4904 ( .B1(n4246), .B2(n4678), .A(n4245), .ZN(n4350) );
  MUX2_X1 U4905 ( .A(n4247), .B(n4350), .S(n4717), .Z(n4248) );
  OAI21_X1 U4906 ( .B1(n4339), .B2(n4353), .A(n4248), .ZN(U3544) );
  AOI21_X1 U4907 ( .B1(n4250), .B2(n4678), .A(n4249), .ZN(n4354) );
  MUX2_X1 U4908 ( .A(n4251), .B(n4354), .S(n4717), .Z(n4252) );
  OAI21_X1 U4909 ( .B1(n4339), .B2(n4357), .A(n4252), .ZN(U3543) );
  AOI21_X1 U4910 ( .B1(n4254), .B2(n4678), .A(n4253), .ZN(n4358) );
  MUX2_X1 U4911 ( .A(n4255), .B(n4358), .S(n4717), .Z(n4256) );
  OAI21_X1 U4912 ( .B1(n4339), .B2(n4361), .A(n4256), .ZN(U3542) );
  INV_X1 U4913 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4259) );
  AOI21_X1 U4914 ( .B1(n4258), .B2(n4678), .A(n4257), .ZN(n4362) );
  MUX2_X1 U4915 ( .A(n4259), .B(n4362), .S(n4717), .Z(n4260) );
  OAI21_X1 U4916 ( .B1(n4339), .B2(n4365), .A(n4260), .ZN(U3541) );
  OR2_X1 U4917 ( .A1(n4261), .A2(n4301), .ZN(n4263) );
  NAND2_X1 U4918 ( .A1(n4263), .A2(n4262), .ZN(n4366) );
  MUX2_X1 U4919 ( .A(n4366), .B(REG1_REG_22__SCAN_IN), .S(n4714), .Z(n4264) );
  INV_X1 U4920 ( .A(n4264), .ZN(n4265) );
  OAI21_X1 U4921 ( .B1(n4339), .B2(n4369), .A(n4265), .ZN(U3540) );
  INV_X1 U4922 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4273) );
  AOI22_X1 U4923 ( .A1(n4267), .A2(n4317), .B1(n4611), .B2(n4266), .ZN(n4268)
         );
  OAI21_X1 U4924 ( .B1(n4269), .B2(n4320), .A(n4268), .ZN(n4270) );
  AOI211_X1 U4925 ( .C1(n4272), .C2(n4678), .A(n4271), .B(n4270), .ZN(n4370)
         );
  MUX2_X1 U4926 ( .A(n4273), .B(n4370), .S(n4717), .Z(n4274) );
  OAI21_X1 U4927 ( .B1(n4339), .B2(n4373), .A(n4274), .ZN(U3539) );
  INV_X1 U4928 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4283) );
  OAI22_X1 U4929 ( .A1(n4276), .A2(n4616), .B1(n4328), .B2(n4275), .ZN(n4277)
         );
  AOI21_X1 U4930 ( .B1(n4613), .B2(n4278), .A(n4277), .ZN(n4279) );
  OAI21_X1 U4931 ( .B1(n4280), .B2(n4333), .A(n4279), .ZN(n4281) );
  AOI21_X1 U4932 ( .B1(n4282), .B2(n4678), .A(n4281), .ZN(n4374) );
  MUX2_X1 U4933 ( .A(n4283), .B(n4374), .S(n4717), .Z(n4284) );
  OAI21_X1 U4934 ( .B1(n4339), .B2(n4377), .A(n4284), .ZN(U3538) );
  AOI21_X1 U4935 ( .B1(n4286), .B2(n4678), .A(n4285), .ZN(n4378) );
  MUX2_X1 U4936 ( .A(n4287), .B(n4378), .S(n4717), .Z(n4288) );
  OAI21_X1 U4937 ( .B1(n4339), .B2(n4381), .A(n4288), .ZN(U3537) );
  OAI211_X1 U4938 ( .C1(n4291), .C2(n4301), .A(n4290), .B(n4289), .ZN(n4382)
         );
  MUX2_X1 U4939 ( .A(REG1_REG_18__SCAN_IN), .B(n4382), .S(n4717), .Z(U3536) );
  AOI22_X1 U4940 ( .A1(n4293), .A2(n4317), .B1(n4611), .B2(n4292), .ZN(n4294)
         );
  OAI211_X1 U4941 ( .C1(n4296), .C2(n4320), .A(n4295), .B(n4294), .ZN(n4297)
         );
  AOI21_X1 U4942 ( .B1(n4298), .B2(n4678), .A(n4297), .ZN(n4383) );
  MUX2_X1 U4943 ( .A(n4299), .B(n4383), .S(n4717), .Z(n4300) );
  OAI21_X1 U4944 ( .B1(n4339), .B2(n4386), .A(n4300), .ZN(U3535) );
  OR2_X1 U4945 ( .A1(n4302), .A2(n4301), .ZN(n4303) );
  NAND2_X1 U4946 ( .A1(n4304), .A2(n4303), .ZN(n4387) );
  MUX2_X1 U4947 ( .A(n4387), .B(REG1_REG_16__SCAN_IN), .S(n4714), .Z(n4305) );
  INV_X1 U4948 ( .A(n4305), .ZN(n4306) );
  OAI21_X1 U4949 ( .B1(n4339), .B2(n4390), .A(n4306), .ZN(U3534) );
  AOI22_X1 U4950 ( .A1(n4308), .A2(n4317), .B1(n4611), .B2(n4307), .ZN(n4309)
         );
  OAI211_X1 U4951 ( .C1(n4329), .C2(n4320), .A(n4310), .B(n4309), .ZN(n4311)
         );
  AOI21_X1 U4952 ( .B1(n4312), .B2(n4678), .A(n4311), .ZN(n4391) );
  MUX2_X1 U4953 ( .A(n4313), .B(n4391), .S(n4717), .Z(n4314) );
  OAI21_X1 U4954 ( .B1(n4339), .B2(n4394), .A(n4314), .ZN(U3533) );
  INV_X1 U4955 ( .A(n4315), .ZN(n4324) );
  AOI22_X1 U4956 ( .A1(n4318), .A2(n4317), .B1(n4611), .B2(n4316), .ZN(n4319)
         );
  OAI21_X1 U4957 ( .B1(n4321), .B2(n4320), .A(n4319), .ZN(n4323) );
  AOI211_X1 U4958 ( .C1(n4689), .C2(n4324), .A(n4323), .B(n4322), .ZN(n4395)
         );
  MUX2_X1 U4959 ( .A(n4325), .B(n4395), .S(n4717), .Z(n4326) );
  OAI21_X1 U4960 ( .B1(n4339), .B2(n4398), .A(n4326), .ZN(U3532) );
  OAI22_X1 U4961 ( .A1(n4329), .A2(n4616), .B1(n4328), .B2(n4327), .ZN(n4330)
         );
  AOI21_X1 U4962 ( .B1(n4613), .B2(n4331), .A(n4330), .ZN(n4332) );
  OAI21_X1 U4963 ( .B1(n4334), .B2(n4333), .A(n4332), .ZN(n4335) );
  AOI21_X1 U4964 ( .B1(n4336), .B2(n4678), .A(n4335), .ZN(n4399) );
  MUX2_X1 U4965 ( .A(n4337), .B(n4399), .S(n4717), .Z(n4338) );
  OAI21_X1 U4966 ( .B1(n4339), .B2(n4403), .A(n4338), .ZN(U3531) );
  MUX2_X1 U4967 ( .A(n4341), .B(n4340), .S(n4701), .Z(n4342) );
  OAI21_X1 U4968 ( .B1(n4343), .B2(n4402), .A(n4342), .ZN(U3517) );
  MUX2_X1 U4969 ( .A(n2878), .B(n4435), .S(n4701), .Z(n4344) );
  OAI21_X1 U4970 ( .B1(n4345), .B2(n4402), .A(n4344), .ZN(U3516) );
  INV_X1 U4971 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4347) );
  MUX2_X1 U4972 ( .A(n4347), .B(n4346), .S(n4701), .Z(n4348) );
  OAI21_X1 U4973 ( .B1(n4349), .B2(n4402), .A(n4348), .ZN(U3513) );
  INV_X1 U4974 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4351) );
  MUX2_X1 U4975 ( .A(n4351), .B(n4350), .S(n4701), .Z(n4352) );
  OAI21_X1 U4976 ( .B1(n4353), .B2(n4402), .A(n4352), .ZN(U3512) );
  INV_X1 U4977 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4355) );
  MUX2_X1 U4978 ( .A(n4355), .B(n4354), .S(n4701), .Z(n4356) );
  OAI21_X1 U4979 ( .B1(n4357), .B2(n4402), .A(n4356), .ZN(U3511) );
  INV_X1 U4980 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4359) );
  MUX2_X1 U4981 ( .A(n4359), .B(n4358), .S(n4701), .Z(n4360) );
  OAI21_X1 U4982 ( .B1(n4361), .B2(n4402), .A(n4360), .ZN(U3510) );
  INV_X1 U4983 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4363) );
  MUX2_X1 U4984 ( .A(n4363), .B(n4362), .S(n4701), .Z(n4364) );
  OAI21_X1 U4985 ( .B1(n4365), .B2(n4402), .A(n4364), .ZN(U3509) );
  MUX2_X1 U4986 ( .A(REG0_REG_22__SCAN_IN), .B(n4366), .S(n4701), .Z(n4367) );
  INV_X1 U4987 ( .A(n4367), .ZN(n4368) );
  OAI21_X1 U4988 ( .B1(n4369), .B2(n4402), .A(n4368), .ZN(U3508) );
  INV_X1 U4989 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4371) );
  MUX2_X1 U4990 ( .A(n4371), .B(n4370), .S(n4701), .Z(n4372) );
  OAI21_X1 U4991 ( .B1(n4373), .B2(n4402), .A(n4372), .ZN(U3507) );
  INV_X1 U4992 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4375) );
  MUX2_X1 U4993 ( .A(n4375), .B(n4374), .S(n4701), .Z(n4376) );
  OAI21_X1 U4994 ( .B1(n4377), .B2(n4402), .A(n4376), .ZN(U3506) );
  INV_X1 U4995 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4379) );
  MUX2_X1 U4996 ( .A(n4379), .B(n4378), .S(n4701), .Z(n4380) );
  OAI21_X1 U4997 ( .B1(n4381), .B2(n4402), .A(n4380), .ZN(U3505) );
  MUX2_X1 U4998 ( .A(REG0_REG_18__SCAN_IN), .B(n4382), .S(n4701), .Z(U3503) );
  INV_X1 U4999 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4384) );
  MUX2_X1 U5000 ( .A(n4384), .B(n4383), .S(n4701), .Z(n4385) );
  OAI21_X1 U5001 ( .B1(n4386), .B2(n4402), .A(n4385), .ZN(U3501) );
  MUX2_X1 U5002 ( .A(n4387), .B(REG0_REG_16__SCAN_IN), .S(n4699), .Z(n4388) );
  INV_X1 U5003 ( .A(n4388), .ZN(n4389) );
  OAI21_X1 U5004 ( .B1(n4390), .B2(n4402), .A(n4389), .ZN(U3499) );
  INV_X1 U5005 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4392) );
  MUX2_X1 U5006 ( .A(n4392), .B(n4391), .S(n4701), .Z(n4393) );
  OAI21_X1 U5007 ( .B1(n4394), .B2(n4402), .A(n4393), .ZN(U3497) );
  INV_X1 U5008 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4396) );
  MUX2_X1 U5009 ( .A(n4396), .B(n4395), .S(n4701), .Z(n4397) );
  OAI21_X1 U5010 ( .B1(n4398), .B2(n4402), .A(n4397), .ZN(U3495) );
  INV_X1 U5011 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4400) );
  MUX2_X1 U5012 ( .A(n4400), .B(n4399), .S(n4701), .Z(n4401) );
  OAI21_X1 U5013 ( .B1(n4403), .B2(n4402), .A(n4401), .ZN(U3493) );
  MUX2_X1 U5014 ( .A(n4404), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5015 ( .A(DATAI_24_), .B(n4405), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U5016 ( .A(DATAI_22_), .B(n4406), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U5017 ( .A(DATAI_20_), .B(n4407), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5018 ( .A(DATAI_4_), .B(n4408), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5019 ( .A(DATAI_3_), .B(n4409), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5020 ( .A(n4410), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5021 ( .A(n4411), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U5022 ( .A(DATAI_28_), .ZN(n4412) );
  AOI22_X1 U5023 ( .A1(STATE_REG_SCAN_IN), .A2(n4413), .B1(n4412), .B2(U3149), 
        .ZN(U3324) );
  NOR2_X1 U5024 ( .A1(STATE_REG_SCAN_IN), .A2(n4414), .ZN(n4563) );
  OAI22_X1 U5025 ( .A1(n4418), .A2(n4417), .B1(n4416), .B2(n4415), .ZN(n4419)
         );
  AOI211_X1 U5026 ( .C1(n4421), .C2(n4420), .A(n4563), .B(n4419), .ZN(n4430)
         );
  OAI21_X1 U5027 ( .B1(n3420), .B2(n4424), .A(n4423), .ZN(n4426) );
  XNOR2_X1 U5028 ( .A(n4426), .B(n4425), .ZN(n4428) );
  NAND2_X1 U5029 ( .A1(n4428), .A2(n4427), .ZN(n4429) );
  OAI211_X1 U5030 ( .C1(n4432), .C2(n4431), .A(n4430), .B(n4429), .ZN(U3223)
         );
  AOI22_X1 U5031 ( .A1(n4433), .A2(n4632), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4626), .ZN(n4434) );
  OAI21_X1 U5032 ( .B1(n4626), .B2(n4435), .A(n4434), .ZN(U3261) );
  OAI211_X1 U5033 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4437), .A(n4439), .B(n4436), 
        .ZN(n4442) );
  AOI22_X1 U5034 ( .A1(n4439), .A2(n4438), .B1(n4585), .B2(n2934), .ZN(n4441)
         );
  AOI22_X1 U5035 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4583), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4440) );
  OAI221_X1 U5036 ( .B1(IR_REG_0__SCAN_IN), .B2(n4442), .C1(n2928), .C2(n4441), 
        .A(n4440), .ZN(U3240) );
  INV_X1 U5037 ( .A(n4585), .ZN(n4453) );
  AOI211_X1 U5038 ( .C1(n4445), .C2(n4444), .A(n4443), .B(n4453), .ZN(n4447)
         );
  AOI211_X1 U5039 ( .C1(n4583), .C2(ADDR_REG_5__SCAN_IN), .A(n4447), .B(n4446), 
        .ZN(n4452) );
  OAI211_X1 U5040 ( .C1(n4450), .C2(n4449), .A(n4528), .B(n4448), .ZN(n4451)
         );
  OAI211_X1 U5041 ( .C1(n4590), .C2(n4657), .A(n4452), .B(n4451), .ZN(U3245)
         );
  AOI211_X1 U5042 ( .C1(n4456), .C2(n4455), .A(n4454), .B(n4453), .ZN(n4458)
         );
  AOI211_X1 U5043 ( .C1(n4583), .C2(ADDR_REG_6__SCAN_IN), .A(n4458), .B(n4457), 
        .ZN(n4462) );
  OAI211_X1 U5044 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4460), .A(n4528), .B(n4459), 
        .ZN(n4461) );
  OAI211_X1 U5045 ( .C1(n4590), .C2(n4656), .A(n4462), .B(n4461), .ZN(U3246)
         );
  NAND2_X1 U5046 ( .A1(n2261), .A2(n4463), .ZN(n4465) );
  OAI21_X1 U5047 ( .B1(n4466), .B2(n4465), .A(n4585), .ZN(n4464) );
  AOI21_X1 U5048 ( .B1(n4466), .B2(n4465), .A(n4464), .ZN(n4468) );
  AOI211_X1 U5049 ( .C1(n4583), .C2(ADDR_REG_7__SCAN_IN), .A(n4468), .B(n4467), 
        .ZN(n4473) );
  OAI211_X1 U5050 ( .C1(n4471), .C2(n4470), .A(n4528), .B(n4469), .ZN(n4472)
         );
  OAI211_X1 U5051 ( .C1(n4590), .C2(n4655), .A(n4473), .B(n4472), .ZN(U3247)
         );
  OAI211_X1 U5052 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4476), .A(n4528), .B(n4475), 
        .ZN(n4478) );
  NAND2_X1 U5053 ( .A1(n4478), .A2(n4477), .ZN(n4479) );
  AOI21_X1 U5054 ( .B1(n4583), .B2(ADDR_REG_8__SCAN_IN), .A(n4479), .ZN(n4483)
         );
  OAI211_X1 U5055 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4481), .A(n4585), .B(n4480), 
        .ZN(n4482) );
  OAI211_X1 U5056 ( .C1(n4590), .C2(n2386), .A(n4483), .B(n4482), .ZN(U3248)
         );
  OAI211_X1 U5057 ( .C1(n4486), .C2(n4485), .A(n4585), .B(n4484), .ZN(n4491)
         );
  OAI211_X1 U5058 ( .C1(n4489), .C2(n4488), .A(n4528), .B(n4487), .ZN(n4490)
         );
  OAI211_X1 U5059 ( .C1(n4590), .C2(n4654), .A(n4491), .B(n4490), .ZN(n4492)
         );
  AOI211_X1 U5060 ( .C1(n4583), .C2(ADDR_REG_9__SCAN_IN), .A(n4493), .B(n4492), 
        .ZN(n4494) );
  INV_X1 U5061 ( .A(n4494), .ZN(U3249) );
  OAI211_X1 U5062 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4497), .A(n4528), .B(n4496), .ZN(n4499) );
  NAND2_X1 U5063 ( .A1(n4499), .A2(n4498), .ZN(n4500) );
  AOI21_X1 U5064 ( .B1(n4583), .B2(ADDR_REG_10__SCAN_IN), .A(n4500), .ZN(n4504) );
  OAI211_X1 U5065 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4502), .A(n4585), .B(n4501), .ZN(n4503) );
  OAI211_X1 U5066 ( .C1(n4590), .C2(n2385), .A(n4504), .B(n4503), .ZN(U3250)
         );
  OAI211_X1 U5067 ( .C1(n4507), .C2(n4506), .A(n4585), .B(n4505), .ZN(n4512)
         );
  OAI211_X1 U5068 ( .C1(n4510), .C2(n4509), .A(n4528), .B(n4508), .ZN(n4511)
         );
  OAI211_X1 U5069 ( .C1(n4590), .C2(n4653), .A(n4512), .B(n4511), .ZN(n4513)
         );
  AOI211_X1 U5070 ( .C1(n4583), .C2(ADDR_REG_11__SCAN_IN), .A(n4514), .B(n4513), .ZN(n4515) );
  INV_X1 U5071 ( .A(n4515), .ZN(U3251) );
  OAI211_X1 U5072 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4518), .A(n4528), .B(n4517), .ZN(n4520) );
  NAND2_X1 U5073 ( .A1(n4520), .A2(n4519), .ZN(n4521) );
  AOI21_X1 U5074 ( .B1(n4583), .B2(ADDR_REG_12__SCAN_IN), .A(n4521), .ZN(n4525) );
  OAI211_X1 U5075 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4523), .A(n4585), .B(n4522), .ZN(n4524) );
  OAI211_X1 U5076 ( .C1(n4590), .C2(n2384), .A(n4525), .B(n4524), .ZN(U3252)
         );
  AOI21_X1 U5077 ( .B1(n4527), .B2(n4651), .A(n4526), .ZN(n4531) );
  OAI21_X1 U5078 ( .B1(n4531), .B2(n4530), .A(n4528), .ZN(n4529) );
  AOI21_X1 U5079 ( .B1(n4531), .B2(n4530), .A(n4529), .ZN(n4532) );
  AOI211_X1 U5080 ( .C1(n4583), .C2(ADDR_REG_13__SCAN_IN), .A(n4533), .B(n4532), .ZN(n4538) );
  OAI211_X1 U5081 ( .C1(n4536), .C2(n4535), .A(n4585), .B(n4534), .ZN(n4537)
         );
  OAI211_X1 U5082 ( .C1(n4590), .C2(n4651), .A(n4538), .B(n4537), .ZN(U3253)
         );
  AOI211_X1 U5083 ( .C1(n4541), .C2(n4540), .A(n4539), .B(n4579), .ZN(n4542)
         );
  AOI211_X1 U5084 ( .C1(n4583), .C2(ADDR_REG_14__SCAN_IN), .A(n4543), .B(n4542), .ZN(n4547) );
  OAI211_X1 U5085 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4545), .A(n4585), .B(n4544), .ZN(n4546) );
  OAI211_X1 U5086 ( .C1(n4590), .C2(n4650), .A(n4547), .B(n4546), .ZN(U3254)
         );
  AOI211_X1 U5087 ( .C1(n4550), .C2(n4549), .A(n4548), .B(n4579), .ZN(n4551)
         );
  AOI211_X1 U5088 ( .C1(n4583), .C2(ADDR_REG_15__SCAN_IN), .A(n4552), .B(n4551), .ZN(n4557) );
  OAI211_X1 U5089 ( .C1(n4555), .C2(n4554), .A(n4585), .B(n4553), .ZN(n4556)
         );
  OAI211_X1 U5090 ( .C1(n4590), .C2(n4558), .A(n4557), .B(n4556), .ZN(U3255)
         );
  AOI221_X1 U5091 ( .B1(n4561), .B2(n4560), .C1(n4559), .C2(n4560), .A(n4579), 
        .ZN(n4562) );
  AOI211_X1 U5092 ( .C1(n4583), .C2(ADDR_REG_16__SCAN_IN), .A(n4563), .B(n4562), .ZN(n4567) );
  OAI221_X1 U5093 ( .B1(n4565), .B2(REG1_REG_16__SCAN_IN), .C1(n4565), .C2(
        n4564), .A(n4585), .ZN(n4566) );
  OAI211_X1 U5094 ( .C1(n4590), .C2(n4647), .A(n4567), .B(n4566), .ZN(U3256)
         );
  AOI221_X1 U5095 ( .B1(n4570), .B2(n4569), .C1(n4568), .C2(n4569), .A(n4579), 
        .ZN(n4571) );
  AOI211_X1 U5096 ( .C1(n4583), .C2(ADDR_REG_17__SCAN_IN), .A(n4572), .B(n4571), .ZN(n4577) );
  OAI221_X1 U5097 ( .B1(n4575), .B2(n4574), .C1(n4575), .C2(n4573), .A(n4585), 
        .ZN(n4576) );
  OAI211_X1 U5098 ( .C1(n4590), .C2(n4645), .A(n4577), .B(n4576), .ZN(U3257)
         );
  NOR2_X1 U5099 ( .A1(STATE_REG_SCAN_IN), .A2(n4578), .ZN(n4582) );
  OAI211_X1 U5100 ( .C1(n4587), .C2(n4586), .A(n4585), .B(n4584), .ZN(n4588)
         );
  OAI211_X1 U5101 ( .C1(n4590), .C2(n4644), .A(n4589), .B(n4588), .ZN(U3258)
         );
  XOR2_X1 U5102 ( .A(n4597), .B(n4591), .Z(n4600) );
  AOI22_X1 U5103 ( .A1(n4593), .A2(n4613), .B1(n4592), .B2(n4611), .ZN(n4594)
         );
  OAI21_X1 U5104 ( .B1(n4595), .B2(n4616), .A(n4594), .ZN(n4599) );
  XOR2_X1 U5105 ( .A(n4597), .B(n4596), .Z(n4696) );
  NOR2_X1 U5106 ( .A1(n4696), .A2(n4621), .ZN(n4598) );
  AOI211_X1 U5107 ( .C1(n4600), .C2(n4625), .A(n4599), .B(n4598), .ZN(n4692)
         );
  INV_X1 U5108 ( .A(n4601), .ZN(n4602) );
  AOI22_X1 U5109 ( .A1(n4602), .A2(n4627), .B1(REG2_REG_11__SCAN_IN), .B2(
        n4626), .ZN(n4608) );
  INV_X1 U5110 ( .A(n4696), .ZN(n4606) );
  OAI21_X1 U5111 ( .B1(n4685), .B2(n4604), .A(n4603), .ZN(n4693) );
  INV_X1 U5112 ( .A(n4693), .ZN(n4605) );
  AOI22_X1 U5113 ( .A1(n4606), .A2(n4633), .B1(n4632), .B2(n4605), .ZN(n4607)
         );
  OAI211_X1 U5114 ( .C1(n4626), .C2(n4692), .A(n4608), .B(n4607), .ZN(U3279)
         );
  INV_X1 U5115 ( .A(n4620), .ZN(n4610) );
  OAI21_X1 U5116 ( .B1(n4610), .B2(n2352), .A(n4609), .ZN(n4624) );
  AOI22_X1 U5117 ( .A1(n4614), .A2(n4613), .B1(n4612), .B2(n4611), .ZN(n4615)
         );
  OAI21_X1 U5118 ( .B1(n4617), .B2(n4616), .A(n4615), .ZN(n4623) );
  OAI21_X1 U5119 ( .B1(n4620), .B2(n4619), .A(n4618), .ZN(n4663) );
  NOR2_X1 U5120 ( .A1(n4663), .A2(n4621), .ZN(n4622) );
  AOI211_X1 U5121 ( .C1(n4625), .C2(n4624), .A(n4623), .B(n4622), .ZN(n4661)
         );
  AOI22_X1 U5122 ( .A1(REG3_REG_1__SCAN_IN), .A2(n4627), .B1(
        REG2_REG_1__SCAN_IN), .B2(n4626), .ZN(n4636) );
  INV_X1 U5123 ( .A(n4663), .ZN(n4634) );
  OAI21_X1 U5124 ( .B1(n4630), .B2(n4629), .A(n4628), .ZN(n4662) );
  INV_X1 U5125 ( .A(n4662), .ZN(n4631) );
  AOI22_X1 U5126 ( .A1(n4634), .A2(n4633), .B1(n4632), .B2(n4631), .ZN(n4635)
         );
  OAI211_X1 U5127 ( .C1(n4626), .C2(n4661), .A(n4636), .B(n4635), .ZN(U3289)
         );
  INV_X1 U5128 ( .A(D_REG_31__SCAN_IN), .ZN(n4997) );
  NOR2_X1 U5129 ( .A1(n4642), .A2(n4997), .ZN(U3291) );
  INV_X1 U5130 ( .A(D_REG_30__SCAN_IN), .ZN(n5020) );
  NOR2_X1 U5131 ( .A1(n4642), .A2(n5020), .ZN(U3292) );
  INV_X1 U5132 ( .A(D_REG_29__SCAN_IN), .ZN(n4840) );
  NOR2_X1 U5133 ( .A1(n4642), .A2(n4840), .ZN(U3293) );
  INV_X1 U5134 ( .A(D_REG_28__SCAN_IN), .ZN(n4828) );
  NOR2_X1 U5135 ( .A1(n4642), .A2(n4828), .ZN(U3294) );
  INV_X1 U5136 ( .A(D_REG_27__SCAN_IN), .ZN(n5036) );
  NOR2_X1 U5137 ( .A1(n4642), .A2(n5036), .ZN(U3295) );
  INV_X1 U5138 ( .A(D_REG_26__SCAN_IN), .ZN(n5031) );
  NOR2_X1 U5139 ( .A1(n4642), .A2(n5031), .ZN(U3296) );
  INV_X1 U5140 ( .A(D_REG_25__SCAN_IN), .ZN(n4875) );
  NOR2_X1 U5141 ( .A1(n4642), .A2(n4875), .ZN(U3297) );
  INV_X1 U5142 ( .A(D_REG_24__SCAN_IN), .ZN(n4795) );
  NOR2_X1 U5143 ( .A1(n4642), .A2(n4795), .ZN(U3298) );
  NOR2_X1 U5144 ( .A1(n4642), .A2(n5034), .ZN(U3299) );
  INV_X1 U5145 ( .A(D_REG_22__SCAN_IN), .ZN(n4844) );
  NOR2_X1 U5146 ( .A1(n4642), .A2(n4844), .ZN(U3300) );
  INV_X1 U5147 ( .A(D_REG_21__SCAN_IN), .ZN(n4845) );
  NOR2_X1 U5148 ( .A1(n4642), .A2(n4845), .ZN(U3301) );
  INV_X1 U5149 ( .A(D_REG_20__SCAN_IN), .ZN(n5023) );
  NOR2_X1 U5150 ( .A1(n4642), .A2(n5023), .ZN(U3302) );
  INV_X1 U5151 ( .A(D_REG_19__SCAN_IN), .ZN(n5014) );
  NOR2_X1 U5152 ( .A1(n4642), .A2(n5014), .ZN(U3303) );
  INV_X1 U5153 ( .A(D_REG_18__SCAN_IN), .ZN(n4805) );
  NOR2_X1 U5154 ( .A1(n4642), .A2(n4805), .ZN(U3304) );
  INV_X1 U5155 ( .A(D_REG_17__SCAN_IN), .ZN(n5024) );
  NOR2_X1 U5156 ( .A1(n4642), .A2(n5024), .ZN(U3305) );
  INV_X1 U5157 ( .A(D_REG_16__SCAN_IN), .ZN(n4771) );
  NOR2_X1 U5158 ( .A1(n4642), .A2(n4771), .ZN(U3306) );
  INV_X1 U5159 ( .A(D_REG_15__SCAN_IN), .ZN(n4637) );
  NOR2_X1 U5160 ( .A1(n4642), .A2(n4637), .ZN(U3307) );
  INV_X1 U5161 ( .A(D_REG_14__SCAN_IN), .ZN(n4638) );
  NOR2_X1 U5162 ( .A1(n4642), .A2(n4638), .ZN(U3308) );
  INV_X1 U5163 ( .A(D_REG_13__SCAN_IN), .ZN(n5018) );
  NOR2_X1 U5164 ( .A1(n4642), .A2(n5018), .ZN(U3309) );
  INV_X1 U5165 ( .A(D_REG_12__SCAN_IN), .ZN(n5033) );
  NOR2_X1 U5166 ( .A1(n4642), .A2(n5033), .ZN(U3310) );
  INV_X1 U5167 ( .A(D_REG_11__SCAN_IN), .ZN(n4639) );
  NOR2_X1 U5168 ( .A1(n4642), .A2(n4639), .ZN(U3311) );
  INV_X1 U5169 ( .A(D_REG_10__SCAN_IN), .ZN(n4743) );
  NOR2_X1 U5170 ( .A1(n4642), .A2(n4743), .ZN(U3312) );
  INV_X1 U5171 ( .A(D_REG_9__SCAN_IN), .ZN(n4640) );
  NOR2_X1 U5172 ( .A1(n4642), .A2(n4640), .ZN(U3313) );
  INV_X1 U5173 ( .A(D_REG_8__SCAN_IN), .ZN(n4641) );
  NOR2_X1 U5174 ( .A1(n4642), .A2(n4641), .ZN(U3314) );
  NOR2_X1 U5175 ( .A1(n4642), .A2(n5017), .ZN(U3315) );
  INV_X1 U5176 ( .A(D_REG_6__SCAN_IN), .ZN(n5015) );
  NOR2_X1 U5177 ( .A1(n4642), .A2(n5015), .ZN(U3316) );
  INV_X1 U5178 ( .A(D_REG_5__SCAN_IN), .ZN(n5021) );
  NOR2_X1 U5179 ( .A1(n4642), .A2(n5021), .ZN(U3317) );
  INV_X1 U5180 ( .A(D_REG_4__SCAN_IN), .ZN(n4842) );
  NOR2_X1 U5181 ( .A1(n4642), .A2(n4842), .ZN(U3318) );
  INV_X1 U5182 ( .A(D_REG_3__SCAN_IN), .ZN(n4998) );
  NOR2_X1 U5183 ( .A1(n4642), .A2(n4998), .ZN(U3319) );
  INV_X1 U5184 ( .A(D_REG_2__SCAN_IN), .ZN(n5030) );
  NOR2_X1 U5185 ( .A1(n4642), .A2(n5030), .ZN(U3320) );
  AOI21_X1 U5186 ( .B1(U3149), .B2(n2753), .A(n4643), .ZN(U3329) );
  INV_X1 U5187 ( .A(DATAI_18_), .ZN(n4855) );
  AOI22_X1 U5188 ( .A1(STATE_REG_SCAN_IN), .A2(n4644), .B1(n4855), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5189 ( .A(DATAI_17_), .ZN(n5043) );
  AOI22_X1 U5190 ( .A1(STATE_REG_SCAN_IN), .A2(n4645), .B1(n5043), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5191 ( .A(DATAI_16_), .ZN(n4646) );
  AOI22_X1 U5192 ( .A1(STATE_REG_SCAN_IN), .A2(n4647), .B1(n4646), .B2(U3149), 
        .ZN(U3336) );
  OAI22_X1 U5193 ( .A1(U3149), .A2(n4648), .B1(DATAI_15_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4649) );
  INV_X1 U5194 ( .A(n4649), .ZN(U3337) );
  INV_X1 U5195 ( .A(DATAI_14_), .ZN(n5057) );
  AOI22_X1 U5196 ( .A1(STATE_REG_SCAN_IN), .A2(n4650), .B1(n5057), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5197 ( .A(DATAI_13_), .ZN(n5002) );
  AOI22_X1 U5198 ( .A1(STATE_REG_SCAN_IN), .A2(n4651), .B1(n5002), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5199 ( .A(DATAI_12_), .ZN(n4878) );
  AOI22_X1 U5200 ( .A1(STATE_REG_SCAN_IN), .A2(n2384), .B1(n4878), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5201 ( .A(DATAI_11_), .ZN(n4652) );
  AOI22_X1 U5202 ( .A1(STATE_REG_SCAN_IN), .A2(n4653), .B1(n4652), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5203 ( .A(DATAI_10_), .ZN(n5046) );
  AOI22_X1 U5204 ( .A1(STATE_REG_SCAN_IN), .A2(n2385), .B1(n5046), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5205 ( .A(DATAI_9_), .ZN(n5001) );
  AOI22_X1 U5206 ( .A1(STATE_REG_SCAN_IN), .A2(n4654), .B1(n5001), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5207 ( .A(DATAI_8_), .ZN(n4860) );
  AOI22_X1 U5208 ( .A1(STATE_REG_SCAN_IN), .A2(n2386), .B1(n4860), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U5209 ( .A(DATAI_7_), .ZN(n4802) );
  AOI22_X1 U5210 ( .A1(STATE_REG_SCAN_IN), .A2(n4655), .B1(n4802), .B2(U3149), 
        .ZN(U3345) );
  INV_X1 U5211 ( .A(DATAI_6_), .ZN(n5055) );
  AOI22_X1 U5212 ( .A1(STATE_REG_SCAN_IN), .A2(n4656), .B1(n5055), .B2(U3149), 
        .ZN(U3346) );
  INV_X1 U5213 ( .A(DATAI_5_), .ZN(n4804) );
  AOI22_X1 U5214 ( .A1(STATE_REG_SCAN_IN), .A2(n4657), .B1(n4804), .B2(U3149), 
        .ZN(U3347) );
  AOI211_X1 U5215 ( .C1(n4689), .C2(n4660), .A(n4659), .B(n4658), .ZN(n4702)
         );
  AOI22_X1 U5216 ( .A1(n4701), .A2(n4702), .B1(n2523), .B2(n4699), .ZN(U3467)
         );
  INV_X1 U5217 ( .A(n4661), .ZN(n4665) );
  OAI22_X1 U5218 ( .A1(n4663), .A2(n4695), .B1(n4694), .B2(n4662), .ZN(n4664)
         );
  NOR2_X1 U5219 ( .A1(n4665), .A2(n4664), .ZN(n4704) );
  AOI22_X1 U5220 ( .A1(n4701), .A2(n4704), .B1(n2529), .B2(n4699), .ZN(U3469)
         );
  AOI21_X1 U5221 ( .B1(n4689), .B2(n4667), .A(n4666), .ZN(n4708) );
  INV_X1 U5222 ( .A(n4668), .ZN(n4706) );
  AOI22_X1 U5223 ( .A1(n4706), .A2(n4669), .B1(REG0_REG_2__SCAN_IN), .B2(n4699), .ZN(n4670) );
  OAI21_X1 U5224 ( .B1(n4708), .B2(n4699), .A(n4670), .ZN(U3471) );
  AND2_X1 U5225 ( .A1(n4671), .A2(n4689), .ZN(n4674) );
  INV_X1 U5226 ( .A(n4672), .ZN(n4673) );
  NOR3_X1 U5227 ( .A1(n4675), .A2(n4674), .A3(n4673), .ZN(n4710) );
  AOI22_X1 U5228 ( .A1(n4701), .A2(n4710), .B1(n2552), .B2(n4699), .ZN(U3475)
         );
  AOI211_X1 U5229 ( .C1(n4679), .C2(n4678), .A(n4677), .B(n4676), .ZN(n4711)
         );
  AOI22_X1 U5230 ( .A1(n4701), .A2(n4711), .B1(n2586), .B2(n4699), .ZN(U3481)
         );
  NOR3_X1 U5231 ( .A1(n4681), .A2(n4680), .A3(n4694), .ZN(n4683) );
  AOI211_X1 U5232 ( .C1(n4684), .C2(n4689), .A(n4683), .B(n4682), .ZN(n4712)
         );
  AOI22_X1 U5233 ( .A1(n4701), .A2(n4712), .B1(n2598), .B2(n4699), .ZN(U3483)
         );
  NOR3_X1 U5234 ( .A1(n4686), .A2(n4685), .A3(n4694), .ZN(n4688) );
  AOI211_X1 U5235 ( .C1(n4690), .C2(n4689), .A(n4688), .B(n4687), .ZN(n4713)
         );
  INV_X1 U5236 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4691) );
  AOI22_X1 U5237 ( .A1(n4701), .A2(n4713), .B1(n4691), .B2(n4699), .ZN(U3487)
         );
  INV_X1 U5238 ( .A(n4692), .ZN(n4698) );
  OAI22_X1 U5239 ( .A1(n4696), .A2(n4695), .B1(n4694), .B2(n4693), .ZN(n4697)
         );
  NOR2_X1 U5240 ( .A1(n4698), .A2(n4697), .ZN(n4716) );
  INV_X1 U5241 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4700) );
  AOI22_X1 U5242 ( .A1(n4701), .A2(n4716), .B1(n4700), .B2(n4699), .ZN(U3489)
         );
  AOI22_X1 U5243 ( .A1(n4717), .A2(n4702), .B1(n2934), .B2(n4714), .ZN(U3518)
         );
  INV_X1 U5244 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4703) );
  AOI22_X1 U5245 ( .A1(n4717), .A2(n4704), .B1(n4703), .B2(n4714), .ZN(U3519)
         );
  AOI22_X1 U5246 ( .A1(n4706), .A2(n4705), .B1(REG1_REG_2__SCAN_IN), .B2(n4714), .ZN(n4707) );
  OAI21_X1 U5247 ( .B1(n4708), .B2(n4714), .A(n4707), .ZN(U3520) );
  AOI22_X1 U5248 ( .A1(n4717), .A2(n4710), .B1(n4709), .B2(n4714), .ZN(U3522)
         );
  AOI22_X1 U5249 ( .A1(n4717), .A2(n4711), .B1(n2587), .B2(n4714), .ZN(U3525)
         );
  AOI22_X1 U5250 ( .A1(n4717), .A2(n4712), .B1(n2599), .B2(n4714), .ZN(U3526)
         );
  AOI22_X1 U5251 ( .A1(n4717), .A2(n4713), .B1(n2625), .B2(n4714), .ZN(U3528)
         );
  AOI22_X1 U5252 ( .A1(n4717), .A2(n4716), .B1(n4715), .B2(n4714), .ZN(U3529)
         );
  OAI22_X1 U5253 ( .A1(IR_REG_30__SCAN_IN), .A2(keyinput_g85), .B1(
        REG3_REG_16__SCAN_IN), .B2(keyinput_g46), .ZN(n4718) );
  AOI221_X1 U5254 ( .B1(IR_REG_30__SCAN_IN), .B2(keyinput_g85), .C1(
        keyinput_g46), .C2(REG3_REG_16__SCAN_IN), .A(n4718), .ZN(n4725) );
  OAI22_X1 U5255 ( .A1(DATAI_20_), .A2(keyinput_g11), .B1(DATAI_15_), .B2(
        keyinput_g16), .ZN(n4719) );
  AOI221_X1 U5256 ( .B1(DATAI_20_), .B2(keyinput_g11), .C1(keyinput_g16), .C2(
        DATAI_15_), .A(n4719), .ZN(n4724) );
  OAI22_X1 U5257 ( .A1(IR_REG_25__SCAN_IN), .A2(keyinput_g80), .B1(
        keyinput_g84), .B2(IR_REG_29__SCAN_IN), .ZN(n4720) );
  AOI221_X1 U5258 ( .B1(IR_REG_25__SCAN_IN), .B2(keyinput_g80), .C1(
        IR_REG_29__SCAN_IN), .C2(keyinput_g84), .A(n4720), .ZN(n4723) );
  OAI22_X1 U5259 ( .A1(D_REG_6__SCAN_IN), .A2(keyinput_g93), .B1(keyinput_g7), 
        .B2(DATAI_24_), .ZN(n4721) );
  AOI221_X1 U5260 ( .B1(D_REG_6__SCAN_IN), .B2(keyinput_g93), .C1(DATAI_24_), 
        .C2(keyinput_g7), .A(n4721), .ZN(n4722) );
  NAND4_X1 U5261 ( .A1(n4725), .A2(n4724), .A3(n4723), .A4(n4722), .ZN(n4756)
         );
  OAI22_X1 U5262 ( .A1(IR_REG_13__SCAN_IN), .A2(keyinput_g68), .B1(
        REG3_REG_19__SCAN_IN), .B2(keyinput_g39), .ZN(n4726) );
  AOI221_X1 U5263 ( .B1(IR_REG_13__SCAN_IN), .B2(keyinput_g68), .C1(
        keyinput_g39), .C2(REG3_REG_19__SCAN_IN), .A(n4726), .ZN(n4733) );
  OAI22_X1 U5264 ( .A1(IR_REG_12__SCAN_IN), .A2(keyinput_g67), .B1(DATAI_10_), 
        .B2(keyinput_g21), .ZN(n4727) );
  AOI221_X1 U5265 ( .B1(IR_REG_12__SCAN_IN), .B2(keyinput_g67), .C1(
        keyinput_g21), .C2(DATAI_10_), .A(n4727), .ZN(n4732) );
  OAI22_X1 U5266 ( .A1(IR_REG_17__SCAN_IN), .A2(keyinput_g72), .B1(
        keyinput_g35), .B2(REG3_REG_14__SCAN_IN), .ZN(n4728) );
  AOI221_X1 U5267 ( .B1(IR_REG_17__SCAN_IN), .B2(keyinput_g72), .C1(
        REG3_REG_14__SCAN_IN), .C2(keyinput_g35), .A(n4728), .ZN(n4731) );
  OAI22_X1 U5268 ( .A1(IR_REG_14__SCAN_IN), .A2(keyinput_g69), .B1(
        keyinput_g102), .B2(D_REG_15__SCAN_IN), .ZN(n4729) );
  AOI221_X1 U5269 ( .B1(IR_REG_14__SCAN_IN), .B2(keyinput_g69), .C1(
        D_REG_15__SCAN_IN), .C2(keyinput_g102), .A(n4729), .ZN(n4730) );
  NAND4_X1 U5270 ( .A1(n4733), .A2(n4732), .A3(n4731), .A4(n4730), .ZN(n4755)
         );
  OAI22_X1 U5271 ( .A1(IR_REG_4__SCAN_IN), .A2(keyinput_g59), .B1(keyinput_g9), 
        .B2(DATAI_22_), .ZN(n4734) );
  AOI221_X1 U5272 ( .B1(IR_REG_4__SCAN_IN), .B2(keyinput_g59), .C1(DATAI_22_), 
        .C2(keyinput_g9), .A(n4734), .ZN(n4741) );
  OAI22_X1 U5273 ( .A1(D_REG_1__SCAN_IN), .A2(keyinput_g88), .B1(keyinput_g95), 
        .B2(D_REG_8__SCAN_IN), .ZN(n4735) );
  AOI221_X1 U5274 ( .B1(D_REG_1__SCAN_IN), .B2(keyinput_g88), .C1(
        D_REG_8__SCAN_IN), .C2(keyinput_g95), .A(n4735), .ZN(n4740) );
  OAI22_X1 U5275 ( .A1(REG0_REG_8__SCAN_IN), .A2(keyinput_g127), .B1(
        REG0_REG_7__SCAN_IN), .B2(keyinput_g126), .ZN(n4736) );
  AOI221_X1 U5276 ( .B1(REG0_REG_8__SCAN_IN), .B2(keyinput_g127), .C1(
        keyinput_g126), .C2(REG0_REG_7__SCAN_IN), .A(n4736), .ZN(n4739) );
  OAI22_X1 U5277 ( .A1(IR_REG_11__SCAN_IN), .A2(keyinput_g66), .B1(
        keyinput_g96), .B2(D_REG_9__SCAN_IN), .ZN(n4737) );
  AOI221_X1 U5278 ( .B1(IR_REG_11__SCAN_IN), .B2(keyinput_g66), .C1(
        D_REG_9__SCAN_IN), .C2(keyinput_g96), .A(n4737), .ZN(n4738) );
  NAND4_X1 U5279 ( .A1(n4741), .A2(n4740), .A3(n4739), .A4(n4738), .ZN(n4754)
         );
  AOI22_X1 U5280 ( .A1(n5058), .A2(keyinput_g54), .B1(n4743), .B2(keyinput_g97), .ZN(n4742) );
  OAI221_X1 U5281 ( .B1(n5058), .B2(keyinput_g54), .C1(n4743), .C2(
        keyinput_g97), .A(n4742), .ZN(n4752) );
  AOI22_X1 U5282 ( .A1(n2545), .A2(keyinput_g122), .B1(keyinput_g42), .B2(
        n2994), .ZN(n4744) );
  OAI221_X1 U5283 ( .B1(n2545), .B2(keyinput_g122), .C1(n2994), .C2(
        keyinput_g42), .A(n4744), .ZN(n4751) );
  AOI22_X1 U5284 ( .A1(n4746), .A2(keyinput_g1), .B1(n2789), .B2(keyinput_g77), 
        .ZN(n4745) );
  OAI221_X1 U5285 ( .B1(n4746), .B2(keyinput_g1), .C1(n2789), .C2(keyinput_g77), .A(n4745), .ZN(n4750) );
  XNOR2_X1 U5286 ( .A(IR_REG_10__SCAN_IN), .B(keyinput_g65), .ZN(n4748) );
  XNOR2_X1 U5287 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_g33), .ZN(n4747) );
  NAND2_X1 U5288 ( .A1(n4748), .A2(n4747), .ZN(n4749) );
  OR4_X1 U5289 ( .A1(n4752), .A2(n4751), .A3(n4750), .A4(n4749), .ZN(n4753) );
  NOR4_X1 U5290 ( .A1(n4756), .A2(n4755), .A3(n4754), .A4(n4753), .ZN(n5083)
         );
  OAI22_X1 U5291 ( .A1(IR_REG_31__SCAN_IN), .A2(keyinput_g86), .B1(
        IR_REG_16__SCAN_IN), .B2(keyinput_g71), .ZN(n4757) );
  AOI221_X1 U5292 ( .B1(IR_REG_31__SCAN_IN), .B2(keyinput_g86), .C1(
        keyinput_g71), .C2(IR_REG_16__SCAN_IN), .A(n4757), .ZN(n4764) );
  OAI22_X1 U5293 ( .A1(IR_REG_15__SCAN_IN), .A2(keyinput_g70), .B1(DATAI_16_), 
        .B2(keyinput_g15), .ZN(n4758) );
  AOI221_X1 U5294 ( .B1(IR_REG_15__SCAN_IN), .B2(keyinput_g70), .C1(
        keyinput_g15), .C2(DATAI_16_), .A(n4758), .ZN(n4763) );
  OAI22_X1 U5295 ( .A1(REG0_REG_0__SCAN_IN), .A2(keyinput_g119), .B1(
        keyinput_g20), .B2(DATAI_11_), .ZN(n4759) );
  AOI221_X1 U5296 ( .B1(REG0_REG_0__SCAN_IN), .B2(keyinput_g119), .C1(
        DATAI_11_), .C2(keyinput_g20), .A(n4759), .ZN(n4762) );
  OAI22_X1 U5297 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(
        keyinput_g125), .B2(REG0_REG_6__SCAN_IN), .ZN(n4760) );
  AOI221_X1 U5298 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(
        REG0_REG_6__SCAN_IN), .C2(keyinput_g125), .A(n4760), .ZN(n4761) );
  NAND4_X1 U5299 ( .A1(n4764), .A2(n4763), .A3(n4762), .A4(n4761), .ZN(n4893)
         );
  OAI22_X1 U5300 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput_g34), .B1(
        keyinput_g3), .B2(DATAI_28_), .ZN(n4765) );
  AOI221_X1 U5301 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput_g34), .C1(
        DATAI_28_), .C2(keyinput_g3), .A(n4765), .ZN(n4791) );
  OAI22_X1 U5302 ( .A1(D_REG_14__SCAN_IN), .A2(keyinput_g101), .B1(
        D_REG_11__SCAN_IN), .B2(keyinput_g98), .ZN(n4766) );
  AOI221_X1 U5303 ( .B1(D_REG_14__SCAN_IN), .B2(keyinput_g101), .C1(
        keyinput_g98), .C2(D_REG_11__SCAN_IN), .A(n4766), .ZN(n4769) );
  OAI22_X1 U5304 ( .A1(REG3_REG_3__SCAN_IN), .A2(keyinput_g38), .B1(
        keyinput_g2), .B2(DATAI_29_), .ZN(n4767) );
  AOI221_X1 U5305 ( .B1(REG3_REG_3__SCAN_IN), .B2(keyinput_g38), .C1(DATAI_29_), .C2(keyinput_g2), .A(n4767), .ZN(n4768) );
  OAI211_X1 U5306 ( .C1(n4771), .C2(keyinput_g103), .A(n4769), .B(n4768), .ZN(
        n4770) );
  AOI21_X1 U5307 ( .B1(n4771), .B2(keyinput_g103), .A(n4770), .ZN(n4790) );
  AOI22_X1 U5308 ( .A1(DATAI_9_), .A2(keyinput_g22), .B1(IR_REG_7__SCAN_IN), 
        .B2(keyinput_g62), .ZN(n4772) );
  OAI221_X1 U5309 ( .B1(DATAI_9_), .B2(keyinput_g22), .C1(IR_REG_7__SCAN_IN), 
        .C2(keyinput_g62), .A(n4772), .ZN(n4779) );
  AOI22_X1 U5310 ( .A1(IR_REG_27__SCAN_IN), .A2(keyinput_g82), .B1(
        IR_REG_20__SCAN_IN), .B2(keyinput_g75), .ZN(n4773) );
  OAI221_X1 U5311 ( .B1(IR_REG_27__SCAN_IN), .B2(keyinput_g82), .C1(
        IR_REG_20__SCAN_IN), .C2(keyinput_g75), .A(n4773), .ZN(n4778) );
  AOI22_X1 U5312 ( .A1(D_REG_30__SCAN_IN), .A2(keyinput_g117), .B1(
        D_REG_3__SCAN_IN), .B2(keyinput_g90), .ZN(n4774) );
  OAI221_X1 U5313 ( .B1(D_REG_30__SCAN_IN), .B2(keyinput_g117), .C1(
        D_REG_3__SCAN_IN), .C2(keyinput_g90), .A(n4774), .ZN(n4777) );
  AOI22_X1 U5314 ( .A1(D_REG_20__SCAN_IN), .A2(keyinput_g107), .B1(
        D_REG_17__SCAN_IN), .B2(keyinput_g104), .ZN(n4775) );
  OAI221_X1 U5315 ( .B1(D_REG_20__SCAN_IN), .B2(keyinput_g107), .C1(
        D_REG_17__SCAN_IN), .C2(keyinput_g104), .A(n4775), .ZN(n4776) );
  NOR4_X1 U5316 ( .A1(n4779), .A2(n4778), .A3(n4777), .A4(n4776), .ZN(n4789)
         );
  AOI22_X1 U5317 ( .A1(D_REG_0__SCAN_IN), .A2(keyinput_g87), .B1(
        D_REG_12__SCAN_IN), .B2(keyinput_g99), .ZN(n4780) );
  OAI221_X1 U5318 ( .B1(D_REG_0__SCAN_IN), .B2(keyinput_g87), .C1(
        D_REG_12__SCAN_IN), .C2(keyinput_g99), .A(n4780), .ZN(n4787) );
  AOI22_X1 U5319 ( .A1(REG3_REG_8__SCAN_IN), .A2(keyinput_g41), .B1(
        IR_REG_8__SCAN_IN), .B2(keyinput_g63), .ZN(n4781) );
  OAI221_X1 U5320 ( .B1(REG3_REG_8__SCAN_IN), .B2(keyinput_g41), .C1(
        IR_REG_8__SCAN_IN), .C2(keyinput_g63), .A(n4781), .ZN(n4786) );
  AOI22_X1 U5321 ( .A1(IR_REG_19__SCAN_IN), .A2(keyinput_g74), .B1(
        IR_REG_24__SCAN_IN), .B2(keyinput_g79), .ZN(n4782) );
  OAI221_X1 U5322 ( .B1(IR_REG_19__SCAN_IN), .B2(keyinput_g74), .C1(
        IR_REG_24__SCAN_IN), .C2(keyinput_g79), .A(n4782), .ZN(n4785) );
  AOI22_X1 U5323 ( .A1(IR_REG_2__SCAN_IN), .A2(keyinput_g57), .B1(
        IR_REG_26__SCAN_IN), .B2(keyinput_g81), .ZN(n4783) );
  OAI221_X1 U5324 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput_g57), .C1(
        IR_REG_26__SCAN_IN), .C2(keyinput_g81), .A(n4783), .ZN(n4784) );
  NOR4_X1 U5325 ( .A1(n4787), .A2(n4786), .A3(n4785), .A4(n4784), .ZN(n4788)
         );
  NAND4_X1 U5326 ( .A1(n4791), .A2(n4790), .A3(n4789), .A4(n4788), .ZN(n4892)
         );
  AOI22_X1 U5327 ( .A1(n5057), .A2(keyinput_g17), .B1(n2499), .B2(keyinput_g6), 
        .ZN(n4792) );
  OAI221_X1 U5328 ( .B1(n5057), .B2(keyinput_g17), .C1(n2499), .C2(keyinput_g6), .A(n4792), .ZN(n4800) );
  AOI22_X1 U5329 ( .A1(n5055), .A2(keyinput_g25), .B1(n4976), .B2(keyinput_g53), .ZN(n4793) );
  OAI221_X1 U5330 ( .B1(n5055), .B2(keyinput_g25), .C1(n4976), .C2(
        keyinput_g53), .A(n4793), .ZN(n4799) );
  AOI22_X1 U5331 ( .A1(n4795), .A2(keyinput_g111), .B1(keyinput_g43), .B2(
        n2735), .ZN(n4794) );
  OAI221_X1 U5332 ( .B1(n4795), .B2(keyinput_g111), .C1(n2735), .C2(
        keyinput_g43), .A(n4794), .ZN(n4798) );
  AOI22_X1 U5333 ( .A1(n2528), .A2(keyinput_g31), .B1(n5030), .B2(keyinput_g89), .ZN(n4796) );
  OAI221_X1 U5334 ( .B1(n2528), .B2(keyinput_g31), .C1(n5030), .C2(
        keyinput_g89), .A(n4796), .ZN(n4797) );
  NOR4_X1 U5335 ( .A1(n4800), .A2(n4799), .A3(n4798), .A4(n4797), .ZN(n4837)
         );
  AOI22_X1 U5336 ( .A1(n4802), .A2(keyinput_g24), .B1(keyinput_g0), .B2(n4975), 
        .ZN(n4801) );
  OAI221_X1 U5337 ( .B1(n4802), .B2(keyinput_g24), .C1(n4975), .C2(keyinput_g0), .A(n4801), .ZN(n4812) );
  AOI22_X1 U5338 ( .A1(n4805), .A2(keyinput_g105), .B1(keyinput_g26), .B2(
        n4804), .ZN(n4803) );
  OAI221_X1 U5339 ( .B1(n4805), .B2(keyinput_g105), .C1(n4804), .C2(
        keyinput_g26), .A(n4803), .ZN(n4811) );
  AOI22_X1 U5340 ( .A1(n5031), .A2(keyinput_g113), .B1(n5036), .B2(
        keyinput_g114), .ZN(n4806) );
  OAI221_X1 U5341 ( .B1(n5031), .B2(keyinput_g113), .C1(n5036), .C2(
        keyinput_g114), .A(n4806), .ZN(n4810) );
  XOR2_X1 U5342 ( .A(n3560), .B(keyinput_g40), .Z(n4808) );
  XNOR2_X1 U5343 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_g60), .ZN(n4807) );
  NAND2_X1 U5344 ( .A1(n4808), .A2(n4807), .ZN(n4809) );
  NOR4_X1 U5345 ( .A1(n4812), .A2(n4811), .A3(n4810), .A4(n4809), .ZN(n4836)
         );
  AOI22_X1 U5346 ( .A1(n3597), .A2(keyinput_g45), .B1(keyinput_g51), .B2(n2610), .ZN(n4813) );
  OAI221_X1 U5347 ( .B1(n3597), .B2(keyinput_g45), .C1(n2610), .C2(
        keyinput_g51), .A(n4813), .ZN(n4822) );
  AOI22_X1 U5348 ( .A1(n2559), .A2(keyinput_g58), .B1(keyinput_g18), .B2(n5002), .ZN(n4814) );
  OAI221_X1 U5349 ( .B1(n2559), .B2(keyinput_g58), .C1(n5002), .C2(
        keyinput_g18), .A(n4814), .ZN(n4821) );
  INV_X1 U5350 ( .A(DATAI_2_), .ZN(n4816) );
  AOI22_X1 U5351 ( .A1(n4816), .A2(keyinput_g29), .B1(n5034), .B2(
        keyinput_g110), .ZN(n4815) );
  OAI221_X1 U5352 ( .B1(n4816), .B2(keyinput_g29), .C1(n5034), .C2(
        keyinput_g110), .A(n4815), .ZN(n4820) );
  XNOR2_X1 U5353 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_g76), .ZN(n4818) );
  XNOR2_X1 U5354 ( .A(DATAI_4_), .B(keyinput_g27), .ZN(n4817) );
  NAND2_X1 U5355 ( .A1(n4818), .A2(n4817), .ZN(n4819) );
  NOR4_X1 U5356 ( .A1(n4822), .A2(n4821), .A3(n4820), .A4(n4819), .ZN(n4835)
         );
  INV_X1 U5357 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4824) );
  AOI22_X1 U5358 ( .A1(n4824), .A2(keyinput_g121), .B1(keyinput_g52), .B2(
        n3010), .ZN(n4823) );
  OAI221_X1 U5359 ( .B1(n4824), .B2(keyinput_g121), .C1(n3010), .C2(
        keyinput_g52), .A(n4823), .ZN(n4833) );
  AOI22_X1 U5360 ( .A1(n4826), .A2(keyinput_g36), .B1(n2394), .B2(keyinput_g56), .ZN(n4825) );
  OAI221_X1 U5361 ( .B1(n4826), .B2(keyinput_g36), .C1(n2394), .C2(
        keyinput_g56), .A(n4825), .ZN(n4832) );
  AOI22_X1 U5362 ( .A1(n2743), .A2(keyinput_g10), .B1(n4828), .B2(
        keyinput_g115), .ZN(n4827) );
  OAI221_X1 U5363 ( .B1(n2743), .B2(keyinput_g10), .C1(n4828), .C2(
        keyinput_g115), .A(n4827), .ZN(n4831) );
  AOI22_X1 U5364 ( .A1(n5043), .A2(keyinput_g14), .B1(keyinput_g123), .B2(
        n2552), .ZN(n4829) );
  OAI221_X1 U5365 ( .B1(n5043), .B2(keyinput_g14), .C1(n2552), .C2(
        keyinput_g123), .A(n4829), .ZN(n4830) );
  NOR4_X1 U5366 ( .A1(n4833), .A2(n4832), .A3(n4831), .A4(n4830), .ZN(n4834)
         );
  NAND4_X1 U5367 ( .A1(n4837), .A2(n4836), .A3(n4835), .A4(n4834), .ZN(n4891)
         );
  AOI22_X1 U5368 ( .A1(n4840), .A2(keyinput_g116), .B1(keyinput_g49), .B2(
        n4839), .ZN(n4838) );
  OAI221_X1 U5369 ( .B1(n4840), .B2(keyinput_g116), .C1(n4839), .C2(
        keyinput_g49), .A(n4838), .ZN(n4850) );
  AOI22_X1 U5370 ( .A1(n4988), .A2(keyinput_g50), .B1(n4842), .B2(keyinput_g91), .ZN(n4841) );
  OAI221_X1 U5371 ( .B1(n4988), .B2(keyinput_g50), .C1(n4842), .C2(
        keyinput_g91), .A(n4841), .ZN(n4849) );
  AOI22_X1 U5372 ( .A1(n4845), .A2(keyinput_g108), .B1(keyinput_g109), .B2(
        n4844), .ZN(n4843) );
  OAI221_X1 U5373 ( .B1(n4845), .B2(keyinput_g108), .C1(n4844), .C2(
        keyinput_g109), .A(n4843), .ZN(n4848) );
  AOI22_X1 U5374 ( .A1(n5045), .A2(keyinput_g37), .B1(n5018), .B2(
        keyinput_g100), .ZN(n4846) );
  OAI221_X1 U5375 ( .B1(n5045), .B2(keyinput_g37), .C1(n5018), .C2(
        keyinput_g100), .A(n4846), .ZN(n4847) );
  NOR4_X1 U5376 ( .A1(n4850), .A2(n4849), .A3(n4848), .A4(n4847), .ZN(n4889)
         );
  AOI22_X1 U5377 ( .A1(n4852), .A2(keyinput_g12), .B1(n4997), .B2(
        keyinput_g118), .ZN(n4851) );
  OAI221_X1 U5378 ( .B1(n4852), .B2(keyinput_g12), .C1(n4997), .C2(
        keyinput_g118), .A(n4851), .ZN(n4858) );
  INV_X1 U5379 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4854) );
  AOI22_X1 U5380 ( .A1(n4855), .A2(keyinput_g13), .B1(n4854), .B2(keyinput_g44), .ZN(n4853) );
  OAI221_X1 U5381 ( .B1(n4855), .B2(keyinput_g13), .C1(n4854), .C2(
        keyinput_g44), .A(n4853), .ZN(n4857) );
  XOR2_X1 U5382 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_g73), .Z(n4856) );
  OR3_X1 U5383 ( .A1(n4858), .A2(n4857), .A3(n4856), .ZN(n4863) );
  AOI22_X1 U5384 ( .A1(n4860), .A2(keyinput_g23), .B1(keyinput_g120), .B2(
        n2529), .ZN(n4859) );
  OAI221_X1 U5385 ( .B1(n4860), .B2(keyinput_g23), .C1(n2529), .C2(
        keyinput_g120), .A(n4859), .ZN(n4862) );
  XNOR2_X1 U5386 ( .A(n5014), .B(keyinput_g106), .ZN(n4861) );
  NOR3_X1 U5387 ( .A1(n4863), .A2(n4862), .A3(n4861), .ZN(n4888) );
  AOI22_X1 U5388 ( .A1(n2399), .A2(keyinput_g30), .B1(n2928), .B2(keyinput_g55), .ZN(n4864) );
  OAI221_X1 U5389 ( .B1(n2399), .B2(keyinput_g30), .C1(n2928), .C2(
        keyinput_g55), .A(n4864), .ZN(n4873) );
  AOI22_X1 U5390 ( .A1(n2698), .A2(keyinput_g48), .B1(n5021), .B2(keyinput_g92), .ZN(n4865) );
  OAI221_X1 U5391 ( .B1(n2698), .B2(keyinput_g48), .C1(n5021), .C2(
        keyinput_g92), .A(n4865), .ZN(n4872) );
  AOI22_X1 U5392 ( .A1(n2773), .A2(keyinput_g4), .B1(n4867), .B2(keyinput_g47), 
        .ZN(n4866) );
  OAI221_X1 U5393 ( .B1(n2773), .B2(keyinput_g4), .C1(n4867), .C2(keyinput_g47), .A(n4866), .ZN(n4871) );
  XNOR2_X1 U5394 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_g83), .ZN(n4869) );
  XNOR2_X1 U5395 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_g64), .ZN(n4868) );
  NAND2_X1 U5396 ( .A1(n4869), .A2(n4868), .ZN(n4870) );
  NOR4_X1 U5397 ( .A1(n4873), .A2(n4872), .A3(n4871), .A4(n4870), .ZN(n4887)
         );
  INV_X1 U5398 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4985) );
  AOI22_X1 U5399 ( .A1(n4985), .A2(keyinput_g124), .B1(n4875), .B2(
        keyinput_g112), .ZN(n4874) );
  OAI221_X1 U5400 ( .B1(n4985), .B2(keyinput_g124), .C1(n4875), .C2(
        keyinput_g112), .A(n4874), .ZN(n4885) );
  AOI22_X1 U5401 ( .A1(n5017), .A2(keyinput_g94), .B1(keyinput_g32), .B2(U3149), .ZN(n4876) );
  OAI221_X1 U5402 ( .B1(n5017), .B2(keyinput_g94), .C1(U3149), .C2(
        keyinput_g32), .A(n4876), .ZN(n4884) );
  AOI22_X1 U5403 ( .A1(n4879), .A2(keyinput_g5), .B1(n4878), .B2(keyinput_g19), 
        .ZN(n4877) );
  OAI221_X1 U5404 ( .B1(n4879), .B2(keyinput_g5), .C1(n4878), .C2(keyinput_g19), .A(n4877), .ZN(n4883) );
  XOR2_X1 U5405 ( .A(n2753), .B(keyinput_g8), .Z(n4881) );
  XNOR2_X1 U5406 ( .A(IR_REG_23__SCAN_IN), .B(keyinput_g78), .ZN(n4880) );
  NAND2_X1 U5407 ( .A1(n4881), .A2(n4880), .ZN(n4882) );
  NOR4_X1 U5408 ( .A1(n4885), .A2(n4884), .A3(n4883), .A4(n4882), .ZN(n4886)
         );
  NAND4_X1 U5409 ( .A1(n4889), .A2(n4888), .A3(n4887), .A4(n4886), .ZN(n4890)
         );
  NOR4_X1 U5410 ( .A1(n4893), .A2(n4892), .A3(n4891), .A4(n4890), .ZN(n5082)
         );
  INV_X1 U5411 ( .A(DATAI_3_), .ZN(n5080) );
  OAI22_X1 U5412 ( .A1(IR_REG_7__SCAN_IN), .A2(keyinput_f62), .B1(keyinput_f33), .B2(REG3_REG_7__SCAN_IN), .ZN(n4894) );
  AOI221_X1 U5413 ( .B1(IR_REG_7__SCAN_IN), .B2(keyinput_f62), .C1(
        REG3_REG_7__SCAN_IN), .C2(keyinput_f33), .A(n4894), .ZN(n4901) );
  OAI22_X1 U5414 ( .A1(IR_REG_12__SCAN_IN), .A2(keyinput_f67), .B1(
        keyinput_f51), .B2(REG3_REG_9__SCAN_IN), .ZN(n4895) );
  AOI221_X1 U5415 ( .B1(IR_REG_12__SCAN_IN), .B2(keyinput_f67), .C1(
        REG3_REG_9__SCAN_IN), .C2(keyinput_f51), .A(n4895), .ZN(n4900) );
  OAI22_X1 U5416 ( .A1(IR_REG_13__SCAN_IN), .A2(keyinput_f68), .B1(
        IR_REG_27__SCAN_IN), .B2(keyinput_f82), .ZN(n4896) );
  AOI221_X1 U5417 ( .B1(IR_REG_13__SCAN_IN), .B2(keyinput_f68), .C1(
        keyinput_f82), .C2(IR_REG_27__SCAN_IN), .A(n4896), .ZN(n4899) );
  OAI22_X1 U5418 ( .A1(IR_REG_20__SCAN_IN), .A2(keyinput_f75), .B1(
        keyinput_f88), .B2(D_REG_1__SCAN_IN), .ZN(n4897) );
  AOI221_X1 U5419 ( .B1(IR_REG_20__SCAN_IN), .B2(keyinput_f75), .C1(
        D_REG_1__SCAN_IN), .C2(keyinput_f88), .A(n4897), .ZN(n4898) );
  NAND4_X1 U5420 ( .A1(n4901), .A2(n4900), .A3(n4899), .A4(n4898), .ZN(n4929)
         );
  OAI22_X1 U5421 ( .A1(IR_REG_18__SCAN_IN), .A2(keyinput_f73), .B1(
        D_REG_28__SCAN_IN), .B2(keyinput_f115), .ZN(n4902) );
  AOI221_X1 U5422 ( .B1(IR_REG_18__SCAN_IN), .B2(keyinput_f73), .C1(
        keyinput_f115), .C2(D_REG_28__SCAN_IN), .A(n4902), .ZN(n4909) );
  OAI22_X1 U5423 ( .A1(D_REG_24__SCAN_IN), .A2(keyinput_f111), .B1(
        D_REG_10__SCAN_IN), .B2(keyinput_f97), .ZN(n4903) );
  AOI221_X1 U5424 ( .B1(D_REG_24__SCAN_IN), .B2(keyinput_f111), .C1(
        keyinput_f97), .C2(D_REG_10__SCAN_IN), .A(n4903), .ZN(n4908) );
  OAI22_X1 U5425 ( .A1(D_REG_25__SCAN_IN), .A2(keyinput_f112), .B1(
        D_REG_16__SCAN_IN), .B2(keyinput_f103), .ZN(n4904) );
  AOI221_X1 U5426 ( .B1(D_REG_25__SCAN_IN), .B2(keyinput_f112), .C1(
        keyinput_f103), .C2(D_REG_16__SCAN_IN), .A(n4904), .ZN(n4907) );
  OAI22_X1 U5427 ( .A1(D_REG_18__SCAN_IN), .A2(keyinput_f105), .B1(
        D_REG_29__SCAN_IN), .B2(keyinput_f116), .ZN(n4905) );
  AOI221_X1 U5428 ( .B1(D_REG_18__SCAN_IN), .B2(keyinput_f105), .C1(
        keyinput_f116), .C2(D_REG_29__SCAN_IN), .A(n4905), .ZN(n4906) );
  NAND4_X1 U5429 ( .A1(n4909), .A2(n4908), .A3(n4907), .A4(n4906), .ZN(n4928)
         );
  OAI22_X1 U5430 ( .A1(D_REG_4__SCAN_IN), .A2(keyinput_f91), .B1(
        D_REG_21__SCAN_IN), .B2(keyinput_f108), .ZN(n4910) );
  AOI221_X1 U5431 ( .B1(D_REG_4__SCAN_IN), .B2(keyinput_f91), .C1(
        keyinput_f108), .C2(D_REG_21__SCAN_IN), .A(n4910), .ZN(n4917) );
  OAI22_X1 U5432 ( .A1(D_REG_22__SCAN_IN), .A2(keyinput_f109), .B1(
        D_REG_0__SCAN_IN), .B2(keyinput_f87), .ZN(n4911) );
  AOI221_X1 U5433 ( .B1(D_REG_22__SCAN_IN), .B2(keyinput_f109), .C1(
        keyinput_f87), .C2(D_REG_0__SCAN_IN), .A(n4911), .ZN(n4916) );
  OAI22_X1 U5434 ( .A1(REG3_REG_25__SCAN_IN), .A2(keyinput_f45), .B1(
        keyinput_f48), .B2(REG3_REG_17__SCAN_IN), .ZN(n4912) );
  AOI221_X1 U5435 ( .B1(REG3_REG_25__SCAN_IN), .B2(keyinput_f45), .C1(
        REG3_REG_17__SCAN_IN), .C2(keyinput_f48), .A(n4912), .ZN(n4915) );
  OAI22_X1 U5436 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput_f46), .B1(
        REG3_REG_8__SCAN_IN), .B2(keyinput_f41), .ZN(n4913) );
  AOI221_X1 U5437 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput_f46), .C1(
        keyinput_f41), .C2(REG3_REG_8__SCAN_IN), .A(n4913), .ZN(n4914) );
  NAND4_X1 U5438 ( .A1(n4917), .A2(n4916), .A3(n4915), .A4(n4914), .ZN(n4927)
         );
  OAI22_X1 U5439 ( .A1(DATAI_12_), .A2(keyinput_f19), .B1(keyinput_f31), .B2(
        DATAI_0_), .ZN(n4918) );
  AOI221_X1 U5440 ( .B1(DATAI_12_), .B2(keyinput_f19), .C1(DATAI_0_), .C2(
        keyinput_f31), .A(n4918), .ZN(n4925) );
  OAI22_X1 U5441 ( .A1(IR_REG_23__SCAN_IN), .A2(keyinput_f78), .B1(
        REG0_REG_2__SCAN_IN), .B2(keyinput_f121), .ZN(n4919) );
  AOI221_X1 U5442 ( .B1(IR_REG_23__SCAN_IN), .B2(keyinput_f78), .C1(
        keyinput_f121), .C2(REG0_REG_2__SCAN_IN), .A(n4919), .ZN(n4924) );
  OAI22_X1 U5443 ( .A1(IR_REG_5__SCAN_IN), .A2(keyinput_f60), .B1(keyinput_f29), .B2(DATAI_2_), .ZN(n4920) );
  AOI221_X1 U5444 ( .B1(IR_REG_5__SCAN_IN), .B2(keyinput_f60), .C1(DATAI_2_), 
        .C2(keyinput_f29), .A(n4920), .ZN(n4923) );
  OAI22_X1 U5445 ( .A1(DATAI_5_), .A2(keyinput_f26), .B1(DATAI_30_), .B2(
        keyinput_f1), .ZN(n4921) );
  AOI221_X1 U5446 ( .B1(DATAI_5_), .B2(keyinput_f26), .C1(keyinput_f1), .C2(
        DATAI_30_), .A(n4921), .ZN(n4922) );
  NAND4_X1 U5447 ( .A1(n4925), .A2(n4924), .A3(n4923), .A4(n4922), .ZN(n4926)
         );
  NOR4_X1 U5448 ( .A1(n4929), .A2(n4928), .A3(n4927), .A4(n4926), .ZN(n5075)
         );
  OAI22_X1 U5449 ( .A1(REG3_REG_24__SCAN_IN), .A2(keyinput_f49), .B1(
        REG3_REG_3__SCAN_IN), .B2(keyinput_f38), .ZN(n4930) );
  AOI221_X1 U5450 ( .B1(REG3_REG_24__SCAN_IN), .B2(keyinput_f49), .C1(
        keyinput_f38), .C2(REG3_REG_3__SCAN_IN), .A(n4930), .ZN(n4937) );
  OAI22_X1 U5451 ( .A1(REG3_REG_14__SCAN_IN), .A2(keyinput_f35), .B1(
        keyinput_f42), .B2(REG3_REG_1__SCAN_IN), .ZN(n4931) );
  AOI221_X1 U5452 ( .B1(REG3_REG_14__SCAN_IN), .B2(keyinput_f35), .C1(
        REG3_REG_1__SCAN_IN), .C2(keyinput_f42), .A(n4931), .ZN(n4936) );
  OAI22_X1 U5453 ( .A1(D_REG_15__SCAN_IN), .A2(keyinput_f102), .B1(
        keyinput_f16), .B2(DATAI_15_), .ZN(n4932) );
  AOI221_X1 U5454 ( .B1(D_REG_15__SCAN_IN), .B2(keyinput_f102), .C1(DATAI_15_), 
        .C2(keyinput_f16), .A(n4932), .ZN(n4935) );
  OAI22_X1 U5455 ( .A1(D_REG_14__SCAN_IN), .A2(keyinput_f101), .B1(
        D_REG_11__SCAN_IN), .B2(keyinput_f98), .ZN(n4933) );
  AOI221_X1 U5456 ( .B1(D_REG_14__SCAN_IN), .B2(keyinput_f101), .C1(
        keyinput_f98), .C2(D_REG_11__SCAN_IN), .A(n4933), .ZN(n4934) );
  NAND4_X1 U5457 ( .A1(n4937), .A2(n4936), .A3(n4935), .A4(n4934), .ZN(n5073)
         );
  AOI22_X1 U5458 ( .A1(D_REG_8__SCAN_IN), .A2(keyinput_f95), .B1(
        D_REG_9__SCAN_IN), .B2(keyinput_f96), .ZN(n4938) );
  OAI221_X1 U5459 ( .B1(D_REG_8__SCAN_IN), .B2(keyinput_f95), .C1(
        D_REG_9__SCAN_IN), .C2(keyinput_f96), .A(n4938), .ZN(n4945) );
  AOI22_X1 U5460 ( .A1(IR_REG_30__SCAN_IN), .A2(keyinput_f85), .B1(
        IR_REG_17__SCAN_IN), .B2(keyinput_f72), .ZN(n4939) );
  OAI221_X1 U5461 ( .B1(IR_REG_30__SCAN_IN), .B2(keyinput_f85), .C1(
        IR_REG_17__SCAN_IN), .C2(keyinput_f72), .A(n4939), .ZN(n4944) );
  AOI22_X1 U5462 ( .A1(IR_REG_15__SCAN_IN), .A2(keyinput_f70), .B1(
        IR_REG_16__SCAN_IN), .B2(keyinput_f71), .ZN(n4940) );
  OAI221_X1 U5463 ( .B1(IR_REG_15__SCAN_IN), .B2(keyinput_f70), .C1(
        IR_REG_16__SCAN_IN), .C2(keyinput_f71), .A(n4940), .ZN(n4943) );
  AOI22_X1 U5464 ( .A1(DATAI_11_), .A2(keyinput_f20), .B1(DATAI_16_), .B2(
        keyinput_f15), .ZN(n4941) );
  OAI221_X1 U5465 ( .B1(DATAI_11_), .B2(keyinput_f20), .C1(DATAI_16_), .C2(
        keyinput_f15), .A(n4941), .ZN(n4942) );
  NOR4_X1 U5466 ( .A1(n4945), .A2(n4944), .A3(n4943), .A4(n4942), .ZN(n4963)
         );
  AOI22_X1 U5467 ( .A1(REG0_REG_3__SCAN_IN), .A2(keyinput_f122), .B1(
        REG0_REG_8__SCAN_IN), .B2(keyinput_f127), .ZN(n4946) );
  OAI221_X1 U5468 ( .B1(REG0_REG_3__SCAN_IN), .B2(keyinput_f122), .C1(
        REG0_REG_8__SCAN_IN), .C2(keyinput_f127), .A(n4946), .ZN(n4953) );
  AOI22_X1 U5469 ( .A1(REG0_REG_4__SCAN_IN), .A2(keyinput_f123), .B1(
        REG0_REG_1__SCAN_IN), .B2(keyinput_f120), .ZN(n4947) );
  OAI221_X1 U5470 ( .B1(REG0_REG_4__SCAN_IN), .B2(keyinput_f123), .C1(
        REG0_REG_1__SCAN_IN), .C2(keyinput_f120), .A(n4947), .ZN(n4952) );
  AOI22_X1 U5471 ( .A1(IR_REG_3__SCAN_IN), .A2(keyinput_f58), .B1(
        IR_REG_4__SCAN_IN), .B2(keyinput_f59), .ZN(n4948) );
  OAI221_X1 U5472 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput_f58), .C1(
        IR_REG_4__SCAN_IN), .C2(keyinput_f59), .A(n4948), .ZN(n4951) );
  AOI22_X1 U5473 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput_f47), .B1(
        IR_REG_6__SCAN_IN), .B2(keyinput_f61), .ZN(n4949) );
  OAI221_X1 U5474 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput_f47), .C1(
        IR_REG_6__SCAN_IN), .C2(keyinput_f61), .A(n4949), .ZN(n4950) );
  NOR4_X1 U5475 ( .A1(n4953), .A2(n4952), .A3(n4951), .A4(n4950), .ZN(n4962)
         );
  OAI22_X1 U5476 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput_f34), .B1(
        REG3_REG_21__SCAN_IN), .B2(keyinput_f43), .ZN(n4954) );
  AOI221_X1 U5477 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput_f34), .C1(
        keyinput_f43), .C2(REG3_REG_21__SCAN_IN), .A(n4954), .ZN(n4960) );
  OAI22_X1 U5478 ( .A1(STATE_REG_SCAN_IN), .A2(keyinput_f32), .B1(DATAI_22_), 
        .B2(keyinput_f9), .ZN(n4955) );
  AOI221_X1 U5479 ( .B1(STATE_REG_SCAN_IN), .B2(keyinput_f32), .C1(keyinput_f9), .C2(DATAI_22_), .A(n4955), .ZN(n4959) );
  OAI22_X1 U5480 ( .A1(DATAI_28_), .A2(keyinput_f3), .B1(DATAI_24_), .B2(
        keyinput_f7), .ZN(n4956) );
  AOI221_X1 U5481 ( .B1(DATAI_28_), .B2(keyinput_f3), .C1(keyinput_f7), .C2(
        DATAI_24_), .A(n4956), .ZN(n4958) );
  XNOR2_X1 U5482 ( .A(IR_REG_10__SCAN_IN), .B(keyinput_f65), .ZN(n4957) );
  AND4_X1 U5483 ( .A1(n4960), .A2(n4959), .A3(n4958), .A4(n4957), .ZN(n4961)
         );
  NAND3_X1 U5484 ( .A1(n4963), .A2(n4962), .A3(n4961), .ZN(n5072) );
  AOI22_X1 U5485 ( .A1(DATAI_25_), .A2(keyinput_f6), .B1(IR_REG_22__SCAN_IN), 
        .B2(keyinput_f77), .ZN(n4964) );
  OAI221_X1 U5486 ( .B1(DATAI_25_), .B2(keyinput_f6), .C1(IR_REG_22__SCAN_IN), 
        .C2(keyinput_f77), .A(n4964), .ZN(n4971) );
  AOI22_X1 U5487 ( .A1(DATAI_19_), .A2(keyinput_f12), .B1(IR_REG_25__SCAN_IN), 
        .B2(keyinput_f80), .ZN(n4965) );
  OAI221_X1 U5488 ( .B1(DATAI_19_), .B2(keyinput_f12), .C1(IR_REG_25__SCAN_IN), 
        .C2(keyinput_f80), .A(n4965), .ZN(n4970) );
  AOI22_X1 U5489 ( .A1(DATAI_18_), .A2(keyinput_f13), .B1(REG3_REG_12__SCAN_IN), .B2(keyinput_f44), .ZN(n4966) );
  OAI221_X1 U5490 ( .B1(DATAI_18_), .B2(keyinput_f13), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput_f44), .A(n4966), .ZN(n4969) );
  AOI22_X1 U5491 ( .A1(DATAI_1_), .A2(keyinput_f30), .B1(DATAI_8_), .B2(
        keyinput_f23), .ZN(n4967) );
  OAI221_X1 U5492 ( .B1(DATAI_1_), .B2(keyinput_f30), .C1(DATAI_8_), .C2(
        keyinput_f23), .A(n4967), .ZN(n4968) );
  NOR4_X1 U5493 ( .A1(n4971), .A2(n4970), .A3(n4969), .A4(n4968), .ZN(n5012)
         );
  AOI22_X1 U5494 ( .A1(DATAI_26_), .A2(keyinput_f5), .B1(IR_REG_9__SCAN_IN), 
        .B2(keyinput_f64), .ZN(n4972) );
  OAI221_X1 U5495 ( .B1(DATAI_26_), .B2(keyinput_f5), .C1(IR_REG_9__SCAN_IN), 
        .C2(keyinput_f64), .A(n4972), .ZN(n4983) );
  AOI22_X1 U5496 ( .A1(n3010), .A2(keyinput_f52), .B1(n3560), .B2(keyinput_f40), .ZN(n4973) );
  OAI221_X1 U5497 ( .B1(n3010), .B2(keyinput_f52), .C1(n3560), .C2(
        keyinput_f40), .A(n4973), .ZN(n4982) );
  AOI22_X1 U5498 ( .A1(n4976), .A2(keyinput_f53), .B1(keyinput_f0), .B2(n4975), 
        .ZN(n4974) );
  OAI221_X1 U5499 ( .B1(n4976), .B2(keyinput_f53), .C1(n4975), .C2(keyinput_f0), .A(n4974), .ZN(n4981) );
  AOI22_X1 U5500 ( .A1(n4979), .A2(keyinput_f2), .B1(keyinput_f11), .B2(n4978), 
        .ZN(n4977) );
  OAI221_X1 U5501 ( .B1(n4979), .B2(keyinput_f2), .C1(n4978), .C2(keyinput_f11), .A(n4977), .ZN(n4980) );
  NOR4_X1 U5502 ( .A1(n4983), .A2(n4982), .A3(n4981), .A4(n4980), .ZN(n5011)
         );
  INV_X1 U5503 ( .A(DATAI_4_), .ZN(n4986) );
  AOI22_X1 U5504 ( .A1(n4986), .A2(keyinput_f27), .B1(n4985), .B2(
        keyinput_f124), .ZN(n4984) );
  OAI221_X1 U5505 ( .B1(n4986), .B2(keyinput_f27), .C1(n4985), .C2(
        keyinput_f124), .A(n4984), .ZN(n4995) );
  AOI22_X1 U5506 ( .A1(n2394), .A2(keyinput_f56), .B1(keyinput_f50), .B2(n4988), .ZN(n4987) );
  OAI221_X1 U5507 ( .B1(n2394), .B2(keyinput_f56), .C1(n4988), .C2(
        keyinput_f50), .A(n4987), .ZN(n4994) );
  XOR2_X1 U5508 ( .A(n2523), .B(keyinput_f119), .Z(n4992) );
  XNOR2_X1 U5509 ( .A(keyinput_f55), .B(IR_REG_0__SCAN_IN), .ZN(n4991) );
  XNOR2_X1 U5510 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_f86), .ZN(n4990) );
  XNOR2_X1 U5511 ( .A(IR_REG_14__SCAN_IN), .B(keyinput_f69), .ZN(n4989) );
  NAND4_X1 U5512 ( .A1(n4992), .A2(n4991), .A3(n4990), .A4(n4989), .ZN(n4993)
         );
  NOR3_X1 U5513 ( .A1(n4995), .A2(n4994), .A3(n4993), .ZN(n5010) );
  AOI22_X1 U5514 ( .A1(n4998), .A2(keyinput_f90), .B1(keyinput_f118), .B2(
        n4997), .ZN(n4996) );
  OAI221_X1 U5515 ( .B1(n4998), .B2(keyinput_f90), .C1(n4997), .C2(
        keyinput_f118), .A(n4996), .ZN(n5008) );
  AOI22_X1 U5516 ( .A1(n2576), .A2(keyinput_f125), .B1(keyinput_f126), .B2(
        n2586), .ZN(n4999) );
  OAI221_X1 U5517 ( .B1(n2576), .B2(keyinput_f125), .C1(n2586), .C2(
        keyinput_f126), .A(n4999), .ZN(n5007) );
  AOI22_X1 U5518 ( .A1(n5001), .A2(keyinput_f22), .B1(n2651), .B2(keyinput_f66), .ZN(n5000) );
  OAI221_X1 U5519 ( .B1(n5001), .B2(keyinput_f22), .C1(n2651), .C2(
        keyinput_f66), .A(n5000), .ZN(n5006) );
  XOR2_X1 U5520 ( .A(n5002), .B(keyinput_f18), .Z(n5004) );
  XNOR2_X1 U5521 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_f83), .ZN(n5003) );
  NAND2_X1 U5522 ( .A1(n5004), .A2(n5003), .ZN(n5005) );
  NOR4_X1 U5523 ( .A1(n5008), .A2(n5007), .A3(n5006), .A4(n5005), .ZN(n5009)
         );
  NAND4_X1 U5524 ( .A1(n5012), .A2(n5011), .A3(n5010), .A4(n5009), .ZN(n5071)
         );
  AOI22_X1 U5525 ( .A1(n5015), .A2(keyinput_f93), .B1(keyinput_f106), .B2(
        n5014), .ZN(n5013) );
  OAI221_X1 U5526 ( .B1(n5015), .B2(keyinput_f93), .C1(n5014), .C2(
        keyinput_f106), .A(n5013), .ZN(n5028) );
  AOI22_X1 U5527 ( .A1(n5018), .A2(keyinput_f100), .B1(keyinput_f94), .B2(
        n5017), .ZN(n5016) );
  OAI221_X1 U5528 ( .B1(n5018), .B2(keyinput_f100), .C1(n5017), .C2(
        keyinput_f94), .A(n5016), .ZN(n5027) );
  AOI22_X1 U5529 ( .A1(n5021), .A2(keyinput_f92), .B1(keyinput_f117), .B2(
        n5020), .ZN(n5019) );
  OAI221_X1 U5530 ( .B1(n5021), .B2(keyinput_f92), .C1(n5020), .C2(
        keyinput_f117), .A(n5019), .ZN(n5026) );
  AOI22_X1 U5531 ( .A1(n5024), .A2(keyinput_f104), .B1(keyinput_f107), .B2(
        n5023), .ZN(n5022) );
  OAI221_X1 U5532 ( .B1(n5024), .B2(keyinput_f104), .C1(n5023), .C2(
        keyinput_f107), .A(n5022), .ZN(n5025) );
  NOR4_X1 U5533 ( .A1(n5028), .A2(n5027), .A3(n5026), .A4(n5025), .ZN(n5069)
         );
  AOI22_X1 U5534 ( .A1(n5031), .A2(keyinput_f113), .B1(keyinput_f89), .B2(
        n5030), .ZN(n5029) );
  OAI221_X1 U5535 ( .B1(n5031), .B2(keyinput_f113), .C1(n5030), .C2(
        keyinput_f89), .A(n5029), .ZN(n5041) );
  AOI22_X1 U5536 ( .A1(n5034), .A2(keyinput_f110), .B1(n5033), .B2(
        keyinput_f99), .ZN(n5032) );
  OAI221_X1 U5537 ( .B1(n5034), .B2(keyinput_f110), .C1(n5033), .C2(
        keyinput_f99), .A(n5032), .ZN(n5040) );
  AOI22_X1 U5538 ( .A1(n5036), .A2(keyinput_f114), .B1(keyinput_f84), .B2(
        n2473), .ZN(n5035) );
  OAI221_X1 U5539 ( .B1(n5036), .B2(keyinput_f114), .C1(n2473), .C2(
        keyinput_f84), .A(n5035), .ZN(n5039) );
  AOI22_X1 U5540 ( .A1(n2753), .A2(keyinput_f8), .B1(n2773), .B2(keyinput_f4), 
        .ZN(n5037) );
  OAI221_X1 U5541 ( .B1(n2753), .B2(keyinput_f8), .C1(n2773), .C2(keyinput_f4), 
        .A(n5037), .ZN(n5038) );
  NOR4_X1 U5542 ( .A1(n5041), .A2(n5040), .A3(n5039), .A4(n5038), .ZN(n5068)
         );
  AOI22_X1 U5543 ( .A1(n5043), .A2(keyinput_f14), .B1(n2743), .B2(keyinput_f10), .ZN(n5042) );
  OAI221_X1 U5544 ( .B1(n5043), .B2(keyinput_f14), .C1(n2743), .C2(
        keyinput_f10), .A(n5042), .ZN(n5053) );
  AOI22_X1 U5545 ( .A1(n5046), .A2(keyinput_f21), .B1(n5045), .B2(keyinput_f37), .ZN(n5044) );
  OAI221_X1 U5546 ( .B1(n5046), .B2(keyinput_f21), .C1(n5045), .C2(
        keyinput_f37), .A(n5044), .ZN(n5052) );
  XNOR2_X1 U5547 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_f39), .ZN(n5050) );
  XNOR2_X1 U5548 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_f79), .ZN(n5049) );
  XNOR2_X1 U5549 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_f76), .ZN(n5048) );
  XNOR2_X1 U5550 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput_f36), .ZN(n5047) );
  NAND4_X1 U5551 ( .A1(n5050), .A2(n5049), .A3(n5048), .A4(n5047), .ZN(n5051)
         );
  NOR3_X1 U5552 ( .A1(n5053), .A2(n5052), .A3(n5051), .ZN(n5067) );
  AOI22_X1 U5553 ( .A1(n5055), .A2(keyinput_f25), .B1(n2784), .B2(keyinput_f74), .ZN(n5054) );
  OAI221_X1 U5554 ( .B1(n5055), .B2(keyinput_f25), .C1(n2784), .C2(
        keyinput_f74), .A(n5054), .ZN(n5065) );
  AOI22_X1 U5555 ( .A1(n5058), .A2(keyinput_f54), .B1(keyinput_f17), .B2(n5057), .ZN(n5056) );
  OAI221_X1 U5556 ( .B1(n5058), .B2(keyinput_f54), .C1(n5057), .C2(
        keyinput_f17), .A(n5056), .ZN(n5064) );
  XOR2_X1 U5557 ( .A(n2618), .B(keyinput_f63), .Z(n5062) );
  XNOR2_X1 U5558 ( .A(IR_REG_26__SCAN_IN), .B(keyinput_f81), .ZN(n5061) );
  XNOR2_X1 U5559 ( .A(DATAI_7_), .B(keyinput_f24), .ZN(n5060) );
  XNOR2_X1 U5560 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_f57), .ZN(n5059) );
  NAND4_X1 U5561 ( .A1(n5062), .A2(n5061), .A3(n5060), .A4(n5059), .ZN(n5063)
         );
  NOR3_X1 U5562 ( .A1(n5065), .A2(n5064), .A3(n5063), .ZN(n5066) );
  NAND4_X1 U5563 ( .A1(n5069), .A2(n5068), .A3(n5067), .A4(n5066), .ZN(n5070)
         );
  NOR4_X1 U5564 ( .A1(n5073), .A2(n5072), .A3(n5071), .A4(n5070), .ZN(n5074)
         );
  NAND2_X1 U5565 ( .A1(n5075), .A2(n5074), .ZN(n5077) );
  AOI21_X1 U5566 ( .B1(keyinput_f28), .B2(n5077), .A(keyinput_g28), .ZN(n5079)
         );
  INV_X1 U5567 ( .A(keyinput_f28), .ZN(n5076) );
  AOI21_X1 U5568 ( .B1(n5077), .B2(n5076), .A(n5080), .ZN(n5078) );
  AOI22_X1 U5569 ( .A1(n5080), .A2(n5079), .B1(keyinput_g28), .B2(n5078), .ZN(
        n5081) );
  AOI21_X1 U5570 ( .B1(n5083), .B2(n5082), .A(n5081), .ZN(n5085) );
  AOI22_X1 U5571 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n5084) );
  XNOR2_X1 U5572 ( .A(n5085), .B(n5084), .ZN(U3352) );
  INV_X4 U3758 ( .A(n3551), .ZN(n3479) );
  INV_X1 U2463 ( .A(n3225), .ZN(n4680) );
endmodule

