

module b17_C_AntiSAT_k_128_5 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9605, n9606, n9607, n9608, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838;

  XNOR2_X1 U11049 ( .A(n12405), .B(n12404), .ZN(n14221) );
  AND2_X1 U11050 ( .A1(n12587), .A2(n12590), .ZN(n13859) );
  NOR2_X1 U11051 ( .A1(n14886), .A2(n12603), .ZN(n14694) );
  NAND2_X1 U11052 ( .A1(n15586), .A2(n12556), .ZN(n13538) );
  OAI21_X1 U11053 ( .B1(n15457), .B2(n15456), .A(n18615), .ZN(n15459) );
  CLKBUF_X1 U11054 ( .A(n10318), .Z(n11155) );
  NAND4_X1 U11055 ( .A1(n10408), .A2(n10407), .A3(n10406), .A4(n10405), .ZN(
        n10448) );
  AOI21_X1 U11056 ( .B1(n19114), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n10398), .ZN(n10406) );
  AND2_X1 U11057 ( .A1(n10332), .A2(n11290), .ZN(n19202) );
  OR2_X1 U11058 ( .A1(n15014), .A2(n18815), .ZN(n10333) );
  NOR2_X1 U11059 ( .A1(n13716), .A2(n13715), .ZN(n16642) );
  NAND2_X1 U11060 ( .A1(n10330), .A2(n10329), .ZN(n11062) );
  CLKBUF_X2 U11061 ( .A(n15201), .Z(n16934) );
  OR2_X2 U11062 ( .A1(n15238), .A2(n15237), .ZN(n17139) );
  BUF_X2 U11063 ( .A(n13772), .Z(n9614) );
  AOI21_X1 U11064 ( .B1(n10295), .B2(n15019), .A(n10296), .ZN(n10300) );
  INV_X2 U11065 ( .A(n16646), .ZN(n16927) );
  CLKBUF_X2 U11066 ( .A(n15225), .Z(n16896) );
  CLKBUF_X3 U11067 ( .A(n13772), .Z(n9613) );
  AND2_X1 U11068 ( .A1(n10371), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10429) );
  INV_X1 U11069 ( .A(n12979), .ZN(n11416) );
  BUF_X1 U11071 ( .A(n9632), .Z(n12315) );
  CLKBUF_X2 U11073 ( .A(n11667), .Z(n12385) );
  CLKBUF_X2 U11074 ( .A(n11681), .Z(n12242) );
  CLKBUF_X2 U11075 ( .A(n11995), .Z(n12314) );
  NAND2_X1 U11076 ( .A1(n10200), .A2(n10199), .ZN(n18965) );
  NAND2_X1 U11077 ( .A1(n10141), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10142) );
  INV_X2 U11078 ( .A(n10247), .ZN(n11600) );
  AND2_X1 U11079 ( .A1(n11613), .A2(n11612), .ZN(n11775) );
  AND2_X1 U11080 ( .A1(n11612), .A2(n11615), .ZN(n11877) );
  AND2_X1 U11081 ( .A1(n11604), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11614) );
  CLKBUF_X2 U11082 ( .A(n10182), .Z(n10221) );
  BUF_X1 U11084 ( .A(n11398), .Z(n9625) );
  INV_X1 U11085 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11606) );
  CLKBUF_X1 U11086 ( .A(n19886), .Z(n9605) );
  NOR2_X1 U11087 ( .A1(n19839), .A2(n19841), .ZN(n19886) );
  CLKBUF_X1 U11088 ( .A(n19885), .Z(n9606) );
  NOR2_X1 U11089 ( .A1(n19841), .A2(n19840), .ZN(n19885) );
  CLKBUF_X1 U11090 ( .A(n18827), .Z(n9607) );
  NOR2_X1 U11091 ( .A1(n18669), .A2(n19582), .ZN(n18827) );
  OR2_X1 U11093 ( .A1(n13065), .A2(n11734), .ZN(n11750) );
  AND2_X1 U11095 ( .A1(n11605), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10098) );
  NAND2_X1 U11096 ( .A1(n11750), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11819) );
  NOR2_X2 U11097 ( .A1(n19863), .A2(n19868), .ZN(n11739) );
  NOR2_X1 U11098 ( .A1(n11922), .A2(n11921), .ZN(n11935) );
  AND2_X1 U11099 ( .A1(n13251), .A2(n9761), .ZN(n9760) );
  AOI22_X1 U11100 ( .A1(n11689), .A2(n9967), .B1(n11690), .B2(n19863), .ZN(
        n9810) );
  NOR2_X2 U11101 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15390) );
  INV_X1 U11102 ( .A(n18965), .ZN(n10254) );
  AND2_X1 U11103 ( .A1(n11290), .A2(n15014), .ZN(n10364) );
  AND4_X1 U11104 ( .A1(n11710), .A2(n11709), .A3(n11708), .A4(n9667), .ZN(
        n19844) );
  NAND2_X1 U11105 ( .A1(n12788), .A2(n9618), .ZN(n13832) );
  INV_X2 U11107 ( .A(n11080), .ZN(n11148) );
  AND2_X1 U11108 ( .A1(n10301), .A2(n10314), .ZN(n10302) );
  NAND2_X1 U11109 ( .A1(n16086), .A2(n10252), .ZN(n15006) );
  AND2_X1 U11110 ( .A1(n10334), .A2(n12893), .ZN(n10468) );
  AND2_X1 U11111 ( .A1(n10334), .A2(n11290), .ZN(n19260) );
  NAND2_X1 U11112 ( .A1(n10364), .A2(n10354), .ZN(n19358) );
  BUF_X1 U11114 ( .A(n9953), .Z(n9947) );
  INV_X1 U11115 ( .A(n13840), .ZN(n13821) );
  INV_X1 U11116 ( .A(n15529), .ZN(n14342) );
  NAND2_X1 U11117 ( .A1(n10099), .A2(n9683), .ZN(n15586) );
  AND2_X1 U11118 ( .A1(n15674), .A2(n19829), .ZN(n15702) );
  NAND2_X1 U11119 ( .A1(n10215), .A2(n10214), .ZN(n10855) );
  NAND2_X1 U11120 ( .A1(n14825), .A2(n9965), .ZN(n9963) );
  INV_X1 U11121 ( .A(n11039), .ZN(n11043) );
  NAND2_X1 U11122 ( .A1(n10306), .A2(n10307), .ZN(n10305) );
  AND2_X1 U11123 ( .A1(n10332), .A2(n12893), .ZN(n10467) );
  INV_X1 U11124 ( .A(n11272), .ZN(n10253) );
  AND3_X1 U11125 ( .A1(n18424), .A2(n18622), .A3(n16323), .ZN(n15457) );
  XNOR2_X1 U11126 ( .A(n15259), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17615) );
  OR2_X1 U11127 ( .A1(n11659), .A2(n11658), .ZN(n11844) );
  XNOR2_X1 U11128 ( .A(n12528), .B(n12527), .ZN(n13251) );
  AND2_X1 U11129 ( .A1(n13081), .A2(n15396), .ZN(n19833) );
  INV_X1 U11130 ( .A(n11290), .ZN(n10350) );
  INV_X2 U11131 ( .A(n12844), .ZN(n18981) );
  BUF_X1 U11132 ( .A(n11290), .Z(n15954) );
  NAND2_X2 U11133 ( .A1(n10304), .A2(n10315), .ZN(n15014) );
  AND2_X1 U11134 ( .A1(n10305), .A2(n10336), .ZN(n18815) );
  INV_X1 U11135 ( .A(n18005), .ZN(n17108) );
  INV_X1 U11136 ( .A(n17534), .ZN(n17516) );
  INV_X1 U11137 ( .A(n15034), .ZN(n15033) );
  INV_X1 U11138 ( .A(n19663), .ZN(n15521) );
  INV_X1 U11139 ( .A(n19703), .ZN(n19731) );
  OAI21_X1 U11140 ( .B1(n14102), .B2(n14104), .A(n14103), .ZN(n15473) );
  INV_X1 U11141 ( .A(n15014), .ZN(n12756) );
  OR2_X1 U11142 ( .A1(n18449), .A2(n18459), .ZN(n16308) );
  OAI21_X1 U11143 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18614), .A(n16308), 
        .ZN(n17625) );
  AND2_X2 U11144 ( .A1(n9867), .A2(n9866), .ZN(n9608) );
  INV_X1 U11145 ( .A(n9615), .ZN(n15190) );
  INV_X4 U11146 ( .A(n17861), .ZN(n17951) );
  AND2_X2 U11147 ( .A1(n11614), .A2(n11613), .ZN(n11667) );
  AND2_X2 U11148 ( .A1(n10098), .A2(n15390), .ZN(n11681) );
  BUF_X4 U11150 ( .A(n10527), .Z(n9610) );
  INV_X2 U11151 ( .A(n10232), .ZN(n10527) );
  NOR2_X2 U11152 ( .A1(n11241), .A2(n14710), .ZN(n11240) );
  XNOR2_X2 U11153 ( .A(n15288), .B(n15287), .ZN(n17545) );
  NAND2_X2 U11154 ( .A1(n12541), .A2(n12540), .ZN(n15594) );
  NAND2_X2 U11155 ( .A1(n10842), .A2(n9687), .ZN(n13600) );
  NAND2_X2 U11157 ( .A1(n9792), .A2(n10847), .ZN(n15905) );
  CLKBUF_X2 U11158 ( .A(n11990), .Z(n9631) );
  NOR3_X2 U11159 ( .A1(n17202), .A2(n17073), .A3(n17039), .ZN(n17035) );
  AOI21_X2 U11160 ( .B1(n10318), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n10294), .ZN(n10299) );
  AND2_X4 U11162 ( .A1(n10377), .A2(n16072), .ZN(n10182) );
  NOR2_X2 U11163 ( .A1(n10625), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10619) );
  NOR2_X2 U11164 ( .A1(n17848), .A2(n18433), .ZN(n18399) );
  NAND2_X2 U11165 ( .A1(n10251), .A2(n10250), .ZN(n10284) );
  AND2_X1 U11166 ( .A1(n11614), .A2(n13210), .ZN(n9611) );
  AND2_X2 U11167 ( .A1(n11614), .A2(n13210), .ZN(n9612) );
  NOR2_X1 U11168 ( .A1(n13688), .A2(n13687), .ZN(n13772) );
  NAND2_X2 U11169 ( .A1(n10143), .A2(n10142), .ZN(n18958) );
  OAI21_X2 U11170 ( .B1(n14591), .B2(n10078), .A(n10077), .ZN(n11474) );
  INV_X2 U11171 ( .A(n12686), .ZN(n12874) );
  INV_X4 U11172 ( .A(n9668), .ZN(n16937) );
  OAI22_X2 U11173 ( .A1(n12631), .A2(n12630), .B1(n10898), .B2(n10897), .ZN(
        n12951) );
  NOR2_X1 U11175 ( .A1(n16689), .A2(n9939), .ZN(n9676) );
  AND2_X1 U11176 ( .A1(n10376), .A2(n9783), .ZN(n9616) );
  INV_X1 U11177 ( .A(n9616), .ZN(n9617) );
  NOR2_X4 U11178 ( .A1(n16191), .A2(n17114), .ZN(n17534) );
  NOR2_X1 U11179 ( .A1(n14603), .A2(n14604), .ZN(n13875) );
  XNOR2_X1 U11180 ( .A(n10850), .B(n10849), .ZN(n11211) );
  NAND2_X1 U11181 ( .A1(n10610), .A2(n9647), .ZN(n15889) );
  NAND2_X1 U11182 ( .A1(n17693), .A2(n17300), .ZN(n17672) );
  AND2_X1 U11183 ( .A1(n11297), .A2(n11317), .ZN(n12890) );
  INV_X1 U11185 ( .A(n14990), .ZN(n12777) );
  OAI21_X1 U11186 ( .B1(n18402), .B2(n15332), .A(n18401), .ZN(n17848) );
  AND3_X1 U11187 ( .A1(n9929), .A2(n9931), .A3(n9928), .ZN(n17594) );
  OAI21_X1 U11188 ( .B1(n11750), .B2(n11744), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11746) );
  AOI211_X1 U11189 ( .C1(n16642), .C2(n15155), .A(n15154), .B(n15153), .ZN(
        n15166) );
  AND3_X1 U11190 ( .A1(n16108), .A2(n10252), .A3(n12876), .ZN(n10262) );
  INV_X2 U11191 ( .A(n11153), .ZN(n11080) );
  NAND2_X2 U11193 ( .A1(n10792), .A2(n10267), .ZN(n11153) );
  NOR2_X1 U11194 ( .A1(n12448), .A2(n12557), .ZN(n12457) );
  INV_X2 U11195 ( .A(n15309), .ZN(n17997) );
  NAND2_X1 U11197 ( .A1(n12465), .A2(n11844), .ZN(n13054) );
  INV_X2 U11198 ( .A(n19844), .ZN(n9618) );
  INV_X1 U11199 ( .A(n15112), .ZN(n15260) );
  CLKBUF_X2 U11200 ( .A(n11682), .Z(n12148) );
  BUF_X2 U11201 ( .A(n11661), .Z(n12384) );
  BUF_X1 U11202 ( .A(n11660), .Z(n9632) );
  BUF_X2 U11203 ( .A(n11662), .Z(n12200) );
  CLKBUF_X2 U11204 ( .A(n13732), .Z(n16946) );
  CLKBUF_X2 U11205 ( .A(n15263), .Z(n16953) );
  CLKBUF_X2 U11206 ( .A(n11769), .Z(n12309) );
  BUF_X2 U11207 ( .A(n10154), .Z(n11567) );
  BUF_X2 U11208 ( .A(n11566), .Z(n11522) );
  AND2_X1 U11209 ( .A1(n10129), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10377) );
  NAND2_X1 U11210 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n13689), .ZN(
        n13687) );
  BUF_X2 U11211 ( .A(n15265), .Z(n9619) );
  AND2_X1 U11212 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12971) );
  INV_X1 U11213 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10131) );
  NAND2_X1 U11214 ( .A1(n12605), .A2(n12604), .ZN(n13874) );
  AND2_X1 U11215 ( .A1(n14682), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14656) );
  AOI21_X1 U11216 ( .B1(n13875), .B2(n13876), .A(n10023), .ZN(n10743) );
  OAI21_X1 U11217 ( .B1(n11211), .B2(n15941), .A(n10084), .ZN(n11219) );
  INV_X1 U11218 ( .A(n14912), .ZN(n14939) );
  AND2_X1 U11219 ( .A1(n10092), .A2(n10090), .ZN(n13912) );
  AOI211_X1 U11220 ( .C1(n14769), .C2(n16033), .A(n14768), .B(n14767), .ZN(
        n14770) );
  NAND2_X1 U11221 ( .A1(n9608), .A2(n9753), .ZN(n14886) );
  AOI211_X1 U11222 ( .C1(n15476), .C2(n19703), .A(n15475), .B(n15474), .ZN(
        n15479) );
  AOI21_X1 U11223 ( .B1(n14000), .B2(n14094), .A(n13999), .ZN(n14273) );
  NOR2_X1 U11224 ( .A1(n14614), .A2(n14613), .ZN(n14615) );
  OAI21_X1 U11225 ( .B1(n12590), .B2(n12588), .A(n12589), .ZN(n14153) );
  CLKBUF_X1 U11226 ( .A(n12587), .Z(n12588) );
  OAI21_X1 U11227 ( .B1(n14276), .B2(n13853), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9777) );
  NOR2_X1 U11228 ( .A1(n13943), .A2(n13944), .ZN(n12587) );
  NAND2_X1 U11229 ( .A1(n12579), .A2(n14342), .ZN(n14276) );
  NAND2_X1 U11230 ( .A1(n12581), .A2(n15529), .ZN(n14275) );
  NAND2_X1 U11231 ( .A1(n14544), .A2(n14543), .ZN(n14542) );
  XNOR2_X1 U11232 ( .A(n11474), .B(n11470), .ZN(n14544) );
  NAND2_X1 U11233 ( .A1(n15937), .A2(n15936), .ZN(n15934) );
  AND2_X1 U11234 ( .A1(n11367), .A2(n10080), .ZN(n11429) );
  OR2_X1 U11235 ( .A1(n13275), .A2(n13276), .ZN(n13364) );
  NOR2_X1 U11236 ( .A1(n10110), .A2(n14342), .ZN(n10109) );
  AND2_X2 U11237 ( .A1(n11325), .A2(n9737), .ZN(n13552) );
  AND3_X1 U11238 ( .A1(n9680), .A2(n14315), .A3(n9811), .ZN(n10110) );
  AND2_X1 U11239 ( .A1(n10550), .A2(n10123), .ZN(n10072) );
  NAND2_X1 U11240 ( .A1(n9791), .A2(n10822), .ZN(n10823) );
  OR2_X1 U11241 ( .A1(n9926), .A2(n17534), .ZN(n9924) );
  AND2_X1 U11242 ( .A1(n14307), .A2(n14304), .ZN(n14305) );
  AND2_X1 U11243 ( .A1(n12566), .A2(n9701), .ZN(n10100) );
  AND2_X1 U11244 ( .A1(n14298), .A2(n10108), .ZN(n10107) );
  AND2_X1 U11245 ( .A1(n17303), .A2(n17648), .ZN(n9926) );
  NAND2_X1 U11246 ( .A1(n11974), .A2(n11973), .ZN(n13392) );
  AND3_X1 U11247 ( .A1(n17319), .A2(n17312), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17304) );
  OR2_X1 U11248 ( .A1(n15529), .A2(n12575), .ZN(n14315) );
  AND2_X1 U11249 ( .A1(n11964), .A2(n11938), .ZN(n12531) );
  XNOR2_X1 U11250 ( .A(n12561), .B(n11967), .ZN(n12547) );
  NAND2_X2 U11251 ( .A1(n12561), .A2(n12560), .ZN(n15529) );
  OR2_X1 U11252 ( .A1(n19842), .A2(n12022), .ZN(n11897) );
  INV_X1 U11253 ( .A(n10396), .ZN(n19167) );
  AOI221_X1 U11254 ( .B1(n17411), .B2(n17338), .C1(n17701), .C2(n17338), .A(
        n17363), .ZN(n17340) );
  NAND2_X1 U11255 ( .A1(n10670), .A2(n10714), .ZN(n10664) );
  OAI211_X1 U11256 ( .C1(n9774), .C2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n9772), .B(n9770), .ZN(n13120) );
  AND4_X1 U11257 ( .A1(n10473), .A2(n10472), .A3(n10471), .A4(n10470), .ZN(
        n10481) );
  NAND2_X1 U11258 ( .A1(n10351), .A2(n10354), .ZN(n10580) );
  AND2_X1 U11259 ( .A1(n10461), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10398) );
  OR2_X1 U11260 ( .A1(n10362), .A2(n10359), .ZN(n10396) );
  NOR2_X1 U11261 ( .A1(n17108), .A2(n17034), .ZN(n17030) );
  OR2_X1 U11262 ( .A1(n10669), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10670) );
  OAI21_X1 U11263 ( .B1(n13225), .B2(n12557), .A(n12498), .ZN(n13121) );
  NAND2_X1 U11264 ( .A1(n10364), .A2(n10363), .ZN(n10476) );
  INV_X1 U11265 ( .A(n10392), .ZN(n18993) );
  AND2_X1 U11266 ( .A1(n15293), .A2(n9937), .ZN(n9936) );
  NAND2_X1 U11267 ( .A1(n10364), .A2(n9955), .ZN(n19332) );
  CLKBUF_X1 U11268 ( .A(n12488), .Z(n14198) );
  AND2_X1 U11269 ( .A1(n15294), .A2(n10125), .ZN(n15293) );
  AND2_X1 U11270 ( .A1(n10641), .A2(n9649), .ZN(n10675) );
  NAND2_X1 U11271 ( .A1(n13081), .A2(n13073), .ZN(n19829) );
  INV_X2 U11272 ( .A(n19747), .ZN(n19776) );
  NAND2_X2 U11273 ( .A1(n14210), .A2(n12963), .ZN(n14209) );
  NAND2_X1 U11274 ( .A1(n10643), .A2(n10714), .ZN(n10641) );
  XNOR2_X1 U11275 ( .A(n12887), .B(n12886), .ZN(n19590) );
  NOR2_X1 U11276 ( .A1(n10333), .A2(n12777), .ZN(n10334) );
  NOR2_X1 U11277 ( .A1(n10333), .A2(n14990), .ZN(n10332) );
  AND2_X1 U11278 ( .A1(n20838), .A2(n17862), .ZN(n9951) );
  NAND2_X1 U11279 ( .A1(n9803), .A2(n11888), .ZN(n11889) );
  CLKBUF_X1 U11280 ( .A(n16682), .Z(n16675) );
  NAND2_X1 U11281 ( .A1(n15424), .A2(n13052), .ZN(n13058) );
  NAND2_X1 U11282 ( .A1(n13201), .A2(n15763), .ZN(n9803) );
  NAND2_X1 U11283 ( .A1(n10338), .A2(n10313), .ZN(n14990) );
  NOR2_X2 U11284 ( .A1(n18959), .A2(n19171), .ZN(n18960) );
  NOR2_X2 U11285 ( .A1(n18966), .A2(n19171), .ZN(n18967) );
  NOR2_X2 U11286 ( .A1(n18945), .A2(n19171), .ZN(n18946) );
  NOR2_X2 U11287 ( .A1(n18951), .A2(n19171), .ZN(n18952) );
  NAND2_X1 U11288 ( .A1(n12459), .A2(n12458), .ZN(n15424) );
  NAND2_X1 U11289 ( .A1(n10031), .A2(n10030), .ZN(n10625) );
  AND2_X1 U11290 ( .A1(n13158), .A2(n10896), .ZN(n12631) );
  INV_X1 U11291 ( .A(n10616), .ZN(n10031) );
  NOR2_X2 U11292 ( .A1(n17188), .A2(n17899), .ZN(n18428) );
  NAND2_X1 U11293 ( .A1(n12456), .A2(n12455), .ZN(n12459) );
  NAND2_X1 U11294 ( .A1(n9835), .A2(n11827), .ZN(n13216) );
  NAND2_X1 U11295 ( .A1(n10310), .A2(n10288), .ZN(n10303) );
  NAND2_X1 U11296 ( .A1(n10105), .A2(n11858), .ZN(n19925) );
  NAND2_X1 U11297 ( .A1(n11061), .A2(n10326), .ZN(n10328) );
  NOR2_X1 U11298 ( .A1(n11816), .A2(n11815), .ZN(n11817) );
  XNOR2_X1 U11299 ( .A(n11816), .B(n11814), .ZN(n11848) );
  NAND2_X1 U11300 ( .A1(n11823), .A2(n11822), .ZN(n9835) );
  OAI21_X1 U11301 ( .B1(n13236), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n9974), 
        .ZN(n11816) );
  AND2_X1 U11302 ( .A1(n11794), .A2(n11793), .ZN(n11768) );
  NAND2_X1 U11303 ( .A1(n11876), .A2(n11875), .ZN(n20003) );
  OAI211_X1 U11304 ( .C1(n15422), .C2(n20148), .A(n11826), .B(n11825), .ZN(
        n11827) );
  NAND3_X1 U11305 ( .A1(n15325), .A2(n15168), .A3(n15162), .ZN(n15332) );
  NOR2_X2 U11306 ( .A1(n18621), .A2(n17249), .ZN(n17241) );
  NAND2_X1 U11307 ( .A1(n11746), .A2(n11745), .ZN(n11824) );
  NAND2_X1 U11308 ( .A1(n10529), .A2(n10528), .ZN(n10555) );
  AND2_X1 U11309 ( .A1(n12856), .A2(n12857), .ZN(n12859) );
  AOI21_X1 U11310 ( .B1(n12903), .B2(n15391), .A(n12895), .ZN(n11753) );
  OR2_X1 U11311 ( .A1(n15329), .A2(n17981), .ZN(n15159) );
  OR2_X1 U11312 ( .A1(n17122), .A2(n15284), .ZN(n15285) );
  INV_X1 U11313 ( .A(n12448), .ZN(n12443) );
  OR2_X1 U11314 ( .A1(n12896), .A2(n13054), .ZN(n13061) );
  CLKBUF_X1 U11315 ( .A(n10273), .Z(n11169) );
  AND2_X1 U11316 ( .A1(n10246), .A2(n11168), .ZN(n11581) );
  AND2_X2 U11317 ( .A1(n12681), .A2(n12876), .ZN(n16086) );
  NOR2_X1 U11318 ( .A1(n17971), .A2(n18005), .ZN(n15161) );
  NAND2_X1 U11319 ( .A1(n11736), .A2(n12466), .ZN(n9809) );
  OR2_X2 U11320 ( .A1(n12414), .A2(n15763), .ZN(n12448) );
  INV_X1 U11321 ( .A(n10615), .ZN(n10030) );
  NAND2_X1 U11322 ( .A1(n13838), .A2(n13821), .ZN(n13829) );
  AND2_X1 U11323 ( .A1(n11735), .A2(n11844), .ZN(n11761) );
  AND2_X1 U11324 ( .A1(n12814), .A2(n12686), .ZN(n10267) );
  AND2_X2 U11325 ( .A1(n10852), .A2(n19582), .ZN(n11039) );
  AND2_X1 U11326 ( .A1(n10254), .A2(n18958), .ZN(n11168) );
  NOR2_X1 U11327 ( .A1(n15308), .A2(n17993), .ZN(n15319) );
  INV_X2 U11328 ( .A(n16642), .ZN(n17971) );
  NOR2_X2 U11329 ( .A1(n13706), .A2(n13705), .ZN(n18621) );
  NOR2_X1 U11330 ( .A1(n18005), .A2(n17985), .ZN(n15326) );
  INV_X1 U11332 ( .A(n18958), .ZN(n11163) );
  AND2_X1 U11333 ( .A1(n11272), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12814) );
  AND2_X1 U11334 ( .A1(n11739), .A2(n12503), .ZN(n12998) );
  INV_X1 U11335 ( .A(n19858), .ZN(n11733) );
  NAND3_X1 U11336 ( .A1(n15274), .A2(n15273), .A3(n15272), .ZN(n17623) );
  NAND2_X1 U11337 ( .A1(n10153), .A2(n9783), .ZN(n9780) );
  NAND2_X1 U11338 ( .A1(n10152), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9781) );
  NAND2_X1 U11339 ( .A1(n10188), .A2(n10187), .ZN(n10247) );
  AND4_X1 U11340 ( .A1(n11710), .A2(n11709), .A3(n11708), .A4(n9667), .ZN(
        n9630) );
  NAND2_X1 U11341 ( .A1(n9671), .A2(n10128), .ZN(n11676) );
  AND4_X1 U11342 ( .A1(n11623), .A2(n11622), .A3(n11621), .A4(n11620), .ZN(
        n11639) );
  AND4_X1 U11343 ( .A1(n11631), .A2(n11630), .A3(n11629), .A4(n11628), .ZN(
        n11637) );
  AND4_X1 U11344 ( .A1(n11694), .A2(n11693), .A3(n11692), .A4(n11691), .ZN(
        n11710) );
  AND4_X1 U11345 ( .A1(n10207), .A2(n10206), .A3(n10205), .A4(n10204), .ZN(
        n10208) );
  AND4_X1 U11346 ( .A1(n11619), .A2(n11618), .A3(n11617), .A4(n11616), .ZN(
        n10128) );
  NAND2_X1 U11347 ( .A1(n10181), .A2(n10180), .ZN(n10188) );
  AND4_X1 U11348 ( .A1(n10151), .A2(n10150), .A3(n10149), .A4(n10148), .ZN(
        n10152) );
  INV_X2 U11349 ( .A(n18302), .ZN(n18000) );
  AND4_X1 U11350 ( .A1(n11715), .A2(n11714), .A3(n11713), .A4(n11712), .ZN(
        n11731) );
  AND4_X1 U11351 ( .A1(n10147), .A2(n10146), .A3(n10145), .A4(n10144), .ZN(
        n10153) );
  AND4_X1 U11352 ( .A1(n11635), .A2(n11634), .A3(n11633), .A4(n11632), .ZN(
        n11636) );
  AND4_X1 U11353 ( .A1(n10179), .A2(n10178), .A3(n10177), .A4(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10181) );
  INV_X2 U11354 ( .A(n16291), .ZN(U215) );
  AND4_X1 U11355 ( .A1(n11627), .A2(n11626), .A3(n11625), .A4(n11624), .ZN(
        n11638) );
  AND4_X1 U11356 ( .A1(n11703), .A2(n11702), .A3(n11701), .A4(n11700), .ZN(
        n11708) );
  AND4_X1 U11357 ( .A1(n11698), .A2(n11697), .A3(n11696), .A4(n11695), .ZN(
        n11709) );
  AND4_X1 U11358 ( .A1(n11723), .A2(n11722), .A3(n11721), .A4(n11720), .ZN(
        n11729) );
  AND4_X1 U11359 ( .A1(n11719), .A2(n11718), .A3(n11717), .A4(n11716), .ZN(
        n11730) );
  AND2_X2 U11360 ( .A1(n11522), .A2(n9783), .ZN(n11417) );
  OR2_X1 U11362 ( .A1(n11252), .A2(n11216), .ZN(n11258) );
  AND2_X2 U11363 ( .A1(n11563), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10794) );
  AND2_X2 U11364 ( .A1(n11563), .A2(n9783), .ZN(n10449) );
  NAND2_X2 U11365 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19627), .ZN(n19569) );
  BUF_X2 U11366 ( .A(n11877), .Z(n11795) );
  NAND2_X2 U11367 ( .A1(n18630), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18553) );
  NOR2_X1 U11368 ( .A1(n9669), .A2(n9916), .ZN(n9915) );
  AND2_X2 U11369 ( .A1(n11613), .A2(n15390), .ZN(n11661) );
  BUF_X2 U11370 ( .A(n11775), .Z(n9621) );
  AND2_X2 U11371 ( .A1(n10377), .A2(n11400), .ZN(n10415) );
  AND2_X2 U11372 ( .A1(n14986), .A2(n11400), .ZN(n10413) );
  AND2_X2 U11373 ( .A1(n10098), .A2(n11612), .ZN(n11682) );
  BUF_X2 U11374 ( .A(n15102), .Z(n16947) );
  CLKBUF_X2 U11375 ( .A(n12221), .Z(n12243) );
  INV_X2 U11376 ( .A(n16295), .ZN(n16297) );
  NOR2_X1 U11377 ( .A1(n13686), .A2(n16689), .ZN(n13770) );
  NOR2_X1 U11378 ( .A1(n18434), .A2(n13686), .ZN(n15225) );
  NOR3_X1 U11379 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n13687), .ZN(n15263) );
  AND2_X2 U11380 ( .A1(n12971), .A2(n16072), .ZN(n10370) );
  OR2_X1 U11381 ( .A1(n18434), .A2(n13688), .ZN(n16646) );
  NAND2_X1 U11382 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18583), .ZN(
        n13680) );
  NOR2_X1 U11383 ( .A1(n9868), .A2(n15872), .ZN(n9866) );
  NAND2_X1 U11384 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18574), .ZN(
        n13686) );
  AND2_X2 U11385 ( .A1(n15004), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11398) );
  AND2_X2 U11386 ( .A1(n15390), .A2(n11615), .ZN(n12221) );
  AND2_X2 U11387 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10795) );
  NOR2_X1 U11388 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10378) );
  BUF_X2 U11389 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n15019) );
  INV_X1 U11390 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18591) );
  NOR2_X2 U11391 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11615) );
  INV_X1 U11392 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16072) );
  NOR2_X2 U11393 ( .A1(n11248), .A2(n11250), .ZN(n11249) );
  NOR2_X1 U11394 ( .A1(n17356), .A2(n17363), .ZN(n17395) );
  NAND2_X1 U11395 ( .A1(n10245), .A2(n10244), .ZN(n12876) );
  XNOR2_X2 U11396 ( .A(n14608), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14757) );
  AND2_X1 U11397 ( .A1(n11613), .A2(n15389), .ZN(n11660) );
  NAND2_X1 U11398 ( .A1(n12983), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9774) );
  MUX2_X1 U11399 ( .A(n14238), .B(n14237), .S(n14342), .Z(n14239) );
  NOR2_X4 U11400 ( .A1(n14607), .A2(n14772), .ZN(n14608) );
  NAND2_X2 U11401 ( .A1(n15846), .A2(n9752), .ZN(n14607) );
  OR2_X1 U11402 ( .A1(n12962), .A2(n11738), .ZN(n15391) );
  NAND2_X2 U11403 ( .A1(n13064), .A2(n12415), .ZN(n11690) );
  NAND2_X1 U11404 ( .A1(n11760), .A2(n12415), .ZN(n12962) );
  AND4_X1 U11405 ( .A1(n12503), .A2(n13064), .A3(n11844), .A4(n11760), .ZN(
        n9828) );
  NOR2_X2 U11406 ( .A1(n16195), .A2(n17628), .ZN(n17452) );
  NOR3_X2 U11407 ( .A1(n13782), .A2(n15165), .A3(n18403), .ZN(n15331) );
  INV_X1 U11408 ( .A(n13343), .ZN(n9767) );
  NAND3_X1 U11409 ( .A1(n10387), .A2(n10448), .A3(n9658), .ZN(n9844) );
  AND2_X4 U11410 ( .A1(n15004), .A2(n10131), .ZN(n10154) );
  NAND2_X1 U11411 ( .A1(n9767), .A2(n15763), .ZN(n9766) );
  NOR2_X2 U11412 ( .A1(n17215), .A2(n17011), .ZN(n17004) );
  AND2_X1 U11413 ( .A1(n12971), .A2(n16072), .ZN(n9623) );
  AND2_X2 U11414 ( .A1(n12971), .A2(n16072), .ZN(n9624) );
  AOI211_X2 U11415 ( .C1(n18934), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n13882), .B(n13881), .ZN(n13883) );
  NAND2_X2 U11416 ( .A1(n9630), .A2(n9633), .ZN(n11756) );
  BUF_X8 U11417 ( .A(n11398), .Z(n9626) );
  NAND2_X2 U11418 ( .A1(n9966), .A2(n11740), .ZN(n12467) );
  BUF_X1 U11419 ( .A(n13787), .Z(n9627) );
  INV_X2 U11420 ( .A(n16912), .ZN(n9628) );
  INV_X2 U11421 ( .A(n11737), .ZN(n13064) );
  NAND4_X1 U11422 ( .A1(n11710), .A2(n11709), .A3(n11708), .A4(n9667), .ZN(
        n9629) );
  AND2_X2 U11423 ( .A1(n11229), .A2(n9662), .ZN(n11217) );
  NOR2_X4 U11424 ( .A1(n11231), .A2(n14629), .ZN(n11229) );
  NOR4_X1 U11425 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n13689), .A4(n18574), .ZN(
        n15265) );
  NAND2_X1 U11426 ( .A1(n9829), .A2(n12526), .ZN(n12528) );
  AOI21_X4 U11427 ( .B1(n11848), .B2(n12499), .A(n11817), .ZN(n11843) );
  AND2_X2 U11428 ( .A1(n11236), .A2(n9910), .ZN(n11232) );
  NOR2_X4 U11429 ( .A1(n11238), .A2(n14683), .ZN(n11236) );
  INV_X1 U11430 ( .A(n19858), .ZN(n9633) );
  AND2_X2 U11431 ( .A1(n13493), .A2(n12007), .ZN(n13546) );
  NOR2_X2 U11432 ( .A1(n13391), .A2(n13494), .ZN(n13493) );
  NOR2_X2 U11433 ( .A1(n14038), .A2(n9976), .ZN(n14110) );
  AND2_X2 U11434 ( .A1(n14110), .A2(n14111), .ZN(n14102) );
  INV_X1 U11435 ( .A(n13264), .ZN(n9634) );
  NAND2_X4 U11436 ( .A1(n9921), .A2(n9923), .ZN(n13264) );
  XNOR2_X1 U11437 ( .A(n11850), .B(n11849), .ZN(n13224) );
  NOR2_X1 U11438 ( .A1(n18621), .A2(n17249), .ZN(n9636) );
  NAND2_X1 U11439 ( .A1(n14342), .A2(n9747), .ZN(n10108) );
  INV_X1 U11440 ( .A(n13331), .ZN(n12397) );
  NAND2_X1 U11441 ( .A1(n20437), .A2(n20334), .ZN(n13331) );
  INV_X1 U11442 ( .A(n9813), .ZN(n9779) );
  AOI21_X1 U11443 ( .B1(n10109), .B2(n10107), .A(n10106), .ZN(n9813) );
  INV_X1 U11444 ( .A(n14293), .ZN(n10106) );
  INV_X1 U11445 ( .A(n11513), .ZN(n11490) );
  INV_X1 U11446 ( .A(n11047), .ZN(n11040) );
  NAND2_X1 U11447 ( .A1(n18981), .A2(n19582), .ZN(n11017) );
  NAND2_X1 U11448 ( .A1(n12839), .A2(n11585), .ZN(n11047) );
  OR2_X1 U11449 ( .A1(n12372), .A2(n12596), .ZN(n13334) );
  AND4_X1 U11450 ( .A1(n10466), .A2(n10465), .A3(n10464), .A4(n10463), .ZN(
        n10482) );
  NAND2_X1 U11451 ( .A1(n11167), .A2(n10254), .ZN(n10241) );
  AND2_X1 U11452 ( .A1(n10603), .A2(n10602), .ZN(n10830) );
  INV_X1 U11453 ( .A(n17544), .ZN(n9953) );
  INV_X1 U11454 ( .A(n9823), .ZN(n13722) );
  OAI21_X1 U11455 ( .B1(n15169), .B2(n15170), .A(n9824), .ZN(n9823) );
  NAND2_X1 U11456 ( .A1(n18413), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9824) );
  AND2_X1 U11458 ( .A1(n12308), .A2(n14104), .ZN(n9985) );
  NOR2_X1 U11459 ( .A1(n9710), .A2(n9972), .ZN(n9971) );
  INV_X1 U11460 ( .A(n11847), .ZN(n9972) );
  NAND2_X1 U11461 ( .A1(n14275), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12584) );
  NAND2_X1 U11462 ( .A1(n11935), .A2(n9800), .ZN(n12561) );
  NOR2_X1 U11463 ( .A1(n9802), .A2(n9801), .ZN(n9800) );
  INV_X1 U11464 ( .A(n11963), .ZN(n9802) );
  NAND2_X1 U11465 ( .A1(n9838), .A2(n13585), .ZN(n9799) );
  INV_X1 U11466 ( .A(n13245), .ZN(n9763) );
  NAND2_X1 U11467 ( .A1(n13840), .A2(n13838), .ZN(n13831) );
  AND3_X1 U11468 ( .A1(n12461), .A2(n11732), .A3(n12460), .ZN(n12916) );
  AND3_X1 U11469 ( .A1(n9715), .A2(n10551), .A3(n10033), .ZN(n10612) );
  NOR2_X1 U11470 ( .A1(n10038), .A2(n10555), .ZN(n10033) );
  INV_X1 U11471 ( .A(n10545), .ZN(n10038) );
  AOI21_X1 U11472 ( .B1(n10289), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10266), .ZN(n10285) );
  INV_X1 U11473 ( .A(n14572), .ZN(n10018) );
  NAND2_X1 U11474 ( .A1(n14533), .A2(n11496), .ZN(n11516) );
  AND2_X1 U11475 ( .A1(n9730), .A2(n13670), .ZN(n10082) );
  NAND2_X1 U11476 ( .A1(n9963), .A2(n9646), .ZN(n10728) );
  AND2_X1 U11477 ( .A1(n9852), .A2(n9851), .ZN(n9850) );
  NOR2_X1 U11478 ( .A1(n13013), .A2(n10016), .ZN(n10015) );
  INV_X1 U11479 ( .A(n12950), .ZN(n10016) );
  NAND2_X1 U11481 ( .A1(n15281), .A2(n15351), .ZN(n15284) );
  NOR2_X1 U11482 ( .A1(n17138), .A2(n15259), .ZN(n15279) );
  OR2_X1 U11483 ( .A1(n15424), .A2(n13191), .ZN(n13000) );
  AND2_X1 U11484 ( .A1(n12375), .A2(n12374), .ZN(n12590) );
  AND2_X1 U11485 ( .A1(n9644), .A2(n12578), .ZN(n9841) );
  NAND2_X1 U11486 ( .A1(n11958), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11968) );
  OAI21_X1 U11487 ( .B1(n13793), .B2(n14342), .A(n13791), .ZN(n14216) );
  NAND2_X1 U11488 ( .A1(n12467), .A2(n9796), .ZN(n13065) );
  NAND2_X1 U11489 ( .A1(n12462), .A2(n13838), .ZN(n9796) );
  AND2_X1 U11490 ( .A1(n11429), .A2(n11452), .ZN(n11430) );
  XNOR2_X1 U11491 ( .A(n11429), .B(n11452), .ZN(n14593) );
  INV_X1 U11492 ( .A(n13139), .ZN(n9991) );
  AND3_X1 U11493 ( .A1(n10890), .A2(n10889), .A3(n10888), .ZN(n13154) );
  AND2_X1 U11494 ( .A1(n10855), .A2(n19582), .ZN(n12839) );
  AND2_X1 U11495 ( .A1(n10055), .A2(n10054), .ZN(n10053) );
  INV_X1 U11496 ( .A(n13549), .ZN(n10054) );
  NAND2_X1 U11497 ( .A1(n9863), .A2(n9862), .ZN(n14674) );
  NOR2_X1 U11498 ( .A1(n14716), .A2(n14670), .ZN(n9862) );
  AOI21_X1 U11499 ( .B1(n14936), .B2(n14933), .A(n14932), .ZN(n14737) );
  AND2_X1 U11500 ( .A1(n10811), .A2(n16106), .ZN(n11182) );
  AND3_X1 U11501 ( .A1(n11206), .A2(n12863), .A3(n10807), .ZN(n10808) );
  NAND2_X1 U11502 ( .A1(n12851), .A2(n11315), .ZN(n12892) );
  XNOR2_X1 U11503 ( .A(n14983), .B(n11309), .ZN(n12887) );
  AOI21_X1 U11504 ( .B1(n14990), .B2(n11308), .A(n11307), .ZN(n12886) );
  NAND2_X1 U11505 ( .A1(n12849), .A2(n12848), .ZN(n12851) );
  NAND2_X1 U11506 ( .A1(n10764), .A2(n10763), .ZN(n16090) );
  CLKBUF_X1 U11507 ( .A(n10247), .Z(n18971) );
  INV_X1 U11508 ( .A(n14927), .ZN(n9788) );
  NAND3_X1 U11509 ( .A1(n9809), .A2(n11761), .A3(n13064), .ZN(n12903) );
  NAND2_X1 U11510 ( .A1(n11935), .A2(n11936), .ZN(n11964) );
  NOR2_X1 U11511 ( .A1(n9768), .A2(n11733), .ZN(n9765) );
  INV_X1 U11512 ( .A(n11430), .ZN(n10079) );
  AND2_X1 U11513 ( .A1(n10496), .A2(n10495), .ZN(n10572) );
  NAND2_X1 U11514 ( .A1(n10575), .A2(n10574), .ZN(n10836) );
  INV_X1 U11515 ( .A(n9844), .ZN(n10575) );
  NOR2_X1 U11516 ( .A1(n10573), .A2(n10821), .ZN(n10574) );
  INV_X1 U11517 ( .A(n10572), .ZN(n10573) );
  INV_X1 U11518 ( .A(n10870), .ZN(n10526) );
  NAND2_X1 U11519 ( .A1(n10240), .A2(n10239), .ZN(n10781) );
  NAND2_X1 U11520 ( .A1(n10232), .A2(n10247), .ZN(n10257) );
  INV_X1 U11521 ( .A(n11168), .ZN(n11166) );
  NAND3_X1 U11522 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n18591), .ZN(n13685) );
  INV_X1 U11523 ( .A(n17981), .ZN(n15308) );
  NAND2_X1 U11524 ( .A1(n13006), .A2(n13005), .ZN(n13093) );
  NOR2_X1 U11525 ( .A1(n14039), .A2(n9980), .ZN(n9979) );
  NAND2_X1 U11526 ( .A1(n13393), .A2(n13392), .ZN(n13391) );
  INV_X1 U11527 ( .A(n11862), .ZN(n12196) );
  NOR2_X1 U11528 ( .A1(n13536), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9836) );
  INV_X1 U11529 ( .A(n15707), .ZN(n9899) );
  NAND2_X1 U11530 ( .A1(n12524), .A2(n10104), .ZN(n9829) );
  NAND2_X1 U11531 ( .A1(n13120), .A2(n13121), .ZN(n12516) );
  NAND2_X1 U11532 ( .A1(n9774), .A2(n12513), .ZN(n12514) );
  NAND2_X1 U11533 ( .A1(n9794), .A2(n11767), .ZN(n19895) );
  AND2_X1 U11534 ( .A1(n11813), .A2(n11812), .ZN(n11814) );
  NOR2_X1 U11535 ( .A1(n9679), .A2(n9975), .ZN(n9974) );
  NOR2_X1 U11536 ( .A1(n12559), .A2(n15763), .ZN(n9975) );
  NAND2_X1 U11537 ( .A1(n11843), .A2(n9973), .ZN(n11890) );
  AND2_X2 U11538 ( .A1(n10234), .A2(n10233), .ZN(n10792) );
  INV_X1 U11539 ( .A(n10257), .ZN(n10233) );
  AND4_X1 U11540 ( .A1(n12844), .A2(n9782), .A3(n18958), .A4(n18965), .ZN(
        n10234) );
  AOI21_X1 U11541 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19588), .A(
        n10540), .ZN(n10745) );
  NOR2_X1 U11542 ( .A1(n10539), .A2(n10538), .ZN(n10540) );
  INV_X1 U11543 ( .A(n10537), .ZN(n10539) );
  INV_X1 U11544 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10041) );
  AND2_X1 U11545 ( .A1(n10664), .A2(n9716), .ZN(n10659) );
  INV_X1 U11546 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10046) );
  NAND2_X1 U11547 ( .A1(n10641), .A2(n10044), .ZN(n10677) );
  INV_X1 U11548 ( .A(n10551), .ZN(n10035) );
  INV_X1 U11549 ( .A(n10556), .ZN(n10037) );
  INV_X1 U11550 ( .A(n10560), .ZN(n10036) );
  NAND2_X1 U11551 ( .A1(n10767), .A2(n9610), .ZN(n10529) );
  AOI21_X1 U11552 ( .B1(n15006), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10249), 
        .ZN(n10250) );
  NOR2_X1 U11553 ( .A1(n15019), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11400) );
  NAND2_X1 U11554 ( .A1(n14542), .A2(n11475), .ZN(n11493) );
  INV_X1 U11555 ( .A(n13553), .ZN(n10075) );
  NOR2_X1 U11556 ( .A1(n14659), .A2(n9912), .ZN(n9911) );
  INV_X1 U11557 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n9912) );
  NOR2_X1 U11558 ( .A1(n10065), .A2(n14495), .ZN(n10064) );
  INV_X1 U11559 ( .A(n13634), .ZN(n10065) );
  NAND2_X1 U11560 ( .A1(n9917), .A2(n9915), .ZN(n11248) );
  INV_X1 U11561 ( .A(n11258), .ZN(n9917) );
  NAND2_X1 U11562 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n9916) );
  INV_X1 U11563 ( .A(n10830), .ZN(n10835) );
  NOR2_X2 U11564 ( .A1(n11254), .A2(n9909), .ZN(n11253) );
  NAND2_X1 U11565 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n9909) );
  NOR2_X1 U11566 ( .A1(n10070), .A2(n10071), .ZN(n10069) );
  INV_X1 U11567 ( .A(n14515), .ZN(n10070) );
  AND4_X1 U11568 ( .A1(n10502), .A2(n10501), .A3(n10500), .A4(n10499), .ZN(
        n10521) );
  NOR2_X1 U11569 ( .A1(n10719), .A2(n9962), .ZN(n9961) );
  INV_X1 U11570 ( .A(n9964), .ZN(n9962) );
  NAND2_X1 U11571 ( .A1(n10718), .A2(n10717), .ZN(n10719) );
  NAND2_X1 U11572 ( .A1(n14823), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9965) );
  AND2_X1 U11573 ( .A1(n10064), .A2(n10063), .ZN(n10062) );
  INV_X1 U11574 ( .A(n12655), .ZN(n10063) );
  INV_X1 U11575 ( .A(n12606), .ZN(n9959) );
  INV_X1 U11576 ( .A(n10318), .ZN(n11144) );
  AND2_X1 U11577 ( .A1(n10058), .A2(n15875), .ZN(n10057) );
  AND2_X1 U11578 ( .A1(n15898), .A2(n10059), .ZN(n10058) );
  INV_X1 U11579 ( .A(n13239), .ZN(n10059) );
  OR2_X1 U11580 ( .A1(n10836), .A2(n10835), .ZN(n10845) );
  NOR2_X1 U11581 ( .A1(n10052), .A2(n12953), .ZN(n10051) );
  INV_X1 U11582 ( .A(n12628), .ZN(n10052) );
  INV_X1 U11583 ( .A(n13302), .ZN(n10050) );
  OR2_X1 U11584 ( .A1(n10600), .A2(n10599), .ZN(n10895) );
  NAND2_X1 U11585 ( .A1(n9844), .A2(n10821), .ZN(n9791) );
  XNOR2_X1 U11586 ( .A(n10284), .B(n10285), .ZN(n10311) );
  NAND2_X1 U11587 ( .A1(n10311), .A2(n10305), .ZN(n10310) );
  NAND2_X1 U11588 ( .A1(n11584), .A2(n11039), .ZN(n10872) );
  NOR2_X1 U11589 ( .A1(n10869), .A2(n10868), .ZN(n10876) );
  NOR2_X1 U11590 ( .A1(n12859), .A2(n10867), .ZN(n10868) );
  NAND2_X1 U11591 ( .A1(n11302), .A2(n11301), .ZN(n11314) );
  INV_X1 U11592 ( .A(n19592), .ZN(n19194) );
  AND4_X1 U11593 ( .A1(n10135), .A2(n10134), .A3(n10133), .A4(n10132), .ZN(
        n10136) );
  AND2_X1 U11594 ( .A1(n9826), .A2(n9825), .ZN(n15169) );
  NAND2_X1 U11595 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9825) );
  NAND2_X1 U11596 ( .A1(n18591), .A2(n18413), .ZN(n9826) );
  NOR3_X1 U11597 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18434), .ZN(n15102) );
  INV_X1 U11598 ( .A(n16190), .ZN(n9934) );
  NOR2_X1 U11599 ( .A1(n17118), .A2(n15285), .ZN(n16194) );
  OAI21_X1 U11600 ( .B1(n15292), .B2(n15291), .A(n17516), .ZN(n15294) );
  NAND2_X1 U11601 ( .A1(n17532), .A2(n15292), .ZN(n17427) );
  XOR2_X1 U11602 ( .A(n17118), .B(n15285), .Z(n15286) );
  INV_X1 U11603 ( .A(n17125), .ZN(n15351) );
  AOI21_X1 U11604 ( .B1(n13722), .B2(n13721), .A(n13720), .ZN(n15314) );
  OR2_X1 U11605 ( .A1(n20623), .A2(n13333), .ZN(n19708) );
  AND2_X1 U11606 ( .A1(n13098), .A2(n13097), .ZN(n13101) );
  INV_X1 U11607 ( .A(n13838), .ZN(n13897) );
  NOR2_X2 U11608 ( .A1(n13364), .A2(n13363), .ZN(n13393) );
  NAND2_X1 U11609 ( .A1(n12998), .A2(n13337), .ZN(n12896) );
  INV_X1 U11610 ( .A(n13223), .ZN(n12401) );
  AND2_X1 U11611 ( .A1(n13334), .A2(n12373), .ZN(n13934) );
  AND2_X1 U11612 ( .A1(n9985), .A2(n9984), .ZN(n9983) );
  INV_X1 U11613 ( .A(n13956), .ZN(n9984) );
  NAND2_X1 U11614 ( .A1(n14102), .A2(n9985), .ZN(n13969) );
  NAND2_X1 U11615 ( .A1(n14284), .A2(n12580), .ZN(n12581) );
  NOR2_X1 U11616 ( .A1(n12069), .A2(n14078), .ZN(n12084) );
  NOR2_X1 U11617 ( .A1(n11941), .A2(n11940), .ZN(n11958) );
  AOI21_X1 U11618 ( .B1(n12524), .B2(n12093), .A(n11917), .ZN(n13282) );
  NAND2_X1 U11619 ( .A1(n13092), .A2(n11870), .ZN(n13165) );
  AOI21_X1 U11620 ( .B1(n9971), .B2(n12022), .A(n9970), .ZN(n9969) );
  NAND2_X1 U11621 ( .A1(n13225), .A2(n9971), .ZN(n9968) );
  INV_X1 U11622 ( .A(n11870), .ZN(n9970) );
  AND2_X1 U11623 ( .A1(n15422), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13052) );
  NOR2_X1 U11624 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n9807), .ZN(
        n9806) );
  INV_X1 U11625 ( .A(n13792), .ZN(n9807) );
  INV_X1 U11626 ( .A(n13791), .ZN(n9759) );
  INV_X1 U11627 ( .A(n10109), .ZN(n9843) );
  AND2_X1 U11628 ( .A1(n10107), .A2(n9751), .ZN(n9644) );
  NAND2_X1 U11629 ( .A1(n14139), .A2(n13653), .ZN(n14069) );
  NAND2_X1 U11630 ( .A1(n9839), .A2(n9793), .ZN(n12567) );
  INV_X1 U11631 ( .A(n9836), .ZN(n9793) );
  INV_X1 U11632 ( .A(n13538), .ZN(n9839) );
  NOR2_X1 U11633 ( .A1(n15750), .A2(n13394), .ZN(n13402) );
  NAND2_X1 U11634 ( .A1(n15594), .A2(n15592), .ZN(n10099) );
  OR2_X1 U11635 ( .A1(n13170), .A2(n9895), .ZN(n15750) );
  NAND2_X1 U11636 ( .A1(n9896), .A2(n13259), .ZN(n9895) );
  NOR2_X1 U11637 ( .A1(n13169), .A2(n15747), .ZN(n9896) );
  OR2_X1 U11638 ( .A1(n13170), .A2(n9893), .ZN(n15748) );
  NAND2_X1 U11639 ( .A1(n13259), .A2(n9894), .ZN(n9893) );
  INV_X1 U11640 ( .A(n13169), .ZN(n9894) );
  NAND2_X1 U11641 ( .A1(n10101), .A2(n10102), .ZN(n19814) );
  AOI21_X1 U11642 ( .B1(n9638), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10103), 
        .ZN(n10102) );
  INV_X1 U11643 ( .A(n12510), .ZN(n10103) );
  AND2_X1 U11644 ( .A1(n11711), .A2(n11733), .ZN(n9966) );
  AND2_X1 U11645 ( .A1(n12922), .A2(n13000), .ZN(n15388) );
  OR2_X1 U11646 ( .A1(n9635), .A2(n19843), .ZN(n20285) );
  AND2_X1 U11647 ( .A1(n12414), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12454) );
  AND2_X1 U11648 ( .A1(n12453), .A2(n12452), .ZN(n12473) );
  OR2_X1 U11649 ( .A1(n12451), .A2(n12450), .ZN(n12453) );
  AOI21_X1 U11650 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n15763), .A(
        n12449), .ZN(n12456) );
  AOI21_X1 U11651 ( .B1(n12471), .B2(n12448), .A(n12447), .ZN(n12449) );
  AND2_X1 U11652 ( .A1(n12446), .A2(n12445), .ZN(n12447) );
  INV_X1 U11653 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n15763) );
  NAND2_X1 U11654 ( .A1(n10230), .A2(n10245), .ZN(n16096) );
  OR2_X1 U11655 ( .A1(n10716), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10124) );
  OR2_X1 U11656 ( .A1(n10618), .A2(n10897), .ZN(n10714) );
  NAND2_X1 U11657 ( .A1(n10697), .A2(n10042), .ZN(n10709) );
  NOR2_X1 U11658 ( .A1(n18681), .A2(n18682), .ZN(n18664) );
  AND2_X1 U11659 ( .A1(n18852), .A2(n13106), .ZN(n11322) );
  AND2_X1 U11660 ( .A1(n13107), .A2(n13105), .ZN(n13106) );
  NAND2_X1 U11661 ( .A1(n10094), .A2(n10093), .ZN(n10092) );
  AND2_X1 U11662 ( .A1(n12674), .A2(n9738), .ZN(n14467) );
  INV_X1 U11663 ( .A(n12645), .ZN(n10017) );
  OR2_X1 U11664 ( .A1(n14529), .A2(n14528), .ZN(n10094) );
  AND2_X1 U11665 ( .A1(n10082), .A2(n10081), .ZN(n10080) );
  INV_X1 U11666 ( .A(n15817), .ZN(n10081) );
  AND2_X1 U11667 ( .A1(n11016), .A2(n11015), .ZN(n14900) );
  NAND2_X1 U11668 ( .A1(n13443), .A2(n13481), .ZN(n14923) );
  AND2_X1 U11669 ( .A1(n11580), .A2(n11579), .ZN(n12870) );
  NOR2_X1 U11670 ( .A1(n15957), .A2(n11218), .ZN(n10086) );
  AND2_X1 U11671 ( .A1(n12642), .A2(n14464), .ZN(n14516) );
  AND2_X1 U11672 ( .A1(n13550), .A2(n14896), .ZN(n14898) );
  CLKBUF_X1 U11673 ( .A(n11241), .Z(n11242) );
  NOR2_X1 U11674 ( .A1(n11258), .A2(n15917), .ZN(n11260) );
  NOR2_X1 U11675 ( .A1(n13320), .A2(n13319), .ZN(n13321) );
  XNOR2_X1 U11676 ( .A(n10844), .B(n16023), .ZN(n15925) );
  NOR2_X1 U11677 ( .A1(n10845), .A2(n10522), .ZN(n10844) );
  XNOR2_X1 U11678 ( .A(n10608), .B(n16013), .ZN(n12634) );
  OR2_X1 U11679 ( .A1(n14538), .A2(n14539), .ZN(n14536) );
  NAND2_X1 U11680 ( .A1(n10069), .A2(n10068), .ZN(n10067) );
  NOR2_X1 U11681 ( .A1(n12643), .A2(n11265), .ZN(n10068) );
  NAND2_X1 U11682 ( .A1(n10124), .A2(n10714), .ZN(n10740) );
  NOR2_X1 U11683 ( .A1(n9685), .A2(n9714), .ZN(n9960) );
  OR2_X1 U11684 ( .A1(n14679), .A2(n10679), .ZN(n10680) );
  AND2_X1 U11685 ( .A1(n14678), .A2(n10691), .ZN(n10695) );
  INV_X1 U11686 ( .A(n9850), .ZN(n9848) );
  OR2_X1 U11687 ( .A1(n9852), .A2(n9851), .ZN(n9849) );
  NAND2_X1 U11688 ( .A1(n9850), .A2(n14677), .ZN(n9847) );
  NAND2_X1 U11689 ( .A1(n14888), .A2(n14675), .ZN(n14891) );
  NOR2_X1 U11690 ( .A1(n14945), .A2(n14944), .ZN(n14946) );
  AOI21_X1 U11691 ( .B1(n9856), .B2(n9857), .A(n9714), .ZN(n9855) );
  OR2_X1 U11692 ( .A1(n15889), .A2(n9858), .ZN(n9854) );
  NAND2_X1 U11693 ( .A1(n9859), .A2(n9857), .ZN(n14743) );
  NAND2_X1 U11694 ( .A1(n15889), .A2(n9860), .ZN(n9859) );
  AND2_X1 U11695 ( .A1(n12951), .A2(n9719), .ZN(n13185) );
  INV_X1 U11696 ( .A(n15987), .ZN(n10014) );
  NAND2_X1 U11697 ( .A1(n9990), .A2(n9989), .ZN(n9988) );
  NAND2_X1 U11698 ( .A1(n10309), .A2(n10308), .ZN(n10336) );
  INV_X1 U11699 ( .A(n11049), .ZN(n10261) );
  OR2_X1 U11700 ( .A1(n10874), .A2(n10873), .ZN(n12933) );
  XNOR2_X1 U11701 ( .A(n11314), .B(n11312), .ZN(n12849) );
  AOI21_X1 U11702 ( .B1(n12887), .B2(n12886), .A(n11311), .ZN(n12848) );
  AND4_X1 U11703 ( .A1(n10254), .A2(n10253), .A3(n11600), .A4(n11163), .ZN(
        n10244) );
  OR2_X1 U11704 ( .A1(n19581), .A2(n19592), .ZN(n19327) );
  NAND2_X1 U11705 ( .A1(n15025), .A2(n15024), .ZN(n19444) );
  NAND2_X1 U11706 ( .A1(n16115), .A2(n18640), .ZN(n15025) );
  INV_X1 U11707 ( .A(n19444), .ZN(n19171) );
  NAND2_X1 U11708 ( .A1(n16978), .A2(P3_EBX_REG_5__SCAN_IN), .ZN(n16968) );
  NOR4_X1 U11709 ( .A1(n18621), .A2(n16642), .A3(n15455), .A4(n18459), .ZN(
        n13787) );
  NOR2_X1 U11710 ( .A1(n13686), .A2(n13687), .ZN(n15264) );
  NAND2_X1 U11711 ( .A1(n18574), .A2(n18583), .ZN(n9939) );
  NAND2_X1 U11712 ( .A1(n9877), .A2(n9875), .ZN(n17378) );
  NOR2_X1 U11713 ( .A1(n9641), .A2(n9876), .ZN(n9875) );
  INV_X1 U11714 ( .A(n16341), .ZN(n9879) );
  INV_X1 U11715 ( .A(n17625), .ZN(n17583) );
  NOR2_X1 U11716 ( .A1(n17363), .A2(n15301), .ZN(n17313) );
  OAI21_X1 U11717 ( .B1(n17411), .B2(n17668), .A(n15299), .ZN(n15300) );
  NAND2_X1 U11718 ( .A1(n9947), .A2(n20838), .ZN(n9948) );
  NAND2_X1 U11719 ( .A1(n17565), .A2(n9940), .ZN(n9941) );
  NAND2_X1 U11720 ( .A1(n9945), .A2(n9944), .ZN(n9943) );
  INV_X1 U11721 ( .A(n17595), .ZN(n9928) );
  NOR2_X1 U11722 ( .A1(n15311), .A2(n15310), .ZN(n16196) );
  INV_X1 U11723 ( .A(n19715), .ZN(n19695) );
  INV_X1 U11724 ( .A(n14210), .ZN(n14206) );
  AND2_X1 U11725 ( .A1(n15603), .A2(n19812), .ZN(n15600) );
  INV_X1 U11726 ( .A(n14290), .ZN(n19841) );
  AND2_X1 U11727 ( .A1(n15410), .A2(n13052), .ZN(n19817) );
  XNOR2_X1 U11728 ( .A(n14216), .B(n10120), .ZN(n14370) );
  NOR2_X1 U11729 ( .A1(n16100), .A2(n19494), .ZN(n18642) );
  AND2_X1 U11730 ( .A1(n13264), .A2(n9922), .ZN(n14507) );
  NAND2_X1 U11731 ( .A1(n18664), .A2(n18665), .ZN(n9922) );
  NAND2_X1 U11732 ( .A1(n18880), .A2(n13440), .ZN(n10022) );
  NOR2_X1 U11733 ( .A1(n10089), .A2(n10087), .ZN(n11577) );
  AND2_X1 U11734 ( .A1(n14596), .A2(n11585), .ZN(n18880) );
  NOR2_X1 U11735 ( .A1(n14983), .A2(n12841), .ZN(n19261) );
  NAND2_X1 U11736 ( .A1(n9863), .A2(n14671), .ZN(n14717) );
  AOI21_X1 U11737 ( .B1(n14917), .B2(n16057), .A(n14916), .ZN(n9785) );
  NAND2_X1 U11738 ( .A1(n9789), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14927) );
  NAND2_X1 U11739 ( .A1(n9673), .A2(n9790), .ZN(n9789) );
  INV_X1 U11740 ( .A(n15963), .ZN(n9790) );
  NAND2_X1 U11741 ( .A1(n12938), .A2(n14910), .ZN(n14973) );
  AND2_X1 U11742 ( .A1(n11182), .A2(n19617), .ZN(n16063) );
  AND2_X1 U11743 ( .A1(n19581), .A2(n19139), .ZN(n19585) );
  INV_X1 U11744 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19588) );
  NOR2_X1 U11745 ( .A1(n9729), .A2(n9997), .ZN(n11479) );
  AND2_X1 U11746 ( .A1(n10027), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n9997) );
  AOI22_X1 U11747 ( .A1(n10027), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9624), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11485) );
  AOI21_X1 U11748 ( .B1(n11567), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n9735), .ZN(n11406) );
  AOI22_X1 U11749 ( .A1(n10027), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10370), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11411) );
  AND4_X1 U11750 ( .A1(n10579), .A2(n10578), .A3(n10577), .A4(n10576), .ZN(
        n10590) );
  OR2_X1 U11751 ( .A1(n11955), .A2(n11954), .ZN(n12549) );
  OR2_X1 U11752 ( .A1(n11932), .A2(n11931), .ZN(n12535) );
  OR2_X1 U11753 ( .A1(n11907), .A2(n11906), .ZN(n12532) );
  OR2_X1 U11754 ( .A1(n11805), .A2(n11804), .ZN(n12500) );
  NAND2_X1 U11755 ( .A1(n9809), .A2(n11761), .ZN(n12898) );
  NAND2_X1 U11756 ( .A1(n10535), .A2(n10534), .ZN(n10537) );
  NOR2_X1 U11757 ( .A1(n10645), .A2(n10045), .ZN(n10044) );
  AND2_X1 U11758 ( .A1(n10619), .A2(n18858), .ZN(n10633) );
  NOR2_X1 U11759 ( .A1(n9743), .A2(n10002), .ZN(n11544) );
  AND2_X1 U11760 ( .A1(n10027), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10002) );
  AOI21_X1 U11761 ( .B1(n11567), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n9992), .ZN(n11540) );
  AND2_X1 U11762 ( .A1(n10027), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n9992) );
  AOI21_X1 U11763 ( .B1(n10182), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n9744), .ZN(n11539) );
  NOR2_X1 U11764 ( .A1(n9741), .A2(n10000), .ZN(n11506) );
  AND2_X1 U11765 ( .A1(n10027), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10000) );
  NOR2_X1 U11766 ( .A1(n9742), .A2(n10001), .ZN(n11500) );
  AND2_X1 U11767 ( .A1(n10027), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10001) );
  NOR2_X1 U11768 ( .A1(n9727), .A2(n9995), .ZN(n11464) );
  AND2_X1 U11769 ( .A1(n10027), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n9995) );
  NOR2_X1 U11770 ( .A1(n9728), .A2(n9996), .ZN(n11458) );
  AND2_X1 U11771 ( .A1(n10027), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n9996) );
  NOR2_X1 U11772 ( .A1(n9745), .A2(n9993), .ZN(n11443) );
  AND2_X1 U11773 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n9993) );
  NOR2_X1 U11774 ( .A1(n9726), .A2(n9994), .ZN(n11437) );
  AND2_X1 U11775 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n9994) );
  AOI21_X1 U11776 ( .B1(n10318), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10321), .ZN(n10323) );
  AOI21_X1 U11777 ( .B1(n10295), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10317), .ZN(n10322) );
  AND3_X1 U11778 ( .A1(n10210), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10209), .ZN(n10211) );
  AND4_X1 U11779 ( .A1(n10517), .A2(n10516), .A3(n10515), .A4(n10514), .ZN(
        n10519) );
  OR2_X1 U11780 ( .A1(n10493), .A2(n10492), .ZN(n10543) );
  NAND2_X1 U11781 ( .A1(n10238), .A2(n10257), .ZN(n10784) );
  NOR2_X1 U11782 ( .A1(n10338), .A2(n10337), .ZN(n10363) );
  AND2_X1 U11783 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n13765) );
  OR2_X1 U11784 ( .A1(n14000), .A2(n14096), .ZN(n13981) );
  NAND2_X1 U11785 ( .A1(n13546), .A2(n9655), .ZN(n14065) );
  OR2_X1 U11786 ( .A1(n11792), .A2(n11791), .ZN(n12562) );
  AND2_X1 U11787 ( .A1(n11846), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11861) );
  NOR2_X1 U11788 ( .A1(n13853), .A2(n14277), .ZN(n9775) );
  NAND2_X1 U11789 ( .A1(n9903), .A2(n14108), .ZN(n9902) );
  NOR2_X1 U11790 ( .A1(n14013), .A2(n9905), .ZN(n9903) );
  INV_X1 U11791 ( .A(n14118), .ZN(n9905) );
  NOR2_X1 U11792 ( .A1(n9812), .A2(n14437), .ZN(n9811) );
  INV_X1 U11793 ( .A(n12572), .ZN(n9812) );
  NOR2_X1 U11794 ( .A1(n14069), .A2(n13658), .ZN(n9885) );
  OR2_X1 U11795 ( .A1(n15529), .A2(n12574), .ZN(n14326) );
  OR2_X1 U11796 ( .A1(n15529), .A2(n15681), .ZN(n14328) );
  NAND2_X1 U11797 ( .A1(n9769), .A2(n12507), .ZN(n12512) );
  NAND2_X1 U11798 ( .A1(n9766), .A2(n9765), .ZN(n9769) );
  NOR2_X1 U11799 ( .A1(n11837), .A2(n11836), .ZN(n12496) );
  NAND2_X1 U11800 ( .A1(n11827), .A2(n15763), .ZN(n9834) );
  NAND2_X1 U11801 ( .A1(n9833), .A2(n9708), .ZN(n9832) );
  INV_X1 U11802 ( .A(n12496), .ZN(n9833) );
  INV_X1 U11803 ( .A(n11890), .ZN(n9804) );
  INV_X1 U11804 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20148) );
  INV_X1 U11805 ( .A(n11889), .ZN(n13228) );
  INV_X1 U11806 ( .A(n11267), .ZN(n10758) );
  NOR2_X1 U11807 ( .A1(n10701), .A2(n10043), .ZN(n10042) );
  INV_X1 U11808 ( .A(n10698), .ZN(n10043) );
  NOR2_X1 U11809 ( .A1(n10650), .A2(n10048), .ZN(n10047) );
  INV_X1 U11810 ( .A(n10663), .ZN(n10048) );
  NAND2_X1 U11811 ( .A1(n10675), .A2(n10673), .ZN(n10669) );
  AND2_X1 U11812 ( .A1(n10723), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10645) );
  NAND2_X1 U11813 ( .A1(n10633), .A2(n18736), .ZN(n10643) );
  NAND2_X1 U11814 ( .A1(n10641), .A2(n10642), .ZN(n10646) );
  NAND2_X1 U11815 ( .A1(n10612), .A2(n10611), .ZN(n10618) );
  NOR2_X1 U11816 ( .A1(n10555), .A2(n10556), .ZN(n10552) );
  NAND2_X1 U11817 ( .A1(n10552), .A2(n10551), .ZN(n10561) );
  NAND2_X1 U11818 ( .A1(n10293), .A2(n10292), .ZN(n10294) );
  INV_X1 U11819 ( .A(n10291), .ZN(n10292) );
  CLKBUF_X1 U11820 ( .A(n10376), .Z(n11559) );
  NOR2_X1 U11821 ( .A1(n9740), .A2(n9999), .ZN(n11530) );
  AND2_X1 U11822 ( .A1(n10027), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n9999) );
  NOR2_X1 U11823 ( .A1(n9739), .A2(n9998), .ZN(n11524) );
  AND2_X1 U11824 ( .A1(n10027), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n9998) );
  INV_X1 U11825 ( .A(n14481), .ZN(n10019) );
  NAND2_X1 U11826 ( .A1(n9725), .A2(n14546), .ZN(n10077) );
  NAND2_X1 U11827 ( .A1(n10079), .A2(n9725), .ZN(n10078) );
  NAND2_X1 U11828 ( .A1(n10011), .A2(n10010), .ZN(n10009) );
  NOR2_X1 U11829 ( .A1(n12658), .A2(n14900), .ZN(n10010) );
  INV_X1 U11830 ( .A(n10012), .ZN(n10011) );
  NAND2_X1 U11831 ( .A1(n14499), .A2(n13614), .ZN(n10012) );
  INV_X1 U11832 ( .A(n15820), .ZN(n10083) );
  AND2_X1 U11833 ( .A1(n11336), .A2(n13475), .ZN(n10076) );
  NOR2_X1 U11834 ( .A1(n15775), .A2(n9914), .ZN(n9913) );
  INV_X1 U11835 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9914) );
  NOR2_X1 U11836 ( .A1(n10056), .A2(n14726), .ZN(n10055) );
  INV_X1 U11837 ( .A(n13476), .ZN(n10056) );
  INV_X1 U11838 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n9918) );
  INV_X1 U11839 ( .A(n10328), .ZN(n10329) );
  OR2_X1 U11840 ( .A1(n10445), .A2(n10446), .ZN(n10870) );
  NOR2_X1 U11841 ( .A1(n10096), .A2(n14779), .ZN(n10095) );
  INV_X1 U11842 ( .A(n10097), .ZN(n10096) );
  NOR2_X1 U11843 ( .A1(n14804), .A2(n14817), .ZN(n10097) );
  OR2_X1 U11844 ( .A1(n14488), .A2(n10522), .ZN(n10730) );
  NAND2_X1 U11845 ( .A1(n10708), .A2(n14830), .ZN(n9964) );
  AOI21_X1 U11846 ( .B1(n9853), .B2(n9639), .A(n14676), .ZN(n9852) );
  NAND2_X1 U11847 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12603) );
  NOR2_X1 U11848 ( .A1(n14943), .A2(n14957), .ZN(n9869) );
  INV_X1 U11849 ( .A(n9860), .ZN(n9856) );
  AND2_X1 U11850 ( .A1(n10632), .A2(n9861), .ZN(n9860) );
  INV_X1 U11851 ( .A(n15881), .ZN(n9861) );
  XNOR2_X1 U11852 ( .A(n10845), .B(n10737), .ZN(n10843) );
  NAND2_X1 U11853 ( .A1(n10838), .A2(n10829), .ZN(n9784) );
  INV_X1 U11854 ( .A(n11017), .ZN(n11044) );
  INV_X1 U11855 ( .A(n13154), .ZN(n9989) );
  OR2_X1 U11856 ( .A1(n10384), .A2(n10383), .ZN(n10882) );
  NAND2_X1 U11857 ( .A1(n10387), .A2(n10386), .ZN(n10549) );
  NAND2_X1 U11858 ( .A1(n10448), .A2(n10447), .ZN(n10548) );
  OAI21_X1 U11859 ( .B1(n10812), .B2(n10737), .A(n13267), .ZN(n10564) );
  NAND2_X1 U11860 ( .A1(n10283), .A2(n10282), .ZN(n10307) );
  INV_X1 U11861 ( .A(n10281), .ZN(n10282) );
  OR2_X1 U11862 ( .A1(n10862), .A2(n10861), .ZN(n10867) );
  CLKBUF_X1 U11863 ( .A(n11049), .Z(n14979) );
  NAND2_X1 U11864 ( .A1(n12756), .A2(n10363), .ZN(n10344) );
  NAND2_X1 U11865 ( .A1(n19613), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10746) );
  NAND2_X1 U11866 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13688) );
  NAND2_X1 U11867 ( .A1(n15303), .A2(n9660), .ZN(n9925) );
  NOR2_X1 U11868 ( .A1(n17411), .A2(n17397), .ZN(n17356) );
  OAI21_X1 U11869 ( .B1(n16194), .B2(n16195), .A(n17516), .ZN(n15287) );
  NOR2_X1 U11870 ( .A1(n15354), .A2(n17562), .ZN(n15356) );
  AND2_X1 U11871 ( .A1(n15337), .A2(n15279), .ZN(n15281) );
  NOR2_X1 U11872 ( .A1(n18402), .A2(n15146), .ZN(n15160) );
  NAND2_X1 U11873 ( .A1(n18632), .A2(n16307), .ZN(n15325) );
  AOI211_X1 U11874 ( .C1(n13727), .C2(n13726), .A(n15314), .B(n15171), .ZN(
        n16126) );
  NAND2_X1 U11875 ( .A1(n12462), .A2(n9618), .ZN(n12785) );
  NOR2_X1 U11876 ( .A1(n14099), .A2(n14001), .ZN(n14003) );
  AND2_X1 U11877 ( .A1(n14003), .A2(n13987), .ZN(n13985) );
  INV_X1 U11878 ( .A(n11844), .ZN(n14147) );
  NAND2_X1 U11879 ( .A1(n12547), .A2(n12093), .ZN(n11974) );
  AND2_X1 U11880 ( .A1(n13927), .A2(n12397), .ZN(n12398) );
  OR2_X1 U11881 ( .A1(n14241), .A2(n13331), .ZN(n12332) );
  AND2_X1 U11882 ( .A1(n12276), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12285) );
  NAND2_X1 U11883 ( .A1(n12285), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12328) );
  OR2_X1 U11884 ( .A1(n14103), .A2(n13981), .ZN(n13998) );
  NOR2_X1 U11885 ( .A1(n12275), .A2(n15471), .ZN(n12305) );
  NAND2_X1 U11886 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n12305), .ZN(
        n12304) );
  OR2_X1 U11887 ( .A1(n14103), .A2(n14096), .ZN(n14094) );
  AND2_X1 U11888 ( .A1(n12216), .A2(n12215), .ZN(n14104) );
  INV_X1 U11889 ( .A(n13980), .ZN(n14103) );
  NAND2_X1 U11890 ( .A1(n9659), .A2(n9977), .ZN(n9976) );
  INV_X1 U11891 ( .A(n14115), .ZN(n9977) );
  AND2_X1 U11892 ( .A1(n12163), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12164) );
  XNOR2_X1 U11893 ( .A(n15529), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14293) );
  OR2_X1 U11894 ( .A1(n12119), .A2(n12118), .ZN(n12132) );
  NAND2_X1 U11895 ( .A1(n12102), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12119) );
  AND2_X1 U11896 ( .A1(n12084), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12102) );
  CLKBUF_X1 U11897 ( .A(n13639), .Z(n13640) );
  OR2_X1 U11898 ( .A1(n12053), .A2(n12039), .ZN(n12069) );
  AND2_X1 U11899 ( .A1(n9982), .A2(n12068), .ZN(n9981) );
  OR2_X1 U11900 ( .A1(n9655), .A2(n9709), .ZN(n9982) );
  AND2_X1 U11901 ( .A1(n12024), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12025) );
  NOR2_X1 U11902 ( .A1(n12019), .A2(n12018), .ZN(n12024) );
  INV_X1 U11903 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12018) );
  AND2_X1 U11904 ( .A1(n13546), .A2(n13565), .ZN(n13621) );
  OR2_X1 U11905 ( .A1(n11989), .A2(n13502), .ZN(n12019) );
  AND4_X1 U11906 ( .A1(n11988), .A2(n11987), .A3(n11986), .A4(n11985), .ZN(
        n13494) );
  AOI21_X1 U11907 ( .B1(n12542), .B2(n12093), .A(n11962), .ZN(n13363) );
  AOI21_X1 U11908 ( .B1(n12531), .B2(n12093), .A(n11945), .ZN(n13276) );
  INV_X1 U11909 ( .A(n13282), .ZN(n11918) );
  INV_X1 U11910 ( .A(n13089), .ZN(n11868) );
  INV_X1 U11911 ( .A(n13899), .ZN(n9891) );
  XNOR2_X1 U11912 ( .A(n9891), .B(n9888), .ZN(n9887) );
  INV_X1 U11913 ( .A(n13896), .ZN(n9888) );
  NOR3_X1 U11914 ( .A1(n13959), .A2(n13937), .A3(n13952), .ZN(n13938) );
  NAND2_X1 U11915 ( .A1(n13985), .A2(n13971), .ZN(n13973) );
  OR2_X1 U11916 ( .A1(n13973), .A2(n13957), .ZN(n13959) );
  NAND2_X1 U11917 ( .A1(n14257), .A2(n9776), .ZN(n14236) );
  AND2_X1 U11918 ( .A1(n14275), .A2(n9775), .ZN(n9778) );
  NAND2_X1 U11919 ( .A1(n9842), .A2(n10107), .ZN(n15431) );
  NOR2_X1 U11920 ( .A1(n14126), .A2(n9901), .ZN(n14116) );
  INV_X1 U11921 ( .A(n9903), .ZN(n9901) );
  OR2_X1 U11922 ( .A1(n14124), .A2(n14123), .ZN(n14126) );
  NOR2_X1 U11923 ( .A1(n14126), .A2(n14013), .ZN(n14119) );
  NAND2_X1 U11924 ( .A1(n9883), .A2(n9882), .ZN(n14124) );
  INV_X1 U11925 ( .A(n14033), .ZN(n9882) );
  INV_X1 U11926 ( .A(n14043), .ZN(n9883) );
  OR2_X1 U11927 ( .A1(n15529), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15551) );
  NAND2_X1 U11928 ( .A1(n14059), .A2(n14044), .ZN(n14043) );
  AND2_X1 U11929 ( .A1(n9885), .A2(n9884), .ZN(n14059) );
  INV_X1 U11930 ( .A(n14056), .ZN(n9884) );
  OR2_X1 U11931 ( .A1(n14316), .A2(n14300), .ZN(n14303) );
  INV_X1 U11932 ( .A(n9885), .ZN(n14057) );
  AND2_X1 U11933 ( .A1(n13084), .A2(n13083), .ZN(n14423) );
  AND2_X1 U11934 ( .A1(n13500), .A2(n9650), .ZN(n14139) );
  NOR2_X1 U11935 ( .A1(n15674), .A2(n13253), .ZN(n15672) );
  INV_X1 U11936 ( .A(n9799), .ZN(n9798) );
  NAND2_X1 U11937 ( .A1(n13500), .A2(n9897), .ZN(n15710) );
  NAND2_X1 U11938 ( .A1(n13500), .A2(n13499), .ZN(n15708) );
  AND2_X1 U11939 ( .A1(n13400), .A2(n13399), .ZN(n13401) );
  AND2_X1 U11940 ( .A1(n13402), .A2(n13401), .ZN(n13500) );
  AND3_X1 U11941 ( .A1(n13370), .A2(n13648), .A3(n13369), .ZN(n13394) );
  INV_X1 U11942 ( .A(n12523), .ZN(n9764) );
  NAND2_X1 U11943 ( .A1(n13100), .A2(n13099), .ZN(n13170) );
  INV_X1 U11944 ( .A(n9881), .ZN(n13100) );
  NOR2_X1 U11945 ( .A1(n13170), .A2(n13169), .ZN(n13260) );
  INV_X1 U11946 ( .A(n13166), .ZN(n13898) );
  NAND2_X1 U11947 ( .A1(n11752), .A2(n11751), .ZN(n11794) );
  AND2_X2 U11948 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13210) );
  OR2_X1 U11949 ( .A1(n13225), .A2(n11889), .ZN(n20111) );
  AND2_X1 U11950 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20010), .ZN(n19887) );
  OR2_X1 U11951 ( .A1(n13225), .A2(n13228), .ZN(n20382) );
  AOI21_X1 U11952 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20639), .A(n19899), 
        .ZN(n20447) );
  OR2_X1 U11953 ( .A1(n16087), .A2(n16086), .ZN(n16100) );
  AOI221_X1 U11954 ( .B1(n10745), .B2(n12878), .C1(n10745), .C2(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n10744), .ZN(n10779) );
  OAI21_X1 U11955 ( .B1(n10870), .B2(n11267), .A(n10039), .ZN(n10767) );
  NAND2_X1 U11956 ( .A1(n11267), .A2(n10776), .ZN(n10039) );
  OR2_X1 U11957 ( .A1(n10725), .A2(n10724), .ZN(n10735) );
  NAND2_X1 U11958 ( .A1(n10740), .A2(n10720), .ZN(n10725) );
  AND2_X1 U11959 ( .A1(n9664), .A2(n20797), .ZN(n10040) );
  NOR2_X1 U11960 ( .A1(n15805), .A2(n15806), .ZN(n15804) );
  NAND2_X1 U11961 ( .A1(n10659), .A2(n14555), .ZN(n10696) );
  NAND2_X1 U11962 ( .A1(n10696), .A2(n10714), .ZN(n10697) );
  NAND2_X1 U11963 ( .A1(n10664), .A2(n10047), .ZN(n10657) );
  NAND2_X1 U11964 ( .A1(n10032), .A2(n9698), .ZN(n10616) );
  INV_X1 U11965 ( .A(n10618), .ZN(n10032) );
  AND2_X1 U11966 ( .A1(n10723), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10615) );
  NOR2_X1 U11967 ( .A1(n18801), .A2(n18803), .ZN(n18784) );
  NAND2_X1 U11968 ( .A1(n13298), .A2(n18943), .ZN(n18801) );
  NOR2_X1 U11969 ( .A1(n10035), .A2(n10555), .ZN(n10034) );
  NOR2_X1 U11970 ( .A1(n13265), .A2(n15947), .ZN(n13298) );
  CLKBUF_X1 U11971 ( .A(n10285), .Z(n10286) );
  NAND2_X1 U11972 ( .A1(n12952), .A2(n9712), .ZN(n13473) );
  AND2_X1 U11973 ( .A1(n11321), .A2(n18861), .ZN(n13105) );
  AND2_X1 U11974 ( .A1(n11062), .A2(n11061), .ZN(n13304) );
  AOI21_X1 U11975 ( .B1(n9626), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A(n9748), 
        .ZN(n11564) );
  OR2_X1 U11976 ( .A1(n10091), .A2(n14528), .ZN(n10088) );
  OAI21_X1 U11977 ( .B1(n10093), .B2(n10091), .A(n11556), .ZN(n10089) );
  AOI21_X1 U11978 ( .B1(n9626), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A(n9749), .ZN(n11557) );
  AOI22_X1 U11979 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10027), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11558) );
  NAND2_X1 U11980 ( .A1(n12674), .A2(n9724), .ZN(n14569) );
  XNOR2_X1 U11981 ( .A(n11493), .B(n11494), .ZN(n14535) );
  NAND2_X1 U11982 ( .A1(n12674), .A2(n9723), .ZN(n14571) );
  AND2_X1 U11983 ( .A1(n11010), .A2(n11009), .ZN(n14924) );
  NAND2_X1 U11984 ( .A1(n11325), .A2(n10076), .ZN(n18832) );
  INV_X1 U11985 ( .A(n10857), .ZN(n11585) );
  AND3_X1 U11986 ( .A1(n10994), .A2(n10993), .A3(n10992), .ZN(n13441) );
  NAND2_X1 U11987 ( .A1(n11229), .A2(n9913), .ZN(n11262) );
  INV_X1 U11988 ( .A(n10069), .ZN(n10066) );
  CLKBUF_X1 U11989 ( .A(n11231), .Z(n11233) );
  AND2_X1 U11990 ( .A1(n9657), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9910) );
  CLKBUF_X1 U11991 ( .A(n11238), .Z(n11239) );
  NAND2_X1 U11992 ( .A1(n14898), .A2(n10062), .ZN(n12657) );
  NAND2_X1 U11993 ( .A1(n14898), .A2(n13634), .ZN(n14496) );
  NAND2_X1 U11994 ( .A1(n14898), .A2(n10064), .ZN(n14498) );
  NAND2_X1 U11995 ( .A1(n14946), .A2(n10055), .ZN(n14729) );
  NOR2_X1 U11996 ( .A1(n14723), .A2(n9865), .ZN(n9864) );
  INV_X1 U11997 ( .A(n14734), .ZN(n9865) );
  INV_X1 U11998 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11215) );
  INV_X1 U11999 ( .A(n10829), .ZN(n10834) );
  INV_X1 U12000 ( .A(n10823), .ZN(n10824) );
  NOR2_X1 U12001 ( .A1(n13302), .A2(n12953), .ZN(n12954) );
  NOR2_X1 U12002 ( .A1(n11254), .A2(n15958), .ZN(n11256) );
  NAND2_X1 U12003 ( .A1(n10025), .A2(n10024), .ZN(n10023) );
  INV_X1 U12004 ( .A(n14605), .ZN(n10025) );
  INV_X1 U12005 ( .A(n13877), .ZN(n10024) );
  INV_X1 U12006 ( .A(n14759), .ZN(n10007) );
  NAND2_X1 U12007 ( .A1(n10728), .A2(n10727), .ZN(n10026) );
  NOR3_X1 U12008 ( .A1(n15776), .A2(n10522), .A3(n14772), .ZN(n14605) );
  NOR2_X1 U12009 ( .A1(n12641), .A2(n10522), .ZN(n14617) );
  AND2_X1 U12010 ( .A1(n9963), .A2(n9961), .ZN(n14614) );
  AND2_X1 U12011 ( .A1(n14815), .A2(n11191), .ZN(n14788) );
  NAND2_X1 U12012 ( .A1(n15846), .A2(n10097), .ZN(n14640) );
  NAND2_X1 U12013 ( .A1(n10028), .A2(n10732), .ZN(n14635) );
  AND2_X1 U12014 ( .A1(n10730), .A2(n14817), .ZN(n14644) );
  INV_X1 U12015 ( .A(n14644), .ZN(n10717) );
  AND2_X1 U12016 ( .A1(n12670), .A2(n14550), .ZN(n14552) );
  AND2_X1 U12017 ( .A1(n14898), .A2(n9718), .ZN(n12672) );
  INV_X1 U12018 ( .A(n12614), .ZN(n10061) );
  AND2_X1 U12019 ( .A1(n12672), .A2(n12671), .ZN(n12670) );
  NAND2_X1 U12020 ( .A1(n9957), .A2(n9956), .ZN(n14658) );
  AOI21_X1 U12021 ( .B1(n9642), .B2(n9959), .A(n9699), .ZN(n9956) );
  AND2_X1 U12022 ( .A1(n9960), .A2(n9959), .ZN(n9958) );
  OR2_X1 U12023 ( .A1(n12668), .A2(n10522), .ZN(n10704) );
  NAND2_X1 U12024 ( .A1(n9608), .A2(n9869), .ZN(n14912) );
  NAND2_X1 U12025 ( .A1(n14946), .A2(n13476), .ZN(n14727) );
  AND2_X1 U12026 ( .A1(n18718), .A2(n10686), .ZN(n14932) );
  NAND2_X1 U12027 ( .A1(n15899), .A2(n9686), .ZN(n14945) );
  INV_X1 U12028 ( .A(n13408), .ZN(n10060) );
  NAND2_X1 U12029 ( .A1(n15899), .A2(n10057), .ZN(n15873) );
  NAND2_X1 U12030 ( .A1(n9608), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14937) );
  NOR2_X1 U12031 ( .A1(n15906), .A2(n9868), .ZN(n15878) );
  AND2_X1 U12032 ( .A1(n15899), .A2(n10058), .ZN(n15874) );
  NAND2_X1 U12033 ( .A1(n9867), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15896) );
  AND2_X1 U12034 ( .A1(n13321), .A2(n13108), .ZN(n15899) );
  NAND2_X1 U12035 ( .A1(n15899), .A2(n15898), .ZN(n15900) );
  AND2_X1 U12036 ( .A1(n16007), .A2(n11185), .ZN(n15977) );
  NAND2_X1 U12037 ( .A1(n12951), .A2(n9697), .ZN(n15988) );
  AND3_X1 U12038 ( .A1(n10914), .A2(n10913), .A3(n10912), .ZN(n13013) );
  AND2_X1 U12039 ( .A1(n12951), .A2(n10015), .ZN(n13126) );
  INV_X1 U12040 ( .A(n13040), .ZN(n10049) );
  NAND2_X1 U12041 ( .A1(n10050), .A2(n10051), .ZN(n13041) );
  NAND2_X1 U12042 ( .A1(n12951), .A2(n12950), .ZN(n13012) );
  NAND2_X1 U12043 ( .A1(n10895), .A2(n10991), .ZN(n10896) );
  NAND2_X1 U12044 ( .A1(n10550), .A2(n9844), .ZN(n10812) );
  NOR2_X1 U12045 ( .A1(n11162), .A2(n11161), .ZN(n16091) );
  OAI21_X1 U12046 ( .B1(n10854), .B2(n9986), .A(n10856), .ZN(n12857) );
  AND2_X1 U12047 ( .A1(n10872), .A2(n10853), .ZN(n10856) );
  INV_X1 U12048 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10130) );
  CLKBUF_X1 U12049 ( .A(n10795), .Z(n15005) );
  AND3_X1 U12050 ( .A1(n12871), .A2(n12870), .A3(n12869), .ZN(n16085) );
  INV_X1 U12051 ( .A(n19045), .ZN(n19043) );
  OR2_X1 U12052 ( .A1(n19221), .A2(n19249), .ZN(n19196) );
  NOR2_X1 U12053 ( .A1(n19590), .A2(n19608), .ZN(n19226) );
  INV_X1 U12054 ( .A(n10361), .ZN(n9955) );
  NAND2_X1 U12055 ( .A1(n10136), .A2(n9783), .ZN(n10143) );
  AND4_X1 U12056 ( .A1(n10140), .A2(n10139), .A3(n10138), .A4(n10137), .ZN(
        n10141) );
  NAND2_X1 U12057 ( .A1(n10193), .A2(n9783), .ZN(n10200) );
  NOR3_X2 U12058 ( .A1(n15034), .A2(n19171), .A3(n19598), .ZN(n18978) );
  NOR3_X2 U12059 ( .A1(n19171), .A2(n15033), .A3(n19598), .ZN(n18979) );
  NOR2_X1 U12060 ( .A1(n19327), .A2(n19599), .ZN(n19448) );
  INV_X1 U12061 ( .A(n18978), .ZN(n18984) );
  INV_X1 U12062 ( .A(n18979), .ZN(n18986) );
  NAND2_X1 U12063 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19444), .ZN(n18980) );
  AOI21_X1 U12064 ( .B1(n15314), .B2(n15172), .A(n15171), .ZN(n18424) );
  AOI22_X1 U12065 ( .A1(n16126), .A2(n18428), .B1(n18426), .B2(n16196), .ZN(
        n18449) );
  NOR2_X1 U12066 ( .A1(n16362), .A2(n16361), .ZN(n16360) );
  NOR2_X1 U12067 ( .A1(n16372), .A2(n16371), .ZN(n16370) );
  NOR2_X1 U12068 ( .A1(n17291), .A2(n16391), .ZN(n16390) );
  NOR2_X1 U12069 ( .A1(n17335), .A2(n16433), .ZN(n16432) );
  INV_X1 U12070 ( .A(n17524), .ZN(n16601) );
  NAND2_X1 U12071 ( .A1(n16756), .A2(n9665), .ZN(n16745) );
  NOR2_X1 U12072 ( .A1(n16417), .A2(n9818), .ZN(n9817) );
  INV_X1 U12073 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n9818) );
  NAND2_X1 U12074 ( .A1(n16820), .A2(n9663), .ZN(n9816) );
  NAND2_X1 U12075 ( .A1(n16967), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n16926) );
  AOI21_X1 U12076 ( .B1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n16937), .A(
        n15231), .ZN(n15232) );
  NAND2_X1 U12077 ( .A1(n17283), .A2(n9656), .ZN(n16128) );
  AND2_X1 U12078 ( .A1(n17283), .A2(n9871), .ZN(n16163) );
  AND2_X1 U12079 ( .A1(n9656), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9871) );
  NOR2_X1 U12080 ( .A1(n17260), .A2(n9873), .ZN(n9872) );
  NAND2_X1 U12081 ( .A1(n17283), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17259) );
  NOR2_X1 U12082 ( .A1(n17296), .A2(n17297), .ZN(n17283) );
  NAND2_X1 U12083 ( .A1(n17323), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17296) );
  NOR2_X1 U12084 ( .A1(n17345), .A2(n17346), .ZN(n17323) );
  NOR2_X1 U12085 ( .A1(n17378), .A2(n17380), .ZN(n17366) );
  INV_X1 U12086 ( .A(n17419), .ZN(n9878) );
  NAND2_X1 U12087 ( .A1(n17823), .A2(n17780), .ZN(n17453) );
  NOR2_X1 U12088 ( .A1(n17526), .A2(n16341), .ZN(n17457) );
  AND2_X1 U12089 ( .A1(n17552), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17524) );
  NAND2_X1 U12090 ( .A1(n9870), .A2(n9689), .ZN(n17484) );
  INV_X1 U12091 ( .A(n17584), .ZN(n9870) );
  INV_X1 U12092 ( .A(n17484), .ZN(n17552) );
  NAND2_X1 U12093 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17584) );
  NOR2_X1 U12094 ( .A1(n16172), .A2(n15440), .ZN(n16134) );
  NAND2_X1 U12095 ( .A1(n9934), .A2(n9932), .ZN(n15440) );
  AND2_X1 U12096 ( .A1(n17534), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9932) );
  NAND2_X1 U12097 ( .A1(n17516), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9935) );
  INV_X1 U12098 ( .A(n15292), .ZN(n17517) );
  INV_X1 U12099 ( .A(n9950), .ZN(n9949) );
  OAI21_X1 U12100 ( .B1(n20838), .B2(n17862), .A(n17534), .ZN(n9950) );
  NOR2_X1 U12101 ( .A1(n17517), .A2(n9640), .ZN(n17533) );
  NOR2_X1 U12102 ( .A1(n17876), .A2(n17551), .ZN(n17550) );
  NOR2_X1 U12103 ( .A1(n17614), .A2(n15275), .ZN(n17606) );
  NAND2_X1 U12104 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17623), .ZN(
        n17622) );
  NAND2_X2 U12105 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18434) );
  NOR2_X1 U12106 ( .A1(n13748), .A2(n13747), .ZN(n17981) );
  NOR2_X1 U12107 ( .A1(n13738), .A2(n13737), .ZN(n17985) );
  INV_X1 U12108 ( .A(n15148), .ZN(n17989) );
  INV_X1 U12109 ( .A(n18253), .ZN(n18227) );
  NAND2_X1 U12110 ( .A1(n13384), .A2(n12799), .ZN(n20623) );
  AND2_X1 U12111 ( .A1(n19708), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19721) );
  NAND2_X1 U12112 ( .A1(n13357), .A2(n13355), .ZN(n19709) );
  AND2_X1 U12113 ( .A1(n13357), .A2(n13340), .ZN(n19700) );
  NAND2_X1 U12114 ( .A1(n13357), .A2(n13356), .ZN(n19715) );
  INV_X1 U12115 ( .A(n19700), .ZN(n19718) );
  INV_X1 U12116 ( .A(n14136), .ZN(n19739) );
  INV_X1 U12117 ( .A(n14146), .ZN(n19738) );
  AND2_X1 U12118 ( .A1(n13001), .A2(n13052), .ZN(n19742) );
  NAND2_X1 U12119 ( .A1(n19742), .A2(n14147), .ZN(n14146) );
  INV_X1 U12120 ( .A(n19739), .ZN(n14144) );
  INV_X1 U12121 ( .A(n14177), .ZN(n14197) );
  NAND2_X1 U12122 ( .A1(n12477), .A2(n12476), .ZN(n14210) );
  OR2_X1 U12123 ( .A1(n14206), .A2(n12963), .ZN(n14213) );
  NAND2_X1 U12124 ( .A1(n19779), .A2(n19760), .ZN(n19747) );
  XOR2_X1 U12125 ( .A(n13860), .B(n13859), .Z(n13923) );
  AOI21_X1 U12126 ( .B1(n9980), .B2(n14028), .A(n14027), .ZN(n15556) );
  NAND2_X1 U12127 ( .A1(n14315), .A2(n12572), .ZN(n14331) );
  OR2_X1 U12128 ( .A1(n19817), .A2(n12592), .ZN(n15603) );
  NAND2_X1 U12129 ( .A1(n9889), .A2(n9886), .ZN(n14350) );
  OR2_X1 U12130 ( .A1(n13938), .A2(n9890), .ZN(n9889) );
  NAND2_X1 U12131 ( .A1(n13938), .A2(n9887), .ZN(n9886) );
  XNOR2_X1 U12132 ( .A(n9891), .B(n13821), .ZN(n9890) );
  NAND2_X1 U12133 ( .A1(n9759), .A2(n9806), .ZN(n9805) );
  XNOR2_X1 U12134 ( .A(n13795), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13866) );
  INV_X1 U12135 ( .A(n14223), .ZN(n14265) );
  AND2_X1 U12136 ( .A1(n9842), .A2(n9644), .ZN(n14285) );
  NAND2_X1 U12137 ( .A1(n12567), .A2(n12566), .ZN(n13587) );
  NAND2_X1 U12138 ( .A1(n10099), .A2(n15591), .ZN(n15584) );
  NAND2_X1 U12139 ( .A1(n9762), .A2(n12523), .ZN(n13252) );
  NAND2_X1 U12140 ( .A1(n13246), .A2(n13245), .ZN(n9762) );
  NAND2_X1 U12141 ( .A1(n13081), .A2(n13077), .ZN(n15733) );
  AND2_X1 U12142 ( .A1(n13081), .A2(n13067), .ZN(n19824) );
  INV_X1 U12143 ( .A(n15733), .ZN(n19826) );
  NAND2_X1 U12144 ( .A1(n11860), .A2(n15763), .ZN(n10105) );
  INV_X1 U12145 ( .A(n12499), .ZN(n11849) );
  NOR2_X1 U12146 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20595) );
  OR2_X1 U12147 ( .A1(n20382), .A2(n20252), .ZN(n20449) );
  OAI221_X1 U12148 ( .B1(n20159), .B2(n20294), .C1(n20159), .C2(n20158), .A(
        n20220), .ZN(n20184) );
  OR2_X1 U12149 ( .A1(n20257), .A2(n20328), .ZN(n20246) );
  OR2_X1 U12150 ( .A1(n20382), .A2(n20285), .ZN(n20337) );
  OAI211_X1 U12151 ( .C1(n20389), .C2(n20388), .A(n20387), .B(n20386), .ZN(
        n20428) );
  INV_X1 U12152 ( .A(n20449), .ZN(n20494) );
  AND2_X1 U12153 ( .A1(n15418), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15422) );
  NOR2_X1 U12154 ( .A1(n10735), .A2(n10734), .ZN(n13893) );
  INV_X1 U12155 ( .A(n9907), .ZN(n15774) );
  INV_X1 U12156 ( .A(n15773), .ZN(n9906) );
  INV_X1 U12157 ( .A(n9908), .ZN(n14461) );
  NOR2_X1 U12158 ( .A1(n14475), .A2(n18785), .ZN(n15786) );
  NOR2_X1 U12159 ( .A1(n15804), .A2(n18785), .ZN(n14476) );
  NOR2_X1 U12160 ( .A1(n14476), .A2(n14651), .ZN(n14475) );
  INV_X1 U12161 ( .A(n9607), .ZN(n18694) );
  NOR2_X1 U12162 ( .A1(n14713), .A2(n9920), .ZN(n9919) );
  INV_X1 U12163 ( .A(n18665), .ZN(n9920) );
  NOR2_X1 U12164 ( .A1(n14507), .A2(n14713), .ZN(n14506) );
  INV_X1 U12165 ( .A(n18810), .ZN(n18669) );
  NAND2_X1 U12166 ( .A1(n18715), .A2(n18716), .ZN(n18703) );
  NOR2_X1 U12167 ( .A1(n13525), .A2(n14748), .ZN(n18715) );
  NAND2_X1 U12168 ( .A1(n18726), .A2(n18728), .ZN(n13525) );
  NOR2_X1 U12169 ( .A1(n18739), .A2(n18741), .ZN(n18726) );
  NAND2_X1 U12170 ( .A1(n18784), .A2(n18787), .ZN(n18769) );
  NAND2_X1 U12171 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n9923) );
  NAND2_X1 U12172 ( .A1(n11275), .A2(n13886), .ZN(n18819) );
  INV_X1 U12173 ( .A(n19499), .ZN(n18779) );
  OR2_X1 U12174 ( .A1(n10937), .A2(n10936), .ZN(n18852) );
  OR2_X1 U12175 ( .A1(n10924), .A2(n10923), .ZN(n13107) );
  INV_X1 U12176 ( .A(n18865), .ZN(n18871) );
  NAND2_X1 U12177 ( .A1(n10092), .A2(n14523), .ZN(n13914) );
  AND2_X1 U12178 ( .A1(n14469), .A2(n14468), .ZN(n14775) );
  NOR2_X1 U12179 ( .A1(n14591), .A2(n11430), .ZN(n14547) );
  NOR3_X1 U12180 ( .A1(n14899), .A2(n14900), .A3(n10013), .ZN(n14500) );
  AND2_X1 U12181 ( .A1(n14601), .A2(n14585), .ZN(n18898) );
  NAND2_X1 U12182 ( .A1(n9987), .A2(n9990), .ZN(n13153) );
  INV_X1 U12183 ( .A(n14601), .ZN(n18885) );
  AND2_X1 U12184 ( .A1(n12813), .A2(n19510), .ZN(n18921) );
  BUF_X1 U12185 ( .A(n18904), .Z(n18930) );
  NOR3_X1 U12186 ( .A1(n9734), .A2(n10086), .A3(n10085), .ZN(n10084) );
  INV_X1 U12187 ( .A(n11210), .ZN(n10085) );
  XNOR2_X1 U12188 ( .A(n14514), .B(n11265), .ZN(n14759) );
  OAI21_X1 U12189 ( .B1(n14516), .B2(n14515), .A(n14514), .ZN(n15780) );
  OR2_X1 U12190 ( .A1(n14516), .A2(n14465), .ZN(n14774) );
  NOR2_X1 U12191 ( .A1(n12642), .A2(n12644), .ZN(n14789) );
  INV_X1 U12192 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15917) );
  AND2_X1 U12193 ( .A1(n10073), .A2(n13600), .ZN(n15926) );
  INV_X1 U12194 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13605) );
  INV_X1 U12195 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15958) );
  AND2_X1 U12196 ( .A1(n15957), .A2(n12782), .ZN(n15948) );
  INV_X1 U12197 ( .A(n15941), .ZN(n18939) );
  INV_X1 U12198 ( .A(n18815), .ZN(n12845) );
  INV_X1 U12199 ( .A(n15957), .ZN(n18934) );
  INV_X1 U12200 ( .A(n15942), .ZN(n18936) );
  XNOR2_X1 U12201 ( .A(n11158), .B(n11157), .ZN(n15813) );
  NOR2_X1 U12202 ( .A1(n14536), .A2(n10067), .ZN(n11158) );
  NAND2_X1 U12203 ( .A1(n18876), .A2(n16057), .ZN(n11053) );
  INV_X1 U12204 ( .A(n10851), .ZN(n11054) );
  OAI21_X1 U12205 ( .B1(n11211), .B2(n16060), .A(n11210), .ZN(n10851) );
  INV_X1 U12206 ( .A(n10004), .ZN(n10003) );
  OAI21_X1 U12207 ( .B1(n14757), .B2(n16060), .A(n10005), .ZN(n10004) );
  AOI21_X1 U12208 ( .B1(n10007), .B2(n16045), .A(n10006), .ZN(n10005) );
  NAND2_X1 U12209 ( .A1(n10113), .A2(n14756), .ZN(n10006) );
  AOI21_X1 U12210 ( .B1(n14743), .B2(n9960), .A(n9642), .ZN(n12608) );
  OR2_X1 U12211 ( .A1(n14891), .A2(n9848), .ZN(n9845) );
  NOR2_X1 U12212 ( .A1(n14915), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9787) );
  NAND2_X1 U12213 ( .A1(n14668), .A2(n14734), .ZN(n14724) );
  NOR2_X1 U12214 ( .A1(n11196), .A2(n16011), .ZN(n16000) );
  NOR2_X1 U12215 ( .A1(n16067), .A2(n16068), .ZN(n16039) );
  NOR2_X1 U12216 ( .A1(n12935), .A2(n10877), .ZN(n13140) );
  AND2_X1 U12217 ( .A1(n11182), .A2(n19618), .ZN(n16033) );
  INV_X1 U12218 ( .A(n19261), .ZN(n19608) );
  INV_X1 U12219 ( .A(n19590), .ZN(n19599) );
  INV_X1 U12220 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19596) );
  INV_X1 U12221 ( .A(n19228), .ZN(n19586) );
  NAND2_X1 U12222 ( .A1(n11304), .A2(n11303), .ZN(n14983) );
  NAND2_X1 U12223 ( .A1(n18815), .A2(n11308), .ZN(n11304) );
  NAND2_X1 U12224 ( .A1(n12851), .A2(n12850), .ZN(n19592) );
  INV_X1 U12225 ( .A(n19105), .ZN(n19074) );
  OAI21_X1 U12226 ( .B1(n19085), .B2(n19082), .A(n19081), .ZN(n19102) );
  INV_X1 U12227 ( .A(n19129), .ZN(n19134) );
  OR3_X1 U12228 ( .A1(n19146), .A2(n19171), .A3(n19145), .ZN(n19164) );
  INV_X1 U12229 ( .A(n19217), .ZN(n19221) );
  OAI21_X1 U12230 ( .B1(n19267), .B2(n19282), .A(n19444), .ZN(n19284) );
  INV_X1 U12231 ( .A(n19453), .ZN(n19388) );
  INV_X1 U12232 ( .A(n19450), .ZN(n19404) );
  INV_X1 U12233 ( .A(n19479), .ZN(n19428) );
  OAI21_X1 U12234 ( .B1(n19401), .B2(n19400), .A(n19399), .ZN(n19432) );
  INV_X1 U12235 ( .A(n19386), .ZN(n19430) );
  INV_X1 U12236 ( .A(n19487), .ZN(n19436) );
  OAI22_X1 U12237 ( .A1(n18948), .A2(n18986), .B1(n18947), .B2(n18984), .ZN(
        n19450) );
  OAI22_X1 U12238 ( .A1(n18954), .A2(n18986), .B1(n18953), .B2(n18984), .ZN(
        n19455) );
  INV_X1 U12239 ( .A(n19412), .ZN(n19460) );
  INV_X1 U12240 ( .A(n19416), .ZN(n19465) );
  INV_X1 U12241 ( .A(n19420), .ZN(n19471) );
  OAI22_X1 U12242 ( .A1(n14176), .A2(n18986), .B1(n13674), .B2(n18984), .ZN(
        n20829) );
  OAI22_X1 U12243 ( .A1(n18974), .A2(n18986), .B1(n18973), .B2(n18984), .ZN(
        n19479) );
  AND2_X1 U12244 ( .A1(n19448), .A2(n19261), .ZN(n19488) );
  OAI22_X1 U12245 ( .A1(n18987), .A2(n18986), .B1(n18985), .B2(n18984), .ZN(
        n19487) );
  OR2_X1 U12246 ( .A1(n11280), .A2(n19606), .ZN(n19494) );
  INV_X1 U12247 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19606) );
  NAND2_X1 U12248 ( .A1(n17971), .A2(n18637), .ZN(n18635) );
  INV_X1 U12249 ( .A(n18624), .ZN(n18632) );
  NOR2_X1 U12250 ( .A1(n17309), .A2(n16411), .ZN(n16410) );
  INV_X1 U12251 ( .A(n16687), .ZN(n16666) );
  NOR2_X1 U12252 ( .A1(n17370), .A2(n16451), .ZN(n16450) );
  NAND2_X1 U12253 ( .A1(n16496), .A2(n9880), .ZN(n16451) );
  NAND2_X1 U12254 ( .A1(n16342), .A2(n16463), .ZN(n9880) );
  INV_X1 U12255 ( .A(n16342), .ZN(n16631) );
  NAND2_X1 U12256 ( .A1(n16342), .A2(n16512), .ZN(n16496) );
  AND4_X1 U12257 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_20__SCAN_IN), 
        .A3(n16809), .A4(n16731), .ZN(n16728) );
  NOR2_X1 U12258 ( .A1(n16745), .A2(n16396), .ZN(n16748) );
  NOR2_X1 U12259 ( .A1(n16437), .A2(n16772), .ZN(n16756) );
  OR2_X1 U12260 ( .A1(n9816), .A2(n16783), .ZN(n16772) );
  NOR2_X1 U12261 ( .A1(n17108), .A2(n9815), .ZN(n9814) );
  INV_X1 U12262 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n9815) );
  AND2_X1 U12263 ( .A1(n16820), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n16809) );
  AND2_X1 U12264 ( .A1(n16835), .A2(P3_EBX_REG_18__SCAN_IN), .ZN(n16820) );
  AND2_X1 U12265 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16858), .ZN(n16823) );
  AND2_X1 U12266 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n16823), .ZN(n16835) );
  NOR3_X1 U12267 ( .A1(n16923), .A2(n9820), .A3(n9819), .ZN(n16860) );
  NAND2_X1 U12268 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .ZN(n9819) );
  AND2_X1 U12269 ( .A1(n16860), .A2(P3_EBX_REG_15__SCAN_IN), .ZN(n16858) );
  NOR3_X1 U12270 ( .A1(n16923), .A2(n9820), .A3(n15136), .ZN(n16874) );
  NAND2_X1 U12271 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .ZN(n9820) );
  NOR2_X1 U12272 ( .A1(n16923), .A2(n16562), .ZN(n16878) );
  NAND2_X1 U12273 ( .A1(n16945), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n16923) );
  NOR2_X1 U12274 ( .A1(n16926), .A2(n15134), .ZN(n16945) );
  NOR2_X1 U12275 ( .A1(n16968), .A2(n9822), .ZN(n16967) );
  NAND2_X1 U12276 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .ZN(n9822) );
  NOR3_X1 U12277 ( .A1(n16983), .A2(n13784), .A3(n13785), .ZN(n16978) );
  INV_X1 U12278 ( .A(n17015), .ZN(n17012) );
  NAND2_X1 U12279 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17012), .ZN(n17011) );
  INV_X1 U12280 ( .A(n17029), .ZN(n17025) );
  NAND2_X1 U12281 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17025), .ZN(n17024) );
  NOR2_X1 U12282 ( .A1(n17196), .A2(n17061), .ZN(n17056) );
  NAND2_X1 U12283 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17077), .ZN(n17073) );
  INV_X1 U12284 ( .A(n17046), .ZN(n17072) );
  INV_X1 U12285 ( .A(n16195), .ZN(n17114) );
  NOR2_X1 U12286 ( .A1(n15188), .A2(n15187), .ZN(n17118) );
  INV_X1 U12287 ( .A(n15338), .ZN(n17122) );
  NOR2_X1 U12288 ( .A1(n15248), .A2(n15247), .ZN(n17125) );
  NOR2_X1 U12289 ( .A1(n15222), .A2(n15221), .ZN(n17138) );
  INV_X1 U12290 ( .A(n17140), .ZN(n17137) );
  NAND2_X1 U12291 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17144), .ZN(n17142) );
  NOR2_X1 U12292 ( .A1(n15458), .A2(n17143), .ZN(n17141) );
  NOR2_X1 U12293 ( .A1(n18408), .A2(n15459), .ZN(n17140) );
  CLKBUF_X1 U12294 ( .A(n17175), .Z(n17181) );
  NOR2_X1 U12295 ( .A1(n16145), .A2(n16144), .ZN(n16146) );
  NOR2_X1 U12296 ( .A1(n17526), .A2(n9641), .ZN(n17401) );
  NAND2_X1 U12297 ( .A1(n9877), .A2(n9672), .ZN(n17414) );
  INV_X1 U12298 ( .A(n17461), .ZN(n17482) );
  NOR2_X2 U12299 ( .A1(n17114), .A2(n17628), .ZN(n17535) );
  AND3_X1 U12300 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17561) );
  INV_X1 U12301 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17586) );
  NOR2_X1 U12302 ( .A1(n17585), .A2(n17583), .ZN(n17621) );
  NOR2_X1 U12303 ( .A1(n16308), .A2(n18621), .ZN(n17617) );
  INV_X1 U12304 ( .A(n17617), .ZN(n17628) );
  INV_X1 U12305 ( .A(n17613), .ZN(n17629) );
  INV_X1 U12306 ( .A(n16202), .ZN(n16206) );
  AOI21_X1 U12307 ( .B1(n16199), .B2(n18428), .A(n16198), .ZN(n16200) );
  NAND2_X1 U12308 ( .A1(n9927), .A2(n17303), .ZN(n17282) );
  AND2_X1 U12309 ( .A1(n9927), .A2(n9926), .ZN(n17281) );
  NAND2_X1 U12310 ( .A1(n15303), .A2(n15302), .ZN(n9927) );
  NAND2_X1 U12311 ( .A1(n9938), .A2(n15293), .ZN(n17403) );
  OR2_X1 U12312 ( .A1(n15295), .A2(n17761), .ZN(n9938) );
  OAI21_X1 U12313 ( .B1(n17766), .B2(n17744), .A(n17952), .ZN(n17857) );
  INV_X1 U12314 ( .A(n9941), .ZN(n17555) );
  NAND2_X1 U12315 ( .A1(n9929), .A2(n9931), .ZN(n17596) );
  INV_X1 U12316 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18412) );
  INV_X1 U12317 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18413) );
  INV_X1 U12318 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18420) );
  INV_X1 U12319 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18569) );
  OR2_X1 U12320 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18482), .ZN(n18608) );
  AND2_X1 U12321 ( .A1(n12487), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n19839)
         );
  NAND2_X1 U12323 ( .A1(n14370), .A2(n19817), .ZN(n12601) );
  OAI21_X1 U12324 ( .B1(n14153), .B2(n19841), .A(n12598), .ZN(n12599) );
  OR2_X1 U12325 ( .A1(n14596), .A2(n11599), .ZN(n10021) );
  OAI211_X1 U12326 ( .C1(n14921), .C2(n14920), .A(n9786), .B(n9690), .ZN(
        P2_U3029) );
  NAND2_X1 U12327 ( .A1(n9788), .A2(n9787), .ZN(n9786) );
  CLKBUF_X3 U12328 ( .A(n15048), .Z(n16929) );
  CLKBUF_X3 U12329 ( .A(n15225), .Z(n16913) );
  INV_X1 U12330 ( .A(n15223), .ZN(n16912) );
  NAND2_X1 U12331 ( .A1(n9608), .A2(n9750), .ZN(n9637) );
  AND2_X1 U12332 ( .A1(n11858), .A2(n10104), .ZN(n9638) );
  AND2_X1 U12333 ( .A1(n12952), .A2(n9661), .ZN(n13406) );
  NAND2_X1 U12334 ( .A1(n11236), .A2(n9657), .ZN(n11234) );
  OAI21_X1 U12335 ( .B1(n11827), .B2(n9835), .A(n13216), .ZN(n13187) );
  INV_X2 U12337 ( .A(n11063), .ZN(n11141) );
  AND2_X1 U12338 ( .A1(n10682), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9639) );
  AND2_X1 U12339 ( .A1(n9948), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9640) );
  OAI21_X2 U12340 ( .B1(n10166), .B2(n10165), .A(n10164), .ZN(n10232) );
  INV_X4 U12341 ( .A(n9610), .ZN(n10723) );
  INV_X2 U12342 ( .A(n15236), .ZN(n15053) );
  NAND2_X1 U12343 ( .A1(n9672), .A2(n9878), .ZN(n9641) );
  NAND2_X1 U12344 ( .A1(n10695), .A2(n10694), .ZN(n9642) );
  NOR2_X1 U12345 ( .A1(n9898), .A2(n13628), .ZN(n9643) );
  AND3_X1 U12346 ( .A1(n9680), .A2(n14315), .A3(n12572), .ZN(n9645) );
  AND2_X1 U12347 ( .A1(n9961), .A2(n9681), .ZN(n9646) );
  AND2_X1 U12348 ( .A1(n10609), .A2(n9696), .ZN(n9647) );
  AND2_X1 U12349 ( .A1(n9990), .A2(n9711), .ZN(n9648) );
  AND2_X1 U12350 ( .A1(n10044), .A2(n9732), .ZN(n9649) );
  AND2_X1 U12351 ( .A1(n9643), .A2(n14137), .ZN(n9650) );
  NAND2_X1 U12352 ( .A1(n9847), .A2(n9849), .ZN(n9651) );
  AND2_X1 U12353 ( .A1(n12952), .A2(n11322), .ZN(n9652) );
  INV_X1 U12354 ( .A(n9900), .ZN(n14097) );
  OR2_X1 U12355 ( .A1(n11258), .A2(n9669), .ZN(n9653) );
  INV_X1 U12356 ( .A(n11936), .ZN(n9801) );
  AND2_X1 U12357 ( .A1(n11367), .A2(n9730), .ZN(n9654) );
  NAND2_X1 U12358 ( .A1(n11236), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11235) );
  AND2_X1 U12359 ( .A1(n13565), .A2(n13620), .ZN(n9655) );
  AND2_X1 U12360 ( .A1(n9872), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9656) );
  AND2_X1 U12361 ( .A1(n9911), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9657) );
  AND2_X1 U12362 ( .A1(n10447), .A2(n10386), .ZN(n9658) );
  AND2_X1 U12363 ( .A1(n9979), .A2(n9707), .ZN(n9659) );
  AND2_X1 U12364 ( .A1(n15302), .A2(n17516), .ZN(n9660) );
  AND2_X1 U12365 ( .A1(n11322), .A2(n9705), .ZN(n9661) );
  AND2_X1 U12366 ( .A1(n9913), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9662) );
  NAND2_X1 U12367 ( .A1(n11229), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11227) );
  INV_X1 U12368 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n18640) );
  INV_X1 U12369 ( .A(n10091), .ZN(n10090) );
  OR2_X1 U12370 ( .A1(n13913), .A2(n11550), .ZN(n10091) );
  AND2_X1 U12371 ( .A1(n11182), .A2(n11160), .ZN(n16045) );
  INV_X1 U12372 ( .A(n16045), .ZN(n16055) );
  AND2_X1 U12373 ( .A1(n9814), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n9663) );
  AND2_X1 U12374 ( .A1(n10042), .A2(n10041), .ZN(n9664) );
  AND2_X1 U12375 ( .A1(n9817), .A2(P3_EBX_REG_25__SCAN_IN), .ZN(n9665) );
  AND2_X2 U12376 ( .A1(n12971), .A2(n11400), .ZN(n10414) );
  OR2_X1 U12377 ( .A1(n14468), .A2(n13915), .ZN(n9666) );
  NOR2_X1 U12378 ( .A1(n16689), .A2(n13688), .ZN(n13700) );
  AND2_X2 U12379 ( .A1(n11400), .A2(n10378), .ZN(n10416) );
  INV_X1 U12380 ( .A(n15265), .ZN(n15236) );
  AND4_X1 U12381 ( .A1(n11707), .A2(n11706), .A3(n11705), .A4(n11704), .ZN(
        n9667) );
  NAND2_X1 U12382 ( .A1(n15846), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14638) );
  OR4_X1 U12383 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(n13689), .ZN(n9668) );
  OR2_X1 U12384 ( .A1(n15917), .A2(n9918), .ZN(n9669) );
  INV_X1 U12385 ( .A(n17139), .ZN(n15259) );
  NAND2_X1 U12386 ( .A1(n9978), .A2(n9979), .ZN(n14010) );
  NAND2_X1 U12387 ( .A1(n10610), .A2(n10609), .ZN(n13602) );
  NAND2_X1 U12388 ( .A1(n9963), .A2(n9964), .ZN(n14633) );
  NOR2_X1 U12389 ( .A1(n14038), .A2(n14039), .ZN(n14026) );
  AND2_X1 U12390 ( .A1(n9978), .A2(n9659), .ZN(n9670) );
  NAND2_X1 U12391 ( .A1(n12567), .A2(n10100), .ZN(n14338) );
  NAND2_X1 U12392 ( .A1(n9953), .A2(n9951), .ZN(n15292) );
  AND4_X1 U12393 ( .A1(n11611), .A2(n11610), .A3(n11609), .A4(n11608), .ZN(
        n9671) );
  AND2_X1 U12394 ( .A1(n17416), .A2(n9879), .ZN(n9672) );
  AOI21_X1 U12395 ( .B1(n10026), .B2(n10116), .A(n14613), .ZN(n14603) );
  XNOR2_X1 U12396 ( .A(n10836), .B(n10830), .ZN(n10829) );
  OR2_X1 U12397 ( .A1(n14912), .A2(n16060), .ZN(n9673) );
  XNOR2_X1 U12398 ( .A(n11794), .B(n11793), .ZN(n13236) );
  NAND2_X1 U12399 ( .A1(n9859), .A2(n10640), .ZN(n15868) );
  AND2_X1 U12400 ( .A1(n10841), .A2(n10840), .ZN(n9674) );
  NOR2_X1 U12401 ( .A1(n15278), .A2(n15277), .ZN(n9675) );
  AND2_X1 U12402 ( .A1(n10697), .A2(n9664), .ZN(n9677) );
  INV_X2 U12403 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9783) );
  AND2_X1 U12404 ( .A1(n15889), .A2(n10632), .ZN(n9678) );
  AND2_X1 U12405 ( .A1(n11855), .A2(n11856), .ZN(n9679) );
  AND2_X1 U12406 ( .A1(n14329), .A2(n14324), .ZN(n9680) );
  NAND2_X1 U12407 ( .A1(n12890), .A2(n12892), .ZN(n12891) );
  OR2_X1 U12408 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n14617), .ZN(
        n9681) );
  AND2_X1 U12409 ( .A1(n15846), .A2(n10095), .ZN(n9682) );
  OR2_X2 U12410 ( .A1(n11688), .A2(n11687), .ZN(n19863) );
  AND2_X1 U12411 ( .A1(n12554), .A2(n15591), .ZN(n9683) );
  AND2_X1 U12412 ( .A1(n10008), .A2(n10003), .ZN(n9684) );
  INV_X1 U12413 ( .A(n14038), .ZN(n9978) );
  OR2_X1 U12414 ( .A1(n14677), .A2(n10680), .ZN(n9685) );
  AND2_X1 U12415 ( .A1(n10057), .A2(n10060), .ZN(n9686) );
  AND2_X1 U12416 ( .A1(n9784), .A2(n10074), .ZN(n9687) );
  OR2_X1 U12417 ( .A1(n14891), .A2(n9639), .ZN(n9688) );
  AND2_X1 U12418 ( .A1(n18815), .A2(n10335), .ZN(n10354) );
  AND2_X1 U12419 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9689) );
  NAND2_X1 U12420 ( .A1(n15905), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15906) );
  XNOR2_X1 U12421 ( .A(n10822), .B(n10572), .ZN(n10827) );
  AND2_X1 U12422 ( .A1(n14919), .A2(n9785), .ZN(n9690) );
  NAND2_X1 U12423 ( .A1(n12674), .A2(n14584), .ZN(n14480) );
  INV_X1 U12424 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18574) );
  AND2_X1 U12425 ( .A1(n10051), .A2(n10049), .ZN(n9691) );
  AND2_X1 U12426 ( .A1(n14861), .A2(n14860), .ZN(n9692) );
  AND2_X1 U12427 ( .A1(n12839), .A2(n9610), .ZN(n10991) );
  INV_X1 U12428 ( .A(n10991), .ZN(n9986) );
  NAND2_X1 U12429 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15286), .ZN(
        n9693) );
  INV_X1 U12430 ( .A(n9898), .ZN(n9897) );
  NAND2_X1 U12431 ( .A1(n13499), .A2(n9899), .ZN(n9898) );
  INV_X1 U12432 ( .A(n9858), .ZN(n9857) );
  NAND2_X1 U12433 ( .A1(n10640), .A2(n9706), .ZN(n9858) );
  INV_X1 U12434 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19603) );
  INV_X1 U12435 ( .A(n12557), .ZN(n10104) );
  NAND2_X1 U12436 ( .A1(n12891), .A2(n11318), .ZN(n12952) );
  NOR2_X1 U12437 ( .A1(n14899), .A2(n14900), .ZN(n13613) );
  NAND2_X1 U12438 ( .A1(n11367), .A2(n10126), .ZN(n13612) );
  NAND2_X1 U12439 ( .A1(n11367), .A2(n10082), .ZN(n13669) );
  NOR2_X1 U12440 ( .A1(n13442), .A2(n13441), .ZN(n13443) );
  NOR3_X1 U12441 ( .A1(n11258), .A2(n9669), .A3(n15888), .ZN(n11251) );
  NOR2_X1 U12442 ( .A1(n11245), .A2(n11247), .ZN(n11246) );
  NOR2_X1 U12443 ( .A1(n11243), .A2(n18676), .ZN(n11244) );
  NOR2_X1 U12444 ( .A1(n14923), .A2(n14924), .ZN(n13592) );
  AND2_X1 U12445 ( .A1(n16756), .A2(n9817), .ZN(n9694) );
  AND2_X1 U12446 ( .A1(n16756), .A2(P3_EBX_REG_23__SCAN_IN), .ZN(n9695) );
  NOR2_X1 U12447 ( .A1(n15921), .A2(n15918), .ZN(n9696) );
  AND2_X1 U12448 ( .A1(n10015), .A2(n13127), .ZN(n9697) );
  AND2_X1 U12449 ( .A1(n14946), .A2(n10053), .ZN(n13550) );
  NOR2_X1 U12450 ( .A1(n13183), .A2(n15968), .ZN(n13288) );
  NAND2_X1 U12451 ( .A1(n10897), .A2(n10614), .ZN(n9698) );
  AND3_X1 U12452 ( .A1(n10700), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n10737), .ZN(n9699) );
  AND2_X1 U12453 ( .A1(n10631), .A2(n15908), .ZN(n9700) );
  OR2_X1 U12454 ( .A1(n15529), .A2(n12568), .ZN(n9701) );
  NOR2_X1 U12455 ( .A1(n14593), .A2(n14592), .ZN(n14591) );
  INV_X1 U12456 ( .A(n10812), .ZN(n15949) );
  NOR2_X1 U12457 ( .A1(n14547), .A2(n14546), .ZN(n9702) );
  NOR2_X1 U12458 ( .A1(n10435), .A2(n10434), .ZN(n10863) );
  OR3_X1 U12459 ( .A1(n14899), .A2(n10012), .A3(n14900), .ZN(n9703) );
  AND2_X1 U12460 ( .A1(n9715), .A2(n10034), .ZN(n9704) );
  AND2_X1 U12461 ( .A1(n18845), .A2(n18844), .ZN(n9705) );
  OR2_X1 U12462 ( .A1(n15869), .A2(n15872), .ZN(n9706) );
  AND2_X1 U12463 ( .A1(n14122), .A2(n14011), .ZN(n9707) );
  NOR3_X1 U12464 ( .A1(n14126), .A2(n9902), .A3(n13819), .ZN(n9904) );
  AND2_X1 U12465 ( .A1(n12466), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9708) );
  AND2_X1 U12466 ( .A1(n13565), .A2(n14064), .ZN(n9709) );
  NOR2_X1 U12467 ( .A1(n14126), .A2(n9902), .ZN(n9900) );
  INV_X1 U12468 ( .A(n14681), .ZN(n9851) );
  INV_X1 U12469 ( .A(n14677), .ZN(n9853) );
  OR2_X1 U12470 ( .A1(n10460), .A2(n10459), .ZN(n10887) );
  AND2_X1 U12471 ( .A1(n11861), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9710) );
  AND2_X1 U12472 ( .A1(n9989), .A2(n13159), .ZN(n9711) );
  AND2_X1 U12473 ( .A1(n9661), .A2(n11323), .ZN(n9712) );
  INV_X1 U12474 ( .A(n9892), .ZN(n13951) );
  NOR2_X1 U12475 ( .A1(n13959), .A2(n13952), .ZN(n9892) );
  AND2_X1 U12476 ( .A1(n16820), .A2(n9814), .ZN(n9713) );
  NAND2_X1 U12477 ( .A1(n14744), .A2(n14742), .ZN(n9714) );
  AND2_X1 U12478 ( .A1(n10037), .A2(n10036), .ZN(n9715) );
  AND2_X2 U12479 ( .A1(n10376), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10504) );
  AND2_X1 U12480 ( .A1(n10047), .A2(n10046), .ZN(n9716) );
  AND2_X1 U12481 ( .A1(n9853), .A2(n14681), .ZN(n9717) );
  AND2_X1 U12482 ( .A1(n10062), .A2(n10061), .ZN(n9718) );
  AND2_X1 U12483 ( .A1(n9697), .A2(n10014), .ZN(n9719) );
  AND2_X1 U12484 ( .A1(n9658), .A2(n10887), .ZN(n9720) );
  AND2_X1 U12485 ( .A1(n9938), .A2(n9936), .ZN(n9721) );
  NOR2_X1 U12486 ( .A1(n10877), .A2(n9991), .ZN(n9990) );
  INV_X1 U12487 ( .A(n14585), .ZN(n18884) );
  NAND2_X1 U12488 ( .A1(n11325), .A2(n13475), .ZN(n13474) );
  NOR2_X1 U12489 ( .A1(n12935), .A2(n9988), .ZN(n13155) );
  AND2_X1 U12490 ( .A1(n11236), .A2(n9911), .ZN(n9722) );
  AND2_X1 U12491 ( .A1(n10019), .A2(n14584), .ZN(n9723) );
  AND2_X1 U12492 ( .A1(n9723), .A2(n10018), .ZN(n9724) );
  NAND2_X1 U12493 ( .A1(n11452), .A2(n11451), .ZN(n9725) );
  AND2_X1 U12494 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n9726) );
  AND2_X1 U12495 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n9727)
         );
  AND2_X1 U12496 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n9728) );
  AND2_X1 U12497 ( .A1(n10370), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n9729) );
  INV_X1 U12498 ( .A(n18938), .ZN(n15859) );
  AND2_X1 U12499 ( .A1(n15957), .A2(n11220), .ZN(n18938) );
  AND2_X1 U12500 ( .A1(n10083), .A2(n10126), .ZN(n9730) );
  XNOR2_X1 U12501 ( .A(n12512), .B(n12511), .ZN(n12983) );
  XNOR2_X1 U12502 ( .A(n12859), .B(n10867), .ZN(n12925) );
  XOR2_X1 U12503 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .Z(n9731) );
  NAND2_X1 U12504 ( .A1(n10723), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n9732) );
  INV_X1 U12505 ( .A(n13614), .ZN(n10013) );
  INV_X2 U12506 ( .A(n13264), .ZN(n18785) );
  INV_X1 U12507 ( .A(n10642), .ZN(n10045) );
  AND2_X1 U12508 ( .A1(n13500), .A2(n9643), .ZN(n9733) );
  NOR2_X1 U12509 ( .A1(n18944), .A2(n11226), .ZN(n9734) );
  INV_X1 U12510 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12878) );
  AND2_X1 U12511 ( .A1(n10370), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n9735) );
  INV_X1 U12512 ( .A(n12462), .ZN(n12910) );
  AND2_X1 U12513 ( .A1(n9828), .A2(n11732), .ZN(n12462) );
  OR2_X1 U12514 ( .A1(n16923), .A2(n9820), .ZN(n9736) );
  AND2_X1 U12515 ( .A1(n10076), .A2(n10075), .ZN(n9737) );
  AND2_X1 U12516 ( .A1(n9724), .A2(n10017), .ZN(n9738) );
  INV_X1 U12517 ( .A(n18933), .ZN(n16010) );
  AND2_X1 U12518 ( .A1(n12591), .A2(n20333), .ZN(n14290) );
  NOR2_X1 U12519 ( .A1(n13695), .A2(n13694), .ZN(n18005) );
  INV_X1 U12520 ( .A(n14025), .ZN(n9980) );
  BUF_X1 U12521 ( .A(n11676), .Z(n12465) );
  AND2_X1 U12522 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n9739) );
  AND2_X1 U12523 ( .A1(n10370), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n9740) );
  AND2_X1 U12524 ( .A1(n10370), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n9741) );
  AND2_X1 U12525 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n9742) );
  AND2_X1 U12526 ( .A1(n10370), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n9743) );
  INV_X1 U12527 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11605) );
  AND2_X1 U12528 ( .A1(n10370), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n9744) );
  INV_X1 U12529 ( .A(n13007), .ZN(n13840) );
  AND2_X1 U12530 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n9745)
         );
  AND2_X1 U12531 ( .A1(n17283), .A2(n9872), .ZN(n9746) );
  NAND4_X1 U12532 ( .A1(n12576), .A2(n14428), .A3(n12575), .A4(n14437), .ZN(
        n9747) );
  AND2_X1 U12533 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n9748)
         );
  AND2_X1 U12534 ( .A1(n10370), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n9749) );
  AND2_X1 U12535 ( .A1(n9869), .A2(n12602), .ZN(n9750) );
  AND2_X1 U12536 ( .A1(n15430), .A2(n15638), .ZN(n9751) );
  NAND2_X1 U12537 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n9868) );
  AND2_X1 U12538 ( .A1(n10095), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9752) );
  NAND2_X1 U12539 ( .A1(n17524), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17526) );
  INV_X1 U12540 ( .A(n17526), .ZN(n9877) );
  INV_X1 U12541 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9873) );
  AND2_X1 U12542 ( .A1(n9750), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9753) );
  INV_X1 U12543 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9876) );
  INV_X1 U12544 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9937) );
  INV_X1 U12545 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9874) );
  NAND2_X2 U12546 ( .A1(n18634), .A2(n18566), .ZN(n17861) );
  NOR2_X1 U12547 ( .A1(n19613), .A2(n19111), .ZN(n9754) );
  INV_X1 U12548 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19613) );
  NOR2_X1 U12549 ( .A1(n16701), .A2(n18569), .ZN(n16682) );
  NOR2_X1 U12550 ( .A1(n18423), .A2(n17186), .ZN(n18637) );
  INV_X1 U12551 ( .A(n20353), .ZN(n9755) );
  INV_X1 U12552 ( .A(n9755), .ZN(n9756) );
  INV_X1 U12553 ( .A(n20488), .ZN(n9757) );
  INV_X1 U12554 ( .A(n9757), .ZN(n9758) );
  AOI22_X2 U12555 ( .A1(DATAI_22_), .A2(n9605), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n9606), .ZN(n20364) );
  AOI22_X2 U12556 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n9606), .B1(DATAI_27_), 
        .B2(n9605), .ZN(n20470) );
  AOI22_X2 U12557 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n9606), .B1(DATAI_20_), 
        .B2(n9605), .ZN(n20357) );
  AOI22_X2 U12558 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n9606), .B1(DATAI_24_), 
        .B2(n9605), .ZN(n20453) );
  AOI22_X2 U12559 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n9606), .B1(DATAI_29_), 
        .B2(n9605), .ZN(n20482) );
  AOI22_X2 U12560 ( .A1(DATAI_17_), .A2(n9605), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n9606), .ZN(n20345) );
  AOI22_X2 U12561 ( .A1(DATAI_31_), .A2(n9605), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n9606), .ZN(n20499) );
  NOR3_X4 U12562 ( .A1(n12415), .A2(n14147), .A3(n14206), .ZN(n14200) );
  AOI22_X2 U12563 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n9606), .B1(DATAI_26_), 
        .B2(n9605), .ZN(n20465) );
  NAND2_X1 U12564 ( .A1(n9759), .A2(n13792), .ZN(n9808) );
  AND2_X2 U12565 ( .A1(n11615), .A2(n15389), .ZN(n11699) );
  AND2_X2 U12566 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15389) );
  NAND2_X1 U12567 ( .A1(n9763), .A2(n12523), .ZN(n9761) );
  OAI21_X1 U12568 ( .B1(n9764), .B2(n13246), .A(n9760), .ZN(n12530) );
  XNOR2_X1 U12569 ( .A(n12522), .B(n12517), .ZN(n13246) );
  AND2_X2 U12570 ( .A1(n9766), .A2(n11782), .ZN(n12499) );
  INV_X1 U12571 ( .A(n11782), .ZN(n9768) );
  NAND2_X1 U12572 ( .A1(n9774), .A2(n9771), .ZN(n9770) );
  AND2_X1 U12573 ( .A1(n12513), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n9771) );
  NAND2_X1 U12574 ( .A1(n9773), .A2(n13844), .ZN(n9772) );
  INV_X1 U12575 ( .A(n12513), .ZN(n9773) );
  NAND2_X1 U12576 ( .A1(n12584), .A2(n14276), .ZN(n14223) );
  NOR2_X1 U12577 ( .A1(n9778), .A2(n9777), .ZN(n9776) );
  NAND2_X1 U12578 ( .A1(n12584), .A2(n15529), .ZN(n14257) );
  AOI21_X2 U12579 ( .B1(n12577), .B2(n10107), .A(n9779), .ZN(n14284) );
  OR2_X2 U12580 ( .A1(n9799), .A2(n9797), .ZN(n12577) );
  NAND4_X2 U12581 ( .A1(n18981), .A2(n10232), .A3(n11600), .A4(n9782), .ZN(
        n11167) );
  NAND2_X2 U12582 ( .A1(n9781), .A2(n9780), .ZN(n9782) );
  AND3_X1 U12583 ( .A1(n9782), .A2(n12844), .A3(n10527), .ZN(n10245) );
  INV_X1 U12584 ( .A(n9784), .ZN(n10839) );
  NAND3_X1 U12585 ( .A1(n10073), .A2(n15925), .A3(n13600), .ZN(n9792) );
  NAND3_X1 U12586 ( .A1(n10841), .A2(n10840), .A3(n16012), .ZN(n10073) );
  INV_X1 U12587 ( .A(n19966), .ZN(n9794) );
  XNOR2_X2 U12588 ( .A(n9795), .B(n11819), .ZN(n19966) );
  NAND2_X1 U12589 ( .A1(n11749), .A2(n11748), .ZN(n9795) );
  INV_X1 U12590 ( .A(n11740), .ZN(n11759) );
  AND3_X2 U12591 ( .A1(n9810), .A2(n11675), .A3(n11763), .ZN(n11740) );
  NAND2_X1 U12592 ( .A1(n12571), .A2(n9837), .ZN(n9797) );
  NAND2_X1 U12593 ( .A1(n9798), .A2(n9837), .ZN(n14297) );
  NAND2_X2 U12594 ( .A1(n9804), .A2(n11889), .ZN(n11922) );
  OAI21_X1 U12595 ( .B1(n14216), .B2(n14215), .A(n9805), .ZN(n14217) );
  NAND2_X1 U12596 ( .A1(n9808), .A2(n13794), .ZN(n13795) );
  INV_X1 U12597 ( .A(n9816), .ZN(n16784) );
  INV_X1 U12598 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n9821) );
  NAND4_X1 U12599 ( .A1(n9828), .A2(n11732), .A3(n9731), .A4(n9618), .ZN(n9827) );
  NAND2_X1 U12600 ( .A1(n9827), .A2(n13061), .ZN(n11734) );
  INV_X1 U12601 ( .A(n12504), .ZN(n11732) );
  XNOR2_X2 U12602 ( .A(n11922), .B(n11920), .ZN(n12524) );
  OAI211_X1 U12603 ( .C1(n9835), .C2(n9834), .A(n9832), .B(n9830), .ZN(n11842)
         );
  NAND2_X1 U12604 ( .A1(n9835), .A2(n9831), .ZN(n9830) );
  NOR2_X1 U12605 ( .A1(n11827), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9831) );
  NAND2_X1 U12606 ( .A1(n10100), .A2(n9836), .ZN(n9837) );
  NAND2_X1 U12607 ( .A1(n13538), .A2(n10100), .ZN(n9838) );
  NAND2_X1 U12608 ( .A1(n9842), .A2(n9841), .ZN(n12579) );
  NAND2_X1 U12609 ( .A1(n9840), .A2(n9843), .ZN(n9842) );
  INV_X1 U12610 ( .A(n12577), .ZN(n9840) );
  NAND2_X1 U12611 ( .A1(n10072), .A2(n9844), .ZN(n15950) );
  OAI21_X1 U12612 ( .B1(n14862), .B2(n16037), .A(n9692), .ZN(P2_U3025) );
  NAND2_X1 U12613 ( .A1(n9846), .A2(n9845), .ZN(n14862) );
  AOI21_X1 U12614 ( .B1(n14891), .B2(n9717), .A(n9651), .ZN(n9846) );
  NAND2_X1 U12615 ( .A1(n9854), .A2(n9855), .ZN(n14665) );
  NAND2_X1 U12616 ( .A1(n14668), .A2(n9864), .ZN(n9863) );
  INV_X1 U12617 ( .A(n15906), .ZN(n9867) );
  NAND3_X1 U12618 ( .A1(n16348), .A2(n16349), .A3(n16347), .ZN(P3_U2640) );
  XNOR2_X2 U12619 ( .A(n16127), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16342) );
  NAND2_X1 U12620 ( .A1(n9881), .A2(n13101), .ZN(n13102) );
  NAND2_X1 U12621 ( .A1(n13094), .A2(n13093), .ZN(n9881) );
  NAND3_X1 U12622 ( .A1(n13840), .A2(n13838), .A3(n13002), .ZN(n13006) );
  INV_X1 U12623 ( .A(n9904), .ZN(n14099) );
  AND2_X2 U12624 ( .A1(n9907), .A2(n9906), .ZN(n15772) );
  OR2_X2 U12625 ( .A1(n14460), .A2(n18785), .ZN(n9907) );
  AND2_X2 U12626 ( .A1(n9908), .A2(n11230), .ZN(n14460) );
  OR2_X2 U12627 ( .A1(n12639), .A2(n18785), .ZN(n9908) );
  AOI21_X2 U12628 ( .B1(n18664), .B2(n9919), .A(n9634), .ZN(n14490) );
  NAND2_X1 U12629 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11254) );
  NAND2_X1 U12630 ( .A1(n11253), .A2(n11214), .ZN(n11252) );
  OR2_X2 U12631 ( .A1(n11226), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9921) );
  NAND3_X1 U12632 ( .A1(n15304), .A2(n9925), .A3(n9924), .ZN(n15305) );
  NOR2_X2 U12633 ( .A1(n15280), .A2(n17594), .ZN(n15282) );
  OR2_X1 U12634 ( .A1(n15278), .A2(n9930), .ZN(n9929) );
  OR2_X1 U12635 ( .A1(n15277), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9930) );
  OAI21_X1 U12636 ( .B1(n15278), .B2(n15277), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n9931) );
  AND2_X1 U12637 ( .A1(n9933), .A2(n16190), .ZN(n17271) );
  INV_X1 U12638 ( .A(n17270), .ZN(n9933) );
  NAND2_X1 U12639 ( .A1(n9934), .A2(n16194), .ZN(n16197) );
  OAI22_X2 U12640 ( .A1(n15295), .A2(n9935), .B1(n9936), .B2(n17534), .ZN(
        n17363) );
  INV_X2 U12641 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13689) );
  AOI21_X1 U12642 ( .B1(n17566), .B2(n9946), .A(n9943), .ZN(n9940) );
  AND2_X2 U12643 ( .A1(n9941), .A2(n9693), .ZN(n15288) );
  NAND2_X1 U12644 ( .A1(n9942), .A2(n17565), .ZN(n17557) );
  OAI21_X1 U12645 ( .B1(n17566), .B2(n17567), .A(n9946), .ZN(n9942) );
  NAND2_X1 U12646 ( .A1(n17567), .A2(n9946), .ZN(n9944) );
  INV_X1 U12647 ( .A(n17556), .ZN(n9945) );
  INV_X1 U12648 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9946) );
  OAI211_X2 U12649 ( .C1(n9947), .C2(n17862), .A(n15292), .B(n9949), .ZN(
        n17532) );
  INV_X1 U12651 ( .A(n10360), .ZN(n9954) );
  NAND2_X1 U12652 ( .A1(n14743), .A2(n9958), .ZN(n9957) );
  NAND3_X1 U12653 ( .A1(n10387), .A2(n10448), .A3(n9720), .ZN(n10822) );
  AND2_X1 U12654 ( .A1(n11740), .A2(n11711), .ZN(n12753) );
  INV_X1 U12655 ( .A(n19863), .ZN(n9967) );
  XNOR2_X1 U12656 ( .A(n11842), .B(n11841), .ZN(n9973) );
  NAND2_X1 U12657 ( .A1(n9968), .A2(n9969), .ZN(n13090) );
  XNOR2_X2 U12658 ( .A(n9973), .B(n11843), .ZN(n13225) );
  NAND2_X1 U12659 ( .A1(n13546), .A2(n9981), .ZN(n13638) );
  NAND2_X1 U12660 ( .A1(n14102), .A2(n9983), .ZN(n13943) );
  AND2_X1 U12661 ( .A1(n14102), .A2(n14104), .ZN(n13980) );
  INV_X1 U12662 ( .A(n12935), .ZN(n9987) );
  NAND2_X1 U12663 ( .A1(n9987), .A2(n9648), .ZN(n13158) );
  NAND2_X1 U12664 ( .A1(n14755), .A2(n16057), .ZN(n10008) );
  NOR2_X2 U12665 ( .A1(n14899), .A2(n10009), .ZN(n12610) );
  AOI21_X1 U12666 ( .B1(n14755), .B2(n18884), .A(n10020), .ZN(n11603) );
  NAND3_X1 U12667 ( .A1(n11602), .A2(n10022), .A3(n10021), .ZN(n10020) );
  CLKBUF_X1 U12668 ( .A(n11563), .Z(n10027) );
  AND2_X2 U12669 ( .A1(n10370), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10424) );
  INV_X1 U12670 ( .A(n10711), .ZN(n15794) );
  INV_X1 U12671 ( .A(n14635), .ZN(n10718) );
  INV_X1 U12672 ( .A(n10029), .ZN(n10028) );
  AOI21_X1 U12673 ( .B1(n10711), .B2(n10737), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10029) );
  NAND2_X1 U12674 ( .A1(n10697), .A2(n10040), .ZN(n10716) );
  NAND2_X1 U12675 ( .A1(n10697), .A2(n10698), .ZN(n10702) );
  NAND2_X1 U12676 ( .A1(n10664), .A2(n10663), .ZN(n10666) );
  NAND2_X1 U12677 ( .A1(n10050), .A2(n9691), .ZN(n13320) );
  NOR2_X1 U12678 ( .A1(n14536), .A2(n12643), .ZN(n12642) );
  OR3_X1 U12679 ( .A1(n14536), .A2(n10066), .A3(n12643), .ZN(n14514) );
  INV_X1 U12680 ( .A(n14464), .ZN(n10071) );
  NOR2_X4 U12681 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15004) );
  INV_X1 U12682 ( .A(n10843), .ZN(n10074) );
  NOR2_X1 U12683 ( .A1(n14529), .A2(n10088), .ZN(n10087) );
  INV_X1 U12684 ( .A(n10094), .ZN(n14527) );
  INV_X1 U12685 ( .A(n14522), .ZN(n10093) );
  AND2_X2 U12686 ( .A1(n10098), .A2(n15389), .ZN(n11769) );
  AND2_X2 U12687 ( .A1(n10098), .A2(n11614), .ZN(n11995) );
  NAND2_X1 U12688 ( .A1(n9638), .A2(n13236), .ZN(n10101) );
  INV_X1 U12689 ( .A(n13236), .ZN(n11860) );
  NAND3_X1 U12690 ( .A1(n14276), .A2(n12584), .A3(n12582), .ZN(n12583) );
  NOR2_X1 U12691 ( .A1(n16133), .A2(n17534), .ZN(n16135) );
  INV_X1 U12692 ( .A(n14694), .ZN(n14704) );
  NAND2_X1 U12693 ( .A1(n14694), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14695) );
  AOI21_X1 U12694 ( .B1(n16184), .B2(n17535), .A(n16146), .ZN(n16147) );
  NAND2_X1 U12695 ( .A1(n13304), .A2(n13303), .ZN(n13302) );
  NAND2_X1 U12696 ( .A1(n13639), .A2(n12101), .ZN(n14038) );
  CLKBUF_X1 U12697 ( .A(n11165), .Z(n14452) );
  NAND2_X1 U12698 ( .A1(n11267), .A2(n10258), .ZN(n11165) );
  AND2_X1 U12699 ( .A1(n10159), .A2(n9783), .ZN(n10162) );
  INV_X1 U12700 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10129) );
  NOR2_X1 U12701 ( .A1(n11202), .A2(n11201), .ZN(n11203) );
  INV_X1 U12702 ( .A(n10580), .ZN(n19114) );
  AOI21_X1 U12703 ( .B1(n14221), .B2(n14290), .A(n14220), .ZN(n14222) );
  NAND2_X1 U12704 ( .A1(n11221), .A2(n18938), .ZN(n11222) );
  CLKBUF_X1 U12705 ( .A(n13343), .Z(n20292) );
  NAND2_X1 U12706 ( .A1(n10831), .A2(n10834), .ZN(n10832) );
  AND2_X1 U12707 ( .A1(n11223), .A2(n11222), .ZN(n11224) );
  NAND2_X1 U12708 ( .A1(n10843), .A2(n10839), .ZN(n10840) );
  NAND2_X1 U12709 ( .A1(n15934), .A2(n15935), .ZN(n10838) );
  NAND2_X1 U12710 ( .A1(n14237), .A2(n12585), .ZN(n13791) );
  AND2_X2 U12711 ( .A1(n15905), .A2(n11197), .ZN(n14826) );
  INV_X1 U12712 ( .A(n19332), .ZN(n19323) );
  INV_X1 U12713 ( .A(n13473), .ZN(n11325) );
  OR3_X1 U12714 ( .A1(n13058), .A2(n13057), .A3(n19863), .ZN(n13059) );
  OAI21_X1 U12715 ( .B1(n11153), .B2(n12761), .A(n10290), .ZN(n10291) );
  INV_X1 U12716 ( .A(n10476), .ZN(n19439) );
  INV_X1 U12717 ( .A(n13611), .ZN(n11367) );
  OAI211_X2 U12718 ( .C1(n10838), .C2(n10834), .A(n10833), .B(n10832), .ZN(
        n12632) );
  NOR2_X2 U12719 ( .A1(n10362), .A2(n10361), .ZN(n10474) );
  NAND2_X1 U12720 ( .A1(n13552), .A2(n15823), .ZN(n13611) );
  INV_X1 U12721 ( .A(n15813), .ZN(n11221) );
  OAI21_X1 U12722 ( .B1(n15813), .B2(n16055), .A(n11200), .ZN(n11201) );
  NAND2_X1 U12723 ( .A1(n14535), .A2(n14534), .ZN(n14533) );
  NAND2_X1 U12724 ( .A1(n10220), .A2(n9783), .ZN(n10228) );
  INV_X1 U12725 ( .A(n10855), .ZN(n10852) );
  AND2_X2 U12726 ( .A1(n9626), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10511) );
  AOI22_X1 U12727 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9625), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U12728 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9626), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10140) );
  AOI22_X1 U12729 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9626), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10172) );
  OR2_X1 U12730 ( .A1(n20759), .A2(n15610), .ZN(n10111) );
  AND2_X1 U12731 ( .A1(n14210), .A2(n14147), .ZN(n10112) );
  INV_X1 U12732 ( .A(n9670), .ZN(n14114) );
  INV_X1 U12733 ( .A(n13640), .ZN(n14051) );
  OR3_X1 U12734 ( .A1(n14780), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14758), .ZN(n10113) );
  OR4_X1 U12735 ( .A1(n14780), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14758), .A4(n14761), .ZN(n10114) );
  NOR2_X1 U12736 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13685), .ZN(
        n15191) );
  CLKBUF_X3 U12737 ( .A(n15263), .Z(n16928) );
  AND3_X1 U12738 ( .A1(n10274), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n11169), 
        .ZN(n10115) );
  INV_X1 U12739 ( .A(n10277), .ZN(n11063) );
  NAND2_X1 U12740 ( .A1(n10729), .A2(n20809), .ZN(n10116) );
  AND4_X1 U12741 ( .A1(n15229), .A2(n15228), .A3(n15227), .A4(n15226), .ZN(
        n10117) );
  AND3_X1 U12742 ( .A1(n10184), .A2(n10183), .A3(n9783), .ZN(n10118) );
  OR2_X1 U12743 ( .A1(n16191), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10119) );
  NAND2_X1 U12744 ( .A1(n11919), .A2(n11918), .ZN(n13275) );
  OR2_X1 U12745 ( .A1(n13792), .A2(n14214), .ZN(n10120) );
  AND2_X1 U12746 ( .A1(n16193), .A2(n17870), .ZN(n10121) );
  AND2_X1 U12747 ( .A1(n17185), .A2(n18460), .ZN(n17244) );
  AND2_X1 U12748 ( .A1(n16196), .A2(n16195), .ZN(n10122) );
  INV_X1 U12749 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n16984) );
  XOR2_X1 U12750 ( .A(n10819), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n10123) );
  OR2_X1 U12751 ( .A1(n17516), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10125) );
  OR2_X1 U12752 ( .A1(n11366), .A2(n11365), .ZN(n10126) );
  AND2_X1 U12753 ( .A1(n12610), .A2(n11024), .ZN(n10127) );
  NAND2_X1 U12754 ( .A1(n19868), .A2(n19858), .ZN(n13007) );
  AND2_X1 U12755 ( .A1(n12454), .A2(n12434), .ZN(n12436) );
  NAND2_X1 U12756 ( .A1(n10277), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10293) );
  NOR2_X1 U12757 ( .A1(n11167), .A2(n11166), .ZN(n10263) );
  AND2_X1 U12758 ( .A1(n10269), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10249) );
  NAND2_X1 U12759 ( .A1(n11584), .A2(n10783), .ZN(n10239) );
  AND2_X1 U12760 ( .A1(n20639), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12420) );
  NAND2_X1 U12761 ( .A1(n10723), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10528) );
  INV_X1 U12762 ( .A(n12611), .ZN(n11024) );
  AND2_X2 U12763 ( .A1(n10263), .A2(n10267), .ZN(n10277) );
  AND2_X1 U12764 ( .A1(n10783), .A2(n12844), .ZN(n10259) );
  OR2_X1 U12765 ( .A1(n13721), .A2(n13722), .ZN(n13717) );
  INV_X1 U12766 ( .A(n12415), .ZN(n12503) );
  INV_X1 U12767 ( .A(n14052), .ZN(n12101) );
  OR2_X1 U12768 ( .A1(n11781), .A2(n11780), .ZN(n12501) );
  NAND2_X1 U12769 ( .A1(n11737), .A2(n9629), .ZN(n12414) );
  INV_X1 U12770 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10849) );
  NOR2_X1 U12771 ( .A1(n9639), .A2(n10690), .ZN(n10691) );
  NAND2_X1 U12772 ( .A1(n10547), .A2(n18796), .ZN(n10569) );
  OAI21_X1 U12773 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18583), .A(
        n13717), .ZN(n13718) );
  NAND2_X1 U12774 ( .A1(n9967), .A2(n19868), .ZN(n12504) );
  INV_X1 U12775 ( .A(n12304), .ZN(n12276) );
  NOR2_X2 U12776 ( .A1(n13638), .A2(n13641), .ZN(n13639) );
  INV_X1 U12777 ( .A(n13163), .ZN(n11919) );
  AND2_X1 U12778 ( .A1(n14326), .A2(n14328), .ZN(n14298) );
  OR2_X1 U12779 ( .A1(n11887), .A2(n11886), .ZN(n12519) );
  AND2_X1 U12780 ( .A1(n11317), .A2(n11316), .ZN(n11318) );
  NAND2_X1 U12781 ( .A1(n15014), .A2(n11308), .ZN(n11302) );
  NAND2_X1 U12782 ( .A1(n11493), .A2(n11495), .ZN(n11496) );
  INV_X1 U12783 ( .A(n10158), .ZN(n10165) );
  NOR2_X1 U12784 ( .A1(n14676), .A2(n14887), .ZN(n10694) );
  NAND2_X1 U12785 ( .A1(n18412), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15170) );
  INV_X1 U12786 ( .A(n19709), .ZN(n14015) );
  AND2_X1 U12787 ( .A1(n13657), .A2(n13656), .ZN(n13658) );
  INV_X1 U12788 ( .A(n13101), .ZN(n13099) );
  NAND2_X1 U12789 ( .A1(n13188), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12368) );
  OR2_X1 U12790 ( .A1(n12330), .A2(n13962), .ZN(n12370) );
  NOR2_X1 U12791 ( .A1(n12182), .A2(n15499), .ZN(n12183) );
  AND2_X1 U12792 ( .A1(n12166), .A2(n12165), .ZN(n14011) );
  INV_X1 U12793 ( .A(n13544), .ZN(n12007) );
  INV_X1 U12794 ( .A(n12022), .ZN(n12093) );
  INV_X1 U12795 ( .A(n15583), .ZN(n12554) );
  INV_X1 U12796 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20217) );
  INV_X1 U12797 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20436) );
  OR2_X1 U12798 ( .A1(n10911), .A2(n10910), .ZN(n18860) );
  OR2_X1 U12799 ( .A1(n11474), .A2(n11473), .ZN(n11475) );
  NAND2_X1 U12800 ( .A1(n10226), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10227) );
  INV_X1 U12801 ( .A(n15934), .ZN(n10831) );
  OR2_X1 U12802 ( .A1(n11193), .A2(n10849), .ZN(n11199) );
  AND2_X1 U12803 ( .A1(n18640), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n11308) );
  OR2_X1 U12804 ( .A1(n17187), .A2(n18621), .ZN(n15168) );
  OAI21_X1 U12805 ( .B1(n17256), .B2(n16201), .A(n16200), .ZN(n16202) );
  INV_X1 U12806 ( .A(n15300), .ZN(n15301) );
  INV_X1 U12807 ( .A(n16194), .ZN(n16191) );
  XNOR2_X1 U12808 ( .A(n15347), .B(n15276), .ZN(n17605) );
  INV_X1 U12809 ( .A(n15332), .ZN(n15330) );
  INV_X1 U12810 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13502) );
  AND2_X1 U12811 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11892) );
  AND2_X1 U12812 ( .A1(n19708), .A2(n13339), .ZN(n13357) );
  AND2_X1 U12813 ( .A1(n13832), .A2(n13821), .ZN(n13166) );
  NAND2_X1 U12814 ( .A1(n12183), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12275) );
  NOR2_X1 U12815 ( .A1(n12132), .A2(n14030), .ZN(n12163) );
  INV_X1 U12816 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11971) );
  AND2_X1 U12817 ( .A1(n15424), .A2(n13062), .ZN(n15410) );
  NAND2_X1 U12818 ( .A1(n13793), .A2(n14214), .ZN(n13794) );
  OR2_X1 U12819 ( .A1(n15570), .A2(n15569), .ZN(n15567) );
  INV_X1 U12820 ( .A(n15696), .ZN(n15689) );
  NAND2_X1 U12821 ( .A1(n13060), .A2(n13059), .ZN(n13081) );
  OAI22_X1 U12822 ( .A1(n15769), .A2(n20620), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n20597), .ZN(n20010) );
  INV_X1 U12823 ( .A(n20015), .ZN(n20035) );
  AND2_X1 U12824 ( .A1(n20116), .A2(n20115), .ZN(n20141) );
  INV_X1 U12825 ( .A(n19925), .ZN(n19843) );
  AND2_X1 U12826 ( .A1(n20377), .A2(n20376), .ZN(n20423) );
  INV_X1 U12827 ( .A(n20288), .ZN(n20442) );
  NAND2_X1 U12828 ( .A1(n10792), .A2(n11272), .ZN(n12681) );
  AOI21_X1 U12829 ( .B1(n11155), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11089), .ZN(n13239) );
  NOR2_X1 U12830 ( .A1(n14463), .A2(n10522), .ZN(n14618) );
  OR2_X1 U12831 ( .A1(n14863), .A2(n15978), .ZN(n14878) );
  AND2_X1 U12832 ( .A1(n11179), .A2(n11178), .ZN(n14978) );
  NAND2_X1 U12833 ( .A1(n19581), .A2(n19592), .ZN(n19023) );
  OR2_X1 U12834 ( .A1(n19023), .A2(n19599), .ZN(n19045) );
  OR2_X1 U12835 ( .A1(n19581), .A2(n19194), .ZN(n19228) );
  OR2_X1 U12836 ( .A1(n19590), .A2(n19261), .ZN(n19326) );
  NAND2_X1 U12837 ( .A1(n15168), .A2(n15176), .ZN(n16323) );
  INV_X1 U12838 ( .A(n16686), .ZN(n16698) );
  NAND2_X1 U12839 ( .A1(n10117), .A2(n15232), .ZN(n15238) );
  INV_X1 U12840 ( .A(n17452), .ZN(n16144) );
  INV_X1 U12841 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17443) );
  NAND2_X1 U12842 ( .A1(n17455), .A2(n17625), .ZN(n17365) );
  INV_X1 U12843 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16204) );
  NOR2_X1 U12844 ( .A1(n17564), .A2(n17563), .ZN(n17562) );
  NAND2_X1 U12845 ( .A1(n18624), .A2(n15331), .ZN(n18406) );
  AND2_X1 U12846 ( .A1(n19708), .A2(n13336), .ZN(n19663) );
  NAND2_X1 U12847 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11892), .ZN(
        n11941) );
  AND2_X1 U12848 ( .A1(n19708), .A2(n13344), .ZN(n19703) );
  INV_X1 U12849 ( .A(n19742), .ZN(n14134) );
  OR2_X1 U12850 ( .A1(n13058), .A2(n12464), .ZN(n12477) );
  NAND2_X1 U12851 ( .A1(n12164), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12182) );
  NAND2_X1 U12852 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n12025), .ZN(
        n12053) );
  OR2_X1 U12853 ( .A1(n11968), .A2(n11971), .ZN(n11989) );
  INV_X1 U12854 ( .A(n15603), .ZN(n19813) );
  INV_X1 U12855 ( .A(n14423), .ZN(n15676) );
  INV_X1 U12856 ( .A(n15702), .ZN(n15722) );
  INV_X1 U12857 ( .A(n15674), .ZN(n15720) );
  INV_X1 U12858 ( .A(n20010), .ZN(n19899) );
  NAND2_X1 U12859 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n15424), .ZN(n20597) );
  INV_X1 U12860 ( .A(n20041), .ZN(n20032) );
  INV_X1 U12861 ( .A(n20067), .ZN(n20070) );
  INV_X1 U12862 ( .A(n20187), .ZN(n20178) );
  INV_X1 U12863 ( .A(n20213), .ZN(n20204) );
  OR2_X1 U12864 ( .A1(n9635), .A2(n19925), .ZN(n20328) );
  OR2_X1 U12865 ( .A1(n19842), .A2(n13226), .ZN(n20257) );
  INV_X1 U12866 ( .A(n20337), .ZN(n20368) );
  INV_X1 U12867 ( .A(n20498), .ZN(n20427) );
  INV_X1 U12868 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n15418) );
  INV_X1 U12869 ( .A(n18795), .ZN(n18818) );
  OR2_X1 U12870 ( .A1(n18642), .A2(n11282), .ZN(n18810) );
  INV_X1 U12871 ( .A(n18789), .ZN(n18814) );
  INV_X1 U12872 ( .A(n19494), .ZN(n16106) );
  INV_X1 U12873 ( .A(n14596), .ZN(n18893) );
  INV_X1 U12874 ( .A(n12811), .ZN(n12750) );
  INV_X1 U12875 ( .A(n11595), .ZN(n15034) );
  INV_X1 U12876 ( .A(n11253), .ZN(n11255) );
  AND2_X1 U12877 ( .A1(n13241), .A2(n13240), .ZN(n18742) );
  INV_X1 U12878 ( .A(n15977), .ZN(n15998) );
  AND2_X1 U12880 ( .A1(n11182), .A2(n11052), .ZN(n16057) );
  AND2_X1 U12881 ( .A1(n16090), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16115) );
  OAI21_X1 U12882 ( .B1(n15029), .B2(n15027), .A(n15022), .ZN(n18988) );
  NOR2_X2 U12883 ( .A1(n19023), .A2(n19326), .ZN(n19016) );
  OR2_X1 U12884 ( .A1(n19028), .A2(n19171), .ZN(n20831) );
  INV_X1 U12885 ( .A(n19072), .ZN(n20830) );
  OAI21_X1 U12886 ( .B1(n19085), .B2(n19084), .A(n19083), .ZN(n19101) );
  INV_X1 U12887 ( .A(n19120), .ZN(n19136) );
  AND2_X1 U12888 ( .A1(n19110), .A2(n19581), .ZN(n19163) );
  AND2_X1 U12889 ( .A1(n19585), .A2(n19608), .ZN(n19190) );
  OAI21_X1 U12890 ( .B1(n19220), .B2(n19199), .A(n19444), .ZN(n19223) );
  NOR2_X1 U12891 ( .A1(n19228), .A2(n19326), .ZN(n19249) );
  NOR2_X2 U12892 ( .A1(n19295), .A2(n19261), .ZN(n19318) );
  NAND2_X1 U12893 ( .A1(n19586), .A2(n19590), .ZN(n19295) );
  INV_X1 U12894 ( .A(n19482), .ZN(n19425) );
  NOR2_X1 U12895 ( .A1(n16324), .A2(n16323), .ZN(n18423) );
  INV_X1 U12896 ( .A(n18406), .ZN(n18438) );
  NOR2_X2 U12897 ( .A1(n18635), .A2(n16326), .ZN(n16687) );
  NOR2_X1 U12898 ( .A1(n17210), .A2(n17024), .ZN(n17019) );
  NOR3_X1 U12899 ( .A1(n17108), .A2(n17073), .A3(n17192), .ZN(n17065) );
  NAND2_X1 U12900 ( .A1(n15258), .A2(n15257), .ZN(n16195) );
  INV_X1 U12901 ( .A(n17184), .ZN(n17166) );
  INV_X1 U12902 ( .A(n18621), .ZN(n17188) );
  NOR2_X1 U12903 ( .A1(n17767), .A2(n17446), .ZN(n17694) );
  INV_X1 U12904 ( .A(n17426), .ZN(n17406) );
  INV_X1 U12905 ( .A(n17522), .ZN(n17499) );
  NAND2_X1 U12906 ( .A1(n18399), .A2(n18406), .ZN(n17899) );
  INV_X1 U12907 ( .A(n17453), .ZN(n17807) );
  INV_X1 U12908 ( .A(n17914), .ZN(n17957) );
  INV_X1 U12909 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18468) );
  OR2_X1 U12910 ( .A1(n13058), .A2(n12785), .ZN(n13384) );
  INV_X1 U12911 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20334) );
  INV_X1 U12912 ( .A(n19721), .ZN(n15525) );
  NAND2_X1 U12913 ( .A1(n19742), .A2(n11844), .ZN(n14136) );
  NOR2_X1 U12914 ( .A1(n12492), .A2(n12491), .ZN(n12493) );
  OR2_X1 U12915 ( .A1(n14143), .A2(n14142), .ZN(n15571) );
  OR2_X1 U12916 ( .A1(n19779), .A2(n9630), .ZN(n19743) );
  OR2_X1 U12917 ( .A1(n13058), .A2(n12806), .ZN(n19779) );
  NOR2_X1 U12918 ( .A1(n13384), .A2(n13383), .ZN(n19799) );
  INV_X1 U12919 ( .A(n12599), .ZN(n12600) );
  INV_X1 U12920 ( .A(n15600), .ZN(n15597) );
  INV_X1 U12921 ( .A(n19817), .ZN(n19637) );
  INV_X1 U12922 ( .A(n19824), .ZN(n15685) );
  INV_X1 U12923 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20639) );
  OR2_X1 U12924 ( .A1(n19970), .A2(n20285), .ZN(n19918) );
  OR2_X1 U12925 ( .A1(n19970), .A2(n20328), .ZN(n19962) );
  OR2_X1 U12926 ( .A1(n19970), .A2(n20381), .ZN(n19997) );
  OR2_X1 U12927 ( .A1(n19970), .A2(n20252), .ZN(n20041) );
  OR2_X1 U12928 ( .A1(n20111), .A2(n20285), .ZN(n20067) );
  OR2_X1 U12929 ( .A1(n20111), .A2(n20328), .ZN(n20105) );
  OR2_X1 U12930 ( .A1(n20111), .A2(n20381), .ZN(n20147) );
  OR2_X1 U12931 ( .A1(n20111), .A2(n20252), .ZN(n20187) );
  OR2_X1 U12932 ( .A1(n20257), .A2(n20285), .ZN(n20213) );
  OR2_X1 U12933 ( .A1(n20257), .A2(n20381), .ZN(n20284) );
  OR2_X1 U12934 ( .A1(n20257), .A2(n20252), .ZN(n20327) );
  NAND2_X1 U12935 ( .A1(n20443), .A2(n20329), .ZN(n20431) );
  OR2_X1 U12936 ( .A1(n20382), .A2(n20381), .ZN(n20498) );
  INV_X1 U12937 ( .A(n20587), .ZN(n20583) );
  AND2_X1 U12938 ( .A1(n11287), .A2(n11286), .ZN(n11288) );
  OR2_X1 U12939 ( .A1(n11279), .A2(n11278), .ZN(n18795) );
  OAI21_X2 U12940 ( .B1(n12890), .B2(n12892), .A(n12891), .ZN(n19581) );
  AND2_X1 U12941 ( .A1(n11583), .A2(n16106), .ZN(n14596) );
  OR2_X1 U12942 ( .A1(n18930), .A2(n18921), .ZN(n18923) );
  OR2_X1 U12943 ( .A1(n12688), .A2(n12686), .ZN(n12811) );
  OR2_X1 U12944 ( .A1(n18645), .A2(n12874), .ZN(n15942) );
  INV_X1 U12945 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15888) );
  INV_X1 U12946 ( .A(n15948), .ZN(n18944) );
  NAND2_X1 U12947 ( .A1(n18645), .A2(n11209), .ZN(n15957) );
  INV_X1 U12948 ( .A(n16063), .ZN(n16037) );
  INV_X1 U12949 ( .A(n16057), .ZN(n16053) );
  INV_X1 U12950 ( .A(n16033), .ZN(n16060) );
  NAND2_X1 U12951 ( .A1(n18995), .A2(n19226), .ZN(n20834) );
  NAND2_X1 U12952 ( .A1(n19043), .A2(n19608), .ZN(n19072) );
  NAND2_X1 U12953 ( .A1(n19043), .A2(n19261), .ZN(n19105) );
  INV_X1 U12954 ( .A(n19163), .ZN(n19142) );
  INV_X1 U12955 ( .A(n19190), .ZN(n19188) );
  NAND2_X1 U12956 ( .A1(n19585), .A2(n19261), .ZN(n19217) );
  INV_X1 U12957 ( .A(n19249), .ZN(n19257) );
  NAND2_X1 U12958 ( .A1(n19586), .A2(n19226), .ZN(n19287) );
  OR2_X1 U12959 ( .A1(n19295), .A2(n19608), .ZN(n19354) );
  OR2_X1 U12960 ( .A1(n19581), .A2(n19355), .ZN(n19386) );
  INV_X1 U12961 ( .A(n20829), .ZN(n19424) );
  NAND2_X1 U12962 ( .A1(n19448), .A2(n19608), .ZN(n19492) );
  INV_X1 U12963 ( .A(n16682), .ZN(n16621) );
  INV_X1 U12964 ( .A(n16693), .ZN(n16697) );
  AND2_X1 U12965 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17091), .ZN(n17094) );
  NOR2_X1 U12966 ( .A1(n17142), .A2(n17081), .ZN(n17112) );
  INV_X1 U12967 ( .A(n17141), .ZN(n17132) );
  NOR2_X1 U12968 ( .A1(n17182), .A2(n17166), .ZN(n17175) );
  NAND2_X1 U12969 ( .A1(n17185), .A2(n17147), .ZN(n17184) );
  NAND2_X1 U12970 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17621), .ZN(n17461) );
  NAND2_X1 U12971 ( .A1(n17412), .A2(n17499), .ZN(n17426) );
  INV_X1 U12972 ( .A(n17535), .ZN(n17508) );
  INV_X1 U12973 ( .A(n17616), .ZN(n17608) );
  INV_X1 U12974 ( .A(n17870), .ZN(n17845) );
  INV_X1 U12975 ( .A(n17952), .ZN(n17938) );
  INV_X1 U12976 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18566) );
  INV_X1 U12977 ( .A(n16254), .ZN(n16259) );
  AOI22_X1 U12978 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9626), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10135) );
  AND2_X4 U12979 ( .A1(n14986), .A2(n15019), .ZN(n11563) );
  AND2_X4 U12980 ( .A1(n10378), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10376) );
  AOI22_X1 U12981 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10134) );
  AOI22_X1 U12982 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10370), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10133) );
  AND2_X4 U12983 ( .A1(n10795), .A2(n10131), .ZN(n11566) );
  AND2_X4 U12984 ( .A1(n10795), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10371) );
  AOI22_X1 U12985 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10132) );
  AOI22_X1 U12986 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10139) );
  AOI22_X1 U12987 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9624), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10138) );
  AOI22_X1 U12988 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10137) );
  AOI22_X1 U12989 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10147) );
  AOI22_X1 U12990 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U12991 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10370), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10145) );
  AOI22_X1 U12992 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10144) );
  AOI22_X1 U12993 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U12994 ( .A1(n10376), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10370), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10150) );
  AOI22_X1 U12995 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U12996 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9625), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U12997 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U12998 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10156) );
  AOI22_X1 U12999 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9623), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10155) );
  NAND4_X1 U13000 ( .A1(n10157), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10156), .A4(n10155), .ZN(n10166) );
  AOI22_X1 U13001 ( .A1(n9625), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U13002 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10159) );
  AOI22_X1 U13003 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9624), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10161) );
  AOI22_X1 U13004 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10160) );
  NAND4_X1 U13005 ( .A1(n10163), .A2(n10162), .A3(n10161), .A4(n10160), .ZN(
        n10164) );
  AOI22_X1 U13006 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10370), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10170) );
  AOI22_X1 U13007 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10169) );
  AOI22_X1 U13008 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9625), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10168) );
  AOI22_X1 U13009 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11566), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10167) );
  NAND4_X1 U13010 ( .A1(n10170), .A2(n10169), .A3(n10168), .A4(n10167), .ZN(
        n10176) );
  AOI22_X1 U13011 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9624), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U13012 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10173) );
  AOI22_X1 U13013 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10171) );
  NAND4_X1 U13014 ( .A1(n10174), .A2(n10173), .A3(n10172), .A4(n10171), .ZN(
        n10175) );
  MUX2_X2 U13015 ( .A(n10176), .B(n10175), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12844) );
  AOI22_X1 U13016 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10370), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10179) );
  AOI22_X1 U13017 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10178) );
  AOI22_X1 U13018 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10177) );
  AOI22_X1 U13019 ( .A1(n10221), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9626), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U13020 ( .A1(n10369), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9626), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10186) );
  AOI22_X1 U13021 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9624), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U13022 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U13023 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10183) );
  NAND3_X1 U13024 ( .A1(n10186), .A2(n10185), .A3(n10118), .ZN(n10187) );
  MUX2_X1 U13025 ( .A(n11600), .B(n12844), .S(n10783), .Z(n10203) );
  AOI22_X1 U13026 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9626), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10192) );
  AOI22_X1 U13027 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10191) );
  AOI22_X1 U13028 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10370), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U13029 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10189) );
  NAND4_X1 U13030 ( .A1(n10192), .A2(n10191), .A3(n10190), .A4(n10189), .ZN(
        n10193) );
  AOI22_X1 U13031 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9626), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10197) );
  AOI22_X1 U13032 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U13033 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9624), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10195) );
  AOI22_X1 U13034 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10194) );
  NAND4_X1 U13035 ( .A1(n10197), .A2(n10196), .A3(n10195), .A4(n10194), .ZN(
        n10198) );
  NAND2_X1 U13036 ( .A1(n10198), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10199) );
  OAI21_X1 U13037 ( .B1(n11163), .B2(n10232), .A(n10254), .ZN(n10201) );
  INV_X1 U13038 ( .A(n11584), .ZN(n10864) );
  NAND2_X1 U13039 ( .A1(n10201), .A2(n10864), .ZN(n10202) );
  OAI211_X1 U13040 ( .C1(n18958), .C2(n10245), .A(n10203), .B(n10202), .ZN(
        n11164) );
  AOI22_X1 U13041 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9624), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10207) );
  AOI22_X1 U13042 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10206) );
  AOI22_X1 U13043 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9626), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10205) );
  AOI22_X1 U13044 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10204) );
  NAND2_X1 U13045 ( .A1(n10208), .A2(n9783), .ZN(n10215) );
  AOI22_X1 U13046 ( .A1(n10369), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9626), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10213) );
  AOI22_X1 U13047 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10370), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10212) );
  AOI22_X1 U13048 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10210) );
  AOI22_X1 U13049 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10209) );
  NAND3_X1 U13050 ( .A1(n10213), .A2(n10212), .A3(n10211), .ZN(n10214) );
  INV_X2 U13051 ( .A(n10855), .ZN(n12686) );
  NAND3_X1 U13052 ( .A1(n10864), .A2(n10855), .A3(n11167), .ZN(n10273) );
  AOI22_X1 U13053 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9626), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10219) );
  AOI22_X1 U13054 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10218) );
  AOI22_X1 U13055 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9624), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10217) );
  AOI22_X1 U13056 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10216) );
  NAND4_X1 U13057 ( .A1(n10219), .A2(n10218), .A3(n10217), .A4(n10216), .ZN(
        n10220) );
  AOI22_X1 U13058 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10370), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10225) );
  AOI22_X1 U13059 ( .A1(n11563), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10224) );
  AOI22_X1 U13060 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10371), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10223) );
  AOI22_X1 U13061 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9625), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10222) );
  NAND4_X1 U13062 ( .A1(n10225), .A2(n10224), .A3(n10223), .A4(n10222), .ZN(
        n10226) );
  NAND2_X2 U13063 ( .A1(n10228), .A2(n10227), .ZN(n11272) );
  NOR2_X1 U13064 ( .A1(n11272), .A2(n18640), .ZN(n10229) );
  OAI21_X1 U13065 ( .B1(n11164), .B2(n10273), .A(n10229), .ZN(n10237) );
  AND3_X1 U13066 ( .A1(n11600), .A2(n18958), .A3(n18965), .ZN(n10230) );
  AND2_X1 U13067 ( .A1(n12686), .A2(n18958), .ZN(n10231) );
  NAND2_X1 U13068 ( .A1(n16096), .A2(n10231), .ZN(n11050) );
  INV_X1 U13069 ( .A(n10792), .ZN(n10235) );
  NAND3_X1 U13070 ( .A1(n11050), .A2(n12814), .A3(n10235), .ZN(n10236) );
  AND2_X2 U13071 ( .A1(n10237), .A2(n10236), .ZN(n10279) );
  NAND2_X1 U13072 ( .A1(n11600), .A2(n9610), .ZN(n10238) );
  NAND2_X1 U13073 ( .A1(n10784), .A2(n9782), .ZN(n10240) );
  NAND2_X1 U13074 ( .A1(n10781), .A2(n12844), .ZN(n11175) );
  NAND2_X1 U13075 ( .A1(n11175), .A2(n18965), .ZN(n10242) );
  NAND2_X1 U13076 ( .A1(n10242), .A2(n10241), .ZN(n10274) );
  NAND2_X1 U13077 ( .A1(n10274), .A2(n10267), .ZN(n10243) );
  NAND2_X2 U13078 ( .A1(n10279), .A2(n10243), .ZN(n10295) );
  NAND2_X1 U13079 ( .A1(n10295), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10251) );
  NAND2_X1 U13080 ( .A1(n10855), .A2(n10253), .ZN(n10258) );
  INV_X1 U13081 ( .A(n10258), .ZN(n10246) );
  NAND2_X1 U13082 ( .A1(n10232), .A2(n12844), .ZN(n10857) );
  NOR2_X1 U13083 ( .A1(n10857), .A2(n18971), .ZN(n10248) );
  NAND2_X1 U13084 ( .A1(n11581), .A2(n10248), .ZN(n10252) );
  NOR2_X1 U13085 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10269) );
  AND2_X1 U13086 ( .A1(n10855), .A2(n11272), .ZN(n14454) );
  NAND2_X1 U13087 ( .A1(n10792), .A2(n14454), .ZN(n16108) );
  NAND2_X1 U13088 ( .A1(n10253), .A2(n10254), .ZN(n10256) );
  NAND2_X1 U13089 ( .A1(n11584), .A2(n18965), .ZN(n10255) );
  OAI21_X1 U13090 ( .B1(n10257), .B2(n10256), .A(n10255), .ZN(n10260) );
  NAND2_X2 U13091 ( .A1(n10852), .A2(n11272), .ZN(n11267) );
  NAND3_X1 U13092 ( .A1(n10260), .A2(n11165), .A3(n10259), .ZN(n11049) );
  NAND2_X2 U13093 ( .A1(n10261), .A2(n11168), .ZN(n12973) );
  AOI21_X2 U13094 ( .B1(n10262), .B2(n12973), .A(n18640), .ZN(n10289) );
  INV_X1 U13095 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n12768) );
  NAND2_X1 U13096 ( .A1(n10277), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10265) );
  NAND2_X1 U13097 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10264) );
  OAI211_X1 U13098 ( .C1(n11153), .C2(n12768), .A(n10265), .B(n10264), .ZN(
        n10266) );
  AND2_X1 U13099 ( .A1(n10267), .A2(n11168), .ZN(n10268) );
  OAI22_X1 U13100 ( .A1(n10295), .A2(n10268), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10277), .ZN(n10272) );
  INV_X1 U13101 ( .A(n10269), .ZN(n10316) );
  OAI22_X1 U13102 ( .A1(n12973), .A2(n18640), .B1(n10316), .B2(n19613), .ZN(
        n10270) );
  INV_X1 U13103 ( .A(n10270), .ZN(n10271) );
  NAND2_X1 U13104 ( .A1(n10272), .A2(n10271), .ZN(n10306) );
  AOI21_X1 U13105 ( .B1(n10289), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n10115), .ZN(n10283) );
  INV_X1 U13106 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n10280) );
  NAND2_X1 U13107 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10275) );
  NAND2_X1 U13108 ( .A1(n10316), .A2(n10275), .ZN(n10276) );
  AOI21_X1 U13109 ( .B1(n10277), .B2(P2_EBX_REG_0__SCAN_IN), .A(n10276), .ZN(
        n10278) );
  OAI211_X1 U13110 ( .C1(n11153), .C2(n10280), .A(n10279), .B(n10278), .ZN(
        n10281) );
  INV_X1 U13111 ( .A(n10284), .ZN(n10287) );
  NAND2_X1 U13112 ( .A1(n10287), .A2(n10286), .ZN(n10288) );
  BUF_X2 U13113 ( .A(n10289), .Z(n10318) );
  INV_X1 U13114 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n12761) );
  NAND2_X1 U13115 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10290) );
  INV_X1 U13116 ( .A(n10299), .ZN(n10298) );
  INV_X1 U13117 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n11065) );
  OAI21_X1 U13118 ( .B1(n19596), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11065), 
        .ZN(n10296) );
  INV_X1 U13119 ( .A(n10300), .ZN(n10297) );
  NAND2_X1 U13120 ( .A1(n10298), .A2(n10297), .ZN(n10301) );
  NAND2_X1 U13121 ( .A1(n10300), .A2(n10299), .ZN(n10314) );
  OR2_X2 U13122 ( .A1(n10303), .A2(n10302), .ZN(n10304) );
  NAND2_X2 U13123 ( .A1(n10303), .A2(n10302), .ZN(n10315) );
  INV_X1 U13124 ( .A(n10306), .ZN(n10309) );
  INV_X1 U13125 ( .A(n10307), .ZN(n10308) );
  BUF_X1 U13126 ( .A(n10310), .Z(n10338) );
  INV_X1 U13127 ( .A(n10305), .ZN(n10312) );
  INV_X1 U13128 ( .A(n10311), .ZN(n10335) );
  NAND2_X1 U13129 ( .A1(n10312), .A2(n10335), .ZN(n10313) );
  NAND2_X2 U13130 ( .A1(n10315), .A2(n10314), .ZN(n10330) );
  INV_X1 U13131 ( .A(n10330), .ZN(n10327) );
  NOR2_X1 U13132 ( .A1(n10316), .A2(n19588), .ZN(n10317) );
  INV_X1 U13133 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n16054) );
  NAND2_X1 U13134 ( .A1(n10277), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10320) );
  NAND2_X1 U13135 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10319) );
  OAI211_X1 U13136 ( .C1(n11148), .C2(n16054), .A(n10320), .B(n10319), .ZN(
        n10321) );
  NAND2_X1 U13137 ( .A1(n10322), .A2(n10323), .ZN(n11061) );
  INV_X1 U13138 ( .A(n10322), .ZN(n10325) );
  INV_X1 U13139 ( .A(n10323), .ZN(n10324) );
  NAND2_X1 U13140 ( .A1(n10325), .A2(n10324), .ZN(n10326) );
  NAND2_X2 U13141 ( .A1(n10327), .A2(n10328), .ZN(n10331) );
  NAND2_X4 U13142 ( .A1(n10331), .A2(n11062), .ZN(n11290) );
  INV_X1 U13143 ( .A(n11290), .ZN(n12893) );
  AOI22_X1 U13144 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10467), .B1(
        n19202), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U13145 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10468), .B1(
        n19260), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10348) );
  INV_X1 U13146 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10340) );
  NAND2_X1 U13147 ( .A1(n12756), .A2(n10354), .ZN(n10342) );
  OR2_X1 U13148 ( .A1(n11290), .A2(n10342), .ZN(n10392) );
  INV_X1 U13149 ( .A(n10336), .ZN(n10337) );
  OR2_X2 U13150 ( .A1(n11290), .A2(n10344), .ZN(n19047) );
  INV_X1 U13151 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10339) );
  OAI22_X1 U13152 ( .A1(n10340), .A2(n10392), .B1(n19047), .B2(n10339), .ZN(
        n10341) );
  INV_X1 U13153 ( .A(n10341), .ZN(n10347) );
  INV_X1 U13154 ( .A(n10342), .ZN(n10343) );
  AND2_X1 U13155 ( .A1(n10343), .A2(n11290), .ZN(n19233) );
  INV_X1 U13156 ( .A(n10344), .ZN(n10345) );
  AND2_X2 U13157 ( .A1(n11290), .A2(n10345), .ZN(n19296) );
  AOI22_X1 U13158 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19233), .B1(
        n19296), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10346) );
  AND4_X1 U13159 ( .A1(n10349), .A2(n10348), .A3(n10347), .A4(n10346), .ZN(
        n10368) );
  NAND2_X2 U13160 ( .A1(n10350), .A2(n15014), .ZN(n10362) );
  INV_X1 U13161 ( .A(n10362), .ZN(n10351) );
  INV_X1 U13162 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10353) );
  INV_X1 U13163 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10352) );
  NAND2_X1 U13164 ( .A1(n12845), .A2(n14990), .ZN(n10360) );
  OAI22_X1 U13165 ( .A1(n10580), .A2(n10353), .B1(n10352), .B2(n19397), .ZN(
        n10358) );
  INV_X1 U13166 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10356) );
  NAND2_X1 U13167 ( .A1(n12777), .A2(n12845), .ZN(n10361) );
  INV_X1 U13168 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10355) );
  OAI22_X1 U13169 ( .A1(n10356), .A2(n19332), .B1(n19358), .B2(n10355), .ZN(
        n10357) );
  NOR2_X1 U13170 ( .A1(n10358), .A2(n10357), .ZN(n10367) );
  INV_X1 U13171 ( .A(n10363), .ZN(n10359) );
  NOR2_X2 U13172 ( .A1(n10362), .A2(n10360), .ZN(n10461) );
  AOI22_X1 U13173 ( .A1(n19167), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n10461), .ZN(n10366) );
  AOI22_X1 U13174 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10474), .B1(
        n19439), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10365) );
  NAND4_X1 U13175 ( .A1(n10368), .A2(n10367), .A3(n10366), .A4(n10365), .ZN(
        n10387) );
  AND2_X2 U13176 ( .A1(n11567), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10901) );
  AOI22_X1 U13177 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n10794), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10375) );
  AOI22_X1 U13178 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10449), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10374) );
  AND2_X2 U13179 ( .A1(n10221), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10483) );
  AOI22_X1 U13180 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10373) );
  INV_X1 U13181 ( .A(n10371), .ZN(n11399) );
  NAND2_X1 U13182 ( .A1(n10371), .A2(n9783), .ZN(n12979) );
  AOI22_X1 U13183 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11417), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10372) );
  NAND4_X1 U13184 ( .A1(n10375), .A2(n10374), .A3(n10373), .A4(n10372), .ZN(
        n10384) );
  AND2_X1 U13185 ( .A1(n10376), .A2(n9783), .ZN(n10417) );
  AOI22_X1 U13186 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10417), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10382) );
  AND2_X2 U13187 ( .A1(n11522), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10454) );
  AOI22_X1 U13188 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10429), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U13189 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10415), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U13190 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10413), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10379) );
  NAND4_X1 U13191 ( .A1(n10382), .A2(n10381), .A3(n10380), .A4(n10379), .ZN(
        n10383) );
  INV_X1 U13192 ( .A(n10882), .ZN(n10385) );
  NAND2_X1 U13193 ( .A1(n10385), .A2(n12874), .ZN(n10386) );
  AOI22_X1 U13194 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19233), .B1(
        n19296), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10391) );
  INV_X1 U13195 ( .A(n19047), .ZN(n10469) );
  AOI22_X1 U13196 ( .A1(n10467), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10469), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10390) );
  NAND2_X1 U13197 ( .A1(n10474), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10389) );
  AOI22_X1 U13198 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10468), .B1(
        n19260), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10388) );
  AND4_X1 U13199 ( .A1(n10391), .A2(n10390), .A3(n10389), .A4(n10388), .ZN(
        n10408) );
  INV_X1 U13200 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10395) );
  AOI21_X1 U13201 ( .B1(n18993), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n12874), .ZN(n10394) );
  NAND2_X1 U13202 ( .A1(n19202), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10393) );
  OAI211_X1 U13203 ( .C1(n10396), .C2(n10395), .A(n10394), .B(n10393), .ZN(
        n10397) );
  INV_X1 U13204 ( .A(n10397), .ZN(n10407) );
  INV_X1 U13205 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10400) );
  INV_X1 U13206 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10399) );
  OAI22_X1 U13207 ( .A1(n10400), .A2(n10476), .B1(n19332), .B2(n10399), .ZN(
        n10404) );
  INV_X1 U13208 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10402) );
  INV_X1 U13209 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10401) );
  OAI22_X1 U13210 ( .A1(n10402), .A2(n19397), .B1(n19358), .B2(n10401), .ZN(
        n10403) );
  NOR2_X1 U13211 ( .A1(n10404), .A2(n10403), .ZN(n10405) );
  AOI22_X1 U13212 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10412) );
  AOI22_X1 U13213 ( .A1(n10454), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10411) );
  AOI22_X1 U13214 ( .A1(n10449), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11417), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10410) );
  AOI22_X1 U13215 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10409) );
  NAND4_X1 U13216 ( .A1(n10412), .A2(n10411), .A3(n10410), .A4(n10409), .ZN(
        n10423) );
  AOI22_X1 U13217 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10421) );
  AOI22_X1 U13218 ( .A1(n10415), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10420) );
  AOI22_X1 U13219 ( .A1(n10417), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10419) );
  AOI22_X1 U13220 ( .A1(n10504), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10418) );
  NAND4_X1 U13221 ( .A1(n10421), .A2(n10420), .A3(n10419), .A4(n10418), .ZN(
        n10422) );
  NOR2_X1 U13222 ( .A1(n10423), .A2(n10422), .ZN(n10854) );
  AOI22_X1 U13223 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11416), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10428) );
  AOI22_X1 U13224 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11417), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10427) );
  AOI22_X1 U13225 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10794), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10426) );
  AOI22_X1 U13226 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10417), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10425) );
  NAND4_X1 U13227 ( .A1(n10428), .A2(n10427), .A3(n10426), .A4(n10425), .ZN(
        n10435) );
  AOI22_X1 U13228 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10415), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U13229 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10413), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U13230 ( .A1(n10449), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10431) );
  AOI22_X1 U13231 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10430) );
  NAND4_X1 U13232 ( .A1(n10433), .A2(n10432), .A3(n10431), .A4(n10430), .ZN(
        n10434) );
  NOR2_X1 U13233 ( .A1(n10854), .A2(n10863), .ZN(n10436) );
  NAND2_X1 U13234 ( .A1(n12874), .A2(n10436), .ZN(n10816) );
  AOI22_X1 U13235 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10417), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10440) );
  AOI22_X1 U13236 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10429), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U13237 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10413), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10438) );
  AOI22_X1 U13238 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10415), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10437) );
  NAND4_X1 U13239 ( .A1(n10440), .A2(n10439), .A3(n10438), .A4(n10437), .ZN(
        n10446) );
  AOI22_X1 U13240 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n10483), .B1(
        n10449), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10444) );
  AOI22_X1 U13241 ( .A1(n10901), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U13242 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n10794), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10442) );
  AOI22_X1 U13243 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11417), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10441) );
  NAND4_X1 U13244 ( .A1(n10444), .A2(n10443), .A3(n10442), .A4(n10441), .ZN(
        n10445) );
  NAND2_X1 U13245 ( .A1(n10816), .A2(n10526), .ZN(n10447) );
  AOI22_X1 U13246 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10449), .B1(
        n10794), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10453) );
  AOI22_X1 U13247 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13248 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n10901), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10451) );
  AOI22_X1 U13249 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11417), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10450) );
  NAND4_X1 U13250 ( .A1(n10453), .A2(n10452), .A3(n10451), .A4(n10450), .ZN(
        n10460) );
  AOI22_X1 U13251 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10504), .B1(
        n10417), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U13252 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10429), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U13253 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10413), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U13254 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10415), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10455) );
  NAND4_X1 U13255 ( .A1(n10458), .A2(n10457), .A3(n10456), .A4(n10455), .ZN(
        n10459) );
  INV_X1 U13256 ( .A(n10887), .ZN(n10821) );
  NAND2_X1 U13257 ( .A1(n19167), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10466) );
  NAND2_X1 U13258 ( .A1(n10461), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10465) );
  INV_X1 U13259 ( .A(n19358), .ZN(n10462) );
  NAND2_X1 U13260 ( .A1(n10462), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10464) );
  NAND2_X1 U13261 ( .A1(n19323), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10463) );
  AOI22_X1 U13262 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n10467), .B1(
        n19202), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10473) );
  AOI22_X1 U13263 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19233), .B1(
        n19296), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13264 ( .A1(n10468), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10469), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10471) );
  AOI22_X1 U13265 ( .A1(n19260), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18993), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10470) );
  AOI22_X1 U13266 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n10474), .B1(
        n19114), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10480) );
  INV_X1 U13267 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10477) );
  INV_X1 U13268 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10475) );
  OAI22_X1 U13269 ( .A1(n10477), .A2(n10476), .B1(n19397), .B2(n10475), .ZN(
        n10478) );
  INV_X1 U13270 ( .A(n10478), .ZN(n10479) );
  NAND4_X1 U13271 ( .A1(n10482), .A2(n10481), .A3(n10480), .A4(n10479), .ZN(
        n10496) );
  AOI22_X1 U13272 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13273 ( .A1(n10449), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13274 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13275 ( .A1(n11417), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10484) );
  NAND4_X1 U13276 ( .A1(n10487), .A2(n10486), .A3(n10485), .A4(n10484), .ZN(
        n10493) );
  AOI22_X1 U13277 ( .A1(n10504), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10417), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10491) );
  AOI22_X1 U13278 ( .A1(n10454), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13279 ( .A1(n10415), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U13280 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10488) );
  NAND4_X1 U13281 ( .A1(n10491), .A2(n10490), .A3(n10489), .A4(n10488), .ZN(
        n10492) );
  INV_X1 U13282 ( .A(n10543), .ZN(n10494) );
  NAND2_X1 U13283 ( .A1(n10494), .A2(n12874), .ZN(n10495) );
  NAND2_X1 U13284 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10502) );
  NAND2_X1 U13285 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10501) );
  INV_X1 U13286 ( .A(n10901), .ZN(n10498) );
  INV_X1 U13287 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10497) );
  OR2_X1 U13288 ( .A1(n10498), .A2(n10497), .ZN(n10500) );
  NAND2_X1 U13289 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10499) );
  AOI22_X1 U13290 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10415), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10510) );
  AOI22_X1 U13291 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10413), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10509) );
  INV_X1 U13292 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10503) );
  OR2_X1 U13293 ( .A1(n9617), .A2(n10503), .ZN(n10508) );
  INV_X1 U13294 ( .A(n10504), .ZN(n10506) );
  INV_X1 U13295 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10505) );
  OR2_X1 U13296 ( .A1(n10506), .A2(n10505), .ZN(n10507) );
  AND4_X1 U13297 ( .A1(n10510), .A2(n10509), .A3(n10508), .A4(n10507), .ZN(
        n10520) );
  NAND2_X1 U13298 ( .A1(n10449), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10517) );
  INV_X1 U13299 ( .A(n10511), .ZN(n10513) );
  INV_X1 U13300 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10512) );
  OR2_X1 U13301 ( .A1(n10513), .A2(n10512), .ZN(n10516) );
  NAND2_X1 U13302 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10515) );
  NAND2_X1 U13303 ( .A1(n10454), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10514) );
  AOI22_X1 U13304 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11417), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10518) );
  NAND4_X1 U13305 ( .A1(n10521), .A2(n10520), .A3(n10519), .A4(n10518), .ZN(
        n10613) );
  INV_X1 U13306 ( .A(n10613), .ZN(n10522) );
  NAND2_X1 U13307 ( .A1(n10827), .A2(n10522), .ZN(n10547) );
  MUX2_X1 U13308 ( .A(n19603), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n10766) );
  INV_X1 U13309 ( .A(n10746), .ZN(n10523) );
  NAND2_X1 U13310 ( .A1(n10766), .A2(n10523), .ZN(n10525) );
  NAND2_X1 U13311 ( .A1(n19603), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10524) );
  NAND2_X1 U13312 ( .A1(n10525), .A2(n10524), .ZN(n10533) );
  XNOR2_X1 U13313 ( .A(n15019), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10532) );
  XNOR2_X1 U13314 ( .A(n10533), .B(n10532), .ZN(n10776) );
  INV_X1 U13315 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n10530) );
  INV_X1 U13316 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n12846) );
  NAND2_X1 U13317 ( .A1(n10530), .A2(n12846), .ZN(n10531) );
  MUX2_X1 U13318 ( .A(n10863), .B(n10531), .S(n10723), .Z(n10556) );
  NAND2_X1 U13319 ( .A1(n10533), .A2(n10532), .ZN(n10535) );
  NAND2_X1 U13320 ( .A1(n19596), .A2(n15019), .ZN(n10534) );
  XNOR2_X1 U13321 ( .A(n9783), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10538) );
  XNOR2_X1 U13322 ( .A(n10537), .B(n10538), .ZN(n10757) );
  MUX2_X1 U13323 ( .A(n10882), .B(n10757), .S(n11267), .Z(n10769) );
  INV_X1 U13324 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10536) );
  MUX2_X1 U13325 ( .A(n10769), .B(n10536), .S(n10723), .Z(n10551) );
  NAND3_X1 U13326 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10745), .A3(
        n12878), .ZN(n10754) );
  INV_X1 U13327 ( .A(n10754), .ZN(n10541) );
  NAND2_X1 U13328 ( .A1(n10541), .A2(n11267), .ZN(n10770) );
  OAI21_X1 U13329 ( .B1(n11267), .B2(n10887), .A(n10770), .ZN(n10542) );
  MUX2_X1 U13330 ( .A(n10542), .B(P2_EBX_REG_4__SCAN_IN), .S(n10723), .Z(
        n10560) );
  NAND2_X1 U13331 ( .A1(n9610), .A2(n10543), .ZN(n10891) );
  INV_X1 U13332 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n18797) );
  NAND2_X1 U13333 ( .A1(n10723), .A2(n18797), .ZN(n10544) );
  NAND2_X1 U13334 ( .A1(n10891), .A2(n10544), .ZN(n10545) );
  NOR2_X1 U13335 ( .A1(n9704), .A2(n10545), .ZN(n10546) );
  OR2_X1 U13336 ( .A1(n10612), .A2(n10546), .ZN(n18796) );
  INV_X1 U13337 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16043) );
  XNOR2_X1 U13338 ( .A(n10569), .B(n16043), .ZN(n15931) );
  NAND2_X1 U13339 ( .A1(n10549), .A2(n10548), .ZN(n10550) );
  INV_X2 U13340 ( .A(n10522), .ZN(n10737) );
  OAI21_X1 U13341 ( .B1(n10552), .B2(n10551), .A(n10561), .ZN(n13267) );
  INV_X1 U13342 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16067) );
  XNOR2_X1 U13343 ( .A(n10564), .B(n16067), .ZN(n15951) );
  INV_X1 U13344 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14992) );
  OAI21_X1 U13345 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19613), .A(
        n10746), .ZN(n10799) );
  MUX2_X1 U13346 ( .A(n10799), .B(n10854), .S(n10758), .Z(n10768) );
  MUX2_X1 U13347 ( .A(n10768), .B(n12846), .S(n10723), .Z(n18816) );
  INV_X1 U13348 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14982) );
  NOR2_X1 U13349 ( .A1(n18816), .A2(n14982), .ZN(n12773) );
  NAND3_X1 U13350 ( .A1(n10723), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n10553) );
  AND2_X1 U13351 ( .A1(n10556), .A2(n10553), .ZN(n13462) );
  NAND2_X1 U13352 ( .A1(n12773), .A2(n13462), .ZN(n10554) );
  NOR2_X1 U13353 ( .A1(n12773), .A2(n13462), .ZN(n12772) );
  AOI21_X1 U13354 ( .B1(n14992), .B2(n10554), .A(n12772), .ZN(n12758) );
  INV_X1 U13355 ( .A(n10555), .ZN(n10557) );
  XNOR2_X1 U13356 ( .A(n10557), .B(n10556), .ZN(n13452) );
  INV_X1 U13357 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11194) );
  XNOR2_X1 U13358 ( .A(n13452), .B(n11194), .ZN(n12757) );
  NAND2_X1 U13359 ( .A1(n12758), .A2(n12757), .ZN(n10559) );
  NAND2_X1 U13360 ( .A1(n13452), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10558) );
  NAND2_X1 U13361 ( .A1(n10559), .A2(n10558), .ZN(n15952) );
  XNOR2_X1 U13362 ( .A(n10561), .B(n10560), .ZN(n13308) );
  XNOR2_X1 U13363 ( .A(n13308), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13516) );
  AND2_X1 U13364 ( .A1(n15952), .A2(n13516), .ZN(n10562) );
  NAND2_X1 U13365 ( .A1(n15951), .A2(n10562), .ZN(n10568) );
  INV_X1 U13366 ( .A(n13308), .ZN(n10563) );
  NAND2_X1 U13367 ( .A1(n10563), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10567) );
  INV_X1 U13368 ( .A(n13516), .ZN(n10565) );
  NAND2_X1 U13369 ( .A1(n10564), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13513) );
  OR2_X1 U13370 ( .A1(n10565), .A2(n13513), .ZN(n10566) );
  NAND3_X1 U13371 ( .A1(n10568), .A2(n10567), .A3(n10566), .ZN(n15932) );
  NAND2_X1 U13372 ( .A1(n15931), .A2(n15932), .ZN(n10571) );
  NAND2_X1 U13373 ( .A1(n10569), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10570) );
  NAND2_X1 U13374 ( .A1(n10571), .A2(n10570), .ZN(n12633) );
  AOI22_X1 U13375 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10467), .B1(
        n19202), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10579) );
  AOI22_X1 U13376 ( .A1(n18993), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n19296), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10578) );
  AOI22_X1 U13377 ( .A1(n19260), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__6__SCAN_IN), .B2(n19233), .ZN(n10577) );
  AOI22_X1 U13378 ( .A1(n10468), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10469), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10576) );
  INV_X1 U13379 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10582) );
  INV_X1 U13380 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10581) );
  OAI22_X1 U13381 ( .A1(n10580), .A2(n10582), .B1(n10581), .B2(n19397), .ZN(
        n10586) );
  INV_X1 U13382 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10584) );
  INV_X1 U13383 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10583) );
  OAI22_X1 U13384 ( .A1(n10584), .A2(n19332), .B1(n19358), .B2(n10583), .ZN(
        n10585) );
  NOR2_X1 U13385 ( .A1(n10586), .A2(n10585), .ZN(n10589) );
  AOI22_X1 U13386 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10474), .B1(
        n19439), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10588) );
  AOI22_X1 U13387 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19167), .B1(
        n10461), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10587) );
  NAND4_X1 U13388 ( .A1(n10590), .A2(n10589), .A3(n10588), .A4(n10587), .ZN(
        n10603) );
  AOI22_X1 U13389 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n10794), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10594) );
  AOI22_X1 U13390 ( .A1(n10449), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U13391 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10592) );
  AOI22_X1 U13392 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11417), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10591) );
  NAND4_X1 U13393 ( .A1(n10594), .A2(n10593), .A3(n10592), .A4(n10591), .ZN(
        n10600) );
  AOI22_X1 U13394 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10417), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10598) );
  AOI22_X1 U13395 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10429), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10597) );
  AOI22_X1 U13396 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10415), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10596) );
  AOI22_X1 U13397 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10413), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10595) );
  NAND4_X1 U13398 ( .A1(n10598), .A2(n10597), .A3(n10596), .A4(n10595), .ZN(
        n10599) );
  INV_X1 U13399 ( .A(n10895), .ZN(n10601) );
  NAND2_X1 U13400 ( .A1(n10601), .A2(n12874), .ZN(n10602) );
  NAND2_X1 U13401 ( .A1(n10829), .A2(n10522), .ZN(n10607) );
  INV_X1 U13402 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n10604) );
  MUX2_X1 U13403 ( .A(n10895), .B(n10604), .S(n10723), .Z(n10611) );
  INV_X1 U13404 ( .A(n10611), .ZN(n10605) );
  XNOR2_X1 U13405 ( .A(n10612), .B(n10605), .ZN(n18781) );
  INV_X1 U13406 ( .A(n18781), .ZN(n10606) );
  NAND2_X1 U13407 ( .A1(n10607), .A2(n10606), .ZN(n10608) );
  INV_X1 U13408 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16013) );
  NAND2_X1 U13409 ( .A1(n12633), .A2(n12634), .ZN(n10610) );
  NAND2_X1 U13410 ( .A1(n10608), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10609) );
  NAND2_X1 U13411 ( .A1(n9610), .A2(n10613), .ZN(n10897) );
  INV_X1 U13412 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13043) );
  NAND2_X1 U13413 ( .A1(n10723), .A2(n13043), .ZN(n10614) );
  NAND2_X1 U13414 ( .A1(n10616), .A2(n10615), .ZN(n10617) );
  NAND2_X1 U13415 ( .A1(n10625), .A2(n10617), .ZN(n13318) );
  NOR2_X1 U13416 ( .A1(n13318), .A2(n10522), .ZN(n10629) );
  AND2_X1 U13417 ( .A1(n10629), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15921) );
  XNOR2_X1 U13418 ( .A(n10618), .B(n9698), .ZN(n18772) );
  AND2_X1 U13419 ( .A1(n18772), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15918) );
  INV_X1 U13420 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n18858) );
  INV_X1 U13421 ( .A(n10633), .ZN(n10623) );
  NOR2_X1 U13422 ( .A1(n10619), .A2(n18858), .ZN(n10620) );
  NAND2_X1 U13423 ( .A1(n10723), .A2(n10620), .ZN(n10621) );
  AND2_X1 U13424 ( .A1(n10714), .A2(n10621), .ZN(n10622) );
  NAND2_X1 U13425 ( .A1(n10623), .A2(n10622), .ZN(n18750) );
  OR2_X1 U13426 ( .A1(n18750), .A2(n10522), .ZN(n10624) );
  INV_X1 U13427 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n20808) );
  NAND2_X1 U13428 ( .A1(n10624), .A2(n20808), .ZN(n15893) );
  NAND2_X1 U13429 ( .A1(n10625), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10626) );
  MUX2_X1 U13430 ( .A(n10626), .B(n10625), .S(n9610), .Z(n10628) );
  INV_X1 U13431 ( .A(n10619), .ZN(n10627) );
  NAND2_X1 U13432 ( .A1(n10628), .A2(n10627), .ZN(n18758) );
  INV_X1 U13433 ( .A(n18758), .ZN(n10637) );
  AOI21_X1 U13434 ( .B1(n10637), .B2(n10737), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15909) );
  INV_X1 U13435 ( .A(n15909), .ZN(n10631) );
  INV_X1 U13436 ( .A(n10629), .ZN(n10630) );
  INV_X1 U13437 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16023) );
  NAND2_X1 U13438 ( .A1(n10630), .A2(n16023), .ZN(n15920) );
  OR2_X1 U13439 ( .A1(n18772), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15919) );
  AND2_X1 U13440 ( .A1(n15920), .A2(n15919), .ZN(n15908) );
  AND2_X1 U13441 ( .A1(n15893), .A2(n9700), .ZN(n10632) );
  INV_X1 U13442 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n18736) );
  AND3_X1 U13443 ( .A1(n10723), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n10623), .ZN(
        n10634) );
  OR2_X1 U13444 ( .A1(n10641), .A2(n10634), .ZN(n18735) );
  INV_X1 U13445 ( .A(n18735), .ZN(n10635) );
  AOI21_X1 U13446 ( .B1(n10635), .B2(n10737), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15881) );
  AND2_X1 U13447 ( .A1(n10737), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10636) );
  NAND2_X1 U13448 ( .A1(n10637), .A2(n10636), .ZN(n15890) );
  NAND2_X1 U13449 ( .A1(n10737), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10638) );
  OR2_X1 U13450 ( .A1(n18750), .A2(n10638), .ZN(n15892) );
  NAND2_X1 U13451 ( .A1(n15890), .A2(n15892), .ZN(n15879) );
  NAND2_X1 U13452 ( .A1(n10737), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10639) );
  NOR2_X1 U13453 ( .A1(n18735), .A2(n10639), .ZN(n15880) );
  NOR2_X1 U13454 ( .A1(n15879), .A2(n15880), .ZN(n10640) );
  NAND2_X1 U13455 ( .A1(n10723), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10642) );
  NAND2_X1 U13456 ( .A1(n10045), .A2(n10643), .ZN(n10644) );
  AND2_X1 U13457 ( .A1(n10646), .A2(n10644), .ZN(n18729) );
  NAND2_X1 U13458 ( .A1(n18729), .A2(n10737), .ZN(n15869) );
  INV_X1 U13459 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15872) );
  NAND2_X1 U13460 ( .A1(n10646), .A2(n10645), .ZN(n10647) );
  NAND2_X1 U13461 ( .A1(n10677), .A2(n10647), .ZN(n13531) );
  INV_X1 U13462 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14957) );
  OAI21_X1 U13463 ( .B1(n13531), .B2(n10522), .A(n14957), .ZN(n14744) );
  NAND2_X1 U13464 ( .A1(n15869), .A2(n15872), .ZN(n14742) );
  NAND2_X1 U13465 ( .A1(n10723), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10673) );
  NAND2_X1 U13466 ( .A1(n10723), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10663) );
  OR2_X1 U13467 ( .A1(n10666), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10653) );
  NAND3_X1 U13468 ( .A1(n10653), .A2(P2_EBX_REG_19__SCAN_IN), .A3(n10723), 
        .ZN(n10651) );
  INV_X1 U13469 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n13635) );
  INV_X1 U13470 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n10648) );
  NAND2_X1 U13471 ( .A1(n13635), .A2(n10648), .ZN(n10649) );
  AND2_X1 U13472 ( .A1(n10723), .A2(n10649), .ZN(n10650) );
  NAND2_X1 U13473 ( .A1(n10651), .A2(n10657), .ZN(n14510) );
  NOR2_X1 U13474 ( .A1(n14510), .A2(n10522), .ZN(n10682) );
  NOR2_X1 U13475 ( .A1(n10682), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14707) );
  NAND2_X1 U13476 ( .A1(n10666), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10652) );
  MUX2_X1 U13477 ( .A(n10652), .B(n10666), .S(n9610), .Z(n10654) );
  NAND2_X1 U13478 ( .A1(n10654), .A2(n10653), .ZN(n18667) );
  INV_X1 U13479 ( .A(n18667), .ZN(n10655) );
  AOI21_X1 U13480 ( .B1(n10655), .B2(n10737), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14890) );
  NOR2_X1 U13481 ( .A1(n14707), .A2(n14890), .ZN(n14689) );
  NAND2_X1 U13482 ( .A1(n10657), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10656) );
  MUX2_X1 U13483 ( .A(n10657), .B(n10656), .S(n10723), .Z(n10658) );
  INV_X1 U13484 ( .A(n10659), .ZN(n10660) );
  NAND2_X1 U13485 ( .A1(n10658), .A2(n10660), .ZN(n14494) );
  INV_X1 U13486 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14697) );
  OAI21_X1 U13487 ( .B1(n14494), .B2(n10522), .A(n14697), .ZN(n14690) );
  NAND2_X1 U13488 ( .A1(n14689), .A2(n14690), .ZN(n14677) );
  INV_X1 U13489 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14555) );
  INV_X1 U13490 ( .A(n10697), .ZN(n10662) );
  NAND3_X1 U13491 ( .A1(n10660), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n10723), 
        .ZN(n10661) );
  NAND2_X1 U13492 ( .A1(n10662), .A2(n10661), .ZN(n12654) );
  INV_X1 U13493 ( .A(n12654), .ZN(n10681) );
  AOI21_X1 U13494 ( .B1(n10681), .B2(n10737), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14679) );
  OR2_X1 U13495 ( .A1(n10664), .A2(n10663), .ZN(n10665) );
  NAND2_X1 U13496 ( .A1(n10666), .A2(n10665), .ZN(n18679) );
  INV_X1 U13497 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14920) );
  OAI21_X1 U13498 ( .B1(n18679), .B2(n10522), .A(n14920), .ZN(n14673) );
  AND2_X1 U13499 ( .A1(n10723), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10668) );
  INV_X1 U13500 ( .A(n10714), .ZN(n10667) );
  AOI21_X1 U13501 ( .B1(n10669), .B2(n10668), .A(n10667), .ZN(n10671) );
  NAND2_X1 U13502 ( .A1(n10671), .A2(n10670), .ZN(n18693) );
  OR2_X1 U13503 ( .A1(n18693), .A2(n10522), .ZN(n10672) );
  XNOR2_X1 U13504 ( .A(n10672), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14669) );
  INV_X1 U13505 ( .A(n10673), .ZN(n10674) );
  XNOR2_X1 U13506 ( .A(n10675), .B(n10674), .ZN(n18706) );
  NAND2_X1 U13507 ( .A1(n18706), .A2(n10737), .ZN(n10676) );
  INV_X1 U13508 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15962) );
  NAND2_X1 U13509 ( .A1(n10676), .A2(n15962), .ZN(n14734) );
  XNOR2_X1 U13510 ( .A(n10677), .B(n9732), .ZN(n18718) );
  NAND2_X1 U13511 ( .A1(n18718), .A2(n10737), .ZN(n10678) );
  INV_X1 U13512 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14943) );
  NAND2_X1 U13513 ( .A1(n10678), .A2(n14943), .ZN(n14933) );
  NAND4_X1 U13514 ( .A1(n14673), .A2(n14669), .A3(n14734), .A4(n14933), .ZN(
        n10679) );
  NAND3_X1 U13515 ( .A1(n10681), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n10737), .ZN(n14678) );
  NAND2_X1 U13516 ( .A1(n10737), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10683) );
  NOR2_X1 U13517 ( .A1(n18693), .A2(n10683), .ZN(n14670) );
  AND2_X1 U13518 ( .A1(n10737), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10684) );
  AND2_X1 U13519 ( .A1(n18706), .A2(n10684), .ZN(n14667) );
  NAND2_X1 U13520 ( .A1(n10737), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10685) );
  NOR2_X1 U13521 ( .A1(n13531), .A2(n10685), .ZN(n14666) );
  AND2_X1 U13522 ( .A1(n10737), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10686) );
  NOR4_X1 U13523 ( .A1(n14670), .A2(n14667), .A3(n14666), .A4(n14932), .ZN(
        n10689) );
  INV_X1 U13524 ( .A(n18679), .ZN(n10688) );
  AND2_X1 U13525 ( .A1(n10737), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10687) );
  NAND2_X1 U13526 ( .A1(n10688), .A2(n10687), .ZN(n14672) );
  NAND2_X1 U13527 ( .A1(n10689), .A2(n14672), .ZN(n10690) );
  NAND2_X1 U13528 ( .A1(n10737), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10692) );
  NOR2_X1 U13529 ( .A1(n14494), .A2(n10692), .ZN(n14676) );
  NAND2_X1 U13530 ( .A1(n10737), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10693) );
  NOR2_X1 U13531 ( .A1(n18667), .A2(n10693), .ZN(n14887) );
  INV_X1 U13532 ( .A(n10696), .ZN(n10699) );
  NAND2_X1 U13533 ( .A1(n10723), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10698) );
  OAI21_X1 U13534 ( .B1(n10699), .B2(n10698), .A(n10702), .ZN(n15383) );
  INV_X1 U13535 ( .A(n15383), .ZN(n10700) );
  AOI21_X1 U13536 ( .B1(n10700), .B2(n10737), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12606) );
  AND2_X1 U13537 ( .A1(n10723), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10701) );
  NAND2_X1 U13538 ( .A1(n10702), .A2(n10701), .ZN(n10703) );
  NAND2_X1 U13539 ( .A1(n10709), .A2(n10703), .ZN(n12668) );
  XNOR2_X1 U13540 ( .A(n10704), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14657) );
  INV_X1 U13541 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14839) );
  NOR3_X1 U13542 ( .A1(n12668), .A2(n10522), .A3(n14839), .ZN(n10705) );
  AOI21_X2 U13543 ( .B1(n14658), .B2(n14657), .A(n10705), .ZN(n14825) );
  INV_X1 U13544 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14830) );
  NAND2_X1 U13545 ( .A1(n10723), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10706) );
  MUX2_X1 U13546 ( .A(P2_EBX_REG_24__SCAN_IN), .B(n10706), .S(n10709), .Z(
        n10707) );
  NAND2_X1 U13547 ( .A1(n10707), .A2(n10714), .ZN(n15799) );
  NOR2_X1 U13548 ( .A1(n15799), .A2(n10522), .ZN(n14823) );
  INV_X1 U13549 ( .A(n14823), .ZN(n10708) );
  INV_X1 U13550 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n20797) );
  AND3_X1 U13551 ( .A1(n10723), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n10716), .ZN(
        n10710) );
  NOR2_X1 U13552 ( .A1(n10740), .A2(n10710), .ZN(n10711) );
  NAND3_X1 U13553 ( .A1(n10711), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n10737), .ZN(n10732) );
  NOR2_X1 U13554 ( .A1(n9677), .A2(n20797), .ZN(n10712) );
  NAND2_X1 U13555 ( .A1(n10723), .A2(n10712), .ZN(n10713) );
  AND2_X1 U13556 ( .A1(n10714), .A2(n10713), .ZN(n10715) );
  NAND2_X1 U13557 ( .A1(n10716), .A2(n10715), .ZN(n14488) );
  INV_X1 U13558 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14817) );
  NAND2_X1 U13559 ( .A1(n10723), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10720) );
  INV_X1 U13560 ( .A(n10720), .ZN(n10721) );
  NAND2_X1 U13561 ( .A1(n10721), .A2(n10124), .ZN(n10722) );
  NAND2_X1 U13562 ( .A1(n10725), .A2(n10722), .ZN(n12641) );
  AND2_X1 U13563 ( .A1(n10723), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10724) );
  NAND2_X1 U13564 ( .A1(n10725), .A2(n10724), .ZN(n10726) );
  NAND2_X1 U13565 ( .A1(n10735), .A2(n10726), .ZN(n14463) );
  OAI21_X1 U13566 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n14618), .ZN(n10727) );
  INV_X1 U13567 ( .A(n14618), .ZN(n10729) );
  INV_X1 U13568 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n20809) );
  INV_X1 U13569 ( .A(n10730), .ZN(n10731) );
  NAND2_X1 U13570 ( .A1(n10731), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14645) );
  NAND2_X1 U13571 ( .A1(n14645), .A2(n10732), .ZN(n14613) );
  AND2_X1 U13572 ( .A1(n10723), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10734) );
  INV_X1 U13573 ( .A(n10734), .ZN(n10733) );
  XNOR2_X1 U13574 ( .A(n10735), .B(n10733), .ZN(n10739) );
  AOI21_X1 U13575 ( .B1(n10739), .B2(n10737), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14604) );
  NAND2_X1 U13576 ( .A1(n10723), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10736) );
  XNOR2_X1 U13577 ( .A(n13893), .B(n10736), .ZN(n11284) );
  INV_X1 U13578 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14761) );
  OAI21_X1 U13579 ( .B1(n11284), .B2(n10522), .A(n14761), .ZN(n13876) );
  NAND2_X1 U13580 ( .A1(n10737), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10738) );
  NOR2_X1 U13581 ( .A1(n11284), .A2(n10738), .ZN(n13877) );
  INV_X1 U13582 ( .A(n10739), .ZN(n15776) );
  INV_X1 U13583 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14772) );
  NOR2_X1 U13584 ( .A1(n10740), .A2(n10897), .ZN(n10741) );
  XOR2_X1 U13585 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n10741), .Z(
        n10742) );
  XNOR2_X1 U13586 ( .A(n10743), .B(n10742), .ZN(n11208) );
  AND2_X1 U13587 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12878), .ZN(
        n10744) );
  NAND2_X1 U13588 ( .A1(n12874), .A2(n10799), .ZN(n10748) );
  XNOR2_X1 U13589 ( .A(n10766), .B(n10746), .ZN(n10777) );
  INV_X1 U13590 ( .A(n10776), .ZN(n10747) );
  AOI22_X1 U13591 ( .A1(n10748), .A2(n10777), .B1(n12874), .B2(n10747), .ZN(
        n10751) );
  INV_X1 U13592 ( .A(n10766), .ZN(n10749) );
  OAI21_X1 U13593 ( .B1(n10799), .B2(n10749), .A(n10758), .ZN(n10750) );
  OAI21_X1 U13594 ( .B1(n10751), .B2(n11272), .A(n10750), .ZN(n10756) );
  INV_X1 U13595 ( .A(n12814), .ZN(n10752) );
  NAND2_X1 U13596 ( .A1(n10752), .A2(n12686), .ZN(n10753) );
  MUX2_X1 U13597 ( .A(n11267), .B(n10753), .S(n10776), .Z(n10755) );
  NAND2_X1 U13598 ( .A1(n10754), .A2(n10757), .ZN(n10775) );
  AOI21_X1 U13599 ( .B1(n10756), .B2(n10755), .A(n10775), .ZN(n10760) );
  OAI21_X1 U13600 ( .B1(n10758), .B2(n10757), .A(n10770), .ZN(n10759) );
  NOR2_X1 U13601 ( .A1(n10760), .A2(n10759), .ZN(n10761) );
  OR2_X1 U13602 ( .A1(n10779), .A2(n10761), .ZN(n10762) );
  MUX2_X1 U13603 ( .A(n10762), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18640), .Z(n10764) );
  NAND2_X1 U13604 ( .A1(n10779), .A2(n12814), .ZN(n10763) );
  NAND2_X1 U13605 ( .A1(n16090), .A2(n12686), .ZN(n12865) );
  NOR2_X1 U13606 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19516) );
  AOI211_X1 U13607 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n19516), .ZN(n19510) );
  NAND2_X1 U13608 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19504) );
  AND2_X1 U13609 ( .A1(n19510), .A2(n19504), .ZN(n12866) );
  NAND2_X1 U13610 ( .A1(n11163), .A2(n12866), .ZN(n10810) );
  AOI21_X1 U13611 ( .B1(n10764), .B2(n10253), .A(n9782), .ZN(n10765) );
  NAND2_X1 U13612 ( .A1(n12865), .A2(n10765), .ZN(n10809) );
  OAI21_X1 U13613 ( .B1(n10768), .B2(n10749), .A(n10767), .ZN(n10772) );
  AND2_X1 U13614 ( .A1(n10770), .A2(n10769), .ZN(n10771) );
  AND2_X1 U13615 ( .A1(n10772), .A2(n10771), .ZN(n10773) );
  NOR2_X1 U13616 ( .A1(n10779), .A2(n10773), .ZN(n19615) );
  INV_X1 U13617 ( .A(n14454), .ZN(n10774) );
  NOR2_X1 U13618 ( .A1(n16096), .A2(n10774), .ZN(n19618) );
  NAND2_X1 U13619 ( .A1(n19615), .A2(n19618), .ZN(n11206) );
  NOR2_X1 U13620 ( .A1(n10776), .A2(n10775), .ZN(n10800) );
  AND2_X1 U13621 ( .A1(n10777), .A2(n10800), .ZN(n10778) );
  OR2_X1 U13622 ( .A1(n10779), .A2(n10778), .ZN(n16087) );
  NAND2_X1 U13623 ( .A1(n10792), .A2(n12866), .ZN(n10780) );
  OR2_X1 U13624 ( .A1(n16087), .A2(n10780), .ZN(n10791) );
  NAND2_X1 U13625 ( .A1(n10781), .A2(n18958), .ZN(n10782) );
  NAND2_X1 U13626 ( .A1(n10782), .A2(n12876), .ZN(n10789) );
  NAND2_X1 U13627 ( .A1(n10783), .A2(n12874), .ZN(n11161) );
  AOI21_X1 U13628 ( .B1(n11161), .B2(n10253), .A(n18981), .ZN(n10786) );
  NAND2_X1 U13629 ( .A1(n10784), .A2(n12844), .ZN(n10785) );
  NAND2_X1 U13630 ( .A1(n10785), .A2(n14454), .ZN(n11176) );
  OAI211_X1 U13631 ( .C1(n10786), .C2(n11163), .A(n11176), .B(n11166), .ZN(
        n10787) );
  INV_X1 U13632 ( .A(n10787), .ZN(n10788) );
  NAND2_X1 U13633 ( .A1(n10789), .A2(n10788), .ZN(n11162) );
  INV_X1 U13634 ( .A(n11162), .ZN(n10790) );
  AND2_X1 U13635 ( .A1(n10791), .A2(n10790), .ZN(n12863) );
  MUX2_X1 U13636 ( .A(n10792), .B(n11163), .S(n12874), .Z(n10793) );
  NAND2_X1 U13637 ( .A1(n10793), .A2(n19504), .ZN(n10805) );
  NAND2_X1 U13638 ( .A1(n15005), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10796) );
  NAND2_X1 U13639 ( .A1(n10796), .A2(n12878), .ZN(n12873) );
  INV_X1 U13640 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n10797) );
  OAI21_X1 U13641 ( .B1(n10794), .B2(n12873), .A(n10797), .ZN(n10798) );
  NAND2_X1 U13642 ( .A1(n10798), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19605) );
  INV_X1 U13643 ( .A(n10799), .ZN(n10801) );
  AOI21_X1 U13644 ( .B1(n10801), .B2(n10800), .A(n16087), .ZN(n10802) );
  NAND2_X1 U13645 ( .A1(n11065), .A2(n10802), .ZN(n10803) );
  NAND2_X1 U13646 ( .A1(n19605), .A2(n10803), .ZN(n16111) );
  NAND2_X1 U13647 ( .A1(n12686), .A2(n16111), .ZN(n10804) );
  OAI22_X1 U13648 ( .A1(n16087), .A2(n10805), .B1(n16096), .B2(n10804), .ZN(
        n10806) );
  INV_X1 U13649 ( .A(n10806), .ZN(n10807) );
  OAI211_X1 U13650 ( .C1(n12865), .C2(n10810), .A(n10809), .B(n10808), .ZN(
        n10811) );
  NAND2_X1 U13651 ( .A1(n11065), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11280) );
  NOR2_X1 U13652 ( .A1(n16096), .A2(n11267), .ZN(n19617) );
  NAND2_X1 U13653 ( .A1(n11208), .A2(n16063), .ZN(n11204) );
  INV_X1 U13654 ( .A(n10854), .ZN(n12779) );
  NOR2_X1 U13655 ( .A1(n12779), .A2(n14982), .ZN(n12778) );
  INV_X1 U13656 ( .A(n12778), .ZN(n10813) );
  NOR2_X1 U13657 ( .A1(n10863), .A2(n10813), .ZN(n10815) );
  NOR2_X1 U13658 ( .A1(n12779), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10814) );
  XNOR2_X1 U13659 ( .A(n10814), .B(n10863), .ZN(n12770) );
  NOR2_X1 U13660 ( .A1(n14992), .A2(n12770), .ZN(n12769) );
  NOR2_X1 U13661 ( .A1(n10815), .A2(n12769), .ZN(n10817) );
  XNOR2_X1 U13662 ( .A(n11194), .B(n10817), .ZN(n12760) );
  XNOR2_X1 U13663 ( .A(n10816), .B(n10870), .ZN(n12759) );
  OR2_X1 U13664 ( .A1(n10817), .A2(n11194), .ZN(n10818) );
  OAI21_X1 U13665 ( .B1(n12760), .B2(n12759), .A(n10818), .ZN(n10819) );
  NAND2_X1 U13666 ( .A1(n10819), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10820) );
  NAND2_X2 U13667 ( .A1(n15950), .A2(n10820), .ZN(n10825) );
  XNOR2_X2 U13668 ( .A(n10825), .B(n10823), .ZN(n13512) );
  INV_X1 U13669 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16042) );
  NOR2_X1 U13670 ( .A1(n10825), .A2(n10824), .ZN(n10826) );
  AOI21_X2 U13671 ( .B1(n13512), .B2(n16042), .A(n10826), .ZN(n15937) );
  INV_X1 U13672 ( .A(n10827), .ZN(n10828) );
  NAND2_X1 U13673 ( .A1(n10828), .A2(n16043), .ZN(n15936) );
  NAND2_X1 U13674 ( .A1(n10827), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15935) );
  INV_X1 U13675 ( .A(n15935), .ZN(n15933) );
  NAND2_X1 U13676 ( .A1(n15933), .A2(n10835), .ZN(n10833) );
  AND2_X1 U13677 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n10843), .ZN(
        n10837) );
  NAND2_X1 U13678 ( .A1(n12632), .A2(n10837), .ZN(n10841) );
  INV_X1 U13679 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16012) );
  NAND2_X1 U13680 ( .A1(n12632), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10842) );
  INV_X1 U13681 ( .A(n10845), .ZN(n10846) );
  NAND3_X1 U13682 ( .A1(n10846), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n10737), .ZN(n10847) );
  AND2_X1 U13683 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15979) );
  AND3_X1 U13684 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14914) );
  NAND3_X1 U13685 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15979), .A3(
        n14914), .ZN(n14908) );
  INV_X1 U13686 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14915) );
  NOR4_X1 U13687 ( .A1(n14920), .A2(n14908), .A3(n15962), .A4(n14915), .ZN(
        n14892) );
  NAND2_X1 U13688 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n14892), .ZN(
        n14863) );
  NAND2_X1 U13689 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12617) );
  NOR2_X1 U13690 ( .A1(n14863), .A2(n12617), .ZN(n14850) );
  NAND2_X1 U13691 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n14850), .ZN(
        n12609) );
  INV_X1 U13692 ( .A(n12609), .ZN(n10848) );
  NAND3_X1 U13693 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n10848), .ZN(n11186) );
  INV_X1 U13694 ( .A(n11186), .ZN(n11197) );
  AND2_X4 U13695 ( .A1(n14826), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15846) );
  INV_X1 U13696 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14804) );
  INV_X1 U13697 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14779) );
  NAND2_X1 U13698 ( .A1(n14608), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10850) );
  NOR2_X2 U13699 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19390) );
  NAND2_X1 U13700 ( .A1(n19390), .A2(n11065), .ZN(n18639) );
  OR2_X1 U13701 ( .A1(n18639), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11181) );
  NAND2_X1 U13702 ( .A1(n18933), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n11210) );
  MUX2_X1 U13703 ( .A(n12844), .B(n19613), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10853) );
  INV_X1 U13704 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19582) );
  NAND2_X1 U13705 ( .A1(n18981), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n10858) );
  OAI211_X1 U13706 ( .C1(n12874), .C2(n14982), .A(n10858), .B(n19582), .ZN(
        n10859) );
  INV_X1 U13707 ( .A(n10859), .ZN(n10860) );
  OAI21_X1 U13708 ( .B1(n11047), .B2(n10280), .A(n10860), .ZN(n12856) );
  NOR2_X1 U13709 ( .A1(n11047), .A2(n12768), .ZN(n10862) );
  INV_X1 U13710 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n18929) );
  OAI22_X1 U13711 ( .A1(n11043), .A2(n14992), .B1(n11017), .B2(n18929), .ZN(
        n10861) );
  OR2_X1 U13712 ( .A1(n10863), .A2(n9986), .ZN(n10866) );
  NAND2_X1 U13713 ( .A1(n10864), .A2(n12844), .ZN(n12854) );
  MUX2_X1 U13714 ( .A(n12854), .B(n19603), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10865) );
  NAND2_X1 U13715 ( .A1(n10866), .A2(n10865), .ZN(n12926) );
  NOR2_X1 U13716 ( .A1(n12925), .A2(n12926), .ZN(n10869) );
  NAND2_X1 U13717 ( .A1(n10991), .A2(n10870), .ZN(n10871) );
  OAI211_X1 U13718 ( .C1(n19582), .C2(n19596), .A(n10872), .B(n10871), .ZN(
        n10875) );
  XNOR2_X1 U13719 ( .A(n10876), .B(n10875), .ZN(n12934) );
  NOR2_X1 U13720 ( .A1(n11047), .A2(n12761), .ZN(n10874) );
  INV_X1 U13721 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n18926) );
  OAI22_X1 U13722 ( .A1(n11043), .A2(n11194), .B1(n11017), .B2(n18926), .ZN(
        n10873) );
  NOR2_X1 U13723 ( .A1(n12934), .A2(n12933), .ZN(n12935) );
  NOR2_X1 U13724 ( .A1(n10876), .A2(n10875), .ZN(n10877) );
  INV_X1 U13725 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n10878) );
  OR2_X1 U13726 ( .A1(n11017), .A2(n10878), .ZN(n10880) );
  NAND2_X1 U13727 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10879) );
  OAI211_X1 U13728 ( .C1(n11043), .C2(n16067), .A(n10880), .B(n10879), .ZN(
        n10881) );
  INV_X1 U13729 ( .A(n10881), .ZN(n10884) );
  NAND2_X1 U13730 ( .A1(n10991), .A2(n10882), .ZN(n10883) );
  OAI211_X1 U13731 ( .C1(n11047), .C2(n16054), .A(n10884), .B(n10883), .ZN(
        n13139) );
  INV_X1 U13732 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n10885) );
  OAI22_X1 U13733 ( .A1(n11043), .A2(n16042), .B1(n11017), .B2(n10885), .ZN(
        n10886) );
  INV_X1 U13734 ( .A(n10886), .ZN(n10890) );
  NAND2_X1 U13735 ( .A1(n11040), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10889) );
  NAND2_X1 U13736 ( .A1(n10991), .A2(n10887), .ZN(n10888) );
  AOI22_X1 U13737 ( .A1(n11039), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n11044), .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n10894) );
  INV_X1 U13738 ( .A(n10891), .ZN(n10892) );
  AOI22_X1 U13739 ( .A1(n11040), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n10892), 
        .B2(n12839), .ZN(n10893) );
  NAND2_X1 U13740 ( .A1(n10894), .A2(n10893), .ZN(n13159) );
  AOI222_X1 U13741 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n11040), .B1(n11039), 
        .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(P2_EAX_REG_6__SCAN_IN), 
        .C2(n11044), .ZN(n12630) );
  INV_X1 U13742 ( .A(n12839), .ZN(n10898) );
  INV_X1 U13743 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n18915) );
  INV_X1 U13744 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19532) );
  OAI222_X1 U13745 ( .A1(n16012), .A2(n11043), .B1(n11017), .B2(n18915), .C1(
        n11047), .C2(n19532), .ZN(n12950) );
  INV_X1 U13746 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n10899) );
  OAI22_X1 U13747 ( .A1(n11043), .A2(n16023), .B1(n11017), .B2(n10899), .ZN(
        n10900) );
  INV_X1 U13748 ( .A(n10900), .ZN(n10914) );
  NAND2_X1 U13749 ( .A1(n11040), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10913) );
  AOI22_X1 U13750 ( .A1(n10449), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10905) );
  AOI22_X1 U13751 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10904) );
  AOI22_X1 U13752 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10903) );
  AOI22_X1 U13753 ( .A1(n10454), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10902) );
  NAND4_X1 U13754 ( .A1(n10905), .A2(n10904), .A3(n10903), .A4(n10902), .ZN(
        n10911) );
  AOI22_X1 U13755 ( .A1(n10504), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9616), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U13756 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11417), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10908) );
  AOI22_X1 U13757 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10907) );
  AOI22_X1 U13758 ( .A1(n10415), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10906) );
  NAND4_X1 U13759 ( .A1(n10909), .A2(n10908), .A3(n10907), .A4(n10906), .ZN(
        n10910) );
  NAND2_X1 U13760 ( .A1(n10991), .A2(n18860), .ZN(n10912) );
  AOI22_X1 U13761 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10794), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10918) );
  AOI22_X1 U13762 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10449), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U13763 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U13764 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11416), .B1(
        n11417), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10915) );
  NAND4_X1 U13765 ( .A1(n10918), .A2(n10917), .A3(n10916), .A4(n10915), .ZN(
        n10924) );
  AOI22_X1 U13766 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9616), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U13767 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10429), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10921) );
  AOI22_X1 U13768 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10415), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10920) );
  AOI22_X1 U13769 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10413), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10919) );
  NAND4_X1 U13770 ( .A1(n10922), .A2(n10921), .A3(n10920), .A4(n10919), .ZN(
        n10923) );
  INV_X1 U13771 ( .A(n13107), .ZN(n10927) );
  AOI22_X1 U13772 ( .A1(n11039), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n11044), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n10926) );
  NAND2_X1 U13773 ( .A1(n11040), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10925) );
  OAI211_X1 U13774 ( .C1(n9986), .C2(n10927), .A(n10926), .B(n10925), .ZN(
        n13127) );
  AOI22_X1 U13775 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n10794), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10931) );
  AOI22_X1 U13776 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10449), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10930) );
  AOI22_X1 U13777 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U13778 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n11416), .B1(
        n11417), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10928) );
  NAND4_X1 U13779 ( .A1(n10931), .A2(n10930), .A3(n10929), .A4(n10928), .ZN(
        n10937) );
  AOI22_X1 U13780 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n9616), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10935) );
  AOI22_X1 U13781 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10429), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U13782 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10415), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U13783 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10413), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10932) );
  NAND4_X1 U13784 ( .A1(n10935), .A2(n10934), .A3(n10933), .A4(n10932), .ZN(
        n10936) );
  INV_X1 U13785 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U13786 ( .A1(n11039), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n11044), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n10938) );
  OAI21_X1 U13787 ( .B1(n11047), .B2(n10939), .A(n10938), .ZN(n10940) );
  AOI21_X1 U13788 ( .B1(n10991), .B2(n18852), .A(n10940), .ZN(n15987) );
  INV_X1 U13789 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n11088) );
  INV_X1 U13790 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15980) );
  OAI22_X1 U13791 ( .A1(n11047), .A2(n11088), .B1(n11043), .B2(n15980), .ZN(
        n10941) );
  INV_X1 U13792 ( .A(n10941), .ZN(n10953) );
  AOI22_X1 U13793 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n10794), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10945) );
  AOI22_X1 U13794 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10449), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U13795 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U13796 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n11416), .B1(
        n11417), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10942) );
  NAND4_X1 U13797 ( .A1(n10945), .A2(n10944), .A3(n10943), .A4(n10942), .ZN(
        n10951) );
  AOI22_X1 U13798 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n9616), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10949) );
  AOI22_X1 U13799 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10454), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U13800 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10415), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10947) );
  AOI22_X1 U13801 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10413), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10946) );
  NAND4_X1 U13802 ( .A1(n10949), .A2(n10948), .A3(n10947), .A4(n10946), .ZN(
        n10950) );
  OR2_X1 U13803 ( .A1(n10951), .A2(n10950), .ZN(n18845) );
  AOI22_X1 U13804 ( .A1(n10991), .A2(n18845), .B1(n11044), .B2(
        P2_EAX_REG_11__SCAN_IN), .ZN(n10952) );
  NAND2_X1 U13805 ( .A1(n10953), .A2(n10952), .ZN(n13184) );
  NAND2_X1 U13806 ( .A1(n13185), .A2(n13184), .ZN(n13183) );
  AOI22_X1 U13807 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U13808 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10449), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10956) );
  AOI22_X1 U13809 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10955) );
  AOI22_X1 U13810 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10454), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10954) );
  NAND4_X1 U13811 ( .A1(n10957), .A2(n10956), .A3(n10955), .A4(n10954), .ZN(
        n10963) );
  AOI22_X1 U13812 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n9616), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U13813 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10429), .B1(
        n11417), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U13814 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10413), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U13815 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10415), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10958) );
  NAND4_X1 U13816 ( .A1(n10961), .A2(n10960), .A3(n10959), .A4(n10958), .ZN(
        n10962) );
  OR2_X1 U13817 ( .A1(n10963), .A2(n10962), .ZN(n18844) );
  INV_X1 U13818 ( .A(n18844), .ZN(n10965) );
  AOI22_X1 U13819 ( .A1(n11039), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n11044), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n10964) );
  OAI21_X1 U13820 ( .B1(n9986), .B2(n10965), .A(n10964), .ZN(n10966) );
  AOI21_X1 U13821 ( .B1(P2_REIP_REG_12__SCAN_IN), .B2(n11040), .A(n10966), 
        .ZN(n15968) );
  AOI22_X1 U13822 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U13823 ( .A1(n10449), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10969) );
  AOI22_X1 U13824 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10968) );
  AOI22_X1 U13825 ( .A1(n11417), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10967) );
  NAND4_X1 U13826 ( .A1(n10970), .A2(n10969), .A3(n10968), .A4(n10967), .ZN(
        n10976) );
  AOI22_X1 U13827 ( .A1(n10504), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9616), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U13828 ( .A1(n10454), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10973) );
  AOI22_X1 U13829 ( .A1(n10415), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10972) );
  AOI22_X1 U13830 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10971) );
  NAND4_X1 U13831 ( .A1(n10974), .A2(n10973), .A3(n10972), .A4(n10971), .ZN(
        n10975) );
  OR2_X1 U13832 ( .A1(n10976), .A2(n10975), .ZN(n18838) );
  AOI22_X1 U13833 ( .A1(n11040), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n10991), 
        .B2(n18838), .ZN(n10978) );
  AOI22_X1 U13834 ( .A1(n11039), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n11044), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n10977) );
  NAND2_X1 U13835 ( .A1(n10978), .A2(n10977), .ZN(n13289) );
  NAND2_X1 U13836 ( .A1(n13288), .A2(n13289), .ZN(n13442) );
  INV_X1 U13837 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n10979) );
  OAI22_X1 U13838 ( .A1(n11043), .A2(n14943), .B1(n11017), .B2(n10979), .ZN(
        n10980) );
  INV_X1 U13839 ( .A(n10980), .ZN(n10994) );
  NAND2_X1 U13840 ( .A1(n11040), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n10993) );
  AOI22_X1 U13841 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10449), .B1(
        n10794), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10984) );
  AOI22_X1 U13842 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10983) );
  AOI22_X1 U13843 ( .A1(n10901), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10982) );
  AOI22_X1 U13844 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n11416), .B1(
        n11417), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10981) );
  NAND4_X1 U13845 ( .A1(n10984), .A2(n10983), .A3(n10982), .A4(n10981), .ZN(
        n10990) );
  AOI22_X1 U13846 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n10504), .B1(
        n9616), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10988) );
  AOI22_X1 U13847 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10429), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10987) );
  AOI22_X1 U13848 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10413), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U13849 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10415), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10985) );
  NAND4_X1 U13850 ( .A1(n10988), .A2(n10987), .A3(n10986), .A4(n10985), .ZN(
        n10989) );
  OR2_X1 U13851 ( .A1(n10990), .A2(n10989), .ZN(n18837) );
  NAND2_X1 U13852 ( .A1(n10991), .A2(n18837), .ZN(n10992) );
  AOI22_X1 U13853 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n10794), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U13854 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10449), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10997) );
  AOI22_X1 U13855 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10996) );
  AOI22_X1 U13856 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11416), .B1(
        n11417), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10995) );
  NAND4_X1 U13857 ( .A1(n10998), .A2(n10997), .A3(n10996), .A4(n10995), .ZN(
        n11004) );
  AOI22_X1 U13858 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n9616), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U13859 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10429), .B1(
        n10454), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11001) );
  AOI22_X1 U13860 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10415), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U13861 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10413), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10999) );
  NAND4_X1 U13862 ( .A1(n11002), .A2(n11001), .A3(n11000), .A4(n10999), .ZN(
        n11003) );
  OR2_X1 U13863 ( .A1(n11004), .A2(n11003), .ZN(n13475) );
  INV_X1 U13864 ( .A(n13475), .ZN(n11324) );
  AOI22_X1 U13865 ( .A1(n11039), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n11044), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n11006) );
  NAND2_X1 U13866 ( .A1(n11040), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11005) );
  OAI211_X1 U13867 ( .C1(n9986), .C2(n11324), .A(n11006), .B(n11005), .ZN(
        n13481) );
  INV_X1 U13868 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n11007) );
  OAI22_X1 U13869 ( .A1(n11043), .A2(n14915), .B1(n11017), .B2(n11007), .ZN(
        n11008) );
  INV_X1 U13870 ( .A(n11008), .ZN(n11010) );
  NAND2_X1 U13871 ( .A1(n11040), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11009) );
  INV_X1 U13872 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19545) );
  NOR2_X1 U13873 ( .A1(n11047), .A2(n19545), .ZN(n11012) );
  INV_X1 U13874 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n12832) );
  OAI22_X1 U13875 ( .A1(n11043), .A2(n14920), .B1(n11017), .B2(n12832), .ZN(
        n11011) );
  OR2_X1 U13876 ( .A1(n11012), .A2(n11011), .ZN(n13593) );
  NAND2_X1 U13877 ( .A1(n13592), .A2(n13593), .ZN(n14899) );
  INV_X1 U13878 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14703) );
  INV_X1 U13879 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n11013) );
  OAI22_X1 U13880 ( .A1(n11043), .A2(n14703), .B1(n11017), .B2(n11013), .ZN(
        n11014) );
  INV_X1 U13881 ( .A(n11014), .ZN(n11016) );
  NAND2_X1 U13882 ( .A1(n11040), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11015) );
  INV_X1 U13883 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19549) );
  INV_X1 U13884 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14877) );
  INV_X1 U13885 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13615) );
  OAI222_X1 U13886 ( .A1(n11047), .A2(n19549), .B1(n11043), .B2(n14877), .C1(
        n11017), .C2(n13615), .ZN(n13614) );
  AOI22_X1 U13887 ( .A1(n11039), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n11044), .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n11019) );
  NAND2_X1 U13888 ( .A1(n11040), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11018) );
  NAND2_X1 U13889 ( .A1(n11019), .A2(n11018), .ZN(n14499) );
  AOI22_X1 U13890 ( .A1(n11039), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n11044), .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n11021) );
  NAND2_X1 U13891 ( .A1(n11040), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11020) );
  AND2_X1 U13892 ( .A1(n11021), .A2(n11020), .ZN(n12658) );
  AOI22_X1 U13893 ( .A1(n11039), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n11044), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n11023) );
  NAND2_X1 U13894 ( .A1(n11040), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11022) );
  AND2_X1 U13895 ( .A1(n11023), .A2(n11022), .ZN(n12611) );
  AOI22_X1 U13896 ( .A1(n11039), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n11044), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n11026) );
  NAND2_X1 U13897 ( .A1(n11040), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11025) );
  NAND2_X1 U13898 ( .A1(n11026), .A2(n11025), .ZN(n12675) );
  AND2_X2 U13899 ( .A1(n10127), .A2(n12675), .ZN(n12674) );
  AOI22_X1 U13900 ( .A1(n11039), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n11044), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U13901 ( .A1(n11040), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11027) );
  NAND2_X1 U13902 ( .A1(n11028), .A2(n11027), .ZN(n14584) );
  AOI22_X1 U13903 ( .A1(n11039), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n11044), .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n11030) );
  NAND2_X1 U13904 ( .A1(n11040), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11029) );
  AND2_X1 U13905 ( .A1(n11030), .A2(n11029), .ZN(n14481) );
  AOI22_X1 U13906 ( .A1(n11039), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n11044), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n11032) );
  NAND2_X1 U13907 ( .A1(n11040), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11031) );
  AND2_X1 U13908 ( .A1(n11032), .A2(n11031), .ZN(n14572) );
  AOI22_X1 U13909 ( .A1(n11039), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n11044), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n11034) );
  NAND2_X1 U13910 ( .A1(n11040), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11033) );
  AND2_X1 U13911 ( .A1(n11034), .A2(n11033), .ZN(n12645) );
  AOI22_X1 U13912 ( .A1(n11039), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n11044), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n11036) );
  NAND2_X1 U13913 ( .A1(n11040), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11035) );
  NAND2_X1 U13914 ( .A1(n11036), .A2(n11035), .ZN(n14466) );
  NAND2_X1 U13915 ( .A1(n14467), .A2(n14466), .ZN(n14468) );
  AOI22_X1 U13916 ( .A1(n11039), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n11044), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n11038) );
  NAND2_X1 U13917 ( .A1(n11040), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11037) );
  AND2_X1 U13918 ( .A1(n11038), .A2(n11037), .ZN(n13915) );
  AOI22_X1 U13919 ( .A1(n11039), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n11044), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n11042) );
  NAND2_X1 U13920 ( .A1(n11040), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11041) );
  AND2_X1 U13921 ( .A1(n11042), .A2(n11041), .ZN(n11270) );
  NOR2_X2 U13922 ( .A1(n9666), .A2(n11270), .ZN(n11269) );
  INV_X1 U13923 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n11152) );
  OR2_X1 U13924 ( .A1(n11043), .A2(n10849), .ZN(n11046) );
  NAND2_X1 U13925 ( .A1(n11044), .A2(P2_EAX_REG_31__SCAN_IN), .ZN(n11045) );
  OAI211_X1 U13926 ( .C1(n11047), .C2(n11152), .A(n11046), .B(n11045), .ZN(
        n11048) );
  XNOR2_X1 U13927 ( .A(n11269), .B(n11048), .ZN(n13890) );
  INV_X1 U13928 ( .A(n13890), .ZN(n18876) );
  NOR2_X1 U13929 ( .A1(n14979), .A2(n11050), .ZN(n16089) );
  NOR2_X1 U13930 ( .A1(n16086), .A2(n12874), .ZN(n11051) );
  OR2_X1 U13931 ( .A1(n16089), .A2(n11051), .ZN(n11052) );
  NAND2_X1 U13932 ( .A1(n11054), .A2(n11053), .ZN(n11202) );
  NAND2_X1 U13933 ( .A1(n11155), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11060) );
  INV_X1 U13934 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n11057) );
  NAND2_X1 U13935 ( .A1(n11141), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11056) );
  NAND2_X1 U13936 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11055) );
  OAI211_X1 U13937 ( .C1(n11148), .C2(n11057), .A(n11056), .B(n11055), .ZN(
        n11058) );
  INV_X1 U13938 ( .A(n11058), .ZN(n11059) );
  NAND2_X1 U13939 ( .A1(n11060), .A2(n11059), .ZN(n12628) );
  INV_X1 U13940 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11066) );
  INV_X1 U13941 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11064) );
  OAI22_X1 U13942 ( .A1(n11148), .A2(n11066), .B1(n11065), .B2(n11064), .ZN(
        n11068) );
  NOR2_X1 U13943 ( .A1(n11144), .A2(n16042), .ZN(n11067) );
  AOI211_X1 U13944 ( .C1(n11141), .C2(P2_EBX_REG_4__SCAN_IN), .A(n11068), .B(
        n11067), .ZN(n11069) );
  INV_X1 U13945 ( .A(n11069), .ZN(n13303) );
  INV_X1 U13946 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n11072) );
  NAND2_X1 U13947 ( .A1(n11141), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11071) );
  NAND2_X1 U13948 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11070) );
  OAI211_X1 U13949 ( .C1(n11153), .C2(n11072), .A(n11071), .B(n11070), .ZN(
        n11073) );
  AOI21_X1 U13950 ( .B1(n11155), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11073), .ZN(n12953) );
  NAND2_X1 U13951 ( .A1(n11141), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11075) );
  NAND2_X1 U13952 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11074) );
  OAI211_X1 U13953 ( .C1(n11148), .C2(n19532), .A(n11075), .B(n11074), .ZN(
        n11076) );
  AOI21_X1 U13954 ( .B1(n11155), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n11076), .ZN(n13040) );
  INV_X1 U13955 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n13323) );
  NAND2_X1 U13956 ( .A1(n11141), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11078) );
  NAND2_X1 U13957 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11077) );
  OAI211_X1 U13958 ( .C1(n11153), .C2(n13323), .A(n11078), .B(n11077), .ZN(
        n11079) );
  AOI21_X1 U13959 ( .B1(n11155), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n11079), .ZN(n13319) );
  INV_X1 U13960 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11083) );
  NAND2_X1 U13961 ( .A1(n11155), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11082) );
  AOI22_X1 U13962 ( .A1(n11080), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11081) );
  OAI211_X1 U13963 ( .C1(n11083), .C2(n11063), .A(n11082), .B(n11081), .ZN(
        n13108) );
  NAND2_X1 U13964 ( .A1(n11155), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11085) );
  AOI22_X1 U13965 ( .A1(n11080), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11084) );
  OAI211_X1 U13966 ( .C1(n11063), .C2(n18858), .A(n11085), .B(n11084), .ZN(
        n15898) );
  NAND2_X1 U13967 ( .A1(n11141), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11087) );
  NAND2_X1 U13968 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11086) );
  OAI211_X1 U13969 ( .C1(n11148), .C2(n11088), .A(n11087), .B(n11086), .ZN(
        n11089) );
  NAND2_X1 U13970 ( .A1(n11155), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11095) );
  INV_X1 U13971 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n11092) );
  NAND2_X1 U13972 ( .A1(n11141), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11091) );
  NAND2_X1 U13973 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11090) );
  OAI211_X1 U13974 ( .C1(n11148), .C2(n11092), .A(n11091), .B(n11090), .ZN(
        n11093) );
  INV_X1 U13975 ( .A(n11093), .ZN(n11094) );
  NAND2_X1 U13976 ( .A1(n11095), .A2(n11094), .ZN(n15875) );
  INV_X1 U13977 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n11098) );
  NAND2_X1 U13978 ( .A1(n11141), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11097) );
  NAND2_X1 U13979 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11096) );
  OAI211_X1 U13980 ( .C1(n11148), .C2(n11098), .A(n11097), .B(n11096), .ZN(
        n11099) );
  AOI21_X1 U13981 ( .B1(n11155), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11099), .ZN(n13408) );
  INV_X1 U13982 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n11102) );
  NAND2_X1 U13983 ( .A1(n11141), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11101) );
  NAND2_X1 U13984 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11100) );
  OAI211_X1 U13985 ( .C1(n11153), .C2(n11102), .A(n11101), .B(n11100), .ZN(
        n11103) );
  AOI21_X1 U13986 ( .B1(n11155), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11103), .ZN(n14944) );
  AOI22_X1 U13987 ( .A1(n11080), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11105) );
  NAND2_X1 U13988 ( .A1(n11141), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11104) );
  OAI211_X1 U13989 ( .C1(n11144), .C2(n15962), .A(n11105), .B(n11104), .ZN(
        n13476) );
  INV_X1 U13990 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n11108) );
  NAND2_X1 U13991 ( .A1(n11141), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11107) );
  NAND2_X1 U13992 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11106) );
  OAI211_X1 U13993 ( .C1(n11148), .C2(n11108), .A(n11107), .B(n11106), .ZN(
        n11109) );
  AOI21_X1 U13994 ( .B1(n11155), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11109), .ZN(n14726) );
  NAND2_X1 U13995 ( .A1(n11141), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11111) );
  NAND2_X1 U13996 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11110) );
  OAI211_X1 U13997 ( .C1(n11153), .C2(n19545), .A(n11111), .B(n11110), .ZN(
        n11112) );
  AOI21_X1 U13998 ( .B1(n11155), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11112), .ZN(n13549) );
  AOI22_X1 U13999 ( .A1(n11080), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11114) );
  NAND2_X1 U14000 ( .A1(n11141), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11113) );
  OAI211_X1 U14001 ( .C1(n11144), .C2(n14703), .A(n11114), .B(n11113), .ZN(
        n14896) );
  AOI22_X1 U14002 ( .A1(n11080), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11116) );
  NAND2_X1 U14003 ( .A1(n11141), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11115) );
  OAI211_X1 U14004 ( .C1(n11144), .C2(n14877), .A(n11116), .B(n11115), .ZN(
        n13634) );
  INV_X1 U14005 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19551) );
  NAND2_X1 U14006 ( .A1(n11141), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11118) );
  NAND2_X1 U14007 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11117) );
  OAI211_X1 U14008 ( .C1(n11148), .C2(n19551), .A(n11118), .B(n11117), .ZN(
        n11119) );
  AOI21_X1 U14009 ( .B1(n11155), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11119), .ZN(n14495) );
  INV_X1 U14010 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19553) );
  NAND2_X1 U14011 ( .A1(n11141), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11121) );
  NAND2_X1 U14012 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11120) );
  OAI211_X1 U14013 ( .C1(n11148), .C2(n19553), .A(n11121), .B(n11120), .ZN(
        n11122) );
  AOI21_X1 U14014 ( .B1(n11155), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11122), .ZN(n12655) );
  INV_X1 U14015 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n12613) );
  NAND2_X1 U14016 ( .A1(n11141), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11124) );
  NAND2_X1 U14017 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11123) );
  OAI211_X1 U14018 ( .C1(n11153), .C2(n12613), .A(n11124), .B(n11123), .ZN(
        n11125) );
  AOI21_X1 U14019 ( .B1(n11155), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n11125), .ZN(n12614) );
  AOI22_X1 U14020 ( .A1(n11080), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11127) );
  NAND2_X1 U14021 ( .A1(n11141), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11126) );
  OAI211_X1 U14022 ( .C1(n11144), .C2(n14839), .A(n11127), .B(n11126), .ZN(
        n12671) );
  AOI22_X1 U14023 ( .A1(n11080), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11129) );
  NAND2_X1 U14024 ( .A1(n11141), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11128) );
  OAI211_X1 U14025 ( .C1(n11144), .C2(n14830), .A(n11129), .B(n11128), .ZN(
        n14550) );
  INV_X1 U14026 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19560) );
  INV_X1 U14027 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14647) );
  OAI22_X1 U14028 ( .A1(n11148), .A2(n19560), .B1(n11065), .B2(n14647), .ZN(
        n11131) );
  NOR2_X1 U14029 ( .A1(n11063), .A2(n20797), .ZN(n11130) );
  NOR2_X1 U14030 ( .A1(n11131), .A2(n11130), .ZN(n11132) );
  OAI21_X1 U14031 ( .B1(n11144), .B2(n14817), .A(n11132), .ZN(n14478) );
  NAND2_X1 U14032 ( .A1(n14552), .A2(n14478), .ZN(n14538) );
  INV_X1 U14033 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n15790) );
  NAND2_X1 U14034 ( .A1(n11141), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11134) );
  NAND2_X1 U14035 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11133) );
  OAI211_X1 U14036 ( .C1(n11148), .C2(n15790), .A(n11134), .B(n11133), .ZN(
        n11135) );
  AOI21_X1 U14037 ( .B1(n11155), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11135), .ZN(n14539) );
  INV_X1 U14038 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20763) );
  NAND2_X1 U14039 ( .A1(n11141), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11137) );
  NAND2_X1 U14040 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11136) );
  OAI211_X1 U14041 ( .C1(n11148), .C2(n20763), .A(n11137), .B(n11136), .ZN(
        n11138) );
  AOI21_X1 U14042 ( .B1(n11155), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11138), .ZN(n12643) );
  AOI22_X1 U14043 ( .A1(n11080), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11140) );
  NAND2_X1 U14044 ( .A1(n11141), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11139) );
  OAI211_X1 U14045 ( .C1(n11144), .C2(n20809), .A(n11140), .B(n11139), .ZN(
        n14464) );
  AOI22_X1 U14046 ( .A1(n11080), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11143) );
  NAND2_X1 U14047 ( .A1(n11141), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11142) );
  OAI211_X1 U14048 ( .C1(n11144), .C2(n14772), .A(n11143), .B(n11142), .ZN(
        n14515) );
  INV_X1 U14049 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n11147) );
  NAND2_X1 U14050 ( .A1(n11141), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11146) );
  NAND2_X1 U14051 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11145) );
  OAI211_X1 U14052 ( .C1(n11148), .C2(n11147), .A(n11146), .B(n11145), .ZN(
        n11149) );
  AOI21_X1 U14053 ( .B1(n11155), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11149), .ZN(n11265) );
  NAND2_X1 U14054 ( .A1(n11141), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n11151) );
  NAND2_X1 U14055 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11150) );
  OAI211_X1 U14056 ( .C1(n11153), .C2(n11152), .A(n11151), .B(n11150), .ZN(
        n11154) );
  AOI21_X1 U14057 ( .B1(n11155), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n11154), .ZN(n11156) );
  INV_X1 U14058 ( .A(n11156), .ZN(n11157) );
  NAND2_X1 U14059 ( .A1(n15006), .A2(n12874), .ZN(n11159) );
  NAND2_X1 U14060 ( .A1(n11159), .A2(n12973), .ZN(n11160) );
  NAND2_X1 U14061 ( .A1(n11182), .A2(n16091), .ZN(n12938) );
  MUX2_X1 U14062 ( .A(n11164), .B(n11163), .S(n11272), .Z(n11174) );
  AOI21_X1 U14063 ( .B1(n9782), .B2(n11166), .A(n14452), .ZN(n11173) );
  AND2_X1 U14064 ( .A1(n11167), .A2(n11168), .ZN(n11170) );
  OAI21_X1 U14065 ( .B1(n11581), .B2(n11170), .A(n11169), .ZN(n11171) );
  INV_X1 U14066 ( .A(n11171), .ZN(n11172) );
  NOR3_X1 U14067 ( .A1(n11174), .A2(n11173), .A3(n11172), .ZN(n11179) );
  NAND2_X1 U14068 ( .A1(n11175), .A2(n12686), .ZN(n14980) );
  NAND2_X1 U14069 ( .A1(n14980), .A2(n11176), .ZN(n11177) );
  NAND2_X1 U14070 ( .A1(n11177), .A2(n18965), .ZN(n11178) );
  NAND2_X1 U14071 ( .A1(n14978), .A2(n11167), .ZN(n11180) );
  NAND2_X1 U14072 ( .A1(n11182), .A2(n11180), .ZN(n14910) );
  NOR2_X1 U14073 ( .A1(n16043), .A2(n16042), .ZN(n16041) );
  INV_X1 U14074 ( .A(n16041), .ZN(n11184) );
  INV_X1 U14075 ( .A(n14973), .ZN(n14940) );
  NOR2_X1 U14077 ( .A1(n11182), .A2(n18933), .ZN(n14968) );
  NAND2_X1 U14078 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14972) );
  NAND2_X1 U14079 ( .A1(n11194), .A2(n14972), .ZN(n12946) );
  NOR2_X1 U14080 ( .A1(n12938), .A2(n12946), .ZN(n12943) );
  INV_X1 U14081 ( .A(n14972), .ZN(n11183) );
  AOI21_X1 U14082 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n11183), .A(
        n14910), .ZN(n12947) );
  NOR3_X1 U14083 ( .A1(n14968), .A2(n12943), .A3(n12947), .ZN(n16066) );
  OAI21_X1 U14084 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14940), .A(
        n16066), .ZN(n16036) );
  AOI21_X1 U14085 ( .B1(n14973), .B2(n11184), .A(n16036), .ZN(n16007) );
  OR3_X1 U14086 ( .A1(n16023), .A2(n16013), .A3(n16012), .ZN(n11196) );
  NAND2_X1 U14087 ( .A1(n14973), .A2(n11196), .ZN(n11185) );
  AOI21_X1 U14088 ( .B1(n14973), .B2(n11186), .A(n14830), .ZN(n11187) );
  AND2_X1 U14089 ( .A1(n15977), .A2(n11187), .ZN(n14828) );
  AND2_X1 U14090 ( .A1(n16007), .A2(n14940), .ZN(n11188) );
  OR2_X1 U14091 ( .A1(n14828), .A2(n11188), .ZN(n14815) );
  INV_X1 U14092 ( .A(n11188), .ZN(n11190) );
  AND2_X1 U14093 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11198) );
  INV_X1 U14094 ( .A(n11198), .ZN(n11189) );
  NAND2_X1 U14095 ( .A1(n11190), .A2(n11189), .ZN(n11191) );
  NAND3_X1 U14096 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14758) );
  NAND2_X1 U14097 ( .A1(n14973), .A2(n14758), .ZN(n11192) );
  NAND2_X1 U14098 ( .A1(n14788), .A2(n11192), .ZN(n14753) );
  AOI21_X1 U14099 ( .B1(n14761), .B2(n14973), .A(n14753), .ZN(n11193) );
  NOR2_X1 U14100 ( .A1(n11194), .A2(n14972), .ZN(n11195) );
  INV_X1 U14101 ( .A(n12938), .ZN(n14907) );
  OAI211_X1 U14102 ( .C1(n11195), .C2(n14907), .A(n12946), .B(n14973), .ZN(
        n16068) );
  NAND2_X1 U14103 ( .A1(n16041), .A2(n16039), .ZN(n16011) );
  NAND2_X1 U14104 ( .A1(n16000), .A2(n11197), .ZN(n14829) );
  NOR2_X1 U14105 ( .A1(n14829), .A2(n14830), .ZN(n14818) );
  NAND2_X1 U14106 ( .A1(n14818), .A2(n11198), .ZN(n14780) );
  AND2_X1 U14107 ( .A1(n11199), .A2(n10114), .ZN(n11200) );
  NAND2_X1 U14108 ( .A1(n11204), .A2(n11203), .ZN(P2_U3015) );
  NAND2_X1 U14109 ( .A1(n19617), .A2(n16111), .ZN(n11205) );
  NAND2_X1 U14110 ( .A1(n11206), .A2(n11205), .ZN(n11207) );
  NAND2_X1 U14111 ( .A1(n11207), .A2(n16106), .ZN(n18645) );
  NAND2_X1 U14112 ( .A1(n11208), .A2(n18936), .ZN(n11225) );
  INV_X1 U14113 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11218) );
  NOR2_X1 U14114 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12980) );
  OR2_X1 U14115 ( .A1(n19390), .A2(n12980), .ZN(n19604) );
  NAND2_X1 U14116 ( .A1(n19604), .A2(n18640), .ZN(n11209) );
  OR2_X1 U14117 ( .A1(n18645), .A2(n12686), .ZN(n15941) );
  INV_X1 U14118 ( .A(n11308), .ZN(n11213) );
  INV_X1 U14119 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19294) );
  NAND2_X1 U14120 ( .A1(n19294), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11212) );
  NAND2_X1 U14121 ( .A1(n11213), .A2(n11212), .ZN(n12782) );
  AND2_X1 U14122 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11214) );
  OR2_X1 U14123 ( .A1(n11215), .A2(n13605), .ZN(n11216) );
  INV_X1 U14124 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11250) );
  NAND2_X1 U14125 ( .A1(n11249), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11245) );
  INV_X1 U14126 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11247) );
  NAND2_X1 U14127 ( .A1(n11246), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11243) );
  INV_X1 U14128 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18676) );
  NAND2_X1 U14129 ( .A1(n11244), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11241) );
  INV_X1 U14130 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14710) );
  NAND2_X1 U14131 ( .A1(n11240), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11238) );
  INV_X1 U14132 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14683) );
  INV_X1 U14133 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14659) );
  NAND2_X1 U14134 ( .A1(n11232), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11231) );
  INV_X1 U14135 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14629) );
  INV_X1 U14136 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15775) );
  INV_X1 U14137 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11261) );
  XNOR2_X1 U14138 ( .A(n11217), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11226) );
  INV_X1 U14139 ( .A(n11219), .ZN(n11223) );
  AND2_X1 U14140 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n11220) );
  NAND2_X1 U14141 ( .A1(n11225), .A2(n11224), .ZN(P2_U2983) );
  INV_X1 U14142 ( .A(n11262), .ZN(n11228) );
  AOI21_X1 U14143 ( .B1(n15775), .B2(n11227), .A(n11228), .ZN(n15773) );
  OAI21_X1 U14144 ( .B1(n11229), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n11227), .ZN(n11230) );
  INV_X1 U14145 ( .A(n11230), .ZN(n14624) );
  AOI21_X1 U14146 ( .B1(n14629), .B2(n11233), .A(n11229), .ZN(n14627) );
  OAI21_X1 U14147 ( .B1(n11232), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n11233), .ZN(n14637) );
  INV_X1 U14148 ( .A(n14637), .ZN(n15787) );
  AOI21_X1 U14149 ( .B1(n14647), .B2(n11234), .A(n11232), .ZN(n14651) );
  OAI21_X1 U14150 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n9722), .A(
        n11234), .ZN(n15854) );
  INV_X1 U14151 ( .A(n15854), .ZN(n15806) );
  AOI21_X1 U14152 ( .B1(n14659), .B2(n11235), .A(n9722), .ZN(n14661) );
  OR2_X1 U14153 ( .A1(n11236), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11237) );
  NAND2_X1 U14154 ( .A1(n11235), .A2(n11237), .ZN(n13869) );
  INV_X1 U14155 ( .A(n13869), .ZN(n15381) );
  AOI21_X1 U14156 ( .B1(n11239), .B2(n14683), .A(n11236), .ZN(n14685) );
  OAI21_X1 U14157 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n11240), .A(
        n11239), .ZN(n14698) );
  INV_X1 U14158 ( .A(n14698), .ZN(n14491) );
  AOI21_X1 U14159 ( .B1(n14710), .B2(n11242), .A(n11240), .ZN(n14713) );
  AOI21_X1 U14160 ( .B1(n18676), .B2(n11243), .A(n11244), .ZN(n18682) );
  AOI21_X1 U14161 ( .B1(n11247), .B2(n11245), .A(n11246), .ZN(n18704) );
  AOI21_X1 U14162 ( .B1(n11250), .B2(n11248), .A(n11249), .ZN(n14748) );
  AOI21_X1 U14163 ( .B1(n15888), .B2(n9653), .A(n11251), .ZN(n18741) );
  AOI21_X1 U14164 ( .B1(n15917), .B2(n11258), .A(n11260), .ZN(n18763) );
  NOR2_X1 U14165 ( .A1(n13605), .A2(n11252), .ZN(n11259) );
  AOI21_X1 U14166 ( .B1(n13605), .B2(n11252), .A(n11259), .ZN(n18770) );
  INV_X1 U14167 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n15946) );
  AND2_X1 U14168 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n11253), .ZN(
        n11257) );
  AOI21_X1 U14169 ( .B1(n15946), .B2(n11255), .A(n11257), .ZN(n18803) );
  AOI21_X1 U14170 ( .B1(n15958), .B2(n11254), .A(n11256), .ZN(n15947) );
  OAI22_X1 U14171 ( .A1(n18640), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n18831) );
  INV_X1 U14172 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13465) );
  OAI22_X1 U14173 ( .A1(n18640), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13465), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13461) );
  AND2_X1 U14174 ( .A1(n18831), .A2(n13461), .ZN(n13447) );
  OAI21_X1 U14175 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n11254), .ZN(n13449) );
  NAND2_X1 U14176 ( .A1(n13447), .A2(n13449), .ZN(n13265) );
  OAI21_X1 U14177 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n11256), .A(
        n11255), .ZN(n18943) );
  OAI21_X1 U14178 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n11257), .A(
        n11252), .ZN(n18787) );
  NOR2_X1 U14179 ( .A1(n18770), .A2(n18769), .ZN(n13315) );
  OAI21_X1 U14180 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n11259), .A(
        n11258), .ZN(n15930) );
  NAND2_X1 U14181 ( .A1(n13315), .A2(n15930), .ZN(n18761) );
  NOR2_X1 U14182 ( .A1(n18763), .A2(n18761), .ZN(n18747) );
  OAI21_X1 U14183 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n11260), .A(
        n9653), .ZN(n18749) );
  NAND2_X1 U14184 ( .A1(n18747), .A2(n18749), .ZN(n18739) );
  OAI21_X1 U14185 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n11251), .A(
        n11248), .ZN(n18728) );
  OAI21_X1 U14186 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n11249), .A(
        n11245), .ZN(n18716) );
  NOR2_X1 U14187 ( .A1(n18704), .A2(n18703), .ZN(n18690) );
  OAI21_X1 U14188 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11246), .A(
        n11243), .ZN(n18691) );
  NAND2_X1 U14189 ( .A1(n18690), .A2(n18691), .ZN(n18681) );
  OAI21_X1 U14190 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n11244), .A(
        n11242), .ZN(n18665) );
  NOR2_X1 U14191 ( .A1(n14491), .A2(n14490), .ZN(n14489) );
  NOR2_X1 U14192 ( .A1(n18785), .A2(n14489), .ZN(n12653) );
  NOR2_X1 U14193 ( .A1(n14685), .A2(n12653), .ZN(n12652) );
  NOR2_X1 U14194 ( .A1(n18785), .A2(n12652), .ZN(n15380) );
  NOR2_X1 U14195 ( .A1(n15381), .A2(n15380), .ZN(n15379) );
  NOR2_X1 U14196 ( .A1(n18785), .A2(n15379), .ZN(n12667) );
  NOR2_X1 U14197 ( .A1(n14661), .A2(n12667), .ZN(n12666) );
  NOR2_X1 U14198 ( .A1(n18785), .A2(n12666), .ZN(n15805) );
  NOR2_X1 U14199 ( .A1(n15787), .A2(n15786), .ZN(n15785) );
  NOR2_X1 U14200 ( .A1(n18785), .A2(n15785), .ZN(n12640) );
  NOR2_X1 U14201 ( .A1(n14627), .A2(n12640), .ZN(n12639) );
  NOR2_X1 U14202 ( .A1(n18785), .A2(n15772), .ZN(n11263) );
  XNOR2_X1 U14203 ( .A(n11262), .B(n11261), .ZN(n13885) );
  XNOR2_X1 U14204 ( .A(n11263), .B(n13885), .ZN(n11264) );
  NOR4_X4 U14205 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n11065), .ZN(n19499) );
  NAND2_X1 U14206 ( .A1(n11264), .A2(n19499), .ZN(n11289) );
  INV_X1 U14207 ( .A(n19504), .ZN(n19520) );
  NOR2_X1 U14208 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19520), .ZN(n11271) );
  INV_X1 U14209 ( .A(n11271), .ZN(n11266) );
  NOR2_X1 U14210 ( .A1(n11267), .A2(n11266), .ZN(n11268) );
  NAND2_X1 U14211 ( .A1(n18642), .A2(n11268), .ZN(n18789) );
  AOI21_X1 U14212 ( .B1(n11270), .B2(n9666), .A(n11269), .ZN(n14755) );
  NAND2_X1 U14213 ( .A1(n18642), .A2(n14454), .ZN(n11274) );
  NAND2_X1 U14214 ( .A1(n19510), .A2(n11271), .ZN(n16107) );
  OR2_X2 U14215 ( .A1(n11274), .A2(n16107), .ZN(n18812) );
  INV_X1 U14216 ( .A(n18812), .ZN(n15802) );
  OAI211_X1 U14217 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n19520), .A(n18642), 
        .B(n11272), .ZN(n11279) );
  OR2_X1 U14218 ( .A1(n11279), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n11275) );
  INV_X1 U14219 ( .A(n16107), .ZN(n11273) );
  OR2_X1 U14220 ( .A1(n11274), .A2(n11273), .ZN(n13886) );
  AOI22_X1 U14221 ( .A1(n14755), .A2(n15802), .B1(P2_EBX_REG_30__SCAN_IN), 
        .B2(n18819), .ZN(n11276) );
  OAI21_X1 U14222 ( .B1(n14759), .B2(n18789), .A(n11276), .ZN(n11277) );
  INV_X1 U14223 ( .A(n11277), .ZN(n11287) );
  NAND2_X1 U14224 ( .A1(n12686), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n11278) );
  NAND2_X1 U14225 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19606), .ZN(n18992) );
  NOR2_X1 U14226 ( .A1(n11280), .A2(n18992), .ZN(n16110) );
  NAND2_X1 U14227 ( .A1(n16010), .A2(n18779), .ZN(n11281) );
  OR2_X1 U14228 ( .A1(n16110), .A2(n11281), .ZN(n11282) );
  AOI22_X1 U14229 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n9607), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n18669), .ZN(n11283) );
  OAI21_X1 U14230 ( .B1(n11284), .B2(n18795), .A(n11283), .ZN(n11285) );
  INV_X1 U14231 ( .A(n11285), .ZN(n11286) );
  NAND2_X1 U14232 ( .A1(n11289), .A2(n11288), .ZN(P2_U2825) );
  NAND2_X1 U14233 ( .A1(n15954), .A2(n11308), .ZN(n11294) );
  OAI21_X1 U14234 ( .B1(n18971), .B2(n18640), .A(n19582), .ZN(n11305) );
  NAND2_X1 U14235 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19387) );
  INV_X1 U14236 ( .A(n19387), .ZN(n19437) );
  AND2_X1 U14237 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19437), .ZN(
        n11291) );
  NAND2_X1 U14238 ( .A1(n11291), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19441) );
  INV_X1 U14239 ( .A(n11291), .ZN(n11298) );
  NAND2_X1 U14240 ( .A1(n19588), .A2(n11298), .ZN(n11292) );
  AND3_X1 U14241 ( .A1(n19441), .A2(n19390), .A3(n11292), .ZN(n19322) );
  AOI21_X1 U14242 ( .B1(n11305), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19322), .ZN(n11293) );
  NAND2_X1 U14243 ( .A1(n11294), .A2(n11293), .ZN(n11296) );
  AND2_X1 U14244 ( .A1(n18971), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12837) );
  NAND2_X1 U14245 ( .A1(n12837), .A2(n12686), .ZN(n11513) );
  INV_X1 U14246 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18970) );
  NOR2_X1 U14247 ( .A1(n11513), .A2(n18970), .ZN(n11295) );
  OR2_X1 U14248 ( .A1(n11296), .A2(n11295), .ZN(n11297) );
  NAND2_X1 U14249 ( .A1(n11296), .A2(n11295), .ZN(n11317) );
  INV_X1 U14250 ( .A(n19390), .ZN(n19393) );
  NAND2_X1 U14251 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19288) );
  NAND2_X1 U14252 ( .A1(n19288), .A2(n19596), .ZN(n11299) );
  NAND2_X1 U14253 ( .A1(n11299), .A2(n11298), .ZN(n19076) );
  NOR2_X1 U14254 ( .A1(n19393), .A2(n19076), .ZN(n11300) );
  AOI21_X1 U14255 ( .B1(n11305), .B2(n15019), .A(n11300), .ZN(n11301) );
  NAND2_X1 U14256 ( .A1(n11490), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11312) );
  AOI22_X1 U14257 ( .A1(n11305), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19390), .B2(n19613), .ZN(n11303) );
  NAND2_X1 U14258 ( .A1(n11490), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11309) );
  NAND2_X1 U14259 ( .A1(n11305), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11306) );
  NAND2_X1 U14260 ( .A1(n19603), .A2(n19613), .ZN(n19195) );
  NAND3_X1 U14261 ( .A1(n19390), .A2(n19195), .A3(n19288), .ZN(n19259) );
  NAND2_X1 U14262 ( .A1(n11306), .A2(n19259), .ZN(n11307) );
  INV_X1 U14263 ( .A(n11309), .ZN(n11310) );
  NOR2_X1 U14264 ( .A1(n14983), .A2(n11310), .ZN(n11311) );
  INV_X1 U14265 ( .A(n11312), .ZN(n11313) );
  NAND2_X1 U14266 ( .A1(n11314), .A2(n11313), .ZN(n11315) );
  NAND2_X1 U14267 ( .A1(n11600), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11316) );
  INV_X1 U14268 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11319) );
  NAND2_X1 U14269 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12967) );
  NOR2_X1 U14270 ( .A1(n11319), .A2(n12967), .ZN(n18862) );
  AND2_X1 U14271 ( .A1(n18860), .A2(n18862), .ZN(n11321) );
  INV_X1 U14272 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11320) );
  NOR2_X1 U14273 ( .A1(n11513), .A2(n11320), .ZN(n18861) );
  AND2_X1 U14274 ( .A1(n18837), .A2(n18838), .ZN(n11323) );
  AOI22_X1 U14275 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11329) );
  AOI22_X1 U14276 ( .A1(n10449), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11328) );
  AOI22_X1 U14277 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11327) );
  AOI22_X1 U14278 ( .A1(n11417), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11326) );
  NAND4_X1 U14279 ( .A1(n11329), .A2(n11328), .A3(n11327), .A4(n11326), .ZN(
        n11335) );
  AOI22_X1 U14280 ( .A1(n10504), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9616), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14281 ( .A1(n10454), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14282 ( .A1(n10415), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14283 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11330) );
  NAND4_X1 U14284 ( .A1(n11333), .A2(n11332), .A3(n11331), .A4(n11330), .ZN(
        n11334) );
  NOR2_X1 U14285 ( .A1(n11335), .A2(n11334), .ZN(n18834) );
  INV_X1 U14286 ( .A(n18834), .ZN(n11336) );
  AOI22_X1 U14287 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10794), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11340) );
  AOI22_X1 U14288 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10449), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11339) );
  AOI22_X1 U14289 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11338) );
  AOI22_X1 U14290 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11417), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11337) );
  NAND4_X1 U14291 ( .A1(n11340), .A2(n11339), .A3(n11338), .A4(n11337), .ZN(
        n11346) );
  AOI22_X1 U14292 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n9616), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11344) );
  AOI22_X1 U14293 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10454), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14294 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10415), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14295 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10413), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11341) );
  NAND4_X1 U14296 ( .A1(n11344), .A2(n11343), .A3(n11342), .A4(n11341), .ZN(
        n11345) );
  NOR2_X1 U14297 ( .A1(n11346), .A2(n11345), .ZN(n13553) );
  AOI22_X1 U14298 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10794), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U14299 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n10449), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11349) );
  AOI22_X1 U14300 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11348) );
  AOI22_X1 U14301 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n11417), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11347) );
  NAND4_X1 U14302 ( .A1(n11350), .A2(n11349), .A3(n11348), .A4(n11347), .ZN(
        n11356) );
  AOI22_X1 U14303 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n9616), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14304 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10454), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14305 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10415), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14306 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10413), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11351) );
  NAND4_X1 U14307 ( .A1(n11354), .A2(n11353), .A3(n11352), .A4(n11351), .ZN(
        n11355) );
  OR2_X1 U14308 ( .A1(n11356), .A2(n11355), .ZN(n15823) );
  AOI22_X1 U14309 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10794), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11360) );
  AOI22_X1 U14310 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10449), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U14311 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14312 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n11417), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11357) );
  NAND4_X1 U14313 ( .A1(n11360), .A2(n11359), .A3(n11358), .A4(n11357), .ZN(
        n11366) );
  AOI22_X1 U14314 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n9616), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U14315 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10454), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14316 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10415), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U14317 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10413), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11361) );
  NAND4_X1 U14318 ( .A1(n11364), .A2(n11363), .A3(n11362), .A4(n11361), .ZN(
        n11365) );
  AOI22_X1 U14319 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10794), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U14320 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10449), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11370) );
  AOI22_X1 U14321 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U14322 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11417), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11368) );
  NAND4_X1 U14323 ( .A1(n11371), .A2(n11370), .A3(n11369), .A4(n11368), .ZN(
        n11377) );
  AOI22_X1 U14324 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n9616), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14325 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10454), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14326 ( .A1(n10415), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11373) );
  AOI22_X1 U14327 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10413), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11372) );
  NAND4_X1 U14328 ( .A1(n11375), .A2(n11374), .A3(n11373), .A4(n11372), .ZN(
        n11376) );
  NOR2_X1 U14329 ( .A1(n11377), .A2(n11376), .ZN(n15820) );
  AOI22_X1 U14330 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11381) );
  AOI22_X1 U14331 ( .A1(n10449), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11380) );
  AOI22_X1 U14332 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11379) );
  AOI22_X1 U14333 ( .A1(n11417), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11378) );
  NAND4_X1 U14334 ( .A1(n11381), .A2(n11380), .A3(n11379), .A4(n11378), .ZN(
        n11387) );
  AOI22_X1 U14335 ( .A1(n10504), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9616), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11385) );
  AOI22_X1 U14336 ( .A1(n10454), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11384) );
  AOI22_X1 U14337 ( .A1(n10415), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14338 ( .A1(n10413), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11382) );
  NAND4_X1 U14339 ( .A1(n11385), .A2(n11384), .A3(n11383), .A4(n11382), .ZN(
        n11386) );
  OR2_X1 U14340 ( .A1(n11387), .A2(n11386), .ZN(n13670) );
  AOI22_X1 U14341 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14342 ( .A1(n10794), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__6__SCAN_IN), .B2(n10901), .ZN(n11390) );
  AOI22_X1 U14343 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n11417), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U14344 ( .A1(n10449), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n10511), .ZN(n11388) );
  NAND4_X1 U14345 ( .A1(n11391), .A2(n11390), .A3(n11389), .A4(n11388), .ZN(
        n11397) );
  AOI22_X1 U14346 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10454), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14347 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10417), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11394) );
  AOI22_X1 U14348 ( .A1(n10415), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n10416), .ZN(n11393) );
  AOI22_X1 U14349 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10413), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11392) );
  NAND4_X1 U14350 ( .A1(n11395), .A2(n11394), .A3(n11393), .A4(n11392), .ZN(
        n11396) );
  NOR2_X1 U14351 ( .A1(n11397), .A2(n11396), .ZN(n15817) );
  AOI22_X1 U14352 ( .A1(n10221), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11563), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11407) );
  INV_X1 U14353 ( .A(n11399), .ZN(n15000) );
  AOI22_X1 U14354 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15000), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11405) );
  AND2_X1 U14355 ( .A1(n15019), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11401) );
  OR2_X1 U14356 ( .A1(n11401), .A2(n11400), .ZN(n11568) );
  INV_X1 U14357 ( .A(n11568), .ZN(n11537) );
  NAND2_X1 U14358 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11403) );
  NAND2_X1 U14359 ( .A1(n11566), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11402) );
  AND3_X1 U14360 ( .A1(n11537), .A2(n11403), .A3(n11402), .ZN(n11404) );
  NAND4_X1 U14361 ( .A1(n11407), .A2(n11406), .A3(n11405), .A4(n11404), .ZN(
        n11415) );
  AOI22_X1 U14362 ( .A1(n10369), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11567), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11413) );
  NAND2_X1 U14363 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11409) );
  NAND2_X1 U14364 ( .A1(n15000), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11408) );
  AND3_X1 U14365 ( .A1(n11409), .A2(n11568), .A3(n11408), .ZN(n11412) );
  AOI22_X1 U14366 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11522), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11410) );
  NAND4_X1 U14367 ( .A1(n11413), .A2(n11412), .A3(n11411), .A4(n11410), .ZN(
        n11414) );
  NAND2_X1 U14368 ( .A1(n11415), .A2(n11414), .ZN(n11450) );
  NOR2_X1 U14369 ( .A1(n12874), .A2(n11450), .ZN(n11428) );
  AOI22_X1 U14370 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10794), .B1(
        n10901), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11421) );
  AOI22_X1 U14371 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10449), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11420) );
  AOI22_X1 U14372 ( .A1(n10483), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14373 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11417), .B1(
        n11416), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11418) );
  NAND4_X1 U14374 ( .A1(n11421), .A2(n11420), .A3(n11419), .A4(n11418), .ZN(
        n11427) );
  AOI22_X1 U14375 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n9616), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14376 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10454), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U14377 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10415), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14378 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10413), .B1(
        n10414), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11422) );
  NAND4_X1 U14379 ( .A1(n11425), .A2(n11424), .A3(n11423), .A4(n11422), .ZN(
        n11426) );
  NOR2_X1 U14380 ( .A1(n11427), .A2(n11426), .ZN(n11431) );
  XNOR2_X1 U14381 ( .A(n11428), .B(n11431), .ZN(n11452) );
  INV_X1 U14382 ( .A(n11450), .ZN(n11432) );
  NAND2_X1 U14383 ( .A1(n12874), .A2(n11432), .ZN(n14592) );
  INV_X1 U14384 ( .A(n11431), .ZN(n11433) );
  NAND2_X1 U14385 ( .A1(n11433), .A2(n11432), .ZN(n11454) );
  NAND2_X1 U14386 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11435) );
  NAND2_X1 U14387 ( .A1(n15000), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11434) );
  AND3_X1 U14388 ( .A1(n11537), .A2(n11435), .A3(n11434), .ZN(n11439) );
  AOI22_X1 U14389 ( .A1(n10369), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11567), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11438) );
  AOI22_X1 U14390 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11522), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11436) );
  NAND4_X1 U14391 ( .A1(n11439), .A2(n11438), .A3(n11437), .A4(n11436), .ZN(
        n11447) );
  AOI22_X1 U14392 ( .A1(n10369), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11567), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11445) );
  NAND2_X1 U14393 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11441) );
  NAND2_X1 U14394 ( .A1(n15000), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11440) );
  AND3_X1 U14395 ( .A1(n11441), .A2(n11568), .A3(n11440), .ZN(n11444) );
  AOI22_X1 U14396 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11522), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11442) );
  NAND4_X1 U14397 ( .A1(n11445), .A2(n11444), .A3(n11443), .A4(n11442), .ZN(
        n11446) );
  NAND2_X1 U14398 ( .A1(n11447), .A2(n11446), .ZN(n11453) );
  XOR2_X1 U14399 ( .A(n11454), .B(n11453), .Z(n11448) );
  NAND2_X1 U14400 ( .A1(n11448), .A2(n11490), .ZN(n14546) );
  INV_X1 U14401 ( .A(n11453), .ZN(n11449) );
  NAND2_X1 U14402 ( .A1(n12874), .A2(n11449), .ZN(n14549) );
  NOR2_X1 U14403 ( .A1(n14549), .A2(n11450), .ZN(n11451) );
  NOR2_X1 U14404 ( .A1(n11454), .A2(n11453), .ZN(n11469) );
  AOI22_X1 U14405 ( .A1(n10369), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11567), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11460) );
  NAND2_X1 U14406 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11456) );
  NAND2_X1 U14407 ( .A1(n15000), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11455) );
  AND3_X1 U14408 ( .A1(n11537), .A2(n11456), .A3(n11455), .ZN(n11459) );
  AOI22_X1 U14409 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11522), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11457) );
  NAND4_X1 U14410 ( .A1(n11460), .A2(n11459), .A3(n11458), .A4(n11457), .ZN(
        n11468) );
  AOI22_X1 U14411 ( .A1(n10221), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11567), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11466) );
  NAND2_X1 U14412 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11462) );
  NAND2_X1 U14413 ( .A1(n15000), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11461) );
  AND3_X1 U14414 ( .A1(n11462), .A2(n11568), .A3(n11461), .ZN(n11465) );
  AOI22_X1 U14415 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11522), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11463) );
  NAND4_X1 U14416 ( .A1(n11466), .A2(n11465), .A3(n11464), .A4(n11463), .ZN(
        n11467) );
  AND2_X1 U14417 ( .A1(n11468), .A2(n11467), .ZN(n11471) );
  NAND2_X1 U14418 ( .A1(n11469), .A2(n11471), .ZN(n11512) );
  OAI211_X1 U14419 ( .C1(n11469), .C2(n11471), .A(n11490), .B(n11512), .ZN(
        n11473) );
  INV_X1 U14420 ( .A(n11473), .ZN(n11470) );
  INV_X1 U14421 ( .A(n11471), .ZN(n11472) );
  NOR2_X1 U14422 ( .A1(n12686), .A2(n11472), .ZN(n14543) );
  AOI22_X1 U14423 ( .A1(n10369), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11567), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11481) );
  NAND2_X1 U14424 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11477) );
  NAND2_X1 U14425 ( .A1(n15000), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11476) );
  AND3_X1 U14426 ( .A1(n11537), .A2(n11477), .A3(n11476), .ZN(n11480) );
  AOI22_X1 U14427 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11522), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11478) );
  NAND4_X1 U14428 ( .A1(n11481), .A2(n11480), .A3(n11479), .A4(n11478), .ZN(
        n11489) );
  AOI22_X1 U14429 ( .A1(n10221), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11567), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11487) );
  NAND2_X1 U14430 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11483) );
  NAND2_X1 U14431 ( .A1(n15000), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11482) );
  AND3_X1 U14432 ( .A1(n11483), .A2(n11568), .A3(n11482), .ZN(n11486) );
  AOI22_X1 U14433 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11484) );
  NAND4_X1 U14434 ( .A1(n11487), .A2(n11486), .A3(n11485), .A4(n11484), .ZN(
        n11488) );
  AND2_X1 U14435 ( .A1(n11489), .A2(n11488), .ZN(n11492) );
  XNOR2_X1 U14436 ( .A(n11512), .B(n11492), .ZN(n11491) );
  NAND2_X1 U14437 ( .A1(n11491), .A2(n11490), .ZN(n11494) );
  INV_X1 U14438 ( .A(n11492), .ZN(n11511) );
  NOR2_X1 U14439 ( .A1(n12686), .A2(n11511), .ZN(n14534) );
  INV_X1 U14440 ( .A(n11494), .ZN(n11495) );
  NAND2_X1 U14441 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11498) );
  NAND2_X1 U14442 ( .A1(n15000), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11497) );
  AND3_X1 U14443 ( .A1(n11537), .A2(n11498), .A3(n11497), .ZN(n11502) );
  AOI22_X1 U14444 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9626), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11501) );
  AOI22_X1 U14445 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11499) );
  NAND4_X1 U14446 ( .A1(n11502), .A2(n11501), .A3(n11500), .A4(n11499), .ZN(
        n11510) );
  AOI22_X1 U14447 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11567), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11508) );
  NAND2_X1 U14448 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11504) );
  NAND2_X1 U14449 ( .A1(n15000), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11503) );
  AND3_X1 U14450 ( .A1(n11504), .A2(n11568), .A3(n11503), .ZN(n11507) );
  AOI22_X1 U14451 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11505) );
  NAND4_X1 U14452 ( .A1(n11508), .A2(n11507), .A3(n11506), .A4(n11505), .ZN(
        n11509) );
  NAND2_X1 U14453 ( .A1(n11510), .A2(n11509), .ZN(n11517) );
  OR2_X1 U14454 ( .A1(n11512), .A2(n11511), .ZN(n11514) );
  NOR2_X1 U14455 ( .A1(n11514), .A2(n11517), .ZN(n14521) );
  AOI211_X1 U14456 ( .C1(n11517), .C2(n11514), .A(n11513), .B(n14521), .ZN(
        n11515) );
  NAND2_X1 U14457 ( .A1(n11516), .A2(n11515), .ZN(n11519) );
  OAI21_X1 U14458 ( .B1(n11516), .B2(n11515), .A(n11519), .ZN(n14529) );
  INV_X1 U14459 ( .A(n11517), .ZN(n11518) );
  NAND2_X1 U14460 ( .A1(n12874), .A2(n11518), .ZN(n14528) );
  INV_X1 U14461 ( .A(n11519), .ZN(n14522) );
  AOI22_X1 U14462 ( .A1(n10369), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11567), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11526) );
  NAND2_X1 U14463 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11521) );
  NAND2_X1 U14464 ( .A1(n15000), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11520) );
  AND3_X1 U14465 ( .A1(n11537), .A2(n11521), .A3(n11520), .ZN(n11525) );
  AOI22_X1 U14466 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11522), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11523) );
  NAND4_X1 U14467 ( .A1(n11526), .A2(n11525), .A3(n11524), .A4(n11523), .ZN(
        n11534) );
  AOI22_X1 U14468 ( .A1(n10221), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11567), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11532) );
  NAND2_X1 U14469 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11528) );
  NAND2_X1 U14470 ( .A1(n15000), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11527) );
  AND3_X1 U14471 ( .A1(n11528), .A2(n11568), .A3(n11527), .ZN(n11531) );
  AOI22_X1 U14472 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11529) );
  NAND4_X1 U14473 ( .A1(n11532), .A2(n11531), .A3(n11530), .A4(n11529), .ZN(
        n11533) );
  AND2_X1 U14474 ( .A1(n11534), .A2(n11533), .ZN(n14523) );
  NAND2_X1 U14475 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11536) );
  NAND2_X1 U14476 ( .A1(n15000), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11535) );
  AND3_X1 U14477 ( .A1(n11537), .A2(n11536), .A3(n11535), .ZN(n11541) );
  AOI22_X1 U14478 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11538) );
  NAND4_X1 U14479 ( .A1(n11541), .A2(n11540), .A3(n11539), .A4(n11538), .ZN(
        n11549) );
  AOI22_X1 U14480 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11567), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11547) );
  NAND2_X1 U14481 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11543) );
  NAND2_X1 U14482 ( .A1(n15000), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11542) );
  AND3_X1 U14483 ( .A1(n11543), .A2(n11568), .A3(n11542), .ZN(n11546) );
  AOI22_X1 U14484 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11545) );
  NAND4_X1 U14485 ( .A1(n11547), .A2(n11546), .A3(n11545), .A4(n11544), .ZN(
        n11548) );
  NAND2_X1 U14486 ( .A1(n11549), .A2(n11548), .ZN(n11552) );
  INV_X1 U14487 ( .A(n11552), .ZN(n11555) );
  INV_X1 U14488 ( .A(n14523), .ZN(n11550) );
  NOR2_X1 U14489 ( .A1(n12874), .A2(n11550), .ZN(n11551) );
  NAND2_X1 U14490 ( .A1(n14521), .A2(n11551), .ZN(n11553) );
  INV_X1 U14491 ( .A(n11553), .ZN(n11554) );
  OR2_X1 U14492 ( .A1(n11553), .A2(n11552), .ZN(n11556) );
  OAI21_X1 U14493 ( .B1(n11555), .B2(n11554), .A(n11556), .ZN(n13913) );
  NAND2_X1 U14494 ( .A1(n11558), .A2(n11557), .ZN(n11575) );
  INV_X1 U14495 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11562) );
  AOI21_X1 U14496 ( .B1(n11559), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n11568), .ZN(n11561) );
  AOI22_X1 U14497 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11560) );
  OAI211_X1 U14498 ( .C1(n11399), .C2(n11562), .A(n11561), .B(n11560), .ZN(
        n11574) );
  AOI22_X1 U14499 ( .A1(n10182), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11563), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11565) );
  NAND2_X1 U14500 ( .A1(n11565), .A2(n11564), .ZN(n11573) );
  AOI22_X1 U14501 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11566), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11571) );
  NAND2_X1 U14502 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11570) );
  NAND2_X1 U14503 ( .A1(n15000), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11569) );
  NAND4_X1 U14504 ( .A1(n11571), .A2(n11570), .A3(n11569), .A4(n11568), .ZN(
        n11572) );
  OAI22_X1 U14505 ( .A1(n11575), .A2(n11574), .B1(n11573), .B2(n11572), .ZN(
        n11576) );
  XNOR2_X1 U14506 ( .A(n11577), .B(n11576), .ZN(n13911) );
  NAND2_X1 U14507 ( .A1(n16090), .A2(n16091), .ZN(n11580) );
  INV_X1 U14508 ( .A(n16100), .ZN(n11578) );
  NAND3_X1 U14509 ( .A1(n11578), .A2(n19504), .A3(n14452), .ZN(n11579) );
  INV_X1 U14510 ( .A(n11167), .ZN(n12842) );
  NAND2_X1 U14511 ( .A1(n11581), .A2(n12842), .ZN(n11582) );
  NAND2_X1 U14512 ( .A1(n12870), .A2(n11582), .ZN(n11583) );
  NAND2_X1 U14513 ( .A1(n14596), .A2(n11584), .ZN(n14601) );
  NOR4_X1 U14514 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n11589) );
  NOR4_X1 U14515 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n11588) );
  NOR4_X1 U14516 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n11587) );
  NOR4_X1 U14517 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n11586) );
  NAND4_X1 U14518 ( .A1(n11589), .A2(n11588), .A3(n11587), .A4(n11586), .ZN(
        n11594) );
  NOR4_X1 U14519 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n11592) );
  NOR4_X1 U14520 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n11591) );
  NOR4_X1 U14521 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n11590) );
  INV_X1 U14522 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19526) );
  NAND4_X1 U14523 ( .A1(n11592), .A2(n11591), .A3(n11590), .A4(n19526), .ZN(
        n11593) );
  OAI21_X1 U14524 ( .B1(n11594), .B2(n11593), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n11595) );
  INV_X1 U14525 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n11596) );
  OR2_X1 U14526 ( .A1(n15033), .A2(n11596), .ZN(n11598) );
  NAND2_X1 U14527 ( .A1(n15033), .A2(BUF2_REG_14__SCAN_IN), .ZN(n11597) );
  NAND2_X1 U14528 ( .A1(n11598), .A2(n11597), .ZN(n13440) );
  NAND2_X1 U14529 ( .A1(n14596), .A2(n18981), .ZN(n14585) );
  INV_X1 U14530 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n11599) );
  NAND3_X1 U14531 ( .A1(n14596), .A2(n11600), .A3(n12844), .ZN(n11601) );
  NOR2_X2 U14532 ( .A1(n11601), .A2(n15033), .ZN(n18882) );
  NOR2_X2 U14533 ( .A1(n11601), .A2(n15034), .ZN(n18881) );
  AOI22_X1 U14534 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n18882), .B1(n18881), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n11602) );
  OAI21_X1 U14535 ( .B1(n13911), .B2(n14601), .A(n11603), .ZN(P2_U2889) );
  INV_X1 U14536 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11604) );
  AND2_X4 U14537 ( .A1(n11614), .A2(n13210), .ZN(n12356) );
  AOI22_X1 U14538 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n12356), .B1(
        n11681), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11611) );
  AND2_X2 U14539 ( .A1(n11606), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11613) );
  INV_X1 U14540 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11607) );
  AND2_X2 U14541 ( .A1(n11607), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11612) );
  AOI22_X1 U14542 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n11775), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U14543 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11995), .B1(
        n12221), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11609) );
  AND2_X2 U14544 ( .A1(n11612), .A2(n13210), .ZN(n11662) );
  AND2_X4 U14545 ( .A1(n13210), .A2(n15389), .ZN(n12379) );
  AOI22_X1 U14546 ( .A1(n11662), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11608) );
  AOI22_X1 U14547 ( .A1(n11661), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11877), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11619) );
  AND2_X2 U14548 ( .A1(n11614), .A2(n11615), .ZN(n11990) );
  AND2_X2 U14549 ( .A1(n15390), .A2(n13210), .ZN(n11668) );
  AOI22_X1 U14550 ( .A1(n11990), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11668), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14551 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11682), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14552 ( .A1(n11667), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11616) );
  INV_X1 U14553 ( .A(n11676), .ZN(n11760) );
  NAND2_X1 U14554 ( .A1(n11667), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11623) );
  NAND2_X1 U14555 ( .A1(n11681), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11622) );
  NAND2_X1 U14556 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11621) );
  NAND2_X1 U14557 ( .A1(n12356), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11620) );
  NAND2_X1 U14558 ( .A1(n11682), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11627) );
  NAND2_X1 U14559 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11626) );
  NAND2_X1 U14560 ( .A1(n11661), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11625) );
  NAND2_X1 U14561 ( .A1(n11877), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11624) );
  NAND2_X1 U14562 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11631) );
  NAND2_X1 U14563 ( .A1(n11775), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11630) );
  NAND2_X1 U14564 ( .A1(n11662), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11629) );
  NAND2_X1 U14565 ( .A1(n12379), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11628) );
  NAND2_X1 U14566 ( .A1(n11990), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11635) );
  NAND2_X1 U14567 ( .A1(n11668), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11634) );
  NAND2_X1 U14568 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11633) );
  NAND2_X1 U14569 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11632) );
  NAND4_X4 U14570 ( .A1(n11639), .A2(n11638), .A3(n11637), .A4(n11636), .ZN(
        n12415) );
  AOI22_X1 U14571 ( .A1(n11775), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11643) );
  AOI22_X1 U14572 ( .A1(n11661), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11642) );
  AOI22_X1 U14573 ( .A1(n11682), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11877), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U14574 ( .A1(n11662), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11640) );
  NAND4_X1 U14575 ( .A1(n11643), .A2(n11642), .A3(n11641), .A4(n11640), .ZN(
        n11649) );
  AOI22_X1 U14576 ( .A1(n12356), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12221), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14577 ( .A1(n11990), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11668), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14578 ( .A1(n11667), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11681), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14579 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11644) );
  NAND4_X1 U14580 ( .A1(n11647), .A2(n11646), .A3(n11645), .A4(n11644), .ZN(
        n11648) );
  NAND2_X1 U14582 ( .A1(n12962), .A2(n19868), .ZN(n11763) );
  AOI22_X1 U14583 ( .A1(n11667), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11681), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14584 ( .A1(n12356), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11775), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14585 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11877), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14586 ( .A1(n11662), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11650) );
  NAND4_X1 U14587 ( .A1(n11653), .A2(n11652), .A3(n11651), .A4(n11650), .ZN(
        n11659) );
  AOI22_X1 U14588 ( .A1(n11682), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11661), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14589 ( .A1(n11990), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11668), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U14590 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12221), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11655) );
  AOI22_X1 U14591 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11654) );
  NAND4_X1 U14592 ( .A1(n11657), .A2(n11656), .A3(n11655), .A4(n11654), .ZN(
        n11658) );
  AOI22_X1 U14593 ( .A1(n11775), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11666) );
  AOI22_X1 U14594 ( .A1(n11661), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11665) );
  AOI22_X1 U14595 ( .A1(n11682), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11877), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14596 ( .A1(n11662), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11663) );
  NAND4_X1 U14597 ( .A1(n11666), .A2(n11665), .A3(n11664), .A4(n11663), .ZN(
        n11674) );
  AOI22_X1 U14598 ( .A1(n11667), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11681), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14599 ( .A1(n11990), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11668), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U14600 ( .A1(n9611), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12221), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U14601 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11669) );
  NAND4_X1 U14602 ( .A1(n11672), .A2(n11671), .A3(n11670), .A4(n11669), .ZN(
        n11673) );
  OR2_X2 U14603 ( .A1(n11674), .A2(n11673), .ZN(n11737) );
  NAND2_X1 U14604 ( .A1(n11737), .A2(n11844), .ZN(n11738) );
  NAND2_X1 U14605 ( .A1(n13054), .A2(n11738), .ZN(n11675) );
  AND2_X1 U14606 ( .A1(n11676), .A2(n12415), .ZN(n11689) );
  AOI22_X1 U14607 ( .A1(n11667), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14608 ( .A1(n11775), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14609 ( .A1(n11990), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11668), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14610 ( .A1(n11662), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11677) );
  NAND4_X1 U14611 ( .A1(n11680), .A2(n11679), .A3(n11678), .A4(n11677), .ZN(
        n11688) );
  AOI22_X1 U14612 ( .A1(n11681), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9612), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U14613 ( .A1(n11661), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11877), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U14614 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12221), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11684) );
  AOI22_X1 U14615 ( .A1(n11682), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11683) );
  NAND4_X1 U14616 ( .A1(n11686), .A2(n11685), .A3(n11684), .A4(n11683), .ZN(
        n11687) );
  NAND2_X1 U14617 ( .A1(n11990), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11694) );
  NAND2_X1 U14618 ( .A1(n11667), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11693) );
  NAND2_X1 U14619 ( .A1(n11681), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11692) );
  NAND2_X1 U14620 ( .A1(n11668), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11691) );
  NAND2_X1 U14621 ( .A1(n11775), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11698) );
  NAND2_X1 U14622 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11697) );
  NAND2_X1 U14623 ( .A1(n11682), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11696) );
  NAND2_X1 U14624 ( .A1(n11877), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11695) );
  NAND2_X1 U14625 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11703) );
  NAND2_X1 U14626 ( .A1(n12356), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11702) );
  NAND2_X1 U14627 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11701) );
  NAND2_X1 U14628 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11700) );
  NAND2_X1 U14629 ( .A1(n11661), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11707) );
  NAND2_X1 U14630 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11706) );
  NAND2_X1 U14631 ( .A1(n11662), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11705) );
  NAND2_X1 U14632 ( .A1(n12379), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11704) );
  NOR2_X1 U14633 ( .A1(n11690), .A2(n9618), .ZN(n11711) );
  NAND2_X1 U14634 ( .A1(n11990), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11715) );
  NAND2_X1 U14635 ( .A1(n11667), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11714) );
  NAND2_X1 U14636 ( .A1(n11681), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11713) );
  NAND2_X1 U14637 ( .A1(n11668), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11712) );
  NAND2_X1 U14638 ( .A1(n12356), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11719) );
  NAND2_X1 U14639 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11718) );
  NAND2_X1 U14640 ( .A1(n11682), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11717) );
  NAND2_X1 U14641 ( .A1(n12221), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11716) );
  NAND2_X1 U14642 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11723) );
  NAND2_X1 U14643 ( .A1(n11775), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11722) );
  NAND2_X1 U14644 ( .A1(n11877), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11721) );
  NAND2_X1 U14645 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11720) );
  NAND2_X1 U14646 ( .A1(n11661), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11727) );
  NAND2_X1 U14647 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11726) );
  NAND2_X1 U14648 ( .A1(n11662), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11725) );
  NAND2_X1 U14649 ( .A1(n12379), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11724) );
  NAND4_X4 U14650 ( .A1(n11731), .A2(n11730), .A3(n11729), .A4(n11728), .ZN(
        n19858) );
  AND2_X4 U14651 ( .A1(n9618), .A2(n19858), .ZN(n13838) );
  NAND2_X1 U14652 ( .A1(n12503), .A2(n12465), .ZN(n11735) );
  INV_X1 U14653 ( .A(n12962), .ZN(n11736) );
  NOR2_X1 U14654 ( .A1(n11690), .A2(n13007), .ZN(n12895) );
  NAND2_X1 U14655 ( .A1(n9630), .A2(n19858), .ZN(n13341) );
  NAND2_X1 U14656 ( .A1(n19863), .A2(n9618), .ZN(n11757) );
  AND2_X1 U14657 ( .A1(n13341), .A2(n11757), .ZN(n11743) );
  INV_X1 U14658 ( .A(n11739), .ZN(n11742) );
  NAND2_X1 U14659 ( .A1(n11759), .A2(n19844), .ZN(n11741) );
  NAND4_X1 U14660 ( .A1(n11753), .A2(n11743), .A3(n11742), .A4(n11741), .ZN(
        n11744) );
  NAND2_X1 U14661 ( .A1(n12443), .A2(n11733), .ZN(n11745) );
  NAND2_X1 U14662 ( .A1(n11824), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11749) );
  NAND2_X1 U14663 ( .A1(n20595), .A2(n15763), .ZN(n12595) );
  NAND2_X1 U14664 ( .A1(n20436), .A2(n20639), .ZN(n20286) );
  NAND2_X1 U14665 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20432) );
  NAND2_X1 U14666 ( .A1(n20286), .A2(n20432), .ZN(n20218) );
  OR2_X1 U14667 ( .A1(n15422), .A2(n20436), .ZN(n11818) );
  OAI21_X1 U14668 ( .B1(n12595), .B2(n20218), .A(n11818), .ZN(n11747) );
  INV_X1 U14669 ( .A(n11747), .ZN(n11748) );
  NAND2_X1 U14670 ( .A1(n11824), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11752) );
  MUX2_X1 U14671 ( .A(n15422), .B(n12595), .S(n20639), .Z(n11751) );
  INV_X1 U14672 ( .A(n11753), .ZN(n11755) );
  NAND2_X1 U14673 ( .A1(n12414), .A2(n11733), .ZN(n11754) );
  NAND2_X1 U14674 ( .A1(n11755), .A2(n11754), .ZN(n11766) );
  INV_X1 U14675 ( .A(n11756), .ZN(n13337) );
  INV_X1 U14676 ( .A(n11757), .ZN(n11758) );
  AOI21_X1 U14677 ( .B1(n11759), .B2(n13337), .A(n11758), .ZN(n12904) );
  NAND2_X1 U14678 ( .A1(n11739), .A2(n11760), .ZN(n13068) );
  AND4_X1 U14679 ( .A1(n13068), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n20595), 
        .A4(n13341), .ZN(n11765) );
  AND2_X1 U14680 ( .A1(n11756), .A2(n13007), .ZN(n12802) );
  INV_X1 U14681 ( .A(n11761), .ZN(n11762) );
  AND2_X1 U14682 ( .A1(n11733), .A2(n9618), .ZN(n13382) );
  AOI22_X1 U14683 ( .A1(n12802), .A2(n11763), .B1(n11762), .B2(n13382), .ZN(
        n11764) );
  NAND4_X1 U14684 ( .A1(n11766), .A2(n12904), .A3(n11765), .A4(n11764), .ZN(
        n11793) );
  INV_X1 U14685 ( .A(n11768), .ZN(n11767) );
  NAND2_X1 U14686 ( .A1(n19966), .A2(n11768), .ZN(n11823) );
  NAND2_X1 U14687 ( .A1(n19895), .A2(n11823), .ZN(n13343) );
  AOI22_X1 U14688 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11774) );
  INV_X1 U14689 ( .A(n11769), .ZN(n11770) );
  AOI22_X1 U14690 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U14691 ( .A1(n12356), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12221), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11772) );
  AOI22_X1 U14692 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11771) );
  NAND4_X1 U14693 ( .A1(n11774), .A2(n11773), .A3(n11772), .A4(n11771), .ZN(
        n11781) );
  AOI22_X1 U14694 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U14695 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11778) );
  AOI22_X1 U14696 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U14697 ( .A1(n12315), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11776) );
  NAND4_X1 U14698 ( .A1(n11779), .A2(n11778), .A3(n11777), .A4(n11776), .ZN(
        n11780) );
  NAND2_X1 U14699 ( .A1(n9708), .A2(n12501), .ZN(n11782) );
  AOI22_X1 U14700 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9632), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U14701 ( .A1(n11661), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U14702 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11784) );
  AOI22_X1 U14703 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11783) );
  NAND4_X1 U14704 ( .A1(n11786), .A2(n11785), .A3(n11784), .A4(n11783), .ZN(
        n11792) );
  AOI22_X1 U14705 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11790) );
  AOI22_X1 U14706 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11789) );
  AOI22_X1 U14707 ( .A1(n12356), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12221), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U14708 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11787) );
  NAND4_X1 U14709 ( .A1(n11790), .A2(n11789), .A3(n11788), .A4(n11787), .ZN(
        n11791) );
  NAND2_X1 U14710 ( .A1(n12466), .A2(n12562), .ZN(n12559) );
  INV_X1 U14711 ( .A(n12562), .ZN(n11811) );
  NAND2_X1 U14712 ( .A1(n12466), .A2(n11811), .ZN(n11806) );
  AOI22_X1 U14713 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U14714 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U14715 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U14716 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11796) );
  NAND4_X1 U14717 ( .A1(n11799), .A2(n11798), .A3(n11797), .A4(n11796), .ZN(
        n11805) );
  AOI22_X1 U14718 ( .A1(n12315), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11803) );
  AOI22_X1 U14719 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U14720 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12221), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U14721 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11800) );
  NAND4_X1 U14722 ( .A1(n11803), .A2(n11802), .A3(n11801), .A4(n11800), .ZN(
        n11804) );
  MUX2_X1 U14723 ( .A(n12559), .B(n11806), .S(n12500), .Z(n11807) );
  NOR2_X1 U14724 ( .A1(n11807), .A2(n15763), .ZN(n11855) );
  INV_X1 U14725 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11809) );
  AOI21_X1 U14726 ( .B1(n9630), .B2(n12500), .A(n15763), .ZN(n11808) );
  OAI211_X1 U14727 ( .C1(n12414), .C2(n11809), .A(n11808), .B(n12559), .ZN(
        n11856) );
  NAND2_X1 U14728 ( .A1(n19844), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11838) );
  INV_X1 U14729 ( .A(n11838), .ZN(n11810) );
  AOI22_X1 U14730 ( .A1(n9708), .A2(n11811), .B1(n11810), .B2(n12501), .ZN(
        n11813) );
  NAND2_X1 U14731 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11812) );
  INV_X1 U14732 ( .A(n11814), .ZN(n11815) );
  INV_X1 U14733 ( .A(n11818), .ZN(n11821) );
  INV_X1 U14734 ( .A(n11819), .ZN(n11820) );
  OAI21_X1 U14735 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11821), .A(
        n11820), .ZN(n11822) );
  NAND2_X1 U14736 ( .A1(n11824), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11826) );
  INV_X1 U14737 ( .A(n12595), .ZN(n11874) );
  XNOR2_X1 U14738 ( .A(n20432), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19853) );
  NAND2_X1 U14739 ( .A1(n11874), .A2(n19853), .ZN(n11825) );
  AOI22_X1 U14740 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U14741 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U14742 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U14743 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11828) );
  NAND4_X1 U14744 ( .A1(n11831), .A2(n11830), .A3(n11829), .A4(n11828), .ZN(
        n11837) );
  AOI22_X1 U14745 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11835) );
  AOI22_X1 U14746 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11834) );
  AOI22_X1 U14747 ( .A1(n12356), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12221), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U14748 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11832) );
  NAND4_X1 U14749 ( .A1(n11835), .A2(n11834), .A3(n11833), .A4(n11832), .ZN(
        n11836) );
  INV_X1 U14750 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11839) );
  OAI22_X1 U14751 ( .A1(n12448), .A2(n11839), .B1(n11838), .B2(n12496), .ZN(
        n11840) );
  INV_X1 U14752 ( .A(n11840), .ZN(n11841) );
  NAND2_X1 U14753 ( .A1(n11760), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12022) );
  INV_X2 U14754 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20437) );
  NOR2_X1 U14755 ( .A1(n11844), .A2(n20437), .ZN(n11862) );
  INV_X1 U14756 ( .A(n12196), .ZN(n12402) );
  INV_X1 U14757 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13345) );
  XNOR2_X1 U14758 ( .A(n13345), .B(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19714) );
  NAND2_X1 U14759 ( .A1(n20437), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13223) );
  OAI21_X1 U14760 ( .B1(n19714), .B2(n13331), .A(n13223), .ZN(n11845) );
  AOI21_X1 U14761 ( .B1(n12402), .B2(P1_EAX_REG_2__SCAN_IN), .A(n11845), .ZN(
        n11847) );
  INV_X1 U14762 ( .A(n13054), .ZN(n11846) );
  NAND2_X1 U14763 ( .A1(n12401), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11870) );
  INV_X1 U14764 ( .A(n13090), .ZN(n11869) );
  INV_X1 U14765 ( .A(n11848), .ZN(n11850) );
  NAND2_X1 U14766 ( .A1(n13224), .A2(n12093), .ZN(n11854) );
  AOI22_X1 U14767 ( .A1(n12402), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20437), .ZN(n11852) );
  NAND2_X1 U14768 ( .A1(n11861), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11851) );
  AND2_X1 U14769 ( .A1(n11852), .A2(n11851), .ZN(n11853) );
  NAND2_X1 U14770 ( .A1(n11854), .A2(n11853), .ZN(n12961) );
  INV_X1 U14771 ( .A(n11855), .ZN(n11857) );
  XNOR2_X1 U14772 ( .A(n11857), .B(n11856), .ZN(n11858) );
  NAND2_X1 U14773 ( .A1(n19925), .A2(n11760), .ZN(n11859) );
  NAND2_X1 U14774 ( .A1(n11859), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13117) );
  INV_X1 U14775 ( .A(n11861), .ZN(n11912) );
  NAND2_X1 U14776 ( .A1(n11862), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11864) );
  NAND2_X1 U14777 ( .A1(n20437), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11863) );
  OAI211_X1 U14778 ( .C1(n11912), .C2(n11607), .A(n11864), .B(n11863), .ZN(
        n11865) );
  AOI21_X1 U14779 ( .B1(n11860), .B2(n12093), .A(n11865), .ZN(n13116) );
  OR2_X1 U14780 ( .A1(n13117), .A2(n13116), .ZN(n13119) );
  INV_X1 U14781 ( .A(n13116), .ZN(n11866) );
  OR2_X1 U14782 ( .A1(n11866), .A2(n13331), .ZN(n11867) );
  NAND2_X1 U14783 ( .A1(n13119), .A2(n11867), .ZN(n12960) );
  NAND2_X1 U14784 ( .A1(n12961), .A2(n12960), .ZN(n13089) );
  NAND2_X1 U14785 ( .A1(n11869), .A2(n11868), .ZN(n13092) );
  NAND2_X1 U14786 ( .A1(n11824), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11876) );
  INV_X1 U14787 ( .A(n20432), .ZN(n19963) );
  NAND2_X1 U14788 ( .A1(n20217), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20074) );
  INV_X1 U14789 ( .A(n20074), .ZN(n11871) );
  NAND2_X1 U14790 ( .A1(n19963), .A2(n11871), .ZN(n20142) );
  OAI21_X1 U14791 ( .B1(n20432), .B2(n20148), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11872) );
  NAND2_X1 U14792 ( .A1(n20142), .A2(n11872), .ZN(n20151) );
  INV_X1 U14793 ( .A(n15422), .ZN(n11873) );
  AOI22_X1 U14794 ( .A1(n20151), .A2(n11874), .B1(n11873), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11875) );
  XNOR2_X2 U14795 ( .A(n13216), .B(n20003), .ZN(n13201) );
  AOI22_X1 U14796 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U14797 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U14798 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U14799 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11878) );
  NAND4_X1 U14800 ( .A1(n11881), .A2(n11880), .A3(n11879), .A4(n11878), .ZN(
        n11887) );
  AOI22_X1 U14801 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11885) );
  AOI22_X1 U14802 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U14803 ( .A1(n12356), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U14804 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11882) );
  NAND4_X1 U14805 ( .A1(n11885), .A2(n11884), .A3(n11883), .A4(n11882), .ZN(
        n11886) );
  AOI22_X1 U14806 ( .A1(n12443), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12454), .B2(n12519), .ZN(n11888) );
  NAND2_X1 U14807 ( .A1(n11890), .A2(n13228), .ZN(n11891) );
  NAND2_X1 U14808 ( .A1(n11922), .A2(n11891), .ZN(n19842) );
  OAI21_X1 U14809 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11892), .A(
        n11941), .ZN(n19702) );
  AOI22_X1 U14810 ( .A1(n12397), .A2(n19702), .B1(n12401), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11894) );
  NAND2_X1 U14811 ( .A1(n12402), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11893) );
  OAI211_X1 U14812 ( .C1(n11912), .C2(n11605), .A(n11894), .B(n11893), .ZN(
        n11895) );
  INV_X1 U14813 ( .A(n11895), .ZN(n11896) );
  NAND2_X1 U14814 ( .A1(n11897), .A2(n11896), .ZN(n13164) );
  NAND2_X1 U14815 ( .A1(n13165), .A2(n13164), .ZN(n13163) );
  INV_X1 U14816 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U14817 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11901) );
  AOI22_X1 U14818 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U14819 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U14820 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11898) );
  NAND4_X1 U14821 ( .A1(n11901), .A2(n11900), .A3(n11899), .A4(n11898), .ZN(
        n11907) );
  AOI22_X1 U14822 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U14823 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U14824 ( .A1(n12356), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11903) );
  AOI22_X1 U14825 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11902) );
  NAND4_X1 U14826 ( .A1(n11905), .A2(n11904), .A3(n11903), .A4(n11902), .ZN(
        n11906) );
  NAND2_X1 U14827 ( .A1(n12454), .A2(n12532), .ZN(n11908) );
  OAI21_X1 U14828 ( .B1(n12448), .B2(n11909), .A(n11908), .ZN(n11920) );
  INV_X1 U14829 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13217) );
  NAND2_X1 U14830 ( .A1(n20437), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11911) );
  NAND2_X1 U14831 ( .A1(n12402), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11910) );
  OAI211_X1 U14832 ( .C1(n11912), .C2(n13217), .A(n11911), .B(n11910), .ZN(
        n11913) );
  NAND2_X1 U14833 ( .A1(n11913), .A2(n13331), .ZN(n11916) );
  INV_X1 U14834 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11914) );
  XNOR2_X1 U14835 ( .A(n11941), .B(n11914), .ZN(n19694) );
  NAND2_X1 U14836 ( .A1(n19694), .A2(n12397), .ZN(n11915) );
  NAND2_X1 U14837 ( .A1(n11916), .A2(n11915), .ZN(n11917) );
  INV_X1 U14838 ( .A(n11920), .ZN(n11921) );
  INV_X1 U14839 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11934) );
  AOI22_X1 U14840 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U14841 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U14842 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U14843 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11923) );
  NAND4_X1 U14844 ( .A1(n11926), .A2(n11925), .A3(n11924), .A4(n11923), .ZN(
        n11932) );
  AOI22_X1 U14845 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U14846 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U14847 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11928) );
  AOI22_X1 U14848 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11927) );
  NAND4_X1 U14849 ( .A1(n11930), .A2(n11929), .A3(n11928), .A4(n11927), .ZN(
        n11931) );
  NAND2_X1 U14850 ( .A1(n12454), .A2(n12535), .ZN(n11933) );
  OAI21_X1 U14851 ( .B1(n12448), .B2(n11934), .A(n11933), .ZN(n11936) );
  INV_X1 U14852 ( .A(n11935), .ZN(n11937) );
  NAND2_X1 U14853 ( .A1(n11937), .A2(n9801), .ZN(n11938) );
  INV_X1 U14854 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11944) );
  INV_X1 U14855 ( .A(n11941), .ZN(n11939) );
  AOI21_X1 U14856 ( .B1(n11939), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11942) );
  NAND2_X1 U14857 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11940) );
  OR2_X1 U14858 ( .A1(n11942), .A2(n11958), .ZN(n19682) );
  AOI22_X1 U14859 ( .A1(n19682), .A2(n12397), .B1(n12401), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11943) );
  OAI21_X1 U14860 ( .B1(n12196), .B2(n11944), .A(n11943), .ZN(n11945) );
  INV_X1 U14861 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U14862 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U14863 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U14864 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U14865 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11946) );
  NAND4_X1 U14866 ( .A1(n11949), .A2(n11948), .A3(n11947), .A4(n11946), .ZN(
        n11955) );
  AOI22_X1 U14867 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U14868 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U14869 ( .A1(n12356), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11951) );
  AOI22_X1 U14870 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11950) );
  NAND4_X1 U14871 ( .A1(n11953), .A2(n11952), .A3(n11951), .A4(n11950), .ZN(
        n11954) );
  NAND2_X1 U14872 ( .A1(n12454), .A2(n12549), .ZN(n11956) );
  OAI21_X1 U14873 ( .B1(n12448), .B2(n11957), .A(n11956), .ZN(n11963) );
  XNOR2_X1 U14874 ( .A(n11964), .B(n11963), .ZN(n12542) );
  INV_X1 U14875 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11961) );
  OR2_X1 U14876 ( .A1(n11958), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11959) );
  NAND2_X1 U14877 ( .A1(n11968), .A2(n11959), .ZN(n19665) );
  AOI22_X1 U14878 ( .A1(n19665), .A2(n12397), .B1(n12401), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11960) );
  OAI21_X1 U14879 ( .B1(n12196), .B2(n11961), .A(n11960), .ZN(n11962) );
  INV_X1 U14880 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11966) );
  NAND2_X1 U14881 ( .A1(n12454), .A2(n12562), .ZN(n11965) );
  OAI21_X1 U14882 ( .B1(n11966), .B2(n12448), .A(n11965), .ZN(n11967) );
  NAND2_X1 U14883 ( .A1(n11968), .A2(n11971), .ZN(n11969) );
  NAND2_X1 U14884 ( .A1(n11989), .A2(n11969), .ZN(n15590) );
  NAND2_X1 U14885 ( .A1(n15590), .A2(n12397), .ZN(n11970) );
  OAI21_X1 U14886 ( .B1(n11971), .B2(n13223), .A(n11970), .ZN(n11972) );
  AOI21_X1 U14887 ( .B1(n12402), .B2(P1_EAX_REG_7__SCAN_IN), .A(n11972), .ZN(
        n11973) );
  AOI22_X1 U14888 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U14889 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U14890 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U14891 ( .A1(n9632), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11975) );
  NAND4_X1 U14892 ( .A1(n11978), .A2(n11977), .A3(n11976), .A4(n11975), .ZN(
        n11984) );
  AOI22_X1 U14893 ( .A1(n9611), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U14894 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11981) );
  AOI22_X1 U14895 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11980) );
  AOI22_X1 U14896 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11979) );
  NAND4_X1 U14897 ( .A1(n11982), .A2(n11981), .A3(n11980), .A4(n11979), .ZN(
        n11983) );
  OAI21_X1 U14898 ( .B1(n11984), .B2(n11983), .A(n12093), .ZN(n11988) );
  NAND2_X1 U14899 ( .A1(n12402), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11987) );
  XNOR2_X1 U14900 ( .A(n11989), .B(n13502), .ZN(n13540) );
  NAND2_X1 U14901 ( .A1(n13540), .A2(n12397), .ZN(n11986) );
  NAND2_X1 U14902 ( .A1(n12401), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11985) );
  XNOR2_X1 U14903 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n12019), .ZN(
        n19657) );
  INV_X1 U14904 ( .A(n19657), .ZN(n12006) );
  AOI22_X1 U14905 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11994) );
  AOI22_X1 U14906 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U14907 ( .A1(n12242), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U14908 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11991) );
  NAND4_X1 U14909 ( .A1(n11994), .A2(n11993), .A3(n11992), .A4(n11991), .ZN(
        n12001) );
  AOI22_X1 U14910 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9612), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U14911 ( .A1(n11995), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U14912 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U14913 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11996) );
  NAND4_X1 U14914 ( .A1(n11999), .A2(n11998), .A3(n11997), .A4(n11996), .ZN(
        n12000) );
  OAI21_X1 U14915 ( .B1(n12001), .B2(n12000), .A(n12093), .ZN(n12004) );
  NAND2_X1 U14916 ( .A1(n12402), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12003) );
  NAND2_X1 U14917 ( .A1(n12401), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12002) );
  NAND3_X1 U14918 ( .A1(n12004), .A2(n12003), .A3(n12002), .ZN(n12005) );
  AOI21_X1 U14919 ( .B1(n12006), .B2(n12397), .A(n12005), .ZN(n13544) );
  AOI22_X1 U14920 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(n9612), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12011) );
  AOI22_X1 U14921 ( .A1(n12315), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U14922 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12009) );
  AOI22_X1 U14923 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12008) );
  NAND4_X1 U14924 ( .A1(n12011), .A2(n12010), .A3(n12009), .A4(n12008), .ZN(
        n12017) );
  AOI22_X1 U14925 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U14926 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U14927 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U14928 ( .A1(n12242), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12012) );
  NAND4_X1 U14929 ( .A1(n12015), .A2(n12014), .A3(n12013), .A4(n12012), .ZN(
        n12016) );
  NOR2_X1 U14930 ( .A1(n12017), .A2(n12016), .ZN(n12023) );
  XNOR2_X1 U14931 ( .A(n12024), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14345) );
  NAND2_X1 U14932 ( .A1(n14345), .A2(n12397), .ZN(n12021) );
  AOI22_X1 U14933 ( .A1(n12402), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12401), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12020) );
  OAI211_X1 U14934 ( .C1(n12023), .C2(n12022), .A(n12021), .B(n12020), .ZN(
        n13565) );
  INV_X1 U14935 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n13631) );
  OR2_X1 U14936 ( .A1(n12196), .A2(n13631), .ZN(n12027) );
  OAI21_X1 U14937 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12025), .A(
        n12053), .ZN(n15582) );
  AOI22_X1 U14938 ( .A1(n12397), .A2(n15582), .B1(n12401), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12026) );
  NAND2_X1 U14939 ( .A1(n12027), .A2(n12026), .ZN(n13620) );
  AOI22_X1 U14940 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U14941 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12030) );
  AOI22_X1 U14942 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U14943 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12028) );
  NAND4_X1 U14944 ( .A1(n12031), .A2(n12030), .A3(n12029), .A4(n12028), .ZN(
        n12037) );
  AOI22_X1 U14945 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9612), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12035) );
  AOI22_X1 U14946 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U14947 ( .A1(n12315), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12033) );
  AOI22_X1 U14948 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12032) );
  NAND4_X1 U14949 ( .A1(n12035), .A2(n12034), .A3(n12033), .A4(n12032), .ZN(
        n12036) );
  OR2_X1 U14950 ( .A1(n12037), .A2(n12036), .ZN(n12038) );
  AND2_X1 U14951 ( .A1(n12093), .A2(n12038), .ZN(n14064) );
  INV_X1 U14952 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12039) );
  XNOR2_X1 U14953 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12069), .ZN(
        n14332) );
  AOI22_X1 U14954 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12043) );
  AOI22_X1 U14955 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U14956 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U14957 ( .A1(n12315), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12040) );
  NAND4_X1 U14958 ( .A1(n12043), .A2(n12042), .A3(n12041), .A4(n12040), .ZN(
        n12049) );
  AOI22_X1 U14959 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12047) );
  AOI22_X1 U14960 ( .A1(n12309), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U14961 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U14962 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12044) );
  NAND4_X1 U14963 ( .A1(n12047), .A2(n12046), .A3(n12045), .A4(n12044), .ZN(
        n12048) );
  OR2_X1 U14964 ( .A1(n12049), .A2(n12048), .ZN(n12050) );
  AOI22_X1 U14965 ( .A1(n12093), .A2(n12050), .B1(n12401), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12052) );
  NAND2_X1 U14966 ( .A1(n11862), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12051) );
  OAI211_X1 U14967 ( .C1(n14332), .C2(n13331), .A(n12052), .B(n12051), .ZN(
        n14068) );
  INV_X1 U14968 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14211) );
  XNOR2_X1 U14969 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12053), .ZN(
        n15573) );
  INV_X1 U14970 ( .A(n15573), .ZN(n12054) );
  AOI22_X1 U14971 ( .A1(n12401), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12397), .B2(n12054), .ZN(n12067) );
  AOI22_X1 U14972 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9632), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U14973 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U14974 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12056) );
  AOI22_X1 U14975 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12055) );
  NAND4_X1 U14976 ( .A1(n12058), .A2(n12057), .A3(n12056), .A4(n12055), .ZN(
        n12064) );
  AOI22_X1 U14977 ( .A1(n12242), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9611), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U14978 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U14979 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U14980 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12059) );
  NAND4_X1 U14981 ( .A1(n12062), .A2(n12061), .A3(n12060), .A4(n12059), .ZN(
        n12063) );
  OR2_X1 U14982 ( .A1(n12064), .A2(n12063), .ZN(n12065) );
  NAND2_X1 U14983 ( .A1(n12093), .A2(n12065), .ZN(n12066) );
  OAI211_X1 U14984 ( .C1(n12196), .C2(n14211), .A(n12067), .B(n12066), .ZN(
        n14140) );
  AND2_X1 U14985 ( .A1(n14068), .A2(n14140), .ZN(n12068) );
  INV_X1 U14986 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14078) );
  XNOR2_X1 U14987 ( .A(n12084), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14320) );
  AOI22_X1 U14988 ( .A1(n12242), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9612), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12073) );
  AOI22_X1 U14989 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9632), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U14990 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12384), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U14991 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11668), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12070) );
  NAND4_X1 U14992 ( .A1(n12073), .A2(n12072), .A3(n12071), .A4(n12070), .ZN(
        n12079) );
  AOI22_X1 U14993 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12077) );
  AOI22_X1 U14994 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12076) );
  AOI22_X1 U14995 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12075) );
  AOI22_X1 U14996 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12074) );
  NAND4_X1 U14997 ( .A1(n12077), .A2(n12076), .A3(n12075), .A4(n12074), .ZN(
        n12078) );
  OAI21_X1 U14998 ( .B1(n12079), .B2(n12078), .A(n12093), .ZN(n12082) );
  NAND2_X1 U14999 ( .A1(n11862), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12081) );
  NAND2_X1 U15000 ( .A1(n12401), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12080) );
  NAND3_X1 U15001 ( .A1(n12082), .A2(n12081), .A3(n12080), .ZN(n12083) );
  AOI21_X1 U15002 ( .B1(n14320), .B2(n12397), .A(n12083), .ZN(n13641) );
  XOR2_X1 U15003 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n12102), .Z(
        n15563) );
  INV_X1 U15004 ( .A(n15563), .ZN(n12100) );
  AOI22_X1 U15005 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9631), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12088) );
  AOI22_X1 U15006 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12087) );
  AOI22_X1 U15007 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U15008 ( .A1(n9632), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12085) );
  NAND4_X1 U15009 ( .A1(n12088), .A2(n12087), .A3(n12086), .A4(n12085), .ZN(
        n12095) );
  AOI22_X1 U15010 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15011 ( .A1(n12242), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11668), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U15012 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12090) );
  AOI22_X1 U15013 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12089) );
  NAND4_X1 U15014 ( .A1(n12092), .A2(n12091), .A3(n12090), .A4(n12089), .ZN(
        n12094) );
  OAI21_X1 U15015 ( .B1(n12095), .B2(n12094), .A(n12093), .ZN(n12098) );
  NAND2_X1 U15016 ( .A1(n11862), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12097) );
  NAND2_X1 U15017 ( .A1(n12401), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12096) );
  NAND3_X1 U15018 ( .A1(n12098), .A2(n12097), .A3(n12096), .ZN(n12099) );
  AOI21_X1 U15019 ( .B1(n12100), .B2(n12397), .A(n12099), .ZN(n14052) );
  XNOR2_X1 U15020 ( .A(n12119), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14309) );
  NAND2_X1 U15021 ( .A1(n14309), .A2(n12397), .ZN(n12117) );
  INV_X1 U15022 ( .A(n15391), .ZN(n13188) );
  AOI22_X1 U15023 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U15024 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9611), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U15025 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U15026 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12103) );
  NAND4_X1 U15027 ( .A1(n12106), .A2(n12105), .A3(n12104), .A4(n12103), .ZN(
        n12112) );
  AOI22_X1 U15028 ( .A1(n9632), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12110) );
  AOI22_X1 U15029 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11668), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15030 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15031 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12107) );
  NAND4_X1 U15032 ( .A1(n12110), .A2(n12109), .A3(n12108), .A4(n12107), .ZN(
        n12111) );
  NOR2_X1 U15033 ( .A1(n12112), .A2(n12111), .ZN(n12115) );
  INV_X1 U15034 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12118) );
  AOI21_X1 U15035 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n12118), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12113) );
  AOI21_X1 U15036 ( .B1(n12402), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12113), .ZN(
        n12114) );
  OAI21_X1 U15037 ( .B1(n12368), .B2(n12115), .A(n12114), .ZN(n12116) );
  NAND2_X1 U15038 ( .A1(n12117), .A2(n12116), .ZN(n14039) );
  XNOR2_X1 U15039 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12132), .ZN(
        n15555) );
  AOI22_X1 U15040 ( .A1(n11862), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n12401), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U15041 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15042 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(n9621), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15043 ( .A1(n11661), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15044 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11668), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12120) );
  NAND4_X1 U15045 ( .A1(n12123), .A2(n12122), .A3(n12121), .A4(n12120), .ZN(
        n12129) );
  AOI22_X1 U15046 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15047 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12126) );
  AOI22_X1 U15048 ( .A1(n12315), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12125) );
  AOI22_X1 U15049 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12124) );
  NAND4_X1 U15050 ( .A1(n12127), .A2(n12126), .A3(n12125), .A4(n12124), .ZN(
        n12128) );
  INV_X1 U15051 ( .A(n12368), .ZN(n12394) );
  OAI21_X1 U15052 ( .B1(n12129), .B2(n12128), .A(n12394), .ZN(n12130) );
  OAI211_X1 U15053 ( .C1(n15555), .C2(n13331), .A(n12131), .B(n12130), .ZN(
        n14025) );
  INV_X1 U15054 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14030) );
  XNOR2_X1 U15055 ( .A(n12163), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15502) );
  NAND2_X1 U15056 ( .A1(n15502), .A2(n12397), .ZN(n12147) );
  AOI22_X1 U15057 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U15058 ( .A1(n12315), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U15059 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U15060 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12133) );
  NAND4_X1 U15061 ( .A1(n12136), .A2(n12135), .A3(n12134), .A4(n12133), .ZN(
        n12142) );
  AOI22_X1 U15062 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12140) );
  AOI22_X1 U15063 ( .A1(n12309), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U15064 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11668), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U15065 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12137) );
  NAND4_X1 U15066 ( .A1(n12140), .A2(n12139), .A3(n12138), .A4(n12137), .ZN(
        n12141) );
  NOR2_X1 U15067 ( .A1(n12142), .A2(n12141), .ZN(n12144) );
  AOI22_X1 U15068 ( .A1(n11862), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20437), .ZN(n12143) );
  OAI21_X1 U15069 ( .B1(n12368), .B2(n12144), .A(n12143), .ZN(n12145) );
  NAND2_X1 U15070 ( .A1(n12145), .A2(n13331), .ZN(n12146) );
  NAND2_X1 U15071 ( .A1(n12147), .A2(n12146), .ZN(n14122) );
  AOI22_X1 U15072 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9611), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15073 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U15074 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U15075 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12149) );
  NAND4_X1 U15076 ( .A1(n12152), .A2(n12151), .A3(n12150), .A4(n12149), .ZN(
        n12158) );
  AOI22_X1 U15077 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9632), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U15078 ( .A1(n11661), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12155) );
  AOI22_X1 U15079 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U15080 ( .A1(n12242), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11668), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12153) );
  NAND4_X1 U15081 ( .A1(n12156), .A2(n12155), .A3(n12154), .A4(n12153), .ZN(
        n12157) );
  NOR2_X1 U15082 ( .A1(n12158), .A2(n12157), .ZN(n12162) );
  OAI21_X1 U15083 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20334), .A(
        n20437), .ZN(n12159) );
  INV_X1 U15084 ( .A(n12159), .ZN(n12160) );
  AOI21_X1 U15085 ( .B1(n11862), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12160), .ZN(
        n12161) );
  OAI21_X1 U15086 ( .B1(n12368), .B2(n12162), .A(n12161), .ZN(n12166) );
  OAI21_X1 U15087 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n12164), .A(
        n12182), .ZN(n15549) );
  OR2_X1 U15088 ( .A1(n13331), .A2(n15549), .ZN(n12165) );
  AOI22_X1 U15089 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12314), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U15090 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15091 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15092 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12167) );
  NAND4_X1 U15093 ( .A1(n12170), .A2(n12169), .A3(n12168), .A4(n12167), .ZN(
        n12176) );
  AOI22_X1 U15094 ( .A1(n12242), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9611), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12174) );
  AOI22_X1 U15095 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12173) );
  AOI22_X1 U15096 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11668), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15097 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12171) );
  NAND4_X1 U15098 ( .A1(n12174), .A2(n12173), .A3(n12172), .A4(n12171), .ZN(
        n12175) );
  NOR2_X1 U15099 ( .A1(n12176), .A2(n12175), .ZN(n12179) );
  INV_X1 U15100 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15499) );
  AOI21_X1 U15101 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15499), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12177) );
  AOI21_X1 U15102 ( .B1(n11862), .B2(P1_EAX_REG_20__SCAN_IN), .A(n12177), .ZN(
        n12178) );
  OAI21_X1 U15103 ( .B1(n12368), .B2(n12179), .A(n12178), .ZN(n12181) );
  XNOR2_X1 U15104 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n12182), .ZN(
        n15489) );
  NAND2_X1 U15105 ( .A1(n12397), .A2(n15489), .ZN(n12180) );
  NAND2_X1 U15106 ( .A1(n12181), .A2(n12180), .ZN(n14115) );
  OR2_X1 U15107 ( .A1(n12183), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12184) );
  NAND2_X1 U15108 ( .A1(n12184), .A2(n12275), .ZN(n15481) );
  INV_X1 U15109 ( .A(n15481), .ZN(n15537) );
  AOI22_X1 U15110 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U15111 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9612), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U15112 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11661), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15113 ( .A1(n9632), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12185) );
  NAND4_X1 U15114 ( .A1(n12188), .A2(n12187), .A3(n12186), .A4(n12185), .ZN(
        n12194) );
  AOI22_X1 U15115 ( .A1(n12309), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U15116 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15117 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11668), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15118 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12189) );
  NAND4_X1 U15119 ( .A1(n12192), .A2(n12191), .A3(n12190), .A4(n12189), .ZN(
        n12193) );
  OR2_X1 U15120 ( .A1(n12194), .A2(n12193), .ZN(n12198) );
  INV_X1 U15121 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14175) );
  NAND2_X1 U15122 ( .A1(n20437), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12195) );
  OAI211_X1 U15123 ( .C1(n12196), .C2(n14175), .A(n13331), .B(n12195), .ZN(
        n12197) );
  AOI21_X1 U15124 ( .B1(n12394), .B2(n12198), .A(n12197), .ZN(n12199) );
  AOI21_X1 U15125 ( .B1(n15537), .B2(n12397), .A(n12199), .ZN(n14111) );
  AOI22_X1 U15126 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U15127 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9632), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15128 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12309), .B1(
        n11661), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12202) );
  AOI22_X1 U15129 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12201) );
  NAND4_X1 U15130 ( .A1(n12204), .A2(n12203), .A3(n12202), .A4(n12201), .ZN(
        n12210) );
  AOI22_X1 U15131 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15132 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15133 ( .A1(n9611), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15134 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n9621), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12205) );
  NAND4_X1 U15135 ( .A1(n12208), .A2(n12207), .A3(n12206), .A4(n12205), .ZN(
        n12209) );
  NOR2_X1 U15136 ( .A1(n12210), .A2(n12209), .ZN(n12214) );
  NAND2_X1 U15137 ( .A1(n20437), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12211) );
  NAND2_X1 U15138 ( .A1(n13331), .A2(n12211), .ZN(n12212) );
  AOI21_X1 U15139 ( .B1(n12402), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12212), .ZN(
        n12213) );
  OAI21_X1 U15140 ( .B1(n12368), .B2(n12214), .A(n12213), .ZN(n12216) );
  XNOR2_X1 U15141 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n12275), .ZN(
        n15476) );
  NAND2_X1 U15142 ( .A1(n15476), .A2(n12397), .ZN(n12215) );
  AOI22_X1 U15143 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9612), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15144 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9632), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12219) );
  AOI22_X1 U15145 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15146 ( .A1(n11662), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12217) );
  NAND4_X1 U15147 ( .A1(n12220), .A2(n12219), .A3(n12218), .A4(n12217), .ZN(
        n12227) );
  AOI22_X1 U15148 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U15149 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15150 ( .A1(n12242), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12223) );
  AOI22_X1 U15151 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12222) );
  NAND4_X1 U15152 ( .A1(n12225), .A2(n12224), .A3(n12223), .A4(n12222), .ZN(
        n12226) );
  NOR2_X1 U15153 ( .A1(n12227), .A2(n12226), .ZN(n12280) );
  AOI22_X1 U15154 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U15155 ( .A1(n12242), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U15156 ( .A1(n12356), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U15157 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12228) );
  NAND4_X1 U15158 ( .A1(n12231), .A2(n12230), .A3(n12229), .A4(n12228), .ZN(
        n12237) );
  AOI22_X1 U15159 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9631), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U15160 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U15161 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12233) );
  AOI22_X1 U15162 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12232) );
  NAND4_X1 U15163 ( .A1(n12235), .A2(n12234), .A3(n12233), .A4(n12232), .ZN(
        n12236) );
  NOR2_X1 U15164 ( .A1(n12237), .A2(n12236), .ZN(n12299) );
  AOI22_X1 U15165 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U15166 ( .A1(n12315), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12240) );
  AOI22_X1 U15167 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U15168 ( .A1(n11662), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12238) );
  NAND4_X1 U15169 ( .A1(n12241), .A2(n12240), .A3(n12239), .A4(n12238), .ZN(
        n12249) );
  AOI22_X1 U15170 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15171 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15172 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U15173 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12244) );
  NAND4_X1 U15174 ( .A1(n12247), .A2(n12246), .A3(n12245), .A4(n12244), .ZN(
        n12248) );
  NOR2_X1 U15175 ( .A1(n12249), .A2(n12248), .ZN(n12298) );
  NOR2_X1 U15176 ( .A1(n12299), .A2(n12298), .ZN(n12291) );
  AOI22_X1 U15177 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15178 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15179 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U15180 ( .A1(n11662), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12250) );
  NAND4_X1 U15181 ( .A1(n12253), .A2(n12252), .A3(n12251), .A4(n12250), .ZN(
        n12260) );
  AOI22_X1 U15182 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12258) );
  AOI22_X1 U15183 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12257) );
  AOI22_X1 U15184 ( .A1(n12356), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12256) );
  AOI22_X1 U15185 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12255) );
  NAND4_X1 U15186 ( .A1(n12258), .A2(n12257), .A3(n12256), .A4(n12255), .ZN(
        n12259) );
  OR2_X1 U15187 ( .A1(n12260), .A2(n12259), .ZN(n12290) );
  NAND2_X1 U15188 ( .A1(n12291), .A2(n12290), .ZN(n12281) );
  NOR2_X1 U15189 ( .A1(n12280), .A2(n12281), .ZN(n12323) );
  AOI22_X1 U15190 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12264) );
  AOI22_X1 U15191 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U15192 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12262) );
  AOI22_X1 U15193 ( .A1(n11662), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12261) );
  NAND4_X1 U15194 ( .A1(n12264), .A2(n12263), .A3(n12262), .A4(n12261), .ZN(
        n12270) );
  AOI22_X1 U15195 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15196 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U15197 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U15198 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12265) );
  NAND4_X1 U15199 ( .A1(n12268), .A2(n12267), .A3(n12266), .A4(n12265), .ZN(
        n12269) );
  OR2_X1 U15200 ( .A1(n12270), .A2(n12269), .ZN(n12322) );
  INV_X1 U15201 ( .A(n12322), .ZN(n12271) );
  XNOR2_X1 U15202 ( .A(n12323), .B(n12271), .ZN(n12272) );
  NAND2_X1 U15203 ( .A1(n12272), .A2(n12394), .ZN(n12279) );
  NAND2_X1 U15204 ( .A1(n20437), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12273) );
  NAND2_X1 U15205 ( .A1(n13331), .A2(n12273), .ZN(n12274) );
  AOI21_X1 U15206 ( .B1(n12402), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12274), .ZN(
        n12278) );
  INV_X1 U15207 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15471) );
  XNOR2_X1 U15208 ( .A(n12328), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14247) );
  AND2_X1 U15209 ( .A1(n14247), .A2(n12397), .ZN(n12277) );
  AOI21_X1 U15210 ( .B1(n12279), .B2(n12278), .A(n12277), .ZN(n13970) );
  XNOR2_X1 U15211 ( .A(n12281), .B(n12280), .ZN(n12284) );
  INV_X1 U15212 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14254) );
  AOI21_X1 U15213 ( .B1(n14254), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12282) );
  AOI21_X1 U15214 ( .B1(n12402), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12282), .ZN(
        n12283) );
  OAI21_X1 U15215 ( .B1(n12284), .B2(n12368), .A(n12283), .ZN(n12289) );
  INV_X1 U15216 ( .A(n12285), .ZN(n12286) );
  NAND2_X1 U15217 ( .A1(n12286), .A2(n14254), .ZN(n12287) );
  AND2_X1 U15218 ( .A1(n12328), .A2(n12287), .ZN(n14256) );
  NAND2_X1 U15219 ( .A1(n14256), .A2(n12397), .ZN(n12288) );
  NAND2_X1 U15220 ( .A1(n12289), .A2(n12288), .ZN(n13983) );
  XNOR2_X1 U15221 ( .A(n12291), .B(n12290), .ZN(n12295) );
  NAND2_X1 U15222 ( .A1(n20437), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12292) );
  NAND2_X1 U15223 ( .A1(n13331), .A2(n12292), .ZN(n12293) );
  AOI21_X1 U15224 ( .B1(n11862), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12293), .ZN(
        n12294) );
  OAI21_X1 U15225 ( .B1(n12295), .B2(n12368), .A(n12294), .ZN(n12297) );
  XNOR2_X1 U15226 ( .A(n12304), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14269) );
  NAND2_X1 U15227 ( .A1(n14269), .A2(n12397), .ZN(n12296) );
  NAND2_X1 U15228 ( .A1(n12297), .A2(n12296), .ZN(n14000) );
  XNOR2_X1 U15229 ( .A(n12299), .B(n12298), .ZN(n12303) );
  NAND2_X1 U15230 ( .A1(n20437), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12300) );
  NAND2_X1 U15231 ( .A1(n13331), .A2(n12300), .ZN(n12301) );
  AOI21_X1 U15232 ( .B1(n11862), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12301), .ZN(
        n12302) );
  OAI21_X1 U15233 ( .B1(n12368), .B2(n12303), .A(n12302), .ZN(n12307) );
  OAI21_X1 U15234 ( .B1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n12305), .A(
        n12304), .ZN(n15534) );
  OR2_X1 U15235 ( .A1(n15534), .A2(n13331), .ZN(n12306) );
  NAND2_X1 U15236 ( .A1(n12307), .A2(n12306), .ZN(n14096) );
  NOR2_X1 U15237 ( .A1(n13983), .A2(n13981), .ZN(n13968) );
  AND2_X1 U15238 ( .A1(n13970), .A2(n13968), .ZN(n12308) );
  AOI22_X1 U15239 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U15240 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15241 ( .A1(n11795), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U15242 ( .A1(n11662), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12310) );
  NAND4_X1 U15243 ( .A1(n12313), .A2(n12312), .A3(n12311), .A4(n12310), .ZN(
        n12321) );
  AOI22_X1 U15244 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12356), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12319) );
  AOI22_X1 U15245 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12318) );
  AOI22_X1 U15246 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U15247 ( .A1(n9632), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12316) );
  NAND4_X1 U15248 ( .A1(n12319), .A2(n12318), .A3(n12317), .A4(n12316), .ZN(
        n12320) );
  NOR2_X1 U15249 ( .A1(n12321), .A2(n12320), .ZN(n12335) );
  NAND2_X1 U15250 ( .A1(n12323), .A2(n12322), .ZN(n12334) );
  XNOR2_X1 U15251 ( .A(n12335), .B(n12334), .ZN(n12327) );
  NAND2_X1 U15252 ( .A1(n20437), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12324) );
  NAND2_X1 U15253 ( .A1(n13331), .A2(n12324), .ZN(n12325) );
  AOI21_X1 U15254 ( .B1(n12402), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12325), .ZN(
        n12326) );
  OAI21_X1 U15255 ( .B1(n12327), .B2(n12368), .A(n12326), .ZN(n12333) );
  INV_X1 U15256 ( .A(n12328), .ZN(n12329) );
  NAND2_X1 U15257 ( .A1(n12329), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12330) );
  INV_X1 U15258 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13962) );
  NAND2_X1 U15259 ( .A1(n12330), .A2(n13962), .ZN(n12331) );
  NAND2_X1 U15260 ( .A1(n12370), .A2(n12331), .ZN(n14241) );
  NAND2_X1 U15261 ( .A1(n12333), .A2(n12332), .ZN(n13956) );
  NOR2_X1 U15262 ( .A1(n12335), .A2(n12334), .ZN(n12364) );
  AOI22_X1 U15263 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15264 ( .A1(n11661), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U15265 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U15266 ( .A1(n11662), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12336) );
  NAND4_X1 U15267 ( .A1(n12339), .A2(n12338), .A3(n12337), .A4(n12336), .ZN(
        n12345) );
  AOI22_X1 U15268 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12343) );
  AOI22_X1 U15269 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12342) );
  AOI22_X1 U15270 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12341) );
  AOI22_X1 U15271 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12340) );
  NAND4_X1 U15272 ( .A1(n12343), .A2(n12342), .A3(n12341), .A4(n12340), .ZN(
        n12344) );
  OR2_X1 U15273 ( .A1(n12345), .A2(n12344), .ZN(n12363) );
  XNOR2_X1 U15274 ( .A(n12364), .B(n12363), .ZN(n12349) );
  INV_X1 U15275 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12346) );
  AOI21_X1 U15276 ( .B1(n12346), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12347) );
  AOI21_X1 U15277 ( .B1(n12402), .B2(P1_EAX_REG_28__SCAN_IN), .A(n12347), .ZN(
        n12348) );
  OAI21_X1 U15278 ( .B1(n12349), .B2(n12368), .A(n12348), .ZN(n12351) );
  XNOR2_X1 U15279 ( .A(n12370), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14230) );
  NAND2_X1 U15280 ( .A1(n14230), .A2(n12397), .ZN(n12350) );
  NAND2_X1 U15281 ( .A1(n12351), .A2(n12350), .ZN(n13944) );
  AOI22_X1 U15282 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n12385), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12355) );
  AOI22_X1 U15283 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n12309), .B1(
        n9632), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12354) );
  AOI22_X1 U15284 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12353) );
  AOI22_X1 U15285 ( .A1(n11662), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12352) );
  NAND4_X1 U15286 ( .A1(n12355), .A2(n12354), .A3(n12353), .A4(n12352), .ZN(
        n12362) );
  AOI22_X1 U15287 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12148), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15288 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n12384), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15289 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12356), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U15290 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12357) );
  NAND4_X1 U15291 ( .A1(n12360), .A2(n12359), .A3(n12358), .A4(n12357), .ZN(
        n12361) );
  NOR2_X1 U15292 ( .A1(n12362), .A2(n12361), .ZN(n12377) );
  NAND2_X1 U15293 ( .A1(n12364), .A2(n12363), .ZN(n12376) );
  XNOR2_X1 U15294 ( .A(n12377), .B(n12376), .ZN(n12369) );
  NAND2_X1 U15295 ( .A1(n20437), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12365) );
  NAND2_X1 U15296 ( .A1(n13331), .A2(n12365), .ZN(n12366) );
  AOI21_X1 U15297 ( .B1(n12402), .B2(P1_EAX_REG_29__SCAN_IN), .A(n12366), .ZN(
        n12367) );
  OAI21_X1 U15298 ( .B1(n12369), .B2(n12368), .A(n12367), .ZN(n12375) );
  INV_X1 U15299 ( .A(n12370), .ZN(n12371) );
  NAND2_X1 U15300 ( .A1(n12371), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12372) );
  INV_X1 U15301 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12596) );
  NAND2_X1 U15302 ( .A1(n12372), .A2(n12596), .ZN(n12373) );
  NAND2_X1 U15303 ( .A1(n13934), .A2(n12397), .ZN(n12374) );
  NOR2_X1 U15304 ( .A1(n12377), .A2(n12376), .ZN(n12393) );
  AOI22_X1 U15305 ( .A1(n12309), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12383) );
  AOI22_X1 U15306 ( .A1(n9612), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12254), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12382) );
  AOI22_X1 U15307 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15308 ( .A1(n11662), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12379), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12380) );
  NAND4_X1 U15309 ( .A1(n12383), .A2(n12382), .A3(n12381), .A4(n12380), .ZN(
        n12391) );
  AOI22_X1 U15310 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12389) );
  AOI22_X1 U15311 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12388) );
  AOI22_X1 U15312 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12387) );
  AOI22_X1 U15313 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12386) );
  NAND4_X1 U15314 ( .A1(n12389), .A2(n12388), .A3(n12387), .A4(n12386), .ZN(
        n12390) );
  NOR2_X1 U15315 ( .A1(n12391), .A2(n12390), .ZN(n12392) );
  XNOR2_X1 U15316 ( .A(n12393), .B(n12392), .ZN(n12395) );
  NAND2_X1 U15317 ( .A1(n12395), .A2(n12394), .ZN(n12400) );
  INV_X1 U15318 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13863) );
  AOI21_X1 U15319 ( .B1(n13863), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12396) );
  AOI21_X1 U15320 ( .B1(n12402), .B2(P1_EAX_REG_30__SCAN_IN), .A(n12396), .ZN(
        n12399) );
  XNOR2_X1 U15321 ( .A(n13334), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13927) );
  AOI21_X1 U15322 ( .B1(n12400), .B2(n12399), .A(n12398), .ZN(n13860) );
  NAND2_X1 U15323 ( .A1(n13859), .A2(n13860), .ZN(n12405) );
  AOI22_X1 U15324 ( .A1(n12402), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12401), .ZN(n12403) );
  INV_X1 U15325 ( .A(n12403), .ZN(n12404) );
  XNOR2_X1 U15326 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12417) );
  NAND2_X1 U15327 ( .A1(n12420), .A2(n12417), .ZN(n12407) );
  NAND2_X1 U15328 ( .A1(n20436), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12406) );
  NAND2_X1 U15329 ( .A1(n12407), .A2(n12406), .ZN(n12433) );
  XNOR2_X1 U15330 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12432) );
  NAND2_X1 U15331 ( .A1(n12433), .A2(n12432), .ZN(n12409) );
  NAND2_X1 U15332 ( .A1(n20148), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12408) );
  NAND2_X1 U15333 ( .A1(n12409), .A2(n12408), .ZN(n12413) );
  MUX2_X1 U15334 ( .A(n20217), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12412) );
  NAND2_X1 U15335 ( .A1(n12413), .A2(n12412), .ZN(n12411) );
  NAND2_X1 U15336 ( .A1(n20217), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12410) );
  NAND2_X1 U15337 ( .A1(n12411), .A2(n12410), .ZN(n12451) );
  INV_X1 U15338 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19838) );
  OR2_X1 U15339 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19838), .ZN(
        n12452) );
  NOR2_X1 U15340 ( .A1(n12451), .A2(n12452), .ZN(n12471) );
  XNOR2_X1 U15341 ( .A(n12413), .B(n12412), .ZN(n12468) );
  INV_X1 U15342 ( .A(n12468), .ZN(n12442) );
  INV_X1 U15343 ( .A(n12414), .ZN(n12416) );
  AOI21_X1 U15344 ( .B1(n12416), .B2(n12415), .A(n15763), .ZN(n12418) );
  NAND2_X1 U15345 ( .A1(n11733), .A2(n12415), .ZN(n12423) );
  XNOR2_X1 U15346 ( .A(n12417), .B(n12420), .ZN(n12470) );
  AOI22_X1 U15347 ( .A1(n12418), .A2(n12423), .B1(n12443), .B2(n12470), .ZN(
        n12427) );
  INV_X1 U15348 ( .A(n12427), .ZN(n12431) );
  NOR2_X1 U15349 ( .A1(n12418), .A2(n11733), .ZN(n12444) );
  INV_X1 U15350 ( .A(n12470), .ZN(n12419) );
  NOR2_X1 U15351 ( .A1(n12444), .A2(n12419), .ZN(n12428) );
  INV_X1 U15352 ( .A(n12428), .ZN(n12430) );
  INV_X1 U15353 ( .A(n12420), .ZN(n12421) );
  OAI21_X1 U15354 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20639), .A(
        n12421), .ZN(n12424) );
  INV_X1 U15355 ( .A(n12424), .ZN(n12422) );
  NAND2_X1 U15356 ( .A1(n19858), .A2(n12415), .ZN(n12557) );
  AOI21_X1 U15357 ( .B1(n12454), .B2(n12422), .A(n12457), .ZN(n12426) );
  INV_X1 U15358 ( .A(n11690), .ZN(n12586) );
  NAND2_X1 U15359 ( .A1(n11756), .A2(n12423), .ZN(n12435) );
  AOI211_X1 U15360 ( .C1(n12586), .C2(n9618), .A(n12424), .B(n12435), .ZN(
        n12425) );
  AOI211_X1 U15361 ( .C1(n12428), .C2(n12427), .A(n12426), .B(n12425), .ZN(
        n12429) );
  AOI21_X1 U15362 ( .B1(n12431), .B2(n12430), .A(n12429), .ZN(n12440) );
  XNOR2_X1 U15363 ( .A(n12433), .B(n12432), .ZN(n12469) );
  INV_X1 U15364 ( .A(n12469), .ZN(n12434) );
  AOI211_X1 U15365 ( .C1(n12443), .C2(n12469), .A(n12435), .B(n12436), .ZN(
        n12439) );
  INV_X1 U15366 ( .A(n12435), .ZN(n12438) );
  INV_X1 U15367 ( .A(n12436), .ZN(n12437) );
  OAI22_X1 U15368 ( .A1(n12440), .A2(n12439), .B1(n12438), .B2(n12437), .ZN(
        n12441) );
  OAI21_X1 U15369 ( .B1(n12443), .B2(n12442), .A(n12441), .ZN(n12446) );
  AOI22_X1 U15370 ( .A1(n12444), .A2(n12471), .B1(n12457), .B2(n12468), .ZN(
        n12445) );
  NOR2_X1 U15371 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13217), .ZN(
        n12450) );
  NAND2_X1 U15372 ( .A1(n12473), .A2(n12454), .ZN(n12455) );
  NAND2_X1 U15373 ( .A1(n12457), .A2(n12473), .ZN(n12458) );
  INV_X1 U15374 ( .A(n12898), .ZN(n12461) );
  NAND2_X1 U15375 ( .A1(n15391), .A2(n9630), .ZN(n12460) );
  NAND2_X1 U15376 ( .A1(n12916), .A2(n13337), .ZN(n13192) );
  NAND2_X1 U15377 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n15448) );
  AND2_X1 U15378 ( .A1(n12462), .A2(n15448), .ZN(n13056) );
  NAND2_X1 U15379 ( .A1(n13056), .A2(n13838), .ZN(n12463) );
  AND2_X1 U15380 ( .A1(n13192), .A2(n12463), .ZN(n12464) );
  NAND3_X1 U15381 ( .A1(n12466), .A2(n14147), .A3(n12465), .ZN(n12996) );
  INV_X1 U15382 ( .A(n12467), .ZN(n12474) );
  NOR4_X1 U15383 ( .A1(n12471), .A2(n12470), .A3(n12469), .A4(n12468), .ZN(
        n12472) );
  NOR2_X1 U15384 ( .A1(n12473), .A2(n12472), .ZN(n12792) );
  AND2_X1 U15385 ( .A1(n12792), .A2(n15448), .ZN(n13047) );
  NAND2_X1 U15386 ( .A1(n12474), .A2(n13047), .ZN(n12919) );
  OAI21_X1 U15387 ( .B1(n12896), .B2(n12996), .A(n12919), .ZN(n12475) );
  NAND2_X1 U15388 ( .A1(n12475), .A2(n13052), .ZN(n12476) );
  NAND2_X1 U15389 ( .A1(n14221), .A2(n10112), .ZN(n12494) );
  NOR4_X1 U15390 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12481) );
  NOR4_X1 U15391 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12480) );
  NOR4_X1 U15392 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12479) );
  NOR4_X1 U15393 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12478) );
  AND4_X1 U15394 ( .A1(n12481), .A2(n12480), .A3(n12479), .A4(n12478), .ZN(
        n12486) );
  NOR4_X1 U15395 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12484) );
  NOR4_X1 U15396 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12483) );
  NOR4_X1 U15397 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12482) );
  INV_X1 U15398 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20520) );
  AND4_X1 U15399 ( .A1(n12484), .A2(n12483), .A3(n12482), .A4(n20520), .ZN(
        n12485) );
  NAND2_X1 U15400 ( .A1(n12486), .A2(n12485), .ZN(n12487) );
  NOR3_X1 U15401 ( .A1(n14206), .A2(n19839), .A3(n13054), .ZN(n12488) );
  AOI22_X1 U15402 ( .A1(n14198), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14206), .ZN(n12489) );
  INV_X1 U15403 ( .A(n12489), .ZN(n12492) );
  INV_X1 U15404 ( .A(n19839), .ZN(n19840) );
  NOR2_X1 U15405 ( .A1(n13054), .A2(n19840), .ZN(n12490) );
  NAND2_X1 U15406 ( .A1(n14210), .A2(n12490), .ZN(n14177) );
  INV_X1 U15407 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20776) );
  NOR2_X1 U15408 ( .A1(n14177), .A2(n20776), .ZN(n12491) );
  NAND2_X1 U15409 ( .A1(n12494), .A2(n12493), .ZN(P1_U2873) );
  NAND2_X1 U15410 ( .A1(n12500), .A2(n12501), .ZN(n12495) );
  NAND2_X1 U15411 ( .A1(n12495), .A2(n12496), .ZN(n12518) );
  OAI21_X1 U15412 ( .B1(n12496), .B2(n12495), .A(n12518), .ZN(n12497) );
  AND2_X1 U15413 ( .A1(n19868), .A2(n9630), .ZN(n12508) );
  AOI21_X1 U15414 ( .B1(n12497), .B2(n13382), .A(n12508), .ZN(n12498) );
  INV_X1 U15415 ( .A(n12500), .ZN(n12509) );
  XNOR2_X1 U15416 ( .A(n12509), .B(n12501), .ZN(n12502) );
  NAND2_X1 U15417 ( .A1(n12502), .A2(n13382), .ZN(n12506) );
  NOR2_X1 U15418 ( .A1(n12504), .A2(n12503), .ZN(n12505) );
  AND2_X1 U15419 ( .A1(n12506), .A2(n12505), .ZN(n12507) );
  AOI21_X1 U15420 ( .B1(n12509), .B2(n13382), .A(n12508), .ZN(n12510) );
  NAND2_X1 U15421 ( .A1(n19814), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12511) );
  INV_X1 U15422 ( .A(n12511), .ZN(n19815) );
  NAND2_X1 U15423 ( .A1(n12512), .A2(n19815), .ZN(n12513) );
  NAND2_X1 U15424 ( .A1(n12514), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12515) );
  NAND2_X1 U15425 ( .A1(n12516), .A2(n12515), .ZN(n12522) );
  INV_X1 U15426 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12517) );
  OR2_X1 U15427 ( .A1(n19842), .A2(n12557), .ZN(n12521) );
  NAND2_X1 U15428 ( .A1(n12518), .A2(n12519), .ZN(n12534) );
  OAI211_X1 U15429 ( .C1(n12519), .C2(n12518), .A(n12534), .B(n13382), .ZN(
        n12520) );
  NAND2_X1 U15430 ( .A1(n12521), .A2(n12520), .ZN(n13245) );
  NAND2_X1 U15431 ( .A1(n12522), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12523) );
  XNOR2_X1 U15432 ( .A(n12534), .B(n12532), .ZN(n12525) );
  NAND2_X1 U15433 ( .A1(n12525), .A2(n13382), .ZN(n12526) );
  INV_X1 U15434 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12527) );
  NAND2_X1 U15435 ( .A1(n12528), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12529) );
  NAND2_X1 U15436 ( .A1(n12530), .A2(n12529), .ZN(n15599) );
  NAND2_X1 U15437 ( .A1(n12531), .A2(n10104), .ZN(n12538) );
  INV_X1 U15438 ( .A(n12532), .ZN(n12533) );
  NOR2_X1 U15439 ( .A1(n12534), .A2(n12533), .ZN(n12536) );
  NAND2_X1 U15440 ( .A1(n12536), .A2(n12535), .ZN(n12548) );
  OAI211_X1 U15441 ( .C1(n12536), .C2(n12535), .A(n12548), .B(n13382), .ZN(
        n12537) );
  NAND2_X1 U15442 ( .A1(n12538), .A2(n12537), .ZN(n12539) );
  INV_X1 U15443 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15758) );
  XNOR2_X1 U15444 ( .A(n12539), .B(n15758), .ZN(n15598) );
  NAND2_X1 U15445 ( .A1(n15599), .A2(n15598), .ZN(n12541) );
  NAND2_X1 U15446 ( .A1(n12539), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12540) );
  NAND2_X1 U15447 ( .A1(n12542), .A2(n10104), .ZN(n12545) );
  XNOR2_X1 U15448 ( .A(n12548), .B(n12549), .ZN(n12543) );
  NAND2_X1 U15449 ( .A1(n12543), .A2(n13382), .ZN(n12544) );
  NAND2_X1 U15450 ( .A1(n12545), .A2(n12544), .ZN(n12546) );
  OR2_X1 U15451 ( .A1(n12546), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15592) );
  NAND2_X1 U15452 ( .A1(n12546), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15591) );
  NAND2_X1 U15453 ( .A1(n12547), .A2(n10104), .ZN(n12553) );
  INV_X1 U15454 ( .A(n12548), .ZN(n12550) );
  NAND2_X1 U15455 ( .A1(n12550), .A2(n12549), .ZN(n12564) );
  XNOR2_X1 U15456 ( .A(n12564), .B(n12562), .ZN(n12551) );
  NAND2_X1 U15457 ( .A1(n12551), .A2(n13382), .ZN(n12552) );
  NAND2_X1 U15458 ( .A1(n12553), .A2(n12552), .ZN(n12555) );
  XNOR2_X1 U15459 ( .A(n12555), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15583) );
  OR2_X1 U15460 ( .A1(n12555), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12556) );
  OR2_X1 U15461 ( .A1(n12557), .A2(n15763), .ZN(n12558) );
  NOR2_X1 U15462 ( .A1(n12559), .A2(n12558), .ZN(n12560) );
  NAND2_X1 U15463 ( .A1(n13382), .A2(n12562), .ZN(n12563) );
  OR2_X1 U15464 ( .A1(n12564), .A2(n12563), .ZN(n12565) );
  NAND2_X1 U15465 ( .A1(n15529), .A2(n12565), .ZN(n13536) );
  NAND2_X1 U15466 ( .A1(n13536), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12566) );
  INV_X1 U15467 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12568) );
  NAND2_X1 U15468 ( .A1(n15529), .A2(n12568), .ZN(n13585) );
  NAND2_X1 U15469 ( .A1(n15529), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12569) );
  NAND2_X1 U15470 ( .A1(n15551), .A2(n12569), .ZN(n14307) );
  INV_X1 U15471 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14428) );
  NAND2_X1 U15472 ( .A1(n15529), .A2(n14428), .ZN(n14304) );
  OAI21_X1 U15473 ( .B1(n14342), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n14305), .ZN(n12570) );
  INV_X1 U15474 ( .A(n12570), .ZN(n12571) );
  INV_X1 U15475 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12575) );
  NAND2_X1 U15476 ( .A1(n15529), .A2(n12575), .ZN(n12572) );
  INV_X1 U15477 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15681) );
  NAND2_X1 U15478 ( .A1(n15529), .A2(n15681), .ZN(n14329) );
  NAND2_X1 U15479 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12573) );
  NAND2_X1 U15480 ( .A1(n15529), .A2(n12573), .ZN(n14324) );
  NOR2_X1 U15481 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12574) );
  NOR2_X1 U15482 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12576) );
  INV_X1 U15483 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14437) );
  INV_X1 U15484 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15430) );
  INV_X1 U15485 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15638) );
  NOR2_X1 U15486 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12578) );
  NAND3_X1 U15487 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13849) );
  INV_X1 U15488 ( .A(n13849), .ZN(n12580) );
  INV_X1 U15489 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15606) );
  INV_X1 U15490 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14260) );
  INV_X1 U15491 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n20803) );
  NAND3_X1 U15492 ( .A1(n15606), .A2(n14260), .A3(n20803), .ZN(n14225) );
  INV_X1 U15493 ( .A(n14225), .ZN(n12582) );
  NAND2_X1 U15494 ( .A1(n12583), .A2(n14342), .ZN(n14249) );
  NAND3_X1 U15495 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14224) );
  AND2_X2 U15496 ( .A1(n14249), .A2(n14236), .ZN(n14237) );
  NAND2_X1 U15497 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14374) );
  NOR2_X2 U15498 ( .A1(n14237), .A2(n14374), .ZN(n13793) );
  NOR2_X1 U15499 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12585) );
  NOR2_X1 U15500 ( .A1(n15529), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13792) );
  AND2_X1 U15501 ( .A1(n15529), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14214) );
  AND2_X1 U15502 ( .A1(n12916), .A2(n12586), .ZN(n13062) );
  INV_X1 U15503 ( .A(n13859), .ZN(n12589) );
  NAND3_X1 U15504 ( .A1(n15763), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15765) );
  INV_X1 U15505 ( .A(n15765), .ZN(n12591) );
  NOR2_X1 U15506 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20288) );
  INV_X1 U15507 ( .A(n20442), .ZN(n20333) );
  NAND2_X1 U15508 ( .A1(n20442), .A2(n12595), .ZN(n20624) );
  AND2_X1 U15509 ( .A1(n20624), .A2(n15763), .ZN(n12592) );
  NAND2_X1 U15510 ( .A1(n20334), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12594) );
  NOR2_X1 U15511 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20437), .ZN(n20626) );
  INV_X1 U15512 ( .A(n20626), .ZN(n12593) );
  NAND2_X1 U15513 ( .A1(n12594), .A2(n12593), .ZN(n19812) );
  OR2_X1 U15514 ( .A1(n12595), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15731) );
  INV_X1 U15515 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20572) );
  NOR2_X1 U15516 ( .A1(n15731), .A2(n20572), .ZN(n14362) );
  NOR2_X1 U15517 ( .A1(n15603), .A2(n12596), .ZN(n12597) );
  AOI211_X1 U15518 ( .C1(n15600), .C2(n13934), .A(n14362), .B(n12597), .ZN(
        n12598) );
  NAND2_X1 U15519 ( .A1(n12601), .A2(n12600), .ZN(P1_U2970) );
  AND2_X1 U15520 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12602) );
  INV_X1 U15521 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14858) );
  NOR2_X2 U15522 ( .A1(n14695), .A2(n14858), .ZN(n14682) );
  INV_X1 U15523 ( .A(n14656), .ZN(n12605) );
  OR2_X1 U15524 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n14682), .ZN(
        n12604) );
  NOR2_X1 U15525 ( .A1(n9699), .A2(n12606), .ZN(n12607) );
  XNOR2_X1 U15526 ( .A(n12608), .B(n12607), .ZN(n13872) );
  AOI21_X1 U15527 ( .B1(n12609), .B2(n14973), .A(n15998), .ZN(n14838) );
  INV_X1 U15528 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12620) );
  INV_X1 U15529 ( .A(n12610), .ZN(n12660) );
  AND2_X1 U15530 ( .A1(n12660), .A2(n12611), .ZN(n12612) );
  NOR2_X1 U15531 ( .A1(n10127), .A2(n12612), .ZN(n15829) );
  NOR2_X1 U15532 ( .A1(n11181), .A2(n12613), .ZN(n13867) );
  AND2_X1 U15533 ( .A1(n12657), .A2(n12614), .ZN(n12615) );
  OR2_X1 U15534 ( .A1(n12615), .A2(n12672), .ZN(n15819) );
  NOR2_X1 U15535 ( .A1(n15819), .A2(n16055), .ZN(n12616) );
  AOI211_X1 U15536 ( .C1(n16057), .C2(n15829), .A(n13867), .B(n12616), .ZN(
        n12619) );
  INV_X1 U15537 ( .A(n16000), .ZN(n15978) );
  NOR2_X1 U15538 ( .A1(n14878), .A2(n12617), .ZN(n14859) );
  NOR2_X1 U15539 ( .A1(n14858), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12618) );
  NAND2_X1 U15540 ( .A1(n14859), .A2(n12618), .ZN(n14837) );
  OAI211_X1 U15541 ( .C1(n14838), .C2(n12620), .A(n12619), .B(n14837), .ZN(
        n12621) );
  AOI21_X1 U15542 ( .B1(n13872), .B2(n16063), .A(n12621), .ZN(n12622) );
  OAI21_X1 U15543 ( .B1(n13874), .B2(n16060), .A(n12622), .ZN(P2_U3024) );
  INV_X1 U15544 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20618) );
  NOR3_X1 U15545 ( .A1(P1_BE_N_REG_3__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20618), .ZN(n12624) );
  NOR4_X1 U15546 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_2__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12623) );
  NAND4_X1 U15547 ( .A1(n19839), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12624), .A4(
        n12623), .ZN(U214) );
  INV_X1 U15548 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19614) );
  NOR2_X1 U15549 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(n19614), .ZN(n12626) );
  NOR4_X1 U15550 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12625) );
  INV_X1 U15551 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20806) );
  NAND4_X1 U15552 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(n12626), .A3(n12625), .A4(
        n20806), .ZN(n12627) );
  NOR2_X1 U15553 ( .A1(n15033), .A2(n12627), .ZN(n16211) );
  NAND2_X1 U15554 ( .A1(n16211), .A2(U214), .ZN(U212) );
  NOR2_X1 U15555 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12627), .ZN(n16293)
         );
  NOR2_X1 U15556 ( .A1(n11057), .A2(n16010), .ZN(n12638) );
  OR2_X1 U15557 ( .A1(n12628), .A2(n12954), .ZN(n12629) );
  AND2_X1 U15558 ( .A1(n12629), .A2(n13041), .ZN(n13556) );
  INV_X1 U15559 ( .A(n13556), .ZN(n18788) );
  OAI22_X1 U15560 ( .A1(n16011), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n18788), .B2(n16055), .ZN(n12637) );
  XNOR2_X1 U15561 ( .A(n12631), .B(n12630), .ZN(n18790) );
  OAI22_X1 U15562 ( .A1(n16007), .A2(n16013), .B1(n16053), .B2(n18790), .ZN(
        n12636) );
  XNOR2_X1 U15563 ( .A(n12632), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13563) );
  XNOR2_X1 U15564 ( .A(n12633), .B(n12634), .ZN(n13560) );
  OAI22_X1 U15565 ( .A1(n13563), .A2(n16060), .B1(n16037), .B2(n13560), .ZN(
        n12635) );
  OR4_X1 U15566 ( .A1(n12638), .A2(n12637), .A3(n12636), .A4(n12635), .ZN(
        P2_U3040) );
  AOI211_X1 U15567 ( .C1(n14627), .C2(n12640), .A(n12639), .B(n18779), .ZN(
        n12651) );
  OAI22_X1 U15568 ( .A1(n20763), .A2(n18810), .B1(n12641), .B2(n18795), .ZN(
        n12650) );
  INV_X1 U15569 ( .A(n18819), .ZN(n18798) );
  INV_X1 U15570 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n20660) );
  OAI22_X1 U15571 ( .A1(n18798), .A2(n20660), .B1(n14629), .B2(n18694), .ZN(
        n12649) );
  AND2_X1 U15572 ( .A1(n14536), .A2(n12643), .ZN(n12644) );
  INV_X1 U15573 ( .A(n14789), .ZN(n12647) );
  AND2_X1 U15574 ( .A1(n14569), .A2(n12645), .ZN(n12646) );
  OR2_X1 U15575 ( .A1(n12646), .A2(n14467), .ZN(n14792) );
  OAI22_X1 U15576 ( .A1(n12647), .A2(n18789), .B1(n14792), .B2(n18812), .ZN(
        n12648) );
  OR4_X1 U15577 ( .A1(n12651), .A2(n12650), .A3(n12649), .A4(n12648), .ZN(
        P2_U2828) );
  AOI211_X1 U15578 ( .C1(n14685), .C2(n12653), .A(n12652), .B(n18779), .ZN(
        n12665) );
  OAI22_X1 U15579 ( .A1(n14683), .A2(n18694), .B1(n19553), .B2(n18810), .ZN(
        n12664) );
  OAI22_X1 U15580 ( .A1(n18798), .A2(n14555), .B1(n12654), .B2(n18795), .ZN(
        n12663) );
  NAND2_X1 U15581 ( .A1(n14498), .A2(n12655), .ZN(n12656) );
  NAND2_X1 U15582 ( .A1(n12657), .A2(n12656), .ZN(n14856) );
  NAND2_X1 U15583 ( .A1(n9703), .A2(n12658), .ZN(n12659) );
  AND2_X1 U15584 ( .A1(n12660), .A2(n12659), .ZN(n14853) );
  INV_X1 U15585 ( .A(n14853), .ZN(n12661) );
  OAI22_X1 U15586 ( .A1(n14856), .A2(n18789), .B1(n12661), .B2(n18812), .ZN(
        n12662) );
  OR4_X1 U15587 ( .A1(n12665), .A2(n12664), .A3(n12663), .A4(n12662), .ZN(
        P2_U2834) );
  AOI211_X1 U15588 ( .C1(n14661), .C2(n12667), .A(n18779), .B(n12666), .ZN(
        n12680) );
  INV_X1 U15589 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19556) );
  OAI22_X1 U15590 ( .A1(n14659), .A2(n18694), .B1(n19556), .B2(n18810), .ZN(
        n12679) );
  INV_X1 U15591 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12669) );
  OAI22_X1 U15592 ( .A1(n18798), .A2(n12669), .B1(n12668), .B2(n18795), .ZN(
        n12678) );
  NOR2_X1 U15593 ( .A1(n12672), .A2(n12671), .ZN(n12673) );
  OR2_X1 U15594 ( .A1(n12670), .A2(n12673), .ZN(n15816) );
  NOR2_X1 U15595 ( .A1(n10127), .A2(n12675), .ZN(n12676) );
  OR2_X1 U15596 ( .A1(n12674), .A2(n12676), .ZN(n14594) );
  OAI22_X1 U15597 ( .A1(n15816), .A2(n18789), .B1(n18812), .B2(n14594), .ZN(
        n12677) );
  OR4_X1 U15598 ( .A1(n12680), .A2(n12679), .A3(n12678), .A4(n12677), .ZN(
        P2_U2832) );
  NOR2_X1 U15599 ( .A1(n16087), .A2(n19494), .ZN(n12683) );
  INV_X1 U15600 ( .A(n12876), .ZN(n12867) );
  NAND2_X1 U15601 ( .A1(n12683), .A2(n12867), .ZN(n13459) );
  INV_X1 U15602 ( .A(n13459), .ZN(n18825) );
  INV_X1 U15603 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19626) );
  INV_X1 U15604 ( .A(n12681), .ZN(n12682) );
  NAND2_X1 U15605 ( .A1(n12683), .A2(n12682), .ZN(n12688) );
  OAI211_X1 U15606 ( .C1(n18825), .C2(n19626), .A(n18639), .B(n12688), .ZN(
        P2_U2814) );
  NOR2_X1 U15607 ( .A1(n18642), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n12685)
         );
  INV_X1 U15608 ( .A(n14452), .ZN(n12684) );
  AOI22_X1 U15609 ( .A1(n12685), .A2(n18639), .B1(n12684), .B2(n18642), .ZN(
        P2_U3612) );
  INV_X1 U15610 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n12816) );
  INV_X1 U15611 ( .A(n12688), .ZN(n12687) );
  OAI21_X1 U15612 ( .B1(n12874), .B2(n19504), .A(n12687), .ZN(n12705) );
  NAND2_X1 U15613 ( .A1(n12705), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12689) );
  OR3_X1 U15614 ( .A1(n12688), .A2(n12874), .A3(n19520), .ZN(n12741) );
  INV_X1 U15615 ( .A(n12741), .ZN(n12737) );
  MUX2_X1 U15616 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n15033), .Z(n18894) );
  NAND2_X1 U15617 ( .A1(n12737), .A2(n18894), .ZN(n12690) );
  OAI211_X1 U15618 ( .C1(n12816), .C2(n12811), .A(n12689), .B(n12690), .ZN(
        P2_U2962) );
  INV_X1 U15619 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n18910) );
  NAND2_X1 U15620 ( .A1(n12705), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12691) );
  OAI211_X1 U15621 ( .C1(n18910), .C2(n12811), .A(n12691), .B(n12690), .ZN(
        P2_U2977) );
  NAND2_X1 U15622 ( .A1(n12705), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12692) );
  NAND2_X1 U15623 ( .A1(n12737), .A2(n13440), .ZN(n12698) );
  OAI211_X1 U15624 ( .C1(n11599), .C2(n12811), .A(n12692), .B(n12698), .ZN(
        P2_U2966) );
  INV_X1 U15625 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n18906) );
  NAND2_X1 U15626 ( .A1(n12705), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12695) );
  INV_X1 U15627 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16238) );
  OR2_X1 U15628 ( .A1(n15033), .A2(n16238), .ZN(n12694) );
  NAND2_X1 U15629 ( .A1(n15033), .A2(BUF2_REG_12__SCAN_IN), .ZN(n12693) );
  NAND2_X1 U15630 ( .A1(n12694), .A2(n12693), .ZN(n18890) );
  NAND2_X1 U15631 ( .A1(n12737), .A2(n18890), .ZN(n12696) );
  OAI211_X1 U15632 ( .C1(n18906), .C2(n12811), .A(n12695), .B(n12696), .ZN(
        P2_U2979) );
  INV_X1 U15633 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n12827) );
  NAND2_X1 U15634 ( .A1(n12705), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12697) );
  OAI211_X1 U15635 ( .C1(n12827), .C2(n12811), .A(n12697), .B(n12696), .ZN(
        P2_U2964) );
  NAND2_X1 U15636 ( .A1(n12705), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n12699) );
  OAI211_X1 U15637 ( .C1(n10979), .C2(n12811), .A(n12699), .B(n12698), .ZN(
        P2_U2981) );
  INV_X1 U15638 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n12818) );
  NAND2_X1 U15639 ( .A1(n12705), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12702) );
  INV_X1 U15640 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16244) );
  OR2_X1 U15641 ( .A1(n15033), .A2(n16244), .ZN(n12701) );
  NAND2_X1 U15642 ( .A1(n15033), .A2(BUF2_REG_8__SCAN_IN), .ZN(n12700) );
  NAND2_X1 U15643 ( .A1(n12701), .A2(n12700), .ZN(n14587) );
  NAND2_X1 U15644 ( .A1(n12737), .A2(n14587), .ZN(n12703) );
  OAI211_X1 U15645 ( .C1(n12818), .C2(n12811), .A(n12702), .B(n12703), .ZN(
        P2_U2960) );
  NAND2_X1 U15646 ( .A1(n12705), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n12704) );
  OAI211_X1 U15647 ( .C1(n10899), .C2(n12811), .A(n12704), .B(n12703), .ZN(
        P2_U2975) );
  INV_X1 U15648 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12707) );
  INV_X1 U15649 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12706) );
  INV_X1 U15650 ( .A(n12705), .ZN(n12712) );
  AOI22_X1 U15651 ( .A1(n15034), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15033), .ZN(n13482) );
  OAI222_X1 U15652 ( .A1(n12707), .A2(n12811), .B1(n12706), .B2(n12712), .C1(
        n12741), .C2(n13482), .ZN(P2_U2982) );
  INV_X1 U15653 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12709) );
  INV_X1 U15654 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n12708) );
  INV_X1 U15655 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16260) );
  INV_X1 U15656 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n17972) );
  AOI22_X1 U15657 ( .A1(n15034), .A2(n16260), .B1(n17972), .B2(n15033), .ZN(
        n18879) );
  INV_X1 U15658 ( .A(n18879), .ZN(n18945) );
  OAI222_X1 U15659 ( .A1(n12811), .A2(n12709), .B1(n12708), .B2(n12712), .C1(
        n12741), .C2(n18945), .ZN(P2_U2967) );
  INV_X1 U15660 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n12710) );
  OAI222_X1 U15661 ( .A1(n12741), .A2(n18945), .B1(n12811), .B2(n11007), .C1(
        n12710), .C2(n12712), .ZN(P2_U2952) );
  INV_X1 U15662 ( .A(n12712), .ZN(n12747) );
  AOI22_X1 U15663 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n12711) );
  MUX2_X1 U15664 ( .A(BUF1_REG_13__SCAN_IN), .B(BUF2_REG_13__SCAN_IN), .S(
        n15033), .Z(n13919) );
  NAND2_X1 U15665 ( .A1(n12737), .A2(n13919), .ZN(n12713) );
  NAND2_X1 U15666 ( .A1(n12711), .A2(n12713), .ZN(P2_U2980) );
  AOI22_X1 U15667 ( .A1(P2_UWORD_REG_13__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n12714) );
  NAND2_X1 U15668 ( .A1(n12714), .A2(n12713), .ZN(P2_U2965) );
  AOI22_X1 U15669 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n12705), .B1(n12750), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n12715) );
  OAI22_X1 U15670 ( .A1(n15033), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n15034), .ZN(n15026) );
  INV_X1 U15671 ( .A(n15026), .ZN(n15834) );
  NAND2_X1 U15672 ( .A1(n12737), .A2(n15834), .ZN(n12743) );
  NAND2_X1 U15673 ( .A1(n12715), .A2(n12743), .ZN(P2_U2956) );
  AOI22_X1 U15674 ( .A1(P2_UWORD_REG_11__SCAN_IN), .A2(n12705), .B1(n12750), 
        .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n12719) );
  INV_X1 U15675 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n12716) );
  OR2_X1 U15676 ( .A1(n15033), .A2(n12716), .ZN(n12718) );
  NAND2_X1 U15677 ( .A1(n15033), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12717) );
  NAND2_X1 U15678 ( .A1(n12718), .A2(n12717), .ZN(n14565) );
  NAND2_X1 U15679 ( .A1(n12737), .A2(n14565), .ZN(n12722) );
  NAND2_X1 U15680 ( .A1(n12719), .A2(n12722), .ZN(P2_U2963) );
  AOI22_X1 U15681 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12720) );
  OAI22_X1 U15682 ( .A1(n15033), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n15034), .ZN(n18972) );
  INV_X1 U15683 ( .A(n18972), .ZN(n15828) );
  NAND2_X1 U15684 ( .A1(n12737), .A2(n15828), .ZN(n12734) );
  NAND2_X1 U15685 ( .A1(n12720), .A2(n12734), .ZN(P2_U2973) );
  AOI22_X1 U15686 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U15687 ( .A1(n15034), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15033), .ZN(n18951) );
  INV_X1 U15688 ( .A(n18951), .ZN(n13594) );
  NAND2_X1 U15689 ( .A1(n12737), .A2(n13594), .ZN(n12728) );
  NAND2_X1 U15690 ( .A1(n12721), .A2(n12728), .ZN(P2_U2953) );
  AOI22_X1 U15691 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n12723) );
  NAND2_X1 U15692 ( .A1(n12723), .A2(n12722), .ZN(P2_U2978) );
  AOI22_X1 U15693 ( .A1(P2_UWORD_REG_9__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n12727) );
  INV_X1 U15694 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n12724) );
  OR2_X1 U15695 ( .A1(n15033), .A2(n12724), .ZN(n12726) );
  NAND2_X1 U15696 ( .A1(n15033), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12725) );
  NAND2_X1 U15697 ( .A1(n12726), .A2(n12725), .ZN(n14580) );
  NAND2_X1 U15698 ( .A1(n12737), .A2(n14580), .ZN(n12730) );
  NAND2_X1 U15699 ( .A1(n12727), .A2(n12730), .ZN(P2_U2961) );
  AOI22_X1 U15700 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12729) );
  NAND2_X1 U15701 ( .A1(n12729), .A2(n12728), .ZN(P2_U2968) );
  AOI22_X1 U15702 ( .A1(P2_LWORD_REG_9__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n12731) );
  NAND2_X1 U15703 ( .A1(n12731), .A2(n12730), .ZN(P2_U2976) );
  AOI22_X1 U15704 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n12733) );
  AOI22_X1 U15705 ( .A1(n15034), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15033), .ZN(n18983) );
  INV_X1 U15706 ( .A(n18983), .ZN(n12732) );
  NAND2_X1 U15707 ( .A1(n12737), .A2(n12732), .ZN(n12751) );
  NAND2_X1 U15708 ( .A1(n12733), .A2(n12751), .ZN(P2_U2974) );
  AOI22_X1 U15709 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n12735) );
  NAND2_X1 U15710 ( .A1(n12735), .A2(n12734), .ZN(P2_U2958) );
  AOI22_X1 U15711 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12736) );
  AOI22_X1 U15712 ( .A1(n15034), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15033), .ZN(n15042) );
  INV_X1 U15713 ( .A(n15042), .ZN(n13671) );
  NAND2_X1 U15714 ( .A1(n12737), .A2(n13671), .ZN(n12739) );
  NAND2_X1 U15715 ( .A1(n12736), .A2(n12739), .ZN(P2_U2957) );
  AOI22_X1 U15716 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12738) );
  AOI22_X1 U15717 ( .A1(n15034), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15033), .ZN(n18966) );
  INV_X1 U15718 ( .A(n18966), .ZN(n13146) );
  NAND2_X1 U15719 ( .A1(n12737), .A2(n13146), .ZN(n12745) );
  NAND2_X1 U15720 ( .A1(n12738), .A2(n12745), .ZN(P2_U2955) );
  AOI22_X1 U15721 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12740) );
  NAND2_X1 U15722 ( .A1(n12740), .A2(n12739), .ZN(P2_U2972) );
  AOI22_X1 U15723 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n12742) );
  INV_X1 U15724 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16253) );
  INV_X1 U15725 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n17980) );
  AOI22_X1 U15726 ( .A1(n15034), .A2(n16253), .B1(n17980), .B2(n15033), .ZN(
        n15840) );
  INV_X1 U15727 ( .A(n15840), .ZN(n18959) );
  OR2_X1 U15728 ( .A1(n12741), .A2(n18959), .ZN(n12748) );
  NAND2_X1 U15729 ( .A1(n12742), .A2(n12748), .ZN(P2_U2954) );
  AOI22_X1 U15730 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12744) );
  NAND2_X1 U15731 ( .A1(n12744), .A2(n12743), .ZN(P2_U2971) );
  AOI22_X1 U15732 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n12746) );
  NAND2_X1 U15733 ( .A1(n12746), .A2(n12745), .ZN(P2_U2970) );
  AOI22_X1 U15734 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12749) );
  NAND2_X1 U15735 ( .A1(n12749), .A2(n12748), .ZN(P2_U2969) );
  AOI22_X1 U15736 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n12747), .B1(n12750), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12752) );
  NAND2_X1 U15737 ( .A1(n12752), .A2(n12751), .ZN(P2_U2959) );
  AND2_X1 U15738 ( .A1(n12792), .A2(n13052), .ZN(n12754) );
  NAND2_X1 U15739 ( .A1(n12753), .A2(n12754), .ZN(n12799) );
  AND2_X1 U15740 ( .A1(n20333), .A2(n15418), .ZN(n13486) );
  AOI21_X1 U15741 ( .B1(n12799), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n13486), 
        .ZN(n12755) );
  NAND2_X1 U15742 ( .A1(n13384), .A2(n12755), .ZN(P1_U2801) );
  XNOR2_X1 U15743 ( .A(n12758), .B(n12757), .ZN(n12940) );
  INV_X1 U15744 ( .A(n12940), .ZN(n12766) );
  XNOR2_X1 U15745 ( .A(n12760), .B(n12759), .ZN(n12941) );
  INV_X1 U15746 ( .A(n13449), .ZN(n13450) );
  NOR2_X1 U15747 ( .A1(n16010), .A2(n12761), .ZN(n12944) );
  INV_X1 U15748 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12762) );
  NOR2_X1 U15749 ( .A1(n15957), .A2(n12762), .ZN(n12763) );
  AOI211_X1 U15750 ( .C1(n15948), .C2(n13450), .A(n12944), .B(n12763), .ZN(
        n12764) );
  OAI21_X1 U15751 ( .B1(n12941), .B2(n15941), .A(n12764), .ZN(n12765) );
  AOI21_X1 U15752 ( .B1(n18936), .B2(n12766), .A(n12765), .ZN(n12767) );
  OAI21_X1 U15753 ( .B1(n12756), .B2(n15859), .A(n12767), .ZN(P2_U3012) );
  NOR2_X1 U15754 ( .A1(n16010), .A2(n12768), .ZN(n14971) );
  AOI21_X1 U15755 ( .B1(n14992), .B2(n12770), .A(n12769), .ZN(n14969) );
  AND2_X1 U15756 ( .A1(n18939), .A2(n14969), .ZN(n12771) );
  AOI211_X1 U15757 ( .C1(n18934), .C2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14971), .B(n12771), .ZN(n12776) );
  AOI21_X1 U15758 ( .B1(n12773), .B2(n13462), .A(n12772), .ZN(n12774) );
  XNOR2_X1 U15759 ( .A(n12774), .B(n14992), .ZN(n14970) );
  AOI22_X1 U15760 ( .A1(n14970), .A2(n18936), .B1(n15948), .B2(n13465), .ZN(
        n12775) );
  OAI211_X1 U15761 ( .C1(n12777), .C2(n15859), .A(n12776), .B(n12775), .ZN(
        P2_U3013) );
  XNOR2_X1 U15762 ( .A(n18816), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12883) );
  NOR2_X1 U15763 ( .A1(n16010), .A2(n10280), .ZN(n12882) );
  AOI21_X1 U15764 ( .B1(n12779), .B2(n14982), .A(n12778), .ZN(n12780) );
  INV_X1 U15765 ( .A(n12780), .ZN(n12880) );
  NOR2_X1 U15766 ( .A1(n15941), .A2(n12880), .ZN(n12781) );
  AOI211_X1 U15767 ( .C1(n18936), .C2(n12883), .A(n12882), .B(n12781), .ZN(
        n12784) );
  OAI21_X1 U15768 ( .B1(n18934), .B2(n12782), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12783) );
  OAI211_X1 U15769 ( .C1(n15859), .C2(n12845), .A(n12784), .B(n12783), .ZN(
        P2_U3014) );
  INV_X1 U15770 ( .A(n15424), .ZN(n12797) );
  INV_X1 U15771 ( .A(n12785), .ZN(n12803) );
  AOI21_X1 U15772 ( .B1(n12753), .B2(n12792), .A(n12803), .ZN(n12786) );
  AOI21_X1 U15773 ( .B1(n12797), .B2(n11756), .A(n12786), .ZN(n19630) );
  INV_X1 U15774 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20504) );
  NAND2_X1 U15775 ( .A1(n9731), .A2(n20504), .ZN(n15450) );
  NAND3_X1 U15776 ( .A1(n13897), .A2(n11756), .A3(n15450), .ZN(n12787) );
  NAND2_X1 U15777 ( .A1(n12787), .A2(n15448), .ZN(n20621) );
  NAND2_X1 U15778 ( .A1(n19630), .A2(n20621), .ZN(n15406) );
  AND2_X1 U15779 ( .A1(n15406), .A2(n13052), .ZN(n19639) );
  INV_X1 U15780 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n15407) );
  INV_X1 U15781 ( .A(n19868), .ZN(n12788) );
  OR2_X1 U15782 ( .A1(n13166), .A2(n11732), .ZN(n12791) );
  INV_X1 U15783 ( .A(n13341), .ZN(n12789) );
  NAND2_X1 U15784 ( .A1(n12789), .A2(n11690), .ZN(n12790) );
  AND2_X1 U15785 ( .A1(n12791), .A2(n12790), .ZN(n12899) );
  NOR2_X1 U15786 ( .A1(n15391), .A2(n11733), .ZN(n13046) );
  NAND2_X1 U15787 ( .A1(n12899), .A2(n13046), .ZN(n13191) );
  INV_X1 U15788 ( .A(n12792), .ZN(n12793) );
  AOI22_X1 U15789 ( .A1(n12797), .A2(n12803), .B1(n12753), .B2(n12793), .ZN(
        n12796) );
  INV_X1 U15790 ( .A(n13192), .ZN(n12794) );
  OAI21_X1 U15791 ( .B1(n12794), .B2(n13062), .A(n12797), .ZN(n12795) );
  OAI211_X1 U15792 ( .C1(n12797), .C2(n13191), .A(n12796), .B(n12795), .ZN(
        n15408) );
  NAND2_X1 U15793 ( .A1(n19639), .A2(n15408), .ZN(n12798) );
  OAI21_X1 U15794 ( .B1(n19639), .B2(n15407), .A(n12798), .ZN(P1_U3484) );
  INV_X1 U15795 ( .A(n20623), .ZN(n12801) );
  OAI21_X1 U15796 ( .B1(n13486), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n12801), 
        .ZN(n12800) );
  OAI21_X1 U15797 ( .B1(n12802), .B2(n12801), .A(n12800), .ZN(P1_U3487) );
  AND2_X1 U15798 ( .A1(n12753), .A2(n19858), .ZN(n15396) );
  INV_X1 U15799 ( .A(n15450), .ZN(n12804) );
  NAND2_X1 U15800 ( .A1(n15396), .A2(n12804), .ZN(n12911) );
  NAND2_X1 U15801 ( .A1(n12803), .A2(n11733), .ZN(n13076) );
  INV_X1 U15802 ( .A(n13076), .ZN(n12805) );
  NAND2_X1 U15803 ( .A1(n12805), .A2(n12804), .ZN(n15416) );
  AND2_X1 U15804 ( .A1(n12911), .A2(n15416), .ZN(n12806) );
  INV_X1 U15805 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12808) );
  NOR2_X1 U15806 ( .A1(n20437), .A2(n15418), .ZN(n15769) );
  NAND2_X1 U15807 ( .A1(n15769), .A2(n15763), .ZN(n19760) );
  INV_X1 U15808 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n20659) );
  INV_X1 U15809 ( .A(P1_UWORD_REG_9__SCAN_IN), .ZN(n12807) );
  OAI222_X1 U15810 ( .A1(n19743), .A2(n12808), .B1(n19747), .B2(n20659), .C1(
        n19760), .C2(n12807), .ZN(P1_U2911) );
  INV_X1 U15811 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12810) );
  INV_X1 U15812 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n20789) );
  INV_X1 U15813 ( .A(P1_UWORD_REG_3__SCAN_IN), .ZN(n12809) );
  OAI222_X1 U15814 ( .A1(n19743), .A2(n12810), .B1(n19747), .B2(n20789), .C1(
        n19760), .C2(n12809), .ZN(P1_U2917) );
  NAND2_X1 U15815 ( .A1(n12867), .A2(n16106), .ZN(n12812) );
  OAI21_X1 U15816 ( .B1(n12865), .B2(n12812), .A(n12811), .ZN(n12813) );
  NAND2_X1 U15817 ( .A1(n18921), .A2(n12814), .ZN(n12836) );
  NOR2_X1 U15818 ( .A1(n19606), .A2(n11065), .ZN(n15023) );
  INV_X1 U15819 ( .A(n15023), .ZN(n12862) );
  NOR2_X1 U15820 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12862), .ZN(n18904) );
  INV_X2 U15821 ( .A(n18923), .ZN(n18927) );
  AOI22_X1 U15822 ( .A1(n18930), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12815) );
  OAI21_X1 U15823 ( .B1(n12816), .B2(n12836), .A(n12815), .ZN(P2_U2925) );
  AOI22_X1 U15824 ( .A1(n18930), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12817) );
  OAI21_X1 U15825 ( .B1(n12818), .B2(n12836), .A(n12817), .ZN(P2_U2927) );
  INV_X1 U15826 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13673) );
  AOI22_X1 U15827 ( .A1(n18904), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12819) );
  OAI21_X1 U15828 ( .B1(n13673), .B2(n12836), .A(n12819), .ZN(P2_U2930) );
  INV_X1 U15829 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U15830 ( .A1(n18904), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n12820) );
  OAI21_X1 U15831 ( .B1(n12821), .B2(n12836), .A(n12820), .ZN(P2_U2929) );
  AOI22_X1 U15832 ( .A1(n18904), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12822) );
  OAI21_X1 U15833 ( .B1(n13615), .B2(n12836), .A(n12822), .ZN(P2_U2932) );
  INV_X1 U15834 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n14595) );
  AOI22_X1 U15835 ( .A1(n18904), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12823) );
  OAI21_X1 U15836 ( .B1(n14595), .B2(n12836), .A(n12823), .ZN(P2_U2928) );
  AOI22_X1 U15837 ( .A1(n18930), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12824) );
  OAI21_X1 U15838 ( .B1(n11599), .B2(n12836), .A(n12824), .ZN(P2_U2921) );
  AOI22_X1 U15839 ( .A1(n18904), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n12825) );
  OAI21_X1 U15840 ( .B1(n11007), .B2(n12836), .A(n12825), .ZN(P2_U2935) );
  AOI22_X1 U15841 ( .A1(n18930), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12826) );
  OAI21_X1 U15842 ( .B1(n12827), .B2(n12836), .A(n12826), .ZN(P2_U2923) );
  INV_X1 U15843 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n12829) );
  AOI22_X1 U15844 ( .A1(n18904), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12828) );
  OAI21_X1 U15845 ( .B1(n12829), .B2(n12836), .A(n12828), .ZN(P2_U2931) );
  AOI22_X1 U15846 ( .A1(n18904), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12830) );
  OAI21_X1 U15847 ( .B1(n11013), .B2(n12836), .A(n12830), .ZN(P2_U2933) );
  AOI22_X1 U15848 ( .A1(n18904), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n12831) );
  OAI21_X1 U15849 ( .B1(n12832), .B2(n12836), .A(n12831), .ZN(P2_U2934) );
  INV_X1 U15850 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13917) );
  AOI22_X1 U15851 ( .A1(n18930), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12833) );
  OAI21_X1 U15852 ( .B1(n13917), .B2(n12836), .A(n12833), .ZN(P2_U2922) );
  INV_X1 U15853 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14563) );
  AOI22_X1 U15854 ( .A1(n18930), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12834) );
  OAI21_X1 U15855 ( .B1(n14563), .B2(n12836), .A(n12834), .ZN(P2_U2924) );
  INV_X1 U15856 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14578) );
  AOI22_X1 U15857 ( .A1(n18930), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12835) );
  OAI21_X1 U15858 ( .B1(n14578), .B2(n12836), .A(n12835), .ZN(P2_U2926) );
  NOR2_X1 U15859 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12838) );
  OAI21_X1 U15860 ( .B1(n12839), .B2(n12838), .A(n12837), .ZN(n12840) );
  INV_X1 U15861 ( .A(n12840), .ZN(n12841) );
  INV_X1 U15862 ( .A(n16090), .ZN(n16092) );
  NAND2_X1 U15863 ( .A1(n16092), .A2(n16089), .ZN(n12864) );
  NAND2_X1 U15864 ( .A1(n14978), .A2(n12842), .ZN(n12974) );
  NAND2_X1 U15865 ( .A1(n12864), .A2(n12974), .ZN(n12843) );
  AND2_X2 U15866 ( .A1(n12843), .A2(n16106), .ZN(n18859) );
  NAND2_X1 U15867 ( .A1(n18859), .A2(n12844), .ZN(n18865) );
  MUX2_X1 U15868 ( .A(n12846), .B(n12845), .S(n18859), .Z(n12847) );
  OAI21_X1 U15869 ( .B1(n19608), .B2(n18865), .A(n12847), .ZN(P2_U2887) );
  OR2_X1 U15870 ( .A1(n12849), .A2(n12848), .ZN(n12850) );
  INV_X1 U15871 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n12852) );
  INV_X2 U15872 ( .A(n18859), .ZN(n18875) );
  MUX2_X1 U15873 ( .A(n12756), .B(n12852), .S(n18875), .Z(n12853) );
  OAI21_X1 U15874 ( .B1(n19592), .B2(n18865), .A(n12853), .ZN(P2_U2885) );
  INV_X1 U15875 ( .A(n12854), .ZN(n12855) );
  NAND2_X1 U15876 ( .A1(n14596), .A2(n12855), .ZN(n13483) );
  NOR2_X1 U15877 ( .A1(n12857), .A2(n12856), .ZN(n12858) );
  NOR2_X1 U15878 ( .A1(n12859), .A2(n12858), .ZN(n18809) );
  NAND2_X1 U15879 ( .A1(n19261), .A2(n18809), .ZN(n12927) );
  OAI211_X1 U15880 ( .C1(n19261), .C2(n18809), .A(n12927), .B(n18885), .ZN(
        n12861) );
  AOI22_X1 U15881 ( .A1(n18884), .A2(n18809), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n18893), .ZN(n12860) );
  OAI211_X1 U15882 ( .C1(n13483), .C2(n18945), .A(n12861), .B(n12860), .ZN(
        P2_U2919) );
  NOR2_X1 U15883 ( .A1(n18640), .A2(n12862), .ZN(n16121) );
  AND2_X1 U15884 ( .A1(n12864), .A2(n12863), .ZN(n12871) );
  INV_X1 U15885 ( .A(n12865), .ZN(n12868) );
  NAND3_X1 U15886 ( .A1(n12868), .A2(n12867), .A3(n12866), .ZN(n12869) );
  OAI22_X1 U15887 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19582), .B1(n16085), 
        .B2(n19494), .ZN(n12872) );
  AOI21_X1 U15888 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16121), .A(n12872), .ZN(
        n15018) );
  INV_X1 U15889 ( .A(n15018), .ZN(n12879) );
  INV_X1 U15890 ( .A(n12980), .ZN(n19496) );
  NAND2_X1 U15891 ( .A1(n12874), .A2(n12873), .ZN(n12875) );
  OR2_X1 U15892 ( .A1(n12876), .A2(n12875), .ZN(n16095) );
  OR3_X1 U15893 ( .A1(n15018), .A2(n19496), .A3(n16095), .ZN(n12877) );
  OAI21_X1 U15894 ( .B1(n12879), .B2(n12878), .A(n12877), .ZN(P2_U3595) );
  INV_X1 U15895 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n18917) );
  OAI222_X1 U15896 ( .A1(n18790), .A2(n18898), .B1(n13483), .B2(n18972), .C1(
        n18917), .C2(n14596), .ZN(P2_U2913) );
  INV_X1 U15897 ( .A(n14968), .ZN(n12937) );
  OAI22_X1 U15898 ( .A1(n12937), .A2(n14982), .B1(n16060), .B2(n12880), .ZN(
        n12881) );
  AOI211_X1 U15899 ( .C1(n16045), .C2(n18815), .A(n12882), .B(n12881), .ZN(
        n12885) );
  AOI22_X1 U15900 ( .A1(n16063), .A2(n12883), .B1(n16057), .B2(n18809), .ZN(
        n12884) );
  OAI211_X1 U15901 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n14940), .A(
        n12885), .B(n12884), .ZN(P2_U3046) );
  NAND2_X1 U15902 ( .A1(n19590), .A2(n18871), .ZN(n12889) );
  NAND2_X1 U15903 ( .A1(n18859), .A2(n14990), .ZN(n12888) );
  OAI211_X1 U15904 ( .C1(n18859), .C2(n10530), .A(n12889), .B(n12888), .ZN(
        P2_U2886) );
  MUX2_X1 U15905 ( .A(n10536), .B(n10350), .S(n18859), .Z(n12894) );
  OAI21_X1 U15906 ( .B1(n19581), .B2(n18865), .A(n12894), .ZN(P2_U2884) );
  INV_X1 U15907 ( .A(n12895), .ZN(n13070) );
  AND3_X1 U15908 ( .A1(n12910), .A2(n12896), .A3(n13070), .ZN(n12897) );
  AND2_X1 U15909 ( .A1(n12467), .A2(n12897), .ZN(n12906) );
  OAI21_X1 U15910 ( .B1(n12898), .B2(n11739), .A(n19858), .ZN(n12900) );
  AND2_X1 U15911 ( .A1(n12900), .A2(n12899), .ZN(n12905) );
  INV_X1 U15912 ( .A(n13382), .ZN(n20619) );
  NAND2_X1 U15913 ( .A1(n12962), .A2(n9618), .ZN(n12901) );
  NAND2_X1 U15914 ( .A1(n20619), .A2(n12901), .ZN(n12902) );
  NAND2_X1 U15915 ( .A1(n12903), .A2(n12902), .ZN(n12915) );
  AND3_X1 U15916 ( .A1(n12905), .A2(n12904), .A3(n12915), .ZN(n13069) );
  AND2_X1 U15917 ( .A1(n12906), .A2(n13069), .ZN(n15394) );
  INV_X1 U15918 ( .A(n15394), .ZN(n12907) );
  AOI22_X1 U15919 ( .A1(n11860), .A2(n12907), .B1(n13188), .B2(n11607), .ZN(
        n15398) );
  INV_X1 U15920 ( .A(n15398), .ZN(n12909) );
  OAI22_X1 U15921 ( .A1(n15418), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20597), .ZN(n12908) );
  AOI21_X1 U15922 ( .B1(n12909), .B2(n20595), .A(n12908), .ZN(n12924) );
  NAND2_X1 U15923 ( .A1(n12911), .A2(n12910), .ZN(n12913) );
  INV_X1 U15924 ( .A(n15448), .ZN(n20507) );
  AOI21_X1 U15925 ( .B1(n13897), .B2(n15450), .A(n20507), .ZN(n12912) );
  NAND2_X1 U15926 ( .A1(n12913), .A2(n12912), .ZN(n12914) );
  NAND2_X1 U15927 ( .A1(n12914), .A2(n13192), .ZN(n12921) );
  INV_X1 U15928 ( .A(n12753), .ZN(n12918) );
  NAND2_X1 U15929 ( .A1(n12916), .A2(n12915), .ZN(n12917) );
  NAND2_X1 U15930 ( .A1(n12918), .A2(n12917), .ZN(n13050) );
  OAI211_X1 U15931 ( .C1(n13341), .C2(n19863), .A(n12919), .B(n13050), .ZN(
        n12920) );
  AOI21_X1 U15932 ( .B1(n15424), .B2(n12921), .A(n12920), .ZN(n12922) );
  INV_X1 U15933 ( .A(n13052), .ZN(n19631) );
  NAND2_X1 U15934 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15769), .ZN(n15770) );
  INV_X1 U15935 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19638) );
  OAI22_X1 U15936 ( .A1(n15388), .A2(n19631), .B1(n15770), .B2(n19638), .ZN(
        n15761) );
  AOI21_X1 U15937 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n15763), .A(n15761), 
        .ZN(n20605) );
  AOI21_X1 U15938 ( .B1(n15396), .B2(n20595), .A(n20605), .ZN(n12923) );
  OAI22_X1 U15939 ( .A1(n12924), .A2(n20605), .B1(n12923), .B2(n11607), .ZN(
        P1_U3474) );
  XNOR2_X1 U15940 ( .A(n12925), .B(n12926), .ZN(n19601) );
  NOR2_X1 U15941 ( .A1(n19590), .A2(n19601), .ZN(n12988) );
  AOI21_X1 U15942 ( .B1(n19601), .B2(n19590), .A(n12988), .ZN(n12928) );
  NAND2_X1 U15943 ( .A1(n12928), .A2(n12927), .ZN(n12990) );
  OAI21_X1 U15944 ( .B1(n12928), .B2(n12927), .A(n12990), .ZN(n12929) );
  NAND2_X1 U15945 ( .A1(n12929), .A2(n18885), .ZN(n12932) );
  OAI22_X1 U15946 ( .A1(n13483), .A2(n18951), .B1(n14596), .B2(n18929), .ZN(
        n12930) );
  AOI21_X1 U15947 ( .B1(n18884), .B2(n19601), .A(n12930), .ZN(n12931) );
  NAND2_X1 U15948 ( .A1(n12932), .A2(n12931), .ZN(P2_U2918) );
  NAND2_X1 U15949 ( .A1(n12934), .A2(n12933), .ZN(n12936) );
  NAND2_X1 U15950 ( .A1(n12936), .A2(n9987), .ZN(n19594) );
  OAI21_X1 U15951 ( .B1(n12938), .B2(n14972), .A(n12937), .ZN(n12939) );
  AOI22_X1 U15952 ( .A1(n19594), .A2(n16057), .B1(n12939), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12949) );
  OAI22_X1 U15953 ( .A1(n16060), .A2(n12941), .B1(n16037), .B2(n12940), .ZN(
        n12942) );
  OR3_X1 U15954 ( .A1(n12944), .A2(n12943), .A3(n12942), .ZN(n12945) );
  AOI21_X1 U15955 ( .B1(n12947), .B2(n12946), .A(n12945), .ZN(n12948) );
  OAI211_X1 U15956 ( .C1(n12756), .C2(n16055), .A(n12949), .B(n12948), .ZN(
        P2_U3044) );
  OAI21_X1 U15957 ( .B1(n12951), .B2(n12950), .A(n13012), .ZN(n18775) );
  OAI222_X1 U15958 ( .A1(n13483), .A2(n18983), .B1(n18775), .B2(n18898), .C1(
        n18915), .C2(n14596), .ZN(P2_U2912) );
  NAND2_X1 U15959 ( .A1(n12952), .A2(n18861), .ZN(n13152) );
  XOR2_X1 U15960 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13152), .Z(n12959)
         );
  NAND2_X1 U15961 ( .A1(n12953), .A2(n13302), .ZN(n12956) );
  INV_X1 U15962 ( .A(n12954), .ZN(n12955) );
  AND2_X1 U15963 ( .A1(n12956), .A2(n12955), .ZN(n18804) );
  NOR2_X1 U15964 ( .A1(n18859), .A2(n18797), .ZN(n12957) );
  AOI21_X1 U15965 ( .B1(n18804), .B2(n18859), .A(n12957), .ZN(n12958) );
  OAI21_X1 U15966 ( .B1(n12959), .B2(n18865), .A(n12958), .ZN(P2_U2882) );
  OAI21_X1 U15967 ( .B1(n12961), .B2(n12960), .A(n13089), .ZN(n13362) );
  NAND2_X1 U15968 ( .A1(n12962), .A2(n11844), .ZN(n12963) );
  NAND2_X1 U15969 ( .A1(n19840), .A2(DATAI_1_), .ZN(n12965) );
  NAND2_X1 U15970 ( .A1(n19839), .A2(BUF1_REG_1__SCAN_IN), .ZN(n12964) );
  AND2_X1 U15971 ( .A1(n12965), .A2(n12964), .ZN(n19860) );
  INV_X1 U15972 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19775) );
  OAI222_X1 U15973 ( .A1(n13362), .A2(n14209), .B1(n14213), .B2(n19860), .C1(
        n14210), .C2(n19775), .ZN(P1_U2903) );
  INV_X1 U15974 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12966) );
  NOR2_X1 U15975 ( .A1(n13152), .A2(n12966), .ZN(n12968) );
  OR2_X1 U15976 ( .A1(n13152), .A2(n12967), .ZN(n13039) );
  OAI211_X1 U15977 ( .C1(n12968), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n18871), .B(n13039), .ZN(n12970) );
  NAND2_X1 U15978 ( .A1(n18859), .A2(n13556), .ZN(n12969) );
  OAI211_X1 U15979 ( .C1(n18859), .C2(n10604), .A(n12970), .B(n12969), .ZN(
        P2_U2881) );
  INV_X1 U15980 ( .A(n19581), .ZN(n13176) );
  OR2_X1 U15981 ( .A1(n16091), .A2(n16089), .ZN(n15009) );
  NOR2_X1 U15982 ( .A1(n12971), .A2(n15019), .ZN(n15001) );
  INV_X1 U15983 ( .A(n15001), .ZN(n12972) );
  AOI22_X1 U15984 ( .A1(n15009), .A2(n12972), .B1(n15005), .B2(n15006), .ZN(
        n12977) );
  NAND2_X1 U15985 ( .A1(n12974), .A2(n12973), .ZN(n15002) );
  INV_X1 U15986 ( .A(n15006), .ZN(n14988) );
  NOR2_X1 U15987 ( .A1(n14988), .A2(n15005), .ZN(n12975) );
  AOI211_X1 U15988 ( .C1(n15002), .C2(n11399), .A(n12975), .B(n15001), .ZN(
        n12976) );
  MUX2_X1 U15989 ( .A(n12977), .B(n12976), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12978) );
  OAI211_X1 U15990 ( .C1(n12893), .C2(n14978), .A(n12979), .B(n12978), .ZN(
        n16070) );
  AOI22_X1 U15991 ( .A1(n13176), .A2(n16115), .B1(n12980), .B2(n16070), .ZN(
        n12982) );
  NAND2_X1 U15992 ( .A1(n15018), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12981) );
  OAI21_X1 U15993 ( .B1(n12982), .B2(n15018), .A(n12981), .ZN(P2_U3596) );
  INV_X1 U15994 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13075) );
  XNOR2_X1 U15995 ( .A(n12983), .B(n13075), .ZN(n13087) );
  INV_X1 U15996 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20609) );
  NOR2_X1 U15997 ( .A1(n15731), .A2(n20609), .ZN(n13078) );
  AOI21_X1 U15998 ( .B1(n19813), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13078), .ZN(n12984) );
  OAI21_X1 U15999 ( .B1(n15597), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n12984), .ZN(n12985) );
  AOI21_X1 U16000 ( .B1(n19817), .B2(n13087), .A(n12985), .ZN(n12986) );
  OAI21_X1 U16001 ( .B1(n19841), .B2(n13362), .A(n12986), .ZN(P1_U2998) );
  INV_X1 U16002 ( .A(n19594), .ZN(n13455) );
  NAND2_X1 U16003 ( .A1(n19592), .A2(n13455), .ZN(n13141) );
  OAI21_X1 U16004 ( .B1(n19592), .B2(n13455), .A(n13141), .ZN(n12987) );
  INV_X1 U16005 ( .A(n12987), .ZN(n12992) );
  INV_X1 U16006 ( .A(n12988), .ZN(n12989) );
  NAND2_X1 U16007 ( .A1(n12990), .A2(n12989), .ZN(n12991) );
  NAND2_X1 U16008 ( .A1(n12991), .A2(n12992), .ZN(n13142) );
  OAI21_X1 U16009 ( .B1(n12992), .B2(n12991), .A(n13142), .ZN(n12993) );
  NAND2_X1 U16010 ( .A1(n12993), .A2(n18885), .ZN(n12995) );
  INV_X1 U16011 ( .A(n13483), .ZN(n18895) );
  AOI22_X1 U16012 ( .A1(n18895), .A2(n15840), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n18893), .ZN(n12994) );
  OAI211_X1 U16013 ( .C1(n13455), .C2(n14585), .A(n12995), .B(n12994), .ZN(
        P2_U2917) );
  NOR2_X1 U16014 ( .A1(n12996), .A2(n13897), .ZN(n12997) );
  NAND2_X1 U16015 ( .A1(n12998), .A2(n12997), .ZN(n12999) );
  NAND2_X1 U16016 ( .A1(n13000), .A2(n12999), .ZN(n13001) );
  NAND2_X1 U16017 ( .A1(n13832), .A2(n13075), .ZN(n13004) );
  INV_X1 U16018 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13002) );
  NAND2_X1 U16019 ( .A1(n13838), .A2(n13002), .ZN(n13003) );
  NAND3_X1 U16020 ( .A1(n13004), .A2(n13007), .A3(n13003), .ZN(n13005) );
  NAND2_X1 U16021 ( .A1(n13832), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13009) );
  INV_X1 U16022 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13373) );
  NAND2_X1 U16023 ( .A1(n13007), .A2(n13373), .ZN(n13008) );
  NAND2_X1 U16024 ( .A1(n13009), .A2(n13008), .ZN(n13115) );
  XNOR2_X1 U16025 ( .A(n13093), .B(n13115), .ZN(n13010) );
  NAND2_X1 U16026 ( .A1(n13010), .A2(n13838), .ZN(n13094) );
  OAI21_X1 U16027 ( .B1(n13010), .B2(n13838), .A(n13094), .ZN(n13360) );
  AOI22_X1 U16028 ( .A1(n19738), .A2(n13360), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14134), .ZN(n13011) );
  OAI21_X1 U16029 ( .B1(n13362), .B2(n14144), .A(n13011), .ZN(P1_U2871) );
  INV_X1 U16030 ( .A(n14587), .ZN(n13015) );
  AOI21_X1 U16031 ( .B1(n13013), .B2(n13012), .A(n13126), .ZN(n16016) );
  INV_X1 U16032 ( .A(n16016), .ZN(n13014) );
  OAI222_X1 U16033 ( .A1(n13483), .A2(n13015), .B1(n13014), .B2(n18898), .C1(
        n10899), .C2(n14596), .ZN(P2_U2911) );
  INV_X1 U16034 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13017) );
  INV_X1 U16035 ( .A(n19760), .ZN(n19771) );
  CLKBUF_X1 U16036 ( .A(n19771), .Z(n19777) );
  AOI22_X1 U16037 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n19777), .B1(n19776), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13016) );
  OAI21_X1 U16038 ( .B1(n13017), .B2(n19743), .A(n13016), .ZN(P1_U2908) );
  INV_X1 U16039 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13019) );
  AOI22_X1 U16040 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n19777), .B1(n19776), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13018) );
  OAI21_X1 U16041 ( .B1(n13019), .B2(n19743), .A(n13018), .ZN(P1_U2916) );
  INV_X1 U16042 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13021) );
  AOI22_X1 U16043 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n19777), .B1(n19776), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13020) );
  OAI21_X1 U16044 ( .B1(n13021), .B2(n19743), .A(n13020), .ZN(P1_U2910) );
  AOI22_X1 U16045 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n19777), .B1(n19776), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13022) );
  OAI21_X1 U16046 ( .B1(n14175), .B2(n19743), .A(n13022), .ZN(P1_U2915) );
  INV_X1 U16047 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13024) );
  AOI22_X1 U16048 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n19777), .B1(n19776), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13023) );
  OAI21_X1 U16049 ( .B1(n13024), .B2(n19743), .A(n13023), .ZN(P1_U2919) );
  INV_X1 U16050 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13026) );
  AOI22_X1 U16051 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n19777), .B1(n19776), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13025) );
  OAI21_X1 U16052 ( .B1(n13026), .B2(n19743), .A(n13025), .ZN(P1_U2913) );
  INV_X1 U16053 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13028) );
  AOI22_X1 U16054 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n19777), .B1(n19776), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13027) );
  OAI21_X1 U16055 ( .B1(n13028), .B2(n19743), .A(n13027), .ZN(P1_U2909) );
  INV_X1 U16056 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13030) );
  AOI22_X1 U16057 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n19777), .B1(n19776), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13029) );
  OAI21_X1 U16058 ( .B1(n13030), .B2(n19743), .A(n13029), .ZN(P1_U2907) );
  INV_X1 U16059 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13032) );
  AOI22_X1 U16060 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n19777), .B1(n19776), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13031) );
  OAI21_X1 U16061 ( .B1(n13032), .B2(n19743), .A(n13031), .ZN(P1_U2918) );
  INV_X1 U16062 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13034) );
  AOI22_X1 U16063 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n19777), .B1(n19776), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13033) );
  OAI21_X1 U16064 ( .B1(n13034), .B2(n19743), .A(n13033), .ZN(P1_U2912) );
  INV_X1 U16065 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13036) );
  AOI22_X1 U16066 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n19777), .B1(n19776), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13035) );
  OAI21_X1 U16067 ( .B1(n13036), .B2(n19743), .A(n13035), .ZN(P1_U2920) );
  INV_X1 U16068 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13038) );
  AOI22_X1 U16069 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n19777), .B1(n19776), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13037) );
  OAI21_X1 U16070 ( .B1(n13038), .B2(n19743), .A(n13037), .ZN(P1_U2914) );
  XOR2_X1 U16071 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n13039), .Z(n13045)
         );
  NAND2_X1 U16072 ( .A1(n13041), .A2(n13040), .ZN(n13042) );
  NAND2_X1 U16073 ( .A1(n13320), .A2(n13042), .ZN(n18774) );
  MUX2_X1 U16074 ( .A(n13043), .B(n18774), .S(n18859), .Z(n13044) );
  OAI21_X1 U16075 ( .B1(n13045), .B2(n18865), .A(n13044), .ZN(P2_U2880) );
  INV_X1 U16076 ( .A(n13046), .ZN(n13051) );
  NAND2_X1 U16077 ( .A1(n19858), .A2(n15450), .ZN(n13048) );
  NAND3_X1 U16078 ( .A1(n13048), .A2(n19863), .A3(n13047), .ZN(n13049) );
  OAI211_X1 U16079 ( .C1(n15424), .C2(n13051), .A(n13050), .B(n13049), .ZN(
        n13053) );
  NAND2_X1 U16080 ( .A1(n13053), .A2(n13052), .ZN(n13060) );
  NAND2_X1 U16081 ( .A1(n11733), .A2(n15450), .ZN(n13352) );
  NAND2_X1 U16082 ( .A1(n13054), .A2(n9618), .ZN(n13055) );
  AOI21_X1 U16083 ( .B1(n13056), .B2(n13352), .A(n13055), .ZN(n13057) );
  INV_X1 U16084 ( .A(n13062), .ZN(n13063) );
  OAI211_X1 U16085 ( .C1(n13064), .C2(n13061), .A(n13063), .B(n13192), .ZN(
        n13066) );
  OR2_X1 U16086 ( .A1(n13066), .A2(n13065), .ZN(n13067) );
  INV_X1 U16087 ( .A(n19833), .ZN(n13072) );
  OAI211_X1 U16088 ( .C1(n13070), .C2(n9618), .A(n13069), .B(n13068), .ZN(
        n13071) );
  NAND2_X1 U16089 ( .A1(n13081), .A2(n13071), .ZN(n19828) );
  AND2_X2 U16090 ( .A1(n13072), .A2(n19828), .ZN(n15674) );
  INV_X1 U16091 ( .A(n13191), .ZN(n13073) );
  NOR2_X1 U16092 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n19833), .ZN(
        n13253) );
  INV_X1 U16093 ( .A(n13253), .ZN(n13074) );
  NAND2_X1 U16094 ( .A1(n13075), .A2(n13074), .ZN(n13080) );
  OAI21_X1 U16095 ( .B1(n13061), .B2(n11737), .A(n13076), .ZN(n13077) );
  AOI21_X1 U16096 ( .B1(n19826), .B2(n13360), .A(n13078), .ZN(n13079) );
  OAI21_X1 U16097 ( .B1(n15702), .B2(n13080), .A(n13079), .ZN(n13086) );
  INV_X1 U16098 ( .A(n19829), .ZN(n14411) );
  INV_X1 U16099 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19830) );
  OR2_X1 U16100 ( .A1(n19828), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13084) );
  INV_X1 U16101 ( .A(n13081), .ZN(n13082) );
  NAND2_X1 U16102 ( .A1(n13082), .A2(n15731), .ZN(n13083) );
  AOI21_X1 U16103 ( .B1(n14411), .B2(n19830), .A(n15676), .ZN(n19827) );
  NOR2_X1 U16104 ( .A1(n19827), .A2(n13075), .ZN(n13085) );
  AOI211_X1 U16105 ( .C1(n19824), .C2(n13087), .A(n13086), .B(n13085), .ZN(
        n13088) );
  INV_X1 U16106 ( .A(n13088), .ZN(P1_U3030) );
  NAND2_X1 U16107 ( .A1(n13090), .A2(n13089), .ZN(n13091) );
  AND2_X1 U16108 ( .A1(n13092), .A2(n13091), .ZN(n19728) );
  INV_X1 U16109 ( .A(n19728), .ZN(n13114) );
  OR2_X1 U16110 ( .A1(n13831), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n13098) );
  NAND2_X1 U16111 ( .A1(n13832), .A2(n13844), .ZN(n13096) );
  INV_X1 U16112 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n19716) );
  NAND2_X1 U16113 ( .A1(n13838), .A2(n19716), .ZN(n13095) );
  NAND3_X1 U16114 ( .A1(n13096), .A2(n13821), .A3(n13095), .ZN(n13097) );
  NAND2_X1 U16115 ( .A1(n13170), .A2(n13102), .ZN(n19717) );
  INV_X1 U16116 ( .A(n19717), .ZN(n13103) );
  AOI22_X1 U16117 ( .A1(n19738), .A2(n13103), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n14134), .ZN(n13104) );
  OAI21_X1 U16118 ( .B1(n13114), .B2(n14136), .A(n13104), .ZN(P1_U2870) );
  AND2_X1 U16119 ( .A1(n12952), .A2(n13105), .ZN(n18864) );
  NAND2_X1 U16120 ( .A1(n12952), .A2(n13106), .ZN(n18853) );
  OAI211_X1 U16121 ( .C1(n18864), .C2(n13107), .A(n18871), .B(n18853), .ZN(
        n13111) );
  NOR2_X1 U16122 ( .A1(n13321), .A2(n13108), .ZN(n13109) );
  OR2_X1 U16123 ( .A1(n15899), .A2(n13109), .ZN(n16001) );
  INV_X1 U16124 ( .A(n16001), .ZN(n18764) );
  NAND2_X1 U16125 ( .A1(n18764), .A2(n18859), .ZN(n13110) );
  OAI211_X1 U16126 ( .C1(n18859), .C2(n11083), .A(n13111), .B(n13110), .ZN(
        P2_U2878) );
  NAND2_X1 U16127 ( .A1(n19840), .A2(DATAI_2_), .ZN(n13113) );
  NAND2_X1 U16128 ( .A1(n19839), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13112) );
  AND2_X1 U16129 ( .A1(n13113), .A2(n13112), .ZN(n19865) );
  INV_X1 U16130 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19773) );
  OAI222_X1 U16131 ( .A1(n13114), .A2(n14209), .B1(n14213), .B2(n19865), .C1(
        n14210), .C2(n19773), .ZN(P1_U2902) );
  OAI21_X1 U16132 ( .B1(n13898), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13115), .ZN(n19822) );
  NAND2_X1 U16133 ( .A1(n13117), .A2(n13116), .ZN(n13118) );
  NAND2_X1 U16134 ( .A1(n13119), .A2(n13118), .ZN(n19821) );
  OAI222_X1 U16135 ( .A1(n19822), .A2(n14146), .B1(n13373), .B2(n19742), .C1(
        n19821), .C2(n14144), .ZN(P1_U2872) );
  XNOR2_X1 U16136 ( .A(n13121), .B(n13120), .ZN(n13138) );
  INV_X1 U16137 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13123) );
  NAND2_X1 U16138 ( .A1(n15600), .A2(n19714), .ZN(n13122) );
  INV_X1 U16139 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n19706) );
  OR2_X1 U16140 ( .A1(n15731), .A2(n19706), .ZN(n13133) );
  OAI211_X1 U16141 ( .C1(n15603), .C2(n13123), .A(n13122), .B(n13133), .ZN(
        n13124) );
  AOI21_X1 U16142 ( .B1(n19728), .B2(n14290), .A(n13124), .ZN(n13125) );
  OAI21_X1 U16143 ( .B1(n19637), .B2(n13138), .A(n13125), .ZN(P1_U2997) );
  INV_X1 U16144 ( .A(n14580), .ZN(n13128) );
  OAI21_X1 U16145 ( .B1(n13127), .B2(n13126), .A(n15988), .ZN(n18768) );
  INV_X1 U16146 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n18912) );
  OAI222_X1 U16147 ( .A1(n13483), .A2(n13128), .B1(n18768), .B2(n18898), .C1(
        n18912), .C2(n14596), .ZN(P2_U2910) );
  NAND2_X1 U16148 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13130) );
  AOI21_X1 U16149 ( .B1(n13075), .B2(n15720), .A(n15676), .ZN(n13129) );
  OAI21_X1 U16150 ( .B1(n19829), .B2(n13130), .A(n13129), .ZN(n13136) );
  AOI21_X1 U16151 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13846) );
  INV_X1 U16152 ( .A(n13846), .ZN(n13131) );
  OR2_X1 U16153 ( .A1(n19829), .A2(n13131), .ZN(n13254) );
  INV_X1 U16154 ( .A(n13254), .ZN(n13135) );
  OR4_X1 U16155 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n15674), .A3(
        n13253), .A4(n13075), .ZN(n13132) );
  OAI211_X1 U16156 ( .C1(n15733), .C2(n19717), .A(n13133), .B(n13132), .ZN(
        n13134) );
  AOI211_X1 U16157 ( .C1(n13136), .C2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n13135), .B(n13134), .ZN(n13137) );
  OAI21_X1 U16158 ( .B1(n15685), .B2(n13138), .A(n13137), .ZN(P1_U3029) );
  XOR2_X1 U16159 ( .A(n13140), .B(n13139), .Z(n16058) );
  INV_X1 U16160 ( .A(n16058), .ZN(n19583) );
  XNOR2_X1 U16161 ( .A(n16058), .B(n19581), .ZN(n13144) );
  NAND2_X1 U16162 ( .A1(n13142), .A2(n13141), .ZN(n13143) );
  NAND2_X1 U16163 ( .A1(n13143), .A2(n13144), .ZN(n13175) );
  OAI21_X1 U16164 ( .B1(n13144), .B2(n13143), .A(n13175), .ZN(n13145) );
  NAND2_X1 U16165 ( .A1(n13145), .A2(n18885), .ZN(n13148) );
  AOI22_X1 U16166 ( .A1(n18895), .A2(n13146), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n18893), .ZN(n13147) );
  OAI211_X1 U16167 ( .C1(n19583), .C2(n14585), .A(n13148), .B(n13147), .ZN(
        P2_U2916) );
  NAND2_X1 U16168 ( .A1(n19840), .A2(DATAI_0_), .ZN(n13150) );
  NAND2_X1 U16169 ( .A1(n19839), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13149) );
  AND2_X1 U16170 ( .A1(n13150), .A2(n13149), .ZN(n19851) );
  INV_X1 U16171 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19780) );
  OAI222_X1 U16172 ( .A1(n19821), .A2(n14209), .B1(n14213), .B2(n19851), .C1(
        n14210), .C2(n19780), .ZN(P1_U2904) );
  INV_X1 U16173 ( .A(n18898), .ZN(n13161) );
  OR2_X1 U16174 ( .A1(n12952), .A2(n18861), .ZN(n13151) );
  NAND2_X1 U16175 ( .A1(n13152), .A2(n13151), .ZN(n13312) );
  INV_X1 U16176 ( .A(n13312), .ZN(n18872) );
  NAND2_X1 U16177 ( .A1(n13154), .A2(n13153), .ZN(n13157) );
  INV_X1 U16178 ( .A(n13155), .ZN(n13156) );
  AND2_X1 U16179 ( .A1(n13157), .A2(n13156), .ZN(n13517) );
  NAND2_X1 U16180 ( .A1(n18872), .A2(n13517), .ZN(n13179) );
  OAI21_X1 U16181 ( .B1(n13155), .B2(n13159), .A(n13158), .ZN(n18808) );
  OAI21_X1 U16182 ( .B1(n13179), .B2(n14601), .A(n18808), .ZN(n13160) );
  AOI222_X1 U16183 ( .A1(n13161), .A2(n13160), .B1(n18893), .B2(
        P2_EAX_REG_5__SCAN_IN), .C1(n13671), .C2(n18895), .ZN(n13162) );
  INV_X1 U16184 ( .A(n13162), .ZN(P2_U2914) );
  OAI21_X1 U16185 ( .B1(n13165), .B2(n13164), .A(n13163), .ZN(n19701) );
  INV_X1 U16186 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13172) );
  NAND2_X1 U16187 ( .A1(n12517), .A2(n13166), .ZN(n13168) );
  MUX2_X1 U16188 ( .A(n13829), .B(n13821), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13167) );
  NAND2_X1 U16189 ( .A1(n13168), .A2(n13167), .ZN(n13169) );
  AND2_X1 U16190 ( .A1(n13170), .A2(n13169), .ZN(n13171) );
  OR2_X1 U16191 ( .A1(n13171), .A2(n13260), .ZN(n19697) );
  OAI222_X1 U16192 ( .A1(n19701), .A2(n14136), .B1(n13172), .B2(n19742), .C1(
        n19697), .C2(n14146), .ZN(P1_U2869) );
  NAND2_X1 U16193 ( .A1(n19840), .A2(DATAI_3_), .ZN(n13174) );
  NAND2_X1 U16194 ( .A1(n19839), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13173) );
  AND2_X1 U16195 ( .A1(n13174), .A2(n13173), .ZN(n19870) );
  INV_X1 U16196 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19770) );
  OAI222_X1 U16197 ( .A1(n19701), .A2(n14209), .B1(n14213), .B2(n19870), .C1(
        n14210), .C2(n19770), .ZN(P1_U2901) );
  OAI21_X1 U16198 ( .B1(n13176), .B2(n16058), .A(n13175), .ZN(n13178) );
  INV_X1 U16199 ( .A(n13517), .ZN(n13177) );
  NAND3_X1 U16200 ( .A1(n13178), .A2(n13177), .A3(n13312), .ZN(n13180) );
  NAND3_X1 U16201 ( .A1(n13180), .A2(n18885), .A3(n13179), .ZN(n13182) );
  AOI22_X1 U16202 ( .A1(n18884), .A2(n13517), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n18893), .ZN(n13181) );
  OAI211_X1 U16203 ( .C1(n15026), .C2(n13483), .A(n13182), .B(n13181), .ZN(
        P2_U2915) );
  INV_X1 U16204 ( .A(n14565), .ZN(n13186) );
  INV_X1 U16205 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n18908) );
  OAI21_X1 U16206 ( .B1(n13185), .B2(n13184), .A(n13183), .ZN(n18746) );
  OAI222_X1 U16207 ( .A1(n13483), .A2(n13186), .B1(n14596), .B2(n18908), .C1(
        n18746), .C2(n18898), .ZN(P2_U2908) );
  NOR2_X1 U16208 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n15418), .ZN(n13221) );
  OR2_X1 U16209 ( .A1(n13187), .A2(n15394), .ZN(n13197) );
  AND2_X1 U16210 ( .A1(n13337), .A2(n11739), .ZN(n13189) );
  NAND2_X1 U16211 ( .A1(n13189), .A2(n13188), .ZN(n13203) );
  INV_X1 U16212 ( .A(n15389), .ZN(n20599) );
  NAND2_X1 U16213 ( .A1(n20599), .A2(n11606), .ZN(n13202) );
  NAND2_X1 U16214 ( .A1(n15389), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13204) );
  NAND2_X1 U16215 ( .A1(n13202), .A2(n13204), .ZN(n14450) );
  XNOR2_X1 U16216 ( .A(n11606), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13190) );
  NAND2_X1 U16217 ( .A1(n15396), .A2(n13190), .ZN(n13194) );
  NAND2_X1 U16218 ( .A1(n13192), .A2(n13191), .ZN(n13208) );
  NAND2_X1 U16219 ( .A1(n13208), .A2(n14450), .ZN(n13193) );
  OAI211_X1 U16220 ( .C1(n13203), .C2(n14450), .A(n13194), .B(n13193), .ZN(
        n13195) );
  INV_X1 U16221 ( .A(n13195), .ZN(n13196) );
  NAND2_X1 U16222 ( .A1(n13197), .A2(n13196), .ZN(n14447) );
  OR2_X1 U16223 ( .A1(n15388), .A2(n14447), .ZN(n13199) );
  NAND2_X1 U16224 ( .A1(n15388), .A2(n11606), .ZN(n13198) );
  NAND2_X1 U16225 ( .A1(n13199), .A2(n13198), .ZN(n15402) );
  INV_X1 U16226 ( .A(n15402), .ZN(n13200) );
  AOI22_X1 U16227 ( .A1(n13221), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n13200), .B2(n15418), .ZN(n13215) );
  INV_X1 U16228 ( .A(n13201), .ZN(n13227) );
  XNOR2_X1 U16229 ( .A(n13202), .B(n11605), .ZN(n13207) );
  INV_X1 U16230 ( .A(n13203), .ZN(n13206) );
  NAND2_X1 U16231 ( .A1(n13204), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13205) );
  NAND2_X1 U16232 ( .A1(n11770), .A2(n13205), .ZN(n20589) );
  AOI22_X1 U16233 ( .A1(n13208), .A2(n13207), .B1(n13206), .B2(n20589), .ZN(
        n13213) );
  NAND2_X1 U16234 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13209) );
  AOI22_X1 U16235 ( .A1(n13210), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n11605), .B2(n13209), .ZN(n13211) );
  NAND2_X1 U16236 ( .A1(n15396), .A2(n13211), .ZN(n13212) );
  OAI211_X1 U16237 ( .C1(n13227), .C2(n15394), .A(n13213), .B(n13212), .ZN(
        n20588) );
  MUX2_X1 U16238 ( .A(n20588), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15388), .Z(n15404) );
  AOI22_X1 U16239 ( .A1(n13221), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n15418), .B2(n15404), .ZN(n13214) );
  NOR2_X1 U16240 ( .A1(n13215), .A2(n13214), .ZN(n15411) );
  INV_X1 U16241 ( .A(n15390), .ZN(n20600) );
  NAND2_X1 U16242 ( .A1(n15411), .A2(n20600), .ZN(n13235) );
  INV_X1 U16243 ( .A(n20003), .ZN(n20291) );
  OR2_X1 U16244 ( .A1(n13216), .A2(n20291), .ZN(n13218) );
  XNOR2_X1 U16245 ( .A(n13218), .B(n13217), .ZN(n19684) );
  NOR2_X1 U16246 ( .A1(n19684), .A2(n12467), .ZN(n15760) );
  NOR2_X1 U16247 ( .A1(n15760), .A2(n15388), .ZN(n13219) );
  AOI211_X1 U16248 ( .C1(n15388), .C2(n13217), .A(P1_STATE2_REG_1__SCAN_IN), 
        .B(n13219), .ZN(n13220) );
  AOI21_X1 U16249 ( .B1(n13221), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13220), .ZN(n15413) );
  AND3_X1 U16250 ( .A1(n13235), .A2(n19638), .A3(n15413), .ZN(n13222) );
  OAI21_X1 U16251 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(
        P1_STATE2_REG_1__SCAN_IN), .A(n15763), .ZN(n20620) );
  OAI21_X1 U16252 ( .B1(n13222), .B2(n15770), .A(n19899), .ZN(n19837) );
  INV_X1 U16253 ( .A(n19837), .ZN(n13234) );
  NOR2_X1 U16254 ( .A1(n13223), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13231) );
  INV_X1 U16255 ( .A(n13225), .ZN(n13226) );
  OAI21_X1 U16256 ( .B1(n9635), .B2(n20382), .A(n20257), .ZN(n13230) );
  NAND2_X1 U16257 ( .A1(n20333), .A2(n20334), .ZN(n20289) );
  INV_X1 U16258 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20294) );
  AND2_X1 U16259 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20294), .ZN(n14445) );
  OAI22_X1 U16260 ( .A1(n19842), .A2(n20289), .B1(n13227), .B2(n14445), .ZN(
        n13229) );
  NAND2_X1 U16261 ( .A1(n9635), .A2(n13231), .ZN(n14443) );
  NOR2_X1 U16262 ( .A1(n20111), .A2(n14443), .ZN(n20118) );
  AOI211_X1 U16263 ( .C1(n13231), .C2(n13230), .A(n13229), .B(n20118), .ZN(
        n13233) );
  OR2_X1 U16264 ( .A1(n19837), .A2(n20217), .ZN(n13232) );
  OAI21_X1 U16265 ( .B1(n13234), .B2(n13233), .A(n13232), .ZN(P1_U3475) );
  AND3_X1 U16266 ( .A1(n13235), .A2(n15413), .A3(n15769), .ZN(n15420) );
  OAI22_X1 U16267 ( .A1(n19925), .A2(n20442), .B1(n13236), .B2(n14445), .ZN(
        n13237) );
  OAI21_X1 U16268 ( .B1(n15420), .B2(n13237), .A(n19837), .ZN(n13238) );
  OAI21_X1 U16269 ( .B1(n19837), .B2(n20639), .A(n13238), .ZN(P1_U3478) );
  XNOR2_X1 U16270 ( .A(n9652), .B(n18845), .ZN(n13244) );
  NAND2_X1 U16271 ( .A1(n13239), .A2(n15900), .ZN(n13241) );
  INV_X1 U16272 ( .A(n15874), .ZN(n13240) );
  NOR2_X1 U16273 ( .A1(n18859), .A2(n18736), .ZN(n13242) );
  AOI21_X1 U16274 ( .B1(n18742), .B2(n18859), .A(n13242), .ZN(n13243) );
  OAI21_X1 U16275 ( .B1(n13244), .B2(n18865), .A(n13243), .ZN(P2_U2876) );
  XOR2_X1 U16276 ( .A(n13246), .B(n13245), .Z(n13296) );
  NAND2_X1 U16277 ( .A1(n13296), .A2(n19817), .ZN(n13250) );
  INV_X2 U16278 ( .A(n15731), .ZN(n19819) );
  NAND2_X1 U16279 ( .A1(n19819), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n13293) );
  INV_X1 U16280 ( .A(n13293), .ZN(n13248) );
  NOR2_X1 U16281 ( .A1(n15597), .A2(n19702), .ZN(n13247) );
  AOI211_X1 U16282 ( .C1(n19813), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13248), .B(n13247), .ZN(n13249) );
  OAI211_X1 U16283 ( .C1(n19841), .C2(n19701), .A(n13250), .B(n13249), .ZN(
        P1_U2996) );
  XNOR2_X1 U16284 ( .A(n13252), .B(n13251), .ZN(n13287) );
  NAND3_X1 U16285 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n15672), .ZN(n15721) );
  NAND2_X1 U16286 ( .A1(n19829), .A2(n15721), .ZN(n15696) );
  NOR2_X1 U16287 ( .A1(n13846), .A2(n15689), .ZN(n15746) );
  NAND2_X1 U16288 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15719) );
  OAI211_X1 U16289 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n15746), .B(n15719), .ZN(n13263) );
  INV_X1 U16290 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13844) );
  AOI221_X1 U16291 ( .B1(n13844), .B2(n15720), .C1(n13075), .C2(n15720), .A(
        n15676), .ZN(n15700) );
  NAND2_X1 U16292 ( .A1(n15700), .A2(n13254), .ZN(n15717) );
  INV_X1 U16293 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20522) );
  NOR2_X1 U16294 ( .A1(n15731), .A2(n20522), .ZN(n13283) );
  MUX2_X1 U16295 ( .A(n13831), .B(n13832), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n13258) );
  INV_X1 U16296 ( .A(n13832), .ZN(n13255) );
  NAND2_X1 U16297 ( .A1(n13255), .A2(n13897), .ZN(n13648) );
  NAND2_X1 U16298 ( .A1(n13897), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13256) );
  AND2_X1 U16299 ( .A1(n13648), .A2(n13256), .ZN(n13257) );
  NAND2_X1 U16300 ( .A1(n13258), .A2(n13257), .ZN(n13259) );
  OAI21_X1 U16301 ( .B1(n13260), .B2(n13259), .A(n15748), .ZN(n19685) );
  NOR2_X1 U16302 ( .A1(n15733), .A2(n19685), .ZN(n13261) );
  AOI211_X1 U16303 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n15717), .A(
        n13283), .B(n13261), .ZN(n13262) );
  OAI211_X1 U16304 ( .C1(n13287), .C2(n15685), .A(n13263), .B(n13262), .ZN(
        P1_U3027) );
  NAND2_X1 U16305 ( .A1(n13264), .A2(n13265), .ZN(n13266) );
  XNOR2_X1 U16306 ( .A(n15947), .B(n13266), .ZN(n13273) );
  NAND2_X1 U16307 ( .A1(n16058), .A2(n15802), .ZN(n13271) );
  OAI22_X1 U16308 ( .A1(n16054), .A2(n18810), .B1(n13267), .B2(n18795), .ZN(
        n13269) );
  OAI22_X1 U16309 ( .A1(n18798), .A2(n10536), .B1(n15958), .B2(n18694), .ZN(
        n13268) );
  AOI211_X1 U16310 ( .C1(n18814), .C2(n15954), .A(n13269), .B(n13268), .ZN(
        n13270) );
  OAI211_X1 U16311 ( .C1(n13459), .C2(n19581), .A(n13271), .B(n13270), .ZN(
        n13272) );
  AOI21_X1 U16312 ( .B1(n13273), .B2(n19499), .A(n13272), .ZN(n13274) );
  INV_X1 U16313 ( .A(n13274), .ZN(P2_U2852) );
  NAND2_X1 U16314 ( .A1(n13275), .A2(n13276), .ZN(n13277) );
  AND2_X1 U16315 ( .A1(n13364), .A2(n13277), .ZN(n19740) );
  INV_X1 U16316 ( .A(n19740), .ZN(n13280) );
  NAND2_X1 U16317 ( .A1(n19840), .A2(DATAI_5_), .ZN(n13279) );
  NAND2_X1 U16318 ( .A1(n19839), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13278) );
  AND2_X1 U16319 ( .A1(n13279), .A2(n13278), .ZN(n19878) );
  OAI222_X1 U16320 ( .A1(n13280), .A2(n14209), .B1(n14213), .B2(n19878), .C1(
        n14210), .C2(n11944), .ZN(P1_U2899) );
  INV_X1 U16321 ( .A(n13275), .ZN(n13281) );
  AOI21_X1 U16322 ( .B1(n13282), .B2(n13163), .A(n13281), .ZN(n19691) );
  AOI21_X1 U16323 ( .B1(n19813), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n13283), .ZN(n13284) );
  OAI21_X1 U16324 ( .B1(n15597), .B2(n19694), .A(n13284), .ZN(n13285) );
  AOI21_X1 U16325 ( .B1(n19691), .B2(n14290), .A(n13285), .ZN(n13286) );
  OAI21_X1 U16326 ( .B1(n19637), .B2(n13287), .A(n13286), .ZN(P1_U2995) );
  XNOR2_X1 U16327 ( .A(n13288), .B(n13289), .ZN(n14963) );
  AOI22_X1 U16328 ( .A1(n18895), .A2(n13919), .B1(P2_EAX_REG_13__SCAN_IN), 
        .B2(n18893), .ZN(n13290) );
  OAI21_X1 U16329 ( .B1(n14963), .B2(n18898), .A(n13290), .ZN(P2_U2906) );
  INV_X1 U16330 ( .A(n19691), .ZN(n13313) );
  NAND2_X1 U16331 ( .A1(n19840), .A2(DATAI_4_), .ZN(n13292) );
  NAND2_X1 U16332 ( .A1(n19839), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13291) );
  AND2_X1 U16333 ( .A1(n13292), .A2(n13291), .ZN(n19874) );
  INV_X1 U16334 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19768) );
  OAI222_X1 U16335 ( .A1(n13313), .A2(n14209), .B1(n14213), .B2(n19874), .C1(
        n14210), .C2(n19768), .ZN(P1_U2900) );
  AOI22_X1 U16336 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15717), .B1(
        n15746), .B2(n12517), .ZN(n13294) );
  OAI211_X1 U16337 ( .C1(n15733), .C2(n19697), .A(n13294), .B(n13293), .ZN(
        n13295) );
  AOI21_X1 U16338 ( .B1(n13296), .B2(n19824), .A(n13295), .ZN(n13297) );
  INV_X1 U16339 ( .A(n13297), .ZN(P1_U3028) );
  INV_X1 U16340 ( .A(n18943), .ZN(n13301) );
  NOR2_X1 U16341 ( .A1(n18785), .A2(n13298), .ZN(n13300) );
  AOI21_X1 U16342 ( .B1(n13301), .B2(n13300), .A(n18779), .ZN(n13299) );
  OAI21_X1 U16343 ( .B1(n13301), .B2(n13300), .A(n13299), .ZN(n13311) );
  OAI21_X1 U16344 ( .B1(n13304), .B2(n13303), .A(n13302), .ZN(n18874) );
  INV_X1 U16345 ( .A(n18874), .ZN(n18937) );
  AOI22_X1 U16346 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n18819), .B1(n15802), .B2(
        n13517), .ZN(n13305) );
  OAI211_X1 U16347 ( .C1(n11064), .C2(n18694), .A(n11181), .B(n13305), .ZN(
        n13306) );
  AOI21_X1 U16348 ( .B1(n18669), .B2(P2_REIP_REG_4__SCAN_IN), .A(n13306), .ZN(
        n13307) );
  OAI21_X1 U16349 ( .B1(n13308), .B2(n18795), .A(n13307), .ZN(n13309) );
  AOI21_X1 U16350 ( .B1(n18937), .B2(n18814), .A(n13309), .ZN(n13310) );
  OAI211_X1 U16351 ( .C1(n13459), .C2(n13312), .A(n13311), .B(n13310), .ZN(
        P2_U2851) );
  INV_X1 U16352 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13314) );
  OAI222_X1 U16353 ( .A1(n19685), .A2(n14146), .B1(n19742), .B2(n13314), .C1(
        n13313), .C2(n14144), .ZN(P1_U2868) );
  NOR2_X1 U16354 ( .A1(n18785), .A2(n13315), .ZN(n13316) );
  XNOR2_X1 U16355 ( .A(n13316), .B(n15930), .ZN(n13328) );
  AOI22_X1 U16356 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(n18819), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n9607), .ZN(n13317) );
  OAI21_X1 U16357 ( .B1(n13318), .B2(n18795), .A(n13317), .ZN(n13327) );
  AND2_X1 U16358 ( .A1(n13320), .A2(n13319), .ZN(n13322) );
  OR2_X1 U16359 ( .A1(n13322), .A2(n13321), .ZN(n18870) );
  OAI21_X1 U16360 ( .B1(n18810), .B2(n13323), .A(n11181), .ZN(n13324) );
  AOI21_X1 U16361 ( .B1(n15802), .B2(n16016), .A(n13324), .ZN(n13325) );
  OAI21_X1 U16362 ( .B1(n18789), .B2(n18870), .A(n13325), .ZN(n13326) );
  AOI211_X1 U16363 ( .C1(n13328), .C2(n19499), .A(n13327), .B(n13326), .ZN(
        n13329) );
  INV_X1 U16364 ( .A(n13329), .ZN(P2_U2847) );
  NAND2_X1 U16365 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n15763), .ZN(n13332) );
  NOR3_X1 U16366 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .A3(n20294), .ZN(n15425) );
  NAND2_X1 U16367 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15425), .ZN(n13330) );
  OAI211_X1 U16368 ( .C1(n13332), .C2(n13331), .A(n15731), .B(n13330), .ZN(
        n13333) );
  NOR2_X1 U16369 ( .A1(n13334), .A2(n13863), .ZN(n13335) );
  XNOR2_X1 U16370 ( .A(n13335), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14219) );
  NOR2_X1 U16371 ( .A1(n14219), .A2(n15418), .ZN(n13336) );
  NAND3_X1 U16372 ( .A1(n19708), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n13337), 
        .ZN(n13338) );
  NAND2_X1 U16373 ( .A1(n15521), .A2(n13338), .ZN(n19727) );
  INV_X1 U16374 ( .A(n19727), .ZN(n13378) );
  AND2_X1 U16375 ( .A1(n9618), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13339) );
  NAND2_X1 U16376 ( .A1(n19858), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13353) );
  NAND2_X1 U16377 ( .A1(n15448), .A2(n20334), .ZN(n15417) );
  INV_X1 U16378 ( .A(n15417), .ZN(n13351) );
  NOR2_X1 U16379 ( .A1(n13353), .A2(n13351), .ZN(n13340) );
  NOR2_X1 U16380 ( .A1(n13341), .A2(n20437), .ZN(n13342) );
  NAND2_X1 U16381 ( .A1(n19708), .A2(n13342), .ZN(n19723) );
  INV_X1 U16382 ( .A(n19723), .ZN(n19696) );
  NAND2_X1 U16383 ( .A1(n19696), .A2(n9622), .ZN(n13350) );
  AND2_X1 U16384 ( .A1(n14219), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13344) );
  NAND2_X1 U16385 ( .A1(n19703), .A2(n13345), .ZN(n13349) );
  NAND2_X1 U16386 ( .A1(n19721), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13348) );
  INV_X1 U16387 ( .A(n19708), .ZN(n13346) );
  NAND2_X1 U16388 ( .A1(n13346), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n13347) );
  NAND4_X1 U16389 ( .A1(n13350), .A2(n13349), .A3(n13348), .A4(n13347), .ZN(
        n13359) );
  AND2_X1 U16390 ( .A1(n13352), .A2(n13351), .ZN(n13355) );
  INV_X1 U16391 ( .A(n13353), .ZN(n13354) );
  NOR2_X1 U16392 ( .A1(n13355), .A2(n13354), .ZN(n13356) );
  OAI22_X1 U16393 ( .A1(n19709), .A2(P1_REIP_REG_1__SCAN_IN), .B1(n19715), 
        .B2(n13002), .ZN(n13358) );
  AOI211_X1 U16394 ( .C1(n19700), .C2(n13360), .A(n13359), .B(n13358), .ZN(
        n13361) );
  OAI21_X1 U16395 ( .B1(n13378), .B2(n13362), .A(n13361), .ZN(P1_U2839) );
  INV_X1 U16396 ( .A(n13363), .ZN(n13365) );
  XNOR2_X1 U16397 ( .A(n13365), .B(n13364), .ZN(n19664) );
  INV_X1 U16398 ( .A(n19664), .ZN(n13381) );
  INV_X1 U16399 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20661) );
  NAND2_X1 U16400 ( .A1(n13838), .A2(n20661), .ZN(n13367) );
  NAND2_X1 U16401 ( .A1(n13821), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13366) );
  NAND3_X1 U16402 ( .A1(n13367), .A2(n13832), .A3(n13366), .ZN(n13368) );
  OAI21_X1 U16403 ( .B1(n13829), .B2(P1_EBX_REG_5__SCAN_IN), .A(n13368), .ZN(
        n15747) );
  MUX2_X1 U16404 ( .A(n13831), .B(n13832), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n13370) );
  NAND2_X1 U16405 ( .A1(n13897), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13369) );
  INV_X1 U16406 ( .A(n13394), .ZN(n13371) );
  XNOR2_X1 U16407 ( .A(n15750), .B(n13371), .ZN(n19667) );
  AOI22_X1 U16408 ( .A1(n19738), .A2(n19667), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14134), .ZN(n13372) );
  OAI21_X1 U16409 ( .B1(n13381), .B2(n14144), .A(n13372), .ZN(P1_U2866) );
  NAND2_X1 U16410 ( .A1(n19709), .A2(n19708), .ZN(n15468) );
  OAI22_X1 U16411 ( .A1(n19718), .A2(n19822), .B1(n13373), .B2(n19715), .ZN(
        n13374) );
  AOI21_X1 U16412 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(n15468), .A(n13374), .ZN(
        n13377) );
  NAND2_X1 U16413 ( .A1(n15525), .A2(n19731), .ZN(n13375) );
  AOI22_X1 U16414 ( .A1(n13375), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n11860), .B2(n19696), .ZN(n13376) );
  OAI211_X1 U16415 ( .C1(n13378), .C2(n19821), .A(n13377), .B(n13376), .ZN(
        P1_U2840) );
  NAND2_X1 U16416 ( .A1(n19840), .A2(DATAI_6_), .ZN(n13380) );
  NAND2_X1 U16417 ( .A1(n19839), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13379) );
  AND2_X1 U16418 ( .A1(n13380), .A2(n13379), .ZN(n19882) );
  OAI222_X1 U16419 ( .A1(n14209), .A2(n13381), .B1(n14213), .B2(n19882), .C1(
        n14210), .C2(n11961), .ZN(P1_U2898) );
  NOR2_X1 U16420 ( .A1(n13382), .A2(n15448), .ZN(n13383) );
  INV_X2 U16421 ( .A(n19799), .ZN(n19804) );
  OR2_X1 U16422 ( .A1(n19804), .A2(n19858), .ZN(n13412) );
  INV_X1 U16423 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n19748) );
  NOR2_X2 U16424 ( .A1(n19804), .A2(n11733), .ZN(n19792) );
  INV_X1 U16425 ( .A(n19792), .ZN(n13387) );
  INV_X1 U16426 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13385) );
  NOR2_X1 U16427 ( .A1(n19840), .A2(n13385), .ZN(n13386) );
  AOI21_X1 U16428 ( .B1(DATAI_15_), .B2(n19840), .A(n13386), .ZN(n14204) );
  INV_X1 U16429 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n19749) );
  OAI222_X1 U16430 ( .A1(n13412), .A2(n19748), .B1(n13387), .B2(n14204), .C1(
        n19799), .C2(n19749), .ZN(P1_U2967) );
  AOI22_X1 U16431 ( .A1(n19809), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n19804), .ZN(n13390) );
  INV_X1 U16432 ( .A(DATAI_9_), .ZN(n13389) );
  NAND2_X1 U16433 ( .A1(n19839), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13388) );
  OAI21_X1 U16434 ( .B1(n19839), .B2(n13389), .A(n13388), .ZN(n14162) );
  NAND2_X1 U16435 ( .A1(n19792), .A2(n14162), .ZN(n19797) );
  NAND2_X1 U16436 ( .A1(n13390), .A2(n19797), .ZN(P1_U2946) );
  OAI21_X1 U16437 ( .B1(n13393), .B2(n13392), .A(n13391), .ZN(n13485) );
  INV_X1 U16438 ( .A(n13829), .ZN(n13395) );
  INV_X1 U16439 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13396) );
  NAND2_X1 U16440 ( .A1(n13395), .A2(n13396), .ZN(n13400) );
  NAND2_X1 U16441 ( .A1(n13838), .A2(n13396), .ZN(n13398) );
  NAND2_X1 U16442 ( .A1(n13821), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13397) );
  NAND3_X1 U16443 ( .A1(n13398), .A2(n13832), .A3(n13397), .ZN(n13399) );
  NOR2_X1 U16444 ( .A1(n13402), .A2(n13401), .ZN(n13403) );
  OR2_X1 U16445 ( .A1(n13500), .A2(n13403), .ZN(n15732) );
  INV_X1 U16446 ( .A(n15732), .ZN(n13404) );
  AOI22_X1 U16447 ( .A1(n19738), .A2(n13404), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n14134), .ZN(n13405) );
  OAI21_X1 U16448 ( .B1(n13485), .B2(n14136), .A(n13405), .ZN(P1_U2865) );
  XNOR2_X1 U16449 ( .A(n13406), .B(n18838), .ZN(n13411) );
  INV_X1 U16450 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n13409) );
  INV_X1 U16451 ( .A(n14945), .ZN(n13407) );
  AOI21_X1 U16452 ( .B1(n13408), .B2(n15873), .A(n13407), .ZN(n14961) );
  INV_X1 U16453 ( .A(n14961), .ZN(n13529) );
  MUX2_X1 U16454 ( .A(n13409), .B(n13529), .S(n18859), .Z(n13410) );
  OAI21_X1 U16455 ( .B1(n13411), .B2(n18865), .A(n13410), .ZN(P2_U2874) );
  INV_X2 U16456 ( .A(n13412), .ZN(n19809) );
  AOI22_X1 U16457 ( .A1(n19809), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n19804), .ZN(n13413) );
  INV_X1 U16458 ( .A(n19860), .ZN(n14193) );
  NAND2_X1 U16459 ( .A1(n19792), .A2(n14193), .ZN(n13434) );
  NAND2_X1 U16460 ( .A1(n13413), .A2(n13434), .ZN(P1_U2938) );
  AOI22_X1 U16461 ( .A1(n19809), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n19804), .ZN(n13416) );
  NAND2_X1 U16462 ( .A1(n19840), .A2(DATAI_7_), .ZN(n13415) );
  NAND2_X1 U16463 ( .A1(n19839), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13414) );
  AND2_X1 U16464 ( .A1(n13415), .A2(n13414), .ZN(n19890) );
  INV_X1 U16465 ( .A(n19890), .ZN(n14168) );
  NAND2_X1 U16466 ( .A1(n19792), .A2(n14168), .ZN(n13419) );
  NAND2_X1 U16467 ( .A1(n13416), .A2(n13419), .ZN(P1_U2944) );
  AOI22_X1 U16468 ( .A1(n19809), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n19804), .ZN(n13417) );
  INV_X1 U16469 ( .A(n19865), .ZN(n14189) );
  NAND2_X1 U16470 ( .A1(n19792), .A2(n14189), .ZN(n13436) );
  NAND2_X1 U16471 ( .A1(n13417), .A2(n13436), .ZN(P1_U2954) );
  AOI22_X1 U16472 ( .A1(n19809), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n19804), .ZN(n13418) );
  INV_X1 U16473 ( .A(n19851), .ZN(n14199) );
  NAND2_X1 U16474 ( .A1(n19792), .A2(n14199), .ZN(n13427) );
  NAND2_X1 U16475 ( .A1(n13418), .A2(n13427), .ZN(P1_U2937) );
  AOI22_X1 U16476 ( .A1(n19809), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n19804), .ZN(n13420) );
  NAND2_X1 U16477 ( .A1(n13420), .A2(n13419), .ZN(P1_U2959) );
  AOI22_X1 U16478 ( .A1(n19809), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n19804), .ZN(n13421) );
  INV_X1 U16479 ( .A(n19874), .ZN(n14182) );
  NAND2_X1 U16480 ( .A1(n19792), .A2(n14182), .ZN(n13423) );
  NAND2_X1 U16481 ( .A1(n13421), .A2(n13423), .ZN(P1_U2941) );
  AOI22_X1 U16482 ( .A1(n19809), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n19804), .ZN(n13422) );
  INV_X1 U16483 ( .A(n19870), .ZN(n14185) );
  NAND2_X1 U16484 ( .A1(n19792), .A2(n14185), .ZN(n13425) );
  NAND2_X1 U16485 ( .A1(n13422), .A2(n13425), .ZN(P1_U2955) );
  AOI22_X1 U16486 ( .A1(n19809), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n19804), .ZN(n13424) );
  NAND2_X1 U16487 ( .A1(n13424), .A2(n13423), .ZN(P1_U2956) );
  AOI22_X1 U16488 ( .A1(n19809), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n19804), .ZN(n13426) );
  NAND2_X1 U16489 ( .A1(n13426), .A2(n13425), .ZN(P1_U2940) );
  AOI22_X1 U16490 ( .A1(n19809), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n19804), .ZN(n13428) );
  NAND2_X1 U16491 ( .A1(n13428), .A2(n13427), .ZN(P1_U2952) );
  AOI22_X1 U16492 ( .A1(n19809), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n19804), .ZN(n13429) );
  INV_X1 U16493 ( .A(n19882), .ZN(n14172) );
  NAND2_X1 U16494 ( .A1(n19792), .A2(n14172), .ZN(n13438) );
  NAND2_X1 U16495 ( .A1(n13429), .A2(n13438), .ZN(P1_U2943) );
  AOI22_X1 U16496 ( .A1(n19809), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n19804), .ZN(n13431) );
  INV_X1 U16497 ( .A(n19878), .ZN(n13430) );
  NAND2_X1 U16498 ( .A1(n19792), .A2(n13430), .ZN(n13432) );
  NAND2_X1 U16499 ( .A1(n13431), .A2(n13432), .ZN(P1_U2942) );
  AOI22_X1 U16500 ( .A1(n19809), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n19804), .ZN(n13433) );
  NAND2_X1 U16501 ( .A1(n13433), .A2(n13432), .ZN(P1_U2957) );
  AOI22_X1 U16502 ( .A1(n19809), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n19804), .ZN(n13435) );
  NAND2_X1 U16503 ( .A1(n13435), .A2(n13434), .ZN(P1_U2953) );
  AOI22_X1 U16504 ( .A1(n19809), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n19804), .ZN(n13437) );
  NAND2_X1 U16505 ( .A1(n13437), .A2(n13436), .ZN(P1_U2939) );
  AOI22_X1 U16506 ( .A1(n19809), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n19804), .ZN(n13439) );
  NAND2_X1 U16507 ( .A1(n13439), .A2(n13438), .ZN(P1_U2958) );
  INV_X1 U16508 ( .A(n13440), .ZN(n13446) );
  NAND2_X1 U16509 ( .A1(n13442), .A2(n13441), .ZN(n13445) );
  INV_X1 U16510 ( .A(n13443), .ZN(n13444) );
  NAND2_X1 U16511 ( .A1(n13445), .A2(n13444), .ZN(n18721) );
  OAI222_X1 U16512 ( .A1(n13483), .A2(n13446), .B1(n18721), .B2(n18898), .C1(
        n10979), .C2(n14596), .ZN(P2_U2905) );
  INV_X1 U16513 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n19764) );
  OAI222_X1 U16514 ( .A1(n13485), .A2(n14209), .B1(n14213), .B2(n19890), .C1(
        n14210), .C2(n19764), .ZN(P1_U2897) );
  NOR2_X1 U16515 ( .A1(n18785), .A2(n13447), .ZN(n13460) );
  INV_X1 U16516 ( .A(n13460), .ZN(n13448) );
  AOI221_X1 U16517 ( .B1(n13450), .B2(n13460), .C1(n13449), .C2(n13448), .A(
        n18779), .ZN(n13451) );
  INV_X1 U16518 ( .A(n13451), .ZN(n13458) );
  AOI22_X1 U16519 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n9607), .B1(
        P2_EBX_REG_2__SCAN_IN), .B2(n18819), .ZN(n13454) );
  AOI22_X1 U16520 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n18669), .B1(n13452), 
        .B2(n18818), .ZN(n13453) );
  OAI211_X1 U16521 ( .C1(n13455), .C2(n18812), .A(n13454), .B(n13453), .ZN(
        n13456) );
  AOI21_X1 U16522 ( .B1(n18814), .B2(n15014), .A(n13456), .ZN(n13457) );
  OAI211_X1 U16523 ( .C1(n19592), .C2(n13459), .A(n13458), .B(n13457), .ZN(
        P2_U2853) );
  OAI21_X1 U16524 ( .B1(n18831), .B2(n13461), .A(n13460), .ZN(n14991) );
  NAND2_X1 U16525 ( .A1(n18819), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n13470) );
  NAND2_X1 U16526 ( .A1(n15802), .A2(n19601), .ZN(n13469) );
  AOI22_X1 U16527 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18669), .B1(n13462), 
        .B2(n18818), .ZN(n13464) );
  NOR2_X1 U16528 ( .A1(n18779), .A2(n13264), .ZN(n18826) );
  NAND2_X1 U16529 ( .A1(n18826), .A2(n13465), .ZN(n13463) );
  OAI211_X1 U16530 ( .C1(n18694), .C2(n13465), .A(n13464), .B(n13463), .ZN(
        n13466) );
  INV_X1 U16531 ( .A(n13466), .ZN(n13468) );
  NAND2_X1 U16532 ( .A1(n14990), .A2(n18814), .ZN(n13467) );
  NAND4_X1 U16533 ( .A1(n13470), .A2(n13469), .A3(n13468), .A4(n13467), .ZN(
        n13471) );
  AOI21_X1 U16534 ( .B1(n19590), .B2(n18825), .A(n13471), .ZN(n13472) );
  OAI21_X1 U16535 ( .B1(n14991), .B2(n18779), .A(n13472), .ZN(P2_U2854) );
  INV_X1 U16536 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n13480) );
  INV_X1 U16537 ( .A(n13473), .ZN(n18840) );
  OAI211_X1 U16538 ( .C1(n18840), .C2(n13475), .A(n18871), .B(n13474), .ZN(
        n13479) );
  OR2_X1 U16539 ( .A1(n14946), .A2(n13476), .ZN(n13477) );
  AND2_X1 U16540 ( .A1(n14727), .A2(n13477), .ZN(n18708) );
  NAND2_X1 U16541 ( .A1(n18708), .A2(n18859), .ZN(n13478) );
  OAI211_X1 U16542 ( .C1(n18859), .C2(n13480), .A(n13479), .B(n13478), .ZN(
        P2_U2872) );
  OAI21_X1 U16543 ( .B1(n13481), .B2(n13443), .A(n14923), .ZN(n18709) );
  OAI222_X1 U16544 ( .A1(n18709), .A2(n18898), .B1(n13483), .B2(n13482), .C1(
        n12707), .C2(n14596), .ZN(P2_U2904) );
  INV_X1 U16545 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20529) );
  NAND2_X1 U16546 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n13484) );
  NAND3_X1 U16547 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n19688) );
  NOR2_X1 U16548 ( .A1(n20522), .A2(n19688), .ZN(n13577) );
  OAI21_X1 U16549 ( .B1(n19709), .B2(n13577), .A(n19708), .ZN(n19690) );
  AOI21_X1 U16550 ( .B1(n13484), .B2(n15468), .A(n19690), .ZN(n19673) );
  INV_X1 U16551 ( .A(n13485), .ZN(n15587) );
  NAND2_X1 U16552 ( .A1(n15587), .A2(n19663), .ZN(n13492) );
  NAND2_X1 U16553 ( .A1(n19708), .A2(n13486), .ZN(n19683) );
  NAND2_X1 U16554 ( .A1(n19721), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13487) );
  OAI211_X1 U16555 ( .C1(n19731), .C2(n15590), .A(n19683), .B(n13487), .ZN(
        n13490) );
  NAND2_X1 U16556 ( .A1(n14015), .A2(n13577), .ZN(n19674) );
  NAND3_X1 U16557 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n20529), .ZN(n13488) );
  OAI22_X1 U16558 ( .A1(n19718), .A2(n15732), .B1(n19674), .B2(n13488), .ZN(
        n13489) );
  AOI211_X1 U16559 ( .C1(n19695), .C2(P1_EBX_REG_7__SCAN_IN), .A(n13490), .B(
        n13489), .ZN(n13491) );
  OAI211_X1 U16560 ( .C1(n20529), .C2(n19673), .A(n13492), .B(n13491), .ZN(
        P1_U2833) );
  INV_X1 U16561 ( .A(n13493), .ZN(n13545) );
  AOI21_X1 U16562 ( .B1(n13494), .B2(n13391), .A(n13493), .ZN(n13542) );
  INV_X1 U16563 ( .A(n13542), .ZN(n13524) );
  INV_X1 U16564 ( .A(n14213), .ZN(n14207) );
  MUX2_X1 U16565 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n19839), .Z(
        n19781) );
  AOI22_X1 U16566 ( .A1(n14207), .A2(n19781), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14206), .ZN(n13495) );
  OAI21_X1 U16567 ( .B1(n13524), .B2(n14209), .A(n13495), .ZN(P1_U2896) );
  NAND3_X1 U16568 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n13503) );
  NOR3_X1 U16569 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n13503), .A3(n19674), .ZN(
        n13510) );
  MUX2_X1 U16570 ( .A(n13831), .B(n13832), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n13498) );
  NAND2_X1 U16571 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n13897), .ZN(
        n13496) );
  AND2_X1 U16572 ( .A1(n13648), .A2(n13496), .ZN(n13497) );
  NAND2_X1 U16573 ( .A1(n13498), .A2(n13497), .ZN(n13499) );
  OR2_X1 U16574 ( .A1(n13500), .A2(n13499), .ZN(n13501) );
  NAND2_X1 U16575 ( .A1(n15708), .A2(n13501), .ZN(n15725) );
  OAI22_X1 U16576 ( .A1(n13502), .A2(n15525), .B1(n19718), .B2(n15725), .ZN(
        n13509) );
  INV_X1 U16577 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13507) );
  INV_X1 U16578 ( .A(n13540), .ZN(n13505) );
  INV_X1 U16579 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20530) );
  NOR2_X1 U16580 ( .A1(n20530), .A2(n13503), .ZN(n13576) );
  NAND3_X1 U16581 ( .A1(n13577), .A2(n13576), .A3(n19708), .ZN(n13574) );
  NAND2_X1 U16582 ( .A1(n15468), .A2(n13574), .ZN(n19654) );
  OAI21_X1 U16583 ( .B1(n20530), .B2(n19654), .A(n19683), .ZN(n13504) );
  AOI21_X1 U16584 ( .B1(n19703), .B2(n13505), .A(n13504), .ZN(n13506) );
  OAI21_X1 U16585 ( .B1(n19715), .B2(n13507), .A(n13506), .ZN(n13508) );
  NOR3_X1 U16586 ( .A1(n13510), .A2(n13509), .A3(n13508), .ZN(n13511) );
  OAI21_X1 U16587 ( .B1(n13524), .B2(n15521), .A(n13511), .ZN(P1_U2832) );
  XNOR2_X1 U16588 ( .A(n13512), .B(n16042), .ZN(n18940) );
  INV_X1 U16589 ( .A(n18940), .ZN(n13523) );
  NAND2_X1 U16590 ( .A1(n15951), .A2(n15952), .ZN(n13514) );
  NAND2_X1 U16591 ( .A1(n13514), .A2(n13513), .ZN(n13515) );
  XOR2_X1 U16592 ( .A(n13516), .B(n13515), .Z(n18935) );
  NAND2_X1 U16593 ( .A1(n18935), .A2(n16063), .ZN(n13522) );
  NAND2_X1 U16594 ( .A1(n16036), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13519) );
  AOI22_X1 U16595 ( .A1(n16057), .A2(n13517), .B1(n18933), .B2(
        P2_REIP_REG_4__SCAN_IN), .ZN(n13518) );
  OAI211_X1 U16596 ( .C1(n18874), .C2(n16055), .A(n13519), .B(n13518), .ZN(
        n13520) );
  AOI21_X1 U16597 ( .B1(n16039), .B2(n16042), .A(n13520), .ZN(n13521) );
  OAI211_X1 U16598 ( .C1(n13523), .C2(n16060), .A(n13522), .B(n13521), .ZN(
        P2_U3042) );
  OAI222_X1 U16599 ( .A1(n13524), .A2(n14136), .B1(n19742), .B2(n13507), .C1(
        n15725), .C2(n14146), .ZN(P1_U2864) );
  NAND2_X1 U16600 ( .A1(n19499), .A2(n13264), .ZN(n18830) );
  AOI211_X1 U16601 ( .C1(n14748), .C2(n13525), .A(n18715), .B(n18830), .ZN(
        n13526) );
  INV_X1 U16602 ( .A(n13526), .ZN(n13535) );
  INV_X1 U16603 ( .A(n18826), .ZN(n13528) );
  INV_X1 U16604 ( .A(n14748), .ZN(n13527) );
  OAI22_X1 U16605 ( .A1(n13529), .A2(n18789), .B1(n13528), .B2(n13527), .ZN(
        n13533) );
  AOI22_X1 U16606 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n9607), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n18669), .ZN(n13530) );
  OAI211_X1 U16607 ( .C1(n13531), .C2(n18795), .A(n13530), .B(n11181), .ZN(
        n13532) );
  AOI211_X1 U16608 ( .C1(P2_EBX_REG_13__SCAN_IN), .C2(n18819), .A(n13533), .B(
        n13532), .ZN(n13534) );
  OAI211_X1 U16609 ( .C1(n14963), .C2(n18812), .A(n13535), .B(n13534), .ZN(
        P2_U2842) );
  XNOR2_X1 U16610 ( .A(n13536), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13537) );
  XNOR2_X1 U16611 ( .A(n13538), .B(n13537), .ZN(n15724) );
  AOI22_X1 U16612 ( .A1(n19813), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19819), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13539) );
  OAI21_X1 U16613 ( .B1(n15597), .B2(n13540), .A(n13539), .ZN(n13541) );
  AOI21_X1 U16614 ( .B1(n13542), .B2(n14290), .A(n13541), .ZN(n13543) );
  OAI21_X1 U16615 ( .B1(n15724), .B2(n19637), .A(n13543), .ZN(P1_U2991) );
  AND2_X1 U16616 ( .A1(n13545), .A2(n13544), .ZN(n13547) );
  OR2_X1 U16617 ( .A1(n13547), .A2(n13546), .ZN(n19656) );
  AOI22_X1 U16618 ( .A1(n14207), .A2(n14162), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14206), .ZN(n13548) );
  OAI21_X1 U16619 ( .B1(n19656), .B2(n14209), .A(n13548), .ZN(P1_U2895) );
  AND2_X1 U16620 ( .A1(n14729), .A2(n13549), .ZN(n13551) );
  OR2_X1 U16621 ( .A1(n13551), .A2(n13550), .ZN(n18683) );
  AOI21_X1 U16622 ( .B1(n13553), .B2(n18832), .A(n13552), .ZN(n13598) );
  NAND2_X1 U16623 ( .A1(n13598), .A2(n18871), .ZN(n13555) );
  NAND2_X1 U16624 ( .A1(n18875), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13554) );
  OAI211_X1 U16625 ( .C1(n18683), .C2(n18875), .A(n13555), .B(n13554), .ZN(
        P2_U2870) );
  AOI22_X1 U16626 ( .A1(n18938), .A2(n13556), .B1(n18934), .B2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13559) );
  OAI22_X1 U16627 ( .A1(n11057), .A2(n16010), .B1(n18944), .B2(n18787), .ZN(
        n13557) );
  INV_X1 U16628 ( .A(n13557), .ZN(n13558) );
  OAI211_X1 U16629 ( .C1(n13560), .C2(n15942), .A(n13559), .B(n13558), .ZN(
        n13561) );
  INV_X1 U16630 ( .A(n13561), .ZN(n13562) );
  OAI21_X1 U16631 ( .B1(n13563), .B2(n15941), .A(n13562), .ZN(P2_U3008) );
  INV_X1 U16632 ( .A(n13621), .ZN(n13564) );
  OAI21_X1 U16633 ( .B1(n13546), .B2(n13565), .A(n13564), .ZN(n14349) );
  INV_X1 U16634 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n19736) );
  NAND2_X1 U16635 ( .A1(n13838), .A2(n19736), .ZN(n13567) );
  NAND2_X1 U16636 ( .A1(n13821), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13566) );
  NAND3_X1 U16637 ( .A1(n13567), .A2(n13832), .A3(n13566), .ZN(n13568) );
  OAI21_X1 U16638 ( .B1(n13829), .B2(P1_EBX_REG_9__SCAN_IN), .A(n13568), .ZN(
        n15707) );
  OR2_X1 U16639 ( .A1(n13831), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n13572) );
  INV_X1 U16640 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14341) );
  NAND2_X1 U16641 ( .A1(n13832), .A2(n14341), .ZN(n13570) );
  INV_X1 U16642 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13579) );
  NAND2_X1 U16643 ( .A1(n13838), .A2(n13579), .ZN(n13569) );
  NAND3_X1 U16644 ( .A1(n13570), .A2(n13821), .A3(n13569), .ZN(n13571) );
  NAND2_X1 U16645 ( .A1(n13572), .A2(n13571), .ZN(n13626) );
  XNOR2_X1 U16646 ( .A(n15710), .B(n13626), .ZN(n15699) );
  AOI22_X1 U16647 ( .A1(n19738), .A2(n15699), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14134), .ZN(n13573) );
  OAI21_X1 U16648 ( .B1(n14349), .B2(n14136), .A(n13573), .ZN(P1_U2862) );
  INV_X1 U16649 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20534) );
  NAND2_X1 U16650 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n15515) );
  OAI21_X1 U16651 ( .B1(n15515), .B2(n13574), .A(n15468), .ZN(n15523) );
  AOI22_X1 U16652 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19721), .B1(
        n19700), .B2(n15699), .ZN(n13575) );
  OAI211_X1 U16653 ( .C1(n20534), .C2(n15523), .A(n13575), .B(n19683), .ZN(
        n13582) );
  NAND2_X1 U16654 ( .A1(n13577), .A2(n13576), .ZN(n13642) );
  NOR2_X1 U16655 ( .A1(n19709), .A2(n13642), .ZN(n19653) );
  NAND2_X1 U16656 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19653), .ZN(n13578) );
  NOR2_X1 U16657 ( .A1(n13578), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n13581) );
  OAI22_X1 U16658 ( .A1(n19731), .A2(n14345), .B1(n19715), .B2(n13579), .ZN(
        n13580) );
  NOR3_X1 U16659 ( .A1(n13582), .A2(n13581), .A3(n13580), .ZN(n13583) );
  OAI21_X1 U16660 ( .B1(n14349), .B2(n15521), .A(n13583), .ZN(P1_U2830) );
  MUX2_X1 U16661 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n19839), .Z(
        n19783) );
  AOI22_X1 U16662 ( .A1(n14207), .A2(n19783), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14206), .ZN(n13584) );
  OAI21_X1 U16663 ( .B1(n14349), .B2(n14209), .A(n13584), .ZN(P1_U2894) );
  NAND2_X1 U16664 ( .A1(n9701), .A2(n13585), .ZN(n13586) );
  XNOR2_X1 U16665 ( .A(n13587), .B(n13586), .ZN(n15713) );
  NAND2_X1 U16666 ( .A1(n15713), .A2(n19817), .ZN(n13591) );
  INV_X1 U16667 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n13588) );
  NOR2_X1 U16668 ( .A1(n15731), .A2(n13588), .ZN(n15711) );
  AND2_X1 U16669 ( .A1(n19813), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13589) );
  AOI211_X1 U16670 ( .C1(n19657), .C2(n15600), .A(n15711), .B(n13589), .ZN(
        n13590) );
  OAI211_X1 U16671 ( .C1(n19841), .C2(n19656), .A(n13591), .B(n13590), .ZN(
        P1_U2990) );
  OAI21_X1 U16672 ( .B1(n13593), .B2(n13592), .A(n14899), .ZN(n18689) );
  AOI22_X1 U16673 ( .A1(n18882), .A2(BUF1_REG_17__SCAN_IN), .B1(n18881), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n13596) );
  AOI22_X1 U16674 ( .A1(n18880), .A2(n13594), .B1(n18893), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n13595) );
  OAI211_X1 U16675 ( .C1(n14585), .C2(n18689), .A(n13596), .B(n13595), .ZN(
        n13597) );
  AOI21_X1 U16676 ( .B1(n13598), .B2(n18885), .A(n13597), .ZN(n13599) );
  INV_X1 U16677 ( .A(n13599), .ZN(P2_U2902) );
  NAND2_X1 U16678 ( .A1(n13600), .A2(n9674), .ZN(n13601) );
  XNOR2_X1 U16679 ( .A(n13601), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16032) );
  INV_X1 U16680 ( .A(n16032), .ZN(n13610) );
  INV_X1 U16681 ( .A(n15918), .ZN(n13603) );
  NAND2_X1 U16682 ( .A1(n13603), .A2(n15919), .ZN(n13604) );
  XNOR2_X1 U16683 ( .A(n13602), .B(n13604), .ZN(n16026) );
  OAI22_X1 U16684 ( .A1(n15957), .A2(n13605), .B1(n19532), .B2(n11181), .ZN(
        n13608) );
  INV_X1 U16685 ( .A(n18770), .ZN(n13606) );
  OAI22_X1 U16686 ( .A1(n15859), .A2(n18774), .B1(n18944), .B2(n13606), .ZN(
        n13607) );
  AOI211_X1 U16687 ( .C1(n16026), .C2(n18936), .A(n13608), .B(n13607), .ZN(
        n13609) );
  OAI21_X1 U16688 ( .B1(n13610), .B2(n15941), .A(n13609), .ZN(P2_U3007) );
  INV_X1 U16689 ( .A(n13611), .ZN(n15824) );
  OAI21_X1 U16690 ( .B1(n15824), .B2(n10126), .A(n13612), .ZN(n13637) );
  XNOR2_X1 U16691 ( .A(n13614), .B(n13613), .ZN(n14879) );
  INV_X1 U16692 ( .A(n14879), .ZN(n13617) );
  INV_X1 U16693 ( .A(n18880), .ZN(n14597) );
  OAI22_X1 U16694 ( .A1(n14597), .A2(n18966), .B1(n14596), .B2(n13615), .ZN(
        n13616) );
  AOI21_X1 U16695 ( .B1(n18884), .B2(n13617), .A(n13616), .ZN(n13619) );
  AOI22_X1 U16696 ( .A1(n18882), .A2(BUF1_REG_19__SCAN_IN), .B1(n18881), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n13618) );
  OAI211_X1 U16697 ( .C1(n13637), .C2(n14601), .A(n13619), .B(n13618), .ZN(
        P2_U2900) );
  OR2_X1 U16698 ( .A1(n13621), .A2(n13620), .ZN(n13622) );
  NAND2_X1 U16699 ( .A1(n14065), .A2(n13622), .ZN(n14067) );
  XNOR2_X1 U16700 ( .A(n14067), .B(n14064), .ZN(n15579) );
  INV_X1 U16701 ( .A(n15579), .ZN(n13633) );
  INV_X1 U16702 ( .A(n15710), .ZN(n13625) );
  MUX2_X1 U16703 ( .A(n13829), .B(n13821), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13624) );
  OR2_X1 U16704 ( .A1(n13898), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13623) );
  AND2_X1 U16705 ( .A1(n13624), .A2(n13623), .ZN(n13627) );
  AOI21_X1 U16706 ( .B1(n13625), .B2(n13626), .A(n13627), .ZN(n13629) );
  NAND2_X1 U16707 ( .A1(n13627), .A2(n13626), .ZN(n13628) );
  NOR2_X1 U16708 ( .A1(n13629), .A2(n9733), .ZN(n15687) );
  AOI22_X1 U16709 ( .A1(n19738), .A2(n15687), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n14134), .ZN(n13630) );
  OAI21_X1 U16710 ( .B1(n13633), .B2(n14136), .A(n13630), .ZN(P1_U2861) );
  MUX2_X1 U16711 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n19839), .Z(
        n19785) );
  INV_X1 U16712 ( .A(n19785), .ZN(n13632) );
  OAI222_X1 U16713 ( .A1(n13633), .A2(n14209), .B1(n14213), .B2(n13632), .C1(
        n13631), .C2(n14210), .ZN(P1_U2893) );
  OAI21_X1 U16714 ( .B1(n14898), .B2(n13634), .A(n14496), .ZN(n14880) );
  MUX2_X1 U16715 ( .A(n13635), .B(n14880), .S(n18859), .Z(n13636) );
  OAI21_X1 U16716 ( .B1(n13637), .B2(n18865), .A(n13636), .ZN(P2_U2868) );
  AOI21_X1 U16717 ( .B1(n13641), .B2(n13638), .A(n13640), .ZN(n14322) );
  INV_X1 U16718 ( .A(n14322), .ZN(n13668) );
  INV_X1 U16719 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20540) );
  INV_X1 U16720 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20538) );
  INV_X1 U16721 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20536) );
  NOR4_X1 U16722 ( .A1(n20538), .A2(n20536), .A3(n13642), .A4(n15515), .ZN(
        n14074) );
  NAND2_X1 U16723 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n14074), .ZN(n13643) );
  NOR2_X1 U16724 ( .A1(n20540), .A2(n13643), .ZN(n14014) );
  NAND2_X1 U16725 ( .A1(n14014), .A2(n19708), .ZN(n13989) );
  NAND2_X1 U16726 ( .A1(n15468), .A2(n13989), .ZN(n14054) );
  AOI221_X1 U16727 ( .B1(n19709), .B2(n20540), .C1(n13643), .C2(n20540), .A(
        n14054), .ZN(n13663) );
  INV_X1 U16728 ( .A(n14320), .ZN(n13644) );
  NAND2_X1 U16729 ( .A1(n19703), .A2(n13644), .ZN(n13646) );
  NAND2_X1 U16730 ( .A1(n19721), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13645) );
  NAND3_X1 U16731 ( .A1(n13646), .A2(n13645), .A3(n19683), .ZN(n13662) );
  MUX2_X1 U16732 ( .A(n13831), .B(n13832), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n13650) );
  NAND2_X1 U16733 ( .A1(n13897), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13647) );
  AND2_X1 U16734 ( .A1(n13648), .A2(n13647), .ZN(n13649) );
  NAND2_X1 U16735 ( .A1(n13650), .A2(n13649), .ZN(n14137) );
  MUX2_X1 U16736 ( .A(n13829), .B(n13821), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n13652) );
  OR2_X1 U16737 ( .A1(n13898), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13651) );
  NAND2_X1 U16738 ( .A1(n13652), .A2(n13651), .ZN(n14072) );
  INV_X1 U16739 ( .A(n14072), .ZN(n13653) );
  OR2_X1 U16740 ( .A1(n13831), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n13657) );
  NAND2_X1 U16741 ( .A1(n13832), .A2(n14437), .ZN(n13655) );
  INV_X1 U16742 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n13660) );
  NAND2_X1 U16743 ( .A1(n13838), .A2(n13660), .ZN(n13654) );
  NAND3_X1 U16744 ( .A1(n13655), .A2(n13821), .A3(n13654), .ZN(n13656) );
  NAND2_X1 U16745 ( .A1(n14069), .A2(n13658), .ZN(n13659) );
  NAND2_X1 U16746 ( .A1(n14057), .A2(n13659), .ZN(n14435) );
  OAI22_X1 U16747 ( .A1(n19718), .A2(n14435), .B1(n13660), .B2(n19715), .ZN(
        n13661) );
  NOR3_X1 U16748 ( .A1(n13663), .A2(n13662), .A3(n13661), .ZN(n13664) );
  OAI21_X1 U16749 ( .B1(n13668), .B2(n15521), .A(n13664), .ZN(P1_U2826) );
  INV_X1 U16750 ( .A(n14435), .ZN(n13665) );
  AOI22_X1 U16751 ( .A1(n13665), .A2(n19738), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n14134), .ZN(n13666) );
  OAI21_X1 U16752 ( .B1(n13668), .B2(n14144), .A(n13666), .ZN(P1_U2858) );
  MUX2_X1 U16753 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n19839), .Z(
        n19791) );
  AOI22_X1 U16754 ( .A1(n14207), .A2(n19791), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14206), .ZN(n13667) );
  OAI21_X1 U16755 ( .B1(n13668), .B2(n14209), .A(n13667), .ZN(P1_U2890) );
  OAI21_X1 U16756 ( .B1(n9654), .B2(n13670), .A(n13669), .ZN(n14557) );
  NAND2_X1 U16757 ( .A1(n18880), .A2(n13671), .ZN(n13672) );
  OAI21_X1 U16758 ( .B1(n14596), .B2(n13673), .A(n13672), .ZN(n13678) );
  INV_X1 U16759 ( .A(n18882), .ZN(n13676) );
  INV_X1 U16760 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n14176) );
  INV_X1 U16761 ( .A(n18881), .ZN(n13675) );
  INV_X1 U16762 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n13674) );
  OAI22_X1 U16763 ( .A1(n13676), .A2(n14176), .B1(n13675), .B2(n13674), .ZN(
        n13677) );
  AOI211_X1 U16764 ( .C1(n18884), .C2(n14853), .A(n13678), .B(n13677), .ZN(
        n13679) );
  OAI21_X1 U16765 ( .B1(n14557), .B2(n14601), .A(n13679), .ZN(P2_U2898) );
  AOI22_X1 U16766 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13684) );
  NOR2_X2 U16767 ( .A1(n13680), .A2(n13687), .ZN(n13732) );
  AOI22_X1 U16768 ( .A1(n13753), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13683) );
  NOR2_X2 U16769 ( .A1(n18434), .A2(n13680), .ZN(n15223) );
  AOI22_X1 U16770 ( .A1(n15223), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13682) );
  NOR2_X2 U16771 ( .A1(n16689), .A2(n13680), .ZN(n15048) );
  AOI22_X1 U16772 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13681) );
  NAND4_X1 U16773 ( .A1(n13684), .A2(n13683), .A3(n13682), .A4(n13681), .ZN(
        n13695) );
  CLKBUF_X3 U16774 ( .A(n15191), .Z(n16935) );
  NOR2_X2 U16775 ( .A1(n18574), .A2(n13685), .ZN(n15201) );
  AOI22_X1 U16776 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13693) );
  AOI22_X1 U16778 ( .A1(n16936), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9613), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13692) );
  AOI22_X1 U16779 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n16895), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13691) );
  INV_X2 U16780 ( .A(n9668), .ZN(n16954) );
  AOI22_X1 U16781 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9619), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13690) );
  NAND4_X1 U16782 ( .A1(n13693), .A2(n13692), .A3(n13691), .A4(n13690), .ZN(
        n13694) );
  INV_X1 U16783 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n15136) );
  INV_X1 U16784 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16562) );
  INV_X1 U16785 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n16971) );
  AOI22_X1 U16786 ( .A1(n15224), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9615), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13699) );
  AOI22_X1 U16787 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13698) );
  AOI22_X1 U16788 ( .A1(n9614), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13697) );
  AOI22_X1 U16789 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13696) );
  NAND4_X1 U16790 ( .A1(n13699), .A2(n13698), .A3(n13697), .A4(n13696), .ZN(
        n13706) );
  AOI22_X1 U16791 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15201), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13704) );
  INV_X1 U16792 ( .A(n13700), .ZN(n15112) );
  INV_X2 U16793 ( .A(n15112), .ZN(n16895) );
  AOI22_X1 U16794 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13703) );
  AOI22_X1 U16795 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13702) );
  AOI22_X1 U16796 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13701) );
  NAND4_X1 U16797 ( .A1(n13704), .A2(n13703), .A3(n13702), .A4(n13701), .ZN(
        n13705) );
  AOI22_X1 U16798 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13710) );
  AOI22_X1 U16799 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13709) );
  AOI22_X1 U16800 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13708) );
  AOI22_X1 U16801 ( .A1(n15223), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13707) );
  NAND4_X1 U16802 ( .A1(n13710), .A2(n13709), .A3(n13708), .A4(n13707), .ZN(
        n13716) );
  AOI22_X1 U16803 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15201), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13714) );
  AOI22_X1 U16804 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9615), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13713) );
  AOI22_X1 U16805 ( .A1(n15224), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13712) );
  AOI22_X1 U16806 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13711) );
  NAND4_X1 U16807 ( .A1(n13714), .A2(n13713), .A3(n13712), .A4(n13711), .ZN(
        n13715) );
  INV_X1 U16808 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18422) );
  OAI22_X1 U16809 ( .A1(n18583), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18420), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13721) );
  OAI22_X1 U16810 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18422), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13718), .ZN(n13724) );
  NOR2_X1 U16811 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18422), .ZN(
        n13719) );
  NAND2_X1 U16812 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13718), .ZN(
        n13723) );
  AOI22_X1 U16813 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13724), .B1(
        n13719), .B2(n13723), .ZN(n13727) );
  OAI21_X1 U16814 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18412), .A(
        n15170), .ZN(n15312) );
  NOR2_X1 U16815 ( .A1(n15169), .A2(n15312), .ZN(n13726) );
  OAI21_X1 U16816 ( .B1(n13722), .B2(n13721), .A(n13727), .ZN(n13720) );
  INV_X1 U16817 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18451) );
  AND2_X1 U16818 ( .A1(n13723), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13725) );
  OAI22_X1 U16819 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18451), .B1(
        n13725), .B2(n13724), .ZN(n15171) );
  AOI22_X1 U16820 ( .A1(n15224), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13731) );
  AOI22_X1 U16821 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13730) );
  AOI22_X1 U16822 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13729) );
  AOI22_X1 U16823 ( .A1(n15223), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16895), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13728) );
  NAND4_X1 U16824 ( .A1(n13731), .A2(n13730), .A3(n13729), .A4(n13728), .ZN(
        n13738) );
  AOI22_X1 U16825 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15201), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13736) );
  AOI22_X1 U16826 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16946), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13735) );
  AOI22_X1 U16827 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13734) );
  AOI22_X1 U16828 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9619), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13733) );
  NAND4_X1 U16829 ( .A1(n13736), .A2(n13735), .A3(n13734), .A4(n13733), .ZN(
        n13737) );
  INV_X1 U16830 ( .A(n15326), .ZN(n13782) );
  AOI22_X1 U16831 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13742) );
  AOI22_X1 U16832 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13741) );
  AOI22_X1 U16833 ( .A1(n15224), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13740) );
  AOI22_X1 U16834 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13739) );
  NAND4_X1 U16835 ( .A1(n13742), .A2(n13741), .A3(n13740), .A4(n13739), .ZN(
        n13748) );
  AOI22_X1 U16836 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15201), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13746) );
  AOI22_X1 U16837 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15223), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13745) );
  AOI22_X1 U16838 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13744) );
  AOI22_X1 U16839 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9619), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13743) );
  NAND4_X1 U16840 ( .A1(n13746), .A2(n13745), .A3(n13744), .A4(n13743), .ZN(
        n13747) );
  AOI22_X1 U16841 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9613), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13752) );
  AOI22_X1 U16842 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16895), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13751) );
  AOI22_X1 U16843 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13750) );
  AOI22_X1 U16844 ( .A1(n15224), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13749) );
  NAND4_X1 U16845 ( .A1(n13752), .A2(n13751), .A3(n13750), .A4(n13749), .ZN(
        n13759) );
  AOI22_X1 U16846 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13757) );
  AOI22_X1 U16847 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13756) );
  AOI22_X1 U16848 ( .A1(n15223), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13755) );
  AOI22_X1 U16849 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9619), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13754) );
  NAND4_X1 U16850 ( .A1(n13757), .A2(n13756), .A3(n13755), .A4(n13754), .ZN(
        n13758) );
  NOR2_X1 U16851 ( .A1(n13759), .A2(n13758), .ZN(n17993) );
  INV_X1 U16852 ( .A(n15319), .ZN(n15165) );
  AOI22_X1 U16853 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n15223), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13769) );
  AOI22_X1 U16854 ( .A1(n13753), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13768) );
  AOI22_X1 U16855 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9619), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13767) );
  AOI22_X1 U16856 ( .A1(n15224), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13763) );
  AOI22_X1 U16857 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13762) );
  AOI22_X1 U16858 ( .A1(n15048), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15260), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13761) );
  AOI22_X1 U16859 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13760) );
  NAND4_X1 U16860 ( .A1(n13763), .A2(n13762), .A3(n13761), .A4(n13760), .ZN(
        n13764) );
  AOI211_X1 U16861 ( .C1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .C2(n15201), .A(
        n13765), .B(n13764), .ZN(n13766) );
  NAND4_X1 U16862 ( .A1(n13769), .A2(n13768), .A3(n13767), .A4(n13766), .ZN(
        n15309) );
  BUF_X2 U16863 ( .A(n13770), .Z(n16948) );
  AOI22_X1 U16864 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13781) );
  AOI22_X1 U16865 ( .A1(n9628), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15260), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13780) );
  INV_X1 U16866 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16976) );
  AOI22_X1 U16867 ( .A1(n16909), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13771) );
  OAI21_X1 U16868 ( .B1(n15190), .B2(n16976), .A(n13771), .ZN(n13778) );
  AOI22_X1 U16869 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13776) );
  AOI22_X1 U16870 ( .A1(n13753), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13775) );
  AOI22_X1 U16871 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13774) );
  AOI22_X1 U16872 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9619), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13773) );
  NAND4_X1 U16873 ( .A1(n13776), .A2(n13775), .A3(n13774), .A4(n13773), .ZN(
        n13777) );
  AOI211_X1 U16874 ( .C1(n16947), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n13778), .B(n13777), .ZN(n13779) );
  NAND3_X1 U16875 ( .A1(n13781), .A2(n13780), .A3(n13779), .ZN(n15148) );
  NAND2_X1 U16876 ( .A1(n17997), .A2(n15148), .ZN(n18403) );
  NAND2_X1 U16877 ( .A1(n17985), .A2(n17981), .ZN(n18402) );
  NAND2_X1 U16878 ( .A1(n17993), .A2(n15309), .ZN(n15146) );
  NOR2_X1 U16879 ( .A1(n17108), .A2(n15148), .ZN(n13783) );
  AOI22_X1 U16880 ( .A1(n16126), .A2(n15331), .B1(n15160), .B2(n13783), .ZN(
        n15455) );
  NOR2_X1 U16881 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18566), .ZN(n18471) );
  NAND2_X1 U16882 ( .A1(n18471), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18459) );
  NAND3_X1 U16883 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(n9627), .ZN(n16983) );
  INV_X1 U16884 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n13785) );
  INV_X1 U16885 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n16644) );
  NAND2_X1 U16886 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_2__SCAN_IN), 
        .ZN(n13784) );
  INV_X1 U16887 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n15134) );
  INV_X1 U16888 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16437) );
  INV_X1 U16889 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16783) );
  NAND2_X1 U16890 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n15047) );
  NAND4_X1 U16891 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .A4(P3_EBX_REG_23__SCAN_IN), .ZN(n13786)
         );
  NOR4_X1 U16892 ( .A1(n16437), .A2(n16783), .A3(n15047), .A4(n13786), .ZN(
        n16731) );
  NAND2_X1 U16893 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16728), .ZN(n13788) );
  NOR2_X1 U16894 ( .A1(n17108), .A2(n13788), .ZN(n13790) );
  INV_X1 U16895 ( .A(n9627), .ZN(n16991) );
  NOR2_X2 U16896 ( .A1(n18005), .A2(n16991), .ZN(n16992) );
  INV_X2 U16897 ( .A(n16992), .ZN(n16986) );
  NAND2_X1 U16898 ( .A1(n16986), .A2(n13788), .ZN(n16729) );
  INV_X1 U16899 ( .A(n16729), .ZN(n13789) );
  MUX2_X1 U16900 ( .A(n13790), .B(n13789), .S(P3_EBX_REG_31__SCAN_IN), .Z(
        P3_U2672) );
  AOI22_X1 U16901 ( .A1(n13898), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n13897), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13896) );
  MUX2_X1 U16902 ( .A(n13829), .B(n13821), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n13796) );
  OAI21_X1 U16903 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n13898), .A(
        n13796), .ZN(n14056) );
  OR2_X1 U16904 ( .A1(n13831), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n13802) );
  INV_X1 U16905 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13797) );
  NAND2_X1 U16906 ( .A1(n13832), .A2(n13797), .ZN(n13800) );
  INV_X1 U16907 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n13798) );
  NAND2_X1 U16908 ( .A1(n13838), .A2(n13798), .ZN(n13799) );
  NAND3_X1 U16909 ( .A1(n13800), .A2(n13821), .A3(n13799), .ZN(n13801) );
  NAND2_X1 U16910 ( .A1(n13802), .A2(n13801), .ZN(n14044) );
  MUX2_X1 U16911 ( .A(n13829), .B(n13821), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n13803) );
  OAI21_X1 U16912 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n13898), .A(
        n13803), .ZN(n14033) );
  OR2_X1 U16913 ( .A1(n13831), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n13807) );
  NAND2_X1 U16914 ( .A1(n13832), .A2(n15638), .ZN(n13805) );
  INV_X1 U16915 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14127) );
  NAND2_X1 U16916 ( .A1(n13838), .A2(n14127), .ZN(n13804) );
  NAND3_X1 U16917 ( .A1(n13805), .A2(n13821), .A3(n13804), .ZN(n13806) );
  AND2_X1 U16918 ( .A1(n13807), .A2(n13806), .ZN(n14123) );
  MUX2_X1 U16919 ( .A(n13829), .B(n13821), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n13808) );
  OAI21_X1 U16920 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n13898), .A(
        n13808), .ZN(n14013) );
  MUX2_X1 U16921 ( .A(n13831), .B(n13832), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n13810) );
  NAND2_X1 U16922 ( .A1(n13897), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13809) );
  NAND2_X1 U16923 ( .A1(n13810), .A2(n13809), .ZN(n14118) );
  MUX2_X1 U16924 ( .A(n13829), .B(n13821), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n13812) );
  OR2_X1 U16925 ( .A1(n13898), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13811) );
  AND2_X1 U16926 ( .A1(n13812), .A2(n13811), .ZN(n14108) );
  MUX2_X1 U16927 ( .A(n13829), .B(n13821), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n13814) );
  OR2_X1 U16928 ( .A1(n13898), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13813) );
  AND2_X1 U16929 ( .A1(n13814), .A2(n13813), .ZN(n14098) );
  OR2_X1 U16930 ( .A1(n13831), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n13818) );
  INV_X1 U16931 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14277) );
  NAND2_X1 U16932 ( .A1(n13832), .A2(n14277), .ZN(n13816) );
  INV_X1 U16933 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15470) );
  NAND2_X1 U16934 ( .A1(n13838), .A2(n15470), .ZN(n13815) );
  NAND3_X1 U16935 ( .A1(n13816), .A2(n13821), .A3(n13815), .ZN(n13817) );
  NAND2_X1 U16936 ( .A1(n13818), .A2(n13817), .ZN(n14105) );
  NAND2_X1 U16937 ( .A1(n14098), .A2(n14105), .ZN(n13819) );
  OR2_X1 U16938 ( .A1(n13831), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n13824) );
  NAND2_X1 U16939 ( .A1(n13832), .A2(n15606), .ZN(n13822) );
  INV_X1 U16940 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14093) );
  NAND2_X1 U16941 ( .A1(n13838), .A2(n14093), .ZN(n13820) );
  NAND3_X1 U16942 ( .A1(n13822), .A2(n13821), .A3(n13820), .ZN(n13823) );
  AND2_X1 U16943 ( .A1(n13824), .A2(n13823), .ZN(n14001) );
  MUX2_X1 U16944 ( .A(n13829), .B(n13821), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n13826) );
  OR2_X1 U16945 ( .A1(n13898), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13825) );
  AND2_X1 U16946 ( .A1(n13826), .A2(n13825), .ZN(n13987) );
  MUX2_X1 U16947 ( .A(n13831), .B(n13832), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n13828) );
  NAND2_X1 U16948 ( .A1(n13897), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13827) );
  NAND2_X1 U16949 ( .A1(n13828), .A2(n13827), .ZN(n13971) );
  MUX2_X1 U16950 ( .A(n13829), .B(n13821), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n13830) );
  OAI21_X1 U16951 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13898), .A(
        n13830), .ZN(n13957) );
  OR2_X1 U16952 ( .A1(n13831), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n13837) );
  INV_X1 U16953 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14377) );
  NAND2_X1 U16954 ( .A1(n13832), .A2(n14377), .ZN(n13835) );
  INV_X1 U16955 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n13833) );
  NAND2_X1 U16956 ( .A1(n13838), .A2(n13833), .ZN(n13834) );
  NAND3_X1 U16957 ( .A1(n13835), .A2(n13821), .A3(n13834), .ZN(n13836) );
  AND2_X1 U16958 ( .A1(n13837), .A2(n13836), .ZN(n13952) );
  OR2_X1 U16959 ( .A1(n13898), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13839) );
  INV_X1 U16960 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14085) );
  NAND2_X1 U16961 ( .A1(n13838), .A2(n14085), .ZN(n13841) );
  NAND2_X1 U16962 ( .A1(n13839), .A2(n13841), .ZN(n13842) );
  MUX2_X1 U16963 ( .A(n13842), .B(n13841), .S(n13840), .Z(n13937) );
  OAI22_X1 U16964 ( .A1(n13938), .A2(n13821), .B1(n13842), .B2(n13951), .ZN(
        n13843) );
  XOR2_X1 U16965 ( .A(n13896), .B(n13843), .Z(n14083) );
  INV_X1 U16966 ( .A(n14083), .ZN(n13931) );
  NAND2_X1 U16967 ( .A1(n19819), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n13861) );
  INV_X1 U16968 ( .A(n13861), .ZN(n13857) );
  NOR2_X1 U16969 ( .A1(n15758), .A2(n15719), .ZN(n15740) );
  NAND4_X1 U16970 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n15740), .ZN(n13845) );
  NAND2_X1 U16971 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15697) );
  NOR4_X1 U16972 ( .A1(n13844), .A2(n13075), .A3(n13845), .A4(n15697), .ZN(
        n15673) );
  NAND3_X1 U16973 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n15673), .ZN(n14421) );
  INV_X1 U16974 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15647) );
  NAND2_X1 U16975 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15649) );
  NOR2_X1 U16976 ( .A1(n15647), .A2(n15649), .ZN(n15640) );
  NAND4_X1 U16977 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(n15640), .ZN(n13850) );
  NOR2_X1 U16978 ( .A1(n14421), .A2(n13850), .ZN(n14408) );
  NAND2_X1 U16979 ( .A1(n14408), .A2(n15672), .ZN(n14399) );
  INV_X1 U16980 ( .A(n13850), .ZN(n13848) );
  INV_X1 U16981 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15694) );
  NOR2_X1 U16982 ( .A1(n13846), .A2(n13845), .ZN(n15701) );
  NAND3_X1 U16983 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n15701), .ZN(n15688) );
  NOR2_X1 U16984 ( .A1(n15694), .A2(n15688), .ZN(n15682) );
  NAND2_X1 U16985 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15682), .ZN(
        n14420) );
  INV_X1 U16986 ( .A(n14421), .ZN(n15667) );
  NAND2_X1 U16987 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15667), .ZN(
        n13847) );
  OAI22_X1 U16988 ( .A1(n19829), .A2(n14420), .B1(n19828), .B2(n13847), .ZN(
        n15666) );
  NAND2_X1 U16989 ( .A1(n13848), .A2(n15666), .ZN(n14412) );
  NAND2_X1 U16990 ( .A1(n14399), .A2(n14412), .ZN(n15436) );
  INV_X1 U16991 ( .A(n15436), .ZN(n15637) );
  NOR3_X1 U16992 ( .A1(n13849), .A2(n14277), .A3(n15637), .ZN(n15618) );
  INV_X1 U16993 ( .A(n15618), .ZN(n15605) );
  NOR2_X1 U16994 ( .A1(n14224), .A2(n15605), .ZN(n14392) );
  NAND2_X1 U16995 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n14392), .ZN(
        n14372) );
  INV_X1 U16996 ( .A(n14372), .ZN(n14383) );
  INV_X1 U16997 ( .A(n14374), .ZN(n14365) );
  NAND3_X1 U16998 ( .A1(n14383), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14365), .ZN(n14352) );
  INV_X1 U16999 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14351) );
  NAND2_X1 U17000 ( .A1(n15702), .A2(n14423), .ZN(n14353) );
  INV_X1 U17001 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n20759) );
  INV_X1 U17002 ( .A(n14224), .ZN(n13853) );
  INV_X1 U17003 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15623) );
  NOR2_X1 U17004 ( .A1(n15623), .A2(n14277), .ZN(n15622) );
  NOR2_X1 U17005 ( .A1(n13850), .A2(n14420), .ZN(n14407) );
  AOI21_X1 U17006 ( .B1(n15674), .B2(n14407), .A(n14408), .ZN(n13852) );
  NAND2_X1 U17007 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n13851) );
  AOI221_X1 U17008 ( .B1(n13852), .B2(n15722), .C1(n13851), .C2(n15722), .A(
        n15676), .ZN(n15630) );
  OAI21_X1 U17009 ( .B1(n15702), .B2(n15622), .A(n15630), .ZN(n15617) );
  AOI21_X1 U17010 ( .B1(n14411), .B2(n20803), .A(n15617), .ZN(n14398) );
  OAI21_X1 U17011 ( .B1(n13853), .B2(n15702), .A(n14398), .ZN(n15610) );
  NAND2_X1 U17012 ( .A1(n14353), .A2(n10111), .ZN(n14386) );
  OR2_X1 U17013 ( .A1(n15702), .A2(n14365), .ZN(n13854) );
  AND2_X1 U17014 ( .A1(n14386), .A2(n13854), .ZN(n14361) );
  OAI211_X1 U17015 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15702), .A(
        n14361), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14354) );
  INV_X1 U17016 ( .A(n14354), .ZN(n13855) );
  AOI21_X1 U17017 ( .B1(n14352), .B2(n14351), .A(n13855), .ZN(n13856) );
  AOI211_X1 U17018 ( .C1(n13931), .C2(n19826), .A(n13857), .B(n13856), .ZN(
        n13858) );
  OAI21_X1 U17019 ( .B1(n13866), .B2(n15685), .A(n13858), .ZN(P1_U3001) );
  NAND2_X1 U17020 ( .A1(n15600), .A2(n13927), .ZN(n13862) );
  OAI211_X1 U17021 ( .C1(n13863), .C2(n15603), .A(n13862), .B(n13861), .ZN(
        n13864) );
  AOI21_X1 U17022 ( .B1(n13923), .B2(n14290), .A(n13864), .ZN(n13865) );
  OAI21_X1 U17023 ( .B1(n13866), .B2(n19637), .A(n13865), .ZN(P1_U2969) );
  NOR2_X1 U17024 ( .A1(n15819), .A2(n15859), .ZN(n13871) );
  AOI21_X1 U17025 ( .B1(n18934), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n13867), .ZN(n13868) );
  OAI21_X1 U17026 ( .B1(n13869), .B2(n18944), .A(n13868), .ZN(n13870) );
  AOI211_X1 U17027 ( .C1(n13872), .C2(n18936), .A(n13871), .B(n13870), .ZN(
        n13873) );
  OAI21_X1 U17028 ( .B1(n13874), .B2(n15941), .A(n13873), .ZN(P2_U2992) );
  NOR2_X1 U17029 ( .A1(n13875), .A2(n14605), .ZN(n13880) );
  INV_X1 U17030 ( .A(n13876), .ZN(n13878) );
  NOR2_X1 U17031 ( .A1(n13878), .A2(n13877), .ZN(n13879) );
  XNOR2_X1 U17032 ( .A(n13880), .B(n13879), .ZN(n14754) );
  NAND2_X1 U17033 ( .A1(n14754), .A2(n18936), .ZN(n13884) );
  NAND2_X1 U17034 ( .A1(n18933), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n14756) );
  OAI21_X1 U17035 ( .B1(n15941), .B2(n14757), .A(n14756), .ZN(n13882) );
  NOR2_X1 U17036 ( .A1(n18944), .A2(n13885), .ZN(n13881) );
  OAI211_X1 U17037 ( .C1(n14759), .C2(n15859), .A(n13884), .B(n13883), .ZN(
        P2_U2984) );
  NAND4_X1 U17038 ( .A1(n15772), .A2(n19499), .A3(n13264), .A4(n13885), .ZN(
        n13895) );
  NOR2_X1 U17039 ( .A1(n18795), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13892) );
  INV_X1 U17040 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n15812) );
  NOR2_X1 U17041 ( .A1(n13886), .A2(n15812), .ZN(n13888) );
  OAI22_X1 U17042 ( .A1(n18810), .A2(n11152), .B1(n11218), .B2(n18694), .ZN(
        n13887) );
  NOR2_X1 U17043 ( .A1(n13888), .A2(n13887), .ZN(n13889) );
  OAI21_X1 U17044 ( .B1(n13890), .B2(n18812), .A(n13889), .ZN(n13891) );
  AOI21_X1 U17045 ( .B1(n13893), .B2(n13892), .A(n13891), .ZN(n13894) );
  OAI211_X1 U17046 ( .C1(n15813), .C2(n18789), .A(n13895), .B(n13894), .ZN(
        P2_U2824) );
  AOI22_X1 U17047 ( .A1(n13898), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n13897), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13899) );
  NAND2_X1 U17048 ( .A1(n14221), .A2(n19663), .ZN(n13908) );
  NAND2_X1 U17049 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n13901) );
  INV_X1 U17050 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20558) );
  INV_X1 U17051 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20557) );
  NAND3_X1 U17052 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .A3(P1_REIP_REG_16__SCAN_IN), .ZN(n14017) );
  NAND3_X1 U17053 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(P1_REIP_REG_18__SCAN_IN), .ZN(n15469) );
  INV_X1 U17054 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20555) );
  INV_X1 U17055 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20553) );
  NOR2_X1 U17056 ( .A1(n20555), .A2(n20553), .ZN(n15461) );
  INV_X1 U17057 ( .A(n15461), .ZN(n15477) );
  NOR4_X1 U17058 ( .A1(n20557), .A2(n14017), .A3(n15469), .A4(n15477), .ZN(
        n13988) );
  NAND2_X1 U17059 ( .A1(n14014), .A2(n13988), .ZN(n14004) );
  NOR2_X1 U17060 ( .A1(n20558), .A2(n14004), .ZN(n13992) );
  NAND3_X1 U17061 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .A3(n13992), .ZN(n13961) );
  INV_X1 U17062 ( .A(n13961), .ZN(n13900) );
  NAND2_X1 U17063 ( .A1(n19708), .A2(n13900), .ZN(n13960) );
  OAI21_X1 U17064 ( .B1(n13901), .B2(n13960), .A(n15468), .ZN(n13933) );
  INV_X1 U17065 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n13904) );
  OAI21_X1 U17066 ( .B1(n20572), .B2(n13904), .A(n14015), .ZN(n13902) );
  NAND2_X1 U17067 ( .A1(n13933), .A2(n13902), .ZN(n13925) );
  INV_X1 U17068 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13903) );
  INV_X1 U17069 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14082) );
  OAI22_X1 U17070 ( .A1(n13903), .A2(n15525), .B1(n19715), .B2(n14082), .ZN(
        n13906) );
  INV_X1 U17071 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20565) );
  NOR3_X1 U17072 ( .A1(n19709), .A2(n20565), .A3(n13961), .ZN(n13945) );
  NAND3_X1 U17073 ( .A1(n13945), .A2(P1_REIP_REG_29__SCAN_IN), .A3(
        P1_REIP_REG_28__SCAN_IN), .ZN(n13924) );
  NOR3_X1 U17074 ( .A1(n13924), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n13904), 
        .ZN(n13905) );
  AOI211_X1 U17075 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n13925), .A(n13906), 
        .B(n13905), .ZN(n13907) );
  OAI211_X1 U17076 ( .C1(n14350), .C2(n19718), .A(n13908), .B(n13907), .ZN(
        P1_U2809) );
  NOR2_X1 U17077 ( .A1(n14759), .A2(n18875), .ZN(n13909) );
  AOI21_X1 U17078 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n18875), .A(n13909), .ZN(
        n13910) );
  OAI21_X1 U17079 ( .B1(n13911), .B2(n18865), .A(n13910), .ZN(P2_U2857) );
  NAND2_X1 U17080 ( .A1(n13914), .A2(n13913), .ZN(n14517) );
  NAND2_X1 U17081 ( .A1(n14517), .A2(n18885), .ZN(n13922) );
  NAND2_X1 U17082 ( .A1(n14468), .A2(n13915), .ZN(n13916) );
  NAND2_X1 U17083 ( .A1(n9666), .A2(n13916), .ZN(n15784) );
  OAI22_X1 U17084 ( .A1(n15784), .A2(n14585), .B1(n14596), .B2(n13917), .ZN(
        n13918) );
  AOI21_X1 U17085 ( .B1(n18880), .B2(n13919), .A(n13918), .ZN(n13921) );
  AOI22_X1 U17086 ( .A1(n18882), .A2(BUF1_REG_29__SCAN_IN), .B1(n18881), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n13920) );
  OAI211_X1 U17087 ( .C1(n13912), .C2(n13922), .A(n13921), .B(n13920), .ZN(
        P2_U2890) );
  INV_X1 U17088 ( .A(n13923), .ZN(n14150) );
  INV_X1 U17089 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14084) );
  INV_X1 U17090 ( .A(n13924), .ZN(n13926) );
  OAI21_X1 U17091 ( .B1(n13926), .B2(P1_REIP_REG_30__SCAN_IN), .A(n13925), 
        .ZN(n13929) );
  AOI22_X1 U17092 ( .A1(n13927), .A2(n19703), .B1(n19721), .B2(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13928) );
  OAI211_X1 U17093 ( .C1(n19715), .C2(n14084), .A(n13929), .B(n13928), .ZN(
        n13930) );
  AOI21_X1 U17094 ( .B1(n13931), .B2(n19700), .A(n13930), .ZN(n13932) );
  OAI21_X1 U17095 ( .B1(n14150), .B2(n15521), .A(n13932), .ZN(P1_U2810) );
  INV_X1 U17096 ( .A(n13933), .ZN(n13950) );
  NAND3_X1 U17097 ( .A1(n13945), .A2(P1_REIP_REG_28__SCAN_IN), .A3(n20572), 
        .ZN(n13936) );
  AOI22_X1 U17098 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19721), .B1(
        n19703), .B2(n13934), .ZN(n13935) );
  OAI211_X1 U17099 ( .C1(n14085), .C2(n19715), .A(n13936), .B(n13935), .ZN(
        n13941) );
  AND2_X1 U17100 ( .A1(n13951), .A2(n13937), .ZN(n13939) );
  OR2_X1 U17101 ( .A1(n13939), .A2(n13938), .ZN(n14368) );
  NOR2_X1 U17102 ( .A1(n14368), .A2(n19718), .ZN(n13940) );
  AOI211_X1 U17103 ( .C1(n13950), .C2(P1_REIP_REG_29__SCAN_IN), .A(n13941), 
        .B(n13940), .ZN(n13942) );
  OAI21_X1 U17104 ( .B1(n14153), .B2(n15521), .A(n13942), .ZN(P1_U2811) );
  AOI21_X1 U17105 ( .B1(n13944), .B2(n13943), .A(n12588), .ZN(n14234) );
  INV_X1 U17106 ( .A(n14234), .ZN(n14156) );
  INV_X1 U17107 ( .A(n13945), .ZN(n13948) );
  AOI22_X1 U17108 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19721), .B1(
        n19703), .B2(n14230), .ZN(n13947) );
  NAND2_X1 U17109 ( .A1(n19695), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n13946) );
  OAI211_X1 U17110 ( .C1(n13948), .C2(P1_REIP_REG_28__SCAN_IN), .A(n13947), 
        .B(n13946), .ZN(n13949) );
  AOI21_X1 U17111 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n13950), .A(n13949), 
        .ZN(n13954) );
  AOI21_X1 U17112 ( .B1(n13952), .B2(n13959), .A(n9892), .ZN(n14379) );
  NAND2_X1 U17113 ( .A1(n14379), .A2(n19700), .ZN(n13953) );
  OAI211_X1 U17114 ( .C1(n14156), .C2(n15521), .A(n13954), .B(n13953), .ZN(
        P1_U2812) );
  INV_X1 U17115 ( .A(n13943), .ZN(n13955) );
  AOI21_X1 U17116 ( .B1(n13956), .B2(n13969), .A(n13955), .ZN(n14243) );
  INV_X1 U17117 ( .A(n14243), .ZN(n14159) );
  NAND2_X1 U17118 ( .A1(n13973), .A2(n13957), .ZN(n13958) );
  AND2_X1 U17119 ( .A1(n13959), .A2(n13958), .ZN(n14388) );
  NAND2_X1 U17120 ( .A1(n15468), .A2(n13960), .ZN(n13974) );
  NOR3_X1 U17121 ( .A1(n19709), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n13961), 
        .ZN(n13964) );
  OAI22_X1 U17122 ( .A1(n13962), .A2(n15525), .B1(n19731), .B2(n14241), .ZN(
        n13963) );
  AOI211_X1 U17123 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n19695), .A(n13964), .B(
        n13963), .ZN(n13965) );
  OAI21_X1 U17124 ( .B1(n20565), .B2(n13974), .A(n13965), .ZN(n13966) );
  AOI21_X1 U17125 ( .B1(n14388), .B2(n19700), .A(n13966), .ZN(n13967) );
  OAI21_X1 U17126 ( .B1(n14159), .B2(n15521), .A(n13967), .ZN(P1_U2813) );
  AND2_X1 U17127 ( .A1(n13980), .A2(n13968), .ZN(n13982) );
  OAI21_X1 U17128 ( .B1(n13982), .B2(n13970), .A(n13969), .ZN(n14253) );
  OR2_X1 U17129 ( .A1(n13985), .A2(n13971), .ZN(n13972) );
  NAND2_X1 U17130 ( .A1(n13973), .A2(n13972), .ZN(n14088) );
  INV_X1 U17131 ( .A(n14088), .ZN(n14394) );
  INV_X1 U17132 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20563) );
  NAND3_X1 U17133 ( .A1(n14015), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n13992), 
        .ZN(n13975) );
  AOI21_X1 U17134 ( .B1(n20563), .B2(n13975), .A(n13974), .ZN(n13978) );
  INV_X1 U17135 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14089) );
  AOI22_X1 U17136 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19721), .B1(
        n19703), .B2(n14247), .ZN(n13976) );
  OAI21_X1 U17137 ( .B1(n19715), .B2(n14089), .A(n13976), .ZN(n13977) );
  AOI211_X1 U17138 ( .C1(n14394), .C2(n19700), .A(n13978), .B(n13977), .ZN(
        n13979) );
  OAI21_X1 U17139 ( .B1(n14253), .B2(n15521), .A(n13979), .ZN(P1_U2814) );
  AOI21_X1 U17140 ( .B1(n13983), .B2(n13998), .A(n13982), .ZN(n13984) );
  INV_X1 U17141 ( .A(n13984), .ZN(n14264) );
  INV_X1 U17142 ( .A(n13985), .ZN(n13986) );
  OAI21_X1 U17143 ( .B1(n13987), .B2(n14003), .A(n13986), .ZN(n14091) );
  INV_X1 U17144 ( .A(n14091), .ZN(n15611) );
  INV_X1 U17145 ( .A(n13988), .ZN(n13990) );
  OAI21_X1 U17146 ( .B1(n13990), .B2(n13989), .A(n15468), .ZN(n15466) );
  INV_X1 U17147 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20561) );
  NOR2_X1 U17148 ( .A1(n15466), .A2(n20561), .ZN(n13996) );
  INV_X1 U17149 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14090) );
  NAND2_X1 U17150 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n13991) );
  OAI211_X1 U17151 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n13992), .A(n14015), 
        .B(n13991), .ZN(n13994) );
  AOI22_X1 U17152 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19721), .B1(
        n19703), .B2(n14256), .ZN(n13993) );
  OAI211_X1 U17153 ( .C1(n14090), .C2(n19715), .A(n13994), .B(n13993), .ZN(
        n13995) );
  AOI211_X1 U17154 ( .C1(n15611), .C2(n19700), .A(n13996), .B(n13995), .ZN(
        n13997) );
  OAI21_X1 U17155 ( .B1(n14264), .B2(n15521), .A(n13997), .ZN(P1_U2815) );
  INV_X1 U17156 ( .A(n13998), .ZN(n13999) );
  NAND2_X1 U17157 ( .A1(n14273), .A2(n19663), .ZN(n14009) );
  AND2_X1 U17158 ( .A1(n14099), .A2(n14001), .ZN(n14002) );
  NOR2_X1 U17159 ( .A1(n14003), .A2(n14002), .ZN(n14092) );
  NOR3_X1 U17160 ( .A1(n19709), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n14004), 
        .ZN(n14007) );
  AOI22_X1 U17161 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19721), .B1(
        n19703), .B2(n14269), .ZN(n14005) );
  OAI21_X1 U17162 ( .B1(n19715), .B2(n14093), .A(n14005), .ZN(n14006) );
  AOI211_X1 U17163 ( .C1(n14092), .C2(n19700), .A(n14007), .B(n14006), .ZN(
        n14008) );
  OAI211_X1 U17164 ( .C1(n15466), .C2(n20558), .A(n14009), .B(n14008), .ZN(
        P1_U2816) );
  INV_X1 U17165 ( .A(n14010), .ZN(n14027) );
  AOI21_X1 U17166 ( .B1(n14027), .B2(n14122), .A(n14011), .ZN(n14012) );
  NOR2_X1 U17167 ( .A1(n14012), .A2(n9670), .ZN(n15546) );
  INV_X1 U17168 ( .A(n15546), .ZN(n14188) );
  AOI21_X1 U17169 ( .B1(n14013), .B2(n14126), .A(n14119), .ZN(n15633) );
  NAND2_X1 U17170 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n14041) );
  NAND2_X1 U17171 ( .A1(n14015), .A2(n14014), .ZN(n14055) );
  NOR2_X1 U17172 ( .A1(n14041), .A2(n14055), .ZN(n14029) );
  NAND2_X1 U17173 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14029), .ZN(n15506) );
  NAND2_X1 U17174 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n15491) );
  OAI21_X1 U17175 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(P1_REIP_REG_18__SCAN_IN), 
        .A(n15491), .ZN(n14016) );
  OAI22_X1 U17176 ( .A1(n15549), .A2(n19731), .B1(n15506), .B2(n14016), .ZN(
        n14023) );
  INV_X1 U17177 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14021) );
  INV_X1 U17178 ( .A(n14017), .ZN(n14019) );
  INV_X1 U17179 ( .A(n15468), .ZN(n14018) );
  OAI21_X1 U17180 ( .B1(n14019), .B2(n14018), .A(n14054), .ZN(n15500) );
  AOI22_X1 U17181 ( .A1(n15500), .A2(P1_REIP_REG_19__SCAN_IN), .B1(n19695), 
        .B2(P1_EBX_REG_19__SCAN_IN), .ZN(n14020) );
  OAI211_X1 U17182 ( .C1(n15525), .C2(n14021), .A(n14020), .B(n19683), .ZN(
        n14022) );
  AOI211_X1 U17183 ( .C1(n15633), .C2(n19700), .A(n14023), .B(n14022), .ZN(
        n14024) );
  OAI21_X1 U17184 ( .B1(n14188), .B2(n15521), .A(n14024), .ZN(P1_U2821) );
  INV_X1 U17185 ( .A(n14026), .ZN(n14028) );
  NAND2_X1 U17186 ( .A1(n15556), .A2(n19663), .ZN(n14037) );
  OAI21_X1 U17187 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n14029), .A(n15500), 
        .ZN(n14036) );
  INV_X1 U17188 ( .A(n19683), .ZN(n19662) );
  NOR2_X1 U17189 ( .A1(n15525), .A2(n14030), .ZN(n14031) );
  AOI211_X1 U17190 ( .C1(n19703), .C2(n15555), .A(n19662), .B(n14031), .ZN(
        n14035) );
  INV_X1 U17191 ( .A(n14124), .ZN(n14032) );
  AOI21_X1 U17192 ( .B1(n14033), .B2(n14043), .A(n14032), .ZN(n15650) );
  AOI22_X1 U17193 ( .A1(n15650), .A2(n19700), .B1(n19695), .B2(
        P1_EBX_REG_17__SCAN_IN), .ZN(n14034) );
  NAND4_X1 U17194 ( .A1(n14037), .A2(n14036), .A3(n14035), .A4(n14034), .ZN(
        P1_U2823) );
  AND2_X1 U17195 ( .A1(n14038), .A2(n14039), .ZN(n14040) );
  NOR2_X1 U17196 ( .A1(n14026), .A2(n14040), .ZN(n14313) );
  INV_X1 U17197 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20545) );
  OAI21_X1 U17198 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(P1_REIP_REG_16__SCAN_IN), 
        .A(n14041), .ZN(n14042) );
  OAI22_X1 U17199 ( .A1(n20545), .A2(n14054), .B1(n14055), .B2(n14042), .ZN(
        n14049) );
  OAI21_X1 U17200 ( .B1(n14059), .B2(n14044), .A(n14043), .ZN(n14427) );
  INV_X1 U17201 ( .A(n14427), .ZN(n14131) );
  AOI22_X1 U17202 ( .A1(n14131), .A2(n19700), .B1(n19695), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n14047) );
  NAND2_X1 U17203 ( .A1(n19703), .A2(n14309), .ZN(n14046) );
  NAND2_X1 U17204 ( .A1(n19721), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14045) );
  NAND4_X1 U17205 ( .A1(n14047), .A2(n19683), .A3(n14046), .A4(n14045), .ZN(
        n14048) );
  AOI211_X1 U17206 ( .C1(n14313), .C2(n19663), .A(n14049), .B(n14048), .ZN(
        n14050) );
  INV_X1 U17207 ( .A(n14050), .ZN(P1_U2824) );
  AOI21_X1 U17208 ( .B1(n14052), .B2(n14051), .A(n9978), .ZN(n15564) );
  INV_X1 U17209 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20542) );
  AOI21_X1 U17210 ( .B1(n19721), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n19662), .ZN(n14053) );
  OAI221_X1 U17211 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n14055), .C1(n20542), 
        .C2(n14054), .A(n14053), .ZN(n14062) );
  AND2_X1 U17212 ( .A1(n14057), .A2(n14056), .ZN(n14058) );
  OR2_X1 U17213 ( .A1(n14059), .A2(n14058), .ZN(n15656) );
  AOI22_X1 U17214 ( .A1(n19695), .A2(P1_EBX_REG_15__SCAN_IN), .B1(n19703), 
        .B2(n15563), .ZN(n14060) );
  OAI21_X1 U17215 ( .B1(n19718), .B2(n15656), .A(n14060), .ZN(n14061) );
  AOI211_X1 U17216 ( .C1(n15564), .C2(n19663), .A(n14062), .B(n14061), .ZN(
        n14063) );
  INV_X1 U17217 ( .A(n14063), .ZN(P1_U2825) );
  INV_X1 U17218 ( .A(n14064), .ZN(n14066) );
  OAI21_X1 U17219 ( .B1(n14067), .B2(n14066), .A(n14065), .ZN(n14141) );
  AND2_X1 U17220 ( .A1(n14141), .A2(n14140), .ZN(n14143) );
  OAI21_X1 U17221 ( .B1(n14143), .B2(n14068), .A(n13638), .ZN(n14335) );
  INV_X1 U17222 ( .A(n14139), .ZN(n14071) );
  INV_X1 U17223 ( .A(n14069), .ZN(n14070) );
  AOI21_X1 U17224 ( .B1(n14072), .B2(n14071), .A(n14070), .ZN(n15663) );
  OAI21_X1 U17225 ( .B1(n14074), .B2(n19709), .A(n19708), .ZN(n15518) );
  AOI22_X1 U17226 ( .A1(n19703), .A2(n14332), .B1(P1_REIP_REG_13__SCAN_IN), 
        .B2(n15518), .ZN(n14073) );
  INV_X1 U17227 ( .A(n14073), .ZN(n14080) );
  INV_X1 U17228 ( .A(n14074), .ZN(n14075) );
  NOR3_X1 U17229 ( .A1(n19709), .A2(P1_REIP_REG_13__SCAN_IN), .A3(n14075), 
        .ZN(n14076) );
  AOI21_X1 U17230 ( .B1(P1_EBX_REG_13__SCAN_IN), .B2(n19695), .A(n14076), .ZN(
        n14077) );
  OAI211_X1 U17231 ( .C1(n15525), .C2(n14078), .A(n14077), .B(n19683), .ZN(
        n14079) );
  AOI211_X1 U17232 ( .C1(n15663), .C2(n19700), .A(n14080), .B(n14079), .ZN(
        n14081) );
  OAI21_X1 U17233 ( .B1(n14335), .B2(n15521), .A(n14081), .ZN(P1_U2827) );
  OAI22_X1 U17234 ( .A1(n14350), .A2(n14146), .B1(n19742), .B2(n14082), .ZN(
        P1_U2841) );
  OAI222_X1 U17235 ( .A1(n14144), .A2(n14150), .B1(n14084), .B2(n19742), .C1(
        n14083), .C2(n14146), .ZN(P1_U2842) );
  OAI222_X1 U17236 ( .A1(n14144), .A2(n14153), .B1(n14085), .B2(n19742), .C1(
        n14368), .C2(n14146), .ZN(P1_U2843) );
  AOI22_X1 U17237 ( .A1(n14379), .A2(n19738), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n14134), .ZN(n14086) );
  OAI21_X1 U17238 ( .B1(n14156), .B2(n14136), .A(n14086), .ZN(P1_U2844) );
  AOI22_X1 U17239 ( .A1(n14388), .A2(n19738), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n14134), .ZN(n14087) );
  OAI21_X1 U17240 ( .B1(n14159), .B2(n14136), .A(n14087), .ZN(P1_U2845) );
  OAI222_X1 U17241 ( .A1(n14144), .A2(n14253), .B1(n14089), .B2(n19742), .C1(
        n14088), .C2(n14146), .ZN(P1_U2846) );
  OAI222_X1 U17242 ( .A1(n14091), .A2(n14146), .B1(n14090), .B2(n19742), .C1(
        n14264), .C2(n14144), .ZN(P1_U2847) );
  INV_X1 U17243 ( .A(n14273), .ZN(n14167) );
  INV_X1 U17244 ( .A(n14092), .ZN(n14401) );
  OAI222_X1 U17245 ( .A1(n14144), .A2(n14167), .B1(n14093), .B2(n19742), .C1(
        n14401), .C2(n14146), .ZN(P1_U2848) );
  INV_X1 U17246 ( .A(n14094), .ZN(n14095) );
  AOI21_X1 U17247 ( .B1(n14096), .B2(n14103), .A(n14095), .ZN(n15531) );
  INV_X1 U17248 ( .A(n15531), .ZN(n14171) );
  AOI21_X1 U17249 ( .B1(n9900), .B2(n14105), .A(n14098), .ZN(n14100) );
  NOR2_X1 U17250 ( .A1(n14100), .A2(n9904), .ZN(n15614) );
  AOI22_X1 U17251 ( .A1(n15614), .A2(n19738), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n14134), .ZN(n14101) );
  OAI21_X1 U17252 ( .B1(n14171), .B2(n14136), .A(n14101), .ZN(P1_U2849) );
  INV_X1 U17253 ( .A(n14105), .ZN(n14106) );
  XNOR2_X1 U17254 ( .A(n14097), .B(n14106), .ZN(n15472) );
  INV_X1 U17255 ( .A(n15472), .ZN(n15626) );
  AOI22_X1 U17256 ( .A1(n15626), .A2(n19738), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n14134), .ZN(n14107) );
  OAI21_X1 U17257 ( .B1(n15473), .B2(n14136), .A(n14107), .ZN(P1_U2850) );
  OR2_X1 U17258 ( .A1(n14116), .A2(n14108), .ZN(n14109) );
  NAND2_X1 U17259 ( .A1(n14097), .A2(n14109), .ZN(n15484) );
  INV_X1 U17260 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14113) );
  NOR2_X1 U17261 ( .A1(n14110), .A2(n14111), .ZN(n14112) );
  OR2_X1 U17262 ( .A1(n14102), .A2(n14112), .ZN(n15539) );
  OAI222_X1 U17263 ( .A1(n15484), .A2(n14146), .B1(n14113), .B2(n19742), .C1(
        n15539), .C2(n14144), .ZN(P1_U2851) );
  AOI21_X1 U17264 ( .B1(n14115), .B2(n14114), .A(n14110), .ZN(n14291) );
  INV_X1 U17265 ( .A(n14291), .ZN(n15493) );
  INV_X1 U17266 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14120) );
  INV_X1 U17267 ( .A(n14116), .ZN(n14117) );
  OAI21_X1 U17268 ( .B1(n14119), .B2(n14118), .A(n14117), .ZN(n15492) );
  OAI222_X1 U17269 ( .A1(n15493), .A2(n14136), .B1(n19742), .B2(n14120), .C1(
        n15492), .C2(n14146), .ZN(P1_U2852) );
  AOI22_X1 U17270 ( .A1(n15633), .A2(n19738), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14134), .ZN(n14121) );
  OAI21_X1 U17271 ( .B1(n14188), .B2(n14144), .A(n14121), .ZN(P1_U2853) );
  XNOR2_X1 U17272 ( .A(n14010), .B(n14122), .ZN(n15508) );
  INV_X1 U17273 ( .A(n15508), .ZN(n14192) );
  NAND2_X1 U17274 ( .A1(n14124), .A2(n14123), .ZN(n14125) );
  NAND2_X1 U17275 ( .A1(n14126), .A2(n14125), .ZN(n15641) );
  OAI22_X1 U17276 ( .A1(n15641), .A2(n14146), .B1(n14127), .B2(n19742), .ZN(
        n14128) );
  INV_X1 U17277 ( .A(n14128), .ZN(n14129) );
  OAI21_X1 U17278 ( .B1(n14192), .B2(n14144), .A(n14129), .ZN(P1_U2854) );
  INV_X1 U17279 ( .A(n15556), .ZN(n14196) );
  AOI22_X1 U17280 ( .A1(n15650), .A2(n19738), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14134), .ZN(n14130) );
  OAI21_X1 U17281 ( .B1(n14196), .B2(n14144), .A(n14130), .ZN(P1_U2855) );
  INV_X1 U17282 ( .A(n14313), .ZN(n14203) );
  AOI22_X1 U17283 ( .A1(n14131), .A2(n19738), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n14134), .ZN(n14132) );
  OAI21_X1 U17284 ( .B1(n14203), .B2(n14144), .A(n14132), .ZN(P1_U2856) );
  INV_X1 U17285 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14133) );
  INV_X1 U17286 ( .A(n15564), .ZN(n14205) );
  OAI222_X1 U17287 ( .A1(n15656), .A2(n14146), .B1(n14133), .B2(n19742), .C1(
        n14205), .C2(n14144), .ZN(P1_U2857) );
  AOI22_X1 U17288 ( .A1(n15663), .A2(n19738), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14134), .ZN(n14135) );
  OAI21_X1 U17289 ( .B1(n14335), .B2(n14136), .A(n14135), .ZN(P1_U2859) );
  NOR2_X1 U17290 ( .A1(n9733), .A2(n14137), .ZN(n14138) );
  OR2_X1 U17291 ( .A1(n14139), .A2(n14138), .ZN(n15678) );
  INV_X1 U17292 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14145) );
  NOR2_X1 U17293 ( .A1(n14141), .A2(n14140), .ZN(n14142) );
  OAI222_X1 U17294 ( .A1(n15678), .A2(n14146), .B1(n19742), .B2(n14145), .C1(
        n15571), .C2(n14144), .ZN(P1_U2860) );
  AOI22_X1 U17295 ( .A1(n14197), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14206), .ZN(n14149) );
  AOI22_X1 U17296 ( .A1(n14200), .A2(n19791), .B1(n14198), .B2(DATAI_30_), 
        .ZN(n14148) );
  OAI211_X1 U17297 ( .C1(n14150), .C2(n14209), .A(n14149), .B(n14148), .ZN(
        P1_U2874) );
  AOI22_X1 U17298 ( .A1(n14197), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14206), .ZN(n14152) );
  MUX2_X1 U17299 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n19839), .Z(
        n19789) );
  AOI22_X1 U17300 ( .A1(n14200), .A2(n19789), .B1(n14198), .B2(DATAI_29_), 
        .ZN(n14151) );
  OAI211_X1 U17301 ( .C1(n14153), .C2(n14209), .A(n14152), .B(n14151), .ZN(
        P1_U2875) );
  AOI22_X1 U17302 ( .A1(n14197), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14206), .ZN(n14155) );
  MUX2_X1 U17303 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n19839), .Z(
        n19787) );
  AOI22_X1 U17304 ( .A1(n14200), .A2(n19787), .B1(n14198), .B2(DATAI_28_), 
        .ZN(n14154) );
  OAI211_X1 U17305 ( .C1(n14156), .C2(n14209), .A(n14155), .B(n14154), .ZN(
        P1_U2876) );
  AOI22_X1 U17306 ( .A1(n14197), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14206), .ZN(n14158) );
  AOI22_X1 U17307 ( .A1(n14200), .A2(n19785), .B1(n14198), .B2(DATAI_27_), 
        .ZN(n14157) );
  OAI211_X1 U17308 ( .C1(n14159), .C2(n14209), .A(n14158), .B(n14157), .ZN(
        P1_U2877) );
  AOI22_X1 U17309 ( .A1(n14197), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n14206), .ZN(n14161) );
  AOI22_X1 U17310 ( .A1(n14200), .A2(n19783), .B1(n14198), .B2(DATAI_26_), 
        .ZN(n14160) );
  OAI211_X1 U17311 ( .C1(n14253), .C2(n14209), .A(n14161), .B(n14160), .ZN(
        P1_U2878) );
  AOI22_X1 U17312 ( .A1(n14197), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14206), .ZN(n14164) );
  AOI22_X1 U17313 ( .A1(n14200), .A2(n14162), .B1(n14198), .B2(DATAI_25_), 
        .ZN(n14163) );
  OAI211_X1 U17314 ( .C1(n14264), .C2(n14209), .A(n14164), .B(n14163), .ZN(
        P1_U2879) );
  AOI22_X1 U17315 ( .A1(n14197), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n14206), .ZN(n14166) );
  AOI22_X1 U17316 ( .A1(n14200), .A2(n19781), .B1(n14198), .B2(DATAI_24_), 
        .ZN(n14165) );
  OAI211_X1 U17317 ( .C1(n14167), .C2(n14209), .A(n14166), .B(n14165), .ZN(
        P1_U2880) );
  AOI22_X1 U17318 ( .A1(n14197), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n14206), .ZN(n14170) );
  AOI22_X1 U17319 ( .A1(n14200), .A2(n14168), .B1(n14198), .B2(DATAI_23_), 
        .ZN(n14169) );
  OAI211_X1 U17320 ( .C1(n14171), .C2(n14209), .A(n14170), .B(n14169), .ZN(
        P1_U2881) );
  AOI22_X1 U17321 ( .A1(n14197), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n14206), .ZN(n14174) );
  AOI22_X1 U17322 ( .A1(n14200), .A2(n14172), .B1(n14198), .B2(DATAI_22_), 
        .ZN(n14173) );
  OAI211_X1 U17323 ( .C1(n15473), .C2(n14209), .A(n14174), .B(n14173), .ZN(
        P1_U2882) );
  OAI22_X1 U17324 ( .A1(n14177), .A2(n14176), .B1(n14175), .B2(n14210), .ZN(
        n14180) );
  INV_X1 U17325 ( .A(n14200), .ZN(n14178) );
  NOR2_X1 U17326 ( .A1(n14178), .A2(n19878), .ZN(n14179) );
  AOI211_X1 U17327 ( .C1(n14198), .C2(DATAI_21_), .A(n14180), .B(n14179), .ZN(
        n14181) );
  OAI21_X1 U17328 ( .B1(n15539), .B2(n14209), .A(n14181), .ZN(P1_U2883) );
  AOI22_X1 U17329 ( .A1(n14197), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n14206), .ZN(n14184) );
  AOI22_X1 U17330 ( .A1(n14200), .A2(n14182), .B1(n14198), .B2(DATAI_20_), 
        .ZN(n14183) );
  OAI211_X1 U17331 ( .C1(n15493), .C2(n14209), .A(n14184), .B(n14183), .ZN(
        P1_U2884) );
  AOI22_X1 U17332 ( .A1(n14197), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14206), .ZN(n14187) );
  AOI22_X1 U17333 ( .A1(n14200), .A2(n14185), .B1(n14198), .B2(DATAI_19_), 
        .ZN(n14186) );
  OAI211_X1 U17334 ( .C1(n14188), .C2(n14209), .A(n14187), .B(n14186), .ZN(
        P1_U2885) );
  AOI22_X1 U17335 ( .A1(n14197), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n14206), .ZN(n14191) );
  AOI22_X1 U17336 ( .A1(n14200), .A2(n14189), .B1(n14198), .B2(DATAI_18_), 
        .ZN(n14190) );
  OAI211_X1 U17337 ( .C1(n14192), .C2(n14209), .A(n14191), .B(n14190), .ZN(
        P1_U2886) );
  AOI22_X1 U17338 ( .A1(n14197), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14206), .ZN(n14195) );
  AOI22_X1 U17339 ( .A1(n14200), .A2(n14193), .B1(n14198), .B2(DATAI_17_), 
        .ZN(n14194) );
  OAI211_X1 U17340 ( .C1(n14196), .C2(n14209), .A(n14195), .B(n14194), .ZN(
        P1_U2887) );
  AOI22_X1 U17341 ( .A1(n14197), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n14206), .ZN(n14202) );
  AOI22_X1 U17342 ( .A1(n14200), .A2(n14199), .B1(n14198), .B2(DATAI_16_), 
        .ZN(n14201) );
  OAI211_X1 U17343 ( .C1(n14203), .C2(n14209), .A(n14202), .B(n14201), .ZN(
        P1_U2888) );
  OAI222_X1 U17344 ( .A1(n14205), .A2(n14209), .B1(n14213), .B2(n14204), .C1(
        n14210), .C2(n19748), .ZN(P1_U2889) );
  AOI22_X1 U17345 ( .A1(n14207), .A2(n19789), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14206), .ZN(n14208) );
  OAI21_X1 U17346 ( .B1(n14335), .B2(n14209), .A(n14208), .ZN(P1_U2891) );
  INV_X1 U17347 ( .A(n19787), .ZN(n14212) );
  OAI222_X1 U17348 ( .A1(n15571), .A2(n14209), .B1(n14213), .B2(n14212), .C1(
        n14211), .C2(n14210), .ZN(P1_U2892) );
  NAND2_X1 U17349 ( .A1(n14214), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14215) );
  XNOR2_X1 U17350 ( .A(n14217), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14360) );
  INV_X1 U17351 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20576) );
  NOR2_X1 U17352 ( .A1(n15731), .A2(n20576), .ZN(n14356) );
  AOI21_X1 U17353 ( .B1(n19813), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14356), .ZN(n14218) );
  OAI21_X1 U17354 ( .B1(n15597), .B2(n14219), .A(n14218), .ZN(n14220) );
  OAI21_X1 U17355 ( .B1(n14360), .B2(n19637), .A(n14222), .ZN(P1_U2968) );
  NAND2_X1 U17356 ( .A1(n15529), .A2(n14224), .ZN(n14248) );
  NAND2_X1 U17357 ( .A1(n14223), .A2(n14248), .ZN(n14228) );
  OAI21_X1 U17358 ( .B1(n14225), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14228), .ZN(n14227) );
  INV_X1 U17359 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14385) );
  MUX2_X1 U17360 ( .A(n14385), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n15529), .Z(n14226) );
  OAI211_X1 U17361 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14228), .A(
        n14227), .B(n14226), .ZN(n14229) );
  XNOR2_X1 U17362 ( .A(n14229), .B(n14377), .ZN(n14381) );
  INV_X1 U17363 ( .A(n14230), .ZN(n14232) );
  INV_X1 U17364 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20568) );
  NOR2_X1 U17365 ( .A1(n15731), .A2(n20568), .ZN(n14373) );
  AOI21_X1 U17366 ( .B1(n19813), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14373), .ZN(n14231) );
  OAI21_X1 U17367 ( .B1(n15597), .B2(n14232), .A(n14231), .ZN(n14233) );
  AOI21_X1 U17368 ( .B1(n14234), .B2(n14290), .A(n14233), .ZN(n14235) );
  OAI21_X1 U17369 ( .B1(n19637), .B2(n14381), .A(n14235), .ZN(P1_U2971) );
  INV_X1 U17370 ( .A(n14236), .ZN(n14238) );
  XNOR2_X1 U17371 ( .A(n14239), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14390) );
  AOI22_X1 U17372 ( .A1(n19813), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        n19819), .B2(P1_REIP_REG_27__SCAN_IN), .ZN(n14240) );
  OAI21_X1 U17373 ( .B1(n15597), .B2(n14241), .A(n14240), .ZN(n14242) );
  AOI21_X1 U17374 ( .B1(n14243), .B2(n14290), .A(n14242), .ZN(n14244) );
  OAI21_X1 U17375 ( .B1(n19637), .B2(n14390), .A(n14244), .ZN(P1_U2972) );
  NOR2_X1 U17376 ( .A1(n15731), .A2(n20563), .ZN(n14393) );
  INV_X1 U17377 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14245) );
  NOR2_X1 U17378 ( .A1(n15603), .A2(n14245), .ZN(n14246) );
  AOI211_X1 U17379 ( .C1(n15600), .C2(n14247), .A(n14393), .B(n14246), .ZN(
        n14252) );
  OAI211_X1 U17380 ( .C1(n14342), .C2(n14223), .A(n14249), .B(n14248), .ZN(
        n14250) );
  XNOR2_X1 U17381 ( .A(n14250), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14391) );
  NAND2_X1 U17382 ( .A1(n14391), .A2(n19817), .ZN(n14251) );
  OAI211_X1 U17383 ( .C1(n14253), .C2(n19841), .A(n14252), .B(n14251), .ZN(
        P1_U2973) );
  OAI22_X1 U17384 ( .A1(n15603), .A2(n14254), .B1(n15731), .B2(n20561), .ZN(
        n14255) );
  AOI21_X1 U17385 ( .B1(n14256), .B2(n15600), .A(n14255), .ZN(n14263) );
  NOR3_X1 U17386 ( .A1(n14223), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14259) );
  NAND2_X1 U17387 ( .A1(n14257), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14266) );
  NOR2_X1 U17388 ( .A1(n14266), .A2(n15606), .ZN(n14258) );
  MUX2_X1 U17389 ( .A(n14259), .B(n14258), .S(n15529), .Z(n14261) );
  XNOR2_X1 U17390 ( .A(n14261), .B(n14260), .ZN(n15609) );
  NAND2_X1 U17391 ( .A1(n15609), .A2(n19817), .ZN(n14262) );
  OAI211_X1 U17392 ( .C1(n14264), .C2(n19841), .A(n14263), .B(n14262), .ZN(
        P1_U2974) );
  NAND2_X1 U17393 ( .A1(n14266), .A2(n14265), .ZN(n14267) );
  MUX2_X1 U17394 ( .A(n14267), .B(n14266), .S(n15529), .Z(n14268) );
  XNOR2_X1 U17395 ( .A(n14268), .B(n15606), .ZN(n14406) );
  INV_X1 U17396 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14271) );
  NAND2_X1 U17397 ( .A1(n15600), .A2(n14269), .ZN(n14270) );
  NAND2_X1 U17398 ( .A1(n19819), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14400) );
  OAI211_X1 U17399 ( .C1(n15603), .C2(n14271), .A(n14270), .B(n14400), .ZN(
        n14272) );
  AOI21_X1 U17400 ( .B1(n14273), .B2(n14290), .A(n14272), .ZN(n14274) );
  OAI21_X1 U17401 ( .B1(n19637), .B2(n14406), .A(n14274), .ZN(P1_U2975) );
  NAND2_X1 U17402 ( .A1(n14276), .A2(n14275), .ZN(n14278) );
  XNOR2_X1 U17403 ( .A(n14278), .B(n14277), .ZN(n15625) );
  INV_X1 U17404 ( .A(n15473), .ZN(n14282) );
  INV_X1 U17405 ( .A(n15476), .ZN(n14280) );
  AOI22_X1 U17406 ( .A1(n19813), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n19819), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n14279) );
  OAI21_X1 U17407 ( .B1(n15597), .B2(n14280), .A(n14279), .ZN(n14281) );
  AOI21_X1 U17408 ( .B1(n14282), .B2(n14290), .A(n14281), .ZN(n14283) );
  OAI21_X1 U17409 ( .B1(n19637), .B2(n15625), .A(n14283), .ZN(P1_U2977) );
  INV_X1 U17410 ( .A(n14284), .ZN(n15429) );
  NOR2_X1 U17411 ( .A1(n15429), .A2(n15430), .ZN(n14286) );
  MUX2_X1 U17412 ( .A(n14286), .B(n14285), .S(n14342), .Z(n14287) );
  XNOR2_X1 U17413 ( .A(n14287), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14419) );
  NAND2_X1 U17414 ( .A1(n15600), .A2(n15489), .ZN(n14288) );
  NAND2_X1 U17415 ( .A1(n19819), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14415) );
  OAI211_X1 U17416 ( .C1(n15603), .C2(n15499), .A(n14288), .B(n14415), .ZN(
        n14289) );
  AOI21_X1 U17417 ( .B1(n14291), .B2(n14290), .A(n14289), .ZN(n14292) );
  OAI21_X1 U17418 ( .B1(n19637), .B2(n14419), .A(n14292), .ZN(P1_U2979) );
  OAI21_X1 U17419 ( .B1(n14293), .B2(n15431), .A(n15429), .ZN(n15642) );
  AOI22_X1 U17420 ( .A1(n19813), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n19819), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14294) );
  OAI21_X1 U17421 ( .B1(n15597), .B2(n15502), .A(n14294), .ZN(n14295) );
  AOI21_X1 U17422 ( .B1(n15508), .B2(n14290), .A(n14295), .ZN(n14296) );
  OAI21_X1 U17423 ( .B1(n19637), .B2(n15642), .A(n14296), .ZN(P1_U2981) );
  NAND2_X1 U17424 ( .A1(n14297), .A2(n14298), .ZN(n14299) );
  NAND2_X1 U17425 ( .A1(n14299), .A2(n9645), .ZN(n14316) );
  AND2_X1 U17426 ( .A1(n15529), .A2(n14437), .ZN(n14300) );
  OR2_X1 U17427 ( .A1(n15529), .A2(n14437), .ZN(n14301) );
  AND2_X1 U17428 ( .A1(n14315), .A2(n14301), .ZN(n14302) );
  NAND2_X1 U17429 ( .A1(n14303), .A2(n14302), .ZN(n15562) );
  NOR2_X1 U17430 ( .A1(n15529), .A2(n14428), .ZN(n15560) );
  NOR2_X1 U17431 ( .A1(n15562), .A2(n15560), .ZN(n15553) );
  INV_X1 U17432 ( .A(n14304), .ZN(n15559) );
  NOR2_X1 U17433 ( .A1(n15553), .A2(n15559), .ZN(n14308) );
  INV_X1 U17434 ( .A(n15553), .ZN(n14306) );
  NAND2_X1 U17435 ( .A1(n14306), .A2(n14305), .ZN(n15550) );
  OAI21_X1 U17436 ( .B1(n14308), .B2(n14307), .A(n15550), .ZN(n14432) );
  INV_X1 U17437 ( .A(n14309), .ZN(n14311) );
  AOI22_X1 U17438 ( .A1(n19813), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n19819), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n14310) );
  OAI21_X1 U17439 ( .B1(n15597), .B2(n14311), .A(n14310), .ZN(n14312) );
  AOI21_X1 U17440 ( .B1(n14313), .B2(n14290), .A(n14312), .ZN(n14314) );
  OAI21_X1 U17441 ( .B1(n14432), .B2(n19637), .A(n14314), .ZN(P1_U2983) );
  NAND2_X1 U17442 ( .A1(n14316), .A2(n14315), .ZN(n14318) );
  XNOR2_X1 U17443 ( .A(n15529), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14317) );
  XNOR2_X1 U17444 ( .A(n14318), .B(n14317), .ZN(n14440) );
  NAND2_X1 U17445 ( .A1(n19819), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n14433) );
  NAND2_X1 U17446 ( .A1(n19813), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14319) );
  OAI211_X1 U17447 ( .C1(n15597), .C2(n14320), .A(n14433), .B(n14319), .ZN(
        n14321) );
  AOI21_X1 U17448 ( .B1(n14322), .B2(n14290), .A(n14321), .ZN(n14323) );
  OAI21_X1 U17449 ( .B1(n14440), .B2(n19637), .A(n14323), .ZN(P1_U2985) );
  INV_X1 U17450 ( .A(n14324), .ZN(n14325) );
  OR2_X1 U17451 ( .A1(n14297), .A2(n14325), .ZN(n14327) );
  NAND2_X1 U17452 ( .A1(n14327), .A2(n14326), .ZN(n15570) );
  NAND2_X1 U17453 ( .A1(n14328), .A2(n14329), .ZN(n15569) );
  NAND2_X1 U17454 ( .A1(n15567), .A2(n14329), .ZN(n14330) );
  XOR2_X1 U17455 ( .A(n14331), .B(n14330), .Z(n15664) );
  AOI22_X1 U17456 ( .A1(n19813), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n19819), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14334) );
  NAND2_X1 U17457 ( .A1(n15600), .A2(n14332), .ZN(n14333) );
  OAI211_X1 U17458 ( .C1(n14335), .C2(n19841), .A(n14334), .B(n14333), .ZN(
        n14336) );
  AOI21_X1 U17459 ( .B1(n15664), .B2(n19817), .A(n14336), .ZN(n14337) );
  INV_X1 U17460 ( .A(n14337), .ZN(P1_U2986) );
  XNOR2_X1 U17461 ( .A(n14297), .B(n14341), .ZN(n14340) );
  NAND2_X1 U17462 ( .A1(n14338), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14339) );
  MUX2_X1 U17463 ( .A(n14340), .B(n14339), .S(n14342), .Z(n14344) );
  INV_X1 U17464 ( .A(n14338), .ZN(n14343) );
  NAND3_X1 U17465 ( .A1(n14343), .A2(n14342), .A3(n14341), .ZN(n15576) );
  NAND2_X1 U17466 ( .A1(n14344), .A2(n15576), .ZN(n15703) );
  NAND2_X1 U17467 ( .A1(n15703), .A2(n19817), .ZN(n14348) );
  NOR2_X1 U17468 ( .A1(n15731), .A2(n20534), .ZN(n15698) );
  NOR2_X1 U17469 ( .A1(n15597), .A2(n14345), .ZN(n14346) );
  AOI211_X1 U17470 ( .C1(n19813), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15698), .B(n14346), .ZN(n14347) );
  OAI211_X1 U17471 ( .C1(n19841), .C2(n14349), .A(n14348), .B(n14347), .ZN(
        P1_U2989) );
  NOR2_X1 U17472 ( .A1(n14350), .A2(n15733), .ZN(n14358) );
  NOR3_X1 U17473 ( .A1(n14352), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14351), .ZN(n14357) );
  AND3_X1 U17474 ( .A1(n14354), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14353), .ZN(n14355) );
  NOR4_X1 U17475 ( .A1(n14358), .A2(n14357), .A3(n14356), .A4(n14355), .ZN(
        n14359) );
  OAI21_X1 U17476 ( .B1(n14360), .B2(n15685), .A(n14359), .ZN(P1_U3000) );
  INV_X1 U17477 ( .A(n14361), .ZN(n14363) );
  AOI21_X1 U17478 ( .B1(n14363), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14362), .ZN(n14367) );
  INV_X1 U17479 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14364) );
  NAND3_X1 U17480 ( .A1(n14383), .A2(n14365), .A3(n14364), .ZN(n14366) );
  OAI211_X1 U17481 ( .C1(n14368), .C2(n15733), .A(n14367), .B(n14366), .ZN(
        n14369) );
  AOI21_X1 U17482 ( .B1(n14370), .B2(n19824), .A(n14369), .ZN(n14371) );
  INV_X1 U17483 ( .A(n14371), .ZN(P1_U3002) );
  AOI21_X1 U17484 ( .B1(n14377), .B2(n14385), .A(n14372), .ZN(n14375) );
  AOI21_X1 U17485 ( .B1(n14375), .B2(n14374), .A(n14373), .ZN(n14376) );
  OAI21_X1 U17486 ( .B1(n14386), .B2(n14377), .A(n14376), .ZN(n14378) );
  AOI21_X1 U17487 ( .B1(n14379), .B2(n19826), .A(n14378), .ZN(n14380) );
  OAI21_X1 U17488 ( .B1(n14381), .B2(n15685), .A(n14380), .ZN(P1_U3003) );
  NOR2_X1 U17489 ( .A1(n15731), .A2(n20565), .ZN(n14382) );
  AOI21_X1 U17490 ( .B1(n14385), .B2(n14383), .A(n14382), .ZN(n14384) );
  OAI21_X1 U17491 ( .B1(n14386), .B2(n14385), .A(n14384), .ZN(n14387) );
  AOI21_X1 U17492 ( .B1(n14388), .B2(n19826), .A(n14387), .ZN(n14389) );
  OAI21_X1 U17493 ( .B1(n14390), .B2(n15685), .A(n14389), .ZN(P1_U3004) );
  INV_X1 U17494 ( .A(n14391), .ZN(n14397) );
  AOI22_X1 U17495 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15610), .B1(
        n14392), .B2(n20759), .ZN(n14396) );
  AOI21_X1 U17496 ( .B1(n14394), .B2(n19826), .A(n14393), .ZN(n14395) );
  OAI211_X1 U17497 ( .C1(n14397), .C2(n15685), .A(n14396), .B(n14395), .ZN(
        P1_U3005) );
  OAI21_X1 U17498 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14399), .A(
        n14398), .ZN(n14404) );
  NOR3_X1 U17499 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n20803), .A3(
        n15605), .ZN(n14403) );
  OAI21_X1 U17500 ( .B1(n14401), .B2(n15733), .A(n14400), .ZN(n14402) );
  AOI211_X1 U17501 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n14404), .A(
        n14403), .B(n14402), .ZN(n14405) );
  OAI21_X1 U17502 ( .B1(n14406), .B2(n15685), .A(n14405), .ZN(P1_U3007) );
  INV_X1 U17503 ( .A(n14407), .ZN(n14410) );
  AOI21_X1 U17504 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n14408), .A(
        n15674), .ZN(n14409) );
  AOI211_X1 U17505 ( .C1(n14411), .C2(n14410), .A(n14409), .B(n15676), .ZN(
        n15631) );
  OAI21_X1 U17506 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n14412), .A(
        n15631), .ZN(n14417) );
  NOR2_X1 U17507 ( .A1(n15637), .A2(n15430), .ZN(n14413) );
  INV_X1 U17508 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15434) );
  NAND2_X1 U17509 ( .A1(n14413), .A2(n15434), .ZN(n14414) );
  OAI211_X1 U17510 ( .C1(n15492), .C2(n15733), .A(n14415), .B(n14414), .ZN(
        n14416) );
  AOI21_X1 U17511 ( .B1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n14417), .A(
        n14416), .ZN(n14418) );
  OAI21_X1 U17512 ( .B1(n14419), .B2(n15685), .A(n14418), .ZN(P1_U3011) );
  NOR3_X1 U17513 ( .A1(n15689), .A2(n14420), .A3(n12575), .ZN(n14438) );
  NAND2_X1 U17514 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n14438), .ZN(
        n15648) );
  NOR2_X1 U17515 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15648), .ZN(
        n15658) );
  INV_X1 U17516 ( .A(n14420), .ZN(n14424) );
  OAI221_X1 U17517 ( .B1(n12575), .B2(n15720), .C1(n12575), .C2(n14421), .A(
        n15722), .ZN(n14422) );
  OAI211_X1 U17518 ( .C1(n14424), .C2(n19829), .A(n14423), .B(n14422), .ZN(
        n15665) );
  AOI21_X1 U17519 ( .B1(n14437), .B2(n15722), .A(n15665), .ZN(n15639) );
  INV_X1 U17520 ( .A(n15639), .ZN(n15659) );
  OAI21_X1 U17521 ( .B1(n15658), .B2(n15659), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14426) );
  OR2_X1 U17522 ( .A1(n15731), .A2(n20545), .ZN(n14425) );
  OAI211_X1 U17523 ( .C1(n15733), .C2(n14427), .A(n14426), .B(n14425), .ZN(
        n14430) );
  NOR3_X1 U17524 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n14428), .A3(
        n15648), .ZN(n14429) );
  NOR2_X1 U17525 ( .A1(n14430), .A2(n14429), .ZN(n14431) );
  OAI21_X1 U17526 ( .B1(n14432), .B2(n15685), .A(n14431), .ZN(P1_U3015) );
  NAND2_X1 U17527 ( .A1(n15665), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14434) );
  OAI211_X1 U17528 ( .C1(n15733), .C2(n14435), .A(n14434), .B(n14433), .ZN(
        n14436) );
  AOI21_X1 U17529 ( .B1(n14438), .B2(n14437), .A(n14436), .ZN(n14439) );
  OAI21_X1 U17530 ( .B1(n14440), .B2(n15685), .A(n14439), .ZN(P1_U3017) );
  AOI21_X1 U17531 ( .B1(n9635), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20442), 
        .ZN(n19969) );
  OAI21_X1 U17532 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n9635), .A(n19969), 
        .ZN(n14441) );
  OAI21_X1 U17533 ( .B1(n14445), .B2(n20292), .A(n14441), .ZN(n14442) );
  MUX2_X1 U17534 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14442), .S(
        n19837), .Z(P1_U3477) );
  INV_X1 U17535 ( .A(n19969), .ZN(n20441) );
  MUX2_X1 U17536 ( .A(n20441), .B(n14443), .S(n13225), .Z(n14444) );
  OAI21_X1 U17537 ( .B1(n14445), .B2(n13187), .A(n14444), .ZN(n14446) );
  MUX2_X1 U17538 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14446), .S(
        n19837), .Z(P1_U3476) );
  INV_X1 U17539 ( .A(n20595), .ZN(n20591) );
  INV_X1 U17540 ( .A(n14447), .ZN(n14449) );
  INV_X1 U17541 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14448) );
  AOI22_X1 U17542 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n13075), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14448), .ZN(n20594) );
  NAND2_X1 U17543 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20604) );
  OAI222_X1 U17544 ( .A1(n14450), .A2(n20597), .B1(n20591), .B2(n14449), .C1(
        n20594), .C2(n20604), .ZN(n14451) );
  MUX2_X1 U17545 ( .A(n14451), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n20605), .Z(P1_U3472) );
  OR2_X1 U17546 ( .A1(n14452), .A2(n19510), .ZN(n16098) );
  INV_X1 U17547 ( .A(n16098), .ZN(n14453) );
  AOI21_X1 U17548 ( .B1(n19294), .B2(n14454), .A(n14453), .ZN(n14456) );
  OAI21_X1 U17549 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .A(n18640), .ZN(n16114) );
  OAI21_X1 U17550 ( .B1(n19520), .B2(n19606), .A(n16114), .ZN(n14455) );
  OAI21_X1 U17551 ( .B1(n14456), .B2(n18640), .A(n14455), .ZN(n14459) );
  NOR4_X1 U17552 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19520), .A3(n19606), 
        .A4(n11065), .ZN(n14457) );
  AOI211_X1 U17553 ( .C1(n19494), .C2(n19604), .A(n14457), .B(n18642), .ZN(
        n14458) );
  MUX2_X1 U17554 ( .A(n14459), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n14458), 
        .Z(P2_U3610) );
  AOI21_X1 U17555 ( .B1(n14461), .B2(n14624), .A(n14460), .ZN(n14473) );
  AOI22_X1 U17556 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n9607), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n18669), .ZN(n14462) );
  OAI21_X1 U17557 ( .B1(n14463), .B2(n18795), .A(n14462), .ZN(n14472) );
  NOR2_X1 U17558 ( .A1(n12642), .A2(n14464), .ZN(n14465) );
  OR2_X1 U17559 ( .A1(n14467), .A2(n14466), .ZN(n14469) );
  AOI22_X1 U17560 ( .A1(n14775), .A2(n15802), .B1(P2_EBX_REG_28__SCAN_IN), 
        .B2(n18819), .ZN(n14470) );
  OAI21_X1 U17561 ( .B1(n14774), .B2(n18789), .A(n14470), .ZN(n14471) );
  AOI211_X1 U17562 ( .C1(n14473), .C2(n19499), .A(n14472), .B(n14471), .ZN(
        n14474) );
  INV_X1 U17563 ( .A(n14474), .ZN(P2_U2827) );
  AOI211_X1 U17564 ( .C1(n14651), .C2(n14476), .A(n14475), .B(n18779), .ZN(
        n14477) );
  INV_X1 U17565 ( .A(n14477), .ZN(n14487) );
  OR2_X1 U17566 ( .A1(n14552), .A2(n14478), .ZN(n14479) );
  AND2_X1 U17567 ( .A1(n14479), .A2(n14538), .ZN(n14813) );
  NAND2_X1 U17568 ( .A1(n14480), .A2(n14481), .ZN(n14482) );
  NAND2_X1 U17569 ( .A1(n14571), .A2(n14482), .ZN(n14811) );
  NAND2_X1 U17570 ( .A1(n18669), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n14484) );
  AOI22_X1 U17571 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n9607), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n18819), .ZN(n14483) );
  OAI211_X1 U17572 ( .C1(n18812), .C2(n14811), .A(n14484), .B(n14483), .ZN(
        n14485) );
  AOI21_X1 U17573 ( .B1(n14813), .B2(n18814), .A(n14485), .ZN(n14486) );
  OAI211_X1 U17574 ( .C1(n18795), .C2(n14488), .A(n14487), .B(n14486), .ZN(
        P2_U2830) );
  AOI211_X1 U17575 ( .C1(n14491), .C2(n14490), .A(n14489), .B(n18779), .ZN(
        n14505) );
  AOI22_X1 U17576 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n9607), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18669), .ZN(n14493) );
  NAND2_X1 U17577 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n18819), .ZN(n14492) );
  OAI211_X1 U17578 ( .C1(n18795), .C2(n14494), .A(n14493), .B(n14492), .ZN(
        n14504) );
  NAND2_X1 U17579 ( .A1(n14496), .A2(n14495), .ZN(n14497) );
  NAND2_X1 U17580 ( .A1(n14498), .A2(n14497), .ZN(n15822) );
  OR2_X1 U17581 ( .A1(n14500), .A2(n14499), .ZN(n14501) );
  AND2_X1 U17582 ( .A1(n9703), .A2(n14501), .ZN(n15835) );
  INV_X1 U17583 ( .A(n15835), .ZN(n14502) );
  OAI22_X1 U17584 ( .A1(n15822), .A2(n18789), .B1(n14502), .B2(n18812), .ZN(
        n14503) );
  OR3_X1 U17585 ( .A1(n14505), .A2(n14504), .A3(n14503), .ZN(P2_U2835) );
  AOI211_X1 U17586 ( .C1(n14713), .C2(n14507), .A(n14506), .B(n18779), .ZN(
        n14513) );
  AOI21_X1 U17587 ( .B1(P2_REIP_REG_19__SCAN_IN), .B2(n18669), .A(n18933), 
        .ZN(n14509) );
  AOI22_X1 U17588 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n9607), .B1(
        P2_EBX_REG_19__SCAN_IN), .B2(n18819), .ZN(n14508) );
  OAI211_X1 U17589 ( .C1(n14510), .C2(n18795), .A(n14509), .B(n14508), .ZN(
        n14512) );
  OAI22_X1 U17590 ( .A1(n14880), .A2(n18789), .B1(n14879), .B2(n18812), .ZN(
        n14511) );
  OR3_X1 U17591 ( .A1(n14513), .A2(n14512), .A3(n14511), .ZN(P2_U2836) );
  INV_X1 U17592 ( .A(n13912), .ZN(n14518) );
  NAND3_X1 U17593 ( .A1(n14518), .A2(n18871), .A3(n14517), .ZN(n14520) );
  NAND2_X1 U17594 ( .A1(n18875), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14519) );
  OAI211_X1 U17595 ( .C1(n18875), .C2(n15780), .A(n14520), .B(n14519), .ZN(
        P2_U2858) );
  NOR2_X1 U17596 ( .A1(n14522), .A2(n14521), .ZN(n14524) );
  XNOR2_X1 U17597 ( .A(n14524), .B(n14523), .ZN(n14558) );
  NAND2_X1 U17598 ( .A1(n14558), .A2(n18871), .ZN(n14526) );
  NAND2_X1 U17599 ( .A1(n18875), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14525) );
  OAI211_X1 U17600 ( .C1(n18875), .C2(n14774), .A(n14526), .B(n14525), .ZN(
        P2_U2859) );
  AOI21_X1 U17601 ( .B1(n14529), .B2(n14528), .A(n14527), .ZN(n14530) );
  INV_X1 U17602 ( .A(n14530), .ZN(n14568) );
  NAND2_X1 U17603 ( .A1(n18875), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14532) );
  NAND2_X1 U17604 ( .A1(n14789), .A2(n18859), .ZN(n14531) );
  OAI211_X1 U17605 ( .C1(n14568), .C2(n18865), .A(n14532), .B(n14531), .ZN(
        P2_U2860) );
  OAI21_X1 U17606 ( .B1(n14535), .B2(n14534), .A(n14533), .ZN(n14577) );
  NAND2_X1 U17607 ( .A1(n18875), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14541) );
  INV_X1 U17608 ( .A(n14536), .ZN(n14537) );
  AOI21_X1 U17609 ( .B1(n14539), .B2(n14538), .A(n14537), .ZN(n15788) );
  NAND2_X1 U17610 ( .A1(n15788), .A2(n18859), .ZN(n14540) );
  OAI211_X1 U17611 ( .C1(n14577), .C2(n18865), .A(n14541), .B(n14540), .ZN(
        P2_U2861) );
  OAI21_X1 U17612 ( .B1(n14544), .B2(n14543), .A(n14542), .ZN(n14583) );
  INV_X1 U17613 ( .A(n14813), .ZN(n14648) );
  MUX2_X1 U17614 ( .A(n14648), .B(n20797), .S(n18875), .Z(n14545) );
  OAI21_X1 U17615 ( .B1(n14583), .B2(n18865), .A(n14545), .ZN(P2_U2862) );
  AOI21_X1 U17616 ( .B1(n14547), .B2(n14546), .A(n9702), .ZN(n14548) );
  XOR2_X1 U17617 ( .A(n14549), .B(n14548), .Z(n14590) );
  NOR2_X1 U17618 ( .A1(n12670), .A2(n14550), .ZN(n14551) );
  OR2_X1 U17619 ( .A1(n14552), .A2(n14551), .ZN(n15848) );
  NOR2_X1 U17620 ( .A1(n15848), .A2(n18875), .ZN(n14553) );
  AOI21_X1 U17621 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n18875), .A(n14553), .ZN(
        n14554) );
  OAI21_X1 U17622 ( .B1(n14590), .B2(n18865), .A(n14554), .ZN(P2_U2863) );
  MUX2_X1 U17623 ( .A(n14856), .B(n14555), .S(n18875), .Z(n14556) );
  OAI21_X1 U17624 ( .B1(n14557), .B2(n18865), .A(n14556), .ZN(P2_U2866) );
  NAND2_X1 U17625 ( .A1(n14558), .A2(n18885), .ZN(n14562) );
  AOI22_X1 U17626 ( .A1(n18880), .A2(n18890), .B1(n18893), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n14561) );
  AOI22_X1 U17627 ( .A1(n18882), .A2(BUF1_REG_28__SCAN_IN), .B1(n18881), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n14560) );
  NAND2_X1 U17628 ( .A1(n14775), .A2(n18884), .ZN(n14559) );
  NAND4_X1 U17629 ( .A1(n14562), .A2(n14561), .A3(n14560), .A4(n14559), .ZN(
        P2_U2891) );
  OAI22_X1 U17630 ( .A1(n14792), .A2(n14585), .B1(n14596), .B2(n14563), .ZN(
        n14564) );
  AOI21_X1 U17631 ( .B1(n18880), .B2(n14565), .A(n14564), .ZN(n14567) );
  AOI22_X1 U17632 ( .A1(n18882), .A2(BUF1_REG_27__SCAN_IN), .B1(n18881), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n14566) );
  OAI211_X1 U17633 ( .C1(n14568), .C2(n14601), .A(n14567), .B(n14566), .ZN(
        P2_U2892) );
  INV_X1 U17634 ( .A(n14569), .ZN(n14570) );
  AOI21_X1 U17635 ( .B1(n14572), .B2(n14571), .A(n14570), .ZN(n15797) );
  INV_X1 U17636 ( .A(n15797), .ZN(n14573) );
  OAI22_X1 U17637 ( .A1(n14573), .A2(n14585), .B1(n14596), .B2(n12816), .ZN(
        n14574) );
  AOI21_X1 U17638 ( .B1(n18880), .B2(n18894), .A(n14574), .ZN(n14576) );
  AOI22_X1 U17639 ( .A1(n18882), .A2(BUF1_REG_26__SCAN_IN), .B1(n18881), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n14575) );
  OAI211_X1 U17640 ( .C1(n14577), .C2(n14601), .A(n14576), .B(n14575), .ZN(
        P2_U2893) );
  OAI22_X1 U17641 ( .A1(n14585), .A2(n14811), .B1(n14596), .B2(n14578), .ZN(
        n14579) );
  AOI21_X1 U17642 ( .B1(n18880), .B2(n14580), .A(n14579), .ZN(n14582) );
  AOI22_X1 U17643 ( .A1(n18882), .A2(BUF1_REG_25__SCAN_IN), .B1(n18881), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n14581) );
  OAI211_X1 U17644 ( .C1(n14583), .C2(n14601), .A(n14582), .B(n14581), .ZN(
        P2_U2894) );
  OAI21_X1 U17645 ( .B1(n12674), .B2(n14584), .A(n14480), .ZN(n14827) );
  OAI22_X1 U17646 ( .A1(n14585), .A2(n14827), .B1(n14596), .B2(n12818), .ZN(
        n14586) );
  AOI21_X1 U17647 ( .B1(n18880), .B2(n14587), .A(n14586), .ZN(n14589) );
  AOI22_X1 U17648 ( .A1(n18882), .A2(BUF1_REG_24__SCAN_IN), .B1(n18881), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n14588) );
  OAI211_X1 U17649 ( .C1(n14590), .C2(n14601), .A(n14589), .B(n14588), .ZN(
        P2_U2895) );
  AOI21_X1 U17650 ( .B1(n14593), .B2(n14592), .A(n14591), .ZN(n15814) );
  INV_X1 U17651 ( .A(n15814), .ZN(n14602) );
  INV_X1 U17652 ( .A(n14594), .ZN(n14841) );
  OAI22_X1 U17653 ( .A1(n14597), .A2(n18983), .B1(n14596), .B2(n14595), .ZN(
        n14598) );
  AOI21_X1 U17654 ( .B1(n18884), .B2(n14841), .A(n14598), .ZN(n14600) );
  AOI22_X1 U17655 ( .A1(n18882), .A2(BUF1_REG_23__SCAN_IN), .B1(n18881), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n14599) );
  OAI211_X1 U17656 ( .C1(n14602), .C2(n14601), .A(n14600), .B(n14599), .ZN(
        P2_U2896) );
  NOR2_X1 U17657 ( .A1(n14605), .A2(n14604), .ZN(n14606) );
  XNOR2_X1 U17658 ( .A(n14603), .B(n14606), .ZN(n14764) );
  NAND2_X1 U17659 ( .A1(n14764), .A2(n18936), .ZN(n14612) );
  AOI21_X1 U17660 ( .B1(n14607), .B2(n14772), .A(n14608), .ZN(n14769) );
  NAND2_X1 U17661 ( .A1(n18939), .A2(n14769), .ZN(n14609) );
  NAND2_X1 U17662 ( .A1(n18933), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n14765) );
  OAI211_X1 U17663 ( .C1(n15957), .C2(n15775), .A(n14609), .B(n14765), .ZN(
        n14610) );
  AOI21_X1 U17664 ( .B1(n15948), .B2(n15773), .A(n14610), .ZN(n14611) );
  OAI211_X1 U17665 ( .C1(n15859), .C2(n15780), .A(n14612), .B(n14611), .ZN(
        P2_U2985) );
  XNOR2_X1 U17666 ( .A(n14615), .B(n14617), .ZN(n14626) );
  INV_X1 U17667 ( .A(n14615), .ZN(n14616) );
  AOI22_X1 U17668 ( .A1(n14626), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n14617), .B2(n14616), .ZN(n14620) );
  XNOR2_X1 U17669 ( .A(n14618), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14619) );
  XNOR2_X1 U17670 ( .A(n14620), .B(n14619), .ZN(n14787) );
  OAI21_X1 U17671 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n9682), .A(
        n14607), .ZN(n14778) );
  NAND2_X1 U17672 ( .A1(n18934), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14621) );
  NAND2_X1 U17673 ( .A1(n18933), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n14776) );
  OAI211_X1 U17674 ( .C1(n15941), .C2(n14778), .A(n14621), .B(n14776), .ZN(
        n14623) );
  NOR2_X1 U17675 ( .A1(n14774), .A2(n15859), .ZN(n14622) );
  AOI211_X1 U17676 ( .C1(n15948), .C2(n14624), .A(n14623), .B(n14622), .ZN(
        n14625) );
  OAI21_X1 U17677 ( .B1(n14787), .B2(n15942), .A(n14625), .ZN(P2_U2986) );
  XNOR2_X1 U17678 ( .A(n14626), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14800) );
  NAND2_X1 U17679 ( .A1(n15948), .A2(n14627), .ZN(n14628) );
  OR2_X1 U17680 ( .A1(n11181), .A2(n20763), .ZN(n14790) );
  OAI211_X1 U17681 ( .C1(n15957), .C2(n14629), .A(n14628), .B(n14790), .ZN(
        n14630) );
  AOI21_X1 U17682 ( .B1(n14789), .B2(n18938), .A(n14630), .ZN(n14632) );
  AOI21_X1 U17683 ( .B1(n14640), .B2(n14779), .A(n9682), .ZN(n14797) );
  NAND2_X1 U17684 ( .A1(n14797), .A2(n18939), .ZN(n14631) );
  OAI211_X1 U17685 ( .C1(n14800), .C2(n15942), .A(n14632), .B(n14631), .ZN(
        P2_U2987) );
  AOI21_X1 U17686 ( .B1(n14633), .B2(n14645), .A(n14644), .ZN(n14634) );
  XOR2_X1 U17687 ( .A(n14635), .B(n14634), .Z(n14810) );
  NOR2_X1 U17688 ( .A1(n11181), .A2(n15790), .ZN(n14801) );
  AOI21_X1 U17689 ( .B1(n18934), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14801), .ZN(n14636) );
  OAI21_X1 U17690 ( .B1(n18944), .B2(n14637), .A(n14636), .ZN(n14642) );
  NAND2_X1 U17691 ( .A1(n14638), .A2(n14804), .ZN(n14639) );
  NAND2_X1 U17692 ( .A1(n14640), .A2(n14639), .ZN(n14805) );
  NOR2_X1 U17693 ( .A1(n14805), .A2(n15941), .ZN(n14641) );
  AOI211_X1 U17694 ( .C1(n15788), .C2(n18938), .A(n14642), .B(n14641), .ZN(
        n14643) );
  OAI21_X1 U17695 ( .B1(n14810), .B2(n15942), .A(n14643), .ZN(P2_U2988) );
  NAND2_X1 U17696 ( .A1(n10717), .A2(n14645), .ZN(n14646) );
  XNOR2_X1 U17697 ( .A(n14633), .B(n14646), .ZN(n14822) );
  OAI22_X1 U17698 ( .A1(n15957), .A2(n14647), .B1(n19560), .B2(n11181), .ZN(
        n14650) );
  NOR2_X1 U17699 ( .A1(n14648), .A2(n15859), .ZN(n14649) );
  AOI211_X1 U17700 ( .C1(n15948), .C2(n14651), .A(n14650), .B(n14649), .ZN(
        n14654) );
  INV_X1 U17701 ( .A(n15846), .ZN(n14652) );
  NAND2_X1 U17702 ( .A1(n14652), .A2(n14817), .ZN(n14819) );
  NAND3_X1 U17703 ( .A1(n14819), .A2(n18939), .A3(n14638), .ZN(n14653) );
  OAI211_X1 U17704 ( .C1(n14822), .C2(n15942), .A(n14654), .B(n14653), .ZN(
        P2_U2989) );
  INV_X1 U17705 ( .A(n14826), .ZN(n14655) );
  OAI21_X1 U17706 ( .B1(n14656), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14655), .ZN(n14848) );
  XOR2_X1 U17707 ( .A(n14658), .B(n14657), .Z(n14846) );
  NOR2_X1 U17708 ( .A1(n11181), .A2(n19556), .ZN(n14840) );
  NOR2_X1 U17709 ( .A1(n15957), .A2(n14659), .ZN(n14660) );
  AOI211_X1 U17710 ( .C1(n14661), .C2(n15948), .A(n14840), .B(n14660), .ZN(
        n14662) );
  OAI21_X1 U17711 ( .B1(n15859), .B2(n15816), .A(n14662), .ZN(n14663) );
  AOI21_X1 U17712 ( .B1(n14846), .B2(n18936), .A(n14663), .ZN(n14664) );
  OAI21_X1 U17713 ( .B1(n14848), .B2(n15941), .A(n14664), .ZN(P2_U2991) );
  INV_X1 U17714 ( .A(n14666), .ZN(n14745) );
  NAND2_X1 U17715 ( .A1(n14665), .A2(n14745), .ZN(n14936) );
  INV_X1 U17716 ( .A(n14667), .ZN(n14735) );
  NAND2_X1 U17717 ( .A1(n14737), .A2(n14735), .ZN(n14668) );
  INV_X1 U17718 ( .A(n14669), .ZN(n14723) );
  INV_X1 U17719 ( .A(n14670), .ZN(n14671) );
  NAND2_X1 U17720 ( .A1(n14673), .A2(n14672), .ZN(n14716) );
  NAND2_X1 U17721 ( .A1(n14674), .A2(n14673), .ZN(n14888) );
  INV_X1 U17722 ( .A(n14887), .ZN(n14675) );
  INV_X1 U17723 ( .A(n14676), .ZN(n14691) );
  INV_X1 U17724 ( .A(n14678), .ZN(n14680) );
  NOR2_X1 U17725 ( .A1(n14680), .A2(n14679), .ZN(n14681) );
  AOI21_X1 U17726 ( .B1(n14858), .B2(n14695), .A(n14682), .ZN(n14849) );
  NOR2_X1 U17727 ( .A1(n11181), .A2(n19553), .ZN(n14852) );
  NOR2_X1 U17728 ( .A1(n15957), .A2(n14683), .ZN(n14684) );
  AOI211_X1 U17729 ( .C1(n14685), .C2(n15948), .A(n14852), .B(n14684), .ZN(
        n14686) );
  OAI21_X1 U17730 ( .B1(n15859), .B2(n14856), .A(n14686), .ZN(n14687) );
  AOI21_X1 U17731 ( .B1(n14849), .B2(n18939), .A(n14687), .ZN(n14688) );
  OAI21_X1 U17732 ( .B1(n14862), .B2(n15942), .A(n14688), .ZN(P2_U2993) );
  NAND2_X1 U17733 ( .A1(n9688), .A2(n14689), .ZN(n14693) );
  NAND2_X1 U17734 ( .A1(n14691), .A2(n14690), .ZN(n14692) );
  XNOR2_X1 U17735 ( .A(n14693), .B(n14692), .ZN(n14873) );
  INV_X1 U17736 ( .A(n14695), .ZN(n14696) );
  AOI21_X1 U17737 ( .B1(n14697), .B2(n14704), .A(n14696), .ZN(n14871) );
  NOR2_X1 U17738 ( .A1(n11181), .A2(n19551), .ZN(n14864) );
  NOR2_X1 U17739 ( .A1(n14698), .A2(n18944), .ZN(n14699) );
  AOI211_X1 U17740 ( .C1(n18934), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n14864), .B(n14699), .ZN(n14700) );
  OAI21_X1 U17741 ( .B1(n15859), .B2(n15822), .A(n14700), .ZN(n14701) );
  AOI21_X1 U17742 ( .B1(n14871), .B2(n18939), .A(n14701), .ZN(n14702) );
  OAI21_X1 U17743 ( .B1(n15942), .B2(n14873), .A(n14702), .ZN(P2_U2994) );
  NOR2_X1 U17744 ( .A1(n14886), .A2(n14703), .ZN(n14705) );
  OAI21_X1 U17745 ( .B1(n14705), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n14704), .ZN(n14875) );
  INV_X1 U17746 ( .A(n14890), .ZN(n14706) );
  NAND2_X1 U17747 ( .A1(n14891), .A2(n14706), .ZN(n14709) );
  NOR2_X1 U17748 ( .A1(n14707), .A2(n9639), .ZN(n14708) );
  XNOR2_X1 U17749 ( .A(n14709), .B(n14708), .ZN(n14874) );
  NAND2_X1 U17750 ( .A1(n14874), .A2(n18936), .ZN(n14715) );
  OAI22_X1 U17751 ( .A1(n15957), .A2(n14710), .B1(n19549), .B2(n11181), .ZN(
        n14712) );
  NOR2_X1 U17752 ( .A1(n14880), .A2(n15859), .ZN(n14711) );
  AOI211_X1 U17753 ( .C1(n15948), .C2(n14713), .A(n14712), .B(n14711), .ZN(
        n14714) );
  OAI211_X1 U17754 ( .C1(n15941), .C2(n14875), .A(n14715), .B(n14714), .ZN(
        P2_U2995) );
  XNOR2_X1 U17755 ( .A(n14717), .B(n14716), .ZN(n14918) );
  AOI22_X1 U17756 ( .A1(n18934), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n15948), .B2(n18682), .ZN(n14718) );
  OR2_X1 U17757 ( .A1(n11181), .A2(n19545), .ZN(n14911) );
  OAI211_X1 U17758 ( .C1(n15859), .C2(n18683), .A(n14718), .B(n14911), .ZN(
        n14721) );
  INV_X1 U17759 ( .A(n14886), .ZN(n14719) );
  AOI211_X1 U17760 ( .C1(n14920), .C2(n9637), .A(n15941), .B(n14719), .ZN(
        n14720) );
  AOI211_X1 U17761 ( .C1(n18936), .C2(n14918), .A(n14721), .B(n14720), .ZN(
        n14722) );
  INV_X1 U17762 ( .A(n14722), .ZN(P2_U2997) );
  XNOR2_X1 U17763 ( .A(n14724), .B(n14723), .ZN(n14931) );
  NOR2_X1 U17764 ( .A1(n14912), .A2(n15962), .ZN(n14725) );
  OAI211_X1 U17765 ( .C1(n14725), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n18939), .B(n9637), .ZN(n14733) );
  NAND2_X1 U17766 ( .A1(n14727), .A2(n14726), .ZN(n14728) );
  NAND2_X1 U17767 ( .A1(n14729), .A2(n14728), .ZN(n18836) );
  INV_X1 U17768 ( .A(n18836), .ZN(n14922) );
  NOR2_X1 U17769 ( .A1(n11108), .A2(n16010), .ZN(n14731) );
  INV_X1 U17770 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18695) );
  OAI22_X1 U17771 ( .A1(n15957), .A2(n18695), .B1(n18944), .B2(n18691), .ZN(
        n14730) );
  AOI211_X1 U17772 ( .C1(n14922), .C2(n18938), .A(n14731), .B(n14730), .ZN(
        n14732) );
  OAI211_X1 U17773 ( .C1(n14931), .C2(n15942), .A(n14733), .B(n14732), .ZN(
        P2_U2998) );
  XNOR2_X1 U17774 ( .A(n14939), .B(n15962), .ZN(n15964) );
  NAND2_X1 U17775 ( .A1(n14735), .A2(n14734), .ZN(n14736) );
  XNOR2_X1 U17776 ( .A(n14737), .B(n14736), .ZN(n15967) );
  AOI22_X1 U17777 ( .A1(n18934), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n15948), .B2(n18704), .ZN(n14739) );
  AOI22_X1 U17778 ( .A1(n18708), .A2(n18938), .B1(n18933), .B2(
        P2_REIP_REG_15__SCAN_IN), .ZN(n14738) );
  OAI211_X1 U17779 ( .C1(n15967), .C2(n15942), .A(n14739), .B(n14738), .ZN(
        n14740) );
  AOI21_X1 U17780 ( .B1(n18939), .B2(n15964), .A(n14740), .ZN(n14741) );
  INV_X1 U17781 ( .A(n14741), .ZN(P2_U2999) );
  OAI21_X1 U17782 ( .B1(n9608), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n14937), .ZN(n14967) );
  AND2_X1 U17783 ( .A1(n14743), .A2(n14742), .ZN(n14747) );
  NAND2_X1 U17784 ( .A1(n14745), .A2(n14744), .ZN(n14746) );
  XNOR2_X1 U17785 ( .A(n14747), .B(n14746), .ZN(n14965) );
  NAND2_X1 U17786 ( .A1(n18938), .A2(n14961), .ZN(n14750) );
  AOI22_X1 U17787 ( .A1(n18934), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n15948), .B2(n14748), .ZN(n14749) );
  OAI211_X1 U17788 ( .C1(n11098), .C2(n11181), .A(n14750), .B(n14749), .ZN(
        n14751) );
  AOI21_X1 U17789 ( .B1(n14965), .B2(n18936), .A(n14751), .ZN(n14752) );
  OAI21_X1 U17790 ( .B1(n14967), .B2(n15941), .A(n14752), .ZN(P2_U3001) );
  INV_X1 U17791 ( .A(n14753), .ZN(n14762) );
  NAND2_X1 U17792 ( .A1(n14754), .A2(n16063), .ZN(n14760) );
  OAI211_X1 U17793 ( .C1(n14762), .C2(n14761), .A(n14760), .B(n9684), .ZN(
        P2_U3016) );
  INV_X1 U17794 ( .A(n14780), .ZN(n14763) );
  NAND2_X1 U17795 ( .A1(n14763), .A2(n14779), .ZN(n14793) );
  NAND2_X1 U17796 ( .A1(n14793), .A2(n14788), .ZN(n14784) );
  AOI21_X1 U17797 ( .B1(n14763), .B2(n20809), .A(n14784), .ZN(n14773) );
  NAND2_X1 U17798 ( .A1(n14764), .A2(n16063), .ZN(n14771) );
  OR4_X1 U17799 ( .A1(n20809), .A2(n14779), .A3(n14780), .A4(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14766) );
  OAI211_X1 U17800 ( .C1(n15784), .C2(n16053), .A(n14766), .B(n14765), .ZN(
        n14768) );
  NOR2_X1 U17801 ( .A1(n15780), .A2(n16055), .ZN(n14767) );
  OAI211_X1 U17802 ( .C1(n14773), .C2(n14772), .A(n14771), .B(n14770), .ZN(
        P2_U3017) );
  INV_X1 U17803 ( .A(n14774), .ZN(n14783) );
  NAND2_X1 U17804 ( .A1(n14775), .A2(n16057), .ZN(n14777) );
  OAI211_X1 U17805 ( .C1(n16060), .C2(n14778), .A(n14777), .B(n14776), .ZN(
        n14782) );
  NOR3_X1 U17806 ( .A1(n14780), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n14779), .ZN(n14781) );
  AOI211_X1 U17807 ( .C1(n14783), .C2(n16045), .A(n14782), .B(n14781), .ZN(
        n14786) );
  NAND2_X1 U17808 ( .A1(n14784), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14785) );
  OAI211_X1 U17809 ( .C1(n14787), .C2(n16037), .A(n14786), .B(n14785), .ZN(
        P2_U3018) );
  INV_X1 U17810 ( .A(n14788), .ZN(n14796) );
  NAND2_X1 U17811 ( .A1(n14789), .A2(n16045), .ZN(n14791) );
  OAI211_X1 U17812 ( .C1(n16053), .C2(n14792), .A(n14791), .B(n14790), .ZN(
        n14795) );
  INV_X1 U17813 ( .A(n14793), .ZN(n14794) );
  AOI211_X1 U17814 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14796), .A(
        n14795), .B(n14794), .ZN(n14799) );
  NAND2_X1 U17815 ( .A1(n14797), .A2(n16033), .ZN(n14798) );
  OAI211_X1 U17816 ( .C1(n14800), .C2(n16037), .A(n14799), .B(n14798), .ZN(
        P2_U3019) );
  XNOR2_X1 U17817 ( .A(n14804), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14808) );
  AOI21_X1 U17818 ( .B1(n15797), .B2(n16057), .A(n14801), .ZN(n14803) );
  NAND2_X1 U17819 ( .A1(n15788), .A2(n16045), .ZN(n14802) );
  OAI211_X1 U17820 ( .C1(n14815), .C2(n14804), .A(n14803), .B(n14802), .ZN(
        n14807) );
  NOR2_X1 U17821 ( .A1(n14805), .A2(n16060), .ZN(n14806) );
  AOI211_X1 U17822 ( .C1(n14818), .C2(n14808), .A(n14807), .B(n14806), .ZN(
        n14809) );
  OAI21_X1 U17823 ( .B1(n14810), .B2(n16037), .A(n14809), .ZN(P2_U3020) );
  OAI22_X1 U17824 ( .A1(n19560), .A2(n11181), .B1(n16053), .B2(n14811), .ZN(
        n14812) );
  AOI21_X1 U17825 ( .B1(n14813), .B2(n16045), .A(n14812), .ZN(n14814) );
  OAI21_X1 U17826 ( .B1(n14815), .B2(n14817), .A(n14814), .ZN(n14816) );
  AOI21_X1 U17827 ( .B1(n14818), .B2(n14817), .A(n14816), .ZN(n14821) );
  NAND3_X1 U17828 ( .A1(n14819), .A2(n16033), .A3(n14638), .ZN(n14820) );
  OAI211_X1 U17829 ( .C1(n14822), .C2(n16037), .A(n14821), .B(n14820), .ZN(
        P2_U3021) );
  XOR2_X1 U17830 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n14823), .Z(
        n14824) );
  XNOR2_X1 U17831 ( .A(n14825), .B(n14824), .ZN(n15851) );
  NOR2_X1 U17832 ( .A1(n14826), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15847) );
  NOR3_X1 U17833 ( .A1(n15847), .A2(n15846), .A3(n16060), .ZN(n14835) );
  INV_X1 U17834 ( .A(n14827), .ZN(n15801) );
  INV_X1 U17835 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19558) );
  NOR2_X1 U17836 ( .A1(n19558), .A2(n16010), .ZN(n14832) );
  AOI21_X1 U17837 ( .B1(n14830), .B2(n14829), .A(n14828), .ZN(n14831) );
  AOI211_X1 U17838 ( .C1(n16057), .C2(n15801), .A(n14832), .B(n14831), .ZN(
        n14833) );
  OAI21_X1 U17839 ( .B1(n15848), .B2(n16055), .A(n14833), .ZN(n14834) );
  AOI211_X1 U17840 ( .C1(n15851), .C2(n16063), .A(n14835), .B(n14834), .ZN(
        n14836) );
  INV_X1 U17841 ( .A(n14836), .ZN(P2_U3022) );
  AOI21_X1 U17842 ( .B1(n14838), .B2(n14837), .A(n14839), .ZN(n14845) );
  NAND4_X1 U17843 ( .A1(n14859), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A4(n14839), .ZN(n14843) );
  AOI21_X1 U17844 ( .B1(n16057), .B2(n14841), .A(n14840), .ZN(n14842) );
  OAI211_X1 U17845 ( .C1(n15816), .C2(n16055), .A(n14843), .B(n14842), .ZN(
        n14844) );
  AOI211_X1 U17846 ( .C1(n14846), .C2(n16063), .A(n14845), .B(n14844), .ZN(
        n14847) );
  OAI21_X1 U17847 ( .B1(n14848), .B2(n16060), .A(n14847), .ZN(P2_U3023) );
  NAND2_X1 U17848 ( .A1(n14849), .A2(n16033), .ZN(n14861) );
  OAI21_X1 U17849 ( .B1(n14940), .B2(n14850), .A(n15977), .ZN(n14851) );
  NAND2_X1 U17850 ( .A1(n14851), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14855) );
  AOI21_X1 U17851 ( .B1(n16057), .B2(n14853), .A(n14852), .ZN(n14854) );
  OAI211_X1 U17852 ( .C1(n14856), .C2(n16055), .A(n14855), .B(n14854), .ZN(
        n14857) );
  AOI21_X1 U17853 ( .B1(n14859), .B2(n14858), .A(n14857), .ZN(n14860) );
  XNOR2_X1 U17854 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14869) );
  AOI21_X1 U17855 ( .B1(n14863), .B2(n14973), .A(n15998), .ZN(n14894) );
  INV_X1 U17856 ( .A(n14894), .ZN(n14867) );
  AOI21_X1 U17857 ( .B1(n16057), .B2(n15835), .A(n14864), .ZN(n14865) );
  OAI21_X1 U17858 ( .B1(n15822), .B2(n16055), .A(n14865), .ZN(n14866) );
  AOI21_X1 U17859 ( .B1(n14867), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14866), .ZN(n14868) );
  OAI21_X1 U17860 ( .B1(n14878), .B2(n14869), .A(n14868), .ZN(n14870) );
  AOI21_X1 U17861 ( .B1(n14871), .B2(n16033), .A(n14870), .ZN(n14872) );
  OAI21_X1 U17862 ( .B1(n16037), .B2(n14873), .A(n14872), .ZN(P2_U3026) );
  INV_X1 U17863 ( .A(n14874), .ZN(n14885) );
  INV_X1 U17864 ( .A(n14875), .ZN(n14883) );
  NAND2_X1 U17865 ( .A1(P2_REIP_REG_19__SCAN_IN), .A2(n18933), .ZN(n14876) );
  OAI221_X1 U17866 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n14878), 
        .C1(n14877), .C2(n14894), .A(n14876), .ZN(n14882) );
  OAI22_X1 U17867 ( .A1(n14880), .A2(n16055), .B1(n14879), .B2(n16053), .ZN(
        n14881) );
  AOI211_X1 U17868 ( .C1(n14883), .C2(n16033), .A(n14882), .B(n14881), .ZN(
        n14884) );
  OAI21_X1 U17869 ( .B1(n16037), .B2(n14885), .A(n14884), .ZN(P2_U3027) );
  XNOR2_X1 U17870 ( .A(n14886), .B(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15856) );
  INV_X1 U17871 ( .A(n15856), .ZN(n14906) );
  NOR2_X1 U17872 ( .A1(n14890), .A2(n14887), .ZN(n14889) );
  OAI22_X1 U17873 ( .A1(n14891), .A2(n14890), .B1(n14889), .B2(n14888), .ZN(
        n15855) );
  NAND2_X1 U17874 ( .A1(n14892), .A2(n16000), .ZN(n14895) );
  NAND2_X1 U17875 ( .A1(P2_REIP_REG_18__SCAN_IN), .A2(n18933), .ZN(n14893) );
  OAI221_X1 U17876 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n14895), 
        .C1(n14703), .C2(n14894), .A(n14893), .ZN(n14904) );
  NOR2_X1 U17877 ( .A1(n13550), .A2(n14896), .ZN(n14897) );
  OR2_X1 U17878 ( .A1(n14898), .A2(n14897), .ZN(n18671) );
  NAND2_X1 U17879 ( .A1(n14900), .A2(n14899), .ZN(n14902) );
  INV_X1 U17880 ( .A(n13613), .ZN(n14901) );
  NAND2_X1 U17881 ( .A1(n14902), .A2(n14901), .ZN(n18670) );
  OAI22_X1 U17882 ( .A1(n18671), .A2(n16055), .B1(n16053), .B2(n18670), .ZN(
        n14903) );
  AOI211_X1 U17883 ( .C1(n15855), .C2(n16063), .A(n14904), .B(n14903), .ZN(
        n14905) );
  OAI21_X1 U17884 ( .B1(n16060), .B2(n14906), .A(n14905), .ZN(P2_U3028) );
  OAI21_X1 U17885 ( .B1(n14907), .B2(n16033), .A(n9637), .ZN(n14909) );
  AOI21_X1 U17886 ( .B1(n14908), .B2(n14973), .A(n15998), .ZN(n15959) );
  OAI211_X1 U17887 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n14910), .A(
        n14909), .B(n15959), .ZN(n14929) );
  AOI21_X1 U17888 ( .B1(n14915), .B2(n14973), .A(n14929), .ZN(n14921) );
  INV_X1 U17889 ( .A(n18689), .ZN(n14917) );
  OAI21_X1 U17890 ( .B1(n18683), .B2(n16055), .A(n14911), .ZN(n14916) );
  NAND3_X1 U17891 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15979), .A3(
        n16000), .ZN(n14948) );
  INV_X1 U17892 ( .A(n14948), .ZN(n14913) );
  AND2_X1 U17893 ( .A1(n14914), .A2(n14913), .ZN(n15963) );
  NAND2_X1 U17894 ( .A1(n14918), .A2(n16063), .ZN(n14919) );
  AOI22_X1 U17895 ( .A1(n14922), .A2(n16045), .B1(P2_REIP_REG_16__SCAN_IN), 
        .B2(n18933), .ZN(n14926) );
  AOI21_X1 U17896 ( .B1(n14924), .B2(n14923), .A(n13592), .ZN(n18883) );
  NAND2_X1 U17897 ( .A1(n16057), .A2(n18883), .ZN(n14925) );
  OAI211_X1 U17898 ( .C1(n14927), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n14926), .B(n14925), .ZN(n14928) );
  AOI21_X1 U17899 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n14929), .A(
        n14928), .ZN(n14930) );
  OAI21_X1 U17900 ( .B1(n16037), .B2(n14931), .A(n14930), .ZN(P2_U3030) );
  INV_X1 U17901 ( .A(n14932), .ZN(n14934) );
  NAND2_X1 U17902 ( .A1(n14934), .A2(n14933), .ZN(n14935) );
  XNOR2_X1 U17903 ( .A(n14936), .B(n14935), .ZN(n15865) );
  INV_X1 U17904 ( .A(n15865), .ZN(n14955) );
  AND2_X1 U17905 ( .A1(n14937), .A2(n14943), .ZN(n14938) );
  NOR2_X1 U17906 ( .A1(n14939), .A2(n14938), .ZN(n15864) );
  NAND2_X1 U17907 ( .A1(n15864), .A2(n16033), .ZN(n14954) );
  NOR2_X1 U17908 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14948), .ZN(
        n15970) );
  INV_X1 U17909 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15999) );
  NOR2_X1 U17910 ( .A1(n15999), .A2(n9868), .ZN(n14941) );
  OAI21_X1 U17911 ( .B1(n14941), .B2(n14940), .A(n15977), .ZN(n15971) );
  NOR2_X1 U17912 ( .A1(n15970), .A2(n15971), .ZN(n14958) );
  OR2_X1 U17913 ( .A1(n14948), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14956) );
  NAND2_X1 U17914 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n18933), .ZN(n14942) );
  OAI221_X1 U17915 ( .B1(n14943), .B2(n14958), .C1(n14943), .C2(n14956), .A(
        n14942), .ZN(n14952) );
  AND2_X1 U17916 ( .A1(n14945), .A2(n14944), .ZN(n14947) );
  OR2_X1 U17917 ( .A1(n14947), .A2(n14946), .ZN(n18843) );
  INV_X1 U17918 ( .A(n18843), .ZN(n15863) );
  NOR4_X1 U17919 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15872), .A3(
        n14957), .A4(n14948), .ZN(n14949) );
  AOI21_X1 U17920 ( .B1(n16045), .B2(n15863), .A(n14949), .ZN(n14950) );
  OAI21_X1 U17921 ( .B1(n18721), .B2(n16053), .A(n14950), .ZN(n14951) );
  NOR2_X1 U17922 ( .A1(n14952), .A2(n14951), .ZN(n14953) );
  OAI211_X1 U17923 ( .C1(n14955), .C2(n16037), .A(n14954), .B(n14953), .ZN(
        P2_U3032) );
  NOR2_X1 U17924 ( .A1(n11098), .A2(n16010), .ZN(n14960) );
  OAI22_X1 U17925 ( .A1(n14958), .A2(n14957), .B1(n15872), .B2(n14956), .ZN(
        n14959) );
  AOI211_X1 U17926 ( .C1(n14961), .C2(n16045), .A(n14960), .B(n14959), .ZN(
        n14962) );
  OAI21_X1 U17927 ( .B1(n16053), .B2(n14963), .A(n14962), .ZN(n14964) );
  AOI21_X1 U17928 ( .B1(n14965), .B2(n16063), .A(n14964), .ZN(n14966) );
  OAI21_X1 U17929 ( .B1(n14967), .B2(n16060), .A(n14966), .ZN(P2_U3033) );
  AOI22_X1 U17930 ( .A1(n14968), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n16057), .B2(n19601), .ZN(n14977) );
  AOI22_X1 U17931 ( .A1(n16063), .A2(n14970), .B1(n16033), .B2(n14969), .ZN(
        n14976) );
  AOI21_X1 U17932 ( .B1(n16045), .B2(n14990), .A(n14971), .ZN(n14975) );
  OAI211_X1 U17933 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n14973), .B(n14972), .ZN(n14974) );
  NAND4_X1 U17934 ( .A1(n14977), .A2(n14976), .A3(n14975), .A4(n14974), .ZN(
        P2_U3045) );
  INV_X1 U17935 ( .A(n16115), .ZN(n15015) );
  INV_X1 U17936 ( .A(n14978), .ZN(n15013) );
  NAND2_X1 U17937 ( .A1(n14980), .A2(n14979), .ZN(n14985) );
  MUX2_X1 U17938 ( .A(n14985), .B(n15006), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n14981) );
  AOI21_X1 U17939 ( .B1(n18815), .B2(n15013), .A(n14981), .ZN(n16074) );
  OAI22_X1 U17940 ( .A1(n13264), .A2(n14982), .B1(n18831), .B2(n18785), .ZN(
        n14994) );
  OAI222_X1 U17941 ( .A1(n15015), .A2(n14983), .B1(n19496), .B2(n16074), .C1(
        n11065), .C2(n14994), .ZN(n14984) );
  MUX2_X1 U17942 ( .A(n14984), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n15018), .Z(P2_U3601) );
  OAI21_X1 U17943 ( .B1(n10377), .B2(n14986), .A(n14985), .ZN(n14987) );
  OAI21_X1 U17944 ( .B1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n14988), .A(
        n14987), .ZN(n14989) );
  AOI21_X1 U17945 ( .B1(n14990), .B2(n15013), .A(n14989), .ZN(n16075) );
  NAND2_X1 U17946 ( .A1(n19590), .A2(n16115), .ZN(n14997) );
  OAI21_X1 U17947 ( .B1(n13264), .B2(n14992), .A(n14991), .ZN(n14993) );
  INV_X1 U17948 ( .A(n14993), .ZN(n15016) );
  INV_X1 U17949 ( .A(n14994), .ZN(n14995) );
  NOR2_X1 U17950 ( .A1(n14995), .A2(n11065), .ZN(n14999) );
  NAND2_X1 U17951 ( .A1(n15016), .A2(n14999), .ZN(n14996) );
  OAI211_X1 U17952 ( .C1(n16075), .C2(n19496), .A(n14997), .B(n14996), .ZN(
        n14998) );
  MUX2_X1 U17953 ( .A(n14998), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15018), .Z(P2_U3600) );
  INV_X1 U17954 ( .A(n14999), .ZN(n15017) );
  NOR2_X1 U17955 ( .A1(n15001), .A2(n15000), .ZN(n15003) );
  NAND2_X1 U17956 ( .A1(n15002), .A2(n15003), .ZN(n15011) );
  INV_X1 U17957 ( .A(n15003), .ZN(n15008) );
  NOR2_X1 U17958 ( .A1(n15005), .A2(n15004), .ZN(n15007) );
  AOI22_X1 U17959 ( .A1(n15009), .A2(n15008), .B1(n15007), .B2(n15006), .ZN(
        n15010) );
  NAND2_X1 U17960 ( .A1(n15011), .A2(n15010), .ZN(n15012) );
  AOI21_X1 U17961 ( .B1(n15014), .B2(n15013), .A(n15012), .ZN(n16073) );
  OAI222_X1 U17962 ( .A1(n15017), .A2(n15016), .B1(n19496), .B2(n16073), .C1(
        n15015), .C2(n19592), .ZN(n15020) );
  MUX2_X1 U17963 ( .A(n15020), .B(n15019), .S(n15018), .Z(P2_U3599) );
  OAI21_X1 U17964 ( .B1(n19488), .B2(n19016), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n15021) );
  NAND2_X1 U17965 ( .A1(n15021), .A2(n19390), .ZN(n15029) );
  NAND2_X1 U17966 ( .A1(n19588), .A2(n19596), .ZN(n19044) );
  NOR2_X1 U17967 ( .A1(n19195), .A2(n19044), .ZN(n18982) );
  INV_X1 U17968 ( .A(n18982), .ZN(n15032) );
  AND2_X1 U17969 ( .A1(n19441), .A2(n15032), .ZN(n15027) );
  OAI21_X1 U17970 ( .B1(n10467), .B2(n18982), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15022) );
  INV_X1 U17971 ( .A(n18988), .ZN(n15040) );
  OR2_X1 U17972 ( .A1(n16114), .A2(n15023), .ZN(n15024) );
  NOR2_X2 U17973 ( .A1(n15026), .A2(n19171), .ZN(n19470) );
  INV_X1 U17974 ( .A(n19470), .ZN(n15039) );
  OAI21_X1 U17975 ( .B1(n10467), .B2(n19606), .A(n19582), .ZN(n15031) );
  INV_X1 U17976 ( .A(n15027), .ZN(n15028) );
  NOR2_X1 U17977 ( .A1(n15029), .A2(n15028), .ZN(n15030) );
  AOI211_X2 U17978 ( .C1(n15032), .C2(n15031), .A(n19171), .B(n15030), .ZN(
        n18991) );
  INV_X1 U17979 ( .A(n18991), .ZN(n15041) );
  INV_X1 U17980 ( .A(n19488), .ZN(n15036) );
  NAND2_X1 U17981 ( .A1(n19390), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19598) );
  AOI22_X1 U17982 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n18979), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n18978), .ZN(n19474) );
  AOI22_X1 U17983 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n18979), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n18978), .ZN(n19420) );
  NOR2_X2 U17984 ( .A1(n9782), .A2(n18980), .ZN(n19469) );
  AOI22_X1 U17985 ( .A1(n19471), .A2(n19016), .B1(n18982), .B2(n19469), .ZN(
        n15035) );
  OAI21_X1 U17986 ( .B1(n15036), .B2(n19474), .A(n15035), .ZN(n15037) );
  AOI21_X1 U17987 ( .B1(n15041), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A(
        n15037), .ZN(n15038) );
  OAI21_X1 U17988 ( .B1(n15040), .B2(n15039), .A(n15038), .ZN(P2_U3052) );
  NAND2_X1 U17989 ( .A1(n15041), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n15046) );
  NOR2_X2 U17990 ( .A1(n10723), .A2(n18980), .ZN(n20826) );
  AOI22_X1 U17991 ( .A1(n20829), .A2(n19016), .B1(n18982), .B2(n20826), .ZN(
        n15045) );
  NOR2_X2 U17992 ( .A1(n15042), .A2(n19171), .ZN(n20827) );
  NAND2_X1 U17993 ( .A1(n18988), .A2(n20827), .ZN(n15044) );
  AOI22_X1 U17994 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18978), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n18979), .ZN(n20835) );
  INV_X1 U17995 ( .A(n20835), .ZN(n19421) );
  NAND2_X1 U17996 ( .A1(n19488), .A2(n19421), .ZN(n15043) );
  NAND4_X1 U17997 ( .A1(n15046), .A2(n15045), .A3(n15044), .A4(n15043), .ZN(
        P2_U3053) );
  INV_X1 U17998 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16396) );
  INV_X1 U17999 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16417) );
  INV_X1 U18000 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16460) );
  NAND2_X1 U18001 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16748), .ZN(n15123) );
  INV_X1 U18002 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16376) );
  NOR2_X1 U18003 ( .A1(n17108), .A2(n16991), .ZN(n16988) );
  NOR2_X1 U18004 ( .A1(n16992), .A2(n16748), .ZN(n16743) );
  AOI21_X1 U18005 ( .B1(n16988), .B2(n15047), .A(n16743), .ZN(n16736) );
  AOI22_X1 U18006 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15260), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15052) );
  AOI22_X1 U18007 ( .A1(n9613), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16946), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15051) );
  AOI22_X1 U18008 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9615), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15050) );
  AOI22_X1 U18009 ( .A1(n15224), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15049) );
  NAND4_X1 U18010 ( .A1(n15052), .A2(n15051), .A3(n15050), .A4(n15049), .ZN(
        n15059) );
  AOI22_X1 U18011 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15057) );
  AOI22_X1 U18012 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15056) );
  AOI22_X1 U18013 ( .A1(n13753), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15055) );
  AOI22_X1 U18014 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15054) );
  NAND4_X1 U18015 ( .A1(n15057), .A2(n15056), .A3(n15055), .A4(n15054), .ZN(
        n15058) );
  NOR2_X1 U18016 ( .A1(n15059), .A2(n15058), .ZN(n16732) );
  AOI22_X1 U18017 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15063) );
  AOI22_X1 U18018 ( .A1(n15048), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16946), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15062) );
  AOI22_X1 U18019 ( .A1(n15224), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15061) );
  AOI22_X1 U18020 ( .A1(n9628), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15060) );
  NAND4_X1 U18021 ( .A1(n15063), .A2(n15062), .A3(n15061), .A4(n15060), .ZN(
        n15069) );
  AOI22_X1 U18022 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15067) );
  AOI22_X1 U18023 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15260), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15066) );
  AOI22_X1 U18024 ( .A1(n9613), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15065) );
  AOI22_X1 U18025 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15064) );
  NAND4_X1 U18026 ( .A1(n15067), .A2(n15066), .A3(n15065), .A4(n15064), .ZN(
        n15068) );
  NOR2_X1 U18027 ( .A1(n15069), .A2(n15068), .ZN(n16746) );
  AOI22_X1 U18028 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n16909), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15073) );
  AOI22_X1 U18029 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15072) );
  AOI22_X1 U18030 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n16928), .ZN(n15071) );
  AOI22_X1 U18031 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n9615), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15070) );
  NAND4_X1 U18032 ( .A1(n15073), .A2(n15072), .A3(n15071), .A4(n15070), .ZN(
        n15079) );
  AOI22_X1 U18033 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15077) );
  AOI22_X1 U18034 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16895), .B1(
        n9613), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15076) );
  AOI22_X1 U18035 ( .A1(n15224), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n16927), .ZN(n15075) );
  AOI22_X1 U18036 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n16937), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n15053), .ZN(n15074) );
  NAND4_X1 U18037 ( .A1(n15077), .A2(n15076), .A3(n15075), .A4(n15074), .ZN(
        n15078) );
  NOR2_X1 U18038 ( .A1(n15079), .A2(n15078), .ZN(n16754) );
  AOI22_X1 U18039 ( .A1(n15224), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15089) );
  AOI22_X1 U18040 ( .A1(n9613), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15088) );
  INV_X1 U18041 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15262) );
  AOI22_X1 U18042 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15080) );
  OAI21_X1 U18043 ( .B1(n15112), .B2(n15262), .A(n15080), .ZN(n15086) );
  AOI22_X1 U18044 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15084) );
  AOI22_X1 U18045 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16946), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15083) );
  AOI22_X1 U18046 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15082) );
  AOI22_X1 U18047 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15081) );
  NAND4_X1 U18048 ( .A1(n15084), .A2(n15083), .A3(n15082), .A4(n15081), .ZN(
        n15085) );
  AOI211_X1 U18049 ( .C1(n16936), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n15086), .B(n15085), .ZN(n15087) );
  NAND3_X1 U18050 ( .A1(n15089), .A2(n15088), .A3(n15087), .ZN(n16758) );
  AOI22_X1 U18051 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9615), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15099) );
  AOI22_X1 U18052 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15098) );
  INV_X1 U18053 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n20778) );
  AOI22_X1 U18054 ( .A1(n15224), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15090) );
  OAI21_X1 U18055 ( .B1(n16646), .B2(n20778), .A(n15090), .ZN(n15096) );
  AOI22_X1 U18056 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15094) );
  AOI22_X1 U18057 ( .A1(n13753), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15093) );
  AOI22_X1 U18058 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15092) );
  AOI22_X1 U18059 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15091) );
  NAND4_X1 U18060 ( .A1(n15094), .A2(n15093), .A3(n15092), .A4(n15091), .ZN(
        n15095) );
  AOI211_X1 U18061 ( .C1(n16929), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n15096), .B(n15095), .ZN(n15097) );
  NAND3_X1 U18062 ( .A1(n15099), .A2(n15098), .A3(n15097), .ZN(n16759) );
  NAND2_X1 U18063 ( .A1(n16758), .A2(n16759), .ZN(n16757) );
  NOR2_X1 U18064 ( .A1(n16754), .A2(n16757), .ZN(n16751) );
  AOI22_X1 U18065 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15110) );
  INV_X1 U18066 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16911) );
  AOI22_X1 U18067 ( .A1(n13753), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15101) );
  AOI22_X1 U18068 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15100) );
  OAI211_X1 U18069 ( .C1(n15236), .C2(n16911), .A(n15101), .B(n15100), .ZN(
        n15108) );
  AOI22_X1 U18070 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15260), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15106) );
  AOI22_X1 U18071 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15105) );
  AOI22_X1 U18072 ( .A1(n16896), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15104) );
  AOI22_X1 U18073 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15103) );
  NAND4_X1 U18074 ( .A1(n15106), .A2(n15105), .A3(n15104), .A4(n15103), .ZN(
        n15107) );
  AOI211_X1 U18075 ( .C1(n16954), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n15108), .B(n15107), .ZN(n15109) );
  NAND2_X1 U18076 ( .A1(n15110), .A2(n15109), .ZN(n16750) );
  NAND2_X1 U18077 ( .A1(n16751), .A2(n16750), .ZN(n16749) );
  NOR2_X1 U18078 ( .A1(n16746), .A2(n16749), .ZN(n16741) );
  AOI22_X1 U18079 ( .A1(n16909), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15121) );
  AOI22_X1 U18080 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15120) );
  AOI22_X1 U18081 ( .A1(n9628), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15111) );
  OAI21_X1 U18082 ( .B1(n15112), .B2(n16976), .A(n15111), .ZN(n15118) );
  AOI22_X1 U18083 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15116) );
  AOI22_X1 U18084 ( .A1(n15048), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15115) );
  AOI22_X1 U18085 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15114) );
  AOI22_X1 U18086 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15113) );
  NAND4_X1 U18087 ( .A1(n15116), .A2(n15115), .A3(n15114), .A4(n15113), .ZN(
        n15117) );
  AOI211_X1 U18088 ( .C1(n9615), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n15118), .B(n15117), .ZN(n15119) );
  NAND3_X1 U18089 ( .A1(n15121), .A2(n15120), .A3(n15119), .ZN(n16740) );
  NAND2_X1 U18090 ( .A1(n16741), .A2(n16740), .ZN(n16739) );
  XOR2_X1 U18091 ( .A(n16732), .B(n16739), .Z(n17010) );
  NAND2_X1 U18092 ( .A1(n16992), .A2(n17010), .ZN(n15122) );
  OAI221_X1 U18093 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n15123), .C1(n16376), 
        .C2(n16736), .A(n15122), .ZN(P3_U2675) );
  AOI22_X1 U18094 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15127) );
  AOI22_X1 U18095 ( .A1(n9628), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15126) );
  AOI22_X1 U18096 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13732), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15125) );
  AOI22_X1 U18097 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15124) );
  NAND4_X1 U18098 ( .A1(n15127), .A2(n15126), .A3(n15125), .A4(n15124), .ZN(
        n15133) );
  AOI22_X1 U18099 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15131) );
  AOI22_X1 U18100 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13772), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15130) );
  AOI22_X1 U18101 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15129) );
  AOI22_X1 U18102 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15128) );
  NAND4_X1 U18103 ( .A1(n15131), .A2(n15130), .A3(n15129), .A4(n15128), .ZN(
        n15132) );
  NOR2_X1 U18104 ( .A1(n15133), .A2(n15132), .ZN(n17087) );
  INV_X1 U18105 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n16545) );
  INV_X1 U18106 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n16576) );
  INV_X1 U18107 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n20811) );
  NOR2_X1 U18108 ( .A1(n17108), .A2(n16968), .ZN(n16969) );
  NAND3_X1 U18109 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(n16969), .ZN(n16962) );
  NOR4_X1 U18110 ( .A1(n16576), .A2(n15134), .A3(n20811), .A4(n16962), .ZN(
        n15135) );
  NAND2_X1 U18111 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n15135), .ZN(n16891) );
  NOR2_X1 U18112 ( .A1(n16545), .A2(n16891), .ZN(n16862) );
  OAI221_X1 U18113 ( .B1(n16862), .B2(P3_EBX_REG_13__SCAN_IN), .C1(n9736), 
        .C2(n15136), .A(n16986), .ZN(n15137) );
  OAI21_X1 U18114 ( .B1(n17087), .B2(n16986), .A(n15137), .ZN(P3_U2690) );
  NOR2_X1 U18115 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18569), .ZN(
        n18228) );
  INV_X1 U18116 ( .A(n18228), .ZN(n15139) );
  NAND3_X1 U18117 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18568)
         );
  NAND2_X1 U18118 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18432) );
  INV_X1 U18119 ( .A(n18432), .ZN(n18436) );
  AOI21_X1 U18120 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18436), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15177) );
  INV_X1 U18121 ( .A(n15177), .ZN(n15138) );
  NOR2_X1 U18122 ( .A1(n16934), .A2(n15138), .ZN(n17962) );
  NAND2_X1 U18123 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n17960) );
  INV_X1 U18124 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18577) );
  NAND2_X1 U18125 ( .A1(n18577), .A2(n18468), .ZN(n18477) );
  NOR2_X1 U18126 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18569), .ZN(
        n18592) );
  AOI21_X1 U18127 ( .B1(n17960), .B2(n18477), .A(n18592), .ZN(n17970) );
  NOR2_X1 U18128 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17970), .ZN(n18253) );
  INV_X1 U18129 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16309) );
  OR2_X1 U18130 ( .A1(n16309), .A2(n18568), .ZN(n15175) );
  OAI211_X1 U18131 ( .C1(n18568), .C2(n17962), .A(n18227), .B(n15175), .ZN(
        n17968) );
  NAND2_X1 U18132 ( .A1(n15139), .A2(n17968), .ZN(n15142) );
  INV_X1 U18133 ( .A(n15142), .ZN(n15141) );
  INV_X1 U18134 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18620) );
  NOR3_X1 U18135 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n18620), .ZN(n18115) );
  INV_X1 U18136 ( .A(n18115), .ZN(n18250) );
  NAND2_X1 U18137 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17523) );
  INV_X1 U18138 ( .A(n17523), .ZN(n17585) );
  NAND2_X1 U18139 ( .A1(n18569), .A2(n17960), .ZN(n18614) );
  OAI22_X1 U18140 ( .A1(n17585), .A2(n18614), .B1(n18412), .B2(n18569), .ZN(
        n15144) );
  NAND3_X1 U18141 ( .A1(n18413), .A2(n17968), .A3(n15144), .ZN(n15140) );
  OAI221_X1 U18142 ( .B1(n18413), .B2(n15141), .C1(n18413), .C2(n18250), .A(
        n15140), .ZN(P3_U2864) );
  NAND2_X1 U18143 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18113) );
  NOR2_X1 U18144 ( .A1(n17585), .A2(n18614), .ZN(n15143) );
  AOI221_X1 U18145 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18113), .C1(n15143), 
        .C2(n18113), .A(n15142), .ZN(n17967) );
  OAI221_X1 U18146 ( .B1(n18115), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18115), .C2(n15144), .A(n17968), .ZN(n17965) );
  AOI22_X1 U18147 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17967), .B1(
        n17965), .B2(n18420), .ZN(P3_U2865) );
  NAND4_X1 U18148 ( .A1(n17985), .A2(n17989), .A3(n15161), .A4(n15151), .ZN(
        n15329) );
  NOR2_X1 U18149 ( .A1(n15309), .A2(n17993), .ZN(n15458) );
  NOR2_X1 U18150 ( .A1(n18621), .A2(n17971), .ZN(n15145) );
  NOR2_X1 U18151 ( .A1(n15145), .A2(n15308), .ZN(n15150) );
  AND2_X1 U18152 ( .A1(n15146), .A2(n15150), .ZN(n15147) );
  OAI211_X1 U18153 ( .C1(n17989), .C2(n15458), .A(n15326), .B(n15147), .ZN(
        n15310) );
  NAND3_X1 U18154 ( .A1(n17981), .A2(n17997), .A3(n17989), .ZN(n15164) );
  NAND2_X1 U18155 ( .A1(n17981), .A2(n15151), .ZN(n15315) );
  NAND2_X1 U18156 ( .A1(n15164), .A2(n15315), .ZN(n15155) );
  INV_X1 U18157 ( .A(n17985), .ZN(n15149) );
  INV_X1 U18158 ( .A(n15458), .ZN(n18408) );
  OAI22_X1 U18159 ( .A1(n15161), .A2(n15149), .B1(n15148), .B2(n18408), .ZN(
        n15154) );
  NOR2_X1 U18160 ( .A1(n18005), .A2(n15151), .ZN(n15152) );
  OAI22_X1 U18161 ( .A1(n17989), .A2(n15152), .B1(n15151), .B2(n15150), .ZN(
        n15153) );
  INV_X1 U18162 ( .A(n15166), .ZN(n15157) );
  NAND2_X1 U18163 ( .A1(n18621), .A2(n17971), .ZN(n15156) );
  AOI21_X1 U18164 ( .B1(n17108), .B2(n18408), .A(n15156), .ZN(n15163) );
  AOI211_X1 U18165 ( .C1(n15159), .C2(n15310), .A(n15157), .B(n15163), .ZN(
        n15324) );
  XNOR2_X1 U18166 ( .A(n18621), .B(n16642), .ZN(n18624) );
  INV_X1 U18167 ( .A(n15164), .ZN(n15158) );
  NAND4_X1 U18168 ( .A1(n15326), .A2(n17993), .A3(n15158), .A4(n17971), .ZN(
        n17187) );
  NAND2_X1 U18169 ( .A1(n17187), .A2(n15159), .ZN(n16307) );
  INV_X1 U18170 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18490) );
  INV_X1 U18171 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18482) );
  INV_X2 U18172 ( .A(n18608), .ZN(n18630) );
  OAI211_X1 U18173 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18490), .B(n18553), .ZN(n18619) );
  NOR2_X1 U18174 ( .A1(n15325), .A2(n18619), .ZN(n17147) );
  NAND3_X1 U18175 ( .A1(n18621), .A2(n15161), .A3(n15160), .ZN(n15162) );
  AOI21_X1 U18176 ( .B1(n15165), .B2(n15164), .A(n15163), .ZN(n15167) );
  OAI21_X1 U18177 ( .B1(n17985), .B2(n15167), .A(n15166), .ZN(n15327) );
  NOR2_X1 U18178 ( .A1(n15329), .A2(n15327), .ZN(n15333) );
  NAND2_X1 U18179 ( .A1(n15330), .A2(n15333), .ZN(n15176) );
  XOR2_X1 U18180 ( .A(n15170), .B(n15169), .Z(n15172) );
  NAND2_X1 U18181 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18622) );
  OAI211_X1 U18182 ( .C1(n17147), .C2(n16323), .A(n18424), .B(n18622), .ZN(
        n15174) );
  NAND2_X1 U18183 ( .A1(n16126), .A2(n15331), .ZN(n15173) );
  NAND3_X1 U18184 ( .A1(n15324), .A2(n15174), .A3(n15173), .ZN(n18450) );
  INV_X1 U18185 ( .A(n18450), .ZN(n18442) );
  NAND2_X1 U18186 ( .A1(n18566), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n17969) );
  OAI211_X1 U18187 ( .C1(n18459), .C2(n18442), .A(n17969), .B(n15175), .ZN(
        n18596) );
  NOR2_X1 U18188 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18594) );
  NOR2_X1 U18189 ( .A1(n15177), .A2(n15176), .ZN(n18453) );
  NAND3_X1 U18190 ( .A1(n18596), .A2(n18594), .A3(n18453), .ZN(n15178) );
  OAI21_X1 U18191 ( .B1(n18596), .B2(n18451), .A(n15178), .ZN(P3_U3284) );
  AOI22_X1 U18192 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15260), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15182) );
  AOI22_X1 U18193 ( .A1(n9628), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9613), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15181) );
  AOI22_X1 U18194 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15180) );
  AOI22_X1 U18195 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15179) );
  NAND4_X1 U18196 ( .A1(n15182), .A2(n15181), .A3(n15180), .A4(n15179), .ZN(
        n15188) );
  AOI22_X1 U18197 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15186) );
  AOI22_X1 U18198 ( .A1(n16896), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15185) );
  AOI22_X1 U18199 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15184) );
  AOI22_X1 U18200 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15183) );
  NAND4_X1 U18201 ( .A1(n15186), .A2(n15185), .A3(n15184), .A4(n15183), .ZN(
        n15187) );
  AOI22_X1 U18202 ( .A1(n13753), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15200) );
  AOI22_X1 U18203 ( .A1(n16896), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15260), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15199) );
  INV_X1 U18204 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n20670) );
  AOI22_X1 U18205 ( .A1(n9628), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9613), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15189) );
  OAI21_X1 U18206 ( .B1(n15190), .B2(n20670), .A(n15189), .ZN(n15197) );
  AOI22_X1 U18207 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15201), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15195) );
  AOI22_X1 U18208 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15194) );
  AOI22_X1 U18209 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15193) );
  AOI22_X1 U18210 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15192) );
  NAND4_X1 U18211 ( .A1(n15195), .A2(n15194), .A3(n15193), .A4(n15192), .ZN(
        n15196) );
  AOI211_X1 U18212 ( .C1(n16929), .C2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n15197), .B(n15196), .ZN(n15198) );
  NAND3_X1 U18213 ( .A1(n15200), .A2(n15199), .A3(n15198), .ZN(n15338) );
  AOI22_X1 U18214 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15201), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15212) );
  INV_X1 U18215 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15204) );
  AOI22_X1 U18216 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15260), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15203) );
  AOI22_X1 U18217 ( .A1(n16909), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15202) );
  OAI211_X1 U18218 ( .C1(n15236), .C2(n15204), .A(n15203), .B(n15202), .ZN(
        n15210) );
  AOI22_X1 U18219 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15223), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15208) );
  AOI22_X1 U18220 ( .A1(n13753), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15207) );
  AOI22_X1 U18221 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n9614), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15206) );
  AOI22_X1 U18222 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15205) );
  NAND4_X1 U18223 ( .A1(n15208), .A2(n15207), .A3(n15206), .A4(n15205), .ZN(
        n15209) );
  AOI211_X1 U18224 ( .C1(n16954), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n15210), .B(n15209), .ZN(n15211) );
  NAND2_X1 U18225 ( .A1(n15212), .A2(n15211), .ZN(n15337) );
  AOI22_X1 U18226 ( .A1(n15223), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15216) );
  AOI22_X1 U18227 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15215) );
  AOI22_X1 U18228 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15260), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15214) );
  AOI22_X1 U18229 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15213) );
  NAND4_X1 U18230 ( .A1(n15216), .A2(n15215), .A3(n15214), .A4(n15213), .ZN(
        n15222) );
  AOI22_X1 U18231 ( .A1(n15191), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15201), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15220) );
  AOI22_X1 U18232 ( .A1(n15048), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15264), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15219) );
  AOI22_X1 U18233 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15218) );
  AOI22_X1 U18234 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9619), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15217) );
  NAND4_X1 U18235 ( .A1(n15220), .A2(n15219), .A3(n15218), .A4(n15217), .ZN(
        n15221) );
  AOI22_X1 U18236 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n13770), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n15264), .ZN(n15229) );
  AOI22_X1 U18237 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n15224), .B1(
        n15223), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15228) );
  AOI22_X1 U18238 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n13700), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n15225), .ZN(n15227) );
  AOI22_X1 U18239 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n15263), .B1(
        n9676), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15226) );
  AOI22_X1 U18240 ( .A1(n15191), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15201), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15230) );
  INV_X1 U18241 ( .A(n15230), .ZN(n15231) );
  INV_X1 U18242 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15235) );
  AOI22_X1 U18243 ( .A1(n15048), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9613), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15234) );
  AOI22_X1 U18244 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16927), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n16946), .ZN(n15233) );
  OAI211_X1 U18245 ( .C1(n15236), .C2(n15235), .A(n15234), .B(n15233), .ZN(
        n15237) );
  AOI22_X1 U18246 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15242) );
  AOI22_X1 U18247 ( .A1(n16896), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15241) );
  AOI22_X1 U18248 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15240) );
  AOI22_X1 U18249 ( .A1(n13753), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15260), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15239) );
  NAND4_X1 U18250 ( .A1(n15242), .A2(n15241), .A3(n15240), .A4(n15239), .ZN(
        n15248) );
  AOI22_X1 U18251 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15246) );
  AOI22_X1 U18252 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15245) );
  AOI22_X1 U18253 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15244) );
  AOI22_X1 U18254 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15243) );
  NAND4_X1 U18255 ( .A1(n15246), .A2(n15245), .A3(n15244), .A4(n15243), .ZN(
        n15247) );
  AOI22_X1 U18256 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15201), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15258) );
  AOI22_X1 U18257 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15260), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15250) );
  AOI22_X1 U18258 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15249) );
  OAI211_X1 U18259 ( .C1(n9668), .C2(n20778), .A(n15250), .B(n15249), .ZN(
        n15256) );
  AOI22_X1 U18260 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15254) );
  AOI22_X1 U18261 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15253) );
  AOI22_X1 U18262 ( .A1(n9614), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15252) );
  AOI22_X1 U18263 ( .A1(n16946), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15251) );
  NAND4_X1 U18264 ( .A1(n15254), .A2(n15253), .A3(n15252), .A4(n15251), .ZN(
        n15255) );
  AOI211_X1 U18265 ( .C1(n15053), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n15256), .B(n15255), .ZN(n15257) );
  INV_X1 U18266 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17905) );
  AOI22_X1 U18267 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15260), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15274) );
  AOI22_X1 U18268 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16946), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15273) );
  AOI22_X1 U18269 ( .A1(n16896), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9613), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15261) );
  OAI21_X1 U18270 ( .B1(n16646), .B2(n15262), .A(n15261), .ZN(n15271) );
  AOI22_X1 U18271 ( .A1(n15191), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15201), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15269) );
  AOI22_X1 U18272 ( .A1(n15223), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15263), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15268) );
  AOI22_X1 U18273 ( .A1(n15048), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15264), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15267) );
  AOI22_X1 U18274 ( .A1(n16937), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9619), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15266) );
  NAND4_X1 U18275 ( .A1(n15269), .A2(n15268), .A3(n15267), .A4(n15266), .ZN(
        n15270) );
  AOI211_X1 U18276 ( .C1(n16936), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n15271), .B(n15270), .ZN(n15272) );
  NOR2_X1 U18277 ( .A1(n17615), .A2(n17622), .ZN(n17614) );
  INV_X1 U18278 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18579) );
  NOR2_X1 U18279 ( .A1(n17139), .A2(n18579), .ZN(n15275) );
  INV_X1 U18280 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n15347) );
  XOR2_X1 U18281 ( .A(n17138), .B(n17139), .Z(n15276) );
  NOR2_X1 U18282 ( .A1(n17606), .A2(n17605), .ZN(n15278) );
  NOR2_X1 U18283 ( .A1(n15347), .A2(n15276), .ZN(n15277) );
  INV_X1 U18284 ( .A(n15337), .ZN(n17129) );
  XOR2_X1 U18285 ( .A(n17129), .B(n15279), .Z(n17595) );
  NOR2_X1 U18286 ( .A1(n9675), .A2(n17905), .ZN(n15280) );
  INV_X1 U18287 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17577) );
  NOR2_X1 U18288 ( .A1(n15282), .A2(n17577), .ZN(n15283) );
  XOR2_X1 U18289 ( .A(n17125), .B(n15281), .Z(n17582) );
  XNOR2_X1 U18290 ( .A(n17577), .B(n15282), .ZN(n17581) );
  NOR2_X1 U18291 ( .A1(n17582), .A2(n17581), .ZN(n17580) );
  NOR2_X2 U18292 ( .A1(n15283), .A2(n17580), .ZN(n17566) );
  XOR2_X1 U18293 ( .A(n15338), .B(n15284), .Z(n17567) );
  NAND2_X1 U18294 ( .A1(n17566), .A2(n17567), .ZN(n17565) );
  XNOR2_X1 U18295 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n15286), .ZN(
        n17556) );
  INV_X1 U18296 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17885) );
  NOR2_X2 U18297 ( .A1(n17545), .A2(n17885), .ZN(n17544) );
  INV_X1 U18299 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17862) );
  NAND2_X1 U18300 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17831) );
  INV_X1 U18301 ( .A(n17831), .ZN(n17801) );
  NAND2_X1 U18302 ( .A1(n17801), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17815) );
  INV_X1 U18303 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17814) );
  NOR2_X1 U18304 ( .A1(n17815), .A2(n17814), .ZN(n17780) );
  INV_X1 U18305 ( .A(n17780), .ZN(n17782) );
  INV_X1 U18306 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17786) );
  NOR2_X1 U18307 ( .A1(n17782), .A2(n17786), .ZN(n17784) );
  AND2_X1 U18308 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17784), .ZN(
        n17759) );
  NAND2_X1 U18309 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17759), .ZN(
        n17745) );
  NOR2_X2 U18310 ( .A1(n17427), .A2(n17745), .ZN(n15295) );
  INV_X1 U18311 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17761) );
  NOR4_X1 U18312 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15290) );
  INV_X1 U18313 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17789) );
  INV_X1 U18314 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17767) );
  NAND4_X1 U18315 ( .A1(n15290), .A2(n17814), .A3(n17789), .A4(n17767), .ZN(
        n15291) );
  INV_X1 U18316 ( .A(n15294), .ZN(n15296) );
  NOR2_X2 U18317 ( .A1(n15296), .A2(n15295), .ZN(n17411) );
  NAND2_X1 U18318 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17397) );
  INV_X1 U18319 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17400) );
  INV_X1 U18320 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17361) );
  NAND2_X1 U18321 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17700) );
  NOR3_X1 U18322 ( .A1(n17400), .A2(n17361), .A3(n17700), .ZN(n17337) );
  NAND2_X1 U18323 ( .A1(n17337), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17679) );
  NOR2_X2 U18324 ( .A1(n17395), .A2(n17679), .ZN(n17319) );
  NOR2_X1 U18325 ( .A1(n17397), .A2(n17679), .ZN(n17300) );
  NAND2_X1 U18326 ( .A1(n17300), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17668) );
  NAND2_X1 U18327 ( .A1(n17400), .A2(n17516), .ZN(n17394) );
  NOR2_X1 U18328 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17394), .ZN(
        n15298) );
  INV_X1 U18329 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15297) );
  NAND2_X1 U18330 ( .A1(n15298), .A2(n15297), .ZN(n17357) );
  NOR2_X1 U18331 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17357), .ZN(
        n17336) );
  INV_X1 U18332 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17339) );
  INV_X1 U18333 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17685) );
  NAND3_X1 U18334 ( .A1(n17336), .A2(n17339), .A3(n17685), .ZN(n15299) );
  INV_X1 U18335 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17654) );
  NAND2_X1 U18336 ( .A1(n17313), .A2(n17654), .ZN(n17312) );
  NAND2_X1 U18337 ( .A1(n17304), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15303) );
  INV_X1 U18338 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17658) );
  NAND2_X1 U18339 ( .A1(n17516), .A2(n17658), .ZN(n15302) );
  NAND2_X1 U18340 ( .A1(n17516), .A2(n17312), .ZN(n17303) );
  INV_X1 U18341 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17648) );
  OR2_X1 U18342 ( .A1(n15303), .A2(n17648), .ZN(n15304) );
  NAND2_X1 U18343 ( .A1(n15305), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16190) );
  NOR2_X2 U18344 ( .A1(n15305), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17270) );
  NOR2_X1 U18345 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17534), .ZN(
        n15306) );
  NAND2_X1 U18346 ( .A1(n17270), .A2(n15306), .ZN(n15441) );
  NAND2_X1 U18347 ( .A1(n15440), .A2(n15441), .ZN(n15307) );
  XNOR2_X1 U18348 ( .A(n15307), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16176) );
  NOR2_X1 U18349 ( .A1(n18621), .A2(n15308), .ZN(n15317) );
  NAND2_X1 U18350 ( .A1(n15317), .A2(n15309), .ZN(n15311) );
  INV_X1 U18351 ( .A(n16196), .ZN(n18425) );
  INV_X1 U18352 ( .A(n15311), .ZN(n15322) );
  INV_X1 U18353 ( .A(n15312), .ZN(n15313) );
  INV_X1 U18354 ( .A(n18424), .ZN(n15318) );
  AOI21_X1 U18355 ( .B1(n15314), .B2(n15313), .A(n15318), .ZN(n18426) );
  INV_X1 U18356 ( .A(n16126), .ZN(n18429) );
  AOI21_X1 U18357 ( .B1(n17989), .B2(n15315), .A(n18429), .ZN(n15321) );
  OAI21_X1 U18358 ( .B1(n17981), .B2(n17188), .A(n18619), .ZN(n15316) );
  OAI21_X1 U18359 ( .B1(n15317), .B2(n15316), .A(n18622), .ZN(n16306) );
  NOR3_X1 U18360 ( .A1(n15319), .A2(n15318), .A3(n16306), .ZN(n15320) );
  AOI211_X1 U18361 ( .C1(n15322), .C2(n18426), .A(n15321), .B(n15320), .ZN(
        n15323) );
  AOI21_X2 U18362 ( .B1(n15324), .B2(n15323), .A(n18459), .ZN(n17952) );
  NOR3_X4 U18363 ( .A1(n17114), .A2(n18425), .A3(n17938), .ZN(n17870) );
  INV_X1 U18364 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16172) );
  INV_X1 U18365 ( .A(n15325), .ZN(n16324) );
  NOR3_X1 U18366 ( .A1(n16324), .A2(n15326), .A3(n18621), .ZN(n15328) );
  NOR2_X1 U18367 ( .A1(n15328), .A2(n15327), .ZN(n18401) );
  NAND2_X1 U18368 ( .A1(n15330), .A2(n15329), .ZN(n18433) );
  NAND2_X1 U18369 ( .A1(n17952), .A2(n17899), .ZN(n17943) );
  NAND2_X1 U18370 ( .A1(n18468), .A2(n18594), .ZN(n16303) );
  INV_X1 U18371 ( .A(n16303), .ZN(n18634) );
  NOR2_X2 U18372 ( .A1(n15333), .A2(n15332), .ZN(n18400) );
  INV_X1 U18373 ( .A(n18400), .ZN(n18411) );
  NOR2_X1 U18374 ( .A1(n18438), .A2(n18411), .ZN(n17841) );
  NOR2_X2 U18375 ( .A1(n17951), .A2(n17952), .ZN(n17936) );
  INV_X1 U18376 ( .A(n17300), .ZN(n17674) );
  NAND2_X1 U18377 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17301) );
  NOR2_X1 U18378 ( .A1(n17658), .A2(n17301), .ZN(n17644) );
  NAND2_X1 U18379 ( .A1(n17644), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15367) );
  NOR2_X1 U18380 ( .A1(n17674), .A2(n15367), .ZN(n16149) );
  NOR3_X1 U18381 ( .A1(n9946), .A2(n17905), .A3(n17577), .ZN(n17865) );
  INV_X1 U18382 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17876) );
  NOR2_X1 U18383 ( .A1(n17885), .A2(n17876), .ZN(n17755) );
  NAND3_X1 U18384 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17865), .A3(
        n17755), .ZN(n17742) );
  INV_X1 U18385 ( .A(n17742), .ZN(n15334) );
  INV_X1 U18386 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18595) );
  OAI21_X1 U18387 ( .B1(n18595), .B2(n18579), .A(n15347), .ZN(n17923) );
  NAND2_X1 U18388 ( .A1(n15334), .A2(n17923), .ZN(n17781) );
  NOR2_X1 U18389 ( .A1(n17745), .A2(n17781), .ZN(n17678) );
  AOI21_X1 U18390 ( .B1(n16149), .B2(n17678), .A(n18406), .ZN(n17631) );
  NAND2_X1 U18391 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17901) );
  NOR2_X1 U18392 ( .A1(n17742), .A2(n17901), .ZN(n17838) );
  NAND2_X1 U18393 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17838), .ZN(
        n17847) );
  NOR2_X1 U18394 ( .A1(n17745), .A2(n17847), .ZN(n15369) );
  INV_X1 U18395 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17279) );
  INV_X1 U18396 ( .A(n16149), .ZN(n17630) );
  NOR2_X1 U18397 ( .A1(n17279), .A2(n17630), .ZN(n16189) );
  INV_X1 U18398 ( .A(n17848), .ZN(n18409) );
  AOI21_X1 U18399 ( .B1(n15369), .B2(n16189), .A(n18409), .ZN(n15336) );
  INV_X1 U18400 ( .A(n17745), .ZN(n17412) );
  NAND2_X1 U18401 ( .A1(n17412), .A2(n17838), .ZN(n15370) );
  INV_X1 U18402 ( .A(n15370), .ZN(n17697) );
  AOI21_X1 U18403 ( .B1(n16149), .B2(n17697), .A(n18400), .ZN(n15335) );
  NOR4_X1 U18404 ( .A1(n17936), .A2(n17631), .A3(n15336), .A4(n15335), .ZN(
        n15443) );
  OAI21_X1 U18405 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17841), .A(
        n15443), .ZN(n16198) );
  NAND2_X1 U18406 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16170) );
  NOR2_X1 U18407 ( .A1(n16170), .A2(n16172), .ZN(n16141) );
  NAND2_X1 U18408 ( .A1(n9640), .A2(n17759), .ZN(n17446) );
  NAND2_X1 U18409 ( .A1(n17694), .A2(n16149), .ZN(n17632) );
  INV_X1 U18410 ( .A(n17632), .ZN(n15373) );
  NAND2_X1 U18411 ( .A1(n16141), .A2(n15373), .ZN(n16161) );
  INV_X1 U18412 ( .A(n16161), .ZN(n16155) );
  NAND2_X1 U18413 ( .A1(n16196), .A2(n17952), .ZN(n17949) );
  NOR2_X1 U18414 ( .A1(n16195), .A2(n17949), .ZN(n17794) );
  INV_X1 U18415 ( .A(n17794), .ZN(n17874) );
  NAND2_X1 U18416 ( .A1(n17623), .A2(n17139), .ZN(n15342) );
  NAND2_X1 U18417 ( .A1(n17138), .A2(n15342), .ZN(n15341) );
  NAND2_X1 U18418 ( .A1(n15341), .A2(n15337), .ZN(n15352) );
  NOR2_X1 U18419 ( .A1(n17125), .A2(n15352), .ZN(n15339) );
  NAND2_X1 U18420 ( .A1(n15339), .A2(n15338), .ZN(n15355) );
  NOR2_X1 U18421 ( .A1(n17118), .A2(n15355), .ZN(n15359) );
  NAND2_X1 U18422 ( .A1(n15359), .A2(n16195), .ZN(n15360) );
  XNOR2_X1 U18423 ( .A(n15339), .B(n17122), .ZN(n15340) );
  AND2_X1 U18424 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15340), .ZN(
        n15354) );
  XNOR2_X1 U18425 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n15340), .ZN(
        n17564) );
  XNOR2_X1 U18426 ( .A(n17129), .B(n15341), .ZN(n15349) );
  AND2_X1 U18427 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15349), .ZN(
        n15350) );
  XOR2_X1 U18428 ( .A(n17138), .B(n15342), .Z(n15346) );
  NOR2_X1 U18429 ( .A1(n15346), .A2(n15347), .ZN(n15348) );
  NOR2_X1 U18430 ( .A1(n15259), .A2(n18595), .ZN(n15345) );
  INV_X1 U18431 ( .A(n17623), .ZN(n15344) );
  NAND3_X1 U18432 ( .A1(n15344), .A2(n15259), .A3(n18595), .ZN(n15343) );
  OAI221_X1 U18433 ( .B1(n15345), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n15344), .C2(n15259), .A(n15343), .ZN(n17604) );
  XNOR2_X1 U18434 ( .A(n15347), .B(n15346), .ZN(n17603) );
  NOR2_X1 U18435 ( .A1(n17604), .A2(n17603), .ZN(n17602) );
  NOR2_X1 U18436 ( .A1(n15348), .A2(n17602), .ZN(n17593) );
  XNOR2_X1 U18437 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n15349), .ZN(
        n17592) );
  NOR2_X1 U18438 ( .A1(n17593), .A2(n17592), .ZN(n17591) );
  NOR2_X1 U18439 ( .A1(n15350), .A2(n17591), .ZN(n17575) );
  XOR2_X1 U18440 ( .A(n15352), .B(n15351), .Z(n17576) );
  NOR2_X1 U18441 ( .A1(n17575), .A2(n17576), .ZN(n15353) );
  NAND2_X1 U18442 ( .A1(n17575), .A2(n17576), .ZN(n17574) );
  OAI21_X1 U18443 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15353), .A(
        n17574), .ZN(n17563) );
  XNOR2_X1 U18444 ( .A(n15355), .B(n17118), .ZN(n15357) );
  NOR2_X1 U18445 ( .A1(n15356), .A2(n15357), .ZN(n15358) );
  XNOR2_X1 U18446 ( .A(n15357), .B(n15356), .ZN(n17551) );
  NOR2_X1 U18447 ( .A1(n15358), .A2(n17550), .ZN(n15361) );
  XNOR2_X1 U18448 ( .A(n15359), .B(n16195), .ZN(n15362) );
  NAND2_X1 U18449 ( .A1(n15361), .A2(n15362), .ZN(n17541) );
  NAND2_X1 U18450 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17541), .ZN(
        n15364) );
  NOR2_X1 U18451 ( .A1(n15360), .A2(n15364), .ZN(n15366) );
  INV_X1 U18452 ( .A(n15360), .ZN(n15365) );
  OR2_X1 U18453 ( .A1(n15362), .A2(n15361), .ZN(n17542) );
  OAI21_X1 U18454 ( .B1(n15365), .B2(n15364), .A(n17542), .ZN(n15363) );
  AOI21_X1 U18455 ( .B1(n15365), .B2(n15364), .A(n15363), .ZN(n17531) );
  NOR2_X1 U18456 ( .A1(n17531), .A2(n17862), .ZN(n17530) );
  OR2_X2 U18457 ( .A1(n15366), .A2(n17530), .ZN(n17823) );
  NAND3_X1 U18458 ( .A1(n17807), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17441) );
  NOR2_X2 U18459 ( .A1(n17441), .A2(n17767), .ZN(n17693) );
  NOR2_X2 U18460 ( .A1(n17672), .A2(n15367), .ZN(n16124) );
  AND2_X1 U18461 ( .A1(n16124), .A2(n16141), .ZN(n16171) );
  NAND2_X1 U18462 ( .A1(n18428), .A2(n17952), .ZN(n17914) );
  OAI22_X1 U18463 ( .A1(n16155), .A2(n17874), .B1(n16171), .B2(n17914), .ZN(
        n15444) );
  AOI21_X1 U18464 ( .B1(n17861), .B2(n16198), .A(n15444), .ZN(n15368) );
  OAI21_X1 U18465 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17943), .A(
        n15368), .ZN(n15375) );
  INV_X1 U18466 ( .A(n16124), .ZN(n17633) );
  INV_X1 U18467 ( .A(n17678), .ZN(n17695) );
  NOR2_X1 U18468 ( .A1(n18406), .A2(n17695), .ZN(n16188) );
  INV_X1 U18469 ( .A(n15369), .ZN(n17757) );
  OAI22_X1 U18470 ( .A1(n18400), .A2(n15370), .B1(n18409), .B2(n17757), .ZN(
        n15371) );
  OAI211_X1 U18471 ( .C1(n16188), .C2(n15371), .A(n17952), .B(n16149), .ZN(
        n16177) );
  OAI21_X1 U18472 ( .B1(n17914), .B2(n17633), .A(n16177), .ZN(n15372) );
  AOI21_X1 U18473 ( .B1(n15373), .B2(n17794), .A(n15372), .ZN(n15447) );
  OAI21_X1 U18474 ( .B1(n16170), .B2(n15447), .A(n16172), .ZN(n15374) );
  OAI21_X1 U18475 ( .B1(n16172), .B2(n15375), .A(n15374), .ZN(n15376) );
  NAND2_X1 U18476 ( .A1(n17951), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16169) );
  OAI211_X1 U18477 ( .C1(n16176), .C2(n17845), .A(n15376), .B(n16169), .ZN(
        P3_U2833) );
  INV_X1 U18478 ( .A(n15829), .ZN(n15377) );
  OAI22_X1 U18479 ( .A1(n15819), .A2(n18789), .B1(n18812), .B2(n15377), .ZN(
        n15378) );
  INV_X1 U18480 ( .A(n15378), .ZN(n15387) );
  AOI211_X1 U18481 ( .C1(n15381), .C2(n15380), .A(n15379), .B(n18779), .ZN(
        n15385) );
  AOI22_X1 U18482 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n9607), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18669), .ZN(n15382) );
  OAI21_X1 U18483 ( .B1(n15383), .B2(n18795), .A(n15382), .ZN(n15384) );
  AOI211_X1 U18484 ( .C1(P2_EBX_REG_22__SCAN_IN), .C2(n18819), .A(n15385), .B(
        n15384), .ZN(n15386) );
  NAND2_X1 U18485 ( .A1(n15387), .A2(n15386), .ZN(P2_U2833) );
  NAND2_X1 U18486 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n15448), .ZN(n15415) );
  INV_X1 U18487 ( .A(n15415), .ZN(n20625) );
  INV_X1 U18488 ( .A(n15388), .ZN(n15395) );
  NOR3_X1 U18489 ( .A1(n15391), .A2(n15390), .A3(n15389), .ZN(n15392) );
  AOI21_X1 U18490 ( .B1(n15396), .B2(n11604), .A(n15392), .ZN(n15393) );
  OAI21_X1 U18491 ( .B1(n20292), .B2(n15394), .A(n15393), .ZN(n20596) );
  NAND2_X1 U18492 ( .A1(n15395), .A2(n20596), .ZN(n15399) );
  INV_X1 U18493 ( .A(n15399), .ZN(n15401) );
  AOI21_X1 U18494 ( .B1(n15396), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n20639), .ZN(n15397) );
  OAI211_X1 U18495 ( .C1(n15399), .C2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15398), .B(n15397), .ZN(n15400) );
  OAI21_X1 U18496 ( .B1(n15401), .B2(n20436), .A(n15400), .ZN(n15403) );
  AOI222_X1 U18497 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n15403), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15402), .C1(n15403), 
        .C2(n15402), .ZN(n15405) );
  AOI222_X1 U18498 ( .A1(n15405), .A2(n20217), .B1(n15405), .B2(n15404), .C1(
        n20217), .C2(n15404), .ZN(n15414) );
  AOI21_X1 U18499 ( .B1(n19638), .B2(n15407), .A(n15406), .ZN(n15409) );
  NOR4_X1 U18500 ( .A1(n15411), .A2(n15410), .A3(n15409), .A4(n15408), .ZN(
        n15412) );
  OAI211_X1 U18501 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n15414), .A(
        n15413), .B(n15412), .ZN(n15421) );
  OR2_X1 U18502 ( .A1(n15422), .A2(n20626), .ZN(n20501) );
  OAI211_X1 U18503 ( .C1(n15417), .C2(n15416), .A(n20501), .B(n15415), .ZN(
        n15768) );
  AOI221_X1 U18504 ( .B1(n15763), .B2(n15418), .C1(n15421), .C2(n15418), .A(
        n15768), .ZN(n15423) );
  NOR2_X1 U18505 ( .A1(n15423), .A2(n15763), .ZN(n15771) );
  INV_X1 U18506 ( .A(n15771), .ZN(n15419) );
  AOI211_X1 U18507 ( .C1(n15422), .C2(n15421), .A(n15420), .B(n15419), .ZN(
        n15428) );
  OAI21_X1 U18508 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20507), .A(n20437), 
        .ZN(n15766) );
  AOI21_X1 U18509 ( .B1(n15425), .B2(n15424), .A(n15423), .ZN(n15426) );
  NOR2_X1 U18510 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15426), .ZN(n15427) );
  AOI221_X1 U18511 ( .B1(n20625), .B2(n15428), .C1(n15766), .C2(n15428), .A(
        n15427), .ZN(P1_U3161) );
  OAI21_X1 U18512 ( .B1(n15529), .B2(n15638), .A(n15429), .ZN(n15545) );
  XNOR2_X1 U18513 ( .A(n15529), .B(n15430), .ZN(n15544) );
  AOI21_X1 U18514 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15434), .A(
        n15544), .ZN(n15433) );
  OAI21_X1 U18515 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15431), .A(
        n15430), .ZN(n15432) );
  OAI211_X1 U18516 ( .C1(n15545), .C2(n15434), .A(n15433), .B(n15432), .ZN(
        n15435) );
  XNOR2_X1 U18517 ( .A(n15435), .B(n15623), .ZN(n15535) );
  INV_X1 U18518 ( .A(n15484), .ZN(n15438) );
  NAND3_X1 U18519 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n15436), .ZN(n15621) );
  NAND2_X1 U18520 ( .A1(n19819), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15541) );
  OAI221_X1 U18521 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n15621), 
        .C1(n15623), .C2(n15630), .A(n15541), .ZN(n15437) );
  AOI21_X1 U18522 ( .B1(n15438), .B2(n19826), .A(n15437), .ZN(n15439) );
  OAI21_X1 U18523 ( .B1(n15685), .B2(n15535), .A(n15439), .ZN(P1_U3010) );
  INV_X1 U18524 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16142) );
  NAND2_X1 U18525 ( .A1(n16141), .A2(n16142), .ZN(n16160) );
  NOR2_X2 U18526 ( .A1(n15441), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16133) );
  NOR2_X1 U18527 ( .A1(n16134), .A2(n16133), .ZN(n15442) );
  XNOR2_X1 U18528 ( .A(n15442), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16156) );
  AOI22_X1 U18529 ( .A1(n17951), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n17870), 
        .B2(n16156), .ZN(n15446) );
  OAI22_X1 U18530 ( .A1(n17951), .A2(n15443), .B1(n16141), .B2(n17943), .ZN(
        n16182) );
  OAI21_X1 U18531 ( .B1(n16182), .B2(n15444), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15445) );
  OAI211_X1 U18532 ( .C1(n15447), .C2(n16160), .A(n15446), .B(n15445), .ZN(
        P3_U2832) );
  INV_X1 U18533 ( .A(HOLD), .ZN(n20782) );
  INV_X1 U18534 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20509) );
  NAND2_X1 U18535 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20509), .ZN(n20506) );
  INV_X1 U18536 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20508) );
  NOR2_X1 U18537 ( .A1(n20504), .A2(n20508), .ZN(n20512) );
  INV_X1 U18538 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20510) );
  NOR2_X1 U18539 ( .A1(n20510), .A2(n15448), .ZN(n15449) );
  AOI221_X1 U18540 ( .B1(n20782), .B2(n20512), .C1(n20509), .C2(n20512), .A(
        n15449), .ZN(n15451) );
  OAI211_X1 U18541 ( .C1(n20782), .C2(n20506), .A(n15451), .B(n15450), .ZN(
        P1_U3195) );
  INV_X1 U18542 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20635) );
  NOR2_X1 U18543 ( .A1(n20635), .A2(n19747), .ZN(P1_U2905) );
  NAND2_X1 U18544 ( .A1(n19504), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19495) );
  INV_X1 U18545 ( .A(n19495), .ZN(n15453) );
  NAND2_X1 U18546 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATEBS16_REG_SCAN_IN), .ZN(n19579) );
  OAI21_X1 U18547 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n19579), .A(n19606), 
        .ZN(n15452) );
  AOI21_X1 U18548 ( .B1(n15453), .B2(P2_STATE2_REG_1__SCAN_IN), .A(n15452), 
        .ZN(n15454) );
  NOR2_X1 U18549 ( .A1(n16121), .A2(n15454), .ZN(P2_U3178) );
  INV_X1 U18550 ( .A(n16111), .ZN(n19616) );
  AOI221_X1 U18551 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16121), .C1(n19616), .C2(
        n16121), .A(n19444), .ZN(n19611) );
  AND2_X1 U18552 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n19611), .ZN(
        P2_U3047) );
  NOR3_X1 U18553 ( .A1(n15455), .A2(n17971), .A3(n17188), .ZN(n15456) );
  INV_X1 U18554 ( .A(n18459), .ZN(n18615) );
  INV_X1 U18555 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17219) );
  NOR2_X2 U18556 ( .A1(n15459), .A2(n17219), .ZN(n17144) );
  OR2_X1 U18557 ( .A1(n17108), .A2(n15459), .ZN(n17040) );
  NOR2_X1 U18558 ( .A1(n15459), .A2(n18005), .ZN(n17134) );
  INV_X2 U18559 ( .A(n17134), .ZN(n17143) );
  AOI22_X1 U18560 ( .A1(n17141), .A2(BUF2_REG_0__SCAN_IN), .B1(n17140), .B2(
        n17623), .ZN(n15460) );
  OAI221_X1 U18561 ( .B1(n17144), .B2(n17219), .C1(n17144), .C2(n17040), .A(
        n15460), .ZN(P3_U2735) );
  NOR2_X1 U18562 ( .A1(n15469), .A2(n15506), .ZN(n15480) );
  AOI21_X1 U18563 ( .B1(n15461), .B2(n15480), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n15467) );
  INV_X1 U18564 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15462) );
  OAI22_X1 U18565 ( .A1(n15462), .A2(n15525), .B1(n19731), .B2(n15534), .ZN(
        n15463) );
  AOI21_X1 U18566 ( .B1(n19695), .B2(P1_EBX_REG_23__SCAN_IN), .A(n15463), .ZN(
        n15465) );
  AOI22_X1 U18567 ( .A1(n15531), .A2(n19663), .B1(n19700), .B2(n15614), .ZN(
        n15464) );
  OAI211_X1 U18568 ( .C1(n15467), .C2(n15466), .A(n15465), .B(n15464), .ZN(
        P1_U2817) );
  AOI21_X1 U18569 ( .B1(n15469), .B2(n15468), .A(n15500), .ZN(n15490) );
  OAI22_X1 U18570 ( .A1(n15471), .A2(n15525), .B1(n19715), .B2(n15470), .ZN(
        n15475) );
  OAI22_X1 U18571 ( .A1(n15473), .A2(n15521), .B1(n15472), .B2(n19718), .ZN(
        n15474) );
  OAI211_X1 U18572 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(P1_REIP_REG_21__SCAN_IN), .A(n15480), .B(n15477), .ZN(n15478) );
  OAI211_X1 U18573 ( .C1(n15490), .C2(n20555), .A(n15479), .B(n15478), .ZN(
        P1_U2818) );
  INV_X1 U18574 ( .A(n15480), .ZN(n15488) );
  INV_X1 U18575 ( .A(n15539), .ZN(n15486) );
  INV_X1 U18576 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15543) );
  OAI22_X1 U18577 ( .A1(n15543), .A2(n15525), .B1(n19731), .B2(n15481), .ZN(
        n15482) );
  AOI21_X1 U18578 ( .B1(n19695), .B2(P1_EBX_REG_21__SCAN_IN), .A(n15482), .ZN(
        n15483) );
  OAI21_X1 U18579 ( .B1(n15484), .B2(n19718), .A(n15483), .ZN(n15485) );
  AOI21_X1 U18580 ( .B1(n15486), .B2(n19663), .A(n15485), .ZN(n15487) );
  OAI221_X1 U18581 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n15488), .C1(n20553), 
        .C2(n15490), .A(n15487), .ZN(P1_U2819) );
  AOI22_X1 U18582 ( .A1(n19695), .A2(P1_EBX_REG_20__SCAN_IN), .B1(n19703), 
        .B2(n15489), .ZN(n15498) );
  INV_X1 U18583 ( .A(n15490), .ZN(n15496) );
  INV_X1 U18584 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20550) );
  OAI21_X1 U18585 ( .B1(n15491), .B2(n15506), .A(n20550), .ZN(n15495) );
  OAI22_X1 U18586 ( .A1(n15493), .A2(n15521), .B1(n19718), .B2(n15492), .ZN(
        n15494) );
  AOI21_X1 U18587 ( .B1(n15496), .B2(n15495), .A(n15494), .ZN(n15497) );
  OAI211_X1 U18588 ( .C1(n15499), .C2(n15525), .A(n15498), .B(n15497), .ZN(
        P1_U2820) );
  NAND2_X1 U18589 ( .A1(n15500), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15505) );
  AOI21_X1 U18590 ( .B1(n19721), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n19662), .ZN(n15501) );
  OAI21_X1 U18591 ( .B1(n15502), .B2(n19731), .A(n15501), .ZN(n15503) );
  AOI21_X1 U18592 ( .B1(n19695), .B2(P1_EBX_REG_18__SCAN_IN), .A(n15503), .ZN(
        n15504) );
  OAI211_X1 U18593 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n15506), .A(n15505), 
        .B(n15504), .ZN(n15507) );
  AOI21_X1 U18594 ( .B1(n15508), .B2(n19663), .A(n15507), .ZN(n15509) );
  OAI21_X1 U18595 ( .B1(n19718), .B2(n15641), .A(n15509), .ZN(P1_U2822) );
  INV_X1 U18596 ( .A(n15678), .ZN(n15510) );
  NAND2_X1 U18597 ( .A1(n19700), .A2(n15510), .ZN(n15513) );
  NAND2_X1 U18598 ( .A1(n19721), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15511) );
  AND2_X1 U18599 ( .A1(n15511), .A2(n19683), .ZN(n15512) );
  OAI211_X1 U18600 ( .C1(n19715), .C2(n14145), .A(n15513), .B(n15512), .ZN(
        n15514) );
  INV_X1 U18601 ( .A(n15514), .ZN(n15520) );
  INV_X1 U18602 ( .A(n15515), .ZN(n15516) );
  NAND2_X1 U18603 ( .A1(n15516), .A2(n19653), .ZN(n15522) );
  OAI21_X1 U18604 ( .B1(n20536), .B2(n15522), .A(n20538), .ZN(n15517) );
  AOI22_X1 U18605 ( .A1(n15573), .A2(n19703), .B1(n15518), .B2(n15517), .ZN(
        n15519) );
  OAI211_X1 U18606 ( .C1(n15521), .C2(n15571), .A(n15520), .B(n15519), .ZN(
        P1_U2828) );
  AOI22_X1 U18607 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15523), .B1(n15522), 
        .B2(n20536), .ZN(n15527) );
  INV_X1 U18608 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n20650) );
  AOI22_X1 U18609 ( .A1(n19695), .A2(P1_EBX_REG_11__SCAN_IN), .B1(n19700), 
        .B2(n15687), .ZN(n15524) );
  OAI211_X1 U18610 ( .C1(n15525), .C2(n20650), .A(n15524), .B(n19683), .ZN(
        n15526) );
  AOI211_X1 U18611 ( .C1(n19663), .C2(n15579), .A(n15527), .B(n15526), .ZN(
        n15528) );
  OAI21_X1 U18612 ( .B1(n15582), .B2(n19731), .A(n15528), .ZN(P1_U2829) );
  AOI22_X1 U18613 ( .A1(n19813), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n19819), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n15533) );
  XNOR2_X1 U18614 ( .A(n15529), .B(n20803), .ZN(n15530) );
  XNOR2_X1 U18615 ( .A(n14223), .B(n15530), .ZN(n15615) );
  AOI22_X1 U18616 ( .A1(n15531), .A2(n14290), .B1(n19817), .B2(n15615), .ZN(
        n15532) );
  OAI211_X1 U18617 ( .C1(n15597), .C2(n15534), .A(n15533), .B(n15532), .ZN(
        P1_U2976) );
  INV_X1 U18618 ( .A(n15535), .ZN(n15536) );
  AOI22_X1 U18619 ( .A1(n15600), .A2(n15537), .B1(n19817), .B2(n15536), .ZN(
        n15538) );
  OAI21_X1 U18620 ( .B1(n15539), .B2(n19841), .A(n15538), .ZN(n15540) );
  INV_X1 U18621 ( .A(n15540), .ZN(n15542) );
  OAI211_X1 U18622 ( .C1(n15543), .C2(n15603), .A(n15542), .B(n15541), .ZN(
        P1_U2978) );
  AOI22_X1 U18623 ( .A1(n19813), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n19819), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15548) );
  XNOR2_X1 U18624 ( .A(n15545), .B(n15544), .ZN(n15634) );
  AOI22_X1 U18625 ( .A1(n15634), .A2(n19817), .B1(n15546), .B2(n14290), .ZN(
        n15547) );
  OAI211_X1 U18626 ( .C1(n15597), .C2(n15549), .A(n15548), .B(n15547), .ZN(
        P1_U2980) );
  INV_X1 U18627 ( .A(n15550), .ZN(n15552) );
  MUX2_X1 U18628 ( .A(n15553), .B(n15552), .S(n15551), .Z(n15554) );
  XNOR2_X1 U18629 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n15554), .ZN(
        n15655) );
  AOI22_X1 U18630 ( .A1(n19813), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n19819), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15558) );
  AOI22_X1 U18631 ( .A1(n15556), .A2(n14290), .B1(n15600), .B2(n15555), .ZN(
        n15557) );
  OAI211_X1 U18632 ( .C1(n19637), .C2(n15655), .A(n15558), .B(n15557), .ZN(
        P1_U2982) );
  NOR2_X1 U18633 ( .A1(n15560), .A2(n15559), .ZN(n15561) );
  XNOR2_X1 U18634 ( .A(n15562), .B(n15561), .ZN(n15662) );
  AOI22_X1 U18635 ( .A1(n19813), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n19819), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15566) );
  AOI22_X1 U18636 ( .A1(n15564), .A2(n14290), .B1(n15600), .B2(n15563), .ZN(
        n15565) );
  OAI211_X1 U18637 ( .C1(n15662), .C2(n19637), .A(n15566), .B(n15565), .ZN(
        P1_U2984) );
  INV_X1 U18638 ( .A(n15567), .ZN(n15568) );
  AOI21_X1 U18639 ( .B1(n15570), .B2(n15569), .A(n15568), .ZN(n15686) );
  AOI22_X1 U18640 ( .A1(n19813), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n19819), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15575) );
  INV_X1 U18641 ( .A(n15571), .ZN(n15572) );
  AOI22_X1 U18642 ( .A1(n15600), .A2(n15573), .B1(n14290), .B2(n15572), .ZN(
        n15574) );
  OAI211_X1 U18643 ( .C1(n15686), .C2(n19637), .A(n15575), .B(n15574), .ZN(
        P1_U2987) );
  AOI22_X1 U18644 ( .A1(n19813), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n19819), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15581) );
  NAND2_X1 U18645 ( .A1(n15529), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15577) );
  OAI21_X1 U18646 ( .B1(n14297), .B2(n15577), .A(n15576), .ZN(n15578) );
  XNOR2_X1 U18647 ( .A(n15578), .B(n15694), .ZN(n15691) );
  AOI22_X1 U18648 ( .A1(n19817), .A2(n15691), .B1(n14290), .B2(n15579), .ZN(
        n15580) );
  OAI211_X1 U18649 ( .C1(n15597), .C2(n15582), .A(n15581), .B(n15580), .ZN(
        P1_U2988) );
  AOI22_X1 U18650 ( .A1(n19813), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n19819), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15589) );
  NAND2_X1 U18651 ( .A1(n15584), .A2(n15583), .ZN(n15585) );
  NAND2_X1 U18652 ( .A1(n15586), .A2(n15585), .ZN(n15735) );
  AOI22_X1 U18653 ( .A1(n15735), .A2(n19817), .B1(n14290), .B2(n15587), .ZN(
        n15588) );
  OAI211_X1 U18654 ( .C1(n15597), .C2(n15590), .A(n15589), .B(n15588), .ZN(
        P1_U2992) );
  AOI22_X1 U18655 ( .A1(n19813), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n19819), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15596) );
  NAND2_X1 U18656 ( .A1(n15592), .A2(n15591), .ZN(n15593) );
  XNOR2_X1 U18657 ( .A(n15594), .B(n15593), .ZN(n15741) );
  AOI22_X1 U18658 ( .A1(n15741), .A2(n19817), .B1(n14290), .B2(n19664), .ZN(
        n15595) );
  OAI211_X1 U18659 ( .C1(n15597), .C2(n19665), .A(n15596), .B(n15595), .ZN(
        P1_U2993) );
  INV_X1 U18660 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n15604) );
  XOR2_X1 U18661 ( .A(n15599), .B(n15598), .Z(n15756) );
  INV_X1 U18662 ( .A(n19682), .ZN(n15601) );
  AOI222_X1 U18663 ( .A1(n15756), .A2(n19817), .B1(n14290), .B2(n19740), .C1(
        n15601), .C2(n15600), .ZN(n15602) );
  NAND2_X1 U18664 ( .A1(n19819), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n15751) );
  OAI211_X1 U18665 ( .C1(n15604), .C2(n15603), .A(n15602), .B(n15751), .ZN(
        P1_U2994) );
  NOR2_X1 U18666 ( .A1(n15731), .A2(n20561), .ZN(n15608) );
  NOR4_X1 U18667 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n20803), .A3(
        n15606), .A4(n15605), .ZN(n15607) );
  AOI211_X1 U18668 ( .C1(n15609), .C2(n19824), .A(n15608), .B(n15607), .ZN(
        n15613) );
  AOI22_X1 U18669 ( .A1(n19826), .A2(n15611), .B1(n15610), .B2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15612) );
  NAND2_X1 U18670 ( .A1(n15613), .A2(n15612), .ZN(P1_U3006) );
  AOI22_X1 U18671 ( .A1(n15615), .A2(n19824), .B1(n19826), .B2(n15614), .ZN(
        n15620) );
  NOR2_X1 U18672 ( .A1(n15731), .A2(n20557), .ZN(n15616) );
  AOI221_X1 U18673 ( .B1(n15618), .B2(n20803), .C1(n15617), .C2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n15616), .ZN(n15619) );
  NAND2_X1 U18674 ( .A1(n15620), .A2(n15619), .ZN(P1_U3008) );
  AOI211_X1 U18675 ( .C1(n15623), .C2(n14277), .A(n15622), .B(n15621), .ZN(
        n15624) );
  AOI21_X1 U18676 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n19819), .A(n15624), 
        .ZN(n15629) );
  INV_X1 U18677 ( .A(n15625), .ZN(n15627) );
  AOI22_X1 U18678 ( .A1(n15627), .A2(n19824), .B1(n19826), .B2(n15626), .ZN(
        n15628) );
  OAI211_X1 U18679 ( .C1(n15630), .C2(n14277), .A(n15629), .B(n15628), .ZN(
        P1_U3009) );
  INV_X1 U18680 ( .A(n15631), .ZN(n15632) );
  AOI22_X1 U18681 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15632), .B1(
        n19819), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15636) );
  AOI22_X1 U18682 ( .A1(n15634), .A2(n19824), .B1(n19826), .B2(n15633), .ZN(
        n15635) );
  OAI211_X1 U18683 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15637), .A(
        n15636), .B(n15635), .ZN(P1_U3012) );
  NAND2_X1 U18684 ( .A1(n15640), .A2(n15638), .ZN(n15646) );
  OAI21_X1 U18685 ( .B1(n15702), .B2(n15640), .A(n15639), .ZN(n15651) );
  OAI22_X1 U18686 ( .A1(n15642), .A2(n15685), .B1(n15733), .B2(n15641), .ZN(
        n15643) );
  AOI21_X1 U18687 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15651), .A(
        n15643), .ZN(n15645) );
  NAND2_X1 U18688 ( .A1(n19819), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15644) );
  OAI211_X1 U18689 ( .C1(n15648), .C2(n15646), .A(n15645), .B(n15644), .ZN(
        P1_U3013) );
  OAI21_X1 U18690 ( .B1(n15649), .B2(n15648), .A(n15647), .ZN(n15652) );
  AOI22_X1 U18691 ( .A1(n15652), .A2(n15651), .B1(n19826), .B2(n15650), .ZN(
        n15654) );
  NAND2_X1 U18692 ( .A1(n19819), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15653) );
  OAI211_X1 U18693 ( .C1(n15655), .C2(n15685), .A(n15654), .B(n15653), .ZN(
        P1_U3014) );
  INV_X1 U18694 ( .A(n15656), .ZN(n15657) );
  AOI22_X1 U18695 ( .A1(n15657), .A2(n19826), .B1(n19819), .B2(
        P1_REIP_REG_15__SCAN_IN), .ZN(n15661) );
  AOI21_X1 U18696 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15659), .A(
        n15658), .ZN(n15660) );
  OAI211_X1 U18697 ( .C1(n15662), .C2(n15685), .A(n15661), .B(n15660), .ZN(
        P1_U3016) );
  AOI22_X1 U18698 ( .A1(n15664), .A2(n19824), .B1(n19826), .B2(n15663), .ZN(
        n15671) );
  NAND2_X1 U18699 ( .A1(n19819), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15670) );
  OAI21_X1 U18700 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15666), .A(
        n15665), .ZN(n15669) );
  NAND3_X1 U18701 ( .A1(n19833), .A2(n15667), .A3(n12575), .ZN(n15668) );
  NAND4_X1 U18702 ( .A1(n15671), .A2(n15670), .A3(n15669), .A4(n15668), .ZN(
        P1_U3018) );
  INV_X1 U18703 ( .A(n15672), .ZN(n15677) );
  OAI22_X1 U18704 ( .A1(n15674), .A2(n15673), .B1(n15682), .B2(n19829), .ZN(
        n15675) );
  NOR2_X1 U18705 ( .A1(n15676), .A2(n15675), .ZN(n15695) );
  OAI21_X1 U18706 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15677), .A(
        n15695), .ZN(n15680) );
  OAI22_X1 U18707 ( .A1(n15733), .A2(n15678), .B1(n20538), .B2(n15731), .ZN(
        n15679) );
  AOI21_X1 U18708 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15680), .A(
        n15679), .ZN(n15684) );
  NAND3_X1 U18709 ( .A1(n15682), .A2(n15681), .A3(n15696), .ZN(n15683) );
  OAI211_X1 U18710 ( .C1(n15686), .C2(n15685), .A(n15684), .B(n15683), .ZN(
        P1_U3019) );
  AOI22_X1 U18711 ( .A1(n19826), .A2(n15687), .B1(n19819), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n15693) );
  NOR3_X1 U18712 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15689), .A3(
        n15688), .ZN(n15690) );
  AOI21_X1 U18713 ( .B1(n15691), .B2(n19824), .A(n15690), .ZN(n15692) );
  OAI211_X1 U18714 ( .C1(n15695), .C2(n15694), .A(n15693), .B(n15692), .ZN(
        P1_U3020) );
  NAND2_X1 U18715 ( .A1(n15701), .A2(n15696), .ZN(n15716) );
  OAI21_X1 U18716 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15697), .ZN(n15706) );
  AOI21_X1 U18717 ( .B1(n19826), .B2(n15699), .A(n15698), .ZN(n15705) );
  OAI21_X1 U18718 ( .B1(n15702), .B2(n15701), .A(n15700), .ZN(n15712) );
  AOI22_X1 U18719 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15712), .B1(
        n19824), .B2(n15703), .ZN(n15704) );
  OAI211_X1 U18720 ( .C1(n15716), .C2(n15706), .A(n15705), .B(n15704), .ZN(
        P1_U3021) );
  NAND2_X1 U18721 ( .A1(n15708), .A2(n15707), .ZN(n15709) );
  AND2_X1 U18722 ( .A1(n15710), .A2(n15709), .ZN(n19733) );
  AOI21_X1 U18723 ( .B1(n19826), .B2(n19733), .A(n15711), .ZN(n15715) );
  AOI22_X1 U18724 ( .A1(n15713), .A2(n19824), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15712), .ZN(n15714) );
  OAI211_X1 U18725 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n15716), .A(
        n15715), .B(n15714), .ZN(P1_U3022) );
  INV_X1 U18726 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15723) );
  OR2_X1 U18727 ( .A1(n15719), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15754) );
  NOR2_X1 U18728 ( .A1(n15740), .A2(n19829), .ZN(n15718) );
  AOI211_X1 U18729 ( .C1(n15720), .C2(n15719), .A(n15718), .B(n15717), .ZN(
        n15759) );
  OAI21_X1 U18730 ( .B1(n15721), .B2(n15754), .A(n15759), .ZN(n15742) );
  AOI21_X1 U18731 ( .B1(n15723), .B2(n15722), .A(n15742), .ZN(n15737) );
  INV_X1 U18732 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15730) );
  INV_X1 U18733 ( .A(n15724), .ZN(n15728) );
  INV_X1 U18734 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15738) );
  NAND3_X1 U18735 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15740), .A3(
        n15746), .ZN(n15739) );
  AOI221_X1 U18736 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n15730), .C2(n15738), .A(
        n15739), .ZN(n15727) );
  OAI22_X1 U18737 ( .A1(n15733), .A2(n15725), .B1(n20530), .B2(n15731), .ZN(
        n15726) );
  AOI211_X1 U18738 ( .C1(n15728), .C2(n19824), .A(n15727), .B(n15726), .ZN(
        n15729) );
  OAI21_X1 U18739 ( .B1(n15737), .B2(n15730), .A(n15729), .ZN(P1_U3023) );
  OAI22_X1 U18740 ( .A1(n15733), .A2(n15732), .B1(n20529), .B2(n15731), .ZN(
        n15734) );
  AOI21_X1 U18741 ( .B1(n15735), .B2(n19824), .A(n15734), .ZN(n15736) );
  OAI221_X1 U18742 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15739), .C1(
        n15738), .C2(n15737), .A(n15736), .ZN(P1_U3024) );
  NAND2_X1 U18743 ( .A1(n15740), .A2(n15746), .ZN(n15745) );
  AOI22_X1 U18744 ( .A1(n19826), .A2(n19667), .B1(n19819), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n15744) );
  AOI22_X1 U18745 ( .A1(n15742), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n19824), .B2(n15741), .ZN(n15743) );
  OAI211_X1 U18746 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n15745), .A(
        n15744), .B(n15743), .ZN(P1_U3025) );
  INV_X1 U18747 ( .A(n15746), .ZN(n15753) );
  NAND2_X1 U18748 ( .A1(n15748), .A2(n15747), .ZN(n15749) );
  AND2_X1 U18749 ( .A1(n15750), .A2(n15749), .ZN(n19737) );
  NAND2_X1 U18750 ( .A1(n19826), .A2(n19737), .ZN(n15752) );
  OAI211_X1 U18751 ( .C1(n15754), .C2(n15753), .A(n15752), .B(n15751), .ZN(
        n15755) );
  AOI21_X1 U18752 ( .B1(n15756), .B2(n19824), .A(n15755), .ZN(n15757) );
  OAI21_X1 U18753 ( .B1(n15759), .B2(n15758), .A(n15757), .ZN(P1_U3026) );
  INV_X1 U18754 ( .A(n20605), .ZN(n20607) );
  NAND3_X1 U18755 ( .A1(n15761), .A2(n15760), .A3(n20595), .ZN(n15762) );
  OAI21_X1 U18756 ( .B1(n20607), .B2(n13217), .A(n15762), .ZN(P1_U3468) );
  NAND3_X1 U18757 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20437), .A3(n20625), 
        .ZN(n15764) );
  NAND2_X1 U18758 ( .A1(n15765), .A2(n15764), .ZN(n20500) );
  AOI21_X1 U18759 ( .B1(n15771), .B2(n15766), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n15767) );
  AOI221_X1 U18760 ( .B1(n15769), .B2(n15768), .C1(n20500), .C2(n15768), .A(
        n15767), .ZN(P1_U3162) );
  OAI21_X1 U18761 ( .B1(n15771), .B2(n20294), .A(n15770), .ZN(P1_U3466) );
  AOI21_X1 U18762 ( .B1(n15774), .B2(n15773), .A(n15772), .ZN(n15782) );
  INV_X1 U18763 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19566) );
  OAI22_X1 U18764 ( .A1(n18810), .A2(n19566), .B1(n15775), .B2(n18694), .ZN(
        n15778) );
  NOR2_X1 U18765 ( .A1(n15776), .A2(n18795), .ZN(n15777) );
  AOI211_X1 U18766 ( .C1(P2_EBX_REG_29__SCAN_IN), .C2(n18819), .A(n15778), .B(
        n15777), .ZN(n15779) );
  OAI21_X1 U18767 ( .B1(n15780), .B2(n18789), .A(n15779), .ZN(n15781) );
  AOI21_X1 U18768 ( .B1(n19499), .B2(n15782), .A(n15781), .ZN(n15783) );
  OAI21_X1 U18769 ( .B1(n15784), .B2(n18812), .A(n15783), .ZN(P2_U2826) );
  AOI211_X1 U18770 ( .C1(n15787), .C2(n15786), .A(n15785), .B(n18779), .ZN(
        n15796) );
  NAND2_X1 U18771 ( .A1(n15788), .A2(n18814), .ZN(n15793) );
  INV_X1 U18772 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15789) );
  OAI22_X1 U18773 ( .A1(n18810), .A2(n15790), .B1(n15789), .B2(n18694), .ZN(
        n15791) );
  AOI21_X1 U18774 ( .B1(n18819), .B2(P2_EBX_REG_26__SCAN_IN), .A(n15791), .ZN(
        n15792) );
  OAI211_X1 U18775 ( .C1(n18795), .C2(n15794), .A(n15793), .B(n15792), .ZN(
        n15795) );
  AOI211_X1 U18776 ( .C1(n15802), .C2(n15797), .A(n15796), .B(n15795), .ZN(
        n15798) );
  INV_X1 U18777 ( .A(n15798), .ZN(P2_U2829) );
  INV_X1 U18778 ( .A(n15799), .ZN(n15800) );
  AOI22_X1 U18779 ( .A1(n15800), .A2(n18818), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n9607), .ZN(n15811) );
  AOI22_X1 U18780 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n18819), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18669), .ZN(n15810) );
  INV_X1 U18781 ( .A(n15848), .ZN(n15803) );
  AOI22_X1 U18782 ( .A1(n15803), .A2(n18814), .B1(n15802), .B2(n15801), .ZN(
        n15809) );
  AOI21_X1 U18783 ( .B1(n15806), .B2(n15805), .A(n15804), .ZN(n15807) );
  NAND2_X1 U18784 ( .A1(n19499), .A2(n15807), .ZN(n15808) );
  NAND4_X1 U18785 ( .A1(n15811), .A2(n15810), .A3(n15809), .A4(n15808), .ZN(
        P2_U2831) );
  AOI22_X1 U18786 ( .A1(n18859), .A2(n15813), .B1(n15812), .B2(n18875), .ZN(
        P2_U2856) );
  AOI22_X1 U18787 ( .A1(n15814), .A2(n18871), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n18875), .ZN(n15815) );
  OAI21_X1 U18788 ( .B1(n18875), .B2(n15816), .A(n15815), .ZN(P2_U2864) );
  AOI21_X1 U18789 ( .B1(n15817), .B2(n13669), .A(n11429), .ZN(n15830) );
  AOI22_X1 U18790 ( .A1(n15830), .A2(n18871), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n18875), .ZN(n15818) );
  OAI21_X1 U18791 ( .B1(n18875), .B2(n15819), .A(n15818), .ZN(P2_U2865) );
  AOI21_X1 U18792 ( .B1(n15820), .B2(n13612), .A(n9654), .ZN(n15836) );
  AOI22_X1 U18793 ( .A1(n15836), .A2(n18871), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n18875), .ZN(n15821) );
  OAI21_X1 U18794 ( .B1(n18875), .B2(n15822), .A(n15821), .ZN(P2_U2867) );
  INV_X1 U18795 ( .A(n15823), .ZN(n15826) );
  INV_X1 U18796 ( .A(n13552), .ZN(n15825) );
  AOI21_X1 U18797 ( .B1(n15826), .B2(n15825), .A(n15824), .ZN(n15842) );
  AOI22_X1 U18798 ( .A1(n15842), .A2(n18871), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n18875), .ZN(n15827) );
  OAI21_X1 U18799 ( .B1(n18875), .B2(n18671), .A(n15827), .ZN(P2_U2869) );
  AOI22_X1 U18800 ( .A1(n18880), .A2(n15828), .B1(n18893), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n15833) );
  AOI22_X1 U18801 ( .A1(n18882), .A2(BUF1_REG_22__SCAN_IN), .B1(n18881), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n15832) );
  AOI22_X1 U18802 ( .A1(n15830), .A2(n18885), .B1(n18884), .B2(n15829), .ZN(
        n15831) );
  NAND3_X1 U18803 ( .A1(n15833), .A2(n15832), .A3(n15831), .ZN(P2_U2897) );
  AOI22_X1 U18804 ( .A1(n18880), .A2(n15834), .B1(n18893), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n15839) );
  AOI22_X1 U18805 ( .A1(n18882), .A2(BUF1_REG_20__SCAN_IN), .B1(n18881), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n15838) );
  AOI22_X1 U18806 ( .A1(n15836), .A2(n18885), .B1(n18884), .B2(n15835), .ZN(
        n15837) );
  NAND3_X1 U18807 ( .A1(n15839), .A2(n15838), .A3(n15837), .ZN(P2_U2899) );
  AOI22_X1 U18808 ( .A1(n18880), .A2(n15840), .B1(n18893), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n15845) );
  AOI22_X1 U18809 ( .A1(n18882), .A2(BUF1_REG_18__SCAN_IN), .B1(n18881), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n15844) );
  INV_X1 U18810 ( .A(n18670), .ZN(n15841) );
  AOI22_X1 U18811 ( .A1(n15842), .A2(n18885), .B1(n18884), .B2(n15841), .ZN(
        n15843) );
  NAND3_X1 U18812 ( .A1(n15845), .A2(n15844), .A3(n15843), .ZN(P2_U2901) );
  AOI22_X1 U18813 ( .A1(n18934), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18933), .ZN(n15853) );
  NOR3_X1 U18814 ( .A1(n15847), .A2(n15846), .A3(n15941), .ZN(n15850) );
  NOR2_X1 U18815 ( .A1(n15848), .A2(n15859), .ZN(n15849) );
  AOI211_X1 U18816 ( .C1(n15851), .C2(n18936), .A(n15850), .B(n15849), .ZN(
        n15852) );
  OAI211_X1 U18817 ( .C1(n18944), .C2(n15854), .A(n15853), .B(n15852), .ZN(
        P2_U2990) );
  AOI22_X1 U18818 ( .A1(n18934), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n18933), .ZN(n15862) );
  NAND2_X1 U18819 ( .A1(n15855), .A2(n18936), .ZN(n15858) );
  NAND2_X1 U18820 ( .A1(n15856), .A2(n18939), .ZN(n15857) );
  OAI211_X1 U18821 ( .C1(n15859), .C2(n18671), .A(n15858), .B(n15857), .ZN(
        n15860) );
  INV_X1 U18822 ( .A(n15860), .ZN(n15861) );
  OAI211_X1 U18823 ( .C1(n18944), .C2(n18665), .A(n15862), .B(n15861), .ZN(
        P2_U2996) );
  AOI22_X1 U18824 ( .A1(n18934), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n18933), .ZN(n15867) );
  AOI222_X1 U18825 ( .A1(n15865), .A2(n18936), .B1(n18939), .B2(n15864), .C1(
        n18938), .C2(n15863), .ZN(n15866) );
  OAI211_X1 U18826 ( .C1(n18944), .C2(n18716), .A(n15867), .B(n15866), .ZN(
        P2_U3000) );
  AOI22_X1 U18827 ( .A1(n18934), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n18933), .ZN(n15877) );
  XNOR2_X1 U18828 ( .A(n15869), .B(n15872), .ZN(n15870) );
  XNOR2_X1 U18829 ( .A(n15868), .B(n15870), .ZN(n15974) );
  INV_X1 U18830 ( .A(n15878), .ZN(n15871) );
  AOI21_X1 U18831 ( .B1(n15872), .B2(n15871), .A(n9608), .ZN(n15973) );
  OAI21_X1 U18832 ( .B1(n15875), .B2(n15874), .A(n15873), .ZN(n18851) );
  INV_X1 U18833 ( .A(n18851), .ZN(n15972) );
  AOI222_X1 U18834 ( .A1(n15974), .A2(n18936), .B1(n18939), .B2(n15973), .C1(
        n18938), .C2(n15972), .ZN(n15876) );
  OAI211_X1 U18835 ( .C1(n18944), .C2(n18728), .A(n15877), .B(n15876), .ZN(
        P2_U3002) );
  AOI22_X1 U18836 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n18933), .B1(n15948), 
        .B2(n18741), .ZN(n15887) );
  AOI21_X1 U18837 ( .B1(n15980), .B2(n15896), .A(n15878), .ZN(n15983) );
  NOR2_X1 U18838 ( .A1(n9678), .A2(n15879), .ZN(n15883) );
  NOR2_X1 U18839 ( .A1(n15881), .A2(n15880), .ZN(n15882) );
  XNOR2_X1 U18840 ( .A(n15883), .B(n15882), .ZN(n15984) );
  AOI22_X1 U18841 ( .A1(n15983), .A2(n18939), .B1(n18936), .B2(n15984), .ZN(
        n15884) );
  INV_X1 U18842 ( .A(n15884), .ZN(n15885) );
  AOI21_X1 U18843 ( .B1(n18938), .B2(n18742), .A(n15885), .ZN(n15886) );
  OAI211_X1 U18844 ( .C1(n15957), .C2(n15888), .A(n15887), .B(n15886), .ZN(
        P2_U3003) );
  AOI22_X1 U18845 ( .A1(n18934), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n18933), .ZN(n15904) );
  AND2_X1 U18846 ( .A1(n15889), .A2(n9700), .ZN(n15891) );
  INV_X1 U18847 ( .A(n15890), .ZN(n15910) );
  NOR2_X1 U18848 ( .A1(n15891), .A2(n15910), .ZN(n15895) );
  NAND2_X1 U18849 ( .A1(n15893), .A2(n15892), .ZN(n15894) );
  XNOR2_X1 U18850 ( .A(n15895), .B(n15894), .ZN(n15996) );
  INV_X1 U18851 ( .A(n15996), .ZN(n15902) );
  INV_X1 U18852 ( .A(n15896), .ZN(n15897) );
  AOI21_X1 U18853 ( .B1(n20808), .B2(n15906), .A(n15897), .ZN(n15993) );
  OR2_X1 U18854 ( .A1(n15899), .A2(n15898), .ZN(n15901) );
  AND2_X1 U18855 ( .A1(n15901), .A2(n15900), .ZN(n18856) );
  AOI222_X1 U18856 ( .A1(n15902), .A2(n18936), .B1(n18939), .B2(n15993), .C1(
        n18938), .C2(n18856), .ZN(n15903) );
  OAI211_X1 U18857 ( .C1(n18944), .C2(n18749), .A(n15904), .B(n15903), .ZN(
        P2_U3004) );
  AOI22_X1 U18858 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n18933), .B1(n15948), 
        .B2(n18763), .ZN(n15916) );
  OR2_X1 U18859 ( .A1(n15905), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15907) );
  AND2_X1 U18860 ( .A1(n15907), .A2(n15906), .ZN(n16004) );
  INV_X1 U18861 ( .A(n16004), .ZN(n15913) );
  NAND2_X1 U18862 ( .A1(n15889), .A2(n15908), .ZN(n15912) );
  OR2_X1 U18863 ( .A1(n15910), .A2(n15909), .ZN(n15911) );
  XNOR2_X1 U18864 ( .A(n15912), .B(n15911), .ZN(n16002) );
  OAI22_X1 U18865 ( .A1(n15913), .A2(n15941), .B1(n15942), .B2(n16002), .ZN(
        n15914) );
  AOI21_X1 U18866 ( .B1(n18938), .B2(n18764), .A(n15914), .ZN(n15915) );
  OAI211_X1 U18867 ( .C1(n15957), .C2(n15917), .A(n15916), .B(n15915), .ZN(
        P2_U3005) );
  AOI22_X1 U18868 ( .A1(n18934), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n18933), .ZN(n15929) );
  AOI21_X1 U18869 ( .B1(n13602), .B2(n15919), .A(n15918), .ZN(n15924) );
  INV_X1 U18870 ( .A(n15920), .ZN(n15922) );
  NOR2_X1 U18871 ( .A1(n15922), .A2(n15921), .ZN(n15923) );
  XNOR2_X1 U18872 ( .A(n15924), .B(n15923), .ZN(n16020) );
  XOR2_X1 U18873 ( .A(n15926), .B(n15925), .Z(n16017) );
  INV_X1 U18874 ( .A(n18870), .ZN(n15927) );
  AOI222_X1 U18875 ( .A1(n16020), .A2(n18936), .B1(n18939), .B2(n16017), .C1(
        n18938), .C2(n15927), .ZN(n15928) );
  OAI211_X1 U18876 ( .C1(n18944), .C2(n15930), .A(n15929), .B(n15928), .ZN(
        P2_U3006) );
  AOI22_X1 U18877 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n18933), .B1(n15948), 
        .B2(n18803), .ZN(n15945) );
  XNOR2_X1 U18878 ( .A(n15931), .B(n15932), .ZN(n16038) );
  OR2_X1 U18879 ( .A1(n15934), .A2(n15933), .ZN(n15940) );
  AND2_X1 U18880 ( .A1(n15936), .A2(n15935), .ZN(n15938) );
  OR2_X1 U18881 ( .A1(n15938), .A2(n15937), .ZN(n15939) );
  NAND2_X1 U18882 ( .A1(n15940), .A2(n15939), .ZN(n16048) );
  OAI22_X1 U18883 ( .A1(n16038), .A2(n15942), .B1(n16048), .B2(n15941), .ZN(
        n15943) );
  AOI21_X1 U18884 ( .B1(n18938), .B2(n18804), .A(n15943), .ZN(n15944) );
  OAI211_X1 U18885 ( .C1(n15957), .C2(n15946), .A(n15945), .B(n15944), .ZN(
        P2_U3009) );
  AOI22_X1 U18886 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n18933), .B1(n15948), 
        .B2(n15947), .ZN(n15956) );
  OAI21_X1 U18887 ( .B1(n15949), .B2(n10123), .A(n15950), .ZN(n16061) );
  INV_X1 U18888 ( .A(n16061), .ZN(n15953) );
  XOR2_X1 U18889 ( .A(n15952), .B(n15951), .Z(n16064) );
  AOI222_X1 U18890 ( .A1(n15954), .A2(n18938), .B1(n18939), .B2(n15953), .C1(
        n16064), .C2(n18936), .ZN(n15955) );
  OAI211_X1 U18891 ( .C1(n15958), .C2(n15957), .A(n15956), .B(n15955), .ZN(
        P2_U3011) );
  INV_X1 U18892 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19542) );
  NOR2_X1 U18893 ( .A1(n19542), .A2(n16010), .ZN(n15961) );
  OAI22_X1 U18894 ( .A1(n15959), .A2(n15962), .B1(n16053), .B2(n18709), .ZN(
        n15960) );
  AOI211_X1 U18895 ( .C1(n15963), .C2(n15962), .A(n15961), .B(n15960), .ZN(
        n15966) );
  AOI22_X1 U18896 ( .A1(n15964), .A2(n16033), .B1(n16045), .B2(n18708), .ZN(
        n15965) );
  OAI211_X1 U18897 ( .C1(n15967), .C2(n16037), .A(n15966), .B(n15965), .ZN(
        P2_U3031) );
  XNOR2_X1 U18898 ( .A(n13183), .B(n15968), .ZN(n18892) );
  NOR2_X1 U18899 ( .A1(n11092), .A2(n16010), .ZN(n15969) );
  AOI211_X1 U18900 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15971), .A(
        n15970), .B(n15969), .ZN(n15976) );
  AOI222_X1 U18901 ( .A1(n15974), .A2(n16063), .B1(n16033), .B2(n15973), .C1(
        n16045), .C2(n15972), .ZN(n15975) );
  OAI211_X1 U18902 ( .C1(n16053), .C2(n18892), .A(n15976), .B(n15975), .ZN(
        P2_U3034) );
  OAI21_X1 U18903 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15978), .A(
        n15977), .ZN(n15992) );
  NOR2_X1 U18904 ( .A1(n11088), .A2(n16010), .ZN(n15982) );
  NAND2_X1 U18905 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16000), .ZN(
        n15989) );
  AOI211_X1 U18906 ( .C1(n20808), .C2(n15980), .A(n15979), .B(n15989), .ZN(
        n15981) );
  AOI211_X1 U18907 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15992), .A(
        n15982), .B(n15981), .ZN(n15986) );
  AOI222_X1 U18908 ( .A1(n15984), .A2(n16063), .B1(n16033), .B2(n15983), .C1(
        n16045), .C2(n18742), .ZN(n15985) );
  OAI211_X1 U18909 ( .C1(n16053), .C2(n18746), .A(n15986), .B(n15985), .ZN(
        P2_U3035) );
  NOR2_X1 U18910 ( .A1(n10939), .A2(n16010), .ZN(n15991) );
  XNOR2_X1 U18911 ( .A(n15988), .B(n15987), .ZN(n18897) );
  OAI22_X1 U18912 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15989), .B1(
        n18897), .B2(n16053), .ZN(n15990) );
  AOI211_X1 U18913 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n15992), .A(
        n15991), .B(n15990), .ZN(n15995) );
  AOI22_X1 U18914 ( .A1(n15993), .A2(n16033), .B1(n16045), .B2(n18856), .ZN(
        n15994) );
  OAI211_X1 U18915 ( .C1(n15996), .C2(n16037), .A(n15995), .B(n15994), .ZN(
        P2_U3036) );
  INV_X1 U18916 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19535) );
  NOR2_X1 U18917 ( .A1(n19535), .A2(n16010), .ZN(n15997) );
  AOI221_X1 U18918 ( .B1(n16000), .B2(n15999), .C1(n15998), .C2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15997), .ZN(n16006) );
  OAI22_X1 U18919 ( .A1(n16002), .A2(n16037), .B1(n16055), .B2(n16001), .ZN(
        n16003) );
  AOI21_X1 U18920 ( .B1(n16004), .B2(n16033), .A(n16003), .ZN(n16005) );
  OAI211_X1 U18921 ( .C1(n16053), .C2(n18768), .A(n16006), .B(n16005), .ZN(
        P2_U3037) );
  INV_X1 U18922 ( .A(n16011), .ZN(n16027) );
  NAND2_X1 U18923 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16009) );
  INV_X1 U18924 ( .A(n16007), .ZN(n16008) );
  AOI21_X1 U18925 ( .B1(n16027), .B2(n16009), .A(n16008), .ZN(n16028) );
  NOR2_X1 U18926 ( .A1(n13323), .A2(n16010), .ZN(n16015) );
  NOR4_X1 U18927 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n16013), .A3(
        n16012), .A4(n16011), .ZN(n16014) );
  AOI211_X1 U18928 ( .C1(n16057), .C2(n16016), .A(n16015), .B(n16014), .ZN(
        n16022) );
  INV_X1 U18929 ( .A(n16017), .ZN(n16018) );
  OAI22_X1 U18930 ( .A1(n16018), .A2(n16060), .B1(n16055), .B2(n18870), .ZN(
        n16019) );
  AOI21_X1 U18931 ( .B1(n16063), .B2(n16020), .A(n16019), .ZN(n16021) );
  OAI211_X1 U18932 ( .C1(n16028), .C2(n16023), .A(n16022), .B(n16021), .ZN(
        P2_U3038) );
  INV_X1 U18933 ( .A(n18774), .ZN(n16025) );
  AOI22_X1 U18934 ( .A1(n16045), .A2(n16025), .B1(n18933), .B2(
        P2_REIP_REG_7__SCAN_IN), .ZN(n16035) );
  INV_X1 U18935 ( .A(n16026), .ZN(n16030) );
  AOI21_X1 U18936 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16027), .A(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16029) );
  OAI22_X1 U18937 ( .A1(n16030), .A2(n16037), .B1(n16029), .B2(n16028), .ZN(
        n16031) );
  AOI21_X1 U18938 ( .B1(n16033), .B2(n16032), .A(n16031), .ZN(n16034) );
  OAI211_X1 U18939 ( .C1(n16053), .C2(n18775), .A(n16035), .B(n16034), .ZN(
        P2_U3039) );
  AOI22_X1 U18940 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16036), .B1(
        P2_REIP_REG_5__SCAN_IN), .B2(n18933), .ZN(n16052) );
  NOR2_X1 U18941 ( .A1(n16038), .A2(n16037), .ZN(n16050) );
  INV_X1 U18942 ( .A(n16039), .ZN(n16040) );
  AOI211_X1 U18943 ( .C1(n16043), .C2(n16042), .A(n16041), .B(n16040), .ZN(
        n16044) );
  INV_X1 U18944 ( .A(n16044), .ZN(n16047) );
  NAND2_X1 U18945 ( .A1(n16045), .A2(n18804), .ZN(n16046) );
  OAI211_X1 U18946 ( .C1(n16048), .C2(n16060), .A(n16047), .B(n16046), .ZN(
        n16049) );
  NOR2_X1 U18947 ( .A1(n16050), .A2(n16049), .ZN(n16051) );
  OAI211_X1 U18948 ( .C1(n16053), .C2(n18808), .A(n16052), .B(n16051), .ZN(
        P2_U3041) );
  OAI22_X1 U18949 ( .A1(n12893), .A2(n16055), .B1(n16054), .B2(n11181), .ZN(
        n16056) );
  AOI21_X1 U18950 ( .B1(n16058), .B2(n16057), .A(n16056), .ZN(n16059) );
  OAI21_X1 U18951 ( .B1(n16061), .B2(n16060), .A(n16059), .ZN(n16062) );
  AOI21_X1 U18952 ( .B1(n16064), .B2(n16063), .A(n16062), .ZN(n16065) );
  OAI221_X1 U18953 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16068), .C1(
        n16067), .C2(n16066), .A(n16065), .ZN(P2_U3043) );
  NAND2_X1 U18954 ( .A1(n16085), .A2(n9783), .ZN(n16069) );
  OAI21_X1 U18955 ( .B1(n16070), .B2(n16085), .A(n16069), .ZN(n16084) );
  INV_X1 U18956 ( .A(n16085), .ZN(n16071) );
  MUX2_X1 U18957 ( .A(n16072), .B(n16073), .S(n16071), .Z(n16083) );
  INV_X1 U18958 ( .A(n19044), .ZN(n19020) );
  INV_X1 U18959 ( .A(n16083), .ZN(n16081) );
  INV_X1 U18960 ( .A(n16073), .ZN(n16078) );
  AOI21_X1 U18961 ( .B1(n16075), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16085), .ZN(n16077) );
  OAI211_X1 U18962 ( .C1(n16075), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16074), .B(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n16076) );
  OAI211_X1 U18963 ( .C1(n16078), .C2(n19596), .A(n16077), .B(n16076), .ZN(
        n16079) );
  AOI222_X1 U18964 ( .A1(n16084), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .B1(n16084), .B2(n16079), .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .C2(n16079), .ZN(n16080) );
  AOI21_X1 U18965 ( .B1(n19020), .B2(n16081), .A(n16080), .ZN(n16082) );
  OAI22_X1 U18966 ( .A1(n16084), .A2(n16083), .B1(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n16082), .ZN(n16105) );
  NAND2_X1 U18967 ( .A1(n16085), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n16103) );
  INV_X1 U18968 ( .A(n16086), .ZN(n16088) );
  AOI22_X1 U18969 ( .A1(n16090), .A2(n16089), .B1(n16088), .B2(n16087), .ZN(
        n16094) );
  NAND2_X1 U18970 ( .A1(n16092), .A2(n16091), .ZN(n16093) );
  AND2_X1 U18971 ( .A1(n16094), .A2(n16093), .ZN(n19621) );
  OAI21_X1 U18972 ( .B1(n16096), .B2(n10253), .A(n16095), .ZN(n16097) );
  INV_X1 U18973 ( .A(n16097), .ZN(n16102) );
  AND2_X1 U18974 ( .A1(n16098), .A2(n19504), .ZN(n16099) );
  NOR2_X1 U18975 ( .A1(n16100), .A2(n16099), .ZN(n18644) );
  OAI21_X1 U18976 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n18644), .ZN(n16101) );
  NAND4_X1 U18977 ( .A1(n16103), .A2(n19621), .A3(n16102), .A4(n16101), .ZN(
        n16104) );
  OR2_X1 U18978 ( .A1(n16105), .A2(n16104), .ZN(n16113) );
  INV_X1 U18979 ( .A(n16113), .ZN(n16119) );
  NAND2_X1 U18980 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19606), .ZN(n19497) );
  OAI21_X1 U18981 ( .B1(n16108), .B2(n16107), .A(n16106), .ZN(n16112) );
  OAI21_X1 U18982 ( .B1(n19504), .B2(n19497), .A(n16112), .ZN(n16109) );
  AOI211_X1 U18983 ( .C1(n16121), .C2(n16111), .A(n16110), .B(n16109), .ZN(
        n16118) );
  NOR2_X1 U18984 ( .A1(n16113), .A2(n16112), .ZN(n16120) );
  NOR2_X1 U18985 ( .A1(n16120), .A2(n18930), .ZN(n19500) );
  OAI21_X1 U18986 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16115), .A(n16114), 
        .ZN(n16116) );
  OAI21_X1 U18987 ( .B1(n19500), .B2(n19504), .A(n16116), .ZN(n16117) );
  OAI211_X1 U18988 ( .C1(n16119), .C2(n19494), .A(n16118), .B(n16117), .ZN(
        P2_U3176) );
  NOR2_X1 U18989 ( .A1(n16120), .A2(n18640), .ZN(n16123) );
  INV_X1 U18990 ( .A(n16121), .ZN(n16122) );
  OAI21_X1 U18991 ( .B1(n16123), .B2(n19582), .A(n16122), .ZN(P2_U3593) );
  NAND3_X1 U18992 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16141), .A3(
        n16124), .ZN(n16125) );
  XOR2_X1 U18993 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n16125), .Z(
        n16187) );
  NOR2_X2 U18994 ( .A1(n17188), .A2(n16308), .ZN(n17613) );
  INV_X1 U18995 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17620) );
  NAND4_X1 U18996 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16341) );
  NAND2_X1 U18997 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17458) );
  NOR2_X1 U18998 ( .A1(n17458), .A2(n17443), .ZN(n17416) );
  NAND2_X1 U18999 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17419) );
  NAND2_X1 U19000 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17380) );
  NAND2_X1 U19001 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17366), .ZN(
        n17345) );
  NAND2_X1 U19002 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17346) );
  NAND2_X1 U19003 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17297) );
  NAND2_X1 U19004 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17260) );
  NAND2_X1 U19005 ( .A1(n16163), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16127) );
  INV_X1 U19006 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18551) );
  NOR2_X1 U19007 ( .A1(n18551), .A2(n17861), .ZN(n16181) );
  NOR2_X1 U19008 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18468), .ZN(n17455) );
  NAND2_X1 U19009 ( .A1(n18253), .A2(n18115), .ZN(n18302) );
  OAI21_X1 U19010 ( .B1(n17620), .B2(n17365), .A(n18302), .ZN(n17417) );
  INV_X1 U19011 ( .A(n17417), .ZN(n17379) );
  OR2_X1 U19012 ( .A1(n16128), .A2(n17379), .ZN(n16153) );
  INV_X1 U19013 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16130) );
  XOR2_X1 U19014 ( .A(n16130), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16131) );
  NOR2_X1 U19015 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17365), .ZN(
        n16164) );
  NOR2_X1 U19016 ( .A1(n17620), .A2(n17259), .ZN(n16334) );
  INV_X1 U19017 ( .A(n16334), .ZN(n16333) );
  NOR2_X1 U19018 ( .A1(n17260), .A2(n16333), .ZN(n16162) );
  INV_X1 U19019 ( .A(n17455), .ZN(n17624) );
  NAND2_X1 U19020 ( .A1(n18000), .A2(n16128), .ZN(n16129) );
  OAI211_X1 U19021 ( .C1(n16162), .C2(n17624), .A(n17625), .B(n16129), .ZN(
        n16165) );
  NOR2_X1 U19022 ( .A1(n16164), .A2(n16165), .ZN(n16151) );
  OAI22_X1 U19023 ( .A1(n16153), .A2(n16131), .B1(n16151), .B2(n16130), .ZN(
        n16132) );
  AOI211_X1 U19024 ( .C1(n17482), .C2(n16342), .A(n16181), .B(n16132), .ZN(
        n16148) );
  INV_X1 U19025 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18578) );
  AOI22_X1 U19026 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17516), .B1(
        n17534), .B2(n18578), .ZN(n16140) );
  OAI22_X1 U19027 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16134), .B1(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16135), .ZN(n16139) );
  NAND2_X1 U19028 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16142), .ZN(
        n16179) );
  OAI21_X1 U19029 ( .B1(n16135), .B2(n16134), .A(n16179), .ZN(n16137) );
  NAND2_X1 U19030 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18578), .ZN(
        n16136) );
  NAND3_X1 U19031 ( .A1(n16140), .A2(n16137), .A3(n16136), .ZN(n16138) );
  OAI21_X1 U19032 ( .B1(n16140), .B2(n16139), .A(n16138), .ZN(n16184) );
  NAND3_X1 U19033 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16141), .A3(
        n18578), .ZN(n16178) );
  OAI21_X1 U19034 ( .B1(n16142), .B2(n16161), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16143) );
  OAI21_X1 U19035 ( .B1(n16178), .B2(n17632), .A(n16143), .ZN(n16183) );
  INV_X1 U19036 ( .A(n16183), .ZN(n16145) );
  OAI211_X1 U19037 ( .C1(n16187), .C2(n17629), .A(n16148), .B(n16147), .ZN(
        P3_U2799) );
  AOI22_X1 U19038 ( .A1(n17823), .A2(n17613), .B1(n17452), .B2(n9640), .ZN(
        n17522) );
  NAND2_X1 U19039 ( .A1(n16149), .A2(n17406), .ZN(n17280) );
  XOR2_X1 U19040 ( .A(n16163), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16354) );
  INV_X1 U19041 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16152) );
  NAND2_X1 U19042 ( .A1(n17951), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16150) );
  OAI221_X1 U19043 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16153), .C1(
        n16152), .C2(n16151), .A(n16150), .ZN(n16154) );
  AOI21_X1 U19044 ( .B1(n17482), .B2(n16354), .A(n16154), .ZN(n16159) );
  OAI22_X1 U19045 ( .A1(n16171), .A2(n17629), .B1(n16155), .B2(n16144), .ZN(
        n16157) );
  AOI22_X1 U19046 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16157), .B1(
        n17535), .B2(n16156), .ZN(n16158) );
  OAI211_X1 U19047 ( .C1(n16160), .C2(n17280), .A(n16159), .B(n16158), .ZN(
        P3_U2800) );
  NOR2_X1 U19048 ( .A1(n16170), .A2(n17632), .ZN(n16203) );
  OAI211_X1 U19049 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16203), .A(
        n17452), .B(n16161), .ZN(n16168) );
  INV_X1 U19050 ( .A(n16162), .ZN(n16331) );
  AOI21_X1 U19051 ( .B1(n9874), .B2(n16331), .A(n16163), .ZN(n16362) );
  OAI21_X1 U19052 ( .B1(n17482), .B2(n16164), .A(n16362), .ZN(n16167) );
  OAI221_X1 U19053 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n9746), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n18000), .A(n16165), .ZN(
        n16166) );
  NAND4_X1 U19054 ( .A1(n16169), .A2(n16168), .A3(n16167), .A4(n16166), .ZN(
        n16174) );
  OR2_X1 U19055 ( .A1(n17633), .A2(n16170), .ZN(n16199) );
  AOI211_X1 U19056 ( .C1(n16172), .C2(n16199), .A(n16171), .B(n17629), .ZN(
        n16173) );
  NOR2_X1 U19057 ( .A1(n16174), .A2(n16173), .ZN(n16175) );
  OAI21_X1 U19058 ( .B1(n16176), .B2(n17508), .A(n16175), .ZN(P3_U2801) );
  OAI22_X1 U19059 ( .A1(n16179), .A2(n17943), .B1(n16178), .B2(n16177), .ZN(
        n16180) );
  AOI211_X1 U19060 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16182), .A(
        n16181), .B(n16180), .ZN(n16186) );
  AOI22_X1 U19061 ( .A1(n17870), .A2(n16184), .B1(n17794), .B2(n16183), .ZN(
        n16185) );
  OAI211_X1 U19062 ( .C1(n16187), .C2(n17914), .A(n16186), .B(n16185), .ZN(
        P3_U2831) );
  NOR2_X1 U19063 ( .A1(n18425), .A2(n16195), .ZN(n17805) );
  AOI22_X1 U19064 ( .A1(n18428), .A2(n17823), .B1(n9640), .B2(n17805), .ZN(
        n17743) );
  AOI21_X1 U19065 ( .B1(n18400), .B2(n18595), .A(n18399), .ZN(n17924) );
  AOI21_X1 U19066 ( .B1(n17697), .B2(n17924), .A(n16188), .ZN(n17653) );
  OAI21_X1 U19067 ( .B1(n17743), .B2(n17745), .A(n17653), .ZN(n17645) );
  NAND2_X1 U19068 ( .A1(n17952), .A2(n17645), .ZN(n17715) );
  NAND2_X1 U19069 ( .A1(n16189), .A2(n16204), .ZN(n17269) );
  AOI21_X1 U19070 ( .B1(n17534), .B2(n16190), .A(n17270), .ZN(n17258) );
  AOI22_X1 U19071 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17516), .B1(
        n17534), .B2(n16204), .ZN(n17257) );
  NOR2_X1 U19072 ( .A1(n17258), .A2(n17257), .ZN(n17256) );
  NAND2_X1 U19073 ( .A1(n17270), .A2(n17257), .ZN(n16192) );
  OAI21_X1 U19074 ( .B1(n17256), .B2(n10119), .A(n16192), .ZN(n16193) );
  NAND2_X1 U19075 ( .A1(n16197), .A2(n10122), .ZN(n16201) );
  INV_X1 U19076 ( .A(n17805), .ZN(n17825) );
  OR2_X1 U19077 ( .A1(n16203), .A2(n17825), .ZN(n16205) );
  AOI211_X1 U19078 ( .C1(n16206), .C2(n16205), .A(n17951), .B(n16204), .ZN(
        n16207) );
  NOR2_X1 U19079 ( .A1(n10121), .A2(n16207), .ZN(n16208) );
  NAND2_X1 U19080 ( .A1(n17951), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17261) );
  OAI211_X1 U19081 ( .C1(n17715), .C2(n17269), .A(n16208), .B(n17261), .ZN(
        P3_U2834) );
  NOR3_X1 U19082 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16210) );
  NOR4_X1 U19083 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16209) );
  NAND4_X1 U19084 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16210), .A3(n16209), .A4(
        U215), .ZN(U213) );
  INV_X1 U19085 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n18899) );
  INV_X2 U19086 ( .A(U214), .ZN(n16256) );
  NOR2_X2 U19087 ( .A1(n16256), .A2(n16211), .ZN(n16254) );
  OAI222_X1 U19088 ( .A1(U212), .A2(n18899), .B1(n16259), .B2(n20776), .C1(
        U214), .C2(n20635), .ZN(U216) );
  INV_X1 U19089 ( .A(U212), .ZN(n16257) );
  AOI222_X1 U19090 ( .A1(n16257), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16254), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n16256), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n16212) );
  INV_X1 U19091 ( .A(n16212), .ZN(U217) );
  INV_X1 U19092 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16214) );
  AOI22_X1 U19093 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16256), .ZN(n16213) );
  OAI21_X1 U19094 ( .B1(n16214), .B2(n16259), .A(n16213), .ZN(U218) );
  INV_X1 U19095 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16216) );
  AOI22_X1 U19096 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16256), .ZN(n16215) );
  OAI21_X1 U19097 ( .B1(n16216), .B2(n16259), .A(n16215), .ZN(U219) );
  INV_X1 U19098 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16218) );
  AOI22_X1 U19099 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16256), .ZN(n16217) );
  OAI21_X1 U19100 ( .B1(n16218), .B2(n16259), .A(n16217), .ZN(U220) );
  INV_X1 U19101 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16220) );
  AOI22_X1 U19102 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16256), .ZN(n16219) );
  OAI21_X1 U19103 ( .B1(n16220), .B2(n16259), .A(n16219), .ZN(U221) );
  AOI222_X1 U19104 ( .A1(n16257), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(n16254), 
        .B2(BUF1_REG_25__SCAN_IN), .C1(n16256), .C2(P1_DATAO_REG_25__SCAN_IN), 
        .ZN(n16221) );
  INV_X1 U19105 ( .A(n16221), .ZN(U222) );
  INV_X1 U19106 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16223) );
  AOI22_X1 U19107 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16256), .ZN(n16222) );
  OAI21_X1 U19108 ( .B1(n16223), .B2(n16259), .A(n16222), .ZN(U223) );
  INV_X1 U19109 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n18987) );
  AOI22_X1 U19110 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16256), .ZN(n16224) );
  OAI21_X1 U19111 ( .B1(n18987), .B2(n16259), .A(n16224), .ZN(U224) );
  INV_X1 U19112 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n18974) );
  AOI22_X1 U19113 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16256), .ZN(n16225) );
  OAI21_X1 U19114 ( .B1(n18974), .B2(n16259), .A(n16225), .ZN(U225) );
  AOI22_X1 U19115 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16256), .ZN(n16226) );
  OAI21_X1 U19116 ( .B1(n14176), .B2(n16259), .A(n16226), .ZN(U226) );
  INV_X1 U19117 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16228) );
  AOI22_X1 U19118 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16256), .ZN(n16227) );
  OAI21_X1 U19119 ( .B1(n16228), .B2(n16259), .A(n16227), .ZN(U227) );
  AOI222_X1 U19120 ( .A1(n16257), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n16254), 
        .B2(BUF1_REG_19__SCAN_IN), .C1(n16256), .C2(P1_DATAO_REG_19__SCAN_IN), 
        .ZN(n16229) );
  INV_X1 U19121 ( .A(n16229), .ZN(U228) );
  INV_X1 U19122 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16231) );
  AOI22_X1 U19123 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16256), .ZN(n16230) );
  OAI21_X1 U19124 ( .B1(n16231), .B2(n16259), .A(n16230), .ZN(U229) );
  INV_X1 U19125 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n18954) );
  AOI22_X1 U19126 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16256), .ZN(n16232) );
  OAI21_X1 U19127 ( .B1(n18954), .B2(n16259), .A(n16232), .ZN(U230) );
  INV_X1 U19128 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n18948) );
  AOI22_X1 U19129 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16256), .ZN(n16233) );
  OAI21_X1 U19130 ( .B1(n18948), .B2(n16259), .A(n16233), .ZN(U231) );
  INV_X1 U19131 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n19746) );
  AOI22_X1 U19132 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n16254), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16257), .ZN(n16234) );
  OAI21_X1 U19133 ( .B1(n19746), .B2(U214), .A(n16234), .ZN(U232) );
  INV_X1 U19134 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16275) );
  AOI22_X1 U19135 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16254), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16256), .ZN(n16235) );
  OAI21_X1 U19136 ( .B1(n16275), .B2(U212), .A(n16235), .ZN(U233) );
  INV_X1 U19137 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16273) );
  AOI22_X1 U19138 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16254), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16256), .ZN(n16236) );
  OAI21_X1 U19139 ( .B1(n16273), .B2(U212), .A(n16236), .ZN(U234) );
  AOI22_X1 U19140 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16256), .ZN(n16237) );
  OAI21_X1 U19141 ( .B1(n16238), .B2(n16259), .A(n16237), .ZN(U235) );
  INV_X1 U19142 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n20646) );
  AOI22_X1 U19143 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16254), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16256), .ZN(n16239) );
  OAI21_X1 U19144 ( .B1(n20646), .B2(U212), .A(n16239), .ZN(U236) );
  INV_X1 U19145 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16241) );
  AOI22_X1 U19146 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16256), .ZN(n16240) );
  OAI21_X1 U19147 ( .B1(n16241), .B2(n16259), .A(n16240), .ZN(U237) );
  INV_X1 U19148 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16269) );
  AOI22_X1 U19149 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16254), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16256), .ZN(n16242) );
  OAI21_X1 U19150 ( .B1(n16269), .B2(U212), .A(n16242), .ZN(U238) );
  AOI22_X1 U19151 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16256), .ZN(n16243) );
  OAI21_X1 U19152 ( .B1(n16244), .B2(n16259), .A(n16243), .ZN(U239) );
  INV_X1 U19153 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16267) );
  AOI22_X1 U19154 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16254), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16256), .ZN(n16245) );
  OAI21_X1 U19155 ( .B1(n16267), .B2(U212), .A(n16245), .ZN(U240) );
  INV_X1 U19156 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16247) );
  AOI22_X1 U19157 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16256), .ZN(n16246) );
  OAI21_X1 U19158 ( .B1(n16247), .B2(n16259), .A(n16246), .ZN(U241) );
  INV_X1 U19159 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16265) );
  AOI22_X1 U19160 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16254), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16256), .ZN(n16248) );
  OAI21_X1 U19161 ( .B1(n16265), .B2(U212), .A(n16248), .ZN(U242) );
  INV_X1 U19162 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16250) );
  AOI22_X1 U19163 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16256), .ZN(n16249) );
  OAI21_X1 U19164 ( .B1(n16250), .B2(n16259), .A(n16249), .ZN(U243) );
  AOI222_X1 U19165 ( .A1(n16256), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n16254), 
        .B2(BUF1_REG_3__SCAN_IN), .C1(n16257), .C2(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n16251) );
  INV_X1 U19166 ( .A(n16251), .ZN(U244) );
  AOI22_X1 U19167 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16256), .ZN(n16252) );
  OAI21_X1 U19168 ( .B1(n16253), .B2(n16259), .A(n16252), .ZN(U245) );
  INV_X1 U19169 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16262) );
  AOI22_X1 U19170 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16254), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16256), .ZN(n16255) );
  OAI21_X1 U19171 ( .B1(n16262), .B2(U212), .A(n16255), .ZN(U246) );
  AOI22_X1 U19172 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n16257), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16256), .ZN(n16258) );
  OAI21_X1 U19173 ( .B1(n16260), .B2(n16259), .A(n16258), .ZN(U247) );
  INV_X1 U19174 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16261) );
  AOI22_X1 U19175 ( .A1(n16291), .A2(n16261), .B1(n17972), .B2(U215), .ZN(U251) );
  INV_X1 U19176 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n17976) );
  AOI22_X1 U19177 ( .A1(n16291), .A2(n16262), .B1(n17976), .B2(U215), .ZN(U252) );
  INV_X1 U19178 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16263) );
  AOI22_X1 U19179 ( .A1(n16291), .A2(n16263), .B1(n17980), .B2(U215), .ZN(U253) );
  INV_X1 U19180 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n18924) );
  INV_X1 U19181 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n17984) );
  AOI22_X1 U19182 ( .A1(n16291), .A2(n18924), .B1(n17984), .B2(U215), .ZN(U254) );
  INV_X1 U19183 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16264) );
  INV_X1 U19184 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n17988) );
  AOI22_X1 U19185 ( .A1(n16291), .A2(n16264), .B1(n17988), .B2(U215), .ZN(U255) );
  INV_X1 U19186 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n17992) );
  AOI22_X1 U19187 ( .A1(n16291), .A2(n16265), .B1(n17992), .B2(U215), .ZN(U256) );
  INV_X1 U19188 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16266) );
  INV_X1 U19189 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n17996) );
  AOI22_X1 U19190 ( .A1(n16293), .A2(n16266), .B1(n17996), .B2(U215), .ZN(U257) );
  INV_X1 U19191 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18002) );
  AOI22_X1 U19192 ( .A1(n16293), .A2(n16267), .B1(n18002), .B2(U215), .ZN(U258) );
  INV_X1 U19193 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16268) );
  INV_X1 U19194 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17113) );
  AOI22_X1 U19195 ( .A1(n16291), .A2(n16268), .B1(n17113), .B2(U215), .ZN(U259) );
  INV_X1 U19196 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17107) );
  AOI22_X1 U19197 ( .A1(n16293), .A2(n16269), .B1(n17107), .B2(U215), .ZN(U260) );
  OAI22_X1 U19198 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16291), .ZN(n16270) );
  INV_X1 U19199 ( .A(n16270), .ZN(U261) );
  INV_X1 U19200 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n16271) );
  AOI22_X1 U19201 ( .A1(n16291), .A2(n20646), .B1(n16271), .B2(U215), .ZN(U262) );
  INV_X1 U19202 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16272) );
  INV_X1 U19203 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17095) );
  AOI22_X1 U19204 ( .A1(n16293), .A2(n16272), .B1(n17095), .B2(U215), .ZN(U263) );
  INV_X1 U19205 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17090) );
  AOI22_X1 U19206 ( .A1(n16291), .A2(n16273), .B1(n17090), .B2(U215), .ZN(U264) );
  INV_X1 U19207 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n16274) );
  AOI22_X1 U19208 ( .A1(n16293), .A2(n16275), .B1(n16274), .B2(U215), .ZN(U265) );
  OAI22_X1 U19209 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16291), .ZN(n16276) );
  INV_X1 U19210 ( .A(n16276), .ZN(U266) );
  INV_X1 U19211 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n16277) );
  INV_X1 U19212 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18947) );
  AOI22_X1 U19213 ( .A1(n16293), .A2(n16277), .B1(n18947), .B2(U215), .ZN(U267) );
  INV_X1 U19214 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n16278) );
  INV_X1 U19215 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n18953) );
  AOI22_X1 U19216 ( .A1(n16291), .A2(n16278), .B1(n18953), .B2(U215), .ZN(U268) );
  OAI22_X1 U19217 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16291), .ZN(n16279) );
  INV_X1 U19218 ( .A(n16279), .ZN(U269) );
  OAI22_X1 U19219 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16293), .ZN(n16280) );
  INV_X1 U19220 ( .A(n16280), .ZN(U270) );
  OAI22_X1 U19221 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16291), .ZN(n16281) );
  INV_X1 U19222 ( .A(n16281), .ZN(U271) );
  INV_X1 U19223 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16282) );
  AOI22_X1 U19224 ( .A1(n16291), .A2(n16282), .B1(n13674), .B2(U215), .ZN(U272) );
  INV_X1 U19225 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16283) );
  INV_X1 U19226 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18973) );
  AOI22_X1 U19227 ( .A1(n16291), .A2(n16283), .B1(n18973), .B2(U215), .ZN(U273) );
  INV_X1 U19228 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n16284) );
  INV_X1 U19229 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n18985) );
  AOI22_X1 U19230 ( .A1(n16291), .A2(n16284), .B1(n18985), .B2(U215), .ZN(U274) );
  OAI22_X1 U19231 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16291), .ZN(n16285) );
  INV_X1 U19232 ( .A(n16285), .ZN(U275) );
  OAI22_X1 U19233 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16293), .ZN(n16286) );
  INV_X1 U19234 ( .A(n16286), .ZN(U276) );
  OAI22_X1 U19235 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16293), .ZN(n16287) );
  INV_X1 U19236 ( .A(n16287), .ZN(U277) );
  OAI22_X1 U19237 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16291), .ZN(n16288) );
  INV_X1 U19238 ( .A(n16288), .ZN(U278) );
  OAI22_X1 U19239 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16291), .ZN(n16289) );
  INV_X1 U19240 ( .A(n16289), .ZN(U279) );
  OAI22_X1 U19241 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16291), .ZN(n16290) );
  INV_X1 U19242 ( .A(n16290), .ZN(U280) );
  OAI22_X1 U19243 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16291), .ZN(n16292) );
  INV_X1 U19244 ( .A(n16292), .ZN(U281) );
  INV_X1 U19245 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18001) );
  AOI22_X1 U19246 ( .A1(n16293), .A2(n18899), .B1(n18001), .B2(U215), .ZN(U282) );
  INV_X1 U19247 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16294) );
  AOI222_X1 U19248 ( .A1(n20635), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n18899), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16294), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16295) );
  INV_X1 U19249 ( .A(n16297), .ZN(n16296) );
  INV_X1 U19250 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18510) );
  INV_X1 U19251 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19537) );
  AOI22_X1 U19252 ( .A1(n16296), .A2(n18510), .B1(n19537), .B2(n16297), .ZN(
        U347) );
  INV_X1 U19253 ( .A(n16297), .ZN(n16298) );
  INV_X1 U19254 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n20762) );
  INV_X1 U19255 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19536) );
  AOI22_X1 U19256 ( .A1(n16298), .A2(n20762), .B1(n19536), .B2(n16297), .ZN(
        U348) );
  INV_X1 U19257 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18506) );
  INV_X1 U19258 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19534) );
  AOI22_X1 U19259 ( .A1(n16296), .A2(n18506), .B1(n19534), .B2(n16297), .ZN(
        U349) );
  INV_X1 U19260 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18505) );
  INV_X1 U19261 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19533) );
  AOI22_X1 U19262 ( .A1(n16296), .A2(n18505), .B1(n19533), .B2(n16297), .ZN(
        U350) );
  INV_X1 U19263 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18503) );
  INV_X1 U19264 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19531) );
  AOI22_X1 U19265 ( .A1(n16296), .A2(n18503), .B1(n19531), .B2(n16297), .ZN(
        U351) );
  INV_X1 U19266 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18501) );
  INV_X1 U19267 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19530) );
  AOI22_X1 U19268 ( .A1(n16296), .A2(n18501), .B1(n19530), .B2(n16297), .ZN(
        U352) );
  INV_X1 U19269 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18500) );
  INV_X1 U19270 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19529) );
  AOI22_X1 U19271 ( .A1(n16298), .A2(n18500), .B1(n19529), .B2(n16297), .ZN(
        U353) );
  INV_X1 U19272 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18498) );
  INV_X1 U19273 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19528) );
  AOI22_X1 U19274 ( .A1(n16296), .A2(n18498), .B1(n19528), .B2(n16297), .ZN(
        U354) );
  INV_X1 U19275 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18552) );
  INV_X1 U19276 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19570) );
  AOI22_X1 U19277 ( .A1(n16296), .A2(n18552), .B1(n19570), .B2(n16297), .ZN(
        U355) );
  INV_X1 U19278 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18549) );
  INV_X1 U19279 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19567) );
  AOI22_X1 U19280 ( .A1(n16296), .A2(n18549), .B1(n19567), .B2(n16297), .ZN(
        U356) );
  INV_X1 U19281 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18546) );
  INV_X1 U19282 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19565) );
  AOI22_X1 U19283 ( .A1(n16296), .A2(n18546), .B1(n19565), .B2(n16297), .ZN(
        U357) );
  INV_X1 U19284 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18545) );
  INV_X1 U19285 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19563) );
  AOI22_X1 U19286 ( .A1(n16296), .A2(n18545), .B1(n19563), .B2(n16297), .ZN(
        U358) );
  INV_X1 U19287 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18543) );
  INV_X1 U19288 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19562) );
  AOI22_X1 U19289 ( .A1(n16296), .A2(n18543), .B1(n19562), .B2(n16297), .ZN(
        U359) );
  INV_X1 U19290 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18540) );
  INV_X1 U19291 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19561) );
  AOI22_X1 U19292 ( .A1(n16296), .A2(n18540), .B1(n19561), .B2(n16297), .ZN(
        U360) );
  INV_X1 U19293 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18538) );
  INV_X1 U19294 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19559) );
  AOI22_X1 U19295 ( .A1(n16296), .A2(n18538), .B1(n19559), .B2(n16297), .ZN(
        U361) );
  INV_X1 U19296 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18535) );
  INV_X1 U19297 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19557) );
  AOI22_X1 U19298 ( .A1(n16296), .A2(n18535), .B1(n19557), .B2(n16297), .ZN(
        U362) );
  INV_X1 U19299 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18534) );
  INV_X1 U19300 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19555) );
  AOI22_X1 U19301 ( .A1(n16296), .A2(n18534), .B1(n19555), .B2(n16297), .ZN(
        U363) );
  INV_X1 U19302 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18532) );
  INV_X1 U19303 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19554) );
  AOI22_X1 U19304 ( .A1(n16296), .A2(n18532), .B1(n19554), .B2(n16297), .ZN(
        U364) );
  INV_X1 U19305 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18496) );
  INV_X1 U19306 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19527) );
  AOI22_X1 U19307 ( .A1(n16296), .A2(n18496), .B1(n19527), .B2(n16297), .ZN(
        U365) );
  INV_X1 U19308 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18529) );
  INV_X1 U19309 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19552) );
  AOI22_X1 U19310 ( .A1(n16296), .A2(n18529), .B1(n19552), .B2(n16297), .ZN(
        U366) );
  INV_X1 U19311 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18528) );
  INV_X1 U19312 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19550) );
  AOI22_X1 U19313 ( .A1(n16296), .A2(n18528), .B1(n19550), .B2(n16297), .ZN(
        U367) );
  INV_X1 U19314 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18526) );
  INV_X1 U19315 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19548) );
  AOI22_X1 U19316 ( .A1(n16296), .A2(n18526), .B1(n19548), .B2(n16297), .ZN(
        U368) );
  INV_X1 U19317 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18523) );
  INV_X1 U19318 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19546) );
  AOI22_X1 U19319 ( .A1(n16296), .A2(n18523), .B1(n19546), .B2(n16297), .ZN(
        U369) );
  INV_X1 U19320 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18522) );
  INV_X1 U19321 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19544) );
  AOI22_X1 U19322 ( .A1(n16296), .A2(n18522), .B1(n19544), .B2(n16297), .ZN(
        U370) );
  INV_X1 U19323 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18520) );
  INV_X1 U19324 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19543) );
  AOI22_X1 U19325 ( .A1(n16298), .A2(n18520), .B1(n19543), .B2(n16297), .ZN(
        U371) );
  INV_X1 U19326 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18518) );
  INV_X1 U19327 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19541) );
  AOI22_X1 U19328 ( .A1(n16298), .A2(n18518), .B1(n19541), .B2(n16297), .ZN(
        U372) );
  INV_X1 U19329 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18516) );
  INV_X1 U19330 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19540) );
  AOI22_X1 U19331 ( .A1(n16298), .A2(n18516), .B1(n19540), .B2(n16297), .ZN(
        U373) );
  INV_X1 U19332 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18514) );
  INV_X1 U19333 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19539) );
  AOI22_X1 U19334 ( .A1(n16298), .A2(n18514), .B1(n19539), .B2(n16297), .ZN(
        U374) );
  INV_X1 U19335 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18512) );
  INV_X1 U19336 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19538) );
  AOI22_X1 U19337 ( .A1(n16298), .A2(n18512), .B1(n19538), .B2(n16297), .ZN(
        U375) );
  INV_X1 U19338 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18494) );
  AOI22_X1 U19339 ( .A1(n16298), .A2(n18494), .B1(n19526), .B2(n16297), .ZN(
        U376) );
  INV_X1 U19340 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16300) );
  INV_X1 U19341 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18493) );
  NAND3_X1 U19342 ( .A1(n18493), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n16299) );
  NAND2_X1 U19343 ( .A1(n18490), .A2(n18482), .ZN(n18478) );
  NAND2_X1 U19344 ( .A1(n16299), .A2(n18478), .ZN(n18565) );
  INV_X1 U19345 ( .A(n18565), .ZN(n18562) );
  OAI21_X1 U19346 ( .B1(n18490), .B2(n16300), .A(n18562), .ZN(P3_U2633) );
  INV_X1 U19347 ( .A(n16307), .ZN(n16301) );
  NAND2_X1 U19348 ( .A1(n18615), .A2(n18424), .ZN(n17186) );
  OAI21_X1 U19349 ( .B1(n16301), .B2(n17186), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16302) );
  OAI21_X1 U19350 ( .B1(n16303), .B2(n18566), .A(n16302), .ZN(P3_U2634) );
  NOR2_X1 U19351 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n16305) );
  AOI22_X1 U19352 ( .A1(P3_D_C_N_REG_SCAN_IN), .A2(n18608), .B1(n16305), .B2(
        n18490), .ZN(n16304) );
  OAI21_X1 U19353 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n18608), .A(n16304), 
        .ZN(P3_U2635) );
  OAI21_X1 U19354 ( .B1(n16305), .B2(BS16), .A(n18565), .ZN(n18563) );
  OAI21_X1 U19355 ( .B1(n18565), .B2(n18620), .A(n18563), .ZN(P3_U2636) );
  AND3_X1 U19356 ( .A1(n18424), .A2(n16307), .A3(n16306), .ZN(n18447) );
  NOR2_X1 U19357 ( .A1(n18447), .A2(n18459), .ZN(n18610) );
  OAI21_X1 U19358 ( .B1(n18610), .B2(n16309), .A(n16308), .ZN(P3_U2637) );
  NOR4_X1 U19359 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16313) );
  NOR4_X1 U19360 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16312) );
  NOR4_X1 U19361 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16311) );
  NOR4_X1 U19362 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16310) );
  NAND4_X1 U19363 ( .A1(n16313), .A2(n16312), .A3(n16311), .A4(n16310), .ZN(
        n16319) );
  NOR4_X1 U19364 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16317) );
  AOI211_X1 U19365 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16316) );
  NOR4_X1 U19366 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16315) );
  NOR4_X1 U19367 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16314) );
  NAND4_X1 U19368 ( .A1(n16317), .A2(n16316), .A3(n16315), .A4(n16314), .ZN(
        n16318) );
  NOR2_X1 U19369 ( .A1(n16319), .A2(n16318), .ZN(n18603) );
  INV_X1 U19370 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18558) );
  NOR3_X1 U19371 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16321) );
  OAI21_X1 U19372 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16321), .A(n18603), .ZN(
        n16320) );
  OAI21_X1 U19373 ( .B1(n18603), .B2(n18558), .A(n16320), .ZN(P3_U2638) );
  INV_X1 U19374 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18599) );
  INV_X1 U19375 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18564) );
  AOI21_X1 U19376 ( .B1(n18599), .B2(n18564), .A(n16321), .ZN(n16322) );
  INV_X1 U19377 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18555) );
  INV_X1 U19378 ( .A(n18603), .ZN(n18606) );
  AOI22_X1 U19379 ( .A1(n18603), .A2(n16322), .B1(n18555), .B2(n18606), .ZN(
        P3_U2639) );
  NAND3_X1 U19380 ( .A1(n18566), .A2(n18468), .A3(n18620), .ZN(n18476) );
  NOR2_X1 U19381 ( .A1(n18577), .A2(n18476), .ZN(n16661) );
  NAND2_X1 U19382 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18468), .ZN(n18469) );
  INV_X1 U19383 ( .A(n18469), .ZN(n18339) );
  AND2_X1 U19384 ( .A1(n18471), .A2(n18339), .ZN(n18463) );
  NOR4_X2 U19385 ( .A1(n17951), .A2(n18637), .A3(n16661), .A4(n18463), .ZN(
        n16701) );
  INV_X1 U19386 ( .A(n18622), .ZN(n18617) );
  AOI211_X1 U19387 ( .C1(n18621), .C2(n18619), .A(n18617), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18461) );
  AOI211_X4 U19388 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n17188), .A(n18461), .B(
        n18635), .ZN(n16693) );
  AOI22_X1 U19389 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n16675), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n16693), .ZN(n16349) );
  NAND2_X1 U19390 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n17188), .ZN(n16325) );
  AOI211_X4 U19391 ( .C1(n18620), .C2(n18622), .A(n18635), .B(n16325), .ZN(
        n16686) );
  NOR2_X1 U19392 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16698), .ZN(n16345) );
  NOR2_X1 U19393 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16685) );
  NAND2_X1 U19394 ( .A1(n16685), .A2(n16984), .ZN(n16670) );
  NOR2_X1 U19395 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n16670), .ZN(n16655) );
  NAND2_X1 U19396 ( .A1(n16655), .A2(n16644), .ZN(n16643) );
  NOR2_X1 U19397 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n16643), .ZN(n16627) );
  NAND2_X1 U19398 ( .A1(n16627), .A2(n16971), .ZN(n16618) );
  NOR2_X1 U19399 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n16618), .ZN(n16609) );
  NAND2_X1 U19400 ( .A1(n16609), .A2(n20811), .ZN(n16593) );
  NOR2_X1 U19401 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16593), .ZN(n16573) );
  NAND2_X1 U19402 ( .A1(n16573), .A2(n16576), .ZN(n16572) );
  NOR2_X1 U19403 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n16572), .ZN(n16552) );
  NAND2_X1 U19404 ( .A1(n16552), .A2(n16545), .ZN(n16544) );
  NOR2_X1 U19405 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16544), .ZN(n16528) );
  NAND2_X1 U19406 ( .A1(n16528), .A2(n9821), .ZN(n16520) );
  NOR2_X1 U19407 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n16520), .ZN(n16509) );
  INV_X1 U19408 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n16499) );
  NAND2_X1 U19409 ( .A1(n16509), .A2(n16499), .ZN(n16498) );
  NOR2_X1 U19410 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n16498), .ZN(n16484) );
  INV_X1 U19411 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16479) );
  NAND2_X1 U19412 ( .A1(n16484), .A2(n16479), .ZN(n16476) );
  NOR2_X1 U19413 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n16476), .ZN(n16468) );
  NAND2_X1 U19414 ( .A1(n16468), .A2(n16460), .ZN(n16457) );
  NOR2_X1 U19415 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16457), .ZN(n16442) );
  NAND2_X1 U19416 ( .A1(n16442), .A2(n16437), .ZN(n16436) );
  NOR2_X1 U19417 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16436), .ZN(n16420) );
  NAND2_X1 U19418 ( .A1(n16420), .A2(n16417), .ZN(n16416) );
  NOR2_X1 U19419 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16416), .ZN(n16400) );
  NAND2_X1 U19420 ( .A1(n16400), .A2(n16396), .ZN(n16395) );
  NOR2_X1 U19421 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16395), .ZN(n16383) );
  NAND2_X1 U19422 ( .A1(n16383), .A2(n16376), .ZN(n16375) );
  NOR2_X1 U19423 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16375), .ZN(n16359) );
  INV_X1 U19424 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18548) );
  NAND2_X1 U19425 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16369) );
  OR2_X1 U19426 ( .A1(n18548), .A2(n16369), .ZN(n16330) );
  INV_X1 U19427 ( .A(n18461), .ZN(n16326) );
  INV_X1 U19428 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18537) );
  INV_X1 U19429 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18536) );
  INV_X1 U19430 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18521) );
  INV_X1 U19431 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18517) );
  INV_X1 U19432 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18499) );
  NAND3_X1 U19433 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16656) );
  NOR2_X1 U19434 ( .A1(n18499), .A2(n16656), .ZN(n16628) );
  NAND2_X1 U19435 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16628), .ZN(n16533) );
  NAND3_X1 U19436 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .A3(P3_REIP_REG_7__SCAN_IN), .ZN(n16534) );
  NOR2_X1 U19437 ( .A1(n16533), .A2(n16534), .ZN(n16531) );
  INV_X1 U19438 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18511) );
  NAND2_X1 U19439 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16567) );
  NOR2_X1 U19440 ( .A1(n18511), .A2(n16567), .ZN(n16532) );
  NAND4_X1 U19441 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(P3_REIP_REG_12__SCAN_IN), 
        .A3(n16531), .A4(n16532), .ZN(n16518) );
  NOR2_X1 U19442 ( .A1(n18517), .A2(n16518), .ZN(n16497) );
  NAND2_X1 U19443 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16497), .ZN(n16502) );
  NOR2_X1 U19444 ( .A1(n18521), .A2(n16502), .ZN(n16487) );
  NAND2_X1 U19445 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16487), .ZN(n16461) );
  NAND3_X1 U19446 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .ZN(n16435) );
  NOR2_X1 U19447 ( .A1(n16461), .A2(n16435), .ZN(n16431) );
  NAND3_X1 U19448 ( .A1(n16431), .A2(P3_REIP_REG_22__SCAN_IN), .A3(
        P3_REIP_REG_21__SCAN_IN), .ZN(n16423) );
  OR2_X1 U19449 ( .A1(n18536), .A2(n16423), .ZN(n16413) );
  NOR2_X1 U19450 ( .A1(n18537), .A2(n16413), .ZN(n16329) );
  INV_X1 U19451 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18539) );
  INV_X1 U19452 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18542) );
  NOR3_X1 U19453 ( .A1(n18539), .A2(n18542), .A3(n16701), .ZN(n16328) );
  INV_X1 U19454 ( .A(n16701), .ZN(n16690) );
  NAND2_X1 U19455 ( .A1(n16666), .A2(n16690), .ZN(n16700) );
  INV_X1 U19456 ( .A(n16700), .ZN(n16327) );
  AOI21_X1 U19457 ( .B1(n16329), .B2(n16328), .A(n16327), .ZN(n16394) );
  AOI21_X1 U19458 ( .B1(n16330), .B2(n16687), .A(n16394), .ZN(n16368) );
  NAND2_X1 U19459 ( .A1(n16687), .A2(n16329), .ZN(n16409) );
  NOR2_X1 U19460 ( .A1(n18539), .A2(n16409), .ZN(n16393) );
  NAND2_X1 U19461 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16393), .ZN(n16380) );
  NOR2_X1 U19462 ( .A1(n16380), .A2(n16330), .ZN(n16346) );
  INV_X1 U19463 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n20804) );
  NAND2_X1 U19464 ( .A1(n16346), .A2(n20804), .ZN(n16355) );
  AOI21_X1 U19465 ( .B1(n16368), .B2(n16355), .A(n18551), .ZN(n16344) );
  INV_X1 U19466 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17276) );
  NOR2_X1 U19467 ( .A1(n17276), .A2(n16333), .ZN(n16332) );
  OAI21_X1 U19468 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16332), .A(
        n16331), .ZN(n17263) );
  INV_X1 U19469 ( .A(n17263), .ZN(n16372) );
  AOI21_X1 U19470 ( .B1(n17276), .B2(n16333), .A(n16332), .ZN(n17273) );
  NAND2_X1 U19471 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17283), .ZN(
        n17255) );
  AOI21_X1 U19472 ( .B1(n9873), .B2(n17255), .A(n16334), .ZN(n17291) );
  INV_X1 U19473 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n20756) );
  AND2_X1 U19474 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17323), .ZN(
        n17294) );
  NAND2_X1 U19475 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17294), .ZN(
        n16336) );
  NOR2_X1 U19476 ( .A1(n20756), .A2(n16336), .ZN(n16335) );
  OAI21_X1 U19477 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16335), .A(
        n17255), .ZN(n17299) );
  INV_X1 U19478 ( .A(n17299), .ZN(n16403) );
  AOI21_X1 U19479 ( .B1(n20756), .B2(n16336), .A(n16335), .ZN(n17309) );
  OAI21_X1 U19480 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17294), .A(
        n16336), .ZN(n16337) );
  INV_X1 U19481 ( .A(n16337), .ZN(n17324) );
  INV_X1 U19482 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16339) );
  INV_X1 U19483 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16453) );
  NOR2_X1 U19484 ( .A1(n17620), .A2(n17378), .ZN(n17377) );
  INV_X1 U19485 ( .A(n17377), .ZN(n16465) );
  NOR2_X1 U19486 ( .A1(n17380), .A2(n16465), .ZN(n17333) );
  INV_X1 U19487 ( .A(n17333), .ZN(n16463) );
  NOR2_X1 U19488 ( .A1(n16453), .A2(n16463), .ZN(n16340) );
  NAND2_X1 U19489 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16340), .ZN(
        n16338) );
  AOI21_X1 U19490 ( .B1(n16339), .B2(n16338), .A(n17294), .ZN(n17335) );
  XOR2_X1 U19491 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n16340), .Z(
        n17350) );
  AOI21_X1 U19492 ( .B1(n16453), .B2(n16463), .A(n16340), .ZN(n17370) );
  NOR2_X1 U19493 ( .A1(n17620), .A2(n17526), .ZN(n16590) );
  INV_X1 U19494 ( .A(n16590), .ZN(n16602) );
  NOR2_X1 U19495 ( .A1(n16341), .A2(n16602), .ZN(n16554) );
  NAND2_X1 U19496 ( .A1(n17416), .A2(n16554), .ZN(n16494) );
  INV_X1 U19497 ( .A(n16494), .ZN(n17415) );
  NAND2_X1 U19498 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17415), .ZN(
        n16507) );
  INV_X1 U19499 ( .A(n16507), .ZN(n16495) );
  INV_X1 U19500 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16702) );
  NAND2_X1 U19501 ( .A1(n16495), .A2(n16702), .ZN(n16512) );
  NOR2_X1 U19502 ( .A1(n16450), .A2(n16631), .ZN(n16445) );
  NOR2_X1 U19503 ( .A1(n17350), .A2(n16445), .ZN(n16444) );
  NOR2_X1 U19504 ( .A1(n16444), .A2(n16631), .ZN(n16433) );
  NOR2_X1 U19505 ( .A1(n16432), .A2(n16631), .ZN(n16422) );
  NOR2_X1 U19506 ( .A1(n17324), .A2(n16422), .ZN(n16421) );
  NOR2_X1 U19507 ( .A1(n16421), .A2(n16631), .ZN(n16411) );
  NOR2_X1 U19508 ( .A1(n16410), .A2(n16631), .ZN(n16402) );
  NOR2_X1 U19509 ( .A1(n16403), .A2(n16402), .ZN(n16401) );
  NOR2_X1 U19510 ( .A1(n16401), .A2(n16631), .ZN(n16391) );
  NOR2_X1 U19511 ( .A1(n16390), .A2(n16631), .ZN(n16382) );
  NOR2_X1 U19512 ( .A1(n17273), .A2(n16382), .ZN(n16381) );
  NOR2_X1 U19513 ( .A1(n16381), .A2(n16631), .ZN(n16371) );
  NOR2_X1 U19514 ( .A1(n16370), .A2(n16631), .ZN(n16361) );
  NOR2_X1 U19515 ( .A1(n16360), .A2(n16631), .ZN(n16353) );
  NAND2_X1 U19516 ( .A1(n16342), .A2(n16661), .ZN(n16615) );
  NOR3_X1 U19517 ( .A1(n16354), .A2(n16353), .A3(n16615), .ZN(n16343) );
  AOI211_X1 U19518 ( .C1(n16345), .C2(n16359), .A(n16344), .B(n16343), .ZN(
        n16348) );
  NAND3_X1 U19519 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16346), .A3(n18551), 
        .ZN(n16347) );
  INV_X1 U19520 ( .A(n16368), .ZN(n16350) );
  AOI22_X1 U19521 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16682), .B1(
        P3_REIP_REG_30__SCAN_IN), .B2(n16350), .ZN(n16358) );
  XNOR2_X1 U19522 ( .A(P3_EBX_REG_30__SCAN_IN), .B(n16359), .ZN(n16351) );
  AOI22_X1 U19523 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16693), .B1(n16686), 
        .B2(n16351), .ZN(n16357) );
  INV_X1 U19524 ( .A(n16661), .ZN(n18474) );
  AOI21_X1 U19525 ( .B1(n16354), .B2(n16353), .A(n18474), .ZN(n16352) );
  OAI21_X1 U19526 ( .B1(n16354), .B2(n16353), .A(n16352), .ZN(n16356) );
  NAND4_X1 U19527 ( .A1(n16358), .A2(n16357), .A3(n16356), .A4(n16355), .ZN(
        P3_U2641) );
  AOI22_X1 U19528 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16675), .B1(
        n16693), .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n16367) );
  AOI211_X1 U19529 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16375), .A(n16359), .B(
        n16698), .ZN(n16365) );
  NOR3_X1 U19530 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16380), .A3(n16369), 
        .ZN(n16364) );
  AOI211_X1 U19531 ( .C1(n16362), .C2(n16361), .A(n16360), .B(n18474), .ZN(
        n16363) );
  NOR3_X1 U19532 ( .A1(n16365), .A2(n16364), .A3(n16363), .ZN(n16366) );
  OAI211_X1 U19533 ( .C1(n16368), .C2(n18548), .A(n16367), .B(n16366), .ZN(
        P3_U2642) );
  OAI21_X1 U19534 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(P3_REIP_REG_27__SCAN_IN), 
        .A(n16369), .ZN(n16379) );
  AOI211_X1 U19535 ( .C1(n16372), .C2(n16371), .A(n16370), .B(n18474), .ZN(
        n16374) );
  INV_X1 U19536 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18547) );
  INV_X1 U19537 ( .A(n16394), .ZN(n16389) );
  OAI22_X1 U19538 ( .A1(n18547), .A2(n16389), .B1(n16697), .B2(n16376), .ZN(
        n16373) );
  AOI211_X1 U19539 ( .C1(n16675), .C2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16374), .B(n16373), .ZN(n16378) );
  OAI211_X1 U19540 ( .C1(n16383), .C2(n16376), .A(n16686), .B(n16375), .ZN(
        n16377) );
  OAI211_X1 U19541 ( .C1(n16380), .C2(n16379), .A(n16378), .B(n16377), .ZN(
        P3_U2643) );
  INV_X1 U19542 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18544) );
  AOI22_X1 U19543 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16682), .B1(
        n16693), .B2(P3_EBX_REG_27__SCAN_IN), .ZN(n16388) );
  INV_X1 U19544 ( .A(n16380), .ZN(n16386) );
  AOI211_X1 U19545 ( .C1(n17273), .C2(n16382), .A(n16381), .B(n18474), .ZN(
        n16385) );
  AOI211_X1 U19546 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16395), .A(n16383), .B(
        n16698), .ZN(n16384) );
  AOI211_X1 U19547 ( .C1(n16386), .C2(n18544), .A(n16385), .B(n16384), .ZN(
        n16387) );
  OAI211_X1 U19548 ( .C1(n18544), .C2(n16389), .A(n16388), .B(n16387), .ZN(
        P3_U2644) );
  AOI22_X1 U19549 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16675), .B1(
        n16693), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16399) );
  AOI211_X1 U19550 ( .C1(n17291), .C2(n16391), .A(n16390), .B(n18474), .ZN(
        n16392) );
  AOI221_X1 U19551 ( .B1(P3_REIP_REG_26__SCAN_IN), .B2(n16394), .C1(n16393), 
        .C2(n16394), .A(n16392), .ZN(n16398) );
  OAI211_X1 U19552 ( .C1(n16400), .C2(n16396), .A(n16686), .B(n16395), .ZN(
        n16397) );
  NAND3_X1 U19553 ( .A1(n16399), .A2(n16398), .A3(n16397), .ZN(P3_U2645) );
  AOI22_X1 U19554 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16682), .B1(
        n16693), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n16408) );
  AOI21_X1 U19555 ( .B1(n16687), .B2(n16413), .A(n16701), .ZN(n16430) );
  OAI21_X1 U19556 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n16666), .A(n16430), 
        .ZN(n16406) );
  AOI211_X1 U19557 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n16416), .A(n16400), .B(
        n16698), .ZN(n16405) );
  AOI211_X1 U19558 ( .C1(n16403), .C2(n16402), .A(n16401), .B(n18474), .ZN(
        n16404) );
  AOI211_X1 U19559 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16406), .A(n16405), 
        .B(n16404), .ZN(n16407) );
  OAI211_X1 U19560 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16409), .A(n16408), 
        .B(n16407), .ZN(P3_U2646) );
  AOI211_X1 U19561 ( .C1(n17309), .C2(n16411), .A(n16410), .B(n18474), .ZN(
        n16415) );
  NAND2_X1 U19562 ( .A1(n16687), .A2(n18537), .ZN(n16412) );
  OAI22_X1 U19563 ( .A1(n16697), .A2(n16417), .B1(n16413), .B2(n16412), .ZN(
        n16414) );
  AOI211_X1 U19564 ( .C1(n16675), .C2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16415), .B(n16414), .ZN(n16419) );
  OAI211_X1 U19565 ( .C1(n16420), .C2(n16417), .A(n16686), .B(n16416), .ZN(
        n16418) );
  OAI211_X1 U19566 ( .C1(n16430), .C2(n18537), .A(n16419), .B(n16418), .ZN(
        P3_U2647) );
  AOI211_X1 U19567 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n16436), .A(n16420), .B(
        n16698), .ZN(n16428) );
  AOI211_X1 U19568 ( .C1(n17324), .C2(n16422), .A(n16421), .B(n18474), .ZN(
        n16427) );
  NOR3_X1 U19569 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16666), .A3(n16423), 
        .ZN(n16426) );
  AOI22_X1 U19570 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n16675), .B1(
        n16693), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n16424) );
  INV_X1 U19571 ( .A(n16424), .ZN(n16425) );
  NOR4_X1 U19572 ( .A1(n16428), .A2(n16427), .A3(n16426), .A4(n16425), .ZN(
        n16429) );
  OAI21_X1 U19573 ( .B1(n18536), .B2(n16430), .A(n16429), .ZN(P3_U2648) );
  AOI22_X1 U19574 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16682), .B1(
        n16693), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16441) );
  OAI21_X1 U19575 ( .B1(n16431), .B2(n16666), .A(n16690), .ZN(n16456) );
  AOI211_X1 U19576 ( .C1(n17335), .C2(n16433), .A(n16432), .B(n18474), .ZN(
        n16434) );
  AOI21_X1 U19577 ( .B1(n16456), .B2(P3_REIP_REG_22__SCAN_IN), .A(n16434), 
        .ZN(n16440) );
  INV_X1 U19578 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18533) );
  INV_X1 U19579 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18531) );
  INV_X1 U19580 ( .A(n16461), .ZN(n16485) );
  NAND2_X1 U19581 ( .A1(n16687), .A2(n16485), .ZN(n16473) );
  NOR2_X1 U19582 ( .A1(n16435), .A2(n16473), .ZN(n16447) );
  OAI221_X1 U19583 ( .B1(P3_REIP_REG_22__SCAN_IN), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n18533), .C2(n18531), .A(n16447), .ZN(n16439) );
  OAI211_X1 U19584 ( .C1(n16442), .C2(n16437), .A(n16686), .B(n16436), .ZN(
        n16438) );
  NAND4_X1 U19585 ( .A1(n16441), .A2(n16440), .A3(n16439), .A4(n16438), .ZN(
        P3_U2649) );
  INV_X1 U19586 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17354) );
  AOI211_X1 U19587 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n16457), .A(n16442), .B(
        n16698), .ZN(n16443) );
  AOI21_X1 U19588 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16693), .A(n16443), .ZN(
        n16449) );
  AOI211_X1 U19589 ( .C1(n17350), .C2(n16445), .A(n16444), .B(n18474), .ZN(
        n16446) );
  AOI221_X1 U19590 ( .B1(n16456), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n16447), 
        .C2(n18531), .A(n16446), .ZN(n16448) );
  OAI211_X1 U19591 ( .C1(n17354), .C2(n16621), .A(n16449), .B(n16448), .ZN(
        P3_U2650) );
  AOI211_X1 U19592 ( .C1(n17370), .C2(n16451), .A(n16450), .B(n18474), .ZN(
        n16455) );
  INV_X1 U19593 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18530) );
  NAND3_X1 U19594 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(n18530), .ZN(n16452) );
  OAI22_X1 U19595 ( .A1(n16453), .A2(n16621), .B1(n16473), .B2(n16452), .ZN(
        n16454) );
  AOI211_X1 U19596 ( .C1(n16456), .C2(P3_REIP_REG_20__SCAN_IN), .A(n16455), 
        .B(n16454), .ZN(n16459) );
  OAI211_X1 U19597 ( .C1(n16468), .C2(n16460), .A(n16686), .B(n16457), .ZN(
        n16458) );
  OAI211_X1 U19598 ( .C1(n16460), .C2(n16697), .A(n16459), .B(n16458), .ZN(
        P3_U2651) );
  AOI21_X1 U19599 ( .B1(n16687), .B2(n16461), .A(n16701), .ZN(n16489) );
  INV_X1 U19600 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18527) );
  INV_X1 U19601 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18525) );
  AOI221_X1 U19602 ( .B1(P3_REIP_REG_19__SCAN_IN), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n18527), .C2(n18525), .A(n16473), .ZN(n16462) );
  AOI211_X1 U19603 ( .C1(n16693), .C2(P3_EBX_REG_19__SCAN_IN), .A(n17951), .B(
        n16462), .ZN(n16472) );
  INV_X1 U19604 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17392) );
  NOR2_X1 U19605 ( .A1(n17392), .A2(n16465), .ZN(n16464) );
  OAI21_X1 U19606 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16464), .A(
        n16463), .ZN(n17383) );
  AOI22_X1 U19607 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16465), .B1(
        n17377), .B2(n17392), .ZN(n17389) );
  NAND2_X1 U19608 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16702), .ZN(
        n16563) );
  OAI21_X1 U19609 ( .B1(n17378), .B2(n16563), .A(n16342), .ZN(n16475) );
  NAND2_X1 U19610 ( .A1(n17389), .A2(n16475), .ZN(n16474) );
  NAND2_X1 U19611 ( .A1(n16342), .A2(n16474), .ZN(n16467) );
  OAI21_X1 U19612 ( .B1(n17383), .B2(n16467), .A(n16661), .ZN(n16466) );
  AOI21_X1 U19613 ( .B1(n17383), .B2(n16467), .A(n16466), .ZN(n16470) );
  AOI211_X1 U19614 ( .C1(P3_EBX_REG_19__SCAN_IN), .C2(n16476), .A(n16468), .B(
        n16698), .ZN(n16469) );
  AOI211_X1 U19615 ( .C1(n16675), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16470), .B(n16469), .ZN(n16471) );
  OAI211_X1 U19616 ( .C1(n16489), .C2(n18527), .A(n16472), .B(n16471), .ZN(
        P3_U2652) );
  OAI22_X1 U19617 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16473), .B1(n17392), 
        .B2(n16621), .ZN(n16481) );
  OAI211_X1 U19618 ( .C1(n17389), .C2(n16475), .A(n16661), .B(n16474), .ZN(
        n16478) );
  OAI211_X1 U19619 ( .C1(n16484), .C2(n16479), .A(n16686), .B(n16476), .ZN(
        n16477) );
  OAI211_X1 U19620 ( .C1(n16479), .C2(n16697), .A(n16478), .B(n16477), .ZN(
        n16480) );
  NOR3_X1 U19621 ( .A1(n17951), .A2(n16481), .A3(n16480), .ZN(n16482) );
  OAI21_X1 U19622 ( .B1(n16489), .B2(n18525), .A(n16482), .ZN(P3_U2653) );
  INV_X1 U19623 ( .A(n16563), .ZN(n16678) );
  AOI21_X1 U19624 ( .B1(n17401), .B2(n16678), .A(n16631), .ZN(n16483) );
  AOI221_X1 U19625 ( .B1(n17419), .B2(n9876), .C1(n16494), .C2(n9876), .A(
        n17377), .ZN(n17402) );
  XNOR2_X1 U19626 ( .A(n16483), .B(n17402), .ZN(n16493) );
  AOI211_X1 U19627 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n16498), .A(n16484), .B(
        n16698), .ZN(n16491) );
  INV_X1 U19628 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18524) );
  NOR2_X1 U19629 ( .A1(n16485), .A2(n16666), .ZN(n16486) );
  AOI22_X1 U19630 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16675), .B1(
        n16487), .B2(n16486), .ZN(n16488) );
  OAI211_X1 U19631 ( .C1(n16489), .C2(n18524), .A(n16488), .B(n17861), .ZN(
        n16490) );
  AOI211_X1 U19632 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n16693), .A(n16491), .B(
        n16490), .ZN(n16492) );
  OAI21_X1 U19633 ( .B1(n18474), .B2(n16493), .A(n16492), .ZN(P3_U2654) );
  OAI22_X1 U19634 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16495), .B1(
        n16494), .B2(n17419), .ZN(n17422) );
  XNOR2_X1 U19635 ( .A(n16496), .B(n17422), .ZN(n16506) );
  AOI22_X1 U19636 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16682), .B1(
        n16693), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n16505) );
  OAI21_X1 U19637 ( .B1(n16497), .B2(n16666), .A(n16690), .ZN(n16524) );
  INV_X1 U19638 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18519) );
  AND3_X1 U19639 ( .A1(n18519), .A2(n16687), .A3(n16497), .ZN(n16511) );
  NAND2_X1 U19640 ( .A1(n16687), .A2(n18521), .ZN(n16501) );
  OAI211_X1 U19641 ( .C1(n16509), .C2(n16499), .A(n16686), .B(n16498), .ZN(
        n16500) );
  OAI211_X1 U19642 ( .C1(n16502), .C2(n16501), .A(n17861), .B(n16500), .ZN(
        n16503) );
  AOI221_X1 U19643 ( .B1(n16524), .B2(P3_REIP_REG_16__SCAN_IN), .C1(n16511), 
        .C2(P3_REIP_REG_16__SCAN_IN), .A(n16503), .ZN(n16504) );
  OAI211_X1 U19644 ( .C1(n18474), .C2(n16506), .A(n16505), .B(n16504), .ZN(
        P3_U2655) );
  AOI22_X1 U19645 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n16675), .B1(
        n16693), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n16516) );
  OAI21_X1 U19646 ( .B1(n16631), .B2(n16702), .A(n16661), .ZN(n16696) );
  OAI21_X1 U19647 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17415), .A(
        n16507), .ZN(n17432) );
  AOI211_X1 U19648 ( .C1(n16342), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16696), .B(n17432), .ZN(n16508) );
  NOR2_X1 U19649 ( .A1(n17951), .A2(n16508), .ZN(n16515) );
  AOI211_X1 U19650 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n16520), .A(n16509), .B(
        n16698), .ZN(n16510) );
  AOI211_X1 U19651 ( .C1(n16524), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16511), 
        .B(n16510), .ZN(n16514) );
  INV_X1 U19652 ( .A(n16615), .ZN(n16683) );
  NAND3_X1 U19653 ( .A1(n16683), .A2(n16512), .A3(n17432), .ZN(n16513) );
  NAND4_X1 U19654 ( .A1(n16516), .A2(n16515), .A3(n16514), .A4(n16513), .ZN(
        P3_U2656) );
  INV_X1 U19655 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17474) );
  INV_X1 U19656 ( .A(n16554), .ZN(n17454) );
  NOR2_X1 U19657 ( .A1(n17474), .A2(n17454), .ZN(n16543) );
  NAND2_X1 U19658 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16543), .ZN(
        n16527) );
  OAI21_X1 U19659 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16527), .A(
        n16342), .ZN(n16517) );
  AOI21_X1 U19660 ( .B1(n17443), .B2(n16527), .A(n17415), .ZN(n17445) );
  XOR2_X1 U19661 ( .A(n16517), .B(n17445), .Z(n16526) );
  NOR3_X1 U19662 ( .A1(n16518), .A2(P3_REIP_REG_14__SCAN_IN), .A3(n16666), 
        .ZN(n16519) );
  AOI211_X1 U19663 ( .C1(n16693), .C2(P3_EBX_REG_14__SCAN_IN), .A(n17951), .B(
        n16519), .ZN(n16522) );
  OAI211_X1 U19664 ( .C1(n16528), .C2(n9821), .A(n16686), .B(n16520), .ZN(
        n16521) );
  OAI211_X1 U19665 ( .C1(n16621), .C2(n17443), .A(n16522), .B(n16521), .ZN(
        n16523) );
  AOI21_X1 U19666 ( .B1(P3_REIP_REG_14__SCAN_IN), .B2(n16524), .A(n16523), 
        .ZN(n16525) );
  OAI21_X1 U19667 ( .B1(n16526), .B2(n18474), .A(n16525), .ZN(P3_U2657) );
  OAI21_X1 U19668 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16543), .A(
        n16527), .ZN(n17460) );
  OAI21_X1 U19669 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16527), .A(
        n17460), .ZN(n16541) );
  AOI211_X1 U19670 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n16544), .A(n16528), .B(
        n16698), .ZN(n16529) );
  AOI211_X1 U19671 ( .C1(n16693), .C2(P3_EBX_REG_13__SCAN_IN), .A(n17951), .B(
        n16529), .ZN(n16540) );
  INV_X1 U19672 ( .A(n16543), .ZN(n16530) );
  AOI211_X1 U19673 ( .C1(n16342), .C2(n16530), .A(n16696), .B(n17460), .ZN(
        n16538) );
  NAND2_X1 U19674 ( .A1(n16687), .A2(n16531), .ZN(n16582) );
  NOR2_X1 U19675 ( .A1(n16567), .A2(n16582), .ZN(n16553) );
  NAND2_X1 U19676 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16553), .ZN(n16551) );
  INV_X1 U19677 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18515) );
  XOR2_X1 U19678 ( .A(n18515), .B(P3_REIP_REG_12__SCAN_IN), .Z(n16536) );
  INV_X1 U19679 ( .A(n16532), .ZN(n16535) );
  OR2_X1 U19680 ( .A1(n16701), .A2(n16533), .ZN(n16600) );
  OAI21_X1 U19681 ( .B1(n16534), .B2(n16600), .A(n16700), .ZN(n16588) );
  INV_X1 U19682 ( .A(n16588), .ZN(n16598) );
  AOI21_X1 U19683 ( .B1(n16535), .B2(n16700), .A(n16598), .ZN(n16558) );
  OAI22_X1 U19684 ( .A1(n16551), .A2(n16536), .B1(n16558), .B2(n18515), .ZN(
        n16537) );
  AOI211_X1 U19685 ( .C1(n16675), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16538), .B(n16537), .ZN(n16539) );
  OAI211_X1 U19686 ( .C1(n16615), .C2(n16541), .A(n16540), .B(n16539), .ZN(
        P3_U2658) );
  INV_X1 U19687 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18513) );
  AOI21_X1 U19688 ( .B1(n17474), .B2(n17454), .A(n16543), .ZN(n17481) );
  OAI21_X1 U19689 ( .B1(n17474), .B2(n16631), .A(n17481), .ZN(n16542) );
  OAI22_X1 U19690 ( .A1(n16696), .A2(n16542), .B1(n17474), .B2(n16621), .ZN(
        n16549) );
  AOI22_X1 U19691 ( .A1(n16543), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n17474), .B2(n17454), .ZN(n16547) );
  OAI211_X1 U19692 ( .C1(n16552), .C2(n16545), .A(n16686), .B(n16544), .ZN(
        n16546) );
  OAI211_X1 U19693 ( .C1(n16547), .C2(n16615), .A(n17861), .B(n16546), .ZN(
        n16548) );
  AOI211_X1 U19694 ( .C1(n16693), .C2(P3_EBX_REG_12__SCAN_IN), .A(n16549), .B(
        n16548), .ZN(n16550) );
  OAI221_X1 U19695 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n16551), .C1(n18513), 
        .C2(n16558), .A(n16550), .ZN(P3_U2659) );
  AOI211_X1 U19696 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n16572), .A(n16552), .B(
        n16698), .ZN(n16560) );
  NOR2_X1 U19697 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16553), .ZN(n16557) );
  INV_X1 U19698 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17485) );
  NAND2_X1 U19699 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16564) );
  NOR2_X1 U19700 ( .A1(n16564), .A2(n16602), .ZN(n16577) );
  NAND2_X1 U19701 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16577), .ZN(
        n16565) );
  AOI21_X1 U19702 ( .B1(n17485), .B2(n16565), .A(n16554), .ZN(n17488) );
  OAI21_X1 U19703 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16565), .A(
        n16342), .ZN(n16555) );
  XOR2_X1 U19704 ( .A(n17488), .B(n16555), .Z(n16556) );
  OAI22_X1 U19705 ( .A1(n16558), .A2(n16557), .B1(n18474), .B2(n16556), .ZN(
        n16559) );
  AOI211_X1 U19706 ( .C1(n16675), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16560), .B(n16559), .ZN(n16561) );
  OAI211_X1 U19707 ( .C1(n16697), .C2(n16562), .A(n16561), .B(n17861), .ZN(
        P3_U2660) );
  NOR2_X1 U19708 ( .A1(n16601), .A2(n16563), .ZN(n16616) );
  AOI21_X1 U19709 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16616), .A(
        n16631), .ZN(n16591) );
  AOI21_X1 U19710 ( .B1(n16342), .B2(n16564), .A(n16591), .ZN(n16581) );
  OAI21_X1 U19711 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16577), .A(
        n16565), .ZN(n17500) );
  OAI21_X1 U19712 ( .B1(n16581), .B2(n17500), .A(n16661), .ZN(n16566) );
  AOI21_X1 U19713 ( .B1(n16581), .B2(n17500), .A(n16566), .ZN(n16571) );
  INV_X1 U19714 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17498) );
  INV_X1 U19715 ( .A(n16582), .ZN(n16568) );
  OAI211_X1 U19716 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n16568), .B(n16567), .ZN(n16569) );
  OAI211_X1 U19717 ( .C1(n17498), .C2(n16621), .A(n17861), .B(n16569), .ZN(
        n16570) );
  AOI211_X1 U19718 ( .C1(n16598), .C2(P3_REIP_REG_10__SCAN_IN), .A(n16571), 
        .B(n16570), .ZN(n16575) );
  OAI211_X1 U19719 ( .C1(n16573), .C2(n16576), .A(n16686), .B(n16572), .ZN(
        n16574) );
  OAI211_X1 U19720 ( .C1(n16576), .C2(n16697), .A(n16575), .B(n16574), .ZN(
        P3_U2661) );
  INV_X1 U19721 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18508) );
  INV_X1 U19722 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17510) );
  NAND2_X1 U19723 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16590), .ZN(
        n16589) );
  AOI21_X1 U19724 ( .B1(n17510), .B2(n16589), .A(n16577), .ZN(n17514) );
  NOR2_X1 U19725 ( .A1(n16342), .A2(n18474), .ZN(n16603) );
  NAND2_X1 U19726 ( .A1(n16686), .A2(n16593), .ZN(n16579) );
  NAND3_X1 U19727 ( .A1(n16661), .A2(n17510), .A3(n16702), .ZN(n16578) );
  OAI22_X1 U19728 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16579), .B1(n16578), .B2(
        n16589), .ZN(n16580) );
  AOI211_X1 U19729 ( .C1(n17514), .C2(n16603), .A(n17951), .B(n16580), .ZN(
        n16587) );
  OAI21_X1 U19730 ( .B1(n16698), .B2(n16593), .A(n16697), .ZN(n16585) );
  NOR3_X1 U19731 ( .A1(n17514), .A2(n16581), .A3(n18474), .ZN(n16584) );
  OAI22_X1 U19732 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16582), .B1(n17510), 
        .B2(n16621), .ZN(n16583) );
  AOI211_X1 U19733 ( .C1(n16585), .C2(P3_EBX_REG_9__SCAN_IN), .A(n16584), .B(
        n16583), .ZN(n16586) );
  OAI211_X1 U19734 ( .C1(n18508), .C2(n16588), .A(n16587), .B(n16586), .ZN(
        P3_U2662) );
  INV_X1 U19735 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17525) );
  NAND2_X1 U19736 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .ZN(n16607) );
  NAND3_X1 U19737 ( .A1(n16687), .A2(P3_REIP_REG_5__SCAN_IN), .A3(n16628), 
        .ZN(n16626) );
  INV_X1 U19738 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18507) );
  OAI21_X1 U19739 ( .B1(n16607), .B2(n16626), .A(n18507), .ZN(n16597) );
  OAI21_X1 U19740 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16590), .A(
        n16589), .ZN(n17527) );
  INV_X1 U19741 ( .A(n17527), .ZN(n16592) );
  INV_X1 U19742 ( .A(n16591), .ZN(n16605) );
  OAI221_X1 U19743 ( .B1(n16592), .B2(n16591), .C1(n17527), .C2(n16605), .A(
        n16661), .ZN(n16595) );
  OAI211_X1 U19744 ( .C1(n16609), .C2(n20811), .A(n16686), .B(n16593), .ZN(
        n16594) );
  OAI211_X1 U19745 ( .C1(n20811), .C2(n16697), .A(n16595), .B(n16594), .ZN(
        n16596) );
  AOI21_X1 U19746 ( .B1(n16598), .B2(n16597), .A(n16596), .ZN(n16599) );
  OAI211_X1 U19747 ( .C1(n17525), .C2(n16621), .A(n16599), .B(n17861), .ZN(
        P3_U2663) );
  INV_X1 U19748 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18504) );
  NAND2_X1 U19749 ( .A1(n16700), .A2(n16600), .ZN(n16633) );
  NOR2_X1 U19750 ( .A1(n17620), .A2(n16601), .ZN(n16614) );
  OAI21_X1 U19751 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16614), .A(
        n16602), .ZN(n17548) );
  INV_X1 U19752 ( .A(n16603), .ZN(n16681) );
  OAI21_X1 U19753 ( .B1(n16616), .B2(n17548), .A(n16661), .ZN(n16604) );
  AOI22_X1 U19754 ( .A1(n17548), .A2(n16605), .B1(n16681), .B2(n16604), .ZN(
        n16606) );
  AOI211_X1 U19755 ( .C1(n16693), .C2(P3_EBX_REG_7__SCAN_IN), .A(n17951), .B(
        n16606), .ZN(n16613) );
  INV_X1 U19756 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20788) );
  INV_X1 U19757 ( .A(n16607), .ZN(n16608) );
  AOI211_X1 U19758 ( .C1(n20788), .C2(n18504), .A(n16608), .B(n16626), .ZN(
        n16611) );
  AOI211_X1 U19759 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n16618), .A(n16609), .B(
        n16698), .ZN(n16610) );
  AOI211_X1 U19760 ( .C1(n16675), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n16611), .B(n16610), .ZN(n16612) );
  OAI211_X1 U19761 ( .C1(n18504), .C2(n16633), .A(n16613), .B(n16612), .ZN(
        P3_U2664) );
  INV_X1 U19762 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20794) );
  NAND2_X1 U19763 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17552), .ZN(
        n16617) );
  AOI21_X1 U19764 ( .B1(n20794), .B2(n16617), .A(n16614), .ZN(n17558) );
  NOR3_X1 U19765 ( .A1(n17558), .A2(n16616), .A3(n16615), .ZN(n16624) );
  INV_X1 U19766 ( .A(n16617), .ZN(n16629) );
  OAI21_X1 U19767 ( .B1(n16629), .B2(n16631), .A(n17558), .ZN(n16620) );
  OAI211_X1 U19768 ( .C1(n16627), .C2(n16971), .A(n16686), .B(n16618), .ZN(
        n16619) );
  OAI21_X1 U19769 ( .B1(n16696), .B2(n16620), .A(n16619), .ZN(n16623) );
  OAI22_X1 U19770 ( .A1(n20794), .A2(n16621), .B1(n16697), .B2(n16971), .ZN(
        n16622) );
  NOR4_X1 U19771 ( .A1(n17951), .A2(n16624), .A3(n16623), .A4(n16622), .ZN(
        n16625) );
  OAI221_X1 U19772 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16626), .C1(n20788), 
        .C2(n16633), .A(n16625), .ZN(P3_U2665) );
  INV_X1 U19773 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16638) );
  AOI211_X1 U19774 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n16643), .A(n16627), .B(
        n16698), .ZN(n16636) );
  AOI21_X1 U19775 ( .B1(n16687), .B2(n16628), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n16634) );
  INV_X1 U19776 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16630) );
  NAND2_X1 U19777 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17561), .ZN(
        n16639) );
  AOI21_X1 U19778 ( .B1(n16630), .B2(n16639), .A(n16629), .ZN(n17569) );
  AOI21_X1 U19779 ( .B1(n17561), .B2(n16678), .A(n16631), .ZN(n16640) );
  XNOR2_X1 U19780 ( .A(n17569), .B(n16640), .ZN(n16632) );
  OAI22_X1 U19781 ( .A1(n16634), .A2(n16633), .B1(n18474), .B2(n16632), .ZN(
        n16635) );
  AOI211_X1 U19782 ( .C1(n16675), .C2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n16636), .B(n16635), .ZN(n16637) );
  OAI211_X1 U19783 ( .C1(n16697), .C2(n16638), .A(n16637), .B(n17861), .ZN(
        P3_U2666) );
  AOI21_X1 U19784 ( .B1(n16687), .B2(n16656), .A(n16701), .ZN(n16665) );
  AOI22_X1 U19785 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16682), .B1(
        n16693), .B2(P3_EBX_REG_4__SCAN_IN), .ZN(n16651) );
  NOR2_X1 U19786 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17584), .ZN(
        n17579) );
  NOR2_X1 U19787 ( .A1(n17620), .A2(n17584), .ZN(n16652) );
  OAI21_X1 U19788 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16652), .A(
        n16639), .ZN(n17587) );
  AOI22_X1 U19789 ( .A1(n16678), .A2(n17579), .B1(n16640), .B2(n17587), .ZN(
        n16641) );
  AOI221_X1 U19790 ( .B1(n16342), .B2(n16641), .C1(n17587), .C2(n16641), .A(
        n18474), .ZN(n16649) );
  NOR3_X1 U19791 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16666), .A3(n16656), .ZN(
        n16648) );
  NAND2_X1 U19792 ( .A1(n16642), .A2(n18637), .ZN(n16705) );
  OAI211_X1 U19793 ( .C1(n16655), .C2(n16644), .A(n16686), .B(n16643), .ZN(
        n16645) );
  OAI221_X1 U19794 ( .B1(n16705), .B2(n16646), .C1(n16705), .C2(n18451), .A(
        n16645), .ZN(n16647) );
  NOR4_X1 U19795 ( .A1(n17951), .A2(n16649), .A3(n16648), .A4(n16647), .ZN(
        n16650) );
  OAI211_X1 U19796 ( .C1(n16665), .C2(n18499), .A(n16651), .B(n16650), .ZN(
        P3_U2667) );
  INV_X1 U19797 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18497) );
  AOI22_X1 U19798 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n16675), .B1(
        n16693), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n16664) );
  INV_X1 U19799 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16653) );
  NAND2_X1 U19800 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16676) );
  AOI21_X1 U19801 ( .B1(n16653), .B2(n16676), .A(n16652), .ZN(n17597) );
  OAI21_X1 U19802 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16676), .A(
        n16342), .ZN(n16654) );
  XNOR2_X1 U19803 ( .A(n17597), .B(n16654), .ZN(n16662) );
  AOI211_X1 U19804 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n16670), .A(n16655), .B(
        n16698), .ZN(n16660) );
  INV_X1 U19805 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18495) );
  NOR2_X1 U19806 ( .A1(n18599), .A2(n18495), .ZN(n16667) );
  AND2_X1 U19807 ( .A1(n16687), .A2(n16656), .ZN(n16657) );
  INV_X1 U19808 ( .A(n16705), .ZN(n16669) );
  NOR2_X1 U19809 ( .A1(n13689), .A2(n18432), .ZN(n16668) );
  INV_X1 U19810 ( .A(n16668), .ZN(n18431) );
  AOI21_X1 U19811 ( .B1(n18574), .B2(n18431), .A(n16927), .ZN(n18571) );
  AOI22_X1 U19812 ( .A1(n16667), .A2(n16657), .B1(n16669), .B2(n18571), .ZN(
        n16658) );
  INV_X1 U19813 ( .A(n16658), .ZN(n16659) );
  AOI211_X1 U19814 ( .C1(n16662), .C2(n16661), .A(n16660), .B(n16659), .ZN(
        n16663) );
  OAI211_X1 U19815 ( .C1(n16665), .C2(n18497), .A(n16664), .B(n16663), .ZN(
        P3_U2668) );
  OAI21_X1 U19816 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16676), .ZN(n17607) );
  AOI211_X1 U19817 ( .C1(n18599), .C2(n18495), .A(n16667), .B(n16666), .ZN(
        n16674) );
  AOI21_X1 U19818 ( .B1(n18583), .B2(n18434), .A(n16668), .ZN(n18580) );
  AOI22_X1 U19819 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n16701), .B1(n18580), 
        .B2(n16669), .ZN(n16672) );
  OAI211_X1 U19820 ( .C1(n16685), .C2(n16984), .A(n16686), .B(n16670), .ZN(
        n16671) );
  OAI211_X1 U19821 ( .C1(n16984), .C2(n16697), .A(n16672), .B(n16671), .ZN(
        n16673) );
  AOI211_X1 U19822 ( .C1(n16675), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n16674), .B(n16673), .ZN(n16680) );
  OR2_X1 U19823 ( .A1(n16676), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16677) );
  OAI211_X1 U19824 ( .C1(n16678), .C2(n17607), .A(n16683), .B(n16677), .ZN(
        n16679) );
  OAI211_X1 U19825 ( .C1(n17607), .C2(n16681), .A(n16680), .B(n16679), .ZN(
        P3_U2669) );
  AOI21_X1 U19826 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16683), .A(
        n16682), .ZN(n16695) );
  NAND2_X1 U19827 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16975) );
  INV_X1 U19828 ( .A(n16975), .ZN(n16684) );
  NOR2_X1 U19829 ( .A1(n16685), .A2(n16684), .ZN(n16989) );
  AOI22_X1 U19830 ( .A1(n18599), .A2(n16687), .B1(n16686), .B2(n16989), .ZN(
        n16688) );
  INV_X1 U19831 ( .A(n16688), .ZN(n16692) );
  NAND2_X1 U19832 ( .A1(n18434), .A2(n16689), .ZN(n18407) );
  OAI22_X1 U19833 ( .A1(n18599), .A2(n16690), .B1(n18407), .B2(n16705), .ZN(
        n16691) );
  AOI211_X1 U19834 ( .C1(n16693), .C2(P3_EBX_REG_1__SCAN_IN), .A(n16692), .B(
        n16691), .ZN(n16694) );
  OAI221_X1 U19835 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16696), .C1(
        n17620), .C2(n16695), .A(n16694), .ZN(P3_U2670) );
  NAND2_X1 U19836 ( .A1(n16698), .A2(n16697), .ZN(n16699) );
  AOI22_X1 U19837 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16700), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n16699), .ZN(n16704) );
  OR3_X1 U19838 ( .A1(n16702), .A2(n18594), .A3(n16701), .ZN(n16703) );
  OAI211_X1 U19839 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n16705), .A(
        n16704), .B(n16703), .ZN(P3_U2671) );
  AOI22_X1 U19840 ( .A1(n9628), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9613), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16709) );
  AOI22_X1 U19841 ( .A1(n16896), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16708) );
  AOI22_X1 U19842 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16946), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16707) );
  AOI22_X1 U19843 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16706) );
  NAND4_X1 U19844 ( .A1(n16709), .A2(n16708), .A3(n16707), .A4(n16706), .ZN(
        n16715) );
  AOI22_X1 U19845 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16713) );
  AOI22_X1 U19846 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16712) );
  AOI22_X1 U19847 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16711) );
  AOI22_X1 U19848 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16710) );
  NAND4_X1 U19849 ( .A1(n16713), .A2(n16712), .A3(n16711), .A4(n16710), .ZN(
        n16714) );
  NOR2_X1 U19850 ( .A1(n16715), .A2(n16714), .ZN(n16727) );
  AOI22_X1 U19851 ( .A1(n13753), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16719) );
  AOI22_X1 U19852 ( .A1(n9613), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16895), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16718) );
  AOI22_X1 U19853 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16717) );
  AOI22_X1 U19854 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16946), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16716) );
  NAND4_X1 U19855 ( .A1(n16719), .A2(n16718), .A3(n16717), .A4(n16716), .ZN(
        n16725) );
  AOI22_X1 U19856 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16723) );
  AOI22_X1 U19857 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16722) );
  AOI22_X1 U19858 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16721) );
  AOI22_X1 U19859 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16720) );
  NAND4_X1 U19860 ( .A1(n16723), .A2(n16722), .A3(n16721), .A4(n16720), .ZN(
        n16724) );
  NOR2_X1 U19861 ( .A1(n16725), .A2(n16724), .ZN(n16733) );
  NOR3_X1 U19862 ( .A1(n16733), .A2(n16739), .A3(n16732), .ZN(n16726) );
  XOR2_X1 U19863 ( .A(n16727), .B(n16726), .Z(n17003) );
  NOR2_X1 U19864 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16728), .ZN(n16730) );
  OAI22_X1 U19865 ( .A1(n17003), .A2(n16986), .B1(n16730), .B2(n16729), .ZN(
        P3_U2673) );
  NAND2_X1 U19866 ( .A1(n16784), .A2(n16731), .ZN(n16738) );
  INV_X1 U19867 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16737) );
  NOR2_X1 U19868 ( .A1(n16739), .A2(n16732), .ZN(n16734) );
  XNOR2_X1 U19869 ( .A(n16734), .B(n16733), .ZN(n17007) );
  NAND2_X1 U19870 ( .A1(n16992), .A2(n17007), .ZN(n16735) );
  OAI221_X1 U19871 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16738), .C1(n16737), 
        .C2(n16736), .A(n16735), .ZN(P3_U2674) );
  OAI21_X1 U19872 ( .B1(n16741), .B2(n16740), .A(n16739), .ZN(n17018) );
  INV_X1 U19873 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16742) );
  AOI22_X1 U19874 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16743), .B1(n16748), 
        .B2(n16742), .ZN(n16744) );
  OAI21_X1 U19875 ( .B1(n16986), .B2(n17018), .A(n16744), .ZN(P3_U2676) );
  INV_X1 U19876 ( .A(n16745), .ZN(n16753) );
  AOI21_X1 U19877 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n16986), .A(n16753), .ZN(
        n16747) );
  XNOR2_X1 U19878 ( .A(n16746), .B(n16749), .ZN(n17023) );
  OAI22_X1 U19879 ( .A1(n16748), .A2(n16747), .B1(n16986), .B2(n17023), .ZN(
        P3_U2677) );
  AOI21_X1 U19880 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16986), .A(n9694), .ZN(
        n16752) );
  OAI21_X1 U19881 ( .B1(n16751), .B2(n16750), .A(n16749), .ZN(n17028) );
  OAI22_X1 U19882 ( .A1(n16753), .A2(n16752), .B1(n16986), .B2(n17028), .ZN(
        P3_U2678) );
  AOI21_X1 U19883 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16986), .A(n9695), .ZN(
        n16755) );
  XNOR2_X1 U19884 ( .A(n16754), .B(n16757), .ZN(n17033) );
  OAI22_X1 U19885 ( .A1(n9694), .A2(n16755), .B1(n16986), .B2(n17033), .ZN(
        P3_U2679) );
  AOI21_X1 U19886 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n16986), .A(n16756), .ZN(
        n16760) );
  OAI21_X1 U19887 ( .B1(n16759), .B2(n16758), .A(n16757), .ZN(n17038) );
  OAI22_X1 U19888 ( .A1(n9695), .A2(n16760), .B1(n16986), .B2(n17038), .ZN(
        P3_U2680) );
  AOI22_X1 U19889 ( .A1(n16896), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16764) );
  AOI22_X1 U19890 ( .A1(n9614), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16763) );
  AOI22_X1 U19891 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16762) );
  AOI22_X1 U19892 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16761) );
  NAND4_X1 U19893 ( .A1(n16764), .A2(n16763), .A3(n16762), .A4(n16761), .ZN(
        n16770) );
  AOI22_X1 U19894 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16768) );
  AOI22_X1 U19895 ( .A1(n16936), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16767) );
  AOI22_X1 U19896 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16895), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16766) );
  AOI22_X1 U19897 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16765) );
  NAND4_X1 U19898 ( .A1(n16768), .A2(n16767), .A3(n16766), .A4(n16765), .ZN(
        n16769) );
  NOR2_X1 U19899 ( .A1(n16770), .A2(n16769), .ZN(n17041) );
  NAND3_X1 U19900 ( .A1(n16772), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n16986), 
        .ZN(n16771) );
  OAI221_X1 U19901 ( .B1(n16772), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n16986), 
        .C2(n17041), .A(n16771), .ZN(P3_U2681) );
  AOI22_X1 U19902 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16776) );
  AOI22_X1 U19903 ( .A1(n16936), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16775) );
  AOI22_X1 U19904 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(n9628), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16774) );
  AOI22_X1 U19905 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9613), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16773) );
  NAND4_X1 U19906 ( .A1(n16776), .A2(n16775), .A3(n16774), .A4(n16773), .ZN(
        n16782) );
  AOI22_X1 U19907 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16780) );
  AOI22_X1 U19908 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16779) );
  AOI22_X1 U19909 ( .A1(n16896), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16778) );
  AOI22_X1 U19910 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9619), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16777) );
  NAND4_X1 U19911 ( .A1(n16780), .A2(n16779), .A3(n16778), .A4(n16777), .ZN(
        n16781) );
  NOR2_X1 U19912 ( .A1(n16782), .A2(n16781), .ZN(n17048) );
  AOI21_X1 U19913 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16809), .A(n16992), .ZN(
        n16796) );
  AOI22_X1 U19914 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16796), .B1(n16784), 
        .B2(n16783), .ZN(n16785) );
  OAI21_X1 U19915 ( .B1(n17048), .B2(n16986), .A(n16785), .ZN(P3_U2682) );
  AOI22_X1 U19916 ( .A1(n15048), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16789) );
  AOI22_X1 U19917 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13732), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16788) );
  AOI22_X1 U19918 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13772), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16787) );
  AOI22_X1 U19919 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16895), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16786) );
  NAND4_X1 U19920 ( .A1(n16789), .A2(n16788), .A3(n16787), .A4(n16786), .ZN(
        n16795) );
  AOI22_X1 U19921 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16793) );
  AOI22_X1 U19922 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16792) );
  AOI22_X1 U19923 ( .A1(n16896), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16791) );
  AOI22_X1 U19924 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9619), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16790) );
  NAND4_X1 U19925 ( .A1(n16793), .A2(n16792), .A3(n16791), .A4(n16790), .ZN(
        n16794) );
  NOR2_X1 U19926 ( .A1(n16795), .A2(n16794), .ZN(n17055) );
  OAI21_X1 U19927 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n9713), .A(n16796), .ZN(
        n16797) );
  OAI21_X1 U19928 ( .B1(n17055), .B2(n16986), .A(n16797), .ZN(P3_U2683) );
  OAI21_X1 U19929 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n16820), .A(n16986), .ZN(
        n16808) );
  AOI22_X1 U19930 ( .A1(n15048), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16895), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16801) );
  AOI22_X1 U19931 ( .A1(n16936), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13732), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16800) );
  AOI22_X1 U19932 ( .A1(n9613), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16799) );
  AOI22_X1 U19933 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16798) );
  NAND4_X1 U19934 ( .A1(n16801), .A2(n16800), .A3(n16799), .A4(n16798), .ZN(
        n16807) );
  AOI22_X1 U19935 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16805) );
  AOI22_X1 U19936 ( .A1(n16896), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16804) );
  AOI22_X1 U19937 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16803) );
  AOI22_X1 U19938 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16802) );
  NAND4_X1 U19939 ( .A1(n16805), .A2(n16804), .A3(n16803), .A4(n16802), .ZN(
        n16806) );
  NOR2_X1 U19940 ( .A1(n16807), .A2(n16806), .ZN(n17060) );
  OAI22_X1 U19941 ( .A1(n16809), .A2(n16808), .B1(n17060), .B2(n16986), .ZN(
        P3_U2684) );
  AOI22_X1 U19942 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16813) );
  AOI22_X1 U19943 ( .A1(n9628), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9614), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16812) );
  AOI22_X1 U19944 ( .A1(n15048), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16811) );
  AOI22_X1 U19945 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16946), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16810) );
  NAND4_X1 U19946 ( .A1(n16813), .A2(n16812), .A3(n16811), .A4(n16810), .ZN(
        n16819) );
  AOI22_X1 U19947 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16817) );
  AOI22_X1 U19948 ( .A1(n16936), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16816) );
  AOI22_X1 U19949 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16815) );
  AOI22_X1 U19950 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16814) );
  NAND4_X1 U19951 ( .A1(n16817), .A2(n16816), .A3(n16815), .A4(n16814), .ZN(
        n16818) );
  NOR2_X1 U19952 ( .A1(n16819), .A2(n16818), .ZN(n17064) );
  INV_X1 U19953 ( .A(n16820), .ZN(n16821) );
  OAI21_X1 U19954 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n16835), .A(n16821), .ZN(
        n16822) );
  AOI22_X1 U19955 ( .A1(n16992), .A2(n17064), .B1(n16822), .B2(n16986), .ZN(
        P3_U2685) );
  OAI21_X1 U19956 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n16823), .A(n16986), .ZN(
        n16834) );
  AOI22_X1 U19957 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n16928), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n9615), .ZN(n16827) );
  AOI22_X1 U19958 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n16909), .B1(
        n16895), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16826) );
  AOI22_X1 U19959 ( .A1(n9614), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16825) );
  AOI22_X1 U19960 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16824) );
  NAND4_X1 U19961 ( .A1(n16827), .A2(n16826), .A3(n16825), .A4(n16824), .ZN(
        n16833) );
  AOI22_X1 U19962 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n16831) );
  AOI22_X1 U19963 ( .A1(n16936), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15048), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16830) );
  AOI22_X1 U19964 ( .A1(n9628), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n16829) );
  AOI22_X1 U19965 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n16937), .B1(
        n9619), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n16828) );
  NAND4_X1 U19966 ( .A1(n16831), .A2(n16830), .A3(n16829), .A4(n16828), .ZN(
        n16832) );
  NOR2_X1 U19967 ( .A1(n16833), .A2(n16832), .ZN(n17070) );
  OAI22_X1 U19968 ( .A1(n16835), .A2(n16834), .B1(n17070), .B2(n16986), .ZN(
        P3_U2686) );
  AOI22_X1 U19969 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9615), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16839) );
  AOI22_X1 U19970 ( .A1(n13732), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n16838) );
  AOI22_X1 U19971 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16837) );
  AOI22_X1 U19972 ( .A1(n9614), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16836) );
  NAND4_X1 U19973 ( .A1(n16839), .A2(n16838), .A3(n16837), .A4(n16836), .ZN(
        n16845) );
  AOI22_X1 U19974 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16843) );
  AOI22_X1 U19975 ( .A1(n16936), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16842) );
  AOI22_X1 U19976 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16841) );
  AOI22_X1 U19977 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16840) );
  NAND4_X1 U19978 ( .A1(n16843), .A2(n16842), .A3(n16841), .A4(n16840), .ZN(
        n16844) );
  NOR2_X1 U19979 ( .A1(n16845), .A2(n16844), .ZN(n17076) );
  OAI22_X1 U19980 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17108), .B1(n16992), 
        .B2(n16858), .ZN(n16846) );
  OAI21_X1 U19981 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n16858), .A(n16846), .ZN(
        n16847) );
  OAI21_X1 U19982 ( .B1(n17076), .B2(n16986), .A(n16847), .ZN(P3_U2687) );
  AOI22_X1 U19983 ( .A1(n15048), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16851) );
  AOI22_X1 U19984 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16850) );
  AOI22_X1 U19985 ( .A1(n16936), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16849) );
  AOI22_X1 U19986 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15225), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16848) );
  NAND4_X1 U19987 ( .A1(n16851), .A2(n16850), .A3(n16849), .A4(n16848), .ZN(
        n16857) );
  AOI22_X1 U19988 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16855) );
  AOI22_X1 U19989 ( .A1(n9613), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16854) );
  AOI22_X1 U19990 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16853) );
  AOI22_X1 U19991 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9619), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16852) );
  NAND4_X1 U19992 ( .A1(n16855), .A2(n16854), .A3(n16853), .A4(n16852), .ZN(
        n16856) );
  NOR2_X1 U19993 ( .A1(n16857), .A2(n16856), .ZN(n17080) );
  NOR2_X1 U19994 ( .A1(n16992), .A2(n16858), .ZN(n16859) );
  OAI21_X1 U19995 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n16860), .A(n16859), .ZN(
        n16861) );
  OAI21_X1 U19996 ( .B1(n17080), .B2(n16986), .A(n16861), .ZN(P3_U2688) );
  NAND2_X1 U19997 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16862), .ZN(n16877) );
  AOI22_X1 U19998 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16873) );
  INV_X1 U19999 ( .A(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16865) );
  AOI22_X1 U20000 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16864) );
  AOI22_X1 U20001 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16863) );
  OAI211_X1 U20002 ( .C1(n15236), .C2(n16865), .A(n16864), .B(n16863), .ZN(
        n16871) );
  AOI22_X1 U20003 ( .A1(n9614), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16895), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16869) );
  AOI22_X1 U20004 ( .A1(n16946), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16868) );
  AOI22_X1 U20005 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16867) );
  AOI22_X1 U20006 ( .A1(n16936), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16866) );
  NAND4_X1 U20007 ( .A1(n16869), .A2(n16868), .A3(n16867), .A4(n16866), .ZN(
        n16870) );
  AOI211_X1 U20008 ( .C1(n16937), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n16871), .B(n16870), .ZN(n16872) );
  NAND2_X1 U20009 ( .A1(n16873), .A2(n16872), .ZN(n17082) );
  OAI21_X1 U20010 ( .B1(n9821), .B2(n16874), .A(n16986), .ZN(n16875) );
  OAI21_X1 U20011 ( .B1(n16986), .B2(n17082), .A(n16875), .ZN(n16876) );
  OAI21_X1 U20012 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n16877), .A(n16876), .ZN(
        P3_U2689) );
  NOR2_X1 U20013 ( .A1(n16992), .A2(n16878), .ZN(n16905) );
  AOI22_X1 U20014 ( .A1(n13732), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16882) );
  AOI22_X1 U20015 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16881) );
  AOI22_X1 U20016 ( .A1(n16936), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16880) );
  AOI22_X1 U20017 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9628), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16879) );
  NAND4_X1 U20018 ( .A1(n16882), .A2(n16881), .A3(n16880), .A4(n16879), .ZN(
        n16888) );
  AOI22_X1 U20019 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16886) );
  AOI22_X1 U20020 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16885) );
  AOI22_X1 U20021 ( .A1(n9614), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16895), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16884) );
  AOI22_X1 U20022 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16883) );
  NAND4_X1 U20023 ( .A1(n16886), .A2(n16885), .A3(n16884), .A4(n16883), .ZN(
        n16887) );
  NOR2_X1 U20024 ( .A1(n16888), .A2(n16887), .ZN(n17092) );
  INV_X1 U20025 ( .A(n17092), .ZN(n16889) );
  AOI22_X1 U20026 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16905), .B1(n16992), 
        .B2(n16889), .ZN(n16890) );
  OAI21_X1 U20027 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n16891), .A(n16890), .ZN(
        P3_U2691) );
  AOI22_X1 U20028 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16904) );
  INV_X1 U20029 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16894) );
  AOI22_X1 U20030 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16893) );
  AOI22_X1 U20031 ( .A1(n16936), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16892) );
  OAI211_X1 U20032 ( .C1(n15236), .C2(n16894), .A(n16893), .B(n16892), .ZN(
        n16902) );
  AOI22_X1 U20033 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16900) );
  AOI22_X1 U20034 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n9628), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16899) );
  AOI22_X1 U20035 ( .A1(n16909), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16898) );
  AOI22_X1 U20036 ( .A1(n16896), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9613), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16897) );
  NAND4_X1 U20037 ( .A1(n16900), .A2(n16899), .A3(n16898), .A4(n16897), .ZN(
        n16901) );
  AOI211_X1 U20038 ( .C1(n16954), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n16902), .B(n16901), .ZN(n16903) );
  NAND2_X1 U20039 ( .A1(n16904), .A2(n16903), .ZN(n17096) );
  INV_X1 U20040 ( .A(n17096), .ZN(n16908) );
  INV_X1 U20041 ( .A(n16923), .ZN(n16906) );
  OAI21_X1 U20042 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n16906), .A(n16905), .ZN(
        n16907) );
  OAI21_X1 U20043 ( .B1(n16908), .B2(n16986), .A(n16907), .ZN(P3_U2692) );
  AOI22_X1 U20044 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16922) );
  AOI22_X1 U20045 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16921) );
  AOI22_X1 U20046 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16910) );
  OAI21_X1 U20047 ( .B1(n16912), .B2(n16911), .A(n16910), .ZN(n16919) );
  AOI22_X1 U20048 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16917) );
  AOI22_X1 U20049 ( .A1(n9614), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16895), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16916) );
  AOI22_X1 U20050 ( .A1(n16913), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16915) );
  AOI22_X1 U20051 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16914) );
  NAND4_X1 U20052 ( .A1(n16917), .A2(n16916), .A3(n16915), .A4(n16914), .ZN(
        n16918) );
  AOI211_X1 U20053 ( .C1(n16936), .C2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n16919), .B(n16918), .ZN(n16920) );
  NAND3_X1 U20054 ( .A1(n16922), .A2(n16921), .A3(n16920), .ZN(n17099) );
  INV_X1 U20055 ( .A(n17099), .ZN(n16925) );
  OAI21_X1 U20056 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n16945), .A(n16923), .ZN(
        n16924) );
  AOI22_X1 U20057 ( .A1(n16992), .A2(n16925), .B1(n16924), .B2(n16986), .ZN(
        P3_U2693) );
  INV_X1 U20058 ( .A(n16926), .ZN(n16961) );
  OAI21_X1 U20059 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n16961), .A(n16986), .ZN(
        n16944) );
  AOI22_X1 U20060 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n9613), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n16927), .ZN(n16933) );
  AOI22_X1 U20061 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n13753), .B1(
        n9615), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16932) );
  AOI22_X1 U20062 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n16928), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n13732), .ZN(n16931) );
  AOI22_X1 U20063 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n16895), .ZN(n16930) );
  NAND4_X1 U20064 ( .A1(n16933), .A2(n16932), .A3(n16931), .A4(n16930), .ZN(
        n16943) );
  AOI22_X1 U20065 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16941) );
  AOI22_X1 U20066 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n16947), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n16940) );
  AOI22_X1 U20067 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n9628), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n16939) );
  AOI22_X1 U20068 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n16937), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n15053), .ZN(n16938) );
  NAND4_X1 U20069 ( .A1(n16941), .A2(n16940), .A3(n16939), .A4(n16938), .ZN(
        n16942) );
  NOR2_X1 U20070 ( .A1(n16943), .A2(n16942), .ZN(n17104) );
  OAI22_X1 U20071 ( .A1(n16945), .A2(n16944), .B1(n17104), .B2(n16986), .ZN(
        P3_U2694) );
  AOI22_X1 U20072 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13753), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16952) );
  AOI22_X1 U20073 ( .A1(n9614), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16895), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16951) );
  AOI22_X1 U20074 ( .A1(n16947), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16946), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16950) );
  AOI22_X1 U20075 ( .A1(n16948), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16913), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16949) );
  NAND4_X1 U20076 ( .A1(n16952), .A2(n16951), .A3(n16950), .A4(n16949), .ZN(
        n16960) );
  AOI22_X1 U20077 ( .A1(n16935), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16958) );
  AOI22_X1 U20078 ( .A1(n9628), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16957) );
  AOI22_X1 U20079 ( .A1(n9615), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16956) );
  AOI22_X1 U20080 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15053), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16955) );
  NAND4_X1 U20081 ( .A1(n16958), .A2(n16957), .A3(n16956), .A4(n16955), .ZN(
        n16959) );
  NOR2_X1 U20082 ( .A1(n16960), .A2(n16959), .ZN(n17110) );
  AOI21_X1 U20083 ( .B1(n20811), .B2(n16962), .A(n16961), .ZN(n16963) );
  INV_X1 U20084 ( .A(n16963), .ZN(n16964) );
  AOI22_X1 U20085 ( .A1(n16992), .A2(n17110), .B1(n16964), .B2(n16986), .ZN(
        P3_U2695) );
  AOI22_X1 U20086 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n16986), .B1(
        P3_EBX_REG_6__SCAN_IN), .B2(n16969), .ZN(n16966) );
  INV_X1 U20087 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16965) );
  OAI22_X1 U20088 ( .A1(n16967), .A2(n16966), .B1(n16965), .B2(n16986), .ZN(
        P3_U2696) );
  NAND2_X1 U20089 ( .A1(n16986), .A2(n16968), .ZN(n16973) );
  AOI22_X1 U20090 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n16992), .B1(
        n16969), .B2(n16971), .ZN(n16970) );
  OAI21_X1 U20091 ( .B1(n16971), .B2(n16973), .A(n16970), .ZN(P3_U2697) );
  NOR2_X1 U20092 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n16978), .ZN(n16974) );
  INV_X1 U20093 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16972) );
  OAI22_X1 U20094 ( .A1(n16974), .A2(n16973), .B1(n16972), .B2(n16986), .ZN(
        P3_U2698) );
  INV_X1 U20095 ( .A(n16988), .ZN(n16994) );
  NOR3_X1 U20096 ( .A1(n16984), .A2(n16975), .A3(n16994), .ZN(n16982) );
  AND2_X1 U20097 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n16982), .ZN(n16981) );
  AOI21_X1 U20098 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n16986), .A(n16981), .ZN(
        n16977) );
  OAI22_X1 U20099 ( .A1(n16978), .A2(n16977), .B1(n16976), .B2(n16986), .ZN(
        P3_U2699) );
  AOI21_X1 U20100 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n16986), .A(n16982), .ZN(
        n16980) );
  INV_X1 U20101 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16979) );
  OAI22_X1 U20102 ( .A1(n16981), .A2(n16980), .B1(n16979), .B2(n16986), .ZN(
        P3_U2700) );
  AOI21_X1 U20103 ( .B1(n16984), .B2(n16983), .A(n16982), .ZN(n16985) );
  OAI22_X1 U20104 ( .A1(n16986), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16985), .B2(n16992), .ZN(n16987) );
  INV_X1 U20105 ( .A(n16987), .ZN(P3_U2701) );
  AOI222_X1 U20106 ( .A1(n16989), .A2(n16988), .B1(P3_EBX_REG_1__SCAN_IN), 
        .B2(n16991), .C1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .C2(n16992), .ZN(
        n16990) );
  INV_X1 U20107 ( .A(n16990), .ZN(P3_U2702) );
  AOI22_X1 U20108 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n16992), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n16991), .ZN(n16993) );
  OAI21_X1 U20109 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n16994), .A(n16993), .ZN(
        P3_U2703) );
  INV_X1 U20110 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17215) );
  INV_X1 U20111 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17210) );
  INV_X1 U20112 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17202) );
  INV_X1 U20113 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17252) );
  INV_X1 U20114 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17227) );
  NAND4_X1 U20115 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(P3_EAX_REG_5__SCAN_IN), .ZN(n16995) );
  NOR2_X1 U20116 ( .A1(n17227), .A2(n16995), .ZN(n17109) );
  NAND3_X1 U20117 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(n17109), .ZN(n17081) );
  AND4_X1 U20118 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n16996)
         );
  NAND4_X1 U20119 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17112), .A3(
        P3_EAX_REG_14__SCAN_IN), .A4(n16996), .ZN(n17083) );
  NOR2_X2 U20120 ( .A1(n17252), .A2(n17083), .ZN(n17077) );
  INV_X1 U20121 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17200) );
  INV_X1 U20122 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17198) );
  NOR2_X1 U20123 ( .A1(n17200), .A2(n17198), .ZN(n16997) );
  NAND4_X1 U20124 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .A4(n16997), .ZN(n17039) );
  NAND2_X1 U20125 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17035), .ZN(n17034) );
  NAND2_X1 U20126 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17030), .ZN(n17029) );
  NAND2_X1 U20127 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17019), .ZN(n17015) );
  NAND2_X1 U20128 ( .A1(n17004), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17000) );
  NOR2_X2 U20129 ( .A1(n17997), .A2(n17143), .ZN(n17071) );
  OAI22_X1 U20130 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17040), .B1(n17134), 
        .B2(n17004), .ZN(n16998) );
  AOI22_X1 U20131 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17071), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n16998), .ZN(n16999) );
  OAI21_X1 U20132 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17000), .A(n16999), .ZN(
        P3_U2704) );
  NAND2_X1 U20133 ( .A1(n17993), .A2(n17134), .ZN(n17046) );
  AOI22_X1 U20134 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17072), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17071), .ZN(n17002) );
  OAI211_X1 U20135 ( .C1(n17004), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17143), .B(
        n17000), .ZN(n17001) );
  OAI211_X1 U20136 ( .C1(n17003), .C2(n17137), .A(n17002), .B(n17001), .ZN(
        P3_U2705) );
  INV_X1 U20137 ( .A(n17004), .ZN(n17006) );
  OAI21_X1 U20138 ( .B1(n17134), .B2(n17215), .A(n17011), .ZN(n17005) );
  AOI22_X1 U20139 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n17071), .B1(n17006), .B2(
        n17005), .ZN(n17009) );
  AOI22_X1 U20140 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17072), .B1(n17007), .B2(
        n17140), .ZN(n17008) );
  NAND2_X1 U20141 ( .A1(n17009), .A2(n17008), .ZN(P3_U2706) );
  AOI22_X1 U20142 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n17071), .B1(n17010), .B2(
        n17140), .ZN(n17014) );
  OAI211_X1 U20143 ( .C1(n17012), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17143), .B(
        n17011), .ZN(n17013) );
  OAI211_X1 U20144 ( .C1(n17046), .C2(n17095), .A(n17014), .B(n17013), .ZN(
        P3_U2707) );
  AOI22_X1 U20145 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17072), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17071), .ZN(n17017) );
  OAI211_X1 U20146 ( .C1(n17019), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17143), .B(
        n17015), .ZN(n17016) );
  OAI211_X1 U20147 ( .C1(n17137), .C2(n17018), .A(n17017), .B(n17016), .ZN(
        P3_U2708) );
  AOI22_X1 U20148 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17072), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17071), .ZN(n17022) );
  AOI211_X1 U20149 ( .C1(n17210), .C2(n17024), .A(n17019), .B(n17134), .ZN(
        n17020) );
  INV_X1 U20150 ( .A(n17020), .ZN(n17021) );
  OAI211_X1 U20151 ( .C1(n17137), .C2(n17023), .A(n17022), .B(n17021), .ZN(
        P3_U2709) );
  AOI22_X1 U20152 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17072), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17071), .ZN(n17027) );
  OAI211_X1 U20153 ( .C1(n17025), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17143), .B(
        n17024), .ZN(n17026) );
  OAI211_X1 U20154 ( .C1(n17137), .C2(n17028), .A(n17027), .B(n17026), .ZN(
        P3_U2710) );
  AOI22_X1 U20155 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17072), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17071), .ZN(n17032) );
  OAI211_X1 U20156 ( .C1(n17030), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17143), .B(
        n17029), .ZN(n17031) );
  OAI211_X1 U20157 ( .C1(n17137), .C2(n17033), .A(n17032), .B(n17031), .ZN(
        P3_U2711) );
  AOI22_X1 U20158 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17072), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17071), .ZN(n17037) );
  OAI211_X1 U20159 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17035), .A(n17143), .B(
        n17034), .ZN(n17036) );
  OAI211_X1 U20160 ( .C1(n17137), .C2(n17038), .A(n17037), .B(n17036), .ZN(
        P3_U2712) );
  NOR3_X1 U20161 ( .A1(n17108), .A2(n17073), .A3(n17039), .ZN(n17044) );
  INV_X1 U20162 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17196) );
  INV_X1 U20163 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17192) );
  NAND2_X1 U20164 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17065), .ZN(n17061) );
  NAND2_X1 U20165 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17056), .ZN(n17052) );
  NAND2_X1 U20166 ( .A1(n17143), .A2(n17052), .ZN(n17051) );
  OAI21_X1 U20167 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17040), .A(n17051), .ZN(
        n17043) );
  INV_X1 U20168 ( .A(n17071), .ZN(n17047) );
  OAI22_X1 U20169 ( .A1(n17041), .A2(n17137), .B1(n18973), .B2(n17047), .ZN(
        n17042) );
  AOI221_X1 U20170 ( .B1(n17044), .B2(n17202), .C1(n17043), .C2(
        P3_EAX_REG_22__SCAN_IN), .A(n17042), .ZN(n17045) );
  OAI21_X1 U20171 ( .B1(n17996), .B2(n17046), .A(n17045), .ZN(P3_U2713) );
  OAI22_X1 U20172 ( .A1(n17048), .A2(n17137), .B1(n13674), .B2(n17047), .ZN(
        n17049) );
  AOI21_X1 U20173 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17072), .A(n17049), .ZN(
        n17050) );
  OAI221_X1 U20174 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17052), .C1(n17200), 
        .C2(n17051), .A(n17050), .ZN(P3_U2714) );
  AOI22_X1 U20175 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17072), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17071), .ZN(n17054) );
  OAI211_X1 U20176 ( .C1(n17056), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17143), .B(
        n17052), .ZN(n17053) );
  OAI211_X1 U20177 ( .C1(n17055), .C2(n17137), .A(n17054), .B(n17053), .ZN(
        P3_U2715) );
  AOI22_X1 U20178 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17072), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17071), .ZN(n17059) );
  AOI211_X1 U20179 ( .C1(n17196), .C2(n17061), .A(n17056), .B(n17134), .ZN(
        n17057) );
  INV_X1 U20180 ( .A(n17057), .ZN(n17058) );
  OAI211_X1 U20181 ( .C1(n17060), .C2(n17137), .A(n17059), .B(n17058), .ZN(
        P3_U2716) );
  AOI22_X1 U20182 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17072), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17071), .ZN(n17063) );
  OAI211_X1 U20183 ( .C1(n17065), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17143), .B(
        n17061), .ZN(n17062) );
  OAI211_X1 U20184 ( .C1(n17064), .C2(n17137), .A(n17063), .B(n17062), .ZN(
        P3_U2717) );
  AOI22_X1 U20185 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17072), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17071), .ZN(n17069) );
  INV_X1 U20186 ( .A(n17073), .ZN(n17067) );
  INV_X1 U20187 ( .A(n17065), .ZN(n17066) );
  OAI211_X1 U20188 ( .C1(n17067), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17143), .B(
        n17066), .ZN(n17068) );
  OAI211_X1 U20189 ( .C1(n17070), .C2(n17137), .A(n17069), .B(n17068), .ZN(
        P3_U2718) );
  AOI22_X1 U20190 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17072), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17071), .ZN(n17075) );
  OAI211_X1 U20191 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17077), .A(n17143), .B(
        n17073), .ZN(n17074) );
  OAI211_X1 U20192 ( .C1(n17076), .C2(n17137), .A(n17075), .B(n17074), .ZN(
        P3_U2719) );
  AOI211_X1 U20193 ( .C1(n17252), .C2(n17083), .A(n17134), .B(n17077), .ZN(
        n17078) );
  AOI21_X1 U20194 ( .B1(n17141), .B2(BUF2_REG_15__SCAN_IN), .A(n17078), .ZN(
        n17079) );
  OAI21_X1 U20195 ( .B1(n17080), .B2(n17137), .A(n17079), .ZN(P3_U2720) );
  INV_X1 U20196 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n20792) );
  NOR3_X1 U20197 ( .A1(n17108), .A2(n17142), .A3(n17081), .ZN(n17103) );
  NAND2_X1 U20198 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17103), .ZN(n17101) );
  INV_X1 U20199 ( .A(n17101), .ZN(n17106) );
  NAND2_X1 U20200 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17106), .ZN(n17098) );
  NOR2_X1 U20201 ( .A1(n20792), .A2(n17098), .ZN(n17091) );
  NAND2_X1 U20202 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17094), .ZN(n17086) );
  AOI22_X1 U20203 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17141), .B1(n17140), .B2(
        n17082), .ZN(n17085) );
  NAND3_X1 U20204 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17143), .A3(n17083), 
        .ZN(n17084) );
  OAI211_X1 U20205 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17086), .A(n17085), .B(
        n17084), .ZN(P3_U2721) );
  INV_X1 U20206 ( .A(n17086), .ZN(n17089) );
  AOI21_X1 U20207 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17143), .A(n17094), .ZN(
        n17088) );
  OAI222_X1 U20208 ( .A1(n17132), .A2(n17090), .B1(n17089), .B2(n17088), .C1(
        n17137), .C2(n17087), .ZN(P3_U2722) );
  AOI21_X1 U20209 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17143), .A(n17091), .ZN(
        n17093) );
  OAI222_X1 U20210 ( .A1(n17132), .A2(n17095), .B1(n17094), .B2(n17093), .C1(
        n17137), .C2(n17092), .ZN(P3_U2723) );
  NAND2_X1 U20211 ( .A1(n17143), .A2(n17098), .ZN(n17102) );
  AOI22_X1 U20212 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17141), .B1(n17140), .B2(
        n17096), .ZN(n17097) );
  OAI221_X1 U20213 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17098), .C1(n20792), 
        .C2(n17102), .A(n17097), .ZN(P3_U2724) );
  INV_X1 U20214 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17239) );
  AOI22_X1 U20215 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17141), .B1(n17140), .B2(
        n17099), .ZN(n17100) );
  OAI221_X1 U20216 ( .B1(n17102), .B2(n17239), .C1(n17102), .C2(n17101), .A(
        n17100), .ZN(P3_U2725) );
  AOI21_X1 U20217 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17143), .A(n17103), .ZN(
        n17105) );
  OAI222_X1 U20218 ( .A1(n17132), .A2(n17107), .B1(n17106), .B2(n17105), .C1(
        n17137), .C2(n17104), .ZN(P3_U2726) );
  NOR2_X1 U20219 ( .A1(n17108), .A2(n17142), .ZN(n17117) );
  AND2_X1 U20220 ( .A1(n17109), .A2(n17117), .ZN(n17120) );
  AOI22_X1 U20221 ( .A1(n17120), .A2(P3_EAX_REG_7__SCAN_IN), .B1(
        P3_EAX_REG_8__SCAN_IN), .B2(n17143), .ZN(n17111) );
  OAI222_X1 U20222 ( .A1(n17132), .A2(n17113), .B1(n17112), .B2(n17111), .C1(
        n17137), .C2(n17110), .ZN(P3_U2727) );
  AND2_X1 U20223 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17120), .ZN(n17116) );
  AOI21_X1 U20224 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17143), .A(n17120), .ZN(
        n17115) );
  OAI222_X1 U20225 ( .A1(n18002), .A2(n17132), .B1(n17116), .B2(n17115), .C1(
        n17137), .C2(n17114), .ZN(P3_U2728) );
  INV_X1 U20226 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17229) );
  INV_X1 U20227 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17225) );
  NAND2_X1 U20228 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17117), .ZN(n17128) );
  NOR2_X1 U20229 ( .A1(n17225), .A2(n17128), .ZN(n17131) );
  NAND2_X1 U20230 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17131), .ZN(n17121) );
  NOR2_X1 U20231 ( .A1(n17229), .A2(n17121), .ZN(n17124) );
  AOI21_X1 U20232 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17143), .A(n17124), .ZN(
        n17119) );
  OAI222_X1 U20233 ( .A1(n17996), .A2(n17132), .B1(n17120), .B2(n17119), .C1(
        n17137), .C2(n17118), .ZN(P3_U2729) );
  INV_X1 U20234 ( .A(n17121), .ZN(n17127) );
  AOI21_X1 U20235 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17143), .A(n17127), .ZN(
        n17123) );
  OAI222_X1 U20236 ( .A1(n17992), .A2(n17132), .B1(n17124), .B2(n17123), .C1(
        n17137), .C2(n17122), .ZN(P3_U2730) );
  AOI21_X1 U20237 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17143), .A(n17131), .ZN(
        n17126) );
  OAI222_X1 U20238 ( .A1(n17988), .A2(n17132), .B1(n17127), .B2(n17126), .C1(
        n17137), .C2(n17125), .ZN(P3_U2731) );
  INV_X1 U20239 ( .A(n17128), .ZN(n17133) );
  AOI21_X1 U20240 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17143), .A(n17133), .ZN(
        n17130) );
  OAI222_X1 U20241 ( .A1(n17984), .A2(n17132), .B1(n17131), .B2(n17130), .C1(
        n17137), .C2(n17129), .ZN(P3_U2732) );
  INV_X1 U20242 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17223) );
  AOI211_X1 U20243 ( .C1(n17142), .C2(n17223), .A(n17134), .B(n17133), .ZN(
        n17135) );
  AOI21_X1 U20244 ( .B1(n17141), .B2(BUF2_REG_2__SCAN_IN), .A(n17135), .ZN(
        n17136) );
  OAI21_X1 U20245 ( .B1(n17138), .B2(n17137), .A(n17136), .ZN(P3_U2733) );
  AOI22_X1 U20246 ( .A1(n17141), .A2(BUF2_REG_1__SCAN_IN), .B1(n17140), .B2(
        n17139), .ZN(n17146) );
  OAI211_X1 U20247 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n17144), .A(n17143), .B(
        n17142), .ZN(n17145) );
  NAND2_X1 U20248 ( .A1(n17146), .A2(n17145), .ZN(P3_U2734) );
  NAND2_X1 U20249 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17455), .ZN(n18616) );
  INV_X2 U20250 ( .A(n18616), .ZN(n17182) );
  INV_X1 U20251 ( .A(n17186), .ZN(n17185) );
  AND2_X1 U20252 ( .A1(n17175), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20253 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17217) );
  NAND2_X1 U20254 ( .A1(n17166), .A2(n17971), .ZN(n17163) );
  AOI22_X1 U20255 ( .A1(n17182), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17148) );
  OAI21_X1 U20256 ( .B1(n17217), .B2(n17163), .A(n17148), .ZN(P3_U2737) );
  AOI22_X1 U20257 ( .A1(n17182), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17149) );
  OAI21_X1 U20258 ( .B1(n17215), .B2(n17163), .A(n17149), .ZN(P3_U2738) );
  INV_X1 U20259 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n20791) );
  AOI22_X1 U20260 ( .A1(n17182), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17175), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17150) );
  OAI21_X1 U20261 ( .B1(n20791), .B2(n17163), .A(n17150), .ZN(P3_U2739) );
  INV_X1 U20262 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17212) );
  AOI22_X1 U20263 ( .A1(n17182), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17175), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17151) );
  OAI21_X1 U20264 ( .B1(n17212), .B2(n17163), .A(n17151), .ZN(P3_U2740) );
  AOI22_X1 U20265 ( .A1(n17182), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17175), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17152) );
  OAI21_X1 U20266 ( .B1(n17210), .B2(n17163), .A(n17152), .ZN(P3_U2741) );
  INV_X1 U20267 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17208) );
  AOI22_X1 U20268 ( .A1(n17182), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17175), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17153) );
  OAI21_X1 U20269 ( .B1(n17208), .B2(n17163), .A(n17153), .ZN(P3_U2742) );
  INV_X1 U20270 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17206) );
  AOI22_X1 U20271 ( .A1(n17182), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17175), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17154) );
  OAI21_X1 U20272 ( .B1(n17206), .B2(n17163), .A(n17154), .ZN(P3_U2743) );
  INV_X1 U20273 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17204) );
  AOI22_X1 U20274 ( .A1(n17182), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17155) );
  OAI21_X1 U20275 ( .B1(n17204), .B2(n17163), .A(n17155), .ZN(P3_U2744) );
  AOI22_X1 U20276 ( .A1(n17182), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17156) );
  OAI21_X1 U20277 ( .B1(n17202), .B2(n17163), .A(n17156), .ZN(P3_U2745) );
  AOI22_X1 U20278 ( .A1(n17182), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17157) );
  OAI21_X1 U20279 ( .B1(n17200), .B2(n17163), .A(n17157), .ZN(P3_U2746) );
  AOI22_X1 U20280 ( .A1(n17182), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17158) );
  OAI21_X1 U20281 ( .B1(n17198), .B2(n17163), .A(n17158), .ZN(P3_U2747) );
  AOI22_X1 U20282 ( .A1(n17182), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17159) );
  OAI21_X1 U20283 ( .B1(n17196), .B2(n17163), .A(n17159), .ZN(P3_U2748) );
  INV_X1 U20284 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17194) );
  AOI22_X1 U20285 ( .A1(n17182), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17160) );
  OAI21_X1 U20286 ( .B1(n17194), .B2(n17163), .A(n17160), .ZN(P3_U2749) );
  AOI22_X1 U20287 ( .A1(n17182), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17161) );
  OAI21_X1 U20288 ( .B1(n17192), .B2(n17163), .A(n17161), .ZN(P3_U2750) );
  INV_X1 U20289 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17190) );
  AOI22_X1 U20290 ( .A1(n17182), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17162) );
  OAI21_X1 U20291 ( .B1(n17190), .B2(n17163), .A(n17162), .ZN(P3_U2751) );
  AOI22_X1 U20292 ( .A1(n17182), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17164) );
  OAI21_X1 U20293 ( .B1(n17252), .B2(n17184), .A(n17164), .ZN(P3_U2752) );
  INV_X1 U20294 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U20295 ( .A1(n17182), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17165) );
  OAI21_X1 U20296 ( .B1(n17248), .B2(n17184), .A(n17165), .ZN(P3_U2753) );
  INV_X1 U20297 ( .A(P3_LWORD_REG_13__SCAN_IN), .ZN(n20757) );
  AOI22_X1 U20298 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17166), .B1(n17181), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17167) );
  OAI21_X1 U20299 ( .B1(n20757), .B2(n18616), .A(n17167), .ZN(P3_U2754) );
  INV_X1 U20300 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17243) );
  AOI22_X1 U20301 ( .A1(n17182), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17168) );
  OAI21_X1 U20302 ( .B1(n17243), .B2(n17184), .A(n17168), .ZN(P3_U2755) );
  AOI22_X1 U20303 ( .A1(n17182), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17169) );
  OAI21_X1 U20304 ( .B1(n20792), .B2(n17184), .A(n17169), .ZN(P3_U2756) );
  AOI22_X1 U20305 ( .A1(P3_LWORD_REG_10__SCAN_IN), .A2(n17182), .B1(n17181), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17170) );
  OAI21_X1 U20306 ( .B1(n17239), .B2(n17184), .A(n17170), .ZN(P3_U2757) );
  INV_X1 U20307 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17237) );
  AOI22_X1 U20308 ( .A1(n17182), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17175), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17171) );
  OAI21_X1 U20309 ( .B1(n17237), .B2(n17184), .A(n17171), .ZN(P3_U2758) );
  INV_X1 U20310 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17235) );
  AOI22_X1 U20311 ( .A1(n17182), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17175), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17172) );
  OAI21_X1 U20312 ( .B1(n17235), .B2(n17184), .A(n17172), .ZN(P3_U2759) );
  INV_X1 U20313 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17233) );
  AOI22_X1 U20314 ( .A1(n17182), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17175), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17173) );
  OAI21_X1 U20315 ( .B1(n17233), .B2(n17184), .A(n17173), .ZN(P3_U2760) );
  INV_X1 U20316 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17231) );
  AOI22_X1 U20317 ( .A1(n17182), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17175), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17174) );
  OAI21_X1 U20318 ( .B1(n17231), .B2(n17184), .A(n17174), .ZN(P3_U2761) );
  AOI22_X1 U20319 ( .A1(n17182), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17175), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17176) );
  OAI21_X1 U20320 ( .B1(n17229), .B2(n17184), .A(n17176), .ZN(P3_U2762) );
  AOI22_X1 U20321 ( .A1(n17182), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17177) );
  OAI21_X1 U20322 ( .B1(n17227), .B2(n17184), .A(n17177), .ZN(P3_U2763) );
  AOI22_X1 U20323 ( .A1(n17182), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17178) );
  OAI21_X1 U20324 ( .B1(n17225), .B2(n17184), .A(n17178), .ZN(P3_U2764) );
  AOI22_X1 U20325 ( .A1(n17182), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17179) );
  OAI21_X1 U20326 ( .B1(n17223), .B2(n17184), .A(n17179), .ZN(P3_U2765) );
  INV_X1 U20327 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17221) );
  AOI22_X1 U20328 ( .A1(n17182), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17180) );
  OAI21_X1 U20329 ( .B1(n17221), .B2(n17184), .A(n17180), .ZN(P3_U2766) );
  AOI22_X1 U20330 ( .A1(n17182), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17181), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17183) );
  OAI21_X1 U20331 ( .B1(n17219), .B2(n17184), .A(n17183), .ZN(P3_U2767) );
  NOR2_X1 U20332 ( .A1(n17188), .A2(n17187), .ZN(n18460) );
  INV_X2 U20333 ( .A(n17244), .ZN(n17251) );
  AOI211_X1 U20334 ( .C1(n17188), .C2(n18617), .A(n17187), .B(n17186), .ZN(
        n17246) );
  INV_X2 U20335 ( .A(n17246), .ZN(n17249) );
  AOI22_X1 U20336 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17241), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17249), .ZN(n17189) );
  OAI21_X1 U20337 ( .B1(n17190), .B2(n17251), .A(n17189), .ZN(P3_U2768) );
  AOI22_X1 U20338 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17241), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17249), .ZN(n17191) );
  OAI21_X1 U20339 ( .B1(n17192), .B2(n17251), .A(n17191), .ZN(P3_U2769) );
  AOI22_X1 U20340 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17241), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17249), .ZN(n17193) );
  OAI21_X1 U20341 ( .B1(n17194), .B2(n17251), .A(n17193), .ZN(P3_U2770) );
  AOI22_X1 U20342 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n9636), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17249), .ZN(n17195) );
  OAI21_X1 U20343 ( .B1(n17196), .B2(n17251), .A(n17195), .ZN(P3_U2771) );
  AOI22_X1 U20344 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n9636), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17249), .ZN(n17197) );
  OAI21_X1 U20345 ( .B1(n17198), .B2(n17251), .A(n17197), .ZN(P3_U2772) );
  AOI22_X1 U20346 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n9636), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17249), .ZN(n17199) );
  OAI21_X1 U20347 ( .B1(n17200), .B2(n17251), .A(n17199), .ZN(P3_U2773) );
  AOI22_X1 U20348 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n9636), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17249), .ZN(n17201) );
  OAI21_X1 U20349 ( .B1(n17202), .B2(n17251), .A(n17201), .ZN(P3_U2774) );
  AOI22_X1 U20350 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n9636), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17249), .ZN(n17203) );
  OAI21_X1 U20351 ( .B1(n17204), .B2(n17251), .A(n17203), .ZN(P3_U2775) );
  AOI22_X1 U20352 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n9636), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17249), .ZN(n17205) );
  OAI21_X1 U20353 ( .B1(n17206), .B2(n17251), .A(n17205), .ZN(P3_U2776) );
  AOI22_X1 U20354 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n9636), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17249), .ZN(n17207) );
  OAI21_X1 U20355 ( .B1(n17208), .B2(n17251), .A(n17207), .ZN(P3_U2777) );
  AOI22_X1 U20356 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n9636), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17249), .ZN(n17209) );
  OAI21_X1 U20357 ( .B1(n17210), .B2(n17251), .A(n17209), .ZN(P3_U2778) );
  AOI22_X1 U20358 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n9636), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17249), .ZN(n17211) );
  OAI21_X1 U20359 ( .B1(n17212), .B2(n17251), .A(n17211), .ZN(P3_U2779) );
  AOI22_X1 U20360 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17241), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17249), .ZN(n17213) );
  OAI21_X1 U20361 ( .B1(n20791), .B2(n17251), .A(n17213), .ZN(P3_U2780) );
  AOI22_X1 U20362 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17241), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17249), .ZN(n17214) );
  OAI21_X1 U20363 ( .B1(n17215), .B2(n17251), .A(n17214), .ZN(P3_U2781) );
  AOI22_X1 U20364 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17241), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17249), .ZN(n17216) );
  OAI21_X1 U20365 ( .B1(n17217), .B2(n17251), .A(n17216), .ZN(P3_U2782) );
  AOI22_X1 U20366 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17241), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17249), .ZN(n17218) );
  OAI21_X1 U20367 ( .B1(n17219), .B2(n17251), .A(n17218), .ZN(P3_U2783) );
  AOI22_X1 U20368 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17241), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17249), .ZN(n17220) );
  OAI21_X1 U20369 ( .B1(n17221), .B2(n17251), .A(n17220), .ZN(P3_U2784) );
  AOI22_X1 U20370 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17241), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17249), .ZN(n17222) );
  OAI21_X1 U20371 ( .B1(n17223), .B2(n17251), .A(n17222), .ZN(P3_U2785) );
  AOI22_X1 U20372 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17241), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17249), .ZN(n17224) );
  OAI21_X1 U20373 ( .B1(n17225), .B2(n17251), .A(n17224), .ZN(P3_U2786) );
  AOI22_X1 U20374 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17241), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17249), .ZN(n17226) );
  OAI21_X1 U20375 ( .B1(n17227), .B2(n17251), .A(n17226), .ZN(P3_U2787) );
  AOI22_X1 U20376 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17241), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17249), .ZN(n17228) );
  OAI21_X1 U20377 ( .B1(n17229), .B2(n17251), .A(n17228), .ZN(P3_U2788) );
  AOI22_X1 U20378 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17241), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17249), .ZN(n17230) );
  OAI21_X1 U20379 ( .B1(n17231), .B2(n17251), .A(n17230), .ZN(P3_U2789) );
  AOI22_X1 U20380 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17241), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17249), .ZN(n17232) );
  OAI21_X1 U20381 ( .B1(n17233), .B2(n17251), .A(n17232), .ZN(P3_U2790) );
  AOI22_X1 U20382 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17241), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17249), .ZN(n17234) );
  OAI21_X1 U20383 ( .B1(n17235), .B2(n17251), .A(n17234), .ZN(P3_U2791) );
  AOI22_X1 U20384 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17241), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17249), .ZN(n17236) );
  OAI21_X1 U20385 ( .B1(n17237), .B2(n17251), .A(n17236), .ZN(P3_U2792) );
  AOI22_X1 U20386 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n9636), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17249), .ZN(n17238) );
  OAI21_X1 U20387 ( .B1(n17239), .B2(n17251), .A(n17238), .ZN(P3_U2793) );
  AOI22_X1 U20388 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17241), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17249), .ZN(n17240) );
  OAI21_X1 U20389 ( .B1(n20792), .B2(n17251), .A(n17240), .ZN(P3_U2794) );
  AOI22_X1 U20390 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n9636), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17249), .ZN(n17242) );
  OAI21_X1 U20391 ( .B1(n17243), .B2(n17251), .A(n17242), .ZN(P3_U2795) );
  AOI22_X1 U20392 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17241), .B1(
        P3_EAX_REG_13__SCAN_IN), .B2(n17244), .ZN(n17245) );
  OAI21_X1 U20393 ( .B1(n17246), .B2(n20757), .A(n17245), .ZN(P3_U2796) );
  AOI22_X1 U20394 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17241), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17249), .ZN(n17247) );
  OAI21_X1 U20395 ( .B1(n17248), .B2(n17251), .A(n17247), .ZN(P3_U2797) );
  AOI22_X1 U20396 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17241), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17249), .ZN(n17250) );
  OAI21_X1 U20397 ( .B1(n17252), .B2(n17251), .A(n17250), .ZN(P3_U2798) );
  INV_X1 U20398 ( .A(n17259), .ZN(n17253) );
  OAI21_X1 U20399 ( .B1(n17253), .B2(n17523), .A(n17625), .ZN(n17254) );
  AOI21_X1 U20400 ( .B1(n17455), .B2(n17255), .A(n17254), .ZN(n17285) );
  OAI21_X1 U20401 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17365), .A(
        n17285), .ZN(n17272) );
  AOI211_X1 U20402 ( .C1(n17258), .C2(n17257), .A(n17256), .B(n17508), .ZN(
        n17265) );
  NOR2_X1 U20403 ( .A1(n17379), .A2(n17259), .ZN(n17277) );
  OAI211_X1 U20404 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17277), .B(n17260), .ZN(n17262) );
  OAI211_X1 U20405 ( .C1(n17461), .C2(n17263), .A(n17262), .B(n17261), .ZN(
        n17264) );
  AOI211_X1 U20406 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17272), .A(
        n17265), .B(n17264), .ZN(n17268) );
  NOR2_X1 U20407 ( .A1(n17613), .A2(n17452), .ZN(n17371) );
  INV_X1 U20408 ( .A(n17371), .ZN(n17341) );
  AOI22_X1 U20409 ( .A1(n17613), .A2(n17633), .B1(n17452), .B2(n17632), .ZN(
        n17286) );
  NAND2_X1 U20410 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17286), .ZN(
        n17266) );
  NAND3_X1 U20411 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17341), .A3(
        n17266), .ZN(n17267) );
  OAI211_X1 U20412 ( .C1(n17426), .C2(n17269), .A(n17268), .B(n17267), .ZN(
        P3_U2802) );
  XNOR2_X1 U20413 ( .A(n17271), .B(n17516), .ZN(n17643) );
  AOI22_X1 U20414 ( .A1(n17482), .A2(n17273), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17272), .ZN(n17274) );
  NAND2_X1 U20415 ( .A1(n17951), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17641) );
  OAI211_X1 U20416 ( .C1(n17643), .C2(n17508), .A(n17274), .B(n17641), .ZN(
        n17275) );
  AOI21_X1 U20417 ( .B1(n17277), .B2(n17276), .A(n17275), .ZN(n17278) );
  OAI221_X1 U20418 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17280), 
        .C1(n17279), .C2(n17286), .A(n17278), .ZN(P3_U2803) );
  AOI21_X1 U20419 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17282), .A(
        n17281), .ZN(n17652) );
  NAND2_X1 U20420 ( .A1(n17461), .A2(n17365), .ZN(n17616) );
  AOI21_X1 U20421 ( .B1(n17283), .B2(n18000), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17284) );
  OAI22_X1 U20422 ( .A1(n17285), .A2(n17284), .B1(n17861), .B2(n18542), .ZN(
        n17290) );
  NAND2_X1 U20423 ( .A1(n17300), .A2(n17644), .ZN(n17634) );
  NOR2_X1 U20424 ( .A1(n17426), .A2(n17634), .ZN(n17288) );
  INV_X1 U20425 ( .A(n17286), .ZN(n17287) );
  MUX2_X1 U20426 ( .A(n17288), .B(n17287), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n17289) );
  AOI211_X1 U20427 ( .C1(n17291), .C2(n17616), .A(n17290), .B(n17289), .ZN(
        n17292) );
  OAI21_X1 U20428 ( .B1(n17652), .B2(n17508), .A(n17292), .ZN(P3_U2804) );
  NOR2_X1 U20429 ( .A1(n17301), .A2(n17672), .ZN(n17293) );
  XNOR2_X1 U20430 ( .A(n17293), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17667) );
  OAI21_X1 U20431 ( .B1(n17294), .B2(n17624), .A(n17625), .ZN(n17295) );
  AOI21_X1 U20432 ( .B1(n18000), .B2(n17296), .A(n17295), .ZN(n17328) );
  OAI21_X1 U20433 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17365), .A(
        n17328), .ZN(n17310) );
  NOR2_X1 U20434 ( .A1(n17379), .A2(n17296), .ZN(n17311) );
  OAI211_X1 U20435 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17311), .B(n17297), .ZN(n17298) );
  NAND2_X1 U20436 ( .A1(n17951), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17661) );
  OAI211_X1 U20437 ( .C1(n17461), .C2(n17299), .A(n17298), .B(n17661), .ZN(
        n17307) );
  NAND2_X1 U20438 ( .A1(n17300), .A2(n17694), .ZN(n17671) );
  NOR2_X1 U20439 ( .A1(n17301), .A2(n17671), .ZN(n17302) );
  XNOR2_X1 U20440 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17302), .ZN(
        n17663) );
  OAI21_X1 U20441 ( .B1(n17516), .B2(n17304), .A(n17303), .ZN(n17305) );
  XNOR2_X1 U20442 ( .A(n17305), .B(n17658), .ZN(n17662) );
  OAI22_X1 U20443 ( .A1(n16144), .A2(n17663), .B1(n17508), .B2(n17662), .ZN(
        n17306) );
  AOI211_X1 U20444 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17310), .A(
        n17307), .B(n17306), .ZN(n17308) );
  OAI21_X1 U20445 ( .B1(n17629), .B2(n17667), .A(n17308), .ZN(P3_U2805) );
  INV_X1 U20446 ( .A(n17309), .ZN(n17318) );
  NOR2_X1 U20447 ( .A1(n17861), .A2(n18537), .ZN(n17669) );
  AOI221_X1 U20448 ( .B1(n17311), .B2(n20756), .C1(n17310), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17669), .ZN(n17317) );
  OAI21_X1 U20449 ( .B1(n17313), .B2(n17654), .A(n17312), .ZN(n17670) );
  NOR3_X1 U20450 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17668), .A3(
        n17426), .ZN(n17315) );
  OAI21_X1 U20451 ( .B1(n17685), .B2(n17671), .A(n17452), .ZN(n17332) );
  OAI21_X1 U20452 ( .B1(n17672), .B2(n17685), .A(n17613), .ZN(n17322) );
  AOI21_X1 U20453 ( .B1(n17332), .B2(n17322), .A(n17654), .ZN(n17314) );
  AOI211_X1 U20454 ( .C1(n17535), .C2(n17670), .A(n17315), .B(n17314), .ZN(
        n17316) );
  OAI211_X1 U20455 ( .C1(n17461), .C2(n17318), .A(n17317), .B(n17316), .ZN(
        P3_U2806) );
  OAI22_X1 U20456 ( .A1(n17534), .A2(n17339), .B1(n17319), .B2(n17336), .ZN(
        n17320) );
  NOR2_X1 U20457 ( .A1(n17320), .A2(n17363), .ZN(n17321) );
  XNOR2_X1 U20458 ( .A(n17321), .B(n17685), .ZN(n17689) );
  AOI21_X1 U20459 ( .B1(n17672), .B2(n17685), .A(n17322), .ZN(n17330) );
  AOI21_X1 U20460 ( .B1(n17323), .B2(n18000), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17327) );
  INV_X1 U20461 ( .A(n17365), .ZN(n17325) );
  OAI21_X1 U20462 ( .B1(n17482), .B2(n17325), .A(n17324), .ZN(n17326) );
  NAND2_X1 U20463 ( .A1(n17951), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17690) );
  OAI211_X1 U20464 ( .C1(n17328), .C2(n17327), .A(n17326), .B(n17690), .ZN(
        n17329) );
  AOI211_X1 U20465 ( .C1(n17535), .C2(n17689), .A(n17330), .B(n17329), .ZN(
        n17331) );
  OAI221_X1 U20466 ( .B1(n17332), .B2(n17685), .C1(n17332), .C2(n17671), .A(
        n17331), .ZN(P3_U2807) );
  OAI21_X1 U20467 ( .B1(n17333), .B2(n17624), .A(n17625), .ZN(n17334) );
  AOI21_X1 U20468 ( .B1(n17585), .B2(n17345), .A(n17334), .ZN(n17368) );
  OAI21_X1 U20469 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17365), .A(
        n17368), .ZN(n17353) );
  AOI22_X1 U20470 ( .A1(n17482), .A2(n17335), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17353), .ZN(n17349) );
  INV_X1 U20471 ( .A(n17336), .ZN(n17338) );
  INV_X1 U20472 ( .A(n17397), .ZN(n17741) );
  NAND2_X1 U20473 ( .A1(n17741), .A2(n17337), .ZN(n17701) );
  XNOR2_X1 U20474 ( .A(n17340), .B(n17339), .ZN(n17706) );
  NOR2_X1 U20475 ( .A1(n17426), .A2(n17701), .ZN(n17343) );
  OAI22_X1 U20476 ( .A1(n17693), .A2(n17629), .B1(n17694), .B2(n16144), .ZN(
        n17388) );
  AOI21_X1 U20477 ( .B1(n17341), .B2(n17701), .A(n17388), .ZN(n17362) );
  INV_X1 U20478 ( .A(n17362), .ZN(n17342) );
  MUX2_X1 U20479 ( .A(n17343), .B(n17342), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17344) );
  AOI21_X1 U20480 ( .B1(n17535), .B2(n17706), .A(n17344), .ZN(n17348) );
  NAND2_X1 U20481 ( .A1(n17951), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17707) );
  NOR2_X1 U20482 ( .A1(n17379), .A2(n17345), .ZN(n17355) );
  OAI211_X1 U20483 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17355), .B(n17346), .ZN(n17347) );
  NAND4_X1 U20484 ( .A1(n17349), .A2(n17348), .A3(n17707), .A4(n17347), .ZN(
        P3_U2808) );
  AOI22_X1 U20485 ( .A1(n17951), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n17482), 
        .B2(n17350), .ZN(n17351) );
  INV_X1 U20486 ( .A(n17351), .ZN(n17352) );
  AOI221_X1 U20487 ( .B1(n17355), .B2(n17354), .C1(n17353), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17352), .ZN(n17360) );
  NAND3_X1 U20488 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17534), .A3(
        n17356), .ZN(n17374) );
  INV_X1 U20489 ( .A(n17395), .ZN(n17375) );
  OAI22_X1 U20490 ( .A1(n17700), .A2(n17374), .B1(n17375), .B2(n17357), .ZN(
        n17358) );
  XNOR2_X1 U20491 ( .A(n17361), .B(n17358), .ZN(n17717) );
  NOR2_X1 U20492 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17700), .ZN(
        n17716) );
  NAND2_X1 U20493 ( .A1(n17741), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17714) );
  NOR2_X1 U20494 ( .A1(n17426), .A2(n17714), .ZN(n17386) );
  AOI22_X1 U20495 ( .A1(n17535), .A2(n17717), .B1(n17716), .B2(n17386), .ZN(
        n17359) );
  OAI211_X1 U20496 ( .C1(n17362), .C2(n17361), .A(n17360), .B(n17359), .ZN(
        P3_U2809) );
  INV_X1 U20497 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17730) );
  AOI221_X1 U20498 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17374), 
        .C1(n17730), .C2(n17394), .A(n17363), .ZN(n17364) );
  XNOR2_X1 U20499 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17364), .ZN(
        n17729) );
  AOI21_X1 U20500 ( .B1(n17366), .B2(n18000), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17367) );
  OAI22_X1 U20501 ( .A1(n17368), .A2(n17367), .B1(n17861), .B2(n18530), .ZN(
        n17369) );
  AOI221_X1 U20502 ( .B1(n17482), .B2(n17370), .C1(n17325), .C2(n17370), .A(
        n17369), .ZN(n17373) );
  NOR2_X1 U20503 ( .A1(n17730), .A2(n17714), .ZN(n17721) );
  INV_X1 U20504 ( .A(n17388), .ZN(n17425) );
  OAI21_X1 U20505 ( .B1(n17371), .B2(n17721), .A(n17425), .ZN(n17385) );
  NOR2_X1 U20506 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17730), .ZN(
        n17720) );
  AOI22_X1 U20507 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17385), .B1(
        n17386), .B2(n17720), .ZN(n17372) );
  OAI211_X1 U20508 ( .C1(n17508), .C2(n17729), .A(n17373), .B(n17372), .ZN(
        P3_U2810) );
  OAI21_X1 U20509 ( .B1(n17394), .B2(n17375), .A(n17374), .ZN(n17376) );
  XNOR2_X1 U20510 ( .A(n17376), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17735) );
  AOI21_X1 U20511 ( .B1(n17585), .B2(n17378), .A(n17583), .ZN(n17409) );
  OAI21_X1 U20512 ( .B1(n17377), .B2(n17624), .A(n17409), .ZN(n17391) );
  AOI22_X1 U20513 ( .A1(n17951), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17391), .ZN(n17382) );
  NOR2_X1 U20514 ( .A1(n17379), .A2(n17378), .ZN(n17393) );
  OAI211_X1 U20515 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17393), .B(n17380), .ZN(n17381) );
  OAI211_X1 U20516 ( .C1(n17461), .C2(n17383), .A(n17382), .B(n17381), .ZN(
        n17384) );
  AOI221_X1 U20517 ( .B1(n17386), .B2(n17730), .C1(n17385), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17384), .ZN(n17387) );
  OAI21_X1 U20518 ( .B1(n17735), .B2(n17508), .A(n17387), .ZN(P3_U2811) );
  AOI21_X1 U20519 ( .B1(n17406), .B2(n17397), .A(n17388), .ZN(n17404) );
  OAI22_X1 U20520 ( .A1(n17861), .A2(n18525), .B1(n17461), .B2(n17389), .ZN(
        n17390) );
  AOI221_X1 U20521 ( .B1(n17393), .B2(n17392), .C1(n17391), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17390), .ZN(n17399) );
  OAI21_X1 U20522 ( .B1(n17400), .B2(n17516), .A(n17394), .ZN(n17396) );
  XNOR2_X1 U20523 ( .A(n17396), .B(n17395), .ZN(n17747) );
  NOR2_X1 U20524 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17397), .ZN(
        n17746) );
  AOI22_X1 U20525 ( .A1(n17535), .A2(n17747), .B1(n17406), .B2(n17746), .ZN(
        n17398) );
  OAI211_X1 U20526 ( .C1(n17404), .C2(n17400), .A(n17399), .B(n17398), .ZN(
        P3_U2812) );
  AOI21_X1 U20527 ( .B1(n17401), .B2(n18000), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17410) );
  AOI22_X1 U20528 ( .A1(n17951), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n17402), 
        .B2(n17616), .ZN(n17408) );
  NOR2_X1 U20529 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17761), .ZN(
        n17750) );
  AOI21_X1 U20530 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17403), .A(
        n9721), .ZN(n17754) );
  OAI22_X1 U20531 ( .A1(n17404), .A2(n9937), .B1(n17754), .B2(n17508), .ZN(
        n17405) );
  AOI21_X1 U20532 ( .B1(n17406), .B2(n17750), .A(n17405), .ZN(n17407) );
  OAI211_X1 U20533 ( .C1(n17410), .C2(n17409), .A(n17408), .B(n17407), .ZN(
        P3_U2813) );
  AND2_X1 U20534 ( .A1(n17534), .A2(n9640), .ZN(n17515) );
  AOI22_X1 U20535 ( .A1(n17515), .A2(n17412), .B1(n17411), .B2(n17516), .ZN(
        n17413) );
  XNOR2_X1 U20536 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17413), .ZN(
        n17763) );
  AOI21_X1 U20537 ( .B1(n17585), .B2(n17414), .A(n17583), .ZN(n17442) );
  OAI21_X1 U20538 ( .B1(n17415), .B2(n17624), .A(n17442), .ZN(n17434) );
  AOI22_X1 U20539 ( .A1(n17951), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17434), .ZN(n17421) );
  INV_X1 U20540 ( .A(n17416), .ZN(n17418) );
  NAND2_X1 U20541 ( .A1(n17457), .A2(n17417), .ZN(n17475) );
  NOR2_X1 U20542 ( .A1(n17418), .A2(n17475), .ZN(n17436) );
  OAI211_X1 U20543 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17436), .B(n17419), .ZN(n17420) );
  OAI211_X1 U20544 ( .C1(n17461), .C2(n17422), .A(n17421), .B(n17420), .ZN(
        n17423) );
  AOI21_X1 U20545 ( .B1(n17535), .B2(n17763), .A(n17423), .ZN(n17424) );
  OAI221_X1 U20546 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17426), 
        .C1(n17761), .C2(n17425), .A(n17424), .ZN(P3_U2814) );
  NOR2_X1 U20547 ( .A1(n17786), .A2(n17789), .ZN(n17429) );
  NOR2_X1 U20548 ( .A1(n17815), .A2(n17427), .ZN(n17463) );
  INV_X1 U20549 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n20633) );
  NAND3_X1 U20550 ( .A1(n17517), .A2(n20633), .A3(n17516), .ZN(n17494) );
  NOR2_X1 U20551 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17494), .ZN(
        n17428) );
  INV_X1 U20552 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17808) );
  NAND2_X1 U20553 ( .A1(n17428), .A2(n17808), .ZN(n17469) );
  NOR2_X1 U20554 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17469), .ZN(
        n17448) );
  AOI21_X1 U20555 ( .B1(n17429), .B2(n17463), .A(n17448), .ZN(n17430) );
  AOI221_X1 U20556 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17814), 
        .C1(n17516), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17430), .ZN(
        n17431) );
  XNOR2_X1 U20557 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17431), .ZN(
        n17774) );
  INV_X1 U20558 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17435) );
  OAI22_X1 U20559 ( .A1(n17861), .A2(n18519), .B1(n17461), .B2(n17432), .ZN(
        n17433) );
  AOI221_X1 U20560 ( .B1(n17436), .B2(n17435), .C1(n17434), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17433), .ZN(n17440) );
  NOR2_X1 U20561 ( .A1(n17694), .A2(n16144), .ZN(n17438) );
  NAND2_X1 U20562 ( .A1(n17767), .A2(n17446), .ZN(n17771) );
  NOR2_X1 U20563 ( .A1(n17693), .A2(n17629), .ZN(n17437) );
  NAND2_X1 U20564 ( .A1(n17441), .A2(n17767), .ZN(n17769) );
  AOI22_X1 U20565 ( .A1(n17438), .A2(n17771), .B1(n17437), .B2(n17769), .ZN(
        n17439) );
  OAI211_X1 U20566 ( .C1(n17508), .C2(n17774), .A(n17440), .B(n17439), .ZN(
        P3_U2815) );
  OAI221_X1 U20567 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17807), .A(n17441), .ZN(
        n17797) );
  NOR2_X1 U20568 ( .A1(n17861), .A2(n18517), .ZN(n17791) );
  NAND2_X1 U20569 ( .A1(n17457), .A2(n18000), .ZN(n17487) );
  AOI221_X1 U20570 ( .B1(n17458), .B2(n17443), .C1(n17487), .C2(n17443), .A(
        n17442), .ZN(n17444) );
  AOI211_X1 U20571 ( .C1(n17445), .C2(n17616), .A(n17791), .B(n17444), .ZN(
        n17451) );
  NAND2_X1 U20572 ( .A1(n17780), .A2(n9640), .ZN(n17804) );
  INV_X1 U20573 ( .A(n17446), .ZN(n17447) );
  AOI221_X1 U20574 ( .B1(n17786), .B2(n17789), .C1(n17804), .C2(n17789), .A(
        n17447), .ZN(n17793) );
  AOI22_X1 U20575 ( .A1(n17515), .A2(n17784), .B1(n17448), .B2(n17814), .ZN(
        n17449) );
  XNOR2_X1 U20576 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17449), .ZN(
        n17792) );
  AOI22_X1 U20577 ( .A1(n17452), .A2(n17793), .B1(n17535), .B2(n17792), .ZN(
        n17450) );
  OAI211_X1 U20578 ( .C1(n17629), .C2(n17797), .A(n17451), .B(n17450), .ZN(
        P3_U2816) );
  AOI22_X1 U20579 ( .A1(n17613), .A2(n17453), .B1(n17452), .B2(n17804), .ZN(
        n17476) );
  AOI21_X1 U20580 ( .B1(n17455), .B2(n17454), .A(n17583), .ZN(n17456) );
  OAI21_X1 U20581 ( .B1(n17457), .B2(n17523), .A(n17456), .ZN(n17471) );
  NOR2_X1 U20582 ( .A1(n17861), .A2(n18515), .ZN(n17799) );
  OAI21_X1 U20583 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17458), .ZN(n17459) );
  OAI22_X1 U20584 ( .A1(n17461), .A2(n17460), .B1(n17475), .B2(n17459), .ZN(
        n17462) );
  AOI211_X1 U20585 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17471), .A(
        n17799), .B(n17462), .ZN(n17468) );
  NOR2_X1 U20586 ( .A1(n17814), .A2(n17516), .ZN(n17465) );
  INV_X1 U20587 ( .A(n17469), .ZN(n17464) );
  OAI22_X1 U20588 ( .A1(n17465), .A2(n17464), .B1(n17463), .B2(n17814), .ZN(
        n17466) );
  XNOR2_X1 U20589 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17466), .ZN(
        n17800) );
  NOR2_X1 U20590 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17782), .ZN(
        n17798) );
  AOI22_X1 U20591 ( .A1(n17535), .A2(n17800), .B1(n17798), .B2(n17499), .ZN(
        n17467) );
  OAI211_X1 U20592 ( .C1(n17476), .C2(n17786), .A(n17468), .B(n17467), .ZN(
        P3_U2817) );
  NAND3_X1 U20593 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n17515), .ZN(n17489) );
  OAI21_X1 U20594 ( .B1(n17808), .B2(n17489), .A(n17469), .ZN(n17470) );
  XNOR2_X1 U20595 ( .A(n17470), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17821) );
  INV_X1 U20596 ( .A(n17471), .ZN(n17473) );
  NAND2_X1 U20597 ( .A1(n17951), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n17472) );
  OAI221_X1 U20598 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17475), .C1(
        n17474), .C2(n17473), .A(n17472), .ZN(n17480) );
  NOR2_X1 U20599 ( .A1(n17522), .A2(n17815), .ZN(n17478) );
  INV_X1 U20600 ( .A(n17476), .ZN(n17477) );
  MUX2_X1 U20601 ( .A(n17478), .B(n17477), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n17479) );
  AOI211_X1 U20602 ( .C1(n17482), .C2(n17481), .A(n17480), .B(n17479), .ZN(
        n17483) );
  OAI21_X1 U20603 ( .B1(n17821), .B2(n17508), .A(n17483), .ZN(P3_U2818) );
  NOR3_X1 U20604 ( .A1(n20794), .A2(n17484), .A3(n18302), .ZN(n17540) );
  NAND3_X1 U20605 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(n17540), .ZN(n17511) );
  NOR2_X1 U20606 ( .A1(n17510), .A2(n17511), .ZN(n17509) );
  NAND2_X1 U20607 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17509), .ZN(
        n17506) );
  OAI21_X1 U20608 ( .B1(n17621), .B2(n17485), .A(n17506), .ZN(n17486) );
  AOI22_X1 U20609 ( .A1(n17488), .A2(n17616), .B1(n17487), .B2(n17486), .ZN(
        n17493) );
  OAI21_X1 U20610 ( .B1(n17494), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17489), .ZN(n17490) );
  XNOR2_X1 U20611 ( .A(n17490), .B(n17808), .ZN(n17822) );
  NAND2_X1 U20612 ( .A1(n17801), .A2(n17808), .ZN(n17836) );
  OAI22_X1 U20613 ( .A1(n9640), .A2(n16144), .B1(n17629), .B2(n17823), .ZN(
        n17519) );
  AOI21_X1 U20614 ( .B1(n17831), .B2(n17499), .A(n17519), .ZN(n17502) );
  OAI22_X1 U20615 ( .A1(n17522), .A2(n17836), .B1(n17502), .B2(n17808), .ZN(
        n17491) );
  AOI21_X1 U20616 ( .B1(n17535), .B2(n17822), .A(n17491), .ZN(n17492) );
  OAI211_X1 U20617 ( .C1(n17861), .C2(n18511), .A(n17493), .B(n17492), .ZN(
        P3_U2819) );
  NAND2_X1 U20618 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17515), .ZN(
        n17495) );
  NAND2_X1 U20619 ( .A1(n17495), .A2(n17494), .ZN(n17496) );
  XNOR2_X1 U20620 ( .A(n17496), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17846) );
  INV_X1 U20621 ( .A(n17509), .ZN(n17497) );
  OAI21_X1 U20622 ( .B1(n17621), .B2(n17498), .A(n17497), .ZN(n17505) );
  INV_X1 U20623 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18509) );
  NOR2_X1 U20624 ( .A1(n17861), .A2(n18509), .ZN(n17504) );
  AOI21_X1 U20625 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17499), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17501) );
  OAI22_X1 U20626 ( .A1(n17502), .A2(n17501), .B1(n17608), .B2(n17500), .ZN(
        n17503) );
  AOI211_X1 U20627 ( .C1(n17506), .C2(n17505), .A(n17504), .B(n17503), .ZN(
        n17507) );
  OAI21_X1 U20628 ( .B1(n17846), .B2(n17508), .A(n17507), .ZN(P3_U2820) );
  AOI211_X1 U20629 ( .C1(n17511), .C2(n17510), .A(n17621), .B(n17509), .ZN(
        n17513) );
  NOR2_X1 U20630 ( .A1(n17861), .A2(n18508), .ZN(n17512) );
  AOI211_X1 U20631 ( .C1(n17514), .C2(n17616), .A(n17513), .B(n17512), .ZN(
        n17521) );
  AOI21_X1 U20632 ( .B1(n17517), .B2(n17516), .A(n17515), .ZN(n17518) );
  XNOR2_X1 U20633 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n17518), .ZN(
        n17854) );
  AOI22_X1 U20634 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17519), .B1(
        n17535), .B2(n17854), .ZN(n17520) );
  OAI211_X1 U20635 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n17522), .A(
        n17521), .B(n17520), .ZN(P3_U2821) );
  INV_X1 U20636 ( .A(n17533), .ZN(n17875) );
  OAI21_X1 U20637 ( .B1(n17524), .B2(n17523), .A(n17625), .ZN(n17538) );
  AOI221_X1 U20638 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C1(n17526), .C2(n17525), .A(n18302), .ZN(n17529) );
  OAI22_X1 U20639 ( .A1(n17608), .A2(n17527), .B1(n17861), .B2(n18507), .ZN(
        n17528) );
  AOI211_X1 U20640 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17538), .A(
        n17529), .B(n17528), .ZN(n17537) );
  AOI21_X1 U20641 ( .B1(n17531), .B2(n17862), .A(n17530), .ZN(n17871) );
  OAI21_X1 U20642 ( .B1(n17534), .B2(n17533), .A(n17532), .ZN(n17869) );
  AOI22_X1 U20643 ( .A1(n17613), .A2(n17871), .B1(n17535), .B2(n17869), .ZN(
        n17536) );
  OAI211_X1 U20644 ( .C1(n16144), .C2(n17875), .A(n17537), .B(n17536), .ZN(
        P3_U2822) );
  INV_X1 U20645 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17539) );
  NOR2_X1 U20646 ( .A1(n17861), .A2(n18504), .ZN(n17878) );
  AOI221_X1 U20647 ( .B1(n17540), .B2(n17539), .C1(n17538), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n17878), .ZN(n17547) );
  NAND2_X1 U20648 ( .A1(n17542), .A2(n17541), .ZN(n17543) );
  XNOR2_X1 U20649 ( .A(n17543), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17880) );
  AOI21_X1 U20650 ( .B1(n17885), .B2(n17545), .A(n17544), .ZN(n17881) );
  AOI22_X1 U20651 ( .A1(n17613), .A2(n17880), .B1(n17617), .B2(n17881), .ZN(
        n17546) );
  OAI211_X1 U20652 ( .C1(n17608), .C2(n17548), .A(n17547), .B(n17546), .ZN(
        P3_U2823) );
  AOI21_X1 U20653 ( .B1(n17552), .B2(n18000), .A(n17621), .ZN(n17549) );
  INV_X1 U20654 ( .A(n17549), .ZN(n17572) );
  AOI21_X1 U20655 ( .B1(n17876), .B2(n17551), .A(n17550), .ZN(n17888) );
  NAND2_X1 U20656 ( .A1(n17552), .A2(n18000), .ZN(n17553) );
  OAI22_X1 U20657 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17553), .B1(
        n17861), .B2(n20788), .ZN(n17554) );
  AOI21_X1 U20658 ( .B1(n17613), .B2(n17888), .A(n17554), .ZN(n17560) );
  AOI21_X1 U20659 ( .B1(n17557), .B2(n17556), .A(n17555), .ZN(n17889) );
  AOI22_X1 U20660 ( .A1(n17617), .A2(n17889), .B1(n17558), .B2(n17616), .ZN(
        n17559) );
  OAI211_X1 U20661 ( .C1(n20794), .C2(n17572), .A(n17560), .B(n17559), .ZN(
        P3_U2824) );
  AOI21_X1 U20662 ( .B1(n17561), .B2(n17625), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17573) );
  AOI21_X1 U20663 ( .B1(n17564), .B2(n17563), .A(n17562), .ZN(n17893) );
  AOI22_X1 U20664 ( .A1(n17613), .A2(n17893), .B1(n17951), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17571) );
  OAI21_X1 U20665 ( .B1(n17567), .B2(n17566), .A(n17565), .ZN(n17568) );
  XNOR2_X1 U20666 ( .A(n17568), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17894) );
  AOI22_X1 U20667 ( .A1(n17617), .A2(n17894), .B1(n17569), .B2(n17616), .ZN(
        n17570) );
  OAI211_X1 U20668 ( .C1(n17573), .C2(n17572), .A(n17571), .B(n17570), .ZN(
        P3_U2825) );
  OAI21_X1 U20669 ( .B1(n17576), .B2(n17575), .A(n17574), .ZN(n17578) );
  XNOR2_X1 U20670 ( .A(n17578), .B(n17577), .ZN(n17913) );
  AOI22_X1 U20671 ( .A1(n17951), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18000), 
        .B2(n17579), .ZN(n17590) );
  AOI21_X1 U20672 ( .B1(n17582), .B2(n17581), .A(n17580), .ZN(n17910) );
  AOI21_X1 U20673 ( .B1(n17585), .B2(n17584), .A(n17583), .ZN(n17601) );
  OAI22_X1 U20674 ( .A1(n17608), .A2(n17587), .B1(n17601), .B2(n17586), .ZN(
        n17588) );
  AOI21_X1 U20675 ( .B1(n17617), .B2(n17910), .A(n17588), .ZN(n17589) );
  OAI211_X1 U20676 ( .C1(n17629), .C2(n17913), .A(n17590), .B(n17589), .ZN(
        P3_U2826) );
  AOI21_X1 U20677 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17625), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17600) );
  AOI21_X1 U20678 ( .B1(n17593), .B2(n17592), .A(n17591), .ZN(n17916) );
  AOI22_X1 U20679 ( .A1(n17613), .A2(n17916), .B1(n17951), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17599) );
  AOI21_X1 U20680 ( .B1(n17596), .B2(n17595), .A(n17594), .ZN(n17917) );
  AOI22_X1 U20681 ( .A1(n17617), .A2(n17917), .B1(n17597), .B2(n17616), .ZN(
        n17598) );
  OAI211_X1 U20682 ( .C1(n17601), .C2(n17600), .A(n17599), .B(n17598), .ZN(
        P3_U2827) );
  INV_X1 U20683 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17611) );
  AOI21_X1 U20684 ( .B1(n17604), .B2(n17603), .A(n17602), .ZN(n17934) );
  NOR2_X1 U20685 ( .A1(n17861), .A2(n18495), .ZN(n17935) );
  XNOR2_X1 U20686 ( .A(n17606), .B(n17605), .ZN(n17922) );
  OAI22_X1 U20687 ( .A1(n17608), .A2(n17607), .B1(n17628), .B2(n17922), .ZN(
        n17609) );
  AOI211_X1 U20688 ( .C1(n17613), .C2(n17934), .A(n17935), .B(n17609), .ZN(
        n17610) );
  OAI221_X1 U20689 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18302), .C1(
        n17611), .C2(n17625), .A(n17610), .ZN(P3_U2828) );
  NOR2_X1 U20690 ( .A1(n17623), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17612) );
  XNOR2_X1 U20691 ( .A(n17612), .B(n17615), .ZN(n17946) );
  AOI22_X1 U20692 ( .A1(n17613), .A2(n17946), .B1(n17951), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17619) );
  AOI21_X1 U20693 ( .B1(n17615), .B2(n17622), .A(n17614), .ZN(n17940) );
  AOI22_X1 U20694 ( .A1(n17617), .A2(n17940), .B1(n17620), .B2(n17616), .ZN(
        n17618) );
  OAI211_X1 U20695 ( .C1(n17621), .C2(n17620), .A(n17619), .B(n17618), .ZN(
        P3_U2829) );
  OAI21_X1 U20696 ( .B1(n17623), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17622), .ZN(n17956) );
  INV_X1 U20697 ( .A(n17956), .ZN(n17954) );
  NAND3_X1 U20698 ( .A1(n18577), .A2(n17625), .A3(n17624), .ZN(n17626) );
  AOI22_X1 U20699 ( .A1(n17951), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17626), .ZN(n17627) );
  OAI221_X1 U20700 ( .B1(n17954), .B2(n17629), .C1(n17956), .C2(n17628), .A(
        n17627), .ZN(P3_U2830) );
  INV_X1 U20701 ( .A(n17645), .ZN(n17692) );
  NOR2_X1 U20702 ( .A1(n17692), .A2(n17630), .ZN(n17639) );
  AOI21_X1 U20703 ( .B1(n17848), .B2(n17648), .A(n17631), .ZN(n17636) );
  AOI22_X1 U20704 ( .A1(n18428), .A2(n17633), .B1(n17805), .B2(n17632), .ZN(
        n17635) );
  NAND2_X1 U20705 ( .A1(n17848), .A2(n18595), .ZN(n17926) );
  NAND2_X1 U20706 ( .A1(n17697), .A2(n17926), .ZN(n17737) );
  INV_X1 U20707 ( .A(n18399), .ZN(n17900) );
  OAI21_X1 U20708 ( .B1(n17737), .B2(n17634), .A(n17900), .ZN(n17655) );
  NAND3_X1 U20709 ( .A1(n17636), .A2(n17635), .A3(n17655), .ZN(n17647) );
  AOI21_X1 U20710 ( .B1(n17648), .B2(n18411), .A(n17647), .ZN(n17637) );
  INV_X1 U20711 ( .A(n17637), .ZN(n17638) );
  MUX2_X1 U20712 ( .A(n17639), .B(n17638), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n17640) );
  AOI22_X1 U20713 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17936), .B1(
        n17952), .B2(n17640), .ZN(n17642) );
  OAI211_X1 U20714 ( .C1(n17643), .C2(n17845), .A(n17642), .B(n17641), .ZN(
        P3_U2835) );
  AOI22_X1 U20715 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17936), .B1(
        n17951), .B2(P3_REIP_REG_26__SCAN_IN), .ZN(n17651) );
  INV_X1 U20716 ( .A(n17644), .ZN(n17646) );
  INV_X1 U20717 ( .A(n17701), .ZN(n17698) );
  NAND3_X1 U20718 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17698), .A3(
        n17645), .ZN(n17686) );
  NOR2_X1 U20719 ( .A1(n17646), .A2(n17686), .ZN(n17649) );
  OAI221_X1 U20720 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17649), 
        .C1(n17648), .C2(n17647), .A(n17952), .ZN(n17650) );
  OAI211_X1 U20721 ( .C1(n17652), .C2(n17845), .A(n17651), .B(n17650), .ZN(
        P3_U2836) );
  NOR3_X1 U20722 ( .A1(n17653), .A2(n17668), .A3(n17654), .ZN(n17659) );
  NOR2_X1 U20723 ( .A1(n17654), .A2(n17668), .ZN(n17656) );
  OAI221_X1 U20724 ( .B1(n18406), .B2(n17678), .C1(n18406), .C2(n17656), .A(
        n17655), .ZN(n17657) );
  OAI221_X1 U20725 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17659), 
        .C1(n17658), .C2(n17657), .A(n17952), .ZN(n17660) );
  NAND2_X1 U20726 ( .A1(n17661), .A2(n17660), .ZN(n17665) );
  OAI22_X1 U20727 ( .A1(n17874), .A2(n17663), .B1(n17845), .B2(n17662), .ZN(
        n17664) );
  AOI211_X1 U20728 ( .C1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n17936), .A(
        n17665), .B(n17664), .ZN(n17666) );
  OAI21_X1 U20729 ( .B1(n17914), .B2(n17667), .A(n17666), .ZN(P3_U2837) );
  OR2_X1 U20730 ( .A1(n17668), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17684) );
  AOI21_X1 U20731 ( .B1(n17870), .B2(n17670), .A(n17669), .ZN(n17683) );
  NOR2_X1 U20732 ( .A1(n17685), .A2(n17671), .ZN(n17677) );
  OR2_X1 U20733 ( .A1(n17672), .A2(n17685), .ZN(n17673) );
  AOI21_X1 U20734 ( .B1(n18428), .B2(n17673), .A(n17936), .ZN(n17676) );
  OAI21_X1 U20735 ( .B1(n17674), .B2(n17737), .A(n17900), .ZN(n17675) );
  OAI211_X1 U20736 ( .C1(n17677), .C2(n17825), .A(n17676), .B(n17675), .ZN(
        n17681) );
  NAND2_X1 U20737 ( .A1(n17741), .A2(n17678), .ZN(n17736) );
  AOI221_X1 U20738 ( .B1(n17679), .B2(n18438), .C1(n17736), .C2(n18438), .A(
        n17681), .ZN(n17680) );
  AOI21_X1 U20739 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17680), .A(
        n17951), .ZN(n17688) );
  OAI211_X1 U20740 ( .C1(n17899), .C2(n17681), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17688), .ZN(n17682) );
  OAI211_X1 U20741 ( .C1(n17684), .C2(n17715), .A(n17683), .B(n17682), .ZN(
        P3_U2838) );
  OAI21_X1 U20742 ( .B1(n17936), .B2(n17686), .A(n17685), .ZN(n17687) );
  AOI22_X1 U20743 ( .A1(n17870), .A2(n17689), .B1(n17688), .B2(n17687), .ZN(
        n17691) );
  NAND2_X1 U20744 ( .A1(n17691), .A2(n17690), .ZN(P3_U2839) );
  NOR2_X1 U20745 ( .A1(n17692), .A2(n17701), .ZN(n17705) );
  INV_X1 U20746 ( .A(n18428), .ZN(n17824) );
  NOR2_X1 U20747 ( .A1(n17693), .A2(n17824), .ZN(n17768) );
  NOR2_X1 U20748 ( .A1(n17694), .A2(n17825), .ZN(n17770) );
  NOR2_X1 U20749 ( .A1(n17768), .A2(n17770), .ZN(n17710) );
  OAI21_X1 U20750 ( .B1(n17695), .B2(n17714), .A(n18438), .ZN(n17696) );
  OAI221_X1 U20751 ( .B1(n18400), .B2(n17697), .C1(n18400), .C2(n17721), .A(
        n17696), .ZN(n17722) );
  NOR2_X1 U20752 ( .A1(n18428), .A2(n17805), .ZN(n17740) );
  OAI22_X1 U20753 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18400), .B1(
        n17698), .B2(n17740), .ZN(n17699) );
  NOR2_X1 U20754 ( .A1(n17722), .A2(n17699), .ZN(n17711) );
  OAI211_X1 U20755 ( .C1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n17841), .A(
        n17710), .B(n17711), .ZN(n17704) );
  INV_X1 U20756 ( .A(n17700), .ZN(n17712) );
  OAI21_X1 U20757 ( .B1(n17757), .B2(n17701), .A(n17848), .ZN(n17702) );
  OAI211_X1 U20758 ( .C1(n17712), .C2(n18406), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17702), .ZN(n17703) );
  OAI22_X1 U20759 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17705), .B1(
        n17704), .B2(n17703), .ZN(n17709) );
  AOI22_X1 U20760 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17936), .B1(
        n17870), .B2(n17706), .ZN(n17708) );
  OAI211_X1 U20761 ( .C1(n17938), .C2(n17709), .A(n17708), .B(n17707), .ZN(
        P3_U2840) );
  NOR2_X1 U20762 ( .A1(n18438), .A2(n17848), .ZN(n17779) );
  NAND2_X1 U20763 ( .A1(n17952), .A2(n17710), .ZN(n17760) );
  AOI221_X1 U20764 ( .B1(n17757), .B2(n17848), .C1(n17714), .C2(n17848), .A(
        n17760), .ZN(n17725) );
  OAI211_X1 U20765 ( .C1(n17712), .C2(n17779), .A(n17725), .B(n17711), .ZN(
        n17713) );
  NAND2_X1 U20766 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17713), .ZN(
        n17719) );
  NOR2_X1 U20767 ( .A1(n17715), .A2(n17714), .ZN(n17731) );
  AOI22_X1 U20768 ( .A1(n17870), .A2(n17717), .B1(n17716), .B2(n17731), .ZN(
        n17718) );
  OAI221_X1 U20769 ( .B1(n17951), .B2(n17719), .C1(n17861), .C2(n18531), .A(
        n17718), .ZN(P3_U2841) );
  AOI22_X1 U20770 ( .A1(n17951), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n17731), 
        .B2(n17720), .ZN(n17728) );
  INV_X1 U20771 ( .A(n17721), .ZN(n17723) );
  INV_X1 U20772 ( .A(n17740), .ZN(n17830) );
  AOI21_X1 U20773 ( .B1(n17723), .B2(n17830), .A(n17722), .ZN(n17724) );
  AOI21_X1 U20774 ( .B1(n17725), .B2(n17724), .A(n17951), .ZN(n17732) );
  NOR3_X1 U20775 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17779), .A3(
        n18468), .ZN(n17726) );
  OAI21_X1 U20776 ( .B1(n17732), .B2(n17726), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17727) );
  OAI211_X1 U20777 ( .C1(n17729), .C2(n17845), .A(n17728), .B(n17727), .ZN(
        P3_U2842) );
  AOI22_X1 U20778 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17732), .B1(
        n17731), .B2(n17730), .ZN(n17734) );
  NAND2_X1 U20779 ( .A1(n17951), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17733) );
  OAI211_X1 U20780 ( .C1(n17735), .C2(n17845), .A(n17734), .B(n17733), .ZN(
        P3_U2843) );
  AOI21_X1 U20781 ( .B1(n18438), .B2(n17736), .A(n17760), .ZN(n17739) );
  OAI21_X1 U20782 ( .B1(n17761), .B2(n17737), .A(n17900), .ZN(n17738) );
  OAI211_X1 U20783 ( .C1(n17741), .C2(n17740), .A(n17739), .B(n17738), .ZN(
        n17751) );
  OAI221_X1 U20784 ( .B1(n17751), .B2(n17900), .C1(n17751), .C2(n9937), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17749) );
  INV_X1 U20785 ( .A(n17901), .ZN(n17756) );
  AOI22_X1 U20786 ( .A1(n18438), .A2(n17923), .B1(n17756), .B2(n17924), .ZN(
        n17864) );
  NOR2_X1 U20787 ( .A1(n17864), .A2(n17742), .ZN(n17766) );
  INV_X1 U20788 ( .A(n17743), .ZN(n17744) );
  NOR2_X1 U20789 ( .A1(n17745), .A2(n17857), .ZN(n17762) );
  AOI22_X1 U20790 ( .A1(n17870), .A2(n17747), .B1(n17746), .B2(n17762), .ZN(
        n17748) );
  OAI221_X1 U20791 ( .B1(n17951), .B2(n17749), .C1(n17861), .C2(n18525), .A(
        n17748), .ZN(P3_U2844) );
  AOI22_X1 U20792 ( .A1(n17951), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n17762), 
        .B2(n17750), .ZN(n17753) );
  NAND3_X1 U20793 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17861), .A3(
        n17751), .ZN(n17752) );
  OAI211_X1 U20794 ( .C1(n17754), .C2(n17845), .A(n17753), .B(n17752), .ZN(
        P3_U2845) );
  INV_X1 U20795 ( .A(n17755), .ZN(n17866) );
  NAND2_X1 U20796 ( .A1(n17865), .A2(n17756), .ZN(n17858) );
  AND2_X1 U20797 ( .A1(n17781), .A2(n18438), .ZN(n17829) );
  AOI221_X1 U20798 ( .B1(n17866), .B2(n18411), .C1(n17858), .C2(n18411), .A(
        n17829), .ZN(n17850) );
  NOR2_X1 U20799 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18400), .ZN(
        n17849) );
  AOI211_X1 U20800 ( .C1(n17757), .C2(n17848), .A(n17767), .B(n17849), .ZN(
        n17758) );
  OAI211_X1 U20801 ( .C1(n17759), .C2(n17841), .A(n17850), .B(n17758), .ZN(
        n17772) );
  OAI221_X1 U20802 ( .B1(n17760), .B2(n17899), .C1(n17760), .C2(n17772), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17765) );
  AOI22_X1 U20803 ( .A1(n17870), .A2(n17763), .B1(n17762), .B2(n17761), .ZN(
        n17764) );
  OAI221_X1 U20804 ( .B1(n17951), .B2(n17765), .C1(n17861), .C2(n18521), .A(
        n17764), .ZN(P3_U2846) );
  NAND2_X1 U20805 ( .A1(n17784), .A2(n17766), .ZN(n17788) );
  OAI21_X1 U20806 ( .B1(n17789), .B2(n17788), .A(n17767), .ZN(n17773) );
  AOI222_X1 U20807 ( .A1(n17773), .A2(n17772), .B1(n17771), .B2(n17770), .C1(
        n17769), .C2(n17768), .ZN(n17778) );
  INV_X1 U20808 ( .A(n17774), .ZN(n17775) );
  AOI22_X1 U20809 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17936), .B1(
        n17870), .B2(n17775), .ZN(n17777) );
  NAND2_X1 U20810 ( .A1(n17951), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n17776) );
  OAI211_X1 U20811 ( .C1(n17778), .C2(n17938), .A(n17777), .B(n17776), .ZN(
        P3_U2847) );
  INV_X1 U20812 ( .A(n17779), .ZN(n17941) );
  INV_X1 U20813 ( .A(n17847), .ZN(n17827) );
  AOI21_X1 U20814 ( .B1(n17780), .B2(n17827), .A(n18409), .ZN(n17803) );
  AOI221_X1 U20815 ( .B1(n17782), .B2(n18438), .C1(n17781), .C2(n18438), .A(
        n17789), .ZN(n17783) );
  OAI221_X1 U20816 ( .B1(n18400), .B2(n17784), .C1(n18400), .C2(n17838), .A(
        n17783), .ZN(n17785) );
  AOI211_X1 U20817 ( .C1(n17786), .C2(n17941), .A(n17803), .B(n17785), .ZN(
        n17787) );
  AOI211_X1 U20818 ( .C1(n17789), .C2(n17788), .A(n17787), .B(n17938), .ZN(
        n17790) );
  AOI211_X1 U20819 ( .C1(n17936), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17791), .B(n17790), .ZN(n17796) );
  AOI22_X1 U20820 ( .A1(n17794), .A2(n17793), .B1(n17870), .B2(n17792), .ZN(
        n17795) );
  OAI211_X1 U20821 ( .C1(n17914), .C2(n17797), .A(n17796), .B(n17795), .ZN(
        P3_U2848) );
  INV_X1 U20822 ( .A(n17798), .ZN(n17812) );
  AOI21_X1 U20823 ( .B1(n17800), .B2(n17870), .A(n17799), .ZN(n17811) );
  AOI21_X1 U20824 ( .B1(n17838), .B2(n17801), .A(n18400), .ZN(n17802) );
  AOI21_X1 U20825 ( .B1(n18438), .B2(n17815), .A(n17802), .ZN(n17832) );
  AOI211_X1 U20826 ( .C1(n17805), .C2(n17804), .A(n17829), .B(n17803), .ZN(
        n17806) );
  OAI211_X1 U20827 ( .C1(n17807), .C2(n17824), .A(n17832), .B(n17806), .ZN(
        n17817) );
  AOI21_X1 U20828 ( .B1(n17808), .B2(n18411), .A(n17814), .ZN(n17813) );
  OAI21_X1 U20829 ( .B1(n17841), .B2(n17813), .A(n17952), .ZN(n17809) );
  OAI211_X1 U20830 ( .C1(n17817), .C2(n17809), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17861), .ZN(n17810) );
  OAI211_X1 U20831 ( .C1(n17812), .C2(n17857), .A(n17811), .B(n17810), .ZN(
        P3_U2849) );
  AOI22_X1 U20832 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17936), .B1(
        n17951), .B2(P3_REIP_REG_12__SCAN_IN), .ZN(n17820) );
  INV_X1 U20833 ( .A(n17813), .ZN(n17818) );
  OAI22_X1 U20834 ( .A1(n17815), .A2(n17857), .B1(n17814), .B2(n17938), .ZN(
        n17816) );
  OAI21_X1 U20835 ( .B1(n17818), .B2(n17817), .A(n17816), .ZN(n17819) );
  OAI211_X1 U20836 ( .C1(n17821), .C2(n17845), .A(n17820), .B(n17819), .ZN(
        P3_U2850) );
  AOI22_X1 U20837 ( .A1(n17951), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17870), 
        .B2(n17822), .ZN(n17835) );
  OAI22_X1 U20838 ( .A1(n9640), .A2(n17825), .B1(n17824), .B2(n17823), .ZN(
        n17826) );
  NOR2_X1 U20839 ( .A1(n17938), .A2(n17826), .ZN(n17851) );
  OAI221_X1 U20840 ( .B1(n18409), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n18409), .C2(n17827), .A(n17851), .ZN(n17828) );
  AOI211_X1 U20841 ( .C1(n17831), .C2(n17830), .A(n17829), .B(n17828), .ZN(
        n17840) );
  OAI211_X1 U20842 ( .C1(n18409), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17832), .B(n17840), .ZN(n17833) );
  NAND3_X1 U20843 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17861), .A3(
        n17833), .ZN(n17834) );
  OAI211_X1 U20844 ( .C1(n17857), .C2(n17836), .A(n17835), .B(n17834), .ZN(
        P3_U2851) );
  NOR3_X1 U20845 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n20633), .A3(
        n17857), .ZN(n17837) );
  AOI21_X1 U20846 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n17951), .A(n17837), 
        .ZN(n17844) );
  OR2_X1 U20847 ( .A1(n17838), .A2(n18400), .ZN(n17839) );
  OAI211_X1 U20848 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n17841), .A(
        n17840), .B(n17839), .ZN(n17842) );
  NAND3_X1 U20849 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17861), .A3(
        n17842), .ZN(n17843) );
  OAI211_X1 U20850 ( .C1(n17846), .C2(n17845), .A(n17844), .B(n17843), .ZN(
        P3_U2852) );
  OAI21_X1 U20851 ( .B1(n17849), .B2(n17848), .A(n17847), .ZN(n17852) );
  NAND3_X1 U20852 ( .A1(n17852), .A2(n17851), .A3(n17850), .ZN(n17853) );
  NAND2_X1 U20853 ( .A1(n17853), .A2(n17861), .ZN(n17856) );
  AOI22_X1 U20854 ( .A1(n17951), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n17870), 
        .B2(n17854), .ZN(n17855) );
  OAI221_X1 U20855 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17857), .C1(
        n20633), .C2(n17856), .A(n17855), .ZN(P3_U2853) );
  INV_X1 U20856 ( .A(n17899), .ZN(n17863) );
  INV_X1 U20857 ( .A(n17936), .ZN(n17942) );
  INV_X1 U20858 ( .A(n17926), .ZN(n17902) );
  OAI21_X1 U20859 ( .B1(n17902), .B2(n17858), .A(n17900), .ZN(n17859) );
  OAI221_X1 U20860 ( .B1(n18406), .B2(n17865), .C1(n18406), .C2(n17923), .A(
        n17859), .ZN(n17886) );
  NOR2_X1 U20861 ( .A1(n17885), .A2(n17886), .ZN(n17877) );
  OAI211_X1 U20862 ( .C1(n17863), .C2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17952), .B(n17877), .ZN(n17860) );
  NAND2_X1 U20863 ( .A1(n17861), .A2(n17860), .ZN(n17884) );
  AOI211_X1 U20864 ( .C1(n17863), .C2(n17942), .A(n17862), .B(n17884), .ZN(
        n17868) );
  NOR2_X1 U20865 ( .A1(n17864), .A2(n17938), .ZN(n17915) );
  NAND2_X1 U20866 ( .A1(n17865), .A2(n17915), .ZN(n17892) );
  NOR3_X1 U20867 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17866), .A3(
        n17892), .ZN(n17867) );
  AOI211_X1 U20868 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n17951), .A(n17868), .B(
        n17867), .ZN(n17873) );
  AOI22_X1 U20869 ( .A1(n17957), .A2(n17871), .B1(n17870), .B2(n17869), .ZN(
        n17872) );
  OAI211_X1 U20870 ( .C1(n17875), .C2(n17874), .A(n17873), .B(n17872), .ZN(
        P3_U2854) );
  NOR3_X1 U20871 ( .A1(n17877), .A2(n17876), .A3(n17892), .ZN(n17879) );
  NOR2_X1 U20872 ( .A1(n17879), .A2(n17878), .ZN(n17883) );
  INV_X1 U20873 ( .A(n17949), .ZN(n17955) );
  AOI22_X1 U20874 ( .A1(n17955), .A2(n17881), .B1(n17957), .B2(n17880), .ZN(
        n17882) );
  OAI211_X1 U20875 ( .C1(n17885), .C2(n17884), .A(n17883), .B(n17882), .ZN(
        P3_U2855) );
  INV_X1 U20876 ( .A(n17886), .ZN(n17887) );
  OAI21_X1 U20877 ( .B1(n17887), .B2(n17938), .A(n17942), .ZN(n17895) );
  AOI22_X1 U20878 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17895), .B1(
        n17951), .B2(P3_REIP_REG_6__SCAN_IN), .ZN(n17891) );
  AOI22_X1 U20879 ( .A1(n17955), .A2(n17889), .B1(n17957), .B2(n17888), .ZN(
        n17890) );
  OAI211_X1 U20880 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n17892), .A(
        n17891), .B(n17890), .ZN(P3_U2856) );
  AOI22_X1 U20881 ( .A1(n17951), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n17957), 
        .B2(n17893), .ZN(n17898) );
  AOI22_X1 U20882 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17895), .B1(
        n17955), .B2(n17894), .ZN(n17897) );
  NAND4_X1 U20883 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n17915), .A4(n9946), .ZN(
        n17896) );
  NAND3_X1 U20884 ( .A1(n17898), .A2(n17897), .A3(n17896), .ZN(P3_U2857) );
  AND2_X1 U20885 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17915), .ZN(
        n17908) );
  NOR2_X1 U20886 ( .A1(n17936), .A2(n17899), .ZN(n17906) );
  OAI21_X1 U20887 ( .B1(n17902), .B2(n17901), .A(n17900), .ZN(n17903) );
  OAI211_X1 U20888 ( .C1(n18406), .C2(n17923), .A(n17952), .B(n17903), .ZN(
        n17904) );
  OAI21_X1 U20889 ( .B1(n17905), .B2(n17904), .A(n17861), .ZN(n17920) );
  NOR2_X1 U20890 ( .A1(n17906), .A2(n17920), .ZN(n17907) );
  MUX2_X1 U20891 ( .A(n17908), .B(n17907), .S(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n17909) );
  AOI21_X1 U20892 ( .B1(n17955), .B2(n17910), .A(n17909), .ZN(n17912) );
  NAND2_X1 U20893 ( .A1(n17951), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n17911) );
  OAI211_X1 U20894 ( .C1(n17914), .C2(n17913), .A(n17912), .B(n17911), .ZN(
        P3_U2858) );
  NOR2_X1 U20895 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17915), .ZN(
        n17921) );
  AOI22_X1 U20896 ( .A1(n17955), .A2(n17917), .B1(n17957), .B2(n17916), .ZN(
        n17919) );
  NAND2_X1 U20897 ( .A1(n17951), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n17918) );
  OAI211_X1 U20898 ( .C1(n17921), .C2(n17920), .A(n17919), .B(n17918), .ZN(
        P3_U2859) );
  OAI22_X1 U20899 ( .A1(n18406), .A2(n17923), .B1(n18425), .B2(n17922), .ZN(
        n17933) );
  INV_X1 U20900 ( .A(n17924), .ZN(n17925) );
  NOR2_X1 U20901 ( .A1(n18579), .A2(n17925), .ZN(n17931) );
  NOR2_X1 U20902 ( .A1(n18595), .A2(n18579), .ZN(n17928) );
  AOI21_X1 U20903 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17926), .A(
        n18399), .ZN(n17927) );
  AOI21_X1 U20904 ( .B1(n17928), .B2(n18438), .A(n17927), .ZN(n17929) );
  INV_X1 U20905 ( .A(n17929), .ZN(n17930) );
  MUX2_X1 U20906 ( .A(n17931), .B(n17930), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n17932) );
  AOI211_X1 U20907 ( .C1(n18428), .C2(n17934), .A(n17933), .B(n17932), .ZN(
        n17939) );
  AOI21_X1 U20908 ( .B1(n17936), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n17935), .ZN(n17937) );
  OAI21_X1 U20909 ( .B1(n17939), .B2(n17938), .A(n17937), .ZN(P3_U2860) );
  INV_X1 U20910 ( .A(n17940), .ZN(n17950) );
  NAND3_X1 U20911 ( .A1(n17952), .A2(n18595), .A3(n17941), .ZN(n17958) );
  AOI21_X1 U20912 ( .B1(n17942), .B2(n17958), .A(n18579), .ZN(n17945) );
  AOI211_X1 U20913 ( .C1(n18400), .C2(n18595), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n17943), .ZN(n17944) );
  AOI211_X1 U20914 ( .C1(n17957), .C2(n17946), .A(n17945), .B(n17944), .ZN(
        n17948) );
  NAND2_X1 U20915 ( .A1(n17951), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n17947) );
  OAI211_X1 U20916 ( .C1(n17950), .C2(n17949), .A(n17948), .B(n17947), .ZN(
        P3_U2861) );
  INV_X1 U20917 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18605) );
  AOI211_X1 U20918 ( .C1(n17952), .C2(n18400), .A(n17951), .B(n18595), .ZN(
        n17953) );
  AOI221_X1 U20919 ( .B1(n17957), .B2(n17956), .C1(n17955), .C2(n17954), .A(
        n17953), .ZN(n17959) );
  OAI211_X1 U20920 ( .C1(n18605), .C2(n17861), .A(n17959), .B(n17958), .ZN(
        P3_U2862) );
  INV_X1 U20921 ( .A(n17960), .ZN(n17961) );
  OAI21_X1 U20922 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n17962), .A(n17961), .ZN(
        n18466) );
  INV_X1 U20923 ( .A(n18466), .ZN(n17963) );
  OAI21_X1 U20924 ( .B1(n17963), .B2(n18228), .A(n17968), .ZN(n17964) );
  OAI221_X1 U20925 ( .B1(n18412), .B2(n18614), .C1(n18412), .C2(n17968), .A(
        n17964), .ZN(P3_U2863) );
  INV_X1 U20926 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18421) );
  NOR2_X1 U20927 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18421), .ZN(
        n18183) );
  NOR2_X1 U20928 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18420), .ZN(
        n18138) );
  NOR2_X1 U20929 ( .A1(n18183), .A2(n18138), .ZN(n17966) );
  OAI22_X1 U20930 ( .A1(n17967), .A2(n18421), .B1(n17966), .B2(n17965), .ZN(
        P3_U2866) );
  NOR2_X1 U20931 ( .A1(n18422), .A2(n17968), .ZN(P3_U2867) );
  NOR2_X1 U20932 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18416) );
  NOR2_X1 U20933 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18048) );
  NAND2_X1 U20934 ( .A1(n18416), .A2(n18048), .ZN(n18063) );
  NOR2_X1 U20935 ( .A1(n17970), .A2(n17969), .ZN(n17977) );
  NAND2_X1 U20936 ( .A1(n17977), .A2(n17971), .ZN(n18348) );
  NAND2_X1 U20937 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18275) );
  INV_X1 U20938 ( .A(n18275), .ZN(n18277) );
  NOR2_X1 U20939 ( .A1(n18412), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18182) );
  NAND2_X1 U20940 ( .A1(n18277), .A2(n18182), .ZN(n18381) );
  INV_X1 U20941 ( .A(n18381), .ZN(n18391) );
  AND2_X1 U20942 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18000), .ZN(n18340) );
  NOR2_X2 U20943 ( .A1(n18227), .A2(n17972), .ZN(n18341) );
  NOR2_X1 U20944 ( .A1(n18421), .A2(n18113), .ZN(n18343) );
  INV_X1 U20945 ( .A(n18343), .ZN(n18338) );
  NOR2_X2 U20946 ( .A1(n18412), .A2(n18338), .ZN(n18393) );
  INV_X1 U20947 ( .A(n18063), .ZN(n18066) );
  NOR2_X1 U20948 ( .A1(n18393), .A2(n18066), .ZN(n18028) );
  NOR2_X1 U20949 ( .A1(n18339), .A2(n18028), .ZN(n18003) );
  AOI22_X1 U20950 ( .A1(n18391), .A2(n18340), .B1(n18341), .B2(n18003), .ZN(
        n17975) );
  AOI21_X1 U20951 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18028), .ZN(n17973) );
  NAND2_X1 U20952 ( .A1(n18343), .A2(n18412), .ZN(n18310) );
  AOI21_X1 U20953 ( .B1(n18310), .B2(n18381), .A(n18227), .ZN(n18305) );
  AOI22_X1 U20954 ( .A1(n18253), .A2(n17973), .B1(n18115), .B2(n18305), .ZN(
        n18006) );
  NOR2_X2 U20955 ( .A1(n18302), .A2(n18947), .ZN(n18345) );
  INV_X1 U20956 ( .A(n18310), .ZN(n18333) );
  AOI22_X1 U20957 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18006), .B1(
        n18345), .B2(n18333), .ZN(n17974) );
  OAI211_X1 U20958 ( .C1(n18063), .C2(n18348), .A(n17975), .B(n17974), .ZN(
        P3_U2868) );
  NAND2_X1 U20959 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18000), .ZN(n18284) );
  NOR2_X2 U20960 ( .A1(n18302), .A2(n18953), .ZN(n18351) );
  NOR2_X2 U20961 ( .A1(n18227), .A2(n17976), .ZN(n18349) );
  AOI22_X1 U20962 ( .A1(n18333), .A2(n18351), .B1(n18003), .B2(n18349), .ZN(
        n17979) );
  INV_X1 U20963 ( .A(n17977), .ZN(n18004) );
  NOR2_X1 U20964 ( .A1(n18621), .A2(n18004), .ZN(n18281) );
  AOI22_X1 U20965 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18006), .B1(
        n18066), .B2(n18281), .ZN(n17978) );
  OAI211_X1 U20966 ( .C1(n18381), .C2(n18284), .A(n17979), .B(n17978), .ZN(
        P3_U2869) );
  NAND2_X1 U20967 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18000), .ZN(n18314) );
  NAND2_X1 U20968 ( .A1(n18000), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18361) );
  INV_X1 U20969 ( .A(n18361), .ZN(n18311) );
  NOR2_X2 U20970 ( .A1(n18227), .A2(n17980), .ZN(n18356) );
  AOI22_X1 U20971 ( .A1(n18333), .A2(n18311), .B1(n18003), .B2(n18356), .ZN(
        n17983) );
  NOR2_X2 U20972 ( .A1(n17981), .A2(n18004), .ZN(n18358) );
  AOI22_X1 U20973 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18006), .B1(
        n18066), .B2(n18358), .ZN(n17982) );
  OAI211_X1 U20974 ( .C1(n18381), .C2(n18314), .A(n17983), .B(n17982), .ZN(
        P3_U2870) );
  NAND2_X1 U20975 ( .A1(n18000), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18367) );
  NAND2_X1 U20976 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18000), .ZN(n18318) );
  INV_X1 U20977 ( .A(n18318), .ZN(n18363) );
  NOR2_X2 U20978 ( .A1(n18227), .A2(n17984), .ZN(n18362) );
  AOI22_X1 U20979 ( .A1(n18391), .A2(n18363), .B1(n18003), .B2(n18362), .ZN(
        n17987) );
  NOR2_X2 U20980 ( .A1(n17985), .A2(n18004), .ZN(n18364) );
  AOI22_X1 U20981 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18006), .B1(
        n18066), .B2(n18364), .ZN(n17986) );
  OAI211_X1 U20982 ( .C1(n18310), .C2(n18367), .A(n17987), .B(n17986), .ZN(
        P3_U2871) );
  NAND2_X1 U20983 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18000), .ZN(n18373) );
  NAND2_X1 U20984 ( .A1(n18000), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18322) );
  INV_X1 U20985 ( .A(n18322), .ZN(n18369) );
  NOR2_X2 U20986 ( .A1(n18227), .A2(n17988), .ZN(n18368) );
  AOI22_X1 U20987 ( .A1(n18333), .A2(n18369), .B1(n18003), .B2(n18368), .ZN(
        n17991) );
  NOR2_X2 U20988 ( .A1(n17989), .A2(n18004), .ZN(n18370) );
  AOI22_X1 U20989 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18006), .B1(
        n18066), .B2(n18370), .ZN(n17990) );
  OAI211_X1 U20990 ( .C1(n18381), .C2(n18373), .A(n17991), .B(n17990), .ZN(
        P3_U2872) );
  NAND2_X1 U20991 ( .A1(n18000), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18380) );
  NAND2_X1 U20992 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18000), .ZN(n18326) );
  INV_X1 U20993 ( .A(n18326), .ZN(n18376) );
  NOR2_X2 U20994 ( .A1(n18227), .A2(n17992), .ZN(n18374) );
  AOI22_X1 U20995 ( .A1(n18391), .A2(n18376), .B1(n18003), .B2(n18374), .ZN(
        n17995) );
  NOR2_X2 U20996 ( .A1(n17993), .A2(n18004), .ZN(n18377) );
  AOI22_X1 U20997 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18006), .B1(
        n18066), .B2(n18377), .ZN(n17994) );
  OAI211_X1 U20998 ( .C1(n18310), .C2(n18380), .A(n17995), .B(n17994), .ZN(
        P3_U2873) );
  NAND2_X1 U20999 ( .A1(n18000), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18331) );
  NAND2_X1 U21000 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18000), .ZN(n18387) );
  INV_X1 U21001 ( .A(n18387), .ZN(n18328) );
  NOR2_X2 U21002 ( .A1(n18227), .A2(n17996), .ZN(n18382) );
  AOI22_X1 U21003 ( .A1(n18391), .A2(n18328), .B1(n18003), .B2(n18382), .ZN(
        n17999) );
  NOR2_X2 U21004 ( .A1(n17997), .A2(n18004), .ZN(n18384) );
  AOI22_X1 U21005 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18006), .B1(
        n18066), .B2(n18384), .ZN(n17998) );
  OAI211_X1 U21006 ( .C1(n18310), .C2(n18331), .A(n17999), .B(n17998), .ZN(
        P3_U2874) );
  NAND2_X1 U21007 ( .A1(n18000), .A2(BUF2_REG_23__SCAN_IN), .ZN(n18301) );
  NOR2_X1 U21008 ( .A1(n18302), .A2(n18001), .ZN(n18297) );
  NOR2_X2 U21009 ( .A1(n18227), .A2(n18002), .ZN(n18389) );
  AOI22_X1 U21010 ( .A1(n18391), .A2(n18297), .B1(n18003), .B2(n18389), .ZN(
        n18008) );
  NOR2_X2 U21011 ( .A1(n18005), .A2(n18004), .ZN(n18392) );
  AOI22_X1 U21012 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18006), .B1(
        n18066), .B2(n18392), .ZN(n18007) );
  OAI211_X1 U21013 ( .C1(n18310), .C2(n18301), .A(n18008), .B(n18007), .ZN(
        P3_U2875) );
  NAND2_X1 U21014 ( .A1(n18048), .A2(n18182), .ZN(n18083) );
  INV_X1 U21015 ( .A(n18048), .ZN(n18027) );
  NAND2_X1 U21016 ( .A1(n18413), .A2(n18469), .ZN(n18274) );
  NOR2_X1 U21017 ( .A1(n18027), .A2(n18274), .ZN(n18023) );
  AOI22_X1 U21018 ( .A1(n18333), .A2(n18340), .B1(n18341), .B2(n18023), .ZN(
        n18010) );
  NOR3_X1 U21019 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18228), .A3(
        n18227), .ZN(n18276) );
  AOI22_X1 U21020 ( .A1(n18000), .A2(n18343), .B1(n18048), .B2(n18276), .ZN(
        n18024) );
  AOI22_X1 U21021 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18024), .B1(
        n18345), .B2(n18393), .ZN(n18009) );
  OAI211_X1 U21022 ( .C1(n18348), .C2(n18083), .A(n18010), .B(n18009), .ZN(
        P3_U2876) );
  INV_X1 U21023 ( .A(n18281), .ZN(n18354) );
  INV_X1 U21024 ( .A(n18284), .ZN(n18350) );
  AOI22_X1 U21025 ( .A1(n18333), .A2(n18350), .B1(n18349), .B2(n18023), .ZN(
        n18012) );
  AOI22_X1 U21026 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18024), .B1(
        n18393), .B2(n18351), .ZN(n18011) );
  OAI211_X1 U21027 ( .C1(n18354), .C2(n18083), .A(n18012), .B(n18011), .ZN(
        P3_U2877) );
  AOI22_X1 U21028 ( .A1(n18393), .A2(n18311), .B1(n18356), .B2(n18023), .ZN(
        n18014) );
  INV_X1 U21029 ( .A(n18083), .ZN(n18087) );
  AOI22_X1 U21030 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18024), .B1(
        n18358), .B2(n18087), .ZN(n18013) );
  OAI211_X1 U21031 ( .C1(n18310), .C2(n18314), .A(n18014), .B(n18013), .ZN(
        P3_U2878) );
  INV_X1 U21032 ( .A(n18393), .ZN(n18355) );
  AOI22_X1 U21033 ( .A1(n18333), .A2(n18363), .B1(n18362), .B2(n18023), .ZN(
        n18016) );
  AOI22_X1 U21034 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18024), .B1(
        n18364), .B2(n18087), .ZN(n18015) );
  OAI211_X1 U21035 ( .C1(n18355), .C2(n18367), .A(n18016), .B(n18015), .ZN(
        P3_U2879) );
  AOI22_X1 U21036 ( .A1(n18393), .A2(n18369), .B1(n18368), .B2(n18023), .ZN(
        n18018) );
  AOI22_X1 U21037 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18024), .B1(
        n18370), .B2(n18087), .ZN(n18017) );
  OAI211_X1 U21038 ( .C1(n18310), .C2(n18373), .A(n18018), .B(n18017), .ZN(
        P3_U2880) );
  INV_X1 U21039 ( .A(n18380), .ZN(n18323) );
  AOI22_X1 U21040 ( .A1(n18393), .A2(n18323), .B1(n18374), .B2(n18023), .ZN(
        n18020) );
  AOI22_X1 U21041 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18024), .B1(
        n18377), .B2(n18087), .ZN(n18019) );
  OAI211_X1 U21042 ( .C1(n18310), .C2(n18326), .A(n18020), .B(n18019), .ZN(
        P3_U2881) );
  INV_X1 U21043 ( .A(n18331), .ZN(n18383) );
  AOI22_X1 U21044 ( .A1(n18393), .A2(n18383), .B1(n18382), .B2(n18023), .ZN(
        n18022) );
  AOI22_X1 U21045 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18024), .B1(
        n18384), .B2(n18087), .ZN(n18021) );
  OAI211_X1 U21046 ( .C1(n18310), .C2(n18387), .A(n18022), .B(n18021), .ZN(
        P3_U2882) );
  AOI22_X1 U21047 ( .A1(n18333), .A2(n18297), .B1(n18389), .B2(n18023), .ZN(
        n18026) );
  AOI22_X1 U21048 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18024), .B1(
        n18392), .B2(n18087), .ZN(n18025) );
  OAI211_X1 U21049 ( .C1(n18355), .C2(n18301), .A(n18026), .B(n18025), .ZN(
        P3_U2883) );
  NOR2_X1 U21050 ( .A1(n18413), .A2(n18027), .ZN(n18092) );
  NAND2_X1 U21051 ( .A1(n18092), .A2(n18412), .ZN(n18112) );
  INV_X1 U21052 ( .A(n18112), .ZN(n18099) );
  NOR2_X1 U21053 ( .A1(n18087), .A2(n18099), .ZN(n18069) );
  NOR2_X1 U21054 ( .A1(n18339), .A2(n18069), .ZN(n18044) );
  AOI22_X1 U21055 ( .A1(n18345), .A2(n18066), .B1(n18341), .B2(n18044), .ZN(
        n18031) );
  OAI21_X1 U21056 ( .B1(n18028), .B2(n18250), .A(n18069), .ZN(n18029) );
  OAI211_X1 U21057 ( .C1(n18099), .C2(n18569), .A(n18253), .B(n18029), .ZN(
        n18045) );
  AOI22_X1 U21058 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18045), .B1(
        n18393), .B2(n18340), .ZN(n18030) );
  OAI211_X1 U21059 ( .C1(n18348), .C2(n18112), .A(n18031), .B(n18030), .ZN(
        P3_U2884) );
  AOI22_X1 U21060 ( .A1(n18393), .A2(n18350), .B1(n18349), .B2(n18044), .ZN(
        n18033) );
  AOI22_X1 U21061 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18045), .B1(
        n18066), .B2(n18351), .ZN(n18032) );
  OAI211_X1 U21062 ( .C1(n18354), .C2(n18112), .A(n18033), .B(n18032), .ZN(
        P3_U2885) );
  AOI22_X1 U21063 ( .A1(n18066), .A2(n18311), .B1(n18356), .B2(n18044), .ZN(
        n18035) );
  AOI22_X1 U21064 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18045), .B1(
        n18358), .B2(n18099), .ZN(n18034) );
  OAI211_X1 U21065 ( .C1(n18355), .C2(n18314), .A(n18035), .B(n18034), .ZN(
        P3_U2886) );
  INV_X1 U21066 ( .A(n18367), .ZN(n18315) );
  AOI22_X1 U21067 ( .A1(n18066), .A2(n18315), .B1(n18362), .B2(n18044), .ZN(
        n18037) );
  AOI22_X1 U21068 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18045), .B1(
        n18364), .B2(n18099), .ZN(n18036) );
  OAI211_X1 U21069 ( .C1(n18355), .C2(n18318), .A(n18037), .B(n18036), .ZN(
        P3_U2887) );
  INV_X1 U21070 ( .A(n18373), .ZN(n18319) );
  AOI22_X1 U21071 ( .A1(n18393), .A2(n18319), .B1(n18368), .B2(n18044), .ZN(
        n18039) );
  AOI22_X1 U21072 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18045), .B1(
        n18370), .B2(n18099), .ZN(n18038) );
  OAI211_X1 U21073 ( .C1(n18063), .C2(n18322), .A(n18039), .B(n18038), .ZN(
        P3_U2888) );
  AOI22_X1 U21074 ( .A1(n18393), .A2(n18376), .B1(n18374), .B2(n18044), .ZN(
        n18041) );
  AOI22_X1 U21075 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18045), .B1(
        n18377), .B2(n18099), .ZN(n18040) );
  OAI211_X1 U21076 ( .C1(n18063), .C2(n18380), .A(n18041), .B(n18040), .ZN(
        P3_U2889) );
  AOI22_X1 U21077 ( .A1(n18066), .A2(n18383), .B1(n18382), .B2(n18044), .ZN(
        n18043) );
  AOI22_X1 U21078 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18045), .B1(
        n18384), .B2(n18099), .ZN(n18042) );
  OAI211_X1 U21079 ( .C1(n18355), .C2(n18387), .A(n18043), .B(n18042), .ZN(
        P3_U2890) );
  INV_X1 U21080 ( .A(n18297), .ZN(n18398) );
  INV_X1 U21081 ( .A(n18301), .ZN(n18390) );
  AOI22_X1 U21082 ( .A1(n18066), .A2(n18390), .B1(n18389), .B2(n18044), .ZN(
        n18047) );
  AOI22_X1 U21083 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18045), .B1(
        n18392), .B2(n18099), .ZN(n18046) );
  OAI211_X1 U21084 ( .C1(n18355), .C2(n18398), .A(n18047), .B(n18046), .ZN(
        P3_U2891) );
  NAND2_X1 U21085 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18092), .ZN(
        n18136) );
  INV_X1 U21086 ( .A(n18136), .ZN(n18129) );
  AOI21_X1 U21087 ( .B1(n18413), .B2(n18250), .A(n18227), .ZN(n18137) );
  OAI211_X1 U21088 ( .C1(n18129), .C2(n18569), .A(n18048), .B(n18137), .ZN(
        n18065) );
  AND2_X1 U21089 ( .A1(n18469), .A2(n18092), .ZN(n18064) );
  AOI22_X1 U21090 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18065), .B1(
        n18341), .B2(n18064), .ZN(n18050) );
  AOI22_X1 U21091 ( .A1(n18345), .A2(n18087), .B1(n18066), .B2(n18340), .ZN(
        n18049) );
  OAI211_X1 U21092 ( .C1(n18348), .C2(n18136), .A(n18050), .B(n18049), .ZN(
        P3_U2892) );
  AOI22_X1 U21093 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18065), .B1(
        n18349), .B2(n18064), .ZN(n18052) );
  AOI22_X1 U21094 ( .A1(n18281), .A2(n18129), .B1(n18351), .B2(n18087), .ZN(
        n18051) );
  OAI211_X1 U21095 ( .C1(n18063), .C2(n18284), .A(n18052), .B(n18051), .ZN(
        P3_U2893) );
  AOI22_X1 U21096 ( .A1(n18311), .A2(n18087), .B1(n18356), .B2(n18064), .ZN(
        n18054) );
  AOI22_X1 U21097 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18065), .B1(
        n18358), .B2(n18129), .ZN(n18053) );
  OAI211_X1 U21098 ( .C1(n18063), .C2(n18314), .A(n18054), .B(n18053), .ZN(
        P3_U2894) );
  AOI22_X1 U21099 ( .A1(n18066), .A2(n18363), .B1(n18362), .B2(n18064), .ZN(
        n18056) );
  AOI22_X1 U21100 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18065), .B1(
        n18364), .B2(n18129), .ZN(n18055) );
  OAI211_X1 U21101 ( .C1(n18367), .C2(n18083), .A(n18056), .B(n18055), .ZN(
        P3_U2895) );
  AOI22_X1 U21102 ( .A1(n18369), .A2(n18087), .B1(n18368), .B2(n18064), .ZN(
        n18058) );
  AOI22_X1 U21103 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18065), .B1(
        n18370), .B2(n18129), .ZN(n18057) );
  OAI211_X1 U21104 ( .C1(n18063), .C2(n18373), .A(n18058), .B(n18057), .ZN(
        P3_U2896) );
  AOI22_X1 U21105 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18065), .B1(
        n18374), .B2(n18064), .ZN(n18060) );
  AOI22_X1 U21106 ( .A1(n18323), .A2(n18087), .B1(n18377), .B2(n18129), .ZN(
        n18059) );
  OAI211_X1 U21107 ( .C1(n18063), .C2(n18326), .A(n18060), .B(n18059), .ZN(
        P3_U2897) );
  AOI22_X1 U21108 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18065), .B1(
        n18382), .B2(n18064), .ZN(n18062) );
  AOI22_X1 U21109 ( .A1(n18383), .A2(n18087), .B1(n18384), .B2(n18129), .ZN(
        n18061) );
  OAI211_X1 U21110 ( .C1(n18063), .C2(n18387), .A(n18062), .B(n18061), .ZN(
        P3_U2898) );
  AOI22_X1 U21111 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18065), .B1(
        n18389), .B2(n18064), .ZN(n18068) );
  AOI22_X1 U21112 ( .A1(n18066), .A2(n18297), .B1(n18392), .B2(n18129), .ZN(
        n18067) );
  OAI211_X1 U21113 ( .C1(n18301), .C2(n18083), .A(n18068), .B(n18067), .ZN(
        P3_U2899) );
  NAND2_X1 U21114 ( .A1(n18416), .A2(n18138), .ZN(n18153) );
  AOI21_X1 U21115 ( .B1(n18136), .B2(n18153), .A(n18339), .ZN(n18086) );
  AOI22_X1 U21116 ( .A1(n18341), .A2(n18086), .B1(n18340), .B2(n18087), .ZN(
        n18072) );
  INV_X1 U21117 ( .A(n18153), .ZN(n18155) );
  AOI21_X1 U21118 ( .B1(n18136), .B2(n18153), .A(n18227), .ZN(n18114) );
  NOR2_X1 U21119 ( .A1(n18069), .A2(n18302), .ZN(n18070) );
  OAI22_X1 U21120 ( .A1(n18155), .A2(n18569), .B1(n18114), .B2(n18070), .ZN(
        n18088) );
  AOI22_X1 U21121 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18088), .B1(
        n18345), .B2(n18099), .ZN(n18071) );
  OAI211_X1 U21122 ( .C1(n18348), .C2(n18153), .A(n18072), .B(n18071), .ZN(
        P3_U2900) );
  AOI22_X1 U21123 ( .A1(n18350), .A2(n18087), .B1(n18349), .B2(n18086), .ZN(
        n18074) );
  AOI22_X1 U21124 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18088), .B1(
        n18351), .B2(n18099), .ZN(n18073) );
  OAI211_X1 U21125 ( .C1(n18354), .C2(n18153), .A(n18074), .B(n18073), .ZN(
        P3_U2901) );
  INV_X1 U21126 ( .A(n18314), .ZN(n18357) );
  AOI22_X1 U21127 ( .A1(n18357), .A2(n18087), .B1(n18356), .B2(n18086), .ZN(
        n18076) );
  AOI22_X1 U21128 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18088), .B1(
        n18358), .B2(n18155), .ZN(n18075) );
  OAI211_X1 U21129 ( .C1(n18361), .C2(n18112), .A(n18076), .B(n18075), .ZN(
        P3_U2902) );
  AOI22_X1 U21130 ( .A1(n18315), .A2(n18099), .B1(n18362), .B2(n18086), .ZN(
        n18078) );
  AOI22_X1 U21131 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18088), .B1(
        n18364), .B2(n18155), .ZN(n18077) );
  OAI211_X1 U21132 ( .C1(n18318), .C2(n18083), .A(n18078), .B(n18077), .ZN(
        P3_U2903) );
  AOI22_X1 U21133 ( .A1(n18319), .A2(n18087), .B1(n18368), .B2(n18086), .ZN(
        n18080) );
  AOI22_X1 U21134 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18088), .B1(
        n18370), .B2(n18155), .ZN(n18079) );
  OAI211_X1 U21135 ( .C1(n18322), .C2(n18112), .A(n18080), .B(n18079), .ZN(
        P3_U2904) );
  AOI22_X1 U21136 ( .A1(n18323), .A2(n18099), .B1(n18374), .B2(n18086), .ZN(
        n18082) );
  AOI22_X1 U21137 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18088), .B1(
        n18377), .B2(n18155), .ZN(n18081) );
  OAI211_X1 U21138 ( .C1(n18326), .C2(n18083), .A(n18082), .B(n18081), .ZN(
        P3_U2905) );
  AOI22_X1 U21139 ( .A1(n18328), .A2(n18087), .B1(n18382), .B2(n18086), .ZN(
        n18085) );
  AOI22_X1 U21140 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18088), .B1(
        n18384), .B2(n18155), .ZN(n18084) );
  OAI211_X1 U21141 ( .C1(n18331), .C2(n18112), .A(n18085), .B(n18084), .ZN(
        P3_U2906) );
  AOI22_X1 U21142 ( .A1(n18297), .A2(n18087), .B1(n18389), .B2(n18086), .ZN(
        n18090) );
  AOI22_X1 U21143 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18088), .B1(
        n18392), .B2(n18155), .ZN(n18089) );
  OAI211_X1 U21144 ( .C1(n18301), .C2(n18112), .A(n18090), .B(n18089), .ZN(
        P3_U2907) );
  NAND2_X1 U21145 ( .A1(n18138), .A2(n18182), .ZN(n18176) );
  INV_X1 U21146 ( .A(n18138), .ZN(n18091) );
  NOR2_X1 U21147 ( .A1(n18091), .A2(n18274), .ZN(n18108) );
  AOI22_X1 U21148 ( .A1(n18345), .A2(n18129), .B1(n18341), .B2(n18108), .ZN(
        n18094) );
  AOI22_X1 U21149 ( .A1(n18000), .A2(n18092), .B1(n18138), .B2(n18276), .ZN(
        n18109) );
  AOI22_X1 U21150 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18109), .B1(
        n18340), .B2(n18099), .ZN(n18093) );
  OAI211_X1 U21151 ( .C1(n18348), .C2(n18176), .A(n18094), .B(n18093), .ZN(
        P3_U2908) );
  AOI22_X1 U21152 ( .A1(n18351), .A2(n18129), .B1(n18349), .B2(n18108), .ZN(
        n18096) );
  AOI22_X1 U21153 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18109), .B1(
        n18350), .B2(n18099), .ZN(n18095) );
  OAI211_X1 U21154 ( .C1(n18354), .C2(n18176), .A(n18096), .B(n18095), .ZN(
        P3_U2909) );
  AOI22_X1 U21155 ( .A1(n18357), .A2(n18099), .B1(n18356), .B2(n18108), .ZN(
        n18098) );
  INV_X1 U21156 ( .A(n18176), .ZN(n18178) );
  AOI22_X1 U21157 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18109), .B1(
        n18358), .B2(n18178), .ZN(n18097) );
  OAI211_X1 U21158 ( .C1(n18361), .C2(n18136), .A(n18098), .B(n18097), .ZN(
        P3_U2910) );
  AOI22_X1 U21159 ( .A1(n18363), .A2(n18099), .B1(n18362), .B2(n18108), .ZN(
        n18101) );
  AOI22_X1 U21160 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18109), .B1(
        n18364), .B2(n18178), .ZN(n18100) );
  OAI211_X1 U21161 ( .C1(n18367), .C2(n18136), .A(n18101), .B(n18100), .ZN(
        P3_U2911) );
  AOI22_X1 U21162 ( .A1(n18369), .A2(n18129), .B1(n18368), .B2(n18108), .ZN(
        n18103) );
  AOI22_X1 U21163 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18109), .B1(
        n18370), .B2(n18178), .ZN(n18102) );
  OAI211_X1 U21164 ( .C1(n18373), .C2(n18112), .A(n18103), .B(n18102), .ZN(
        P3_U2912) );
  AOI22_X1 U21165 ( .A1(n18323), .A2(n18129), .B1(n18374), .B2(n18108), .ZN(
        n18105) );
  AOI22_X1 U21166 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18109), .B1(
        n18377), .B2(n18178), .ZN(n18104) );
  OAI211_X1 U21167 ( .C1(n18326), .C2(n18112), .A(n18105), .B(n18104), .ZN(
        P3_U2913) );
  AOI22_X1 U21168 ( .A1(n18383), .A2(n18129), .B1(n18382), .B2(n18108), .ZN(
        n18107) );
  AOI22_X1 U21169 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18109), .B1(
        n18384), .B2(n18178), .ZN(n18106) );
  OAI211_X1 U21170 ( .C1(n18387), .C2(n18112), .A(n18107), .B(n18106), .ZN(
        P3_U2914) );
  AOI22_X1 U21171 ( .A1(n18390), .A2(n18129), .B1(n18389), .B2(n18108), .ZN(
        n18111) );
  AOI22_X1 U21172 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18109), .B1(
        n18392), .B2(n18178), .ZN(n18110) );
  OAI211_X1 U21173 ( .C1(n18398), .C2(n18112), .A(n18111), .B(n18110), .ZN(
        P3_U2915) );
  NOR2_X1 U21174 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18113), .ZN(
        n18184) );
  NAND2_X1 U21175 ( .A1(n18184), .A2(n18412), .ZN(n18199) );
  AOI21_X1 U21176 ( .B1(n18176), .B2(n18199), .A(n18339), .ZN(n18132) );
  AOI22_X1 U21177 ( .A1(n18341), .A2(n18132), .B1(n18340), .B2(n18129), .ZN(
        n18118) );
  INV_X1 U21178 ( .A(n18199), .ZN(n18200) );
  AOI21_X1 U21179 ( .B1(n18176), .B2(n18199), .A(n18227), .ZN(n18159) );
  AND2_X1 U21180 ( .A1(n18115), .A2(n18114), .ZN(n18116) );
  OAI22_X1 U21181 ( .A1(n18200), .A2(n18569), .B1(n18159), .B2(n18116), .ZN(
        n18133) );
  AOI22_X1 U21182 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18133), .B1(
        n18345), .B2(n18155), .ZN(n18117) );
  OAI211_X1 U21183 ( .C1(n18348), .C2(n18199), .A(n18118), .B(n18117), .ZN(
        P3_U2916) );
  AOI22_X1 U21184 ( .A1(n18351), .A2(n18155), .B1(n18349), .B2(n18132), .ZN(
        n18120) );
  AOI22_X1 U21185 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18133), .B1(
        n18281), .B2(n18200), .ZN(n18119) );
  OAI211_X1 U21186 ( .C1(n18284), .C2(n18136), .A(n18120), .B(n18119), .ZN(
        P3_U2917) );
  AOI22_X1 U21187 ( .A1(n18357), .A2(n18129), .B1(n18356), .B2(n18132), .ZN(
        n18122) );
  AOI22_X1 U21188 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18133), .B1(
        n18358), .B2(n18200), .ZN(n18121) );
  OAI211_X1 U21189 ( .C1(n18361), .C2(n18153), .A(n18122), .B(n18121), .ZN(
        P3_U2918) );
  AOI22_X1 U21190 ( .A1(n18363), .A2(n18129), .B1(n18362), .B2(n18132), .ZN(
        n18124) );
  AOI22_X1 U21191 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18133), .B1(
        n18364), .B2(n18200), .ZN(n18123) );
  OAI211_X1 U21192 ( .C1(n18367), .C2(n18153), .A(n18124), .B(n18123), .ZN(
        P3_U2919) );
  AOI22_X1 U21193 ( .A1(n18319), .A2(n18129), .B1(n18368), .B2(n18132), .ZN(
        n18126) );
  AOI22_X1 U21194 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18133), .B1(
        n18370), .B2(n18200), .ZN(n18125) );
  OAI211_X1 U21195 ( .C1(n18322), .C2(n18153), .A(n18126), .B(n18125), .ZN(
        P3_U2920) );
  AOI22_X1 U21196 ( .A1(n18376), .A2(n18129), .B1(n18374), .B2(n18132), .ZN(
        n18128) );
  AOI22_X1 U21197 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18133), .B1(
        n18377), .B2(n18200), .ZN(n18127) );
  OAI211_X1 U21198 ( .C1(n18380), .C2(n18153), .A(n18128), .B(n18127), .ZN(
        P3_U2921) );
  AOI22_X1 U21199 ( .A1(n18328), .A2(n18129), .B1(n18382), .B2(n18132), .ZN(
        n18131) );
  AOI22_X1 U21200 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18133), .B1(
        n18384), .B2(n18200), .ZN(n18130) );
  OAI211_X1 U21201 ( .C1(n18331), .C2(n18153), .A(n18131), .B(n18130), .ZN(
        P3_U2922) );
  AOI22_X1 U21202 ( .A1(n18390), .A2(n18155), .B1(n18389), .B2(n18132), .ZN(
        n18135) );
  AOI22_X1 U21203 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18133), .B1(
        n18392), .B2(n18200), .ZN(n18134) );
  OAI211_X1 U21204 ( .C1(n18398), .C2(n18136), .A(n18135), .B(n18134), .ZN(
        P3_U2923) );
  NAND2_X1 U21205 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18184), .ZN(
        n18221) );
  INV_X1 U21206 ( .A(n18221), .ZN(n18223) );
  OAI211_X1 U21207 ( .C1(n18223), .C2(n18569), .A(n18138), .B(n18137), .ZN(
        n18156) );
  AND2_X1 U21208 ( .A1(n18469), .A2(n18184), .ZN(n18154) );
  AOI22_X1 U21209 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18156), .B1(
        n18341), .B2(n18154), .ZN(n18140) );
  AOI22_X1 U21210 ( .A1(n18345), .A2(n18178), .B1(n18340), .B2(n18155), .ZN(
        n18139) );
  OAI211_X1 U21211 ( .C1(n18348), .C2(n18221), .A(n18140), .B(n18139), .ZN(
        P3_U2924) );
  AOI22_X1 U21212 ( .A1(n18351), .A2(n18178), .B1(n18349), .B2(n18154), .ZN(
        n18142) );
  AOI22_X1 U21213 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18156), .B1(
        n18281), .B2(n18223), .ZN(n18141) );
  OAI211_X1 U21214 ( .C1(n18284), .C2(n18153), .A(n18142), .B(n18141), .ZN(
        P3_U2925) );
  AOI22_X1 U21215 ( .A1(n18357), .A2(n18155), .B1(n18356), .B2(n18154), .ZN(
        n18144) );
  AOI22_X1 U21216 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18156), .B1(
        n18358), .B2(n18223), .ZN(n18143) );
  OAI211_X1 U21217 ( .C1(n18361), .C2(n18176), .A(n18144), .B(n18143), .ZN(
        P3_U2926) );
  AOI22_X1 U21218 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18156), .B1(
        n18362), .B2(n18154), .ZN(n18146) );
  AOI22_X1 U21219 ( .A1(n18315), .A2(n18178), .B1(n18364), .B2(n18223), .ZN(
        n18145) );
  OAI211_X1 U21220 ( .C1(n18318), .C2(n18153), .A(n18146), .B(n18145), .ZN(
        P3_U2927) );
  AOI22_X1 U21221 ( .A1(n18369), .A2(n18178), .B1(n18368), .B2(n18154), .ZN(
        n18148) );
  AOI22_X1 U21222 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18156), .B1(
        n18370), .B2(n18223), .ZN(n18147) );
  OAI211_X1 U21223 ( .C1(n18373), .C2(n18153), .A(n18148), .B(n18147), .ZN(
        P3_U2928) );
  AOI22_X1 U21224 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18156), .B1(
        n18374), .B2(n18154), .ZN(n18150) );
  AOI22_X1 U21225 ( .A1(n18377), .A2(n18223), .B1(n18376), .B2(n18155), .ZN(
        n18149) );
  OAI211_X1 U21226 ( .C1(n18380), .C2(n18176), .A(n18150), .B(n18149), .ZN(
        P3_U2929) );
  AOI22_X1 U21227 ( .A1(n18383), .A2(n18178), .B1(n18382), .B2(n18154), .ZN(
        n18152) );
  AOI22_X1 U21228 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18156), .B1(
        n18384), .B2(n18223), .ZN(n18151) );
  OAI211_X1 U21229 ( .C1(n18387), .C2(n18153), .A(n18152), .B(n18151), .ZN(
        P3_U2930) );
  AOI22_X1 U21230 ( .A1(n18297), .A2(n18155), .B1(n18389), .B2(n18154), .ZN(
        n18158) );
  AOI22_X1 U21231 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18156), .B1(
        n18392), .B2(n18223), .ZN(n18157) );
  OAI211_X1 U21232 ( .C1(n18301), .C2(n18176), .A(n18158), .B(n18157), .ZN(
        P3_U2931) );
  NAND2_X1 U21233 ( .A1(n18416), .A2(n18183), .ZN(n18244) );
  INV_X1 U21234 ( .A(n18244), .ZN(n18246) );
  NOR2_X1 U21235 ( .A1(n18223), .A2(n18246), .ZN(n18205) );
  NOR2_X1 U21236 ( .A1(n18339), .A2(n18205), .ZN(n18177) );
  AOI22_X1 U21237 ( .A1(n18341), .A2(n18177), .B1(n18340), .B2(n18178), .ZN(
        n18163) );
  INV_X1 U21238 ( .A(n18159), .ZN(n18160) );
  OAI22_X1 U21239 ( .A1(n18205), .A2(n18227), .B1(n18250), .B2(n18160), .ZN(
        n18161) );
  OAI21_X1 U21240 ( .B1(n18246), .B2(n18569), .A(n18161), .ZN(n18179) );
  AOI22_X1 U21241 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18179), .B1(
        n18345), .B2(n18200), .ZN(n18162) );
  OAI211_X1 U21242 ( .C1(n18348), .C2(n18244), .A(n18163), .B(n18162), .ZN(
        P3_U2932) );
  AOI22_X1 U21243 ( .A1(n18351), .A2(n18200), .B1(n18349), .B2(n18177), .ZN(
        n18165) );
  AOI22_X1 U21244 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18179), .B1(
        n18281), .B2(n18246), .ZN(n18164) );
  OAI211_X1 U21245 ( .C1(n18284), .C2(n18176), .A(n18165), .B(n18164), .ZN(
        P3_U2933) );
  AOI22_X1 U21246 ( .A1(n18357), .A2(n18178), .B1(n18356), .B2(n18177), .ZN(
        n18167) );
  AOI22_X1 U21247 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18179), .B1(
        n18358), .B2(n18246), .ZN(n18166) );
  OAI211_X1 U21248 ( .C1(n18361), .C2(n18199), .A(n18167), .B(n18166), .ZN(
        P3_U2934) );
  AOI22_X1 U21249 ( .A1(n18315), .A2(n18200), .B1(n18362), .B2(n18177), .ZN(
        n18169) );
  AOI22_X1 U21250 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18179), .B1(
        n18364), .B2(n18246), .ZN(n18168) );
  OAI211_X1 U21251 ( .C1(n18318), .C2(n18176), .A(n18169), .B(n18168), .ZN(
        P3_U2935) );
  AOI22_X1 U21252 ( .A1(n18369), .A2(n18200), .B1(n18368), .B2(n18177), .ZN(
        n18171) );
  AOI22_X1 U21253 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18179), .B1(
        n18370), .B2(n18246), .ZN(n18170) );
  OAI211_X1 U21254 ( .C1(n18373), .C2(n18176), .A(n18171), .B(n18170), .ZN(
        P3_U2936) );
  AOI22_X1 U21255 ( .A1(n18376), .A2(n18178), .B1(n18374), .B2(n18177), .ZN(
        n18173) );
  AOI22_X1 U21256 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18179), .B1(
        n18377), .B2(n18246), .ZN(n18172) );
  OAI211_X1 U21257 ( .C1(n18380), .C2(n18199), .A(n18173), .B(n18172), .ZN(
        P3_U2937) );
  AOI22_X1 U21258 ( .A1(n18383), .A2(n18200), .B1(n18382), .B2(n18177), .ZN(
        n18175) );
  AOI22_X1 U21259 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18179), .B1(
        n18384), .B2(n18246), .ZN(n18174) );
  OAI211_X1 U21260 ( .C1(n18387), .C2(n18176), .A(n18175), .B(n18174), .ZN(
        P3_U2938) );
  AOI22_X1 U21261 ( .A1(n18297), .A2(n18178), .B1(n18389), .B2(n18177), .ZN(
        n18181) );
  AOI22_X1 U21262 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18179), .B1(
        n18392), .B2(n18246), .ZN(n18180) );
  OAI211_X1 U21263 ( .C1(n18301), .C2(n18199), .A(n18181), .B(n18180), .ZN(
        P3_U2939) );
  NAND2_X1 U21264 ( .A1(n18183), .A2(n18182), .ZN(n18273) );
  INV_X1 U21265 ( .A(n18183), .ZN(n18204) );
  NOR2_X1 U21266 ( .A1(n18204), .A2(n18274), .ZN(n18229) );
  AOI22_X1 U21267 ( .A1(n18341), .A2(n18229), .B1(n18340), .B2(n18200), .ZN(
        n18186) );
  AOI22_X1 U21268 ( .A1(n18000), .A2(n18184), .B1(n18183), .B2(n18276), .ZN(
        n18201) );
  AOI22_X1 U21269 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18201), .B1(
        n18345), .B2(n18223), .ZN(n18185) );
  OAI211_X1 U21270 ( .C1(n18348), .C2(n18273), .A(n18186), .B(n18185), .ZN(
        P3_U2940) );
  AOI22_X1 U21271 ( .A1(n18350), .A2(n18200), .B1(n18349), .B2(n18229), .ZN(
        n18188) );
  AOI22_X1 U21272 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18201), .B1(
        n18351), .B2(n18223), .ZN(n18187) );
  OAI211_X1 U21273 ( .C1(n18354), .C2(n18273), .A(n18188), .B(n18187), .ZN(
        P3_U2941) );
  AOI22_X1 U21274 ( .A1(n18311), .A2(n18223), .B1(n18356), .B2(n18229), .ZN(
        n18190) );
  INV_X1 U21275 ( .A(n18273), .ZN(n18266) );
  AOI22_X1 U21276 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18201), .B1(
        n18358), .B2(n18266), .ZN(n18189) );
  OAI211_X1 U21277 ( .C1(n18314), .C2(n18199), .A(n18190), .B(n18189), .ZN(
        P3_U2942) );
  AOI22_X1 U21278 ( .A1(n18363), .A2(n18200), .B1(n18362), .B2(n18229), .ZN(
        n18192) );
  AOI22_X1 U21279 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18201), .B1(
        n18364), .B2(n18266), .ZN(n18191) );
  OAI211_X1 U21280 ( .C1(n18367), .C2(n18221), .A(n18192), .B(n18191), .ZN(
        P3_U2943) );
  AOI22_X1 U21281 ( .A1(n18369), .A2(n18223), .B1(n18368), .B2(n18229), .ZN(
        n18194) );
  AOI22_X1 U21282 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18201), .B1(
        n18370), .B2(n18266), .ZN(n18193) );
  OAI211_X1 U21283 ( .C1(n18373), .C2(n18199), .A(n18194), .B(n18193), .ZN(
        P3_U2944) );
  AOI22_X1 U21284 ( .A1(n18323), .A2(n18223), .B1(n18374), .B2(n18229), .ZN(
        n18196) );
  AOI22_X1 U21285 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18201), .B1(
        n18377), .B2(n18266), .ZN(n18195) );
  OAI211_X1 U21286 ( .C1(n18326), .C2(n18199), .A(n18196), .B(n18195), .ZN(
        P3_U2945) );
  AOI22_X1 U21287 ( .A1(n18383), .A2(n18223), .B1(n18382), .B2(n18229), .ZN(
        n18198) );
  AOI22_X1 U21288 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18201), .B1(
        n18384), .B2(n18266), .ZN(n18197) );
  OAI211_X1 U21289 ( .C1(n18387), .C2(n18199), .A(n18198), .B(n18197), .ZN(
        P3_U2946) );
  AOI22_X1 U21290 ( .A1(n18297), .A2(n18200), .B1(n18389), .B2(n18229), .ZN(
        n18203) );
  AOI22_X1 U21291 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18201), .B1(
        n18392), .B2(n18266), .ZN(n18202) );
  OAI211_X1 U21292 ( .C1(n18301), .C2(n18221), .A(n18203), .B(n18202), .ZN(
        P3_U2947) );
  NOR2_X1 U21293 ( .A1(n18413), .A2(n18204), .ZN(n18278) );
  NAND2_X1 U21294 ( .A1(n18278), .A2(n18412), .ZN(n18293) );
  INV_X1 U21295 ( .A(n18293), .ZN(n18296) );
  NOR2_X1 U21296 ( .A1(n18266), .A2(n18296), .ZN(n18251) );
  NOR2_X1 U21297 ( .A1(n18339), .A2(n18251), .ZN(n18222) );
  AOI22_X1 U21298 ( .A1(n18341), .A2(n18222), .B1(n18340), .B2(n18223), .ZN(
        n18208) );
  OAI21_X1 U21299 ( .B1(n18205), .B2(n18250), .A(n18251), .ZN(n18206) );
  OAI211_X1 U21300 ( .C1(n18296), .C2(n18569), .A(n18253), .B(n18206), .ZN(
        n18224) );
  AOI22_X1 U21301 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18224), .B1(
        n18345), .B2(n18246), .ZN(n18207) );
  OAI211_X1 U21302 ( .C1(n18348), .C2(n18293), .A(n18208), .B(n18207), .ZN(
        P3_U2948) );
  AOI22_X1 U21303 ( .A1(n18351), .A2(n18246), .B1(n18349), .B2(n18222), .ZN(
        n18210) );
  AOI22_X1 U21304 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18224), .B1(
        n18281), .B2(n18296), .ZN(n18209) );
  OAI211_X1 U21305 ( .C1(n18284), .C2(n18221), .A(n18210), .B(n18209), .ZN(
        P3_U2949) );
  AOI22_X1 U21306 ( .A1(n18357), .A2(n18223), .B1(n18356), .B2(n18222), .ZN(
        n18212) );
  AOI22_X1 U21307 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18224), .B1(
        n18358), .B2(n18296), .ZN(n18211) );
  OAI211_X1 U21308 ( .C1(n18361), .C2(n18244), .A(n18212), .B(n18211), .ZN(
        P3_U2950) );
  AOI22_X1 U21309 ( .A1(n18363), .A2(n18223), .B1(n18362), .B2(n18222), .ZN(
        n18214) );
  AOI22_X1 U21310 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18224), .B1(
        n18364), .B2(n18296), .ZN(n18213) );
  OAI211_X1 U21311 ( .C1(n18367), .C2(n18244), .A(n18214), .B(n18213), .ZN(
        P3_U2951) );
  AOI22_X1 U21312 ( .A1(n18319), .A2(n18223), .B1(n18368), .B2(n18222), .ZN(
        n18216) );
  AOI22_X1 U21313 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18224), .B1(
        n18370), .B2(n18296), .ZN(n18215) );
  OAI211_X1 U21314 ( .C1(n18322), .C2(n18244), .A(n18216), .B(n18215), .ZN(
        P3_U2952) );
  AOI22_X1 U21315 ( .A1(n18376), .A2(n18223), .B1(n18374), .B2(n18222), .ZN(
        n18218) );
  AOI22_X1 U21316 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18224), .B1(
        n18377), .B2(n18296), .ZN(n18217) );
  OAI211_X1 U21317 ( .C1(n18380), .C2(n18244), .A(n18218), .B(n18217), .ZN(
        P3_U2953) );
  AOI22_X1 U21318 ( .A1(n18383), .A2(n18246), .B1(n18382), .B2(n18222), .ZN(
        n18220) );
  AOI22_X1 U21319 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18224), .B1(
        n18384), .B2(n18296), .ZN(n18219) );
  OAI211_X1 U21320 ( .C1(n18387), .C2(n18221), .A(n18220), .B(n18219), .ZN(
        P3_U2954) );
  AOI22_X1 U21321 ( .A1(n18297), .A2(n18223), .B1(n18389), .B2(n18222), .ZN(
        n18226) );
  AOI22_X1 U21322 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18224), .B1(
        n18392), .B2(n18296), .ZN(n18225) );
  OAI211_X1 U21323 ( .C1(n18301), .C2(n18244), .A(n18226), .B(n18225), .ZN(
        P3_U2955) );
  NAND2_X1 U21324 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18278), .ZN(
        n18337) );
  AND2_X1 U21325 ( .A1(n18469), .A2(n18278), .ZN(n18245) );
  AOI22_X1 U21326 ( .A1(n18341), .A2(n18245), .B1(n18340), .B2(n18246), .ZN(
        n18231) );
  NOR2_X1 U21327 ( .A1(n18228), .A2(n18227), .ZN(n18342) );
  AOI22_X1 U21328 ( .A1(n18000), .A2(n18229), .B1(n18342), .B2(n18278), .ZN(
        n18247) );
  AOI22_X1 U21329 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18247), .B1(
        n18345), .B2(n18266), .ZN(n18230) );
  OAI211_X1 U21330 ( .C1(n18348), .C2(n18337), .A(n18231), .B(n18230), .ZN(
        P3_U2956) );
  AOI22_X1 U21331 ( .A1(n18351), .A2(n18266), .B1(n18349), .B2(n18245), .ZN(
        n18233) );
  AOI22_X1 U21332 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18247), .B1(
        n18350), .B2(n18246), .ZN(n18232) );
  OAI211_X1 U21333 ( .C1(n18354), .C2(n18337), .A(n18233), .B(n18232), .ZN(
        P3_U2957) );
  AOI22_X1 U21334 ( .A1(n18357), .A2(n18246), .B1(n18356), .B2(n18245), .ZN(
        n18235) );
  INV_X1 U21335 ( .A(n18337), .ZN(n18327) );
  AOI22_X1 U21336 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18247), .B1(
        n18358), .B2(n18327), .ZN(n18234) );
  OAI211_X1 U21337 ( .C1(n18361), .C2(n18273), .A(n18235), .B(n18234), .ZN(
        P3_U2958) );
  AOI22_X1 U21338 ( .A1(n18363), .A2(n18246), .B1(n18362), .B2(n18245), .ZN(
        n18237) );
  AOI22_X1 U21339 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18247), .B1(
        n18364), .B2(n18327), .ZN(n18236) );
  OAI211_X1 U21340 ( .C1(n18367), .C2(n18273), .A(n18237), .B(n18236), .ZN(
        P3_U2959) );
  AOI22_X1 U21341 ( .A1(n18369), .A2(n18266), .B1(n18368), .B2(n18245), .ZN(
        n18239) );
  AOI22_X1 U21342 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18247), .B1(
        n18370), .B2(n18327), .ZN(n18238) );
  OAI211_X1 U21343 ( .C1(n18373), .C2(n18244), .A(n18239), .B(n18238), .ZN(
        P3_U2960) );
  AOI22_X1 U21344 ( .A1(n18376), .A2(n18246), .B1(n18374), .B2(n18245), .ZN(
        n18241) );
  AOI22_X1 U21345 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18247), .B1(
        n18377), .B2(n18327), .ZN(n18240) );
  OAI211_X1 U21346 ( .C1(n18380), .C2(n18273), .A(n18241), .B(n18240), .ZN(
        P3_U2961) );
  AOI22_X1 U21347 ( .A1(n18383), .A2(n18266), .B1(n18382), .B2(n18245), .ZN(
        n18243) );
  AOI22_X1 U21348 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18247), .B1(
        n18384), .B2(n18327), .ZN(n18242) );
  OAI211_X1 U21349 ( .C1(n18387), .C2(n18244), .A(n18243), .B(n18242), .ZN(
        P3_U2962) );
  AOI22_X1 U21350 ( .A1(n18297), .A2(n18246), .B1(n18389), .B2(n18245), .ZN(
        n18249) );
  AOI22_X1 U21351 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18247), .B1(
        n18392), .B2(n18327), .ZN(n18248) );
  OAI211_X1 U21352 ( .C1(n18301), .C2(n18273), .A(n18249), .B(n18248), .ZN(
        P3_U2963) );
  NAND2_X1 U21353 ( .A1(n18416), .A2(n18277), .ZN(n18397) );
  INV_X1 U21354 ( .A(n18397), .ZN(n18375) );
  NOR2_X1 U21355 ( .A1(n18327), .A2(n18375), .ZN(n18303) );
  NOR2_X1 U21356 ( .A1(n18339), .A2(n18303), .ZN(n18269) );
  AOI22_X1 U21357 ( .A1(n18341), .A2(n18269), .B1(n18340), .B2(n18266), .ZN(
        n18255) );
  OAI21_X1 U21358 ( .B1(n18251), .B2(n18250), .A(n18303), .ZN(n18252) );
  OAI211_X1 U21359 ( .C1(n18375), .C2(n18569), .A(n18253), .B(n18252), .ZN(
        n18270) );
  AOI22_X1 U21360 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18270), .B1(
        n18345), .B2(n18296), .ZN(n18254) );
  OAI211_X1 U21361 ( .C1(n18348), .C2(n18397), .A(n18255), .B(n18254), .ZN(
        P3_U2964) );
  AOI22_X1 U21362 ( .A1(n18350), .A2(n18266), .B1(n18349), .B2(n18269), .ZN(
        n18257) );
  AOI22_X1 U21363 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18270), .B1(
        n18351), .B2(n18296), .ZN(n18256) );
  OAI211_X1 U21364 ( .C1(n18354), .C2(n18397), .A(n18257), .B(n18256), .ZN(
        P3_U2965) );
  AOI22_X1 U21365 ( .A1(n18357), .A2(n18266), .B1(n18356), .B2(n18269), .ZN(
        n18259) );
  AOI22_X1 U21366 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18270), .B1(
        n18358), .B2(n18375), .ZN(n18258) );
  OAI211_X1 U21367 ( .C1(n18361), .C2(n18293), .A(n18259), .B(n18258), .ZN(
        P3_U2966) );
  AOI22_X1 U21368 ( .A1(n18315), .A2(n18296), .B1(n18362), .B2(n18269), .ZN(
        n18261) );
  AOI22_X1 U21369 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18270), .B1(
        n18364), .B2(n18375), .ZN(n18260) );
  OAI211_X1 U21370 ( .C1(n18318), .C2(n18273), .A(n18261), .B(n18260), .ZN(
        P3_U2967) );
  AOI22_X1 U21371 ( .A1(n18369), .A2(n18296), .B1(n18368), .B2(n18269), .ZN(
        n18263) );
  AOI22_X1 U21372 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18270), .B1(
        n18370), .B2(n18375), .ZN(n18262) );
  OAI211_X1 U21373 ( .C1(n18373), .C2(n18273), .A(n18263), .B(n18262), .ZN(
        P3_U2968) );
  AOI22_X1 U21374 ( .A1(n18323), .A2(n18296), .B1(n18374), .B2(n18269), .ZN(
        n18265) );
  AOI22_X1 U21375 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18270), .B1(
        n18377), .B2(n18375), .ZN(n18264) );
  OAI211_X1 U21376 ( .C1(n18326), .C2(n18273), .A(n18265), .B(n18264), .ZN(
        P3_U2969) );
  AOI22_X1 U21377 ( .A1(n18328), .A2(n18266), .B1(n18382), .B2(n18269), .ZN(
        n18268) );
  AOI22_X1 U21378 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18270), .B1(
        n18384), .B2(n18375), .ZN(n18267) );
  OAI211_X1 U21379 ( .C1(n18331), .C2(n18293), .A(n18268), .B(n18267), .ZN(
        P3_U2970) );
  AOI22_X1 U21380 ( .A1(n18390), .A2(n18296), .B1(n18389), .B2(n18269), .ZN(
        n18272) );
  AOI22_X1 U21381 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18270), .B1(
        n18392), .B2(n18375), .ZN(n18271) );
  OAI211_X1 U21382 ( .C1(n18398), .C2(n18273), .A(n18272), .B(n18271), .ZN(
        P3_U2971) );
  NOR2_X1 U21383 ( .A1(n18275), .A2(n18274), .ZN(n18344) );
  AOI22_X1 U21384 ( .A1(n18341), .A2(n18344), .B1(n18340), .B2(n18296), .ZN(
        n18280) );
  AOI22_X1 U21385 ( .A1(n18000), .A2(n18278), .B1(n18277), .B2(n18276), .ZN(
        n18298) );
  AOI22_X1 U21386 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18298), .B1(
        n18345), .B2(n18327), .ZN(n18279) );
  OAI211_X1 U21387 ( .C1(n18381), .C2(n18348), .A(n18280), .B(n18279), .ZN(
        P3_U2972) );
  AOI22_X1 U21388 ( .A1(n18351), .A2(n18327), .B1(n18349), .B2(n18344), .ZN(
        n18283) );
  AOI22_X1 U21389 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18298), .B1(
        n18391), .B2(n18281), .ZN(n18282) );
  OAI211_X1 U21390 ( .C1(n18284), .C2(n18293), .A(n18283), .B(n18282), .ZN(
        P3_U2973) );
  AOI22_X1 U21391 ( .A1(n18357), .A2(n18296), .B1(n18356), .B2(n18344), .ZN(
        n18286) );
  AOI22_X1 U21392 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18298), .B1(
        n18391), .B2(n18358), .ZN(n18285) );
  OAI211_X1 U21393 ( .C1(n18361), .C2(n18337), .A(n18286), .B(n18285), .ZN(
        P3_U2974) );
  AOI22_X1 U21394 ( .A1(n18315), .A2(n18327), .B1(n18362), .B2(n18344), .ZN(
        n18288) );
  AOI22_X1 U21395 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18298), .B1(
        n18391), .B2(n18364), .ZN(n18287) );
  OAI211_X1 U21396 ( .C1(n18318), .C2(n18293), .A(n18288), .B(n18287), .ZN(
        P3_U2975) );
  AOI22_X1 U21397 ( .A1(n18369), .A2(n18327), .B1(n18368), .B2(n18344), .ZN(
        n18290) );
  AOI22_X1 U21398 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18298), .B1(
        n18391), .B2(n18370), .ZN(n18289) );
  OAI211_X1 U21399 ( .C1(n18373), .C2(n18293), .A(n18290), .B(n18289), .ZN(
        P3_U2976) );
  AOI22_X1 U21400 ( .A1(n18323), .A2(n18327), .B1(n18374), .B2(n18344), .ZN(
        n18292) );
  AOI22_X1 U21401 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18298), .B1(
        n18391), .B2(n18377), .ZN(n18291) );
  OAI211_X1 U21402 ( .C1(n18326), .C2(n18293), .A(n18292), .B(n18291), .ZN(
        P3_U2977) );
  AOI22_X1 U21403 ( .A1(n18328), .A2(n18296), .B1(n18382), .B2(n18344), .ZN(
        n18295) );
  AOI22_X1 U21404 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18298), .B1(
        n18391), .B2(n18384), .ZN(n18294) );
  OAI211_X1 U21405 ( .C1(n18331), .C2(n18337), .A(n18295), .B(n18294), .ZN(
        P3_U2978) );
  AOI22_X1 U21406 ( .A1(n18297), .A2(n18296), .B1(n18389), .B2(n18344), .ZN(
        n18300) );
  AOI22_X1 U21407 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18298), .B1(
        n18391), .B2(n18392), .ZN(n18299) );
  OAI211_X1 U21408 ( .C1(n18301), .C2(n18337), .A(n18300), .B(n18299), .ZN(
        P3_U2979) );
  AOI21_X1 U21409 ( .B1(n18310), .B2(n18381), .A(n18339), .ZN(n18332) );
  AOI22_X1 U21410 ( .A1(n18341), .A2(n18332), .B1(n18340), .B2(n18327), .ZN(
        n18307) );
  NOR2_X1 U21411 ( .A1(n18303), .A2(n18302), .ZN(n18304) );
  OAI22_X1 U21412 ( .A1(n18333), .A2(n18569), .B1(n18305), .B2(n18304), .ZN(
        n18334) );
  AOI22_X1 U21413 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18334), .B1(
        n18345), .B2(n18375), .ZN(n18306) );
  OAI211_X1 U21414 ( .C1(n18310), .C2(n18348), .A(n18307), .B(n18306), .ZN(
        P3_U2980) );
  AOI22_X1 U21415 ( .A1(n18350), .A2(n18327), .B1(n18349), .B2(n18332), .ZN(
        n18309) );
  AOI22_X1 U21416 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18334), .B1(
        n18351), .B2(n18375), .ZN(n18308) );
  OAI211_X1 U21417 ( .C1(n18310), .C2(n18354), .A(n18309), .B(n18308), .ZN(
        P3_U2981) );
  AOI22_X1 U21418 ( .A1(n18311), .A2(n18375), .B1(n18356), .B2(n18332), .ZN(
        n18313) );
  AOI22_X1 U21419 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18334), .B1(
        n18333), .B2(n18358), .ZN(n18312) );
  OAI211_X1 U21420 ( .C1(n18314), .C2(n18337), .A(n18313), .B(n18312), .ZN(
        P3_U2982) );
  AOI22_X1 U21421 ( .A1(n18315), .A2(n18375), .B1(n18362), .B2(n18332), .ZN(
        n18317) );
  AOI22_X1 U21422 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18334), .B1(
        n18333), .B2(n18364), .ZN(n18316) );
  OAI211_X1 U21423 ( .C1(n18318), .C2(n18337), .A(n18317), .B(n18316), .ZN(
        P3_U2983) );
  AOI22_X1 U21424 ( .A1(n18319), .A2(n18327), .B1(n18368), .B2(n18332), .ZN(
        n18321) );
  AOI22_X1 U21425 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18334), .B1(
        n18333), .B2(n18370), .ZN(n18320) );
  OAI211_X1 U21426 ( .C1(n18322), .C2(n18397), .A(n18321), .B(n18320), .ZN(
        P3_U2984) );
  AOI22_X1 U21427 ( .A1(n18323), .A2(n18375), .B1(n18374), .B2(n18332), .ZN(
        n18325) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18334), .B1(
        n18333), .B2(n18377), .ZN(n18324) );
  OAI211_X1 U21429 ( .C1(n18326), .C2(n18337), .A(n18325), .B(n18324), .ZN(
        P3_U2985) );
  AOI22_X1 U21430 ( .A1(n18328), .A2(n18327), .B1(n18382), .B2(n18332), .ZN(
        n18330) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18334), .B1(
        n18333), .B2(n18384), .ZN(n18329) );
  OAI211_X1 U21432 ( .C1(n18331), .C2(n18397), .A(n18330), .B(n18329), .ZN(
        P3_U2986) );
  AOI22_X1 U21433 ( .A1(n18390), .A2(n18375), .B1(n18389), .B2(n18332), .ZN(
        n18336) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18334), .B1(
        n18333), .B2(n18392), .ZN(n18335) );
  OAI211_X1 U21435 ( .C1(n18398), .C2(n18337), .A(n18336), .B(n18335), .ZN(
        P3_U2987) );
  NOR2_X1 U21436 ( .A1(n18339), .A2(n18338), .ZN(n18388) );
  AOI22_X1 U21437 ( .A1(n18341), .A2(n18388), .B1(n18340), .B2(n18375), .ZN(
        n18347) );
  AOI22_X1 U21438 ( .A1(n18000), .A2(n18344), .B1(n18343), .B2(n18342), .ZN(
        n18394) );
  AOI22_X1 U21439 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18394), .B1(
        n18345), .B2(n18391), .ZN(n18346) );
  OAI211_X1 U21440 ( .C1(n18355), .C2(n18348), .A(n18347), .B(n18346), .ZN(
        P3_U2988) );
  AOI22_X1 U21441 ( .A1(n18350), .A2(n18375), .B1(n18349), .B2(n18388), .ZN(
        n18353) );
  AOI22_X1 U21442 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18394), .B1(
        n18391), .B2(n18351), .ZN(n18352) );
  OAI211_X1 U21443 ( .C1(n18355), .C2(n18354), .A(n18353), .B(n18352), .ZN(
        P3_U2989) );
  AOI22_X1 U21444 ( .A1(n18357), .A2(n18375), .B1(n18356), .B2(n18388), .ZN(
        n18360) );
  AOI22_X1 U21445 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18358), .ZN(n18359) );
  OAI211_X1 U21446 ( .C1(n18381), .C2(n18361), .A(n18360), .B(n18359), .ZN(
        P3_U2990) );
  AOI22_X1 U21447 ( .A1(n18363), .A2(n18375), .B1(n18362), .B2(n18388), .ZN(
        n18366) );
  AOI22_X1 U21448 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18364), .ZN(n18365) );
  OAI211_X1 U21449 ( .C1(n18381), .C2(n18367), .A(n18366), .B(n18365), .ZN(
        P3_U2991) );
  AOI22_X1 U21450 ( .A1(n18391), .A2(n18369), .B1(n18368), .B2(n18388), .ZN(
        n18372) );
  AOI22_X1 U21451 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18370), .ZN(n18371) );
  OAI211_X1 U21452 ( .C1(n18373), .C2(n18397), .A(n18372), .B(n18371), .ZN(
        P3_U2992) );
  AOI22_X1 U21453 ( .A1(n18376), .A2(n18375), .B1(n18374), .B2(n18388), .ZN(
        n18379) );
  AOI22_X1 U21454 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18377), .ZN(n18378) );
  OAI211_X1 U21455 ( .C1(n18381), .C2(n18380), .A(n18379), .B(n18378), .ZN(
        P3_U2993) );
  AOI22_X1 U21456 ( .A1(n18391), .A2(n18383), .B1(n18382), .B2(n18388), .ZN(
        n18386) );
  AOI22_X1 U21457 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18384), .ZN(n18385) );
  OAI211_X1 U21458 ( .C1(n18387), .C2(n18397), .A(n18386), .B(n18385), .ZN(
        P3_U2994) );
  AOI22_X1 U21459 ( .A1(n18391), .A2(n18390), .B1(n18389), .B2(n18388), .ZN(
        n18396) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18392), .ZN(n18395) );
  OAI211_X1 U21461 ( .C1(n18398), .C2(n18397), .A(n18396), .B(n18395), .ZN(
        P3_U2995) );
  AOI21_X1 U21462 ( .B1(n18400), .B2(n13689), .A(n18399), .ZN(n18437) );
  OAI211_X1 U21463 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18437), .B(n18432), .ZN(
        n18405) );
  OAI21_X1 U21464 ( .B1(n18403), .B2(n18402), .A(n18401), .ZN(n18430) );
  NAND3_X1 U21465 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18434), .A3(
        n18430), .ZN(n18404) );
  OAI211_X1 U21466 ( .C1(n18580), .C2(n18406), .A(n18405), .B(n18404), .ZN(
        n18581) );
  MUX2_X1 U21467 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n18581), .S(
        n18450), .Z(n18419) );
  INV_X1 U21468 ( .A(n18419), .ZN(n18445) );
  INV_X1 U21469 ( .A(n18407), .ZN(n18588) );
  NAND2_X1 U21470 ( .A1(n18409), .A2(n18408), .ZN(n18410) );
  AOI22_X1 U21471 ( .A1(n18588), .A2(n18410), .B1(n18437), .B2(n18591), .ZN(
        n18584) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18411), .B1(
        n18410), .B2(n13689), .ZN(n18414) );
  INV_X1 U21473 ( .A(n18414), .ZN(n18593) );
  NOR3_X1 U21474 ( .A1(n18413), .A2(n18412), .A3(n18593), .ZN(n18415) );
  OAI22_X1 U21475 ( .A1(n18584), .A2(n18415), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18414), .ZN(n18417) );
  AOI21_X1 U21476 ( .B1(n18417), .B2(n18450), .A(n18416), .ZN(n18418) );
  AOI21_X1 U21477 ( .B1(n18445), .B2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n18418), .ZN(n18444) );
  AOI21_X1 U21478 ( .B1(n18420), .B2(n18419), .A(n18444), .ZN(n18458) );
  NAND2_X1 U21479 ( .A1(n18422), .A2(n18421), .ZN(n18457) );
  OAI22_X1 U21480 ( .A1(n18426), .A2(n18425), .B1(n18424), .B2(n18423), .ZN(
        n18427) );
  AOI221_X1 U21481 ( .B1(n18438), .B2(n18429), .C1(n18428), .C2(n18429), .A(
        n18427), .ZN(n18612) );
  AOI22_X1 U21482 ( .A1(n18433), .A2(n18432), .B1(n18431), .B2(n18430), .ZN(
        n18435) );
  NAND2_X1 U21483 ( .A1(n18583), .A2(n18434), .ZN(n18439) );
  NAND2_X1 U21484 ( .A1(n18435), .A2(n18439), .ZN(n18573) );
  NOR2_X1 U21485 ( .A1(n18573), .A2(n18442), .ZN(n18443) );
  AOI22_X1 U21486 ( .A1(n18439), .A2(n18438), .B1(n18437), .B2(n18436), .ZN(
        n18440) );
  NOR2_X1 U21487 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18440), .ZN(
        n18572) );
  INV_X1 U21488 ( .A(n18572), .ZN(n18441) );
  OAI22_X1 U21489 ( .A1(n18574), .A2(n18443), .B1(n18442), .B2(n18441), .ZN(
        n18455) );
  INV_X1 U21490 ( .A(n18444), .ZN(n18446) );
  OAI221_X1 U21491 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n18446), .A(n18445), .ZN(
        n18454) );
  OAI21_X1 U21492 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18447), .ZN(n18448) );
  OAI211_X1 U21493 ( .C1(n18451), .C2(n18450), .A(n18449), .B(n18448), .ZN(
        n18452) );
  AOI211_X1 U21494 ( .C1(n18455), .C2(n18454), .A(n18453), .B(n18452), .ZN(
        n18456) );
  OAI211_X1 U21495 ( .C1(n18458), .C2(n18457), .A(n18612), .B(n18456), .ZN(
        n18464) );
  AOI211_X1 U21496 ( .C1(n18461), .C2(n18460), .A(n18459), .B(n18464), .ZN(
        n18567) );
  AOI21_X1 U21497 ( .B1(n18617), .B2(n18468), .A(n18567), .ZN(n18470) );
  INV_X1 U21498 ( .A(n18477), .ZN(n18625) );
  NOR2_X1 U21499 ( .A1(n18622), .A2(n18616), .ZN(n18467) );
  AOI211_X1 U21500 ( .C1(n18592), .C2(n18625), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n18467), .ZN(n18462) );
  AOI211_X1 U21501 ( .C1(n18615), .C2(n18464), .A(n18463), .B(n18462), .ZN(
        n18465) );
  OAI221_X1 U21502 ( .B1(n18566), .B2(n18470), .C1(n18566), .C2(n18466), .A(
        n18465), .ZN(P3_U2996) );
  INV_X1 U21503 ( .A(n18467), .ZN(n18473) );
  NAND4_X1 U21504 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n18617), .A4(n18468), .ZN(n18475) );
  NAND3_X1 U21505 ( .A1(n18471), .A2(n18470), .A3(n18469), .ZN(n18472) );
  NAND4_X1 U21506 ( .A1(n18474), .A2(n18473), .A3(n18475), .A4(n18472), .ZN(
        P3_U2997) );
  AND4_X1 U21507 ( .A1(n18477), .A2(n18476), .A3(n18475), .A4(n18568), .ZN(
        P3_U2998) );
  AND2_X1 U21508 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18562), .ZN(
        P3_U2999) );
  AND2_X1 U21509 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18562), .ZN(
        P3_U3000) );
  AND2_X1 U21510 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18562), .ZN(
        P3_U3001) );
  AND2_X1 U21511 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18562), .ZN(
        P3_U3002) );
  AND2_X1 U21512 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18562), .ZN(
        P3_U3003) );
  AND2_X1 U21513 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18562), .ZN(
        P3_U3004) );
  AND2_X1 U21514 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18562), .ZN(
        P3_U3005) );
  AND2_X1 U21515 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18562), .ZN(
        P3_U3006) );
  AND2_X1 U21516 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18562), .ZN(
        P3_U3007) );
  AND2_X1 U21517 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18562), .ZN(
        P3_U3008) );
  AND2_X1 U21518 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18562), .ZN(
        P3_U3009) );
  AND2_X1 U21519 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18562), .ZN(
        P3_U3010) );
  AND2_X1 U21520 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18562), .ZN(
        P3_U3011) );
  AND2_X1 U21521 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18562), .ZN(
        P3_U3012) );
  AND2_X1 U21522 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18562), .ZN(
        P3_U3013) );
  AND2_X1 U21523 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18562), .ZN(
        P3_U3014) );
  AND2_X1 U21524 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18562), .ZN(
        P3_U3015) );
  AND2_X1 U21525 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18562), .ZN(
        P3_U3016) );
  AND2_X1 U21526 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18562), .ZN(
        P3_U3017) );
  AND2_X1 U21527 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18562), .ZN(
        P3_U3018) );
  AND2_X1 U21528 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18562), .ZN(
        P3_U3019) );
  AND2_X1 U21529 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18562), .ZN(
        P3_U3020) );
  AND2_X1 U21530 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18562), .ZN(P3_U3021) );
  AND2_X1 U21531 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18562), .ZN(P3_U3022) );
  AND2_X1 U21532 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18562), .ZN(P3_U3023) );
  AND2_X1 U21533 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18562), .ZN(P3_U3024) );
  AND2_X1 U21534 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18562), .ZN(P3_U3025) );
  AND2_X1 U21535 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18562), .ZN(P3_U3026) );
  AND2_X1 U21536 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18562), .ZN(P3_U3027) );
  AND2_X1 U21537 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18562), .ZN(P3_U3028) );
  NOR2_X1 U21538 ( .A1(n18493), .A2(n20782), .ZN(n18488) );
  INV_X1 U21539 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18481) );
  AOI211_X1 U21540 ( .C1(HOLD), .C2(P3_STATE_REG_1__SCAN_IN), .A(n18488), .B(
        n18481), .ZN(n18480) );
  NAND2_X1 U21541 ( .A1(n18617), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18486) );
  AND2_X1 U21542 ( .A1(n18486), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18492) );
  INV_X1 U21543 ( .A(NA), .ZN(n20513) );
  OAI21_X1 U21544 ( .B1(n20513), .B2(n18478), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18491) );
  INV_X1 U21545 ( .A(n18491), .ZN(n18479) );
  OAI22_X1 U21546 ( .A1(n18630), .A2(n18480), .B1(n18492), .B2(n18479), .ZN(
        P3_U3029) );
  NOR2_X1 U21547 ( .A1(n18488), .A2(n18481), .ZN(n18484) );
  NOR2_X1 U21548 ( .A1(n18482), .A2(n20782), .ZN(n18483) );
  AOI22_X1 U21549 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18484), .B1(n18483), 
        .B2(n18493), .ZN(n18485) );
  NAND3_X1 U21550 ( .A1(n18485), .A2(n18619), .A3(n18486), .ZN(P3_U3030) );
  OAI22_X1 U21551 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18486), .ZN(n18487) );
  OAI22_X1 U21552 ( .A1(n18488), .A2(n18487), .B1(HOLD), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18489) );
  OAI22_X1 U21553 ( .A1(n18492), .A2(n18491), .B1(n18490), .B2(n18489), .ZN(
        P3_U3031) );
  NAND2_X1 U21554 ( .A1(n18630), .A2(n18493), .ZN(n18541) );
  CLKBUF_X1 U21555 ( .A(n18541), .Z(n18550) );
  OAI222_X1 U21556 ( .A1(n18599), .A2(n18553), .B1(n18494), .B2(n18630), .C1(
        n18495), .C2(n18550), .ZN(P3_U3032) );
  OAI222_X1 U21557 ( .A1(n18541), .A2(n18497), .B1(n18496), .B2(n18630), .C1(
        n18495), .C2(n18553), .ZN(P3_U3033) );
  OAI222_X1 U21558 ( .A1(n18541), .A2(n18499), .B1(n18498), .B2(n18630), .C1(
        n18497), .C2(n18553), .ZN(P3_U3034) );
  INV_X1 U21559 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18502) );
  OAI222_X1 U21560 ( .A1(n18541), .A2(n18502), .B1(n18500), .B2(n18630), .C1(
        n18499), .C2(n18553), .ZN(P3_U3035) );
  OAI222_X1 U21561 ( .A1(n18502), .A2(n18553), .B1(n18501), .B2(n18630), .C1(
        n20788), .C2(n18550), .ZN(P3_U3036) );
  OAI222_X1 U21562 ( .A1(n20788), .A2(n18553), .B1(n18503), .B2(n18630), .C1(
        n18504), .C2(n18550), .ZN(P3_U3037) );
  OAI222_X1 U21563 ( .A1(n18541), .A2(n18507), .B1(n18505), .B2(n18630), .C1(
        n18504), .C2(n18553), .ZN(P3_U3038) );
  OAI222_X1 U21564 ( .A1(n18507), .A2(n18553), .B1(n18506), .B2(n18630), .C1(
        n18508), .C2(n18550), .ZN(P3_U3039) );
  OAI222_X1 U21565 ( .A1(n18541), .A2(n18509), .B1(n20762), .B2(n18630), .C1(
        n18508), .C2(n18553), .ZN(P3_U3040) );
  OAI222_X1 U21566 ( .A1(n18541), .A2(n18511), .B1(n18510), .B2(n18630), .C1(
        n18509), .C2(n18553), .ZN(P3_U3041) );
  OAI222_X1 U21567 ( .A1(n18550), .A2(n18513), .B1(n18512), .B2(n18630), .C1(
        n18511), .C2(n18553), .ZN(P3_U3042) );
  OAI222_X1 U21568 ( .A1(n18550), .A2(n18515), .B1(n18514), .B2(n18630), .C1(
        n18513), .C2(n18553), .ZN(P3_U3043) );
  OAI222_X1 U21569 ( .A1(n18550), .A2(n18517), .B1(n18516), .B2(n18630), .C1(
        n18515), .C2(n18553), .ZN(P3_U3044) );
  OAI222_X1 U21570 ( .A1(n18550), .A2(n18519), .B1(n18518), .B2(n18630), .C1(
        n18517), .C2(n18553), .ZN(P3_U3045) );
  OAI222_X1 U21571 ( .A1(n18550), .A2(n18521), .B1(n18520), .B2(n18630), .C1(
        n18519), .C2(n18553), .ZN(P3_U3046) );
  OAI222_X1 U21572 ( .A1(n18550), .A2(n18524), .B1(n18522), .B2(n18630), .C1(
        n18521), .C2(n18553), .ZN(P3_U3047) );
  OAI222_X1 U21573 ( .A1(n18524), .A2(n18553), .B1(n18523), .B2(n18630), .C1(
        n18525), .C2(n18550), .ZN(P3_U3048) );
  OAI222_X1 U21574 ( .A1(n18541), .A2(n18527), .B1(n18526), .B2(n18630), .C1(
        n18525), .C2(n18553), .ZN(P3_U3049) );
  OAI222_X1 U21575 ( .A1(n18541), .A2(n18530), .B1(n18528), .B2(n18630), .C1(
        n18527), .C2(n18553), .ZN(P3_U3050) );
  OAI222_X1 U21576 ( .A1(n18530), .A2(n18553), .B1(n18529), .B2(n18630), .C1(
        n18531), .C2(n18550), .ZN(P3_U3051) );
  OAI222_X1 U21577 ( .A1(n18541), .A2(n18533), .B1(n18532), .B2(n18630), .C1(
        n18531), .C2(n18553), .ZN(P3_U3052) );
  OAI222_X1 U21578 ( .A1(n18541), .A2(n18536), .B1(n18534), .B2(n18630), .C1(
        n18533), .C2(n18553), .ZN(P3_U3053) );
  OAI222_X1 U21579 ( .A1(n18536), .A2(n18553), .B1(n18535), .B2(n18630), .C1(
        n18537), .C2(n18550), .ZN(P3_U3054) );
  OAI222_X1 U21580 ( .A1(n18541), .A2(n18539), .B1(n18538), .B2(n18630), .C1(
        n18537), .C2(n18553), .ZN(P3_U3055) );
  OAI222_X1 U21581 ( .A1(n18541), .A2(n18542), .B1(n18540), .B2(n18630), .C1(
        n18539), .C2(n18553), .ZN(P3_U3056) );
  OAI222_X1 U21582 ( .A1(n18550), .A2(n18544), .B1(n18543), .B2(n18630), .C1(
        n18542), .C2(n18553), .ZN(P3_U3057) );
  OAI222_X1 U21583 ( .A1(n18550), .A2(n18547), .B1(n18545), .B2(n18630), .C1(
        n18544), .C2(n18553), .ZN(P3_U3058) );
  OAI222_X1 U21584 ( .A1(n18547), .A2(n18553), .B1(n18546), .B2(n18630), .C1(
        n18548), .C2(n18550), .ZN(P3_U3059) );
  OAI222_X1 U21585 ( .A1(n18550), .A2(n20804), .B1(n18549), .B2(n18630), .C1(
        n18548), .C2(n18553), .ZN(P3_U3060) );
  OAI222_X1 U21586 ( .A1(n18553), .A2(n20804), .B1(n18552), .B2(n18630), .C1(
        n18551), .C2(n18550), .ZN(P3_U3061) );
  INV_X1 U21587 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18554) );
  AOI22_X1 U21588 ( .A1(n18630), .A2(n18555), .B1(n18554), .B2(n18608), .ZN(
        P3_U3274) );
  INV_X1 U21589 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18601) );
  INV_X1 U21590 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18556) );
  AOI22_X1 U21591 ( .A1(n18630), .A2(n18601), .B1(n18556), .B2(n18608), .ZN(
        P3_U3275) );
  INV_X1 U21592 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18557) );
  AOI22_X1 U21593 ( .A1(n18630), .A2(n18558), .B1(n18557), .B2(n18608), .ZN(
        P3_U3276) );
  INV_X1 U21594 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18607) );
  INV_X1 U21595 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18559) );
  AOI22_X1 U21596 ( .A1(n18630), .A2(n18607), .B1(n18559), .B2(n18608), .ZN(
        P3_U3277) );
  INV_X1 U21597 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18561) );
  INV_X1 U21598 ( .A(n18563), .ZN(n18560) );
  AOI21_X1 U21599 ( .B1(n18562), .B2(n18561), .A(n18560), .ZN(P3_U3280) );
  OAI21_X1 U21600 ( .B1(n18565), .B2(n18564), .A(n18563), .ZN(P3_U3281) );
  NOR2_X1 U21601 ( .A1(n18567), .A2(n18566), .ZN(n18570) );
  OAI21_X1 U21602 ( .B1(n18570), .B2(n18569), .A(n18568), .ZN(P3_U3282) );
  INV_X1 U21603 ( .A(n18596), .ZN(n18598) );
  AOI22_X1 U21604 ( .A1(n18594), .A2(n18572), .B1(n18592), .B2(n18571), .ZN(
        n18576) );
  AOI21_X1 U21605 ( .B1(n18594), .B2(n18573), .A(n18598), .ZN(n18575) );
  OAI22_X1 U21606 ( .A1(n18598), .A2(n18576), .B1(n18575), .B2(n18574), .ZN(
        P3_U3285) );
  NOR2_X1 U21607 ( .A1(n18577), .A2(n18595), .ZN(n18586) );
  AOI22_X1 U21608 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18579), .B2(n18578), .ZN(
        n18585) );
  AOI222_X1 U21609 ( .A1(n18581), .A2(n18594), .B1(n18586), .B2(n18585), .C1(
        n18592), .C2(n18580), .ZN(n18582) );
  AOI22_X1 U21610 ( .A1(n18598), .A2(n18583), .B1(n18582), .B2(n18596), .ZN(
        P3_U3288) );
  INV_X1 U21611 ( .A(n18584), .ZN(n18589) );
  INV_X1 U21612 ( .A(n18585), .ZN(n18587) );
  AOI222_X1 U21613 ( .A1(n18589), .A2(n18594), .B1(n18592), .B2(n18588), .C1(
        n18587), .C2(n18586), .ZN(n18590) );
  AOI22_X1 U21614 ( .A1(n18598), .A2(n18591), .B1(n18590), .B2(n18596), .ZN(
        P3_U3289) );
  AOI222_X1 U21615 ( .A1(n18595), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18594), 
        .B2(n18593), .C1(n13689), .C2(n18592), .ZN(n18597) );
  AOI22_X1 U21616 ( .A1(n18598), .A2(n13689), .B1(n18597), .B2(n18596), .ZN(
        P3_U3290) );
  AOI21_X1 U21617 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18600) );
  AOI22_X1 U21618 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18600), .B2(n18599), .ZN(n18602) );
  AOI22_X1 U21619 ( .A1(n18603), .A2(n18602), .B1(n18601), .B2(n18606), .ZN(
        P3_U3292) );
  NOR2_X1 U21620 ( .A1(n18606), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18604) );
  AOI22_X1 U21621 ( .A1(n18607), .A2(n18606), .B1(n18605), .B2(n18604), .ZN(
        P3_U3293) );
  INV_X1 U21622 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18609) );
  AOI22_X1 U21623 ( .A1(n18630), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18609), 
        .B2(n18608), .ZN(P3_U3294) );
  INV_X1 U21624 ( .A(n18610), .ZN(n18613) );
  NAND2_X1 U21625 ( .A1(n18613), .A2(P3_MORE_REG_SCAN_IN), .ZN(n18611) );
  OAI21_X1 U21626 ( .B1(n18613), .B2(n18612), .A(n18611), .ZN(P3_U3295) );
  OAI22_X1 U21627 ( .A1(n18617), .A2(n18616), .B1(n18615), .B2(n18614), .ZN(
        n18618) );
  NOR2_X1 U21628 ( .A1(n18637), .A2(n18618), .ZN(n18629) );
  AOI21_X1 U21629 ( .B1(n18621), .B2(n18620), .A(n18619), .ZN(n18623) );
  OAI211_X1 U21630 ( .C1(n18624), .C2(n18623), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18622), .ZN(n18626) );
  AOI21_X1 U21631 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18626), .A(n18625), 
        .ZN(n18628) );
  NAND2_X1 U21632 ( .A1(n18629), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18627) );
  OAI21_X1 U21633 ( .B1(n18629), .B2(n18628), .A(n18627), .ZN(P3_U3296) );
  MUX2_X1 U21634 ( .A(P3_M_IO_N_REG_SCAN_IN), .B(P3_MEMORYFETCH_REG_SCAN_IN), 
        .S(n18630), .Z(P3_U3297) );
  INV_X1 U21635 ( .A(n18637), .ZN(n18633) );
  OAI21_X1 U21636 ( .B1(n18634), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n18633), 
        .ZN(n18631) );
  OAI21_X1 U21637 ( .B1(n18633), .B2(n18632), .A(n18631), .ZN(P3_U3298) );
  NOR2_X1 U21638 ( .A1(n18634), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18636)
         );
  OAI21_X1 U21639 ( .B1(n18637), .B2(n18636), .A(n18635), .ZN(P3_U3299) );
  INV_X1 U21640 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19505) );
  INV_X1 U21641 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18638) );
  INV_X1 U21642 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19525) );
  NAND2_X1 U21643 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19525), .ZN(n19513) );
  AOI22_X1 U21644 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19513), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n19505), .ZN(n19578) );
  INV_X1 U21645 ( .A(n19578), .ZN(n19503) );
  OAI21_X1 U21646 ( .B1(n19505), .B2(n18638), .A(n19503), .ZN(P2_U2815) );
  INV_X1 U21647 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18641) );
  OAI22_X1 U21648 ( .A1(n18642), .A2(n18641), .B1(n18640), .B2(n18639), .ZN(
        P2_U2816) );
  INV_X1 U21649 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19517) );
  OR2_X1 U21650 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19517), .ZN(n19624) );
  INV_X2 U21651 ( .A(n19624), .ZN(n19627) );
  OR2_X1 U21652 ( .A1(n19516), .A2(n19627), .ZN(n19508) );
  AOI21_X1 U21653 ( .B1(n19505), .B2(n19508), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18643) );
  AOI21_X1 U21654 ( .B1(n19627), .B2(P2_CODEFETCH_REG_SCAN_IN), .A(n18643), 
        .ZN(P2_U2817) );
  OAI21_X1 U21655 ( .B1(n19516), .B2(BS16), .A(n19578), .ZN(n19576) );
  OAI21_X1 U21656 ( .B1(n19578), .B2(n19294), .A(n19576), .ZN(P2_U2818) );
  NOR2_X1 U21657 ( .A1(n18644), .A2(n19494), .ZN(n19622) );
  OAI21_X1 U21658 ( .B1(n19622), .B2(n10797), .A(n18645), .ZN(P2_U2819) );
  NOR4_X1 U21659 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18649) );
  NOR4_X1 U21660 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18648) );
  NOR4_X1 U21661 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18647) );
  NOR4_X1 U21662 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18646) );
  NAND4_X1 U21663 ( .A1(n18649), .A2(n18648), .A3(n18647), .A4(n18646), .ZN(
        n18655) );
  NOR4_X1 U21664 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18653) );
  AOI211_X1 U21665 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n18652) );
  NOR4_X1 U21666 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18651) );
  NOR4_X1 U21667 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18650) );
  NAND4_X1 U21668 ( .A1(n18653), .A2(n18652), .A3(n18651), .A4(n18650), .ZN(
        n18654) );
  NOR2_X1 U21669 ( .A1(n18655), .A2(n18654), .ZN(n18663) );
  INV_X1 U21670 ( .A(n18663), .ZN(n18656) );
  NOR2_X1 U21671 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18656), .ZN(n18658) );
  INV_X1 U21672 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19574) );
  AOI22_X1 U21673 ( .A1(n18658), .A2(n10280), .B1(n18656), .B2(n19574), .ZN(
        P2_U2820) );
  NOR2_X1 U21674 ( .A1(n18663), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18657)
         );
  OR4_X1 U21675 ( .A1(n18656), .A2(P2_REIP_REG_0__SCAN_IN), .A3(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A4(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18662) );
  OAI21_X1 U21676 ( .B1(n18658), .B2(n18657), .A(n18662), .ZN(P2_U2821) );
  INV_X1 U21677 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19577) );
  NAND2_X1 U21678 ( .A1(n18658), .A2(n19577), .ZN(n18661) );
  OAI21_X1 U21679 ( .B1(n10280), .B2(n12768), .A(n18663), .ZN(n18659) );
  OAI21_X1 U21680 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18663), .A(n18659), 
        .ZN(n18660) );
  OAI221_X1 U21681 ( .B1(n18661), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18661), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18660), .ZN(P2_U2822) );
  INV_X1 U21682 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19573) );
  OAI211_X1 U21683 ( .C1(n18663), .C2(n19573), .A(n18662), .B(n18661), .ZN(
        P2_U2823) );
  NOR2_X1 U21684 ( .A1(n18785), .A2(n18664), .ZN(n18686) );
  XOR2_X1 U21685 ( .A(n18686), .B(n18665), .Z(n18675) );
  AOI22_X1 U21686 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(n18819), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n9607), .ZN(n18666) );
  OAI21_X1 U21687 ( .B1(n18667), .B2(n18795), .A(n18666), .ZN(n18668) );
  AOI211_X1 U21688 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n18669), .A(n18933), 
        .B(n18668), .ZN(n18674) );
  OAI22_X1 U21689 ( .A1(n18671), .A2(n18789), .B1(n18812), .B2(n18670), .ZN(
        n18672) );
  INV_X1 U21690 ( .A(n18672), .ZN(n18673) );
  OAI211_X1 U21691 ( .C1(n18779), .C2(n18675), .A(n18674), .B(n18673), .ZN(
        P2_U2837) );
  OAI22_X1 U21692 ( .A1(n18676), .A2(n18694), .B1(n19545), .B2(n18810), .ZN(
        n18677) );
  AOI211_X1 U21693 ( .C1(n18682), .C2(n18826), .A(n18933), .B(n18677), .ZN(
        n18678) );
  OAI21_X1 U21694 ( .B1(n18679), .B2(n18795), .A(n18678), .ZN(n18680) );
  AOI21_X1 U21695 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n18819), .A(n18680), .ZN(
        n18688) );
  AOI21_X1 U21696 ( .B1(n18682), .B2(n18681), .A(n18779), .ZN(n18685) );
  INV_X1 U21697 ( .A(n18683), .ZN(n18684) );
  AOI22_X1 U21698 ( .A1(n18686), .A2(n18685), .B1(n18814), .B2(n18684), .ZN(
        n18687) );
  OAI211_X1 U21699 ( .C1(n18689), .C2(n18812), .A(n18688), .B(n18687), .ZN(
        P2_U2838) );
  NOR2_X1 U21700 ( .A1(n18785), .A2(n18690), .ZN(n18692) );
  XOR2_X1 U21701 ( .A(n18692), .B(n18691), .Z(n18702) );
  OAI21_X1 U21702 ( .B1(n11108), .B2(n18810), .A(n11181), .ZN(n18697) );
  OAI22_X1 U21703 ( .A1(n18695), .A2(n18694), .B1(n18693), .B2(n18795), .ZN(
        n18696) );
  AOI211_X1 U21704 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n18819), .A(n18697), .B(
        n18696), .ZN(n18701) );
  INV_X1 U21705 ( .A(n18883), .ZN(n18698) );
  OAI22_X1 U21706 ( .A1(n18836), .A2(n18789), .B1(n18812), .B2(n18698), .ZN(
        n18699) );
  INV_X1 U21707 ( .A(n18699), .ZN(n18700) );
  OAI211_X1 U21708 ( .C1(n18779), .C2(n18702), .A(n18701), .B(n18700), .ZN(
        P2_U2839) );
  NAND2_X1 U21709 ( .A1(n13264), .A2(n18703), .ZN(n18705) );
  XOR2_X1 U21710 ( .A(n18705), .B(n18704), .Z(n18714) );
  AOI22_X1 U21711 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n9607), .B1(
        n18706), .B2(n18818), .ZN(n18707) );
  OAI211_X1 U21712 ( .C1(n19542), .C2(n18810), .A(n18707), .B(n11181), .ZN(
        n18712) );
  INV_X1 U21713 ( .A(n18708), .ZN(n18710) );
  OAI22_X1 U21714 ( .A1(n18710), .A2(n18789), .B1(n18812), .B2(n18709), .ZN(
        n18711) );
  AOI211_X1 U21715 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n18819), .A(n18712), .B(
        n18711), .ZN(n18713) );
  OAI21_X1 U21716 ( .B1(n18714), .B2(n18779), .A(n18713), .ZN(P2_U2840) );
  NOR2_X1 U21717 ( .A1(n18785), .A2(n18715), .ZN(n18717) );
  XOR2_X1 U21718 ( .A(n18717), .B(n18716), .Z(n18725) );
  AOI22_X1 U21719 ( .A1(P2_EBX_REG_14__SCAN_IN), .A2(n18819), .B1(n18718), 
        .B2(n18818), .ZN(n18719) );
  OAI211_X1 U21720 ( .C1(n11102), .C2(n18810), .A(n18719), .B(n16010), .ZN(
        n18720) );
  AOI21_X1 U21721 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n9607), .A(
        n18720), .ZN(n18724) );
  OAI22_X1 U21722 ( .A1(n18721), .A2(n18812), .B1(n18789), .B2(n18843), .ZN(
        n18722) );
  INV_X1 U21723 ( .A(n18722), .ZN(n18723) );
  OAI211_X1 U21724 ( .C1(n18779), .C2(n18725), .A(n18724), .B(n18723), .ZN(
        P2_U2841) );
  NOR2_X1 U21725 ( .A1(n18785), .A2(n18726), .ZN(n18727) );
  XOR2_X1 U21726 ( .A(n18728), .B(n18727), .Z(n18734) );
  AOI22_X1 U21727 ( .A1(P2_EBX_REG_12__SCAN_IN), .A2(n18819), .B1(n18729), 
        .B2(n18818), .ZN(n18730) );
  OAI211_X1 U21728 ( .C1(n11092), .C2(n18810), .A(n18730), .B(n16010), .ZN(
        n18732) );
  OAI22_X1 U21729 ( .A1(n18892), .A2(n18812), .B1(n18789), .B2(n18851), .ZN(
        n18731) );
  AOI211_X1 U21730 ( .C1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n9607), .A(
        n18732), .B(n18731), .ZN(n18733) );
  OAI21_X1 U21731 ( .B1(n18779), .B2(n18734), .A(n18733), .ZN(P2_U2843) );
  OAI21_X1 U21732 ( .B1(n11088), .B2(n18810), .A(n11181), .ZN(n18738) );
  OAI22_X1 U21733 ( .A1(n18798), .A2(n18736), .B1(n18735), .B2(n18795), .ZN(
        n18737) );
  AOI211_X1 U21734 ( .C1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n9607), .A(
        n18738), .B(n18737), .ZN(n18745) );
  NAND2_X1 U21735 ( .A1(n13264), .A2(n18739), .ZN(n18740) );
  XNOR2_X1 U21736 ( .A(n18741), .B(n18740), .ZN(n18743) );
  AOI22_X1 U21737 ( .A1(n18743), .A2(n19499), .B1(n18814), .B2(n18742), .ZN(
        n18744) );
  OAI211_X1 U21738 ( .C1(n18746), .C2(n18812), .A(n18745), .B(n18744), .ZN(
        P2_U2844) );
  NOR2_X1 U21739 ( .A1(n18785), .A2(n18747), .ZN(n18748) );
  XOR2_X1 U21740 ( .A(n18749), .B(n18748), .Z(n18757) );
  INV_X1 U21741 ( .A(n18750), .ZN(n18751) );
  AOI22_X1 U21742 ( .A1(n18751), .A2(n18818), .B1(P2_EBX_REG_10__SCAN_IN), 
        .B2(n18819), .ZN(n18752) );
  OAI211_X1 U21743 ( .C1(n10939), .C2(n18810), .A(n18752), .B(n11181), .ZN(
        n18755) );
  INV_X1 U21744 ( .A(n18856), .ZN(n18753) );
  OAI22_X1 U21745 ( .A1(n18753), .A2(n18789), .B1(n18812), .B2(n18897), .ZN(
        n18754) );
  AOI211_X1 U21746 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n9607), .A(
        n18755), .B(n18754), .ZN(n18756) );
  OAI21_X1 U21747 ( .B1(n18779), .B2(n18757), .A(n18756), .ZN(P2_U2845) );
  OAI21_X1 U21748 ( .B1(n19535), .B2(n18810), .A(n11181), .ZN(n18760) );
  OAI22_X1 U21749 ( .A1(n18758), .A2(n18795), .B1(n18798), .B2(n11083), .ZN(
        n18759) );
  AOI211_X1 U21750 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n9607), .A(
        n18760), .B(n18759), .ZN(n18767) );
  NAND2_X1 U21751 ( .A1(n13264), .A2(n18761), .ZN(n18762) );
  XNOR2_X1 U21752 ( .A(n18763), .B(n18762), .ZN(n18765) );
  AOI22_X1 U21753 ( .A1(n18765), .A2(n19499), .B1(n18814), .B2(n18764), .ZN(
        n18766) );
  OAI211_X1 U21754 ( .C1(n18768), .C2(n18812), .A(n18767), .B(n18766), .ZN(
        P2_U2846) );
  NAND2_X1 U21755 ( .A1(n13264), .A2(n18769), .ZN(n18771) );
  XOR2_X1 U21756 ( .A(n18771), .B(n18770), .Z(n18780) );
  AOI22_X1 U21757 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n9607), .B1(
        n18772), .B2(n18818), .ZN(n18773) );
  OAI211_X1 U21758 ( .C1(n19532), .C2(n18810), .A(n18773), .B(n16010), .ZN(
        n18777) );
  OAI22_X1 U21759 ( .A1(n18775), .A2(n18812), .B1(n18789), .B2(n18774), .ZN(
        n18776) );
  AOI211_X1 U21760 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n18819), .A(n18777), .B(
        n18776), .ZN(n18778) );
  OAI21_X1 U21761 ( .B1(n18780), .B2(n18779), .A(n18778), .ZN(P2_U2848) );
  AOI22_X1 U21762 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n9607), .B1(
        n18781), .B2(n18818), .ZN(n18782) );
  OAI211_X1 U21763 ( .C1(n11057), .C2(n18810), .A(n11181), .B(n18782), .ZN(
        n18783) );
  INV_X1 U21764 ( .A(n18783), .ZN(n18794) );
  NOR2_X1 U21765 ( .A1(n18785), .A2(n18784), .ZN(n18786) );
  XNOR2_X1 U21766 ( .A(n18787), .B(n18786), .ZN(n18792) );
  OAI22_X1 U21767 ( .A1(n18790), .A2(n18812), .B1(n18789), .B2(n18788), .ZN(
        n18791) );
  AOI21_X1 U21768 ( .B1(n18792), .B2(n19499), .A(n18791), .ZN(n18793) );
  OAI211_X1 U21769 ( .C1(n18798), .C2(n10604), .A(n18794), .B(n18793), .ZN(
        P2_U2849) );
  OAI21_X1 U21770 ( .B1(n11072), .B2(n18810), .A(n11181), .ZN(n18800) );
  OAI22_X1 U21771 ( .A1(n18798), .A2(n18797), .B1(n18796), .B2(n18795), .ZN(
        n18799) );
  AOI211_X1 U21772 ( .C1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n9607), .A(
        n18800), .B(n18799), .ZN(n18807) );
  NAND2_X1 U21773 ( .A1(n13264), .A2(n18801), .ZN(n18802) );
  XNOR2_X1 U21774 ( .A(n18803), .B(n18802), .ZN(n18805) );
  AOI22_X1 U21775 ( .A1(n18805), .A2(n19499), .B1(n18814), .B2(n18804), .ZN(
        n18806) );
  OAI211_X1 U21776 ( .C1(n18812), .C2(n18808), .A(n18807), .B(n18806), .ZN(
        P2_U2850) );
  INV_X1 U21777 ( .A(n18809), .ZN(n18811) );
  OAI22_X1 U21778 ( .A1(n18812), .A2(n18811), .B1(n10280), .B2(n18810), .ZN(
        n18813) );
  INV_X1 U21779 ( .A(n18813), .ZN(n18823) );
  NAND2_X1 U21780 ( .A1(n18815), .A2(n18814), .ZN(n18822) );
  INV_X1 U21781 ( .A(n18816), .ZN(n18817) );
  NAND2_X1 U21782 ( .A1(n18818), .A2(n18817), .ZN(n18821) );
  NAND2_X1 U21783 ( .A1(n18819), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n18820) );
  NAND4_X1 U21784 ( .A1(n18823), .A2(n18822), .A3(n18821), .A4(n18820), .ZN(
        n18824) );
  AOI21_X1 U21785 ( .B1(n19261), .B2(n18825), .A(n18824), .ZN(n18829) );
  OAI21_X1 U21786 ( .B1(n9607), .B2(n18826), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18828) );
  OAI211_X1 U21787 ( .C1(n18831), .C2(n18830), .A(n18829), .B(n18828), .ZN(
        P2_U2855) );
  INV_X1 U21788 ( .A(n18832), .ZN(n18833) );
  AOI21_X1 U21789 ( .B1(n18834), .B2(n13474), .A(n18833), .ZN(n18886) );
  AOI22_X1 U21790 ( .A1(n18886), .A2(n18871), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n18875), .ZN(n18835) );
  OAI21_X1 U21791 ( .B1(n18875), .B2(n18836), .A(n18835), .ZN(P2_U2871) );
  AOI21_X1 U21792 ( .B1(n13406), .B2(n18838), .A(n18837), .ZN(n18839) );
  NOR3_X1 U21793 ( .A1(n18840), .A2(n18839), .A3(n18865), .ZN(n18841) );
  AOI21_X1 U21794 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n18875), .A(n18841), .ZN(
        n18842) );
  OAI21_X1 U21795 ( .B1(n18843), .B2(n18875), .A(n18842), .ZN(P2_U2873) );
  INV_X1 U21796 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n18848) );
  AOI21_X1 U21797 ( .B1(n9652), .B2(n18845), .A(n18844), .ZN(n18846) );
  OR3_X1 U21798 ( .A1(n13406), .A2(n18846), .A3(n18865), .ZN(n18847) );
  OAI21_X1 U21799 ( .B1(n18859), .B2(n18848), .A(n18847), .ZN(n18849) );
  INV_X1 U21800 ( .A(n18849), .ZN(n18850) );
  OAI21_X1 U21801 ( .B1(n18851), .B2(n18875), .A(n18850), .ZN(P2_U2875) );
  INV_X1 U21802 ( .A(n18852), .ZN(n18854) );
  AOI211_X1 U21803 ( .C1(n18854), .C2(n18853), .A(n18865), .B(n9652), .ZN(
        n18855) );
  AOI21_X1 U21804 ( .B1(n18856), .B2(n18859), .A(n18855), .ZN(n18857) );
  OAI21_X1 U21805 ( .B1(n18859), .B2(n18858), .A(n18857), .ZN(P2_U2877) );
  INV_X1 U21806 ( .A(n18860), .ZN(n18867) );
  AND2_X1 U21807 ( .A1(n12952), .A2(n18861), .ZN(n18863) );
  NAND2_X1 U21808 ( .A1(n18863), .A2(n18862), .ZN(n18866) );
  AOI211_X1 U21809 ( .C1(n18867), .C2(n18866), .A(n18865), .B(n18864), .ZN(
        n18868) );
  AOI21_X1 U21810 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n18875), .A(n18868), .ZN(
        n18869) );
  OAI21_X1 U21811 ( .B1(n18870), .B2(n18875), .A(n18869), .ZN(P2_U2879) );
  AOI22_X1 U21812 ( .A1(n18872), .A2(n18871), .B1(P2_EBX_REG_4__SCAN_IN), .B2(
        n18875), .ZN(n18873) );
  OAI21_X1 U21813 ( .B1(n18875), .B2(n18874), .A(n18873), .ZN(P2_U2883) );
  AOI22_X1 U21814 ( .A1(n18876), .A2(n18884), .B1(n18881), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n18878) );
  AOI22_X1 U21815 ( .A1(n18882), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n18893), .ZN(n18877) );
  NAND2_X1 U21816 ( .A1(n18878), .A2(n18877), .ZN(P2_U2888) );
  AOI22_X1 U21817 ( .A1(n18880), .A2(n18879), .B1(n18893), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n18889) );
  AOI22_X1 U21818 ( .A1(n18882), .A2(BUF1_REG_16__SCAN_IN), .B1(n18881), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n18888) );
  AOI22_X1 U21819 ( .A1(n18886), .A2(n18885), .B1(n18884), .B2(n18883), .ZN(
        n18887) );
  NAND3_X1 U21820 ( .A1(n18889), .A2(n18888), .A3(n18887), .ZN(P2_U2903) );
  AOI22_X1 U21821 ( .A1(n18895), .A2(n18890), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n18893), .ZN(n18891) );
  OAI21_X1 U21822 ( .B1(n18898), .B2(n18892), .A(n18891), .ZN(P2_U2907) );
  AOI22_X1 U21823 ( .A1(n18895), .A2(n18894), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n18893), .ZN(n18896) );
  OAI21_X1 U21824 ( .B1(n18898), .B2(n18897), .A(n18896), .ZN(P2_U2909) );
  NOR2_X1 U21825 ( .A1(n18923), .A2(n18899), .ZN(P2_U2920) );
  INV_X1 U21826 ( .A(n18921), .ZN(n18932) );
  AOI22_X1 U21827 ( .A1(n18930), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n18900) );
  OAI21_X1 U21828 ( .B1(n12707), .B2(n18932), .A(n18900), .ZN(P2_U2936) );
  AOI22_X1 U21829 ( .A1(n18930), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n18901) );
  OAI21_X1 U21830 ( .B1(n10979), .B2(n18932), .A(n18901), .ZN(P2_U2937) );
  INV_X1 U21831 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n18903) );
  AOI22_X1 U21832 ( .A1(n18904), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n18902) );
  OAI21_X1 U21833 ( .B1(n18903), .B2(n18932), .A(n18902), .ZN(P2_U2938) );
  AOI22_X1 U21834 ( .A1(n18904), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n18905) );
  OAI21_X1 U21835 ( .B1(n18906), .B2(n18932), .A(n18905), .ZN(P2_U2939) );
  AOI22_X1 U21836 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n18927), .B1(n18930), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n18907) );
  OAI21_X1 U21837 ( .B1(n18908), .B2(n18932), .A(n18907), .ZN(P2_U2940) );
  AOI22_X1 U21838 ( .A1(n18930), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n18909) );
  OAI21_X1 U21839 ( .B1(n18910), .B2(n18932), .A(n18909), .ZN(P2_U2941) );
  AOI22_X1 U21840 ( .A1(n18930), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n18911) );
  OAI21_X1 U21841 ( .B1(n18912), .B2(n18932), .A(n18911), .ZN(P2_U2942) );
  AOI22_X1 U21842 ( .A1(n18930), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n18913) );
  OAI21_X1 U21843 ( .B1(n10899), .B2(n18932), .A(n18913), .ZN(P2_U2943) );
  AOI22_X1 U21844 ( .A1(n18930), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n18914) );
  OAI21_X1 U21845 ( .B1(n18915), .B2(n18932), .A(n18914), .ZN(P2_U2944) );
  AOI22_X1 U21846 ( .A1(n18930), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n18916) );
  OAI21_X1 U21847 ( .B1(n18917), .B2(n18932), .A(n18916), .ZN(P2_U2945) );
  INV_X1 U21848 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n18919) );
  AOI22_X1 U21849 ( .A1(n18930), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n18918) );
  OAI21_X1 U21850 ( .B1(n18919), .B2(n18932), .A(n18918), .ZN(P2_U2946) );
  AOI22_X1 U21851 ( .A1(n18930), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n18920) );
  OAI21_X1 U21852 ( .B1(n10885), .B2(n18932), .A(n18920), .ZN(P2_U2947) );
  AOI22_X1 U21853 ( .A1(P2_EAX_REG_3__SCAN_IN), .A2(n18921), .B1(n18930), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n18922) );
  OAI21_X1 U21854 ( .B1(n18924), .B2(n18923), .A(n18922), .ZN(P2_U2948) );
  AOI22_X1 U21855 ( .A1(n18930), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n18925) );
  OAI21_X1 U21856 ( .B1(n18926), .B2(n18932), .A(n18925), .ZN(P2_U2949) );
  AOI22_X1 U21857 ( .A1(n18930), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n18928) );
  OAI21_X1 U21858 ( .B1(n18929), .B2(n18932), .A(n18928), .ZN(P2_U2950) );
  AOI22_X1 U21859 ( .A1(n18930), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n18927), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n18931) );
  OAI21_X1 U21860 ( .B1(n12709), .B2(n18932), .A(n18931), .ZN(P2_U2951) );
  AOI22_X1 U21861 ( .A1(n18934), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n18933), .ZN(n18942) );
  AOI222_X1 U21862 ( .A1(n18940), .A2(n18939), .B1(n18938), .B2(n18937), .C1(
        n18936), .C2(n18935), .ZN(n18941) );
  OAI211_X1 U21863 ( .C1(n18944), .C2(n18943), .A(n18942), .B(n18941), .ZN(
        P2_U3010) );
  INV_X1 U21864 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20760) );
  AOI22_X1 U21865 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18978), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n18979), .ZN(n19453) );
  NOR2_X2 U21866 ( .A1(n10253), .A2(n18980), .ZN(n19442) );
  AOI22_X1 U21867 ( .A1(n19488), .A2(n19388), .B1(n18982), .B2(n19442), .ZN(
        n18950) );
  AOI22_X1 U21868 ( .A1(n18946), .A2(n18988), .B1(n19016), .B2(n19450), .ZN(
        n18949) );
  OAI211_X1 U21869 ( .C1(n18991), .C2(n20760), .A(n18950), .B(n18949), .ZN(
        P2_U3048) );
  INV_X1 U21870 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18957) );
  AOI22_X1 U21871 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n18979), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18978), .ZN(n19458) );
  INV_X1 U21872 ( .A(n19458), .ZN(n19405) );
  NOR2_X2 U21873 ( .A1(n12874), .A2(n18980), .ZN(n19454) );
  AOI22_X1 U21874 ( .A1(n19488), .A2(n19405), .B1(n18982), .B2(n19454), .ZN(
        n18956) );
  AOI22_X1 U21875 ( .A1(n18952), .A2(n18988), .B1(n19016), .B2(n19455), .ZN(
        n18955) );
  OAI211_X1 U21876 ( .C1(n18991), .C2(n18957), .A(n18956), .B(n18955), .ZN(
        P2_U3049) );
  INV_X1 U21877 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18963) );
  AOI22_X1 U21878 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n18979), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18978), .ZN(n19463) );
  INV_X1 U21879 ( .A(n19463), .ZN(n19409) );
  NOR2_X2 U21880 ( .A1(n18958), .A2(n18980), .ZN(n19459) );
  AOI22_X1 U21881 ( .A1(n19488), .A2(n19409), .B1(n18982), .B2(n19459), .ZN(
        n18962) );
  AOI22_X1 U21882 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n18979), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18978), .ZN(n19412) );
  AOI22_X1 U21883 ( .A1(n18960), .A2(n18988), .B1(n19016), .B2(n19460), .ZN(
        n18961) );
  OAI211_X1 U21884 ( .C1(n18991), .C2(n18963), .A(n18962), .B(n18961), .ZN(
        P2_U3050) );
  AOI22_X1 U21885 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n18979), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18978), .ZN(n19468) );
  INV_X1 U21886 ( .A(n19468), .ZN(n19413) );
  INV_X1 U21887 ( .A(n18980), .ZN(n18964) );
  AND2_X1 U21888 ( .A1(n18965), .A2(n18964), .ZN(n19464) );
  AOI22_X1 U21889 ( .A1(n19488), .A2(n19413), .B1(n18982), .B2(n19464), .ZN(
        n18969) );
  AOI22_X1 U21890 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n18979), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18978), .ZN(n19416) );
  AOI22_X1 U21891 ( .A1(n18967), .A2(n18988), .B1(n19016), .B2(n19465), .ZN(
        n18968) );
  OAI211_X1 U21892 ( .C1(n18991), .C2(n18970), .A(n18969), .B(n18968), .ZN(
        P2_U3051) );
  INV_X1 U21893 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18977) );
  AOI22_X1 U21894 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18978), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n18979), .ZN(n19482) );
  NOR2_X2 U21895 ( .A1(n18971), .A2(n18980), .ZN(n19477) );
  AOI22_X1 U21896 ( .A1(n19488), .A2(n19425), .B1(n18982), .B2(n19477), .ZN(
        n18976) );
  NOR2_X2 U21897 ( .A1(n18972), .A2(n19171), .ZN(n19478) );
  AOI22_X1 U21898 ( .A1(n19478), .A2(n18988), .B1(n19016), .B2(n19479), .ZN(
        n18975) );
  OAI211_X1 U21899 ( .C1(n18991), .C2(n18977), .A(n18976), .B(n18975), .ZN(
        P2_U3054) );
  AOI22_X1 U21900 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n18979), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n18978), .ZN(n19493) );
  INV_X1 U21901 ( .A(n19493), .ZN(n19431) );
  NOR2_X2 U21902 ( .A1(n18981), .A2(n18980), .ZN(n19483) );
  AOI22_X1 U21903 ( .A1(n19488), .A2(n19431), .B1(n18982), .B2(n19483), .ZN(
        n18990) );
  NOR2_X2 U21904 ( .A1(n18983), .A2(n19171), .ZN(n19485) );
  AOI22_X1 U21905 ( .A1(n19485), .A2(n18988), .B1(n19016), .B2(n19487), .ZN(
        n18989) );
  OAI211_X1 U21906 ( .C1(n18991), .C2(n11319), .A(n18990), .B(n18989), .ZN(
        P2_U3055) );
  INV_X1 U21907 ( .A(n19023), .ZN(n18995) );
  NAND2_X1 U21908 ( .A1(n19020), .A2(n19603), .ZN(n18997) );
  INV_X1 U21909 ( .A(n18992), .ZN(n19168) );
  NOR2_X1 U21910 ( .A1(n19613), .A2(n18997), .ZN(n19014) );
  NOR3_X1 U21911 ( .A1(n18993), .A2(n19014), .A3(n19606), .ZN(n18996) );
  AOI211_X2 U21912 ( .C1(n18997), .C2(n19606), .A(n19168), .B(n18996), .ZN(
        n19015) );
  AOI22_X1 U21913 ( .A1(n19015), .A2(n18946), .B1(n19442), .B2(n19014), .ZN(
        n19001) );
  OR2_X1 U21914 ( .A1(n19590), .A2(n19294), .ZN(n19227) );
  INV_X1 U21915 ( .A(n19227), .ZN(n18994) );
  NAND2_X1 U21916 ( .A1(n18995), .A2(n18994), .ZN(n18998) );
  AOI21_X1 U21917 ( .B1(n18998), .B2(n18997), .A(n18996), .ZN(n18999) );
  OAI211_X1 U21918 ( .C1(n19014), .C2(n19582), .A(n18999), .B(n19444), .ZN(
        n19017) );
  AOI22_X1 U21919 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19017), .B1(
        n19016), .B2(n19388), .ZN(n19000) );
  OAI211_X1 U21920 ( .C1(n19404), .C2(n20834), .A(n19001), .B(n19000), .ZN(
        P2_U3056) );
  INV_X1 U21921 ( .A(n19455), .ZN(n19408) );
  AOI22_X1 U21922 ( .A1(n19015), .A2(n18952), .B1(n19454), .B2(n19014), .ZN(
        n19003) );
  AOI22_X1 U21923 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19017), .B1(
        n19016), .B2(n19405), .ZN(n19002) );
  OAI211_X1 U21924 ( .C1(n19408), .C2(n20834), .A(n19003), .B(n19002), .ZN(
        P2_U3057) );
  AOI22_X1 U21925 ( .A1(n19015), .A2(n18960), .B1(n19459), .B2(n19014), .ZN(
        n19005) );
  AOI22_X1 U21926 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19017), .B1(
        n19016), .B2(n19409), .ZN(n19004) );
  OAI211_X1 U21927 ( .C1(n19412), .C2(n20834), .A(n19005), .B(n19004), .ZN(
        P2_U3058) );
  AOI22_X1 U21928 ( .A1(n19015), .A2(n18967), .B1(n19464), .B2(n19014), .ZN(
        n19007) );
  AOI22_X1 U21929 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19017), .B1(
        n19016), .B2(n19413), .ZN(n19006) );
  OAI211_X1 U21930 ( .C1(n19416), .C2(n20834), .A(n19007), .B(n19006), .ZN(
        P2_U3059) );
  AOI22_X1 U21931 ( .A1(n19015), .A2(n19470), .B1(n19469), .B2(n19014), .ZN(
        n19009) );
  INV_X1 U21932 ( .A(n19474), .ZN(n19417) );
  AOI22_X1 U21933 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19017), .B1(
        n19016), .B2(n19417), .ZN(n19008) );
  OAI211_X1 U21934 ( .C1(n19420), .C2(n20834), .A(n19009), .B(n19008), .ZN(
        P2_U3060) );
  AOI22_X1 U21935 ( .A1(n19015), .A2(n20827), .B1(n20826), .B2(n19014), .ZN(
        n19011) );
  AOI22_X1 U21936 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19017), .B1(
        n19016), .B2(n19421), .ZN(n19010) );
  OAI211_X1 U21937 ( .C1(n19424), .C2(n20834), .A(n19011), .B(n19010), .ZN(
        P2_U3061) );
  AOI22_X1 U21938 ( .A1(n19015), .A2(n19478), .B1(n19477), .B2(n19014), .ZN(
        n19013) );
  AOI22_X1 U21939 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19017), .B1(
        n19016), .B2(n19425), .ZN(n19012) );
  OAI211_X1 U21940 ( .C1(n19428), .C2(n20834), .A(n19013), .B(n19012), .ZN(
        P2_U3062) );
  AOI22_X1 U21941 ( .A1(n19015), .A2(n19485), .B1(n19483), .B2(n19014), .ZN(
        n19019) );
  AOI22_X1 U21942 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19017), .B1(
        n19016), .B2(n19431), .ZN(n19018) );
  OAI211_X1 U21943 ( .C1(n19436), .C2(n20834), .A(n19019), .B(n19018), .ZN(
        P2_U3063) );
  NAND2_X1 U21944 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19020), .ZN(
        n19051) );
  NOR2_X1 U21945 ( .A1(n19051), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20825) );
  OAI21_X1 U21946 ( .B1(n10468), .B2(n20825), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19022) );
  NOR2_X1 U21947 ( .A1(n19259), .A2(n19044), .ZN(n19024) );
  INV_X1 U21948 ( .A(n19024), .ZN(n19021) );
  NAND2_X1 U21949 ( .A1(n19022), .A2(n19021), .ZN(n20828) );
  AOI22_X1 U21950 ( .A1(n20828), .A2(n18946), .B1(n19442), .B2(n20825), .ZN(
        n19030) );
  AOI21_X1 U21951 ( .B1(n10468), .B2(n19582), .A(n20825), .ZN(n19027) );
  AOI21_X1 U21952 ( .B1(n19072), .B2(n20834), .A(n19294), .ZN(n19025) );
  NOR2_X1 U21953 ( .A1(n19025), .A2(n19024), .ZN(n19026) );
  MUX2_X1 U21954 ( .A(n19027), .B(n19026), .S(n19390), .Z(n19028) );
  AOI22_X1 U21955 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20831), .B1(
        n20830), .B2(n19450), .ZN(n19029) );
  OAI211_X1 U21956 ( .C1(n19453), .C2(n20834), .A(n19030), .B(n19029), .ZN(
        P2_U3064) );
  AOI22_X1 U21957 ( .A1(n20828), .A2(n18952), .B1(n19454), .B2(n20825), .ZN(
        n19032) );
  AOI22_X1 U21958 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20831), .B1(
        n20830), .B2(n19455), .ZN(n19031) );
  OAI211_X1 U21959 ( .C1(n19458), .C2(n20834), .A(n19032), .B(n19031), .ZN(
        P2_U3065) );
  AOI22_X1 U21960 ( .A1(n20828), .A2(n18960), .B1(n19459), .B2(n20825), .ZN(
        n19034) );
  AOI22_X1 U21961 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20831), .B1(
        n20830), .B2(n19460), .ZN(n19033) );
  OAI211_X1 U21962 ( .C1(n19463), .C2(n20834), .A(n19034), .B(n19033), .ZN(
        P2_U3066) );
  AOI22_X1 U21963 ( .A1(n20828), .A2(n18967), .B1(n19464), .B2(n20825), .ZN(
        n19036) );
  AOI22_X1 U21964 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20831), .B1(
        n20830), .B2(n19465), .ZN(n19035) );
  OAI211_X1 U21965 ( .C1(n19468), .C2(n20834), .A(n19036), .B(n19035), .ZN(
        P2_U3067) );
  AOI22_X1 U21966 ( .A1(n20828), .A2(n19470), .B1(n19469), .B2(n20825), .ZN(
        n19038) );
  AOI22_X1 U21967 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20831), .B1(
        n20830), .B2(n19471), .ZN(n19037) );
  OAI211_X1 U21968 ( .C1(n19474), .C2(n20834), .A(n19038), .B(n19037), .ZN(
        P2_U3068) );
  AOI22_X1 U21969 ( .A1(n20828), .A2(n19478), .B1(n19477), .B2(n20825), .ZN(
        n19040) );
  AOI22_X1 U21970 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20831), .B1(
        n20830), .B2(n19479), .ZN(n19039) );
  OAI211_X1 U21971 ( .C1(n19482), .C2(n20834), .A(n19040), .B(n19039), .ZN(
        P2_U3070) );
  AOI22_X1 U21972 ( .A1(n20828), .A2(n19485), .B1(n19483), .B2(n20825), .ZN(
        n19042) );
  AOI22_X1 U21973 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20831), .B1(
        n20830), .B2(n19487), .ZN(n19041) );
  OAI211_X1 U21974 ( .C1(n19493), .C2(n20834), .A(n19042), .B(n19041), .ZN(
        P2_U3071) );
  NOR2_X1 U21975 ( .A1(n19288), .A2(n19044), .ZN(n19067) );
  AOI22_X1 U21976 ( .A1(n20830), .A2(n19388), .B1(n19067), .B2(n19442), .ZN(
        n19054) );
  OAI21_X1 U21977 ( .B1(n19045), .B2(n19294), .A(n19390), .ZN(n19052) );
  INV_X1 U21978 ( .A(n19051), .ZN(n19049) );
  INV_X1 U21979 ( .A(n19067), .ZN(n19046) );
  OAI211_X1 U21980 ( .C1(n19047), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19046), 
        .B(n19393), .ZN(n19048) );
  OAI211_X1 U21981 ( .C1(n19052), .C2(n19049), .A(n19444), .B(n19048), .ZN(
        n19069) );
  OAI21_X1 U21982 ( .B1(n10469), .B2(n19067), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19050) );
  OAI21_X1 U21983 ( .B1(n19052), .B2(n19051), .A(n19050), .ZN(n19068) );
  AOI22_X1 U21984 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19069), .B1(
        n18946), .B2(n19068), .ZN(n19053) );
  OAI211_X1 U21985 ( .C1(n19404), .C2(n19105), .A(n19054), .B(n19053), .ZN(
        P2_U3072) );
  AOI22_X1 U21986 ( .A1(n20830), .A2(n19405), .B1(n19067), .B2(n19454), .ZN(
        n19056) );
  AOI22_X1 U21987 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19069), .B1(
        n18952), .B2(n19068), .ZN(n19055) );
  OAI211_X1 U21988 ( .C1(n19408), .C2(n19105), .A(n19056), .B(n19055), .ZN(
        P2_U3073) );
  AOI22_X1 U21989 ( .A1(n19074), .A2(n19460), .B1(n19067), .B2(n19459), .ZN(
        n19058) );
  AOI22_X1 U21990 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19069), .B1(
        n18960), .B2(n19068), .ZN(n19057) );
  OAI211_X1 U21991 ( .C1(n19463), .C2(n19072), .A(n19058), .B(n19057), .ZN(
        P2_U3074) );
  AOI22_X1 U21992 ( .A1(n19074), .A2(n19465), .B1(n19067), .B2(n19464), .ZN(
        n19060) );
  AOI22_X1 U21993 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19069), .B1(
        n18967), .B2(n19068), .ZN(n19059) );
  OAI211_X1 U21994 ( .C1(n19468), .C2(n19072), .A(n19060), .B(n19059), .ZN(
        P2_U3075) );
  AOI22_X1 U21995 ( .A1(n19074), .A2(n19471), .B1(n19469), .B2(n19067), .ZN(
        n19062) );
  AOI22_X1 U21996 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19069), .B1(
        n19470), .B2(n19068), .ZN(n19061) );
  OAI211_X1 U21997 ( .C1(n19474), .C2(n19072), .A(n19062), .B(n19061), .ZN(
        P2_U3076) );
  AOI22_X1 U21998 ( .A1(n19074), .A2(n20829), .B1(n20826), .B2(n19067), .ZN(
        n19064) );
  AOI22_X1 U21999 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19069), .B1(
        n20827), .B2(n19068), .ZN(n19063) );
  OAI211_X1 U22000 ( .C1(n20835), .C2(n19072), .A(n19064), .B(n19063), .ZN(
        P2_U3077) );
  AOI22_X1 U22001 ( .A1(n19074), .A2(n19479), .B1(n19067), .B2(n19477), .ZN(
        n19066) );
  AOI22_X1 U22002 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19069), .B1(
        n19478), .B2(n19068), .ZN(n19065) );
  OAI211_X1 U22003 ( .C1(n19482), .C2(n19072), .A(n19066), .B(n19065), .ZN(
        P2_U3078) );
  AOI22_X1 U22004 ( .A1(n19074), .A2(n19487), .B1(n19067), .B2(n19483), .ZN(
        n19071) );
  AOI22_X1 U22005 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19069), .B1(
        n19485), .B2(n19068), .ZN(n19070) );
  OAI211_X1 U22006 ( .C1(n19493), .C2(n19072), .A(n19071), .B(n19070), .ZN(
        P2_U3079) );
  NOR2_X1 U22007 ( .A1(n19592), .A2(n19326), .ZN(n19073) );
  NAND2_X1 U22008 ( .A1(n19581), .A2(n19073), .ZN(n19129) );
  NAND3_X1 U22009 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19588), .A3(
        n19603), .ZN(n19111) );
  NOR2_X1 U22010 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19111), .ZN(
        n19100) );
  AOI22_X1 U22011 ( .A1(n19450), .A2(n19134), .B1(n19442), .B2(n19100), .ZN(
        n19087) );
  NOR2_X1 U22012 ( .A1(n19074), .A2(n19134), .ZN(n19075) );
  OAI21_X1 U22013 ( .B1(n19075), .B2(n19294), .A(n19390), .ZN(n19085) );
  INV_X1 U22014 ( .A(n19076), .ZN(n19078) );
  NAND2_X1 U22015 ( .A1(n19288), .A2(n19195), .ZN(n19077) );
  NAND2_X1 U22016 ( .A1(n19078), .A2(n19077), .ZN(n19330) );
  NOR2_X1 U22017 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19330), .ZN(
        n19082) );
  OAI21_X1 U22018 ( .B1(n10474), .B2(n19606), .A(n19582), .ZN(n19080) );
  INV_X1 U22019 ( .A(n19100), .ZN(n19079) );
  AOI21_X1 U22020 ( .B1(n19080), .B2(n19079), .A(n19171), .ZN(n19081) );
  INV_X1 U22021 ( .A(n19082), .ZN(n19084) );
  OAI21_X1 U22022 ( .B1(n10474), .B2(n19100), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19083) );
  AOI22_X1 U22023 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19102), .B1(
        n18946), .B2(n19101), .ZN(n19086) );
  OAI211_X1 U22024 ( .C1(n19453), .C2(n19105), .A(n19087), .B(n19086), .ZN(
        P2_U3080) );
  AOI22_X1 U22025 ( .A1(n19455), .A2(n19134), .B1(n19454), .B2(n19100), .ZN(
        n19089) );
  AOI22_X1 U22026 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19102), .B1(
        n18952), .B2(n19101), .ZN(n19088) );
  OAI211_X1 U22027 ( .C1(n19458), .C2(n19105), .A(n19089), .B(n19088), .ZN(
        P2_U3081) );
  AOI22_X1 U22028 ( .A1(n19460), .A2(n19134), .B1(n19459), .B2(n19100), .ZN(
        n19091) );
  AOI22_X1 U22029 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19102), .B1(
        n18960), .B2(n19101), .ZN(n19090) );
  OAI211_X1 U22030 ( .C1(n19463), .C2(n19105), .A(n19091), .B(n19090), .ZN(
        P2_U3082) );
  AOI22_X1 U22031 ( .A1(n19465), .A2(n19134), .B1(n19464), .B2(n19100), .ZN(
        n19093) );
  AOI22_X1 U22032 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19102), .B1(
        n18967), .B2(n19101), .ZN(n19092) );
  OAI211_X1 U22033 ( .C1(n19468), .C2(n19105), .A(n19093), .B(n19092), .ZN(
        P2_U3083) );
  AOI22_X1 U22034 ( .A1(n19471), .A2(n19134), .B1(n19469), .B2(n19100), .ZN(
        n19095) );
  AOI22_X1 U22035 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19102), .B1(
        n19470), .B2(n19101), .ZN(n19094) );
  OAI211_X1 U22036 ( .C1(n19474), .C2(n19105), .A(n19095), .B(n19094), .ZN(
        P2_U3084) );
  AOI22_X1 U22037 ( .A1(n20829), .A2(n19134), .B1(n20826), .B2(n19100), .ZN(
        n19097) );
  AOI22_X1 U22038 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19102), .B1(
        n20827), .B2(n19101), .ZN(n19096) );
  OAI211_X1 U22039 ( .C1(n20835), .C2(n19105), .A(n19097), .B(n19096), .ZN(
        P2_U3085) );
  AOI22_X1 U22040 ( .A1(n19479), .A2(n19134), .B1(n19477), .B2(n19100), .ZN(
        n19099) );
  AOI22_X1 U22041 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19102), .B1(
        n19478), .B2(n19101), .ZN(n19098) );
  OAI211_X1 U22042 ( .C1(n19482), .C2(n19105), .A(n19099), .B(n19098), .ZN(
        P2_U3086) );
  AOI22_X1 U22043 ( .A1(n19487), .A2(n19134), .B1(n19483), .B2(n19100), .ZN(
        n19104) );
  AOI22_X1 U22044 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19102), .B1(
        n19485), .B2(n19101), .ZN(n19103) );
  OAI211_X1 U22045 ( .C1(n19493), .C2(n19105), .A(n19104), .B(n19103), .ZN(
        P2_U3087) );
  NOR2_X1 U22046 ( .A1(n19613), .A2(n19111), .ZN(n19144) );
  INV_X1 U22047 ( .A(n19144), .ZN(n19106) );
  OAI21_X1 U22048 ( .B1(n10580), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19106), 
        .ZN(n19108) );
  NOR2_X1 U22049 ( .A1(n19592), .A2(n19227), .ZN(n19360) );
  NAND2_X1 U22050 ( .A1(n19581), .A2(n19360), .ZN(n19113) );
  NAND2_X1 U22051 ( .A1(n19113), .A2(n19111), .ZN(n19107) );
  MUX2_X1 U22052 ( .A(n19108), .B(n19107), .S(n19390), .Z(n19109) );
  AND2_X1 U22053 ( .A1(n19109), .A2(n19444), .ZN(n19120) );
  INV_X1 U22054 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n19119) );
  NAND2_X1 U22055 ( .A1(n19194), .A2(n19226), .ZN(n19355) );
  INV_X1 U22056 ( .A(n19355), .ZN(n19110) );
  AOI22_X1 U22057 ( .A1(n19450), .A2(n19163), .B1(n19442), .B2(n9754), .ZN(
        n19118) );
  INV_X1 U22058 ( .A(n19111), .ZN(n19112) );
  NAND3_X1 U22059 ( .A1(n19113), .A2(n19390), .A3(n19112), .ZN(n19116) );
  OAI21_X1 U22060 ( .B1(n19114), .B2(n9754), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19115) );
  NAND2_X1 U22061 ( .A1(n19116), .A2(n19115), .ZN(n19135) );
  AOI22_X1 U22062 ( .A1(n18946), .A2(n19135), .B1(n19134), .B2(n19388), .ZN(
        n19117) );
  OAI211_X1 U22063 ( .C1(n19120), .C2(n19119), .A(n19118), .B(n19117), .ZN(
        P2_U3088) );
  AOI22_X1 U22064 ( .A1(n19455), .A2(n19163), .B1(n19454), .B2(n9754), .ZN(
        n19122) );
  AOI22_X1 U22065 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19136), .B1(
        n18952), .B2(n19135), .ZN(n19121) );
  OAI211_X1 U22066 ( .C1(n19458), .C2(n19129), .A(n19122), .B(n19121), .ZN(
        P2_U3089) );
  AOI22_X1 U22067 ( .A1(n19460), .A2(n19163), .B1(n19459), .B2(n9754), .ZN(
        n19124) );
  AOI22_X1 U22068 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19136), .B1(
        n18960), .B2(n19135), .ZN(n19123) );
  OAI211_X1 U22069 ( .C1(n19463), .C2(n19129), .A(n19124), .B(n19123), .ZN(
        P2_U3090) );
  AOI22_X1 U22070 ( .A1(n19465), .A2(n19163), .B1(n19464), .B2(n9754), .ZN(
        n19126) );
  AOI22_X1 U22071 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19136), .B1(
        n18967), .B2(n19135), .ZN(n19125) );
  OAI211_X1 U22072 ( .C1(n19468), .C2(n19129), .A(n19126), .B(n19125), .ZN(
        P2_U3091) );
  AOI22_X1 U22073 ( .A1(n19471), .A2(n19163), .B1(n19469), .B2(n9754), .ZN(
        n19128) );
  AOI22_X1 U22074 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19136), .B1(
        n19470), .B2(n19135), .ZN(n19127) );
  OAI211_X1 U22075 ( .C1(n19474), .C2(n19129), .A(n19128), .B(n19127), .ZN(
        P2_U3092) );
  AOI22_X1 U22076 ( .A1(n19421), .A2(n19134), .B1(n20826), .B2(n9754), .ZN(
        n19131) );
  AOI22_X1 U22077 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19136), .B1(
        n20827), .B2(n19135), .ZN(n19130) );
  OAI211_X1 U22078 ( .C1(n19424), .C2(n19142), .A(n19131), .B(n19130), .ZN(
        P2_U3093) );
  AOI22_X1 U22079 ( .A1(n19425), .A2(n19134), .B1(n19477), .B2(n9754), .ZN(
        n19133) );
  AOI22_X1 U22080 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19136), .B1(
        n19478), .B2(n19135), .ZN(n19132) );
  OAI211_X1 U22081 ( .C1(n19428), .C2(n19142), .A(n19133), .B(n19132), .ZN(
        P2_U3094) );
  AOI22_X1 U22082 ( .A1(n19431), .A2(n19134), .B1(n19483), .B2(n9754), .ZN(
        n19138) );
  AOI22_X1 U22083 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19136), .B1(
        n19485), .B2(n19135), .ZN(n19137) );
  OAI211_X1 U22084 ( .C1(n19436), .C2(n19142), .A(n19138), .B(n19137), .ZN(
        P2_U3095) );
  NOR2_X1 U22085 ( .A1(n19592), .A2(n19599), .ZN(n19139) );
  NOR2_X1 U22086 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19387), .ZN(
        n19173) );
  INV_X1 U22087 ( .A(n19173), .ZN(n19169) );
  NOR2_X1 U22088 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19169), .ZN(
        n19161) );
  NOR2_X1 U22089 ( .A1(n19161), .A2(n19144), .ZN(n19140) );
  OR2_X1 U22090 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19140), .ZN(n19141) );
  NOR3_X1 U22091 ( .A1(n10461), .A2(n19161), .A3(n19606), .ZN(n19145) );
  AOI21_X1 U22092 ( .B1(n19606), .B2(n19141), .A(n19145), .ZN(n19162) );
  AOI22_X1 U22093 ( .A1(n19162), .A2(n18946), .B1(n19442), .B2(n19161), .ZN(
        n19148) );
  AOI21_X1 U22094 ( .B1(n19188), .B2(n19142), .A(n19294), .ZN(n19143) );
  AOI221_X1 U22095 ( .B1(n19582), .B2(n19144), .C1(n19582), .C2(n19143), .A(
        n19161), .ZN(n19146) );
  AOI22_X1 U22096 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19164), .B1(
        n19163), .B2(n19388), .ZN(n19147) );
  OAI211_X1 U22097 ( .C1(n19404), .C2(n19188), .A(n19148), .B(n19147), .ZN(
        P2_U3096) );
  AOI22_X1 U22098 ( .A1(n19162), .A2(n18952), .B1(n19454), .B2(n19161), .ZN(
        n19150) );
  AOI22_X1 U22099 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19164), .B1(
        n19163), .B2(n19405), .ZN(n19149) );
  OAI211_X1 U22100 ( .C1(n19408), .C2(n19188), .A(n19150), .B(n19149), .ZN(
        P2_U3097) );
  AOI22_X1 U22101 ( .A1(n19162), .A2(n18960), .B1(n19459), .B2(n19161), .ZN(
        n19152) );
  AOI22_X1 U22102 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19164), .B1(
        n19163), .B2(n19409), .ZN(n19151) );
  OAI211_X1 U22103 ( .C1(n19412), .C2(n19188), .A(n19152), .B(n19151), .ZN(
        P2_U3098) );
  AOI22_X1 U22104 ( .A1(n19162), .A2(n18967), .B1(n19464), .B2(n19161), .ZN(
        n19154) );
  AOI22_X1 U22105 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19164), .B1(
        n19163), .B2(n19413), .ZN(n19153) );
  OAI211_X1 U22106 ( .C1(n19416), .C2(n19188), .A(n19154), .B(n19153), .ZN(
        P2_U3099) );
  AOI22_X1 U22107 ( .A1(n19162), .A2(n19470), .B1(n19469), .B2(n19161), .ZN(
        n19156) );
  AOI22_X1 U22108 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19164), .B1(
        n19163), .B2(n19417), .ZN(n19155) );
  OAI211_X1 U22109 ( .C1(n19420), .C2(n19188), .A(n19156), .B(n19155), .ZN(
        P2_U3100) );
  AOI22_X1 U22110 ( .A1(n19162), .A2(n20827), .B1(n20826), .B2(n19161), .ZN(
        n19158) );
  AOI22_X1 U22111 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19164), .B1(
        n19163), .B2(n19421), .ZN(n19157) );
  OAI211_X1 U22112 ( .C1(n19424), .C2(n19188), .A(n19158), .B(n19157), .ZN(
        P2_U3101) );
  AOI22_X1 U22113 ( .A1(n19162), .A2(n19478), .B1(n19477), .B2(n19161), .ZN(
        n19160) );
  AOI22_X1 U22114 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19164), .B1(
        n19163), .B2(n19425), .ZN(n19159) );
  OAI211_X1 U22115 ( .C1(n19428), .C2(n19188), .A(n19160), .B(n19159), .ZN(
        P2_U3102) );
  AOI22_X1 U22116 ( .A1(n19162), .A2(n19485), .B1(n19483), .B2(n19161), .ZN(
        n19166) );
  AOI22_X1 U22117 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19164), .B1(
        n19163), .B2(n19431), .ZN(n19165) );
  OAI211_X1 U22118 ( .C1(n19436), .C2(n19188), .A(n19166), .B(n19165), .ZN(
        P2_U3103) );
  NAND2_X1 U22119 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19173), .ZN(
        n19198) );
  INV_X1 U22120 ( .A(n19198), .ZN(n19201) );
  NOR3_X1 U22121 ( .A1(n19167), .A2(n19201), .A3(n19606), .ZN(n19170) );
  AOI211_X2 U22122 ( .C1(n19169), .C2(n19606), .A(n19168), .B(n19170), .ZN(
        n19189) );
  AOI22_X1 U22123 ( .A1(n19189), .A2(n18946), .B1(n19442), .B2(n19201), .ZN(
        n19175) );
  AOI211_X1 U22124 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19198), .A(n19171), 
        .B(n19170), .ZN(n19172) );
  OAI221_X1 U22125 ( .B1(n19173), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19173), 
        .C2(n19585), .A(n19172), .ZN(n19191) );
  AOI22_X1 U22126 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19191), .B1(
        n19190), .B2(n19388), .ZN(n19174) );
  OAI211_X1 U22127 ( .C1(n19404), .C2(n19217), .A(n19175), .B(n19174), .ZN(
        P2_U3104) );
  AOI22_X1 U22128 ( .A1(n19189), .A2(n18952), .B1(n19454), .B2(n19201), .ZN(
        n19177) );
  AOI22_X1 U22129 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19191), .B1(
        n19221), .B2(n19455), .ZN(n19176) );
  OAI211_X1 U22130 ( .C1(n19458), .C2(n19188), .A(n19177), .B(n19176), .ZN(
        P2_U3105) );
  AOI22_X1 U22131 ( .A1(n19189), .A2(n18960), .B1(n19459), .B2(n19201), .ZN(
        n19179) );
  AOI22_X1 U22132 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19191), .B1(
        n19190), .B2(n19409), .ZN(n19178) );
  OAI211_X1 U22133 ( .C1(n19412), .C2(n19217), .A(n19179), .B(n19178), .ZN(
        P2_U3106) );
  AOI22_X1 U22134 ( .A1(n19189), .A2(n18967), .B1(n19464), .B2(n19201), .ZN(
        n19181) );
  AOI22_X1 U22135 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19191), .B1(
        n19190), .B2(n19413), .ZN(n19180) );
  OAI211_X1 U22136 ( .C1(n19416), .C2(n19217), .A(n19181), .B(n19180), .ZN(
        P2_U3107) );
  AOI22_X1 U22137 ( .A1(n19189), .A2(n19470), .B1(n19469), .B2(n19201), .ZN(
        n19183) );
  AOI22_X1 U22138 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19191), .B1(
        n19221), .B2(n19471), .ZN(n19182) );
  OAI211_X1 U22139 ( .C1(n19474), .C2(n19188), .A(n19183), .B(n19182), .ZN(
        P2_U3108) );
  AOI22_X1 U22140 ( .A1(n19189), .A2(n20827), .B1(n20826), .B2(n19201), .ZN(
        n19185) );
  AOI22_X1 U22141 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19191), .B1(
        n19190), .B2(n19421), .ZN(n19184) );
  OAI211_X1 U22142 ( .C1(n19424), .C2(n19217), .A(n19185), .B(n19184), .ZN(
        P2_U3109) );
  AOI22_X1 U22143 ( .A1(n19189), .A2(n19478), .B1(n19477), .B2(n19201), .ZN(
        n19187) );
  AOI22_X1 U22144 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19191), .B1(
        n19221), .B2(n19479), .ZN(n19186) );
  OAI211_X1 U22145 ( .C1(n19482), .C2(n19188), .A(n19187), .B(n19186), .ZN(
        P2_U3110) );
  AOI22_X1 U22146 ( .A1(n19189), .A2(n19485), .B1(n19483), .B2(n19201), .ZN(
        n19193) );
  AOI22_X1 U22147 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19191), .B1(
        n19190), .B2(n19431), .ZN(n19192) );
  OAI211_X1 U22148 ( .C1(n19436), .C2(n19217), .A(n19193), .B(n19192), .ZN(
        P2_U3111) );
  NAND2_X1 U22149 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19596), .ZN(
        n19289) );
  NOR2_X1 U22150 ( .A1(n19195), .A2(n19289), .ZN(n19220) );
  AOI22_X1 U22151 ( .A1(n19450), .A2(n19249), .B1(n19442), .B2(n19220), .ZN(
        n19206) );
  AOI21_X1 U22152 ( .B1(n19196), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19393), 
        .ZN(n19200) );
  OAI21_X1 U22153 ( .B1(n19202), .B2(n19606), .A(n19582), .ZN(n19197) );
  AOI21_X1 U22154 ( .B1(n19200), .B2(n19198), .A(n19197), .ZN(n19199) );
  OAI21_X1 U22155 ( .B1(n19220), .B2(n19201), .A(n19200), .ZN(n19204) );
  OAI21_X1 U22156 ( .B1(n19202), .B2(n19220), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19203) );
  NAND2_X1 U22157 ( .A1(n19204), .A2(n19203), .ZN(n19222) );
  AOI22_X1 U22158 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19223), .B1(
        n18946), .B2(n19222), .ZN(n19205) );
  OAI211_X1 U22159 ( .C1(n19453), .C2(n19217), .A(n19206), .B(n19205), .ZN(
        P2_U3112) );
  AOI22_X1 U22160 ( .A1(n19455), .A2(n19249), .B1(n19454), .B2(n19220), .ZN(
        n19208) );
  AOI22_X1 U22161 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19223), .B1(
        n18952), .B2(n19222), .ZN(n19207) );
  OAI211_X1 U22162 ( .C1(n19458), .C2(n19217), .A(n19208), .B(n19207), .ZN(
        P2_U3113) );
  AOI22_X1 U22163 ( .A1(n19460), .A2(n19249), .B1(n19459), .B2(n19220), .ZN(
        n19210) );
  AOI22_X1 U22164 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19223), .B1(
        n18960), .B2(n19222), .ZN(n19209) );
  OAI211_X1 U22165 ( .C1(n19463), .C2(n19217), .A(n19210), .B(n19209), .ZN(
        P2_U3114) );
  AOI22_X1 U22166 ( .A1(n19413), .A2(n19221), .B1(n19464), .B2(n19220), .ZN(
        n19212) );
  AOI22_X1 U22167 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19223), .B1(
        n18967), .B2(n19222), .ZN(n19211) );
  OAI211_X1 U22168 ( .C1(n19416), .C2(n19257), .A(n19212), .B(n19211), .ZN(
        P2_U3115) );
  AOI22_X1 U22169 ( .A1(n19417), .A2(n19221), .B1(n19469), .B2(n19220), .ZN(
        n19214) );
  AOI22_X1 U22170 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19223), .B1(
        n19470), .B2(n19222), .ZN(n19213) );
  OAI211_X1 U22171 ( .C1(n19420), .C2(n19257), .A(n19214), .B(n19213), .ZN(
        P2_U3116) );
  AOI22_X1 U22172 ( .A1(n20829), .A2(n19249), .B1(n20826), .B2(n19220), .ZN(
        n19216) );
  AOI22_X1 U22173 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19223), .B1(
        n20827), .B2(n19222), .ZN(n19215) );
  OAI211_X1 U22174 ( .C1(n20835), .C2(n19217), .A(n19216), .B(n19215), .ZN(
        P2_U3117) );
  AOI22_X1 U22175 ( .A1(n19221), .A2(n19425), .B1(n19477), .B2(n19220), .ZN(
        n19219) );
  AOI22_X1 U22176 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19223), .B1(
        n19478), .B2(n19222), .ZN(n19218) );
  OAI211_X1 U22177 ( .C1(n19428), .C2(n19257), .A(n19219), .B(n19218), .ZN(
        P2_U3118) );
  AOI22_X1 U22178 ( .A1(n19431), .A2(n19221), .B1(n19483), .B2(n19220), .ZN(
        n19225) );
  AOI22_X1 U22179 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19223), .B1(
        n19485), .B2(n19222), .ZN(n19224) );
  OAI211_X1 U22180 ( .C1(n19436), .C2(n19257), .A(n19225), .B(n19224), .ZN(
        P2_U3119) );
  NOR3_X2 U22181 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19613), .A3(
        n19289), .ZN(n19263) );
  AOI22_X1 U22182 ( .A1(n19249), .A2(n19388), .B1(n19442), .B2(n19263), .ZN(
        n19238) );
  OAI21_X1 U22183 ( .B1(n19228), .B2(n19227), .A(n19390), .ZN(n19236) );
  NOR2_X1 U22184 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19289), .ZN(
        n19232) );
  INV_X1 U22185 ( .A(n19233), .ZN(n19230) );
  INV_X1 U22186 ( .A(n19263), .ZN(n19229) );
  OAI211_X1 U22187 ( .C1(n19230), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19229), 
        .B(n19393), .ZN(n19231) );
  OAI211_X1 U22188 ( .C1(n19236), .C2(n19232), .A(n19444), .B(n19231), .ZN(
        n19254) );
  INV_X1 U22189 ( .A(n19232), .ZN(n19235) );
  OAI21_X1 U22190 ( .B1(n19233), .B2(n19263), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19234) );
  OAI21_X1 U22191 ( .B1(n19236), .B2(n19235), .A(n19234), .ZN(n19253) );
  AOI22_X1 U22192 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19254), .B1(
        n18946), .B2(n19253), .ZN(n19237) );
  OAI211_X1 U22193 ( .C1(n19404), .C2(n19287), .A(n19238), .B(n19237), .ZN(
        P2_U3120) );
  AOI22_X1 U22194 ( .A1(n19405), .A2(n19249), .B1(n19454), .B2(n19263), .ZN(
        n19240) );
  AOI22_X1 U22195 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19254), .B1(
        n18952), .B2(n19253), .ZN(n19239) );
  OAI211_X1 U22196 ( .C1(n19408), .C2(n19287), .A(n19240), .B(n19239), .ZN(
        P2_U3121) );
  AOI22_X1 U22197 ( .A1(n19409), .A2(n19249), .B1(n19459), .B2(n19263), .ZN(
        n19242) );
  AOI22_X1 U22198 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19254), .B1(
        n18960), .B2(n19253), .ZN(n19241) );
  OAI211_X1 U22199 ( .C1(n19412), .C2(n19287), .A(n19242), .B(n19241), .ZN(
        P2_U3122) );
  INV_X1 U22200 ( .A(n19287), .ZN(n19252) );
  AOI22_X1 U22201 ( .A1(n19252), .A2(n19465), .B1(n19464), .B2(n19263), .ZN(
        n19244) );
  AOI22_X1 U22202 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19254), .B1(
        n18967), .B2(n19253), .ZN(n19243) );
  OAI211_X1 U22203 ( .C1(n19468), .C2(n19257), .A(n19244), .B(n19243), .ZN(
        P2_U3123) );
  AOI22_X1 U22204 ( .A1(n19417), .A2(n19249), .B1(n19469), .B2(n19263), .ZN(
        n19246) );
  AOI22_X1 U22205 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19254), .B1(
        n19470), .B2(n19253), .ZN(n19245) );
  OAI211_X1 U22206 ( .C1(n19420), .C2(n19287), .A(n19246), .B(n19245), .ZN(
        P2_U3124) );
  AOI22_X1 U22207 ( .A1(n20829), .A2(n19252), .B1(n20826), .B2(n19263), .ZN(
        n19248) );
  AOI22_X1 U22208 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19254), .B1(
        n20827), .B2(n19253), .ZN(n19247) );
  OAI211_X1 U22209 ( .C1(n20835), .C2(n19257), .A(n19248), .B(n19247), .ZN(
        P2_U3125) );
  AOI22_X1 U22210 ( .A1(n19249), .A2(n19425), .B1(n19477), .B2(n19263), .ZN(
        n19251) );
  AOI22_X1 U22211 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19254), .B1(
        n19478), .B2(n19253), .ZN(n19250) );
  OAI211_X1 U22212 ( .C1(n19428), .C2(n19287), .A(n19251), .B(n19250), .ZN(
        P2_U3126) );
  AOI22_X1 U22213 ( .A1(n19487), .A2(n19252), .B1(n19483), .B2(n19263), .ZN(
        n19256) );
  AOI22_X1 U22214 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19254), .B1(
        n19485), .B2(n19253), .ZN(n19255) );
  OAI211_X1 U22215 ( .C1(n19493), .C2(n19257), .A(n19256), .B(n19255), .ZN(
        P2_U3127) );
  NOR3_X2 U22216 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19603), .A3(
        n19289), .ZN(n19282) );
  OAI21_X1 U22217 ( .B1(n19260), .B2(n19282), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19258) );
  OAI21_X1 U22218 ( .B1(n19289), .B2(n19259), .A(n19258), .ZN(n19283) );
  AOI22_X1 U22219 ( .A1(n19283), .A2(n18946), .B1(n19442), .B2(n19282), .ZN(
        n19269) );
  INV_X1 U22220 ( .A(n19260), .ZN(n19266) );
  INV_X1 U22221 ( .A(n19318), .ZN(n19262) );
  NAND2_X1 U22222 ( .A1(n19262), .A2(n19287), .ZN(n19264) );
  AOI21_X1 U22223 ( .B1(n19264), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19263), 
        .ZN(n19265) );
  AOI211_X1 U22224 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19266), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19265), .ZN(n19267) );
  AOI22_X1 U22225 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19284), .B1(
        n19318), .B2(n19450), .ZN(n19268) );
  OAI211_X1 U22226 ( .C1(n19453), .C2(n19287), .A(n19269), .B(n19268), .ZN(
        P2_U3128) );
  AOI22_X1 U22227 ( .A1(n19283), .A2(n18952), .B1(n19454), .B2(n19282), .ZN(
        n19271) );
  AOI22_X1 U22228 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19284), .B1(
        n19318), .B2(n19455), .ZN(n19270) );
  OAI211_X1 U22229 ( .C1(n19458), .C2(n19287), .A(n19271), .B(n19270), .ZN(
        P2_U3129) );
  AOI22_X1 U22230 ( .A1(n19283), .A2(n18960), .B1(n19459), .B2(n19282), .ZN(
        n19273) );
  AOI22_X1 U22231 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19284), .B1(
        n19318), .B2(n19460), .ZN(n19272) );
  OAI211_X1 U22232 ( .C1(n19463), .C2(n19287), .A(n19273), .B(n19272), .ZN(
        P2_U3130) );
  AOI22_X1 U22233 ( .A1(n19283), .A2(n18967), .B1(n19464), .B2(n19282), .ZN(
        n19275) );
  AOI22_X1 U22234 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19284), .B1(
        n19318), .B2(n19465), .ZN(n19274) );
  OAI211_X1 U22235 ( .C1(n19468), .C2(n19287), .A(n19275), .B(n19274), .ZN(
        P2_U3131) );
  AOI22_X1 U22236 ( .A1(n19283), .A2(n19470), .B1(n19469), .B2(n19282), .ZN(
        n19277) );
  AOI22_X1 U22237 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19284), .B1(
        n19318), .B2(n19471), .ZN(n19276) );
  OAI211_X1 U22238 ( .C1(n19474), .C2(n19287), .A(n19277), .B(n19276), .ZN(
        P2_U3132) );
  AOI22_X1 U22239 ( .A1(n19283), .A2(n20827), .B1(n20826), .B2(n19282), .ZN(
        n19279) );
  AOI22_X1 U22240 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19284), .B1(
        n19318), .B2(n20829), .ZN(n19278) );
  OAI211_X1 U22241 ( .C1(n20835), .C2(n19287), .A(n19279), .B(n19278), .ZN(
        P2_U3133) );
  AOI22_X1 U22242 ( .A1(n19283), .A2(n19478), .B1(n19477), .B2(n19282), .ZN(
        n19281) );
  AOI22_X1 U22243 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19284), .B1(
        n19318), .B2(n19479), .ZN(n19280) );
  OAI211_X1 U22244 ( .C1(n19482), .C2(n19287), .A(n19281), .B(n19280), .ZN(
        P2_U3134) );
  AOI22_X1 U22245 ( .A1(n19283), .A2(n19485), .B1(n19483), .B2(n19282), .ZN(
        n19286) );
  AOI22_X1 U22246 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19284), .B1(
        n19318), .B2(n19487), .ZN(n19285) );
  OAI211_X1 U22247 ( .C1(n19493), .C2(n19287), .A(n19286), .B(n19285), .ZN(
        P2_U3135) );
  NOR2_X1 U22248 ( .A1(n19603), .A2(n19289), .ZN(n19300) );
  INV_X1 U22249 ( .A(n19300), .ZN(n19293) );
  INV_X1 U22250 ( .A(n19288), .ZN(n19291) );
  INV_X1 U22251 ( .A(n19289), .ZN(n19290) );
  NAND2_X1 U22252 ( .A1(n19291), .A2(n19290), .ZN(n19297) );
  INV_X1 U22253 ( .A(n19297), .ZN(n19316) );
  OAI21_X1 U22254 ( .B1(n19296), .B2(n19316), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19292) );
  OAI21_X1 U22255 ( .B1(n19293), .B2(n19393), .A(n19292), .ZN(n19317) );
  AOI22_X1 U22256 ( .A1(n19317), .A2(n18946), .B1(n19442), .B2(n19316), .ZN(
        n19303) );
  NOR2_X1 U22257 ( .A1(n19295), .A2(n19294), .ZN(n19301) );
  INV_X1 U22258 ( .A(n19296), .ZN(n19298) );
  OAI211_X1 U22259 ( .C1(n19298), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19297), 
        .B(n19393), .ZN(n19299) );
  OAI211_X1 U22260 ( .C1(n19301), .C2(n19300), .A(n19444), .B(n19299), .ZN(
        n19319) );
  AOI22_X1 U22261 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19319), .B1(
        n19318), .B2(n19388), .ZN(n19302) );
  OAI211_X1 U22262 ( .C1(n19404), .C2(n19354), .A(n19303), .B(n19302), .ZN(
        P2_U3136) );
  AOI22_X1 U22263 ( .A1(n19317), .A2(n18952), .B1(n19454), .B2(n19316), .ZN(
        n19305) );
  AOI22_X1 U22264 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19319), .B1(
        n19318), .B2(n19405), .ZN(n19304) );
  OAI211_X1 U22265 ( .C1(n19408), .C2(n19354), .A(n19305), .B(n19304), .ZN(
        P2_U3137) );
  AOI22_X1 U22266 ( .A1(n19317), .A2(n18960), .B1(n19459), .B2(n19316), .ZN(
        n19307) );
  AOI22_X1 U22267 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19319), .B1(
        n19318), .B2(n19409), .ZN(n19306) );
  OAI211_X1 U22268 ( .C1(n19412), .C2(n19354), .A(n19307), .B(n19306), .ZN(
        P2_U3138) );
  AOI22_X1 U22269 ( .A1(n19317), .A2(n18967), .B1(n19464), .B2(n19316), .ZN(
        n19309) );
  AOI22_X1 U22270 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19319), .B1(
        n19318), .B2(n19413), .ZN(n19308) );
  OAI211_X1 U22271 ( .C1(n19416), .C2(n19354), .A(n19309), .B(n19308), .ZN(
        P2_U3139) );
  AOI22_X1 U22272 ( .A1(n19317), .A2(n19470), .B1(n19469), .B2(n19316), .ZN(
        n19311) );
  AOI22_X1 U22273 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19319), .B1(
        n19318), .B2(n19417), .ZN(n19310) );
  OAI211_X1 U22274 ( .C1(n19420), .C2(n19354), .A(n19311), .B(n19310), .ZN(
        P2_U3140) );
  AOI22_X1 U22275 ( .A1(n19317), .A2(n20827), .B1(n20826), .B2(n19316), .ZN(
        n19313) );
  AOI22_X1 U22276 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19319), .B1(
        n19318), .B2(n19421), .ZN(n19312) );
  OAI211_X1 U22277 ( .C1(n19424), .C2(n19354), .A(n19313), .B(n19312), .ZN(
        P2_U3141) );
  AOI22_X1 U22278 ( .A1(n19317), .A2(n19478), .B1(n19477), .B2(n19316), .ZN(
        n19315) );
  AOI22_X1 U22279 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19319), .B1(
        n19318), .B2(n19425), .ZN(n19314) );
  OAI211_X1 U22280 ( .C1(n19428), .C2(n19354), .A(n19315), .B(n19314), .ZN(
        P2_U3142) );
  AOI22_X1 U22281 ( .A1(n19317), .A2(n19485), .B1(n19483), .B2(n19316), .ZN(
        n19321) );
  AOI22_X1 U22282 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19319), .B1(
        n19318), .B2(n19431), .ZN(n19320) );
  OAI211_X1 U22283 ( .C1(n19436), .C2(n19354), .A(n19321), .B(n19320), .ZN(
        P2_U3143) );
  INV_X1 U22284 ( .A(n19322), .ZN(n19325) );
  NOR3_X1 U22285 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19596), .A3(
        n19588), .ZN(n19356) );
  INV_X1 U22286 ( .A(n19356), .ZN(n19361) );
  NOR2_X1 U22287 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19361), .ZN(
        n19349) );
  OAI21_X1 U22288 ( .B1(n19323), .B2(n19349), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19324) );
  OAI21_X1 U22289 ( .B1(n19325), .B2(n19330), .A(n19324), .ZN(n19350) );
  AOI22_X1 U22290 ( .A1(n19350), .A2(n18946), .B1(n19442), .B2(n19349), .ZN(
        n19336) );
  INV_X1 U22291 ( .A(n19354), .ZN(n19328) );
  NOR2_X2 U22292 ( .A1(n19327), .A2(n19326), .ZN(n19382) );
  OAI21_X1 U22293 ( .B1(n19328), .B2(n19382), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19329) );
  OAI21_X1 U22294 ( .B1(n19330), .B2(n19588), .A(n19329), .ZN(n19334) );
  INV_X1 U22295 ( .A(n19349), .ZN(n19331) );
  OAI211_X1 U22296 ( .C1(n19332), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19331), 
        .B(n19393), .ZN(n19333) );
  NAND3_X1 U22297 ( .A1(n19334), .A2(n19444), .A3(n19333), .ZN(n19351) );
  AOI22_X1 U22298 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19351), .B1(
        n19382), .B2(n19450), .ZN(n19335) );
  OAI211_X1 U22299 ( .C1(n19453), .C2(n19354), .A(n19336), .B(n19335), .ZN(
        P2_U3144) );
  AOI22_X1 U22300 ( .A1(n19350), .A2(n18952), .B1(n19454), .B2(n19349), .ZN(
        n19338) );
  AOI22_X1 U22301 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19351), .B1(
        n19382), .B2(n19455), .ZN(n19337) );
  OAI211_X1 U22302 ( .C1(n19458), .C2(n19354), .A(n19338), .B(n19337), .ZN(
        P2_U3145) );
  AOI22_X1 U22303 ( .A1(n19350), .A2(n18960), .B1(n19459), .B2(n19349), .ZN(
        n19340) );
  AOI22_X1 U22304 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19351), .B1(
        n19382), .B2(n19460), .ZN(n19339) );
  OAI211_X1 U22305 ( .C1(n19463), .C2(n19354), .A(n19340), .B(n19339), .ZN(
        P2_U3146) );
  AOI22_X1 U22306 ( .A1(n19350), .A2(n18967), .B1(n19464), .B2(n19349), .ZN(
        n19342) );
  AOI22_X1 U22307 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19351), .B1(
        n19382), .B2(n19465), .ZN(n19341) );
  OAI211_X1 U22308 ( .C1(n19468), .C2(n19354), .A(n19342), .B(n19341), .ZN(
        P2_U3147) );
  AOI22_X1 U22309 ( .A1(n19350), .A2(n19470), .B1(n19469), .B2(n19349), .ZN(
        n19344) );
  AOI22_X1 U22310 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19351), .B1(
        n19382), .B2(n19471), .ZN(n19343) );
  OAI211_X1 U22311 ( .C1(n19474), .C2(n19354), .A(n19344), .B(n19343), .ZN(
        P2_U3148) );
  AOI22_X1 U22312 ( .A1(n19350), .A2(n20827), .B1(n20826), .B2(n19349), .ZN(
        n19346) );
  AOI22_X1 U22313 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19351), .B1(
        n19382), .B2(n20829), .ZN(n19345) );
  OAI211_X1 U22314 ( .C1(n20835), .C2(n19354), .A(n19346), .B(n19345), .ZN(
        P2_U3149) );
  AOI22_X1 U22315 ( .A1(n19350), .A2(n19478), .B1(n19477), .B2(n19349), .ZN(
        n19348) );
  AOI22_X1 U22316 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19351), .B1(
        n19382), .B2(n19479), .ZN(n19347) );
  OAI211_X1 U22317 ( .C1(n19482), .C2(n19354), .A(n19348), .B(n19347), .ZN(
        P2_U3150) );
  AOI22_X1 U22318 ( .A1(n19350), .A2(n19485), .B1(n19483), .B2(n19349), .ZN(
        n19353) );
  AOI22_X1 U22319 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19351), .B1(
        n19382), .B2(n19487), .ZN(n19352) );
  OAI211_X1 U22320 ( .C1(n19493), .C2(n19354), .A(n19353), .B(n19352), .ZN(
        P2_U3151) );
  NAND2_X1 U22321 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19356), .ZN(
        n19363) );
  AND2_X1 U22322 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19363), .ZN(n19357) );
  NAND2_X1 U22323 ( .A1(n19358), .A2(n19357), .ZN(n19365) );
  OAI21_X1 U22324 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19361), .A(n19606), 
        .ZN(n19359) );
  AND2_X1 U22325 ( .A1(n19365), .A2(n19359), .ZN(n19381) );
  INV_X1 U22326 ( .A(n19363), .ZN(n19392) );
  AOI22_X1 U22327 ( .A1(n19381), .A2(n18946), .B1(n19442), .B2(n19392), .ZN(
        n19368) );
  INV_X1 U22328 ( .A(n19360), .ZN(n19362) );
  OAI21_X1 U22329 ( .B1(n19362), .B2(n19581), .A(n19361), .ZN(n19366) );
  NAND2_X1 U22330 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19363), .ZN(n19364) );
  NAND4_X1 U22331 ( .A1(n19366), .A2(n19444), .A3(n19365), .A4(n19364), .ZN(
        n19383) );
  AOI22_X1 U22332 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19383), .B1(
        n19382), .B2(n19388), .ZN(n19367) );
  OAI211_X1 U22333 ( .C1(n19404), .C2(n19386), .A(n19368), .B(n19367), .ZN(
        P2_U3152) );
  AOI22_X1 U22334 ( .A1(n19381), .A2(n18952), .B1(n19454), .B2(n19392), .ZN(
        n19370) );
  AOI22_X1 U22335 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19383), .B1(
        n19382), .B2(n19405), .ZN(n19369) );
  OAI211_X1 U22336 ( .C1(n19408), .C2(n19386), .A(n19370), .B(n19369), .ZN(
        P2_U3153) );
  AOI22_X1 U22337 ( .A1(n19381), .A2(n18960), .B1(n19459), .B2(n19392), .ZN(
        n19372) );
  AOI22_X1 U22338 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19383), .B1(
        n19382), .B2(n19409), .ZN(n19371) );
  OAI211_X1 U22339 ( .C1(n19412), .C2(n19386), .A(n19372), .B(n19371), .ZN(
        P2_U3154) );
  AOI22_X1 U22340 ( .A1(n19381), .A2(n18967), .B1(n19464), .B2(n19392), .ZN(
        n19374) );
  AOI22_X1 U22341 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19383), .B1(
        n19382), .B2(n19413), .ZN(n19373) );
  OAI211_X1 U22342 ( .C1(n19416), .C2(n19386), .A(n19374), .B(n19373), .ZN(
        P2_U3155) );
  AOI22_X1 U22343 ( .A1(n19381), .A2(n19470), .B1(n19469), .B2(n19392), .ZN(
        n19376) );
  AOI22_X1 U22344 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19383), .B1(
        n19382), .B2(n19417), .ZN(n19375) );
  OAI211_X1 U22345 ( .C1(n19420), .C2(n19386), .A(n19376), .B(n19375), .ZN(
        P2_U3156) );
  AOI22_X1 U22346 ( .A1(n19381), .A2(n20827), .B1(n20826), .B2(n19392), .ZN(
        n19378) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19383), .B1(
        n19382), .B2(n19421), .ZN(n19377) );
  OAI211_X1 U22348 ( .C1(n19424), .C2(n19386), .A(n19378), .B(n19377), .ZN(
        P2_U3157) );
  AOI22_X1 U22349 ( .A1(n19381), .A2(n19478), .B1(n19477), .B2(n19392), .ZN(
        n19380) );
  AOI22_X1 U22350 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19383), .B1(
        n19382), .B2(n19425), .ZN(n19379) );
  OAI211_X1 U22351 ( .C1(n19428), .C2(n19386), .A(n19380), .B(n19379), .ZN(
        P2_U3158) );
  AOI22_X1 U22352 ( .A1(n19381), .A2(n19485), .B1(n19483), .B2(n19392), .ZN(
        n19385) );
  AOI22_X1 U22353 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19383), .B1(
        n19382), .B2(n19431), .ZN(n19384) );
  OAI211_X1 U22354 ( .C1(n19436), .C2(n19386), .A(n19385), .B(n19384), .ZN(
        P2_U3159) );
  NOR3_X2 U22355 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19588), .A3(
        n19387), .ZN(n19429) );
  AOI22_X1 U22356 ( .A1(n19388), .A2(n19430), .B1(n19442), .B2(n19429), .ZN(
        n19403) );
  INV_X1 U22357 ( .A(n19492), .ZN(n19389) );
  NOR2_X1 U22358 ( .A1(n19389), .A2(n19430), .ZN(n19391) );
  OAI21_X1 U22359 ( .B1(n19391), .B2(n19294), .A(n19390), .ZN(n19401) );
  NOR2_X1 U22360 ( .A1(n19429), .A2(n19392), .ZN(n19400) );
  INV_X1 U22361 ( .A(n19400), .ZN(n19396) );
  INV_X1 U22362 ( .A(n19429), .ZN(n19394) );
  OAI211_X1 U22363 ( .C1(n19397), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19394), 
        .B(n19393), .ZN(n19395) );
  OAI211_X1 U22364 ( .C1(n19401), .C2(n19396), .A(n19444), .B(n19395), .ZN(
        n19433) );
  INV_X1 U22365 ( .A(n19397), .ZN(n19398) );
  OAI21_X1 U22366 ( .B1(n19398), .B2(n19429), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19399) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19433), .B1(
        n18946), .B2(n19432), .ZN(n19402) );
  OAI211_X1 U22368 ( .C1(n19404), .C2(n19492), .A(n19403), .B(n19402), .ZN(
        P2_U3160) );
  AOI22_X1 U22369 ( .A1(n19405), .A2(n19430), .B1(n19454), .B2(n19429), .ZN(
        n19407) );
  AOI22_X1 U22370 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19433), .B1(
        n18952), .B2(n19432), .ZN(n19406) );
  OAI211_X1 U22371 ( .C1(n19408), .C2(n19492), .A(n19407), .B(n19406), .ZN(
        P2_U3161) );
  AOI22_X1 U22372 ( .A1(n19409), .A2(n19430), .B1(n19459), .B2(n19429), .ZN(
        n19411) );
  AOI22_X1 U22373 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19433), .B1(
        n18960), .B2(n19432), .ZN(n19410) );
  OAI211_X1 U22374 ( .C1(n19412), .C2(n19492), .A(n19411), .B(n19410), .ZN(
        P2_U3162) );
  AOI22_X1 U22375 ( .A1(n19413), .A2(n19430), .B1(n19464), .B2(n19429), .ZN(
        n19415) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19433), .B1(
        n18967), .B2(n19432), .ZN(n19414) );
  OAI211_X1 U22377 ( .C1(n19416), .C2(n19492), .A(n19415), .B(n19414), .ZN(
        P2_U3163) );
  AOI22_X1 U22378 ( .A1(n19417), .A2(n19430), .B1(n19469), .B2(n19429), .ZN(
        n19419) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19433), .B1(
        n19470), .B2(n19432), .ZN(n19418) );
  OAI211_X1 U22380 ( .C1(n19420), .C2(n19492), .A(n19419), .B(n19418), .ZN(
        P2_U3164) );
  AOI22_X1 U22381 ( .A1(n19421), .A2(n19430), .B1(n20826), .B2(n19429), .ZN(
        n19423) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19433), .B1(
        n20827), .B2(n19432), .ZN(n19422) );
  OAI211_X1 U22383 ( .C1(n19424), .C2(n19492), .A(n19423), .B(n19422), .ZN(
        P2_U3165) );
  AOI22_X1 U22384 ( .A1(n19425), .A2(n19430), .B1(n19477), .B2(n19429), .ZN(
        n19427) );
  AOI22_X1 U22385 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19433), .B1(
        n19478), .B2(n19432), .ZN(n19426) );
  OAI211_X1 U22386 ( .C1(n19428), .C2(n19492), .A(n19427), .B(n19426), .ZN(
        P2_U3166) );
  AOI22_X1 U22387 ( .A1(n19431), .A2(n19430), .B1(n19483), .B2(n19429), .ZN(
        n19435) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19433), .B1(
        n19485), .B2(n19432), .ZN(n19434) );
  OAI211_X1 U22389 ( .C1(n19436), .C2(n19492), .A(n19435), .B(n19434), .ZN(
        P2_U3167) );
  NAND2_X1 U22390 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19437), .ZN(
        n19443) );
  OR2_X1 U22391 ( .A1(n19443), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19440) );
  NAND2_X1 U22392 ( .A1(n19441), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19438) );
  NOR2_X1 U22393 ( .A1(n19439), .A2(n19438), .ZN(n19446) );
  AOI21_X1 U22394 ( .B1(n19606), .B2(n19440), .A(n19446), .ZN(n19486) );
  INV_X1 U22395 ( .A(n19441), .ZN(n19484) );
  AOI22_X1 U22396 ( .A1(n19486), .A2(n18946), .B1(n19484), .B2(n19442), .ZN(
        n19452) );
  INV_X1 U22397 ( .A(n19443), .ZN(n19449) );
  OAI21_X1 U22398 ( .B1(n19484), .B2(n19582), .A(n19444), .ZN(n19445) );
  NOR2_X1 U22399 ( .A1(n19446), .A2(n19445), .ZN(n19447) );
  OAI221_X1 U22400 ( .B1(n19449), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19449), 
        .C2(n19448), .A(n19447), .ZN(n19489) );
  AOI22_X1 U22401 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19489), .B1(
        n19488), .B2(n19450), .ZN(n19451) );
  OAI211_X1 U22402 ( .C1(n19453), .C2(n19492), .A(n19452), .B(n19451), .ZN(
        P2_U3168) );
  AOI22_X1 U22403 ( .A1(n19486), .A2(n18952), .B1(n19484), .B2(n19454), .ZN(
        n19457) );
  AOI22_X1 U22404 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19489), .B1(
        n19488), .B2(n19455), .ZN(n19456) );
  OAI211_X1 U22405 ( .C1(n19458), .C2(n19492), .A(n19457), .B(n19456), .ZN(
        P2_U3169) );
  AOI22_X1 U22406 ( .A1(n19486), .A2(n18960), .B1(n19484), .B2(n19459), .ZN(
        n19462) );
  AOI22_X1 U22407 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19489), .B1(
        n19488), .B2(n19460), .ZN(n19461) );
  OAI211_X1 U22408 ( .C1(n19463), .C2(n19492), .A(n19462), .B(n19461), .ZN(
        P2_U3170) );
  AOI22_X1 U22409 ( .A1(n19486), .A2(n18967), .B1(n19484), .B2(n19464), .ZN(
        n19467) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19489), .B1(
        n19488), .B2(n19465), .ZN(n19466) );
  OAI211_X1 U22411 ( .C1(n19468), .C2(n19492), .A(n19467), .B(n19466), .ZN(
        P2_U3171) );
  AOI22_X1 U22412 ( .A1(n19486), .A2(n19470), .B1(n19484), .B2(n19469), .ZN(
        n19473) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19489), .B1(
        n19488), .B2(n19471), .ZN(n19472) );
  OAI211_X1 U22414 ( .C1(n19474), .C2(n19492), .A(n19473), .B(n19472), .ZN(
        P2_U3172) );
  AOI22_X1 U22415 ( .A1(n19486), .A2(n20827), .B1(n19484), .B2(n20826), .ZN(
        n19476) );
  AOI22_X1 U22416 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19489), .B1(
        n19488), .B2(n20829), .ZN(n19475) );
  OAI211_X1 U22417 ( .C1(n20835), .C2(n19492), .A(n19476), .B(n19475), .ZN(
        P2_U3173) );
  AOI22_X1 U22418 ( .A1(n19486), .A2(n19478), .B1(n19484), .B2(n19477), .ZN(
        n19481) );
  AOI22_X1 U22419 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19489), .B1(
        n19488), .B2(n19479), .ZN(n19480) );
  OAI211_X1 U22420 ( .C1(n19482), .C2(n19492), .A(n19481), .B(n19480), .ZN(
        P2_U3174) );
  AOI22_X1 U22421 ( .A1(n19486), .A2(n19485), .B1(n19484), .B2(n19483), .ZN(
        n19491) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19489), .B1(
        n19488), .B2(n19487), .ZN(n19490) );
  OAI211_X1 U22423 ( .C1(n19493), .C2(n19492), .A(n19491), .B(n19490), .ZN(
        P2_U3175) );
  OAI21_X1 U22424 ( .B1(n19496), .B2(n19495), .A(n19494), .ZN(n19501) );
  AOI211_X1 U22425 ( .C1(n19497), .C2(n19500), .A(n19504), .B(n11065), .ZN(
        n19498) );
  AOI211_X1 U22426 ( .C1(n19501), .C2(n19500), .A(n19499), .B(n19498), .ZN(
        n19502) );
  INV_X1 U22427 ( .A(n19502), .ZN(P2_U3177) );
  AND2_X1 U22428 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19503), .ZN(
        P2_U3179) );
  AND2_X1 U22429 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19503), .ZN(
        P2_U3180) );
  AND2_X1 U22430 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19503), .ZN(
        P2_U3181) );
  AND2_X1 U22431 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19503), .ZN(
        P2_U3182) );
  AND2_X1 U22432 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19503), .ZN(
        P2_U3183) );
  AND2_X1 U22433 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19503), .ZN(
        P2_U3184) );
  AND2_X1 U22434 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19503), .ZN(
        P2_U3185) );
  AND2_X1 U22435 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19503), .ZN(
        P2_U3186) );
  AND2_X1 U22436 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19503), .ZN(
        P2_U3187) );
  AND2_X1 U22437 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19503), .ZN(
        P2_U3188) );
  AND2_X1 U22438 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19503), .ZN(
        P2_U3189) );
  AND2_X1 U22439 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19503), .ZN(
        P2_U3190) );
  AND2_X1 U22440 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19503), .ZN(
        P2_U3191) );
  AND2_X1 U22441 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19503), .ZN(
        P2_U3192) );
  AND2_X1 U22442 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19503), .ZN(
        P2_U3193) );
  AND2_X1 U22443 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19503), .ZN(
        P2_U3194) );
  AND2_X1 U22444 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19503), .ZN(
        P2_U3195) );
  AND2_X1 U22445 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19503), .ZN(
        P2_U3196) );
  AND2_X1 U22446 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19503), .ZN(
        P2_U3197) );
  AND2_X1 U22447 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19503), .ZN(
        P2_U3198) );
  AND2_X1 U22448 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19503), .ZN(
        P2_U3199) );
  AND2_X1 U22449 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19503), .ZN(
        P2_U3200) );
  AND2_X1 U22450 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19503), .ZN(P2_U3201) );
  AND2_X1 U22451 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19503), .ZN(P2_U3202) );
  AND2_X1 U22452 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19503), .ZN(P2_U3203) );
  AND2_X1 U22453 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19503), .ZN(P2_U3204) );
  AND2_X1 U22454 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19503), .ZN(P2_U3205) );
  AND2_X1 U22455 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19503), .ZN(P2_U3206) );
  AND2_X1 U22456 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19503), .ZN(P2_U3207) );
  AND2_X1 U22457 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19503), .ZN(P2_U3208) );
  INV_X1 U22458 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19515) );
  NOR2_X1 U22459 ( .A1(n19517), .A2(n19504), .ZN(n19514) );
  OR3_X1 U22460 ( .A1(n19515), .A2(n19505), .A3(n19514), .ZN(n19506) );
  NOR3_X1 U22461 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n20513), .ZN(n19522) );
  AOI21_X1 U22462 ( .B1(n19525), .B2(n19506), .A(n19522), .ZN(n19507) );
  OAI221_X1 U22463 ( .B1(n19508), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .C1(
        n19508), .C2(n20782), .A(n19507), .ZN(P2_U3209) );
  AOI21_X1 U22464 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20782), .A(n19525), 
        .ZN(n19518) );
  NOR3_X1 U22465 ( .A1(n19518), .A2(n19515), .A3(n19505), .ZN(n19509) );
  NOR2_X1 U22466 ( .A1(n19509), .A2(n19514), .ZN(n19512) );
  INV_X1 U22467 ( .A(n19510), .ZN(n19511) );
  OAI211_X1 U22468 ( .C1(n20782), .C2(n19513), .A(n19512), .B(n19511), .ZN(
        P2_U3210) );
  AOI22_X1 U22469 ( .A1(n19516), .A2(n19515), .B1(n19514), .B2(n20513), .ZN(
        n19524) );
  OAI21_X1 U22470 ( .B1(HOLD), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n19523) );
  NOR2_X1 U22471 ( .A1(n19517), .A2(n19525), .ZN(n19519) );
  AOI21_X1 U22472 ( .B1(n19520), .B2(n19519), .A(n19518), .ZN(n19521) );
  OAI22_X1 U22473 ( .A1(n19524), .A2(n19523), .B1(n19522), .B2(n19521), .ZN(
        P2_U3211) );
  NAND2_X1 U22474 ( .A1(n19627), .A2(n19525), .ZN(n19571) );
  CLKBUF_X1 U22475 ( .A(n19571), .Z(n19568) );
  OAI222_X1 U22476 ( .A1(n19568), .A2(n12761), .B1(n19526), .B2(n19627), .C1(
        n12768), .C2(n19569), .ZN(P2_U3212) );
  OAI222_X1 U22477 ( .A1(n19571), .A2(n16054), .B1(n19527), .B2(n19627), .C1(
        n12761), .C2(n19569), .ZN(P2_U3213) );
  OAI222_X1 U22478 ( .A1(n19571), .A2(n11066), .B1(n19528), .B2(n19627), .C1(
        n16054), .C2(n19569), .ZN(P2_U3214) );
  OAI222_X1 U22479 ( .A1(n19571), .A2(n11072), .B1(n19529), .B2(n19627), .C1(
        n11066), .C2(n19569), .ZN(P2_U3215) );
  OAI222_X1 U22480 ( .A1(n19571), .A2(n11057), .B1(n19530), .B2(n19627), .C1(
        n11072), .C2(n19569), .ZN(P2_U3216) );
  OAI222_X1 U22481 ( .A1(n19571), .A2(n19532), .B1(n19531), .B2(n19627), .C1(
        n11057), .C2(n19569), .ZN(P2_U3217) );
  OAI222_X1 U22482 ( .A1(n19568), .A2(n13323), .B1(n19533), .B2(n19627), .C1(
        n19532), .C2(n19569), .ZN(P2_U3218) );
  OAI222_X1 U22483 ( .A1(n19568), .A2(n19535), .B1(n19534), .B2(n19627), .C1(
        n13323), .C2(n19569), .ZN(P2_U3219) );
  OAI222_X1 U22484 ( .A1(n19568), .A2(n10939), .B1(n19536), .B2(n19627), .C1(
        n19535), .C2(n19569), .ZN(P2_U3220) );
  OAI222_X1 U22485 ( .A1(n19568), .A2(n11088), .B1(n19537), .B2(n19627), .C1(
        n10939), .C2(n19569), .ZN(P2_U3221) );
  OAI222_X1 U22486 ( .A1(n19568), .A2(n11092), .B1(n19538), .B2(n19627), .C1(
        n11088), .C2(n19569), .ZN(P2_U3222) );
  OAI222_X1 U22487 ( .A1(n19568), .A2(n11098), .B1(n19539), .B2(n19627), .C1(
        n11092), .C2(n19569), .ZN(P2_U3223) );
  OAI222_X1 U22488 ( .A1(n19571), .A2(n11102), .B1(n19540), .B2(n19627), .C1(
        n11098), .C2(n19569), .ZN(P2_U3224) );
  OAI222_X1 U22489 ( .A1(n19571), .A2(n19542), .B1(n19541), .B2(n19627), .C1(
        n11102), .C2(n19569), .ZN(P2_U3225) );
  OAI222_X1 U22490 ( .A1(n19571), .A2(n11108), .B1(n19543), .B2(n19627), .C1(
        n19542), .C2(n19569), .ZN(P2_U3226) );
  OAI222_X1 U22491 ( .A1(n19571), .A2(n19545), .B1(n19544), .B2(n19627), .C1(
        n11108), .C2(n19569), .ZN(P2_U3227) );
  INV_X1 U22492 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19547) );
  OAI222_X1 U22493 ( .A1(n19571), .A2(n19547), .B1(n19546), .B2(n19627), .C1(
        n19545), .C2(n19569), .ZN(P2_U3228) );
  OAI222_X1 U22494 ( .A1(n19571), .A2(n19549), .B1(n19548), .B2(n19627), .C1(
        n19547), .C2(n19569), .ZN(P2_U3229) );
  OAI222_X1 U22495 ( .A1(n19568), .A2(n19551), .B1(n19550), .B2(n19627), .C1(
        n19549), .C2(n19569), .ZN(P2_U3230) );
  OAI222_X1 U22496 ( .A1(n19568), .A2(n19553), .B1(n19552), .B2(n19627), .C1(
        n19551), .C2(n19569), .ZN(P2_U3231) );
  OAI222_X1 U22497 ( .A1(n19568), .A2(n12613), .B1(n19554), .B2(n19627), .C1(
        n19553), .C2(n19569), .ZN(P2_U3232) );
  OAI222_X1 U22498 ( .A1(n19568), .A2(n19556), .B1(n19555), .B2(n19627), .C1(
        n12613), .C2(n19569), .ZN(P2_U3233) );
  OAI222_X1 U22499 ( .A1(n19568), .A2(n19558), .B1(n19557), .B2(n19627), .C1(
        n19556), .C2(n19569), .ZN(P2_U3234) );
  OAI222_X1 U22500 ( .A1(n19568), .A2(n19560), .B1(n19559), .B2(n19627), .C1(
        n19558), .C2(n19569), .ZN(P2_U3235) );
  OAI222_X1 U22501 ( .A1(n19568), .A2(n15790), .B1(n19561), .B2(n19627), .C1(
        n19560), .C2(n19569), .ZN(P2_U3236) );
  OAI222_X1 U22502 ( .A1(n19568), .A2(n20763), .B1(n19562), .B2(n19627), .C1(
        n15790), .C2(n19569), .ZN(P2_U3237) );
  INV_X1 U22503 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19564) );
  OAI222_X1 U22504 ( .A1(n19569), .A2(n20763), .B1(n19563), .B2(n19627), .C1(
        n19564), .C2(n19568), .ZN(P2_U3238) );
  OAI222_X1 U22505 ( .A1(n19568), .A2(n19566), .B1(n19565), .B2(n19627), .C1(
        n19564), .C2(n19569), .ZN(P2_U3239) );
  OAI222_X1 U22506 ( .A1(n19568), .A2(n11147), .B1(n19567), .B2(n19627), .C1(
        n19566), .C2(n19569), .ZN(P2_U3240) );
  OAI222_X1 U22507 ( .A1(n19571), .A2(n11152), .B1(n19570), .B2(n19627), .C1(
        n11147), .C2(n19569), .ZN(P2_U3241) );
  INV_X1 U22508 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19572) );
  AOI22_X1 U22509 ( .A1(n19627), .A2(n19573), .B1(n19572), .B2(n19624), .ZN(
        P2_U3585) );
  MUX2_X1 U22510 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19627), .Z(P2_U3586) );
  MUX2_X1 U22511 ( .A(P2_BE_N_REG_1__SCAN_IN), .B(P2_BYTEENABLE_REG_1__SCAN_IN), .S(n19627), .Z(P2_U3587) );
  AOI22_X1 U22512 ( .A1(n19627), .A2(n19574), .B1(n20806), .B2(n19624), .ZN(
        P2_U3588) );
  OAI21_X1 U22513 ( .B1(n19578), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19576), 
        .ZN(n19575) );
  INV_X1 U22514 ( .A(n19575), .ZN(P2_U3591) );
  OAI21_X1 U22515 ( .B1(n19578), .B2(n19577), .A(n19576), .ZN(P2_U3592) );
  INV_X1 U22516 ( .A(n19598), .ZN(n19589) );
  NAND2_X1 U22517 ( .A1(n19590), .A2(n11220), .ZN(n19580) );
  NAND2_X1 U22518 ( .A1(n19580), .A2(n19604), .ZN(n19597) );
  OAI22_X1 U22519 ( .A1(n19583), .A2(n19582), .B1(n19581), .B2(n19597), .ZN(
        n19584) );
  AOI221_X1 U22520 ( .B1(n19586), .B2(n19589), .C1(n19585), .C2(n19589), .A(
        n19584), .ZN(n19587) );
  INV_X1 U22521 ( .A(n19611), .ZN(n19612) );
  AOI22_X1 U22522 ( .A1(n19611), .A2(n19588), .B1(n19587), .B2(n19612), .ZN(
        P2_U3602) );
  NAND3_X1 U22523 ( .A1(n19592), .A2(n19590), .A3(n19589), .ZN(n19591) );
  OAI21_X1 U22524 ( .B1(n19592), .B2(n19597), .A(n19591), .ZN(n19593) );
  AOI21_X1 U22525 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19594), .A(n19593), 
        .ZN(n19595) );
  AOI22_X1 U22526 ( .A1(n19611), .A2(n19596), .B1(n19595), .B2(n19612), .ZN(
        P2_U3603) );
  AOI21_X1 U22527 ( .B1(n19599), .B2(n19598), .A(n19597), .ZN(n19600) );
  AOI21_X1 U22528 ( .B1(n19601), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19600), 
        .ZN(n19602) );
  AOI22_X1 U22529 ( .A1(n19611), .A2(n19603), .B1(n19602), .B2(n19612), .ZN(
        P2_U3604) );
  INV_X1 U22530 ( .A(n19604), .ZN(n19607) );
  OAI22_X1 U22531 ( .A1(n19608), .A2(n19607), .B1(n19606), .B2(n19605), .ZN(
        n19609) );
  AOI21_X1 U22532 ( .B1(n19613), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19609), 
        .ZN(n19610) );
  OAI22_X1 U22533 ( .A1(n19613), .A2(n19612), .B1(n19611), .B2(n19610), .ZN(
        P2_U3605) );
  AOI22_X1 U22534 ( .A1(n19627), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19614), 
        .B2(n19624), .ZN(P2_U3608) );
  INV_X1 U22535 ( .A(n19615), .ZN(n19619) );
  AOI22_X1 U22536 ( .A1(n19619), .A2(n19618), .B1(n19617), .B2(n19616), .ZN(
        n19620) );
  NAND2_X1 U22537 ( .A1(n19621), .A2(n19620), .ZN(n19623) );
  MUX2_X1 U22538 ( .A(P2_MORE_REG_SCAN_IN), .B(n19623), .S(n19622), .Z(
        P2_U3609) );
  INV_X1 U22539 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n19625) );
  AOI22_X1 U22540 ( .A1(n19627), .A2(n19626), .B1(n19625), .B2(n19624), .ZN(
        P2_U3611) );
  AND2_X1 U22541 ( .A1(n20506), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n19629) );
  INV_X1 U22542 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19628) );
  OR2_X1 U22543 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20510), .ZN(n20617) );
  INV_X2 U22544 ( .A(n20617), .ZN(n20630) );
  AOI21_X1 U22545 ( .B1(n19629), .B2(n19628), .A(n20630), .ZN(P1_U2802) );
  NAND2_X1 U22546 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20595), .ZN(n19634) );
  INV_X1 U22547 ( .A(n19630), .ZN(n19632) );
  OAI21_X1 U22548 ( .B1(n19632), .B2(n19631), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19633) );
  OAI21_X1 U22549 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n19634), .A(n19633), 
        .ZN(P1_U2803) );
  NOR2_X1 U22550 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19636) );
  OAI21_X1 U22551 ( .B1(n19636), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20617), .ZN(
        n19635) );
  OAI21_X1 U22552 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20617), .A(n19635), 
        .ZN(P1_U2804) );
  AOI21_X1 U22553 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20506), .A(n20630), 
        .ZN(n20587) );
  OAI21_X1 U22554 ( .B1(BS16), .B2(n19636), .A(n20587), .ZN(n20585) );
  OAI21_X1 U22555 ( .B1(n20587), .B2(n20334), .A(n20585), .ZN(P1_U2805) );
  OAI21_X1 U22556 ( .B1(n19639), .B2(n19638), .A(n19637), .ZN(P1_U2806) );
  NOR4_X1 U22557 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19643) );
  NOR4_X1 U22558 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19642) );
  NOR4_X1 U22559 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19641) );
  NOR4_X1 U22560 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19640) );
  NAND4_X1 U22561 ( .A1(n19643), .A2(n19642), .A3(n19641), .A4(n19640), .ZN(
        n19649) );
  NOR4_X1 U22562 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19647) );
  AOI211_X1 U22563 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_20__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19646) );
  NOR4_X1 U22564 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19645) );
  NOR4_X1 U22565 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19644) );
  NAND4_X1 U22566 ( .A1(n19647), .A2(n19646), .A3(n19645), .A4(n19644), .ZN(
        n19648) );
  NOR2_X1 U22567 ( .A1(n19649), .A2(n19648), .ZN(n20616) );
  INV_X1 U22568 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20580) );
  NOR3_X1 U22569 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19651) );
  OAI21_X1 U22570 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19651), .A(n20616), .ZN(
        n19650) );
  OAI21_X1 U22571 ( .B1(n20616), .B2(n20580), .A(n19650), .ZN(P1_U2807) );
  INV_X1 U22572 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20586) );
  AOI21_X1 U22573 ( .B1(n20609), .B2(n20586), .A(n19651), .ZN(n19652) );
  INV_X1 U22574 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20577) );
  INV_X1 U22575 ( .A(n20616), .ZN(n20611) );
  AOI22_X1 U22576 ( .A1(n20616), .A2(n19652), .B1(n20577), .B2(n20611), .ZN(
        P1_U2808) );
  AOI22_X1 U22577 ( .A1(n19700), .A2(n19733), .B1(n19653), .B2(n13588), .ZN(
        n19660) );
  OAI22_X1 U22578 ( .A1(n19654), .A2(n13588), .B1(n19736), .B2(n19715), .ZN(
        n19655) );
  AOI211_X1 U22579 ( .C1(n19721), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n19662), .B(n19655), .ZN(n19659) );
  INV_X1 U22580 ( .A(n19656), .ZN(n19734) );
  AOI22_X1 U22581 ( .A1(n19734), .A2(n19663), .B1(n19703), .B2(n19657), .ZN(
        n19658) );
  NAND3_X1 U22582 ( .A1(n19660), .A2(n19659), .A3(n19658), .ZN(P1_U2831) );
  INV_X1 U22583 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20527) );
  INV_X1 U22584 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20525) );
  NOR3_X1 U22585 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20525), .A3(n19674), .ZN(
        n19661) );
  AOI211_X1 U22586 ( .C1(n19721), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n19662), .B(n19661), .ZN(n19671) );
  NAND2_X1 U22587 ( .A1(n19664), .A2(n19663), .ZN(n19670) );
  INV_X1 U22588 ( .A(n19665), .ZN(n19666) );
  AOI22_X1 U22589 ( .A1(n19695), .A2(P1_EBX_REG_6__SCAN_IN), .B1(n19666), .B2(
        n19703), .ZN(n19669) );
  NAND2_X1 U22590 ( .A1(n19700), .A2(n19667), .ZN(n19668) );
  AND4_X1 U22591 ( .A1(n19671), .A2(n19670), .A3(n19669), .A4(n19668), .ZN(
        n19672) );
  OAI21_X1 U22592 ( .B1(n19673), .B2(n20527), .A(n19672), .ZN(P1_U2834) );
  INV_X1 U22593 ( .A(n19674), .ZN(n19675) );
  AOI22_X1 U22594 ( .A1(n19700), .A2(n19737), .B1(n19675), .B2(n20525), .ZN(
        n19681) );
  NAND2_X1 U22595 ( .A1(n19690), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n19678) );
  NAND2_X1 U22596 ( .A1(n19695), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n19677) );
  NAND2_X1 U22597 ( .A1(n19721), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n19676) );
  NAND4_X1 U22598 ( .A1(n19678), .A2(n19683), .A3(n19677), .A4(n19676), .ZN(
        n19679) );
  AOI21_X1 U22599 ( .B1(n19740), .B2(n19727), .A(n19679), .ZN(n19680) );
  OAI211_X1 U22600 ( .C1(n19682), .C2(n19731), .A(n19681), .B(n19680), .ZN(
        P1_U2835) );
  OAI21_X1 U22601 ( .B1(n19723), .B2(n19684), .A(n19683), .ZN(n19687) );
  OAI22_X1 U22602 ( .A1(n19718), .A2(n19685), .B1(n13314), .B2(n19715), .ZN(
        n19686) );
  AOI211_X1 U22603 ( .C1(n19721), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n19687), .B(n19686), .ZN(n19693) );
  OAI21_X1 U22604 ( .B1(n19709), .B2(n19688), .A(n20522), .ZN(n19689) );
  AOI22_X1 U22605 ( .A1(n19691), .A2(n19727), .B1(n19690), .B2(n19689), .ZN(
        n19692) );
  OAI211_X1 U22606 ( .C1(n19694), .C2(n19731), .A(n19693), .B(n19692), .ZN(
        P1_U2836) );
  AOI222_X1 U22607 ( .A1(n13201), .A2(n19696), .B1(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n19721), .C1(n19695), .C2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n19713) );
  INV_X1 U22608 ( .A(n19697), .ZN(n19699) );
  NOR3_X1 U22609 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n20609), .A3(n19709), .ZN(
        n19698) );
  AOI22_X1 U22610 ( .A1(n19700), .A2(n19699), .B1(P1_REIP_REG_2__SCAN_IN), 
        .B2(n19698), .ZN(n19712) );
  INV_X1 U22611 ( .A(n19701), .ZN(n19705) );
  INV_X1 U22612 ( .A(n19702), .ZN(n19704) );
  AOI22_X1 U22613 ( .A1(n19705), .A2(n19727), .B1(n19704), .B2(n19703), .ZN(
        n19711) );
  NAND2_X1 U22614 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n19706), .ZN(n19707) );
  NOR2_X1 U22615 ( .A1(n19709), .A2(n19707), .ZN(n19725) );
  OAI21_X1 U22616 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19709), .A(n19708), .ZN(
        n19720) );
  OAI21_X1 U22617 ( .B1(n19725), .B2(n19720), .A(P1_REIP_REG_3__SCAN_IN), .ZN(
        n19710) );
  NAND4_X1 U22618 ( .A1(n19713), .A2(n19712), .A3(n19711), .A4(n19710), .ZN(
        P1_U2837) );
  INV_X1 U22619 ( .A(n19714), .ZN(n19732) );
  OAI22_X1 U22620 ( .A1(n19718), .A2(n19717), .B1(n19716), .B2(n19715), .ZN(
        n19719) );
  AOI21_X1 U22621 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(n19720), .A(n19719), .ZN(
        n19730) );
  NAND2_X1 U22622 ( .A1(n19721), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19722) );
  OAI21_X1 U22623 ( .B1(n13187), .B2(n19723), .A(n19722), .ZN(n19724) );
  OR2_X1 U22624 ( .A1(n19725), .A2(n19724), .ZN(n19726) );
  AOI21_X1 U22625 ( .B1(n19728), .B2(n19727), .A(n19726), .ZN(n19729) );
  OAI211_X1 U22626 ( .C1(n19732), .C2(n19731), .A(n19730), .B(n19729), .ZN(
        P1_U2838) );
  AOI22_X1 U22627 ( .A1(n19734), .A2(n19739), .B1(n19738), .B2(n19733), .ZN(
        n19735) );
  OAI21_X1 U22628 ( .B1(n19742), .B2(n19736), .A(n19735), .ZN(P1_U2863) );
  AOI22_X1 U22629 ( .A1(n19740), .A2(n19739), .B1(n19738), .B2(n19737), .ZN(
        n19741) );
  OAI21_X1 U22630 ( .B1(n19742), .B2(n20661), .A(n19741), .ZN(P1_U2867) );
  INV_X1 U22631 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n20812) );
  INV_X1 U22632 ( .A(n19743), .ZN(n19744) );
  AOI22_X1 U22633 ( .A1(n19744), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n19777), .ZN(n19745) );
  OAI21_X1 U22634 ( .B1(n20812), .B2(n19747), .A(n19745), .ZN(P1_U2906) );
  OAI222_X1 U22635 ( .A1(n19760), .A2(n19749), .B1(n19779), .B2(n19748), .C1(
        n19747), .C2(n19746), .ZN(P1_U2921) );
  INV_X1 U22636 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n19751) );
  AOI22_X1 U22637 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n19777), .B1(n19776), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19750) );
  OAI21_X1 U22638 ( .B1(n19751), .B2(n19779), .A(n19750), .ZN(P1_U2922) );
  INV_X1 U22639 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n19753) );
  AOI22_X1 U22640 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n19777), .B1(n19776), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19752) );
  OAI21_X1 U22641 ( .B1(n19753), .B2(n19779), .A(n19752), .ZN(P1_U2923) );
  AOI22_X1 U22642 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n19771), .B1(n19776), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19754) );
  OAI21_X1 U22643 ( .B1(n14211), .B2(n19779), .A(n19754), .ZN(P1_U2924) );
  AOI22_X1 U22644 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n19771), .B1(n19776), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19755) );
  OAI21_X1 U22645 ( .B1(n13631), .B2(n19779), .A(n19755), .ZN(P1_U2925) );
  INV_X1 U22646 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n19757) );
  AOI22_X1 U22647 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n19771), .B1(n19776), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19756) );
  OAI21_X1 U22648 ( .B1(n19757), .B2(n19779), .A(n19756), .ZN(P1_U2926) );
  INV_X1 U22649 ( .A(P1_LWORD_REG_9__SCAN_IN), .ZN(n20632) );
  INV_X1 U22650 ( .A(n19779), .ZN(n19758) );
  AOI22_X1 U22651 ( .A1(P1_EAX_REG_9__SCAN_IN), .A2(n19758), .B1(n19776), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n19759) );
  OAI21_X1 U22652 ( .B1(n20632), .B2(n19760), .A(n19759), .ZN(P1_U2927) );
  INV_X1 U22653 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n19762) );
  AOI22_X1 U22654 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n19771), .B1(n19776), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19761) );
  OAI21_X1 U22655 ( .B1(n19762), .B2(n19779), .A(n19761), .ZN(P1_U2928) );
  AOI22_X1 U22656 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n19771), .B1(n19776), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19763) );
  OAI21_X1 U22657 ( .B1(n19764), .B2(n19779), .A(n19763), .ZN(P1_U2929) );
  AOI22_X1 U22658 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n19771), .B1(n19776), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19765) );
  OAI21_X1 U22659 ( .B1(n11961), .B2(n19779), .A(n19765), .ZN(P1_U2930) );
  AOI22_X1 U22660 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n19771), .B1(n19776), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19766) );
  OAI21_X1 U22661 ( .B1(n11944), .B2(n19779), .A(n19766), .ZN(P1_U2931) );
  AOI22_X1 U22662 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n19771), .B1(n19776), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19767) );
  OAI21_X1 U22663 ( .B1(n19768), .B2(n19779), .A(n19767), .ZN(P1_U2932) );
  AOI22_X1 U22664 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n19771), .B1(n19776), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19769) );
  OAI21_X1 U22665 ( .B1(n19770), .B2(n19779), .A(n19769), .ZN(P1_U2933) );
  AOI22_X1 U22666 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n19771), .B1(n19776), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19772) );
  OAI21_X1 U22667 ( .B1(n19773), .B2(n19779), .A(n19772), .ZN(P1_U2934) );
  AOI22_X1 U22668 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n19777), .B1(n19776), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19774) );
  OAI21_X1 U22669 ( .B1(n19775), .B2(n19779), .A(n19774), .ZN(P1_U2935) );
  AOI22_X1 U22670 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n19777), .B1(n19776), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19778) );
  OAI21_X1 U22671 ( .B1(n19780), .B2(n19779), .A(n19778), .ZN(P1_U2936) );
  AOI22_X1 U22672 ( .A1(n19809), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n19804), .ZN(n19782) );
  NAND2_X1 U22673 ( .A1(n19792), .A2(n19781), .ZN(n19794) );
  NAND2_X1 U22674 ( .A1(n19782), .A2(n19794), .ZN(P1_U2945) );
  AOI22_X1 U22675 ( .A1(n19809), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n19804), .ZN(n19784) );
  NAND2_X1 U22676 ( .A1(n19792), .A2(n19783), .ZN(n19800) );
  NAND2_X1 U22677 ( .A1(n19784), .A2(n19800), .ZN(P1_U2947) );
  AOI22_X1 U22678 ( .A1(n19809), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n19804), .ZN(n19786) );
  NAND2_X1 U22679 ( .A1(n19792), .A2(n19785), .ZN(n19802) );
  NAND2_X1 U22680 ( .A1(n19786), .A2(n19802), .ZN(P1_U2948) );
  AOI22_X1 U22681 ( .A1(n19809), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n19804), .ZN(n19788) );
  NAND2_X1 U22682 ( .A1(n19792), .A2(n19787), .ZN(n19805) );
  NAND2_X1 U22683 ( .A1(n19788), .A2(n19805), .ZN(P1_U2949) );
  AOI22_X1 U22684 ( .A1(n19809), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n19804), .ZN(n19790) );
  NAND2_X1 U22685 ( .A1(n19792), .A2(n19789), .ZN(n19807) );
  NAND2_X1 U22686 ( .A1(n19790), .A2(n19807), .ZN(P1_U2950) );
  AOI22_X1 U22687 ( .A1(n19809), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n19804), .ZN(n19793) );
  NAND2_X1 U22688 ( .A1(n19792), .A2(n19791), .ZN(n19810) );
  NAND2_X1 U22689 ( .A1(n19793), .A2(n19810), .ZN(P1_U2951) );
  AOI22_X1 U22690 ( .A1(n19809), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n19804), .ZN(n19795) );
  NAND2_X1 U22691 ( .A1(n19795), .A2(n19794), .ZN(P1_U2960) );
  NAND2_X1 U22692 ( .A1(n19809), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n19796) );
  AND2_X1 U22693 ( .A1(n19797), .A2(n19796), .ZN(n19798) );
  OAI21_X1 U22694 ( .B1(n19799), .B2(n20632), .A(n19798), .ZN(P1_U2961) );
  AOI22_X1 U22695 ( .A1(n19809), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n19804), .ZN(n19801) );
  NAND2_X1 U22696 ( .A1(n19801), .A2(n19800), .ZN(P1_U2962) );
  AOI22_X1 U22697 ( .A1(n19809), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n19804), .ZN(n19803) );
  NAND2_X1 U22698 ( .A1(n19803), .A2(n19802), .ZN(P1_U2963) );
  AOI22_X1 U22699 ( .A1(n19809), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n19804), .ZN(n19806) );
  NAND2_X1 U22700 ( .A1(n19806), .A2(n19805), .ZN(P1_U2964) );
  AOI22_X1 U22701 ( .A1(n19809), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n19804), .ZN(n19808) );
  NAND2_X1 U22702 ( .A1(n19808), .A2(n19807), .ZN(P1_U2965) );
  AOI22_X1 U22703 ( .A1(n19809), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n19804), .ZN(n19811) );
  NAND2_X1 U22704 ( .A1(n19811), .A2(n19810), .ZN(P1_U2966) );
  OR2_X1 U22705 ( .A1(n19813), .A2(n19812), .ZN(n19818) );
  INV_X1 U22706 ( .A(n19814), .ZN(n19816) );
  AOI21_X1 U22707 ( .B1(n19816), .B2(n19830), .A(n19815), .ZN(n19823) );
  AOI22_X1 U22708 ( .A1(n19818), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19817), .B2(n19823), .ZN(n19820) );
  NAND2_X1 U22709 ( .A1(n19819), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n19835) );
  OAI211_X1 U22710 ( .C1(n19821), .C2(n19841), .A(n19820), .B(n19835), .ZN(
        P1_U2999) );
  INV_X1 U22711 ( .A(n19822), .ZN(n19825) );
  AOI22_X1 U22712 ( .A1(n19826), .A2(n19825), .B1(n19824), .B2(n19823), .ZN(
        n19836) );
  INV_X1 U22713 ( .A(n19827), .ZN(n19832) );
  NAND3_X1 U22714 ( .A1(n19830), .A2(n19829), .A3(n19828), .ZN(n19831) );
  OAI21_X1 U22715 ( .B1(n19833), .B2(n19832), .A(n19831), .ZN(n19834) );
  NAND3_X1 U22716 ( .A1(n19836), .A2(n19835), .A3(n19834), .ZN(P1_U3031) );
  NOR2_X1 U22717 ( .A1(n19838), .A2(n19837), .ZN(P1_U3032) );
  AOI22_X1 U22718 ( .A1(DATAI_16_), .A2(n9605), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n9606), .ZN(n20341) );
  NAND2_X1 U22719 ( .A1(n19842), .A2(n13225), .ZN(n19970) );
  NAND2_X1 U22720 ( .A1(n9635), .A2(n19843), .ZN(n20252) );
  NAND2_X1 U22721 ( .A1(n19887), .A2(n9618), .ZN(n20379) );
  NOR2_X1 U22722 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19964) );
  INV_X1 U22723 ( .A(n19964), .ZN(n19845) );
  NOR2_X1 U22724 ( .A1(n19845), .A2(n20286), .ZN(n19850) );
  INV_X1 U22725 ( .A(n19850), .ZN(n19888) );
  OAI22_X1 U22726 ( .A1(n20449), .A2(n20453), .B1(n20379), .B2(n19888), .ZN(
        n19846) );
  INV_X1 U22727 ( .A(n19846), .ZN(n19857) );
  NAND2_X1 U22728 ( .A1(n19853), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20298) );
  AND2_X1 U22729 ( .A1(n20010), .A2(n20298), .ZN(n20220) );
  NAND3_X1 U22730 ( .A1(n19918), .A2(n20288), .A3(n20449), .ZN(n19847) );
  NAND2_X1 U22731 ( .A1(n19847), .A2(n20289), .ZN(n19852) );
  INV_X1 U22732 ( .A(n13187), .ZN(n19848) );
  OR2_X1 U22733 ( .A1(n13201), .A2(n19848), .ZN(n19928) );
  OR2_X1 U22734 ( .A1(n19928), .A2(n9622), .ZN(n19854) );
  INV_X1 U22735 ( .A(n20218), .ZN(n19933) );
  OR2_X1 U22736 ( .A1(n19933), .A2(n20151), .ZN(n20004) );
  AOI22_X1 U22737 ( .A1(n19852), .A2(n19854), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20004), .ZN(n19849) );
  OAI211_X1 U22738 ( .C1(n19850), .C2(n20294), .A(n20220), .B(n19849), .ZN(
        n19892) );
  NOR2_X2 U22739 ( .A1(n19851), .A2(n19899), .ZN(n20439) );
  INV_X1 U22740 ( .A(n19852), .ZN(n19855) );
  OR2_X1 U22741 ( .A1(n19853), .A2(n20437), .ZN(n20222) );
  OAI22_X1 U22742 ( .A1(n19855), .A2(n19854), .B1(n20222), .B2(n20004), .ZN(
        n19891) );
  AOI22_X1 U22743 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19892), .B1(
        n20439), .B2(n19891), .ZN(n19856) );
  OAI211_X1 U22744 ( .C1(n20341), .C2(n19918), .A(n19857), .B(n19856), .ZN(
        P1_U3033) );
  AOI22_X1 U22745 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n9606), .B1(DATAI_25_), 
        .B2(n9605), .ZN(n20459) );
  NAND2_X1 U22746 ( .A1(n19887), .A2(n19858), .ZN(n20393) );
  OAI22_X1 U22747 ( .A1(n20449), .A2(n20459), .B1(n20393), .B2(n19888), .ZN(
        n19859) );
  INV_X1 U22748 ( .A(n19859), .ZN(n19862) );
  NOR2_X2 U22749 ( .A1(n19860), .A2(n19899), .ZN(n20454) );
  AOI22_X1 U22750 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19892), .B1(
        n20454), .B2(n19891), .ZN(n19861) );
  OAI211_X1 U22751 ( .C1(n20345), .C2(n19918), .A(n19862), .B(n19861), .ZN(
        P1_U3034) );
  AOI22_X1 U22752 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n9606), .B1(DATAI_18_), 
        .B2(n9605), .ZN(n20349) );
  NAND2_X1 U22753 ( .A1(n19887), .A2(n19863), .ZN(n20398) );
  OAI22_X1 U22754 ( .A1(n20449), .A2(n20465), .B1(n20398), .B2(n19888), .ZN(
        n19864) );
  INV_X1 U22755 ( .A(n19864), .ZN(n19867) );
  NOR2_X2 U22756 ( .A1(n19865), .A2(n19899), .ZN(n20460) );
  AOI22_X1 U22757 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19892), .B1(
        n20460), .B2(n19891), .ZN(n19866) );
  OAI211_X1 U22758 ( .C1(n20349), .C2(n19918), .A(n19867), .B(n19866), .ZN(
        P1_U3035) );
  AOI22_X1 U22759 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n9606), .B1(DATAI_19_), 
        .B2(n9605), .ZN(n20353) );
  NAND2_X1 U22760 ( .A1(n19887), .A2(n19868), .ZN(n20403) );
  OAI22_X1 U22761 ( .A1(n20449), .A2(n20470), .B1(n20403), .B2(n19888), .ZN(
        n19869) );
  INV_X1 U22762 ( .A(n19869), .ZN(n19872) );
  NOR2_X2 U22763 ( .A1(n19870), .A2(n19899), .ZN(n20466) );
  AOI22_X1 U22764 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19892), .B1(
        n20466), .B2(n19891), .ZN(n19871) );
  OAI211_X1 U22765 ( .C1(n9756), .C2(n19918), .A(n19872), .B(n19871), .ZN(
        P1_U3036) );
  AOI22_X1 U22766 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n9606), .B1(DATAI_28_), 
        .B2(n9605), .ZN(n20476) );
  NAND2_X1 U22767 ( .A1(n19887), .A2(n11737), .ZN(n20408) );
  OAI22_X1 U22768 ( .A1(n20449), .A2(n20476), .B1(n20408), .B2(n19888), .ZN(
        n19873) );
  INV_X1 U22769 ( .A(n19873), .ZN(n19876) );
  NOR2_X2 U22770 ( .A1(n19874), .A2(n19899), .ZN(n20471) );
  AOI22_X1 U22771 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19892), .B1(
        n20471), .B2(n19891), .ZN(n19875) );
  OAI211_X1 U22772 ( .C1(n20357), .C2(n19918), .A(n19876), .B(n19875), .ZN(
        P1_U3037) );
  AOI22_X1 U22773 ( .A1(DATAI_21_), .A2(n9605), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n9606), .ZN(n20361) );
  NAND2_X1 U22774 ( .A1(n19887), .A2(n12415), .ZN(n20413) );
  OAI22_X1 U22775 ( .A1(n20449), .A2(n20482), .B1(n20413), .B2(n19888), .ZN(
        n19877) );
  INV_X1 U22776 ( .A(n19877), .ZN(n19880) );
  NOR2_X2 U22777 ( .A1(n19878), .A2(n19899), .ZN(n20477) );
  AOI22_X1 U22778 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19892), .B1(
        n20477), .B2(n19891), .ZN(n19879) );
  OAI211_X1 U22779 ( .C1(n20361), .C2(n19918), .A(n19880), .B(n19879), .ZN(
        P1_U3038) );
  AOI22_X1 U22780 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n9606), .B1(DATAI_30_), 
        .B2(n9605), .ZN(n20488) );
  NAND2_X1 U22781 ( .A1(n19887), .A2(n12465), .ZN(n20418) );
  OAI22_X1 U22782 ( .A1(n20449), .A2(n9758), .B1(n20418), .B2(n19888), .ZN(
        n19881) );
  INV_X1 U22783 ( .A(n19881), .ZN(n19884) );
  NOR2_X2 U22784 ( .A1(n19882), .A2(n19899), .ZN(n20483) );
  AOI22_X1 U22785 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19892), .B1(
        n20483), .B2(n19891), .ZN(n19883) );
  OAI211_X1 U22786 ( .C1(n20364), .C2(n19918), .A(n19884), .B(n19883), .ZN(
        P1_U3039) );
  AOI22_X1 U22787 ( .A1(DATAI_23_), .A2(n9605), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n9606), .ZN(n20372) );
  NAND2_X1 U22788 ( .A1(n19887), .A2(n11844), .ZN(n20425) );
  OAI22_X1 U22789 ( .A1(n20449), .A2(n20499), .B1(n20425), .B2(n19888), .ZN(
        n19889) );
  INV_X1 U22790 ( .A(n19889), .ZN(n19894) );
  NOR2_X2 U22791 ( .A1(n19890), .A2(n19899), .ZN(n20490) );
  AOI22_X1 U22792 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19892), .B1(
        n20490), .B2(n19891), .ZN(n19893) );
  OAI211_X1 U22793 ( .C1(n20372), .C2(n19918), .A(n19894), .B(n19893), .ZN(
        P1_U3040) );
  INV_X1 U22794 ( .A(n20379), .ZN(n20440) );
  NAND2_X1 U22795 ( .A1(n19964), .A2(n20436), .ZN(n19896) );
  NOR2_X1 U22796 ( .A1(n20639), .A2(n19896), .ZN(n19920) );
  INV_X1 U22797 ( .A(n19928), .ZN(n19968) );
  INV_X1 U22798 ( .A(n19895), .ZN(n20330) );
  AOI21_X1 U22799 ( .B1(n19968), .B2(n20330), .A(n19920), .ZN(n19900) );
  OR2_X1 U22800 ( .A1(n19900), .A2(n20442), .ZN(n19898) );
  INV_X1 U22801 ( .A(n19896), .ZN(n19902) );
  NAND2_X1 U22802 ( .A1(n19902), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n19897) );
  NAND2_X1 U22803 ( .A1(n19898), .A2(n19897), .ZN(n19919) );
  AOI22_X1 U22804 ( .A1(n20440), .A2(n19920), .B1(n20439), .B2(n19919), .ZN(
        n19904) );
  OAI211_X1 U22805 ( .C1(n19970), .C2(n20334), .A(n20333), .B(n19900), .ZN(
        n19901) );
  OAI211_X1 U22806 ( .C1(n20288), .C2(n19902), .A(n20447), .B(n19901), .ZN(
        n19922) );
  INV_X1 U22807 ( .A(n19962), .ZN(n19915) );
  INV_X1 U22808 ( .A(n20341), .ZN(n20450) );
  AOI22_X1 U22809 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19922), .B1(
        n19915), .B2(n20450), .ZN(n19903) );
  OAI211_X1 U22810 ( .C1(n20453), .C2(n19918), .A(n19904), .B(n19903), .ZN(
        P1_U3041) );
  INV_X1 U22811 ( .A(n20393), .ZN(n20455) );
  AOI22_X1 U22812 ( .A1(n20455), .A2(n19920), .B1(n20454), .B2(n19919), .ZN(
        n19906) );
  INV_X1 U22813 ( .A(n20345), .ZN(n20456) );
  AOI22_X1 U22814 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19922), .B1(
        n19915), .B2(n20456), .ZN(n19905) );
  OAI211_X1 U22815 ( .C1(n20459), .C2(n19918), .A(n19906), .B(n19905), .ZN(
        P1_U3042) );
  INV_X1 U22816 ( .A(n20398), .ZN(n20461) );
  AOI22_X1 U22817 ( .A1(n20461), .A2(n19920), .B1(n20460), .B2(n19919), .ZN(
        n19908) );
  INV_X1 U22818 ( .A(n20349), .ZN(n20462) );
  AOI22_X1 U22819 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19922), .B1(
        n19915), .B2(n20462), .ZN(n19907) );
  OAI211_X1 U22820 ( .C1(n20465), .C2(n19918), .A(n19908), .B(n19907), .ZN(
        P1_U3043) );
  INV_X1 U22821 ( .A(n20403), .ZN(n20467) );
  AOI22_X1 U22822 ( .A1(n20467), .A2(n19920), .B1(n20466), .B2(n19919), .ZN(
        n19910) );
  AOI22_X1 U22823 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19922), .B1(
        n19915), .B2(n9755), .ZN(n19909) );
  OAI211_X1 U22824 ( .C1(n20470), .C2(n19918), .A(n19910), .B(n19909), .ZN(
        P1_U3044) );
  INV_X1 U22825 ( .A(n20408), .ZN(n20472) );
  AOI22_X1 U22826 ( .A1(n20472), .A2(n19920), .B1(n20471), .B2(n19919), .ZN(
        n19912) );
  INV_X1 U22827 ( .A(n19918), .ZN(n19921) );
  INV_X1 U22828 ( .A(n20476), .ZN(n20354) );
  AOI22_X1 U22829 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19922), .B1(
        n19921), .B2(n20354), .ZN(n19911) );
  OAI211_X1 U22830 ( .C1(n20357), .C2(n19962), .A(n19912), .B(n19911), .ZN(
        P1_U3045) );
  INV_X1 U22831 ( .A(n20413), .ZN(n20478) );
  AOI22_X1 U22832 ( .A1(n20478), .A2(n19920), .B1(n20477), .B2(n19919), .ZN(
        n19914) );
  INV_X1 U22833 ( .A(n20482), .ZN(n20358) );
  AOI22_X1 U22834 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19922), .B1(
        n19921), .B2(n20358), .ZN(n19913) );
  OAI211_X1 U22835 ( .C1(n20361), .C2(n19962), .A(n19914), .B(n19913), .ZN(
        P1_U3046) );
  INV_X1 U22836 ( .A(n20418), .ZN(n20484) );
  AOI22_X1 U22837 ( .A1(n20484), .A2(n19920), .B1(n20483), .B2(n19919), .ZN(
        n19917) );
  INV_X1 U22838 ( .A(n20364), .ZN(n20485) );
  AOI22_X1 U22839 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19922), .B1(
        n19915), .B2(n20485), .ZN(n19916) );
  OAI211_X1 U22840 ( .C1(n9758), .C2(n19918), .A(n19917), .B(n19916), .ZN(
        P1_U3047) );
  INV_X1 U22841 ( .A(n20425), .ZN(n20492) );
  AOI22_X1 U22842 ( .A1(n20492), .A2(n19920), .B1(n20490), .B2(n19919), .ZN(
        n19924) );
  INV_X1 U22843 ( .A(n20499), .ZN(n20367) );
  AOI22_X1 U22844 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19922), .B1(
        n19921), .B2(n20367), .ZN(n19923) );
  OAI211_X1 U22845 ( .C1(n20372), .C2(n19962), .A(n19924), .B(n19923), .ZN(
        P1_U3048) );
  NAND2_X1 U22846 ( .A1(n9635), .A2(n19925), .ZN(n20381) );
  NAND2_X1 U22847 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19964), .ZN(
        n19973) );
  NOR2_X1 U22848 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19973), .ZN(
        n19929) );
  INV_X1 U22849 ( .A(n19929), .ZN(n19956) );
  OAI22_X1 U22850 ( .A1(n19997), .A2(n20341), .B1(n20379), .B2(n19956), .ZN(
        n19926) );
  INV_X1 U22851 ( .A(n19926), .ZN(n19937) );
  NAND2_X1 U22852 ( .A1(n19997), .A2(n19962), .ZN(n19927) );
  AOI21_X1 U22853 ( .B1(n19927), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20442), 
        .ZN(n19932) );
  OR2_X1 U22854 ( .A1(n19928), .A2(n20292), .ZN(n19934) );
  NOR2_X1 U22855 ( .A1(n19929), .A2(n20294), .ZN(n19930) );
  AOI21_X1 U22856 ( .B1(n19932), .B2(n19934), .A(n19930), .ZN(n19931) );
  OAI21_X1 U22857 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20218), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20078) );
  NAND3_X1 U22858 ( .A1(n20220), .A2(n19931), .A3(n20078), .ZN(n19959) );
  INV_X1 U22859 ( .A(n19932), .ZN(n19935) );
  NAND2_X1 U22860 ( .A1(n19933), .A2(n20217), .ZN(n20081) );
  OAI22_X1 U22861 ( .A1(n19935), .A2(n19934), .B1(n20222), .B2(n20081), .ZN(
        n19958) );
  AOI22_X1 U22862 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19959), .B1(
        n20439), .B2(n19958), .ZN(n19936) );
  OAI211_X1 U22863 ( .C1(n20453), .C2(n19962), .A(n19937), .B(n19936), .ZN(
        P1_U3049) );
  OAI22_X1 U22864 ( .A1(n19962), .A2(n20459), .B1(n19956), .B2(n20393), .ZN(
        n19938) );
  INV_X1 U22865 ( .A(n19938), .ZN(n19940) );
  AOI22_X1 U22866 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19959), .B1(
        n20454), .B2(n19958), .ZN(n19939) );
  OAI211_X1 U22867 ( .C1(n20345), .C2(n19997), .A(n19940), .B(n19939), .ZN(
        P1_U3050) );
  OAI22_X1 U22868 ( .A1(n19997), .A2(n20349), .B1(n19956), .B2(n20398), .ZN(
        n19941) );
  INV_X1 U22869 ( .A(n19941), .ZN(n19943) );
  AOI22_X1 U22870 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19959), .B1(
        n20460), .B2(n19958), .ZN(n19942) );
  OAI211_X1 U22871 ( .C1(n20465), .C2(n19962), .A(n19943), .B(n19942), .ZN(
        P1_U3051) );
  OAI22_X1 U22872 ( .A1(n19962), .A2(n20470), .B1(n19956), .B2(n20403), .ZN(
        n19944) );
  INV_X1 U22873 ( .A(n19944), .ZN(n19946) );
  AOI22_X1 U22874 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19959), .B1(
        n20466), .B2(n19958), .ZN(n19945) );
  OAI211_X1 U22875 ( .C1(n9756), .C2(n19997), .A(n19946), .B(n19945), .ZN(
        P1_U3052) );
  OAI22_X1 U22876 ( .A1(n19962), .A2(n20476), .B1(n19956), .B2(n20408), .ZN(
        n19947) );
  INV_X1 U22877 ( .A(n19947), .ZN(n19949) );
  AOI22_X1 U22878 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19959), .B1(
        n20471), .B2(n19958), .ZN(n19948) );
  OAI211_X1 U22879 ( .C1(n20357), .C2(n19997), .A(n19949), .B(n19948), .ZN(
        P1_U3053) );
  OAI22_X1 U22880 ( .A1(n19997), .A2(n20361), .B1(n19956), .B2(n20413), .ZN(
        n19950) );
  INV_X1 U22881 ( .A(n19950), .ZN(n19952) );
  AOI22_X1 U22882 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19959), .B1(
        n20477), .B2(n19958), .ZN(n19951) );
  OAI211_X1 U22883 ( .C1(n20482), .C2(n19962), .A(n19952), .B(n19951), .ZN(
        P1_U3054) );
  OAI22_X1 U22884 ( .A1(n19962), .A2(n9758), .B1(n19956), .B2(n20418), .ZN(
        n19953) );
  INV_X1 U22885 ( .A(n19953), .ZN(n19955) );
  AOI22_X1 U22886 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19959), .B1(
        n20483), .B2(n19958), .ZN(n19954) );
  OAI211_X1 U22887 ( .C1(n20364), .C2(n19997), .A(n19955), .B(n19954), .ZN(
        P1_U3055) );
  OAI22_X1 U22888 ( .A1(n19997), .A2(n20372), .B1(n19956), .B2(n20425), .ZN(
        n19957) );
  INV_X1 U22889 ( .A(n19957), .ZN(n19961) );
  AOI22_X1 U22890 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19959), .B1(
        n20490), .B2(n19958), .ZN(n19960) );
  OAI211_X1 U22891 ( .C1(n20499), .C2(n19962), .A(n19961), .B(n19960), .ZN(
        P1_U3056) );
  NAND2_X1 U22892 ( .A1(n19964), .A2(n19963), .ZN(n19996) );
  OAI22_X1 U22893 ( .A1(n20041), .A2(n20341), .B1(n20379), .B2(n19996), .ZN(
        n19965) );
  INV_X1 U22894 ( .A(n19965), .ZN(n19977) );
  AND2_X1 U22895 ( .A1(n19966), .A2(n11860), .ZN(n20433) );
  INV_X1 U22896 ( .A(n19996), .ZN(n19967) );
  AOI21_X1 U22897 ( .B1(n19968), .B2(n20433), .A(n19967), .ZN(n19975) );
  AOI21_X1 U22898 ( .B1(n19970), .B2(n20288), .A(n19969), .ZN(n19974) );
  INV_X1 U22899 ( .A(n19974), .ZN(n19971) );
  AOI22_X1 U22900 ( .A1(n19975), .A2(n19971), .B1(n20442), .B2(n19973), .ZN(
        n19972) );
  NAND2_X1 U22901 ( .A1(n20447), .A2(n19972), .ZN(n20000) );
  OAI22_X1 U22902 ( .A1(n19975), .A2(n19974), .B1(n20437), .B2(n19973), .ZN(
        n19999) );
  AOI22_X1 U22903 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20000), .B1(
        n20439), .B2(n19999), .ZN(n19976) );
  OAI211_X1 U22904 ( .C1(n20453), .C2(n19997), .A(n19977), .B(n19976), .ZN(
        P1_U3057) );
  OAI22_X1 U22905 ( .A1(n19997), .A2(n20459), .B1(n20393), .B2(n19996), .ZN(
        n19978) );
  INV_X1 U22906 ( .A(n19978), .ZN(n19980) );
  AOI22_X1 U22907 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20000), .B1(
        n20454), .B2(n19999), .ZN(n19979) );
  OAI211_X1 U22908 ( .C1(n20345), .C2(n20041), .A(n19980), .B(n19979), .ZN(
        P1_U3058) );
  OAI22_X1 U22909 ( .A1(n20041), .A2(n20349), .B1(n20398), .B2(n19996), .ZN(
        n19981) );
  INV_X1 U22910 ( .A(n19981), .ZN(n19983) );
  AOI22_X1 U22911 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20000), .B1(
        n20460), .B2(n19999), .ZN(n19982) );
  OAI211_X1 U22912 ( .C1(n20465), .C2(n19997), .A(n19983), .B(n19982), .ZN(
        P1_U3059) );
  OAI22_X1 U22913 ( .A1(n19997), .A2(n20470), .B1(n19996), .B2(n20403), .ZN(
        n19984) );
  INV_X1 U22914 ( .A(n19984), .ZN(n19986) );
  AOI22_X1 U22915 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20000), .B1(
        n20466), .B2(n19999), .ZN(n19985) );
  OAI211_X1 U22916 ( .C1(n9756), .C2(n20041), .A(n19986), .B(n19985), .ZN(
        P1_U3060) );
  OAI22_X1 U22917 ( .A1(n20041), .A2(n20357), .B1(n19996), .B2(n20408), .ZN(
        n19987) );
  INV_X1 U22918 ( .A(n19987), .ZN(n19989) );
  AOI22_X1 U22919 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20000), .B1(
        n20471), .B2(n19999), .ZN(n19988) );
  OAI211_X1 U22920 ( .C1(n20476), .C2(n19997), .A(n19989), .B(n19988), .ZN(
        P1_U3061) );
  OAI22_X1 U22921 ( .A1(n19997), .A2(n20482), .B1(n20413), .B2(n19996), .ZN(
        n19990) );
  INV_X1 U22922 ( .A(n19990), .ZN(n19992) );
  AOI22_X1 U22923 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20000), .B1(
        n20477), .B2(n19999), .ZN(n19991) );
  OAI211_X1 U22924 ( .C1(n20361), .C2(n20041), .A(n19992), .B(n19991), .ZN(
        P1_U3062) );
  OAI22_X1 U22925 ( .A1(n20041), .A2(n20364), .B1(n19996), .B2(n20418), .ZN(
        n19993) );
  INV_X1 U22926 ( .A(n19993), .ZN(n19995) );
  AOI22_X1 U22927 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20000), .B1(
        n20483), .B2(n19999), .ZN(n19994) );
  OAI211_X1 U22928 ( .C1(n9758), .C2(n19997), .A(n19995), .B(n19994), .ZN(
        P1_U3063) );
  OAI22_X1 U22929 ( .A1(n19997), .A2(n20499), .B1(n20425), .B2(n19996), .ZN(
        n19998) );
  INV_X1 U22930 ( .A(n19998), .ZN(n20002) );
  AOI22_X1 U22931 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20000), .B1(
        n20490), .B2(n19999), .ZN(n20001) );
  OAI211_X1 U22932 ( .C1(n20372), .C2(n20041), .A(n20002), .B(n20001), .ZN(
        P1_U3064) );
  OR2_X1 U22933 ( .A1(n20286), .A2(n20074), .ZN(n20036) );
  INV_X1 U22934 ( .A(n20036), .ZN(n20012) );
  NOR2_X1 U22935 ( .A1(n13187), .A2(n20003), .ZN(n20112) );
  AND2_X1 U22936 ( .A1(n20292), .A2(n20333), .ZN(n20149) );
  NAND2_X1 U22937 ( .A1(n20112), .A2(n20149), .ZN(n20007) );
  INV_X1 U22938 ( .A(n20004), .ZN(n20005) );
  INV_X1 U22939 ( .A(n20298), .ZN(n20375) );
  NAND2_X1 U22940 ( .A1(n20005), .A2(n20375), .ZN(n20006) );
  NAND2_X1 U22941 ( .A1(n20007), .A2(n20006), .ZN(n20015) );
  AOI22_X1 U22942 ( .A1(n20440), .A2(n20012), .B1(n20439), .B2(n20015), .ZN(
        n20014) );
  INV_X1 U22943 ( .A(n20112), .ZN(n20009) );
  OAI21_X1 U22944 ( .B1(n20032), .B2(n20070), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20008) );
  OAI21_X1 U22945 ( .B1(n9622), .B2(n20009), .A(n20008), .ZN(n20011) );
  AND2_X1 U22946 ( .A1(n20010), .A2(n20222), .ZN(n20387) );
  OAI221_X1 U22947 ( .B1(n20012), .B2(n20294), .C1(n20012), .C2(n20011), .A(
        n20387), .ZN(n20038) );
  AOI22_X1 U22948 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20038), .B1(
        n20070), .B2(n20450), .ZN(n20013) );
  OAI211_X1 U22949 ( .C1(n20453), .C2(n20041), .A(n20014), .B(n20013), .ZN(
        P1_U3065) );
  INV_X1 U22950 ( .A(n20454), .ZN(n20392) );
  OAI22_X1 U22951 ( .A1(n20393), .A2(n20036), .B1(n20035), .B2(n20392), .ZN(
        n20016) );
  INV_X1 U22952 ( .A(n20016), .ZN(n20018) );
  INV_X1 U22953 ( .A(n20459), .ZN(n20342) );
  AOI22_X1 U22954 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20038), .B1(
        n20032), .B2(n20342), .ZN(n20017) );
  OAI211_X1 U22955 ( .C1(n20345), .C2(n20067), .A(n20018), .B(n20017), .ZN(
        P1_U3066) );
  INV_X1 U22956 ( .A(n20460), .ZN(n20397) );
  OAI22_X1 U22957 ( .A1(n20398), .A2(n20036), .B1(n20035), .B2(n20397), .ZN(
        n20019) );
  INV_X1 U22958 ( .A(n20019), .ZN(n20021) );
  AOI22_X1 U22959 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20038), .B1(
        n20070), .B2(n20462), .ZN(n20020) );
  OAI211_X1 U22960 ( .C1(n20465), .C2(n20041), .A(n20021), .B(n20020), .ZN(
        P1_U3067) );
  INV_X1 U22961 ( .A(n20466), .ZN(n20402) );
  OAI22_X1 U22962 ( .A1(n20403), .A2(n20036), .B1(n20035), .B2(n20402), .ZN(
        n20022) );
  INV_X1 U22963 ( .A(n20022), .ZN(n20024) );
  INV_X1 U22964 ( .A(n20470), .ZN(n20350) );
  AOI22_X1 U22965 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20038), .B1(
        n20032), .B2(n20350), .ZN(n20023) );
  OAI211_X1 U22966 ( .C1(n9756), .C2(n20067), .A(n20024), .B(n20023), .ZN(
        P1_U3068) );
  INV_X1 U22967 ( .A(n20471), .ZN(n20407) );
  OAI22_X1 U22968 ( .A1(n20408), .A2(n20036), .B1(n20035), .B2(n20407), .ZN(
        n20025) );
  INV_X1 U22969 ( .A(n20025), .ZN(n20027) );
  AOI22_X1 U22970 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20038), .B1(
        n20032), .B2(n20354), .ZN(n20026) );
  OAI211_X1 U22971 ( .C1(n20357), .C2(n20067), .A(n20027), .B(n20026), .ZN(
        P1_U3069) );
  INV_X1 U22972 ( .A(n20477), .ZN(n20412) );
  OAI22_X1 U22973 ( .A1(n20413), .A2(n20036), .B1(n20035), .B2(n20412), .ZN(
        n20028) );
  INV_X1 U22974 ( .A(n20028), .ZN(n20030) );
  INV_X1 U22975 ( .A(n20361), .ZN(n20479) );
  AOI22_X1 U22976 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20038), .B1(
        n20070), .B2(n20479), .ZN(n20029) );
  OAI211_X1 U22977 ( .C1(n20482), .C2(n20041), .A(n20030), .B(n20029), .ZN(
        P1_U3070) );
  INV_X1 U22978 ( .A(n20483), .ZN(n20417) );
  OAI22_X1 U22979 ( .A1(n20418), .A2(n20036), .B1(n20035), .B2(n20417), .ZN(
        n20031) );
  INV_X1 U22980 ( .A(n20031), .ZN(n20034) );
  AOI22_X1 U22981 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20038), .B1(
        n20032), .B2(n9757), .ZN(n20033) );
  OAI211_X1 U22982 ( .C1(n20364), .C2(n20067), .A(n20034), .B(n20033), .ZN(
        P1_U3071) );
  INV_X1 U22983 ( .A(n20490), .ZN(n20422) );
  OAI22_X1 U22984 ( .A1(n20425), .A2(n20036), .B1(n20035), .B2(n20422), .ZN(
        n20037) );
  INV_X1 U22985 ( .A(n20037), .ZN(n20040) );
  INV_X1 U22986 ( .A(n20372), .ZN(n20493) );
  AOI22_X1 U22987 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20038), .B1(
        n20070), .B2(n20493), .ZN(n20039) );
  OAI211_X1 U22988 ( .C1(n20499), .C2(n20041), .A(n20040), .B(n20039), .ZN(
        P1_U3072) );
  NOR2_X1 U22989 ( .A1(n20074), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20051) );
  INV_X1 U22990 ( .A(n20051), .ZN(n20042) );
  NOR2_X1 U22991 ( .A1(n20639), .A2(n20042), .ZN(n20069) );
  NAND2_X1 U22992 ( .A1(n20112), .A2(n20330), .ZN(n20044) );
  INV_X1 U22993 ( .A(n20069), .ZN(n20043) );
  NAND2_X1 U22994 ( .A1(n20044), .A2(n20043), .ZN(n20047) );
  NAND2_X1 U22995 ( .A1(n20047), .A2(n20333), .ZN(n20046) );
  NAND2_X1 U22996 ( .A1(n20051), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20045) );
  NAND2_X1 U22997 ( .A1(n20046), .A2(n20045), .ZN(n20068) );
  AOI22_X1 U22998 ( .A1(n20440), .A2(n20069), .B1(n20439), .B2(n20068), .ZN(
        n20053) );
  INV_X1 U22999 ( .A(n20289), .ZN(n20049) );
  INV_X1 U23000 ( .A(n20047), .ZN(n20048) );
  OAI21_X1 U23001 ( .B1(n20111), .B2(n20049), .A(n20048), .ZN(n20050) );
  OAI211_X1 U23002 ( .C1(n20288), .C2(n20051), .A(n20447), .B(n20050), .ZN(
        n20071) );
  INV_X1 U23003 ( .A(n20105), .ZN(n20064) );
  AOI22_X1 U23004 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20071), .B1(
        n20064), .B2(n20450), .ZN(n20052) );
  OAI211_X1 U23005 ( .C1(n20453), .C2(n20067), .A(n20053), .B(n20052), .ZN(
        P1_U3073) );
  AOI22_X1 U23006 ( .A1(n20455), .A2(n20069), .B1(n20454), .B2(n20068), .ZN(
        n20055) );
  AOI22_X1 U23007 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20071), .B1(
        n20070), .B2(n20342), .ZN(n20054) );
  OAI211_X1 U23008 ( .C1(n20345), .C2(n20105), .A(n20055), .B(n20054), .ZN(
        P1_U3074) );
  AOI22_X1 U23009 ( .A1(n20461), .A2(n20069), .B1(n20460), .B2(n20068), .ZN(
        n20057) );
  AOI22_X1 U23010 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20071), .B1(
        n20064), .B2(n20462), .ZN(n20056) );
  OAI211_X1 U23011 ( .C1(n20465), .C2(n20067), .A(n20057), .B(n20056), .ZN(
        P1_U3075) );
  AOI22_X1 U23012 ( .A1(n20467), .A2(n20069), .B1(n20466), .B2(n20068), .ZN(
        n20059) );
  AOI22_X1 U23013 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20071), .B1(
        n20064), .B2(n9755), .ZN(n20058) );
  OAI211_X1 U23014 ( .C1(n20470), .C2(n20067), .A(n20059), .B(n20058), .ZN(
        P1_U3076) );
  AOI22_X1 U23015 ( .A1(n20472), .A2(n20069), .B1(n20471), .B2(n20068), .ZN(
        n20061) );
  AOI22_X1 U23016 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20071), .B1(
        n20070), .B2(n20354), .ZN(n20060) );
  OAI211_X1 U23017 ( .C1(n20357), .C2(n20105), .A(n20061), .B(n20060), .ZN(
        P1_U3077) );
  AOI22_X1 U23018 ( .A1(n20478), .A2(n20069), .B1(n20477), .B2(n20068), .ZN(
        n20063) );
  AOI22_X1 U23019 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20071), .B1(
        n20070), .B2(n20358), .ZN(n20062) );
  OAI211_X1 U23020 ( .C1(n20361), .C2(n20105), .A(n20063), .B(n20062), .ZN(
        P1_U3078) );
  AOI22_X1 U23021 ( .A1(n20484), .A2(n20069), .B1(n20483), .B2(n20068), .ZN(
        n20066) );
  AOI22_X1 U23022 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20071), .B1(
        n20064), .B2(n20485), .ZN(n20065) );
  OAI211_X1 U23023 ( .C1(n9758), .C2(n20067), .A(n20066), .B(n20065), .ZN(
        P1_U3079) );
  AOI22_X1 U23024 ( .A1(n20492), .A2(n20069), .B1(n20490), .B2(n20068), .ZN(
        n20073) );
  AOI22_X1 U23025 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20071), .B1(
        n20070), .B2(n20367), .ZN(n20072) );
  OAI211_X1 U23026 ( .C1(n20372), .C2(n20105), .A(n20073), .B(n20072), .ZN(
        P1_U3080) );
  NOR2_X1 U23027 ( .A1(n20436), .A2(n20074), .ZN(n20119) );
  INV_X1 U23028 ( .A(n20119), .ZN(n20075) );
  OR2_X1 U23029 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20075), .ZN(
        n20104) );
  OAI22_X1 U23030 ( .A1(n20147), .A2(n20341), .B1(n20379), .B2(n20104), .ZN(
        n20076) );
  INV_X1 U23031 ( .A(n20076), .ZN(n20085) );
  NAND3_X1 U23032 ( .A1(n20147), .A2(n20105), .A3(n20288), .ZN(n20077) );
  NAND2_X1 U23033 ( .A1(n20077), .A2(n20289), .ZN(n20080) );
  NAND2_X1 U23034 ( .A1(n20112), .A2(n9622), .ZN(n20082) );
  AOI22_X1 U23035 ( .A1(n20080), .A2(n20082), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20104), .ZN(n20079) );
  NAND3_X1 U23036 ( .A1(n20387), .A2(n20079), .A3(n20078), .ZN(n20108) );
  INV_X1 U23037 ( .A(n20080), .ZN(n20083) );
  OAI22_X1 U23038 ( .A1(n20083), .A2(n20082), .B1(n20081), .B2(n20298), .ZN(
        n20107) );
  AOI22_X1 U23039 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20108), .B1(
        n20439), .B2(n20107), .ZN(n20084) );
  OAI211_X1 U23040 ( .C1(n20453), .C2(n20105), .A(n20085), .B(n20084), .ZN(
        P1_U3081) );
  OAI22_X1 U23041 ( .A1(n20105), .A2(n20459), .B1(n20393), .B2(n20104), .ZN(
        n20086) );
  INV_X1 U23042 ( .A(n20086), .ZN(n20088) );
  AOI22_X1 U23043 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20108), .B1(
        n20454), .B2(n20107), .ZN(n20087) );
  OAI211_X1 U23044 ( .C1(n20345), .C2(n20147), .A(n20088), .B(n20087), .ZN(
        P1_U3082) );
  OAI22_X1 U23045 ( .A1(n20105), .A2(n20465), .B1(n20398), .B2(n20104), .ZN(
        n20089) );
  INV_X1 U23046 ( .A(n20089), .ZN(n20091) );
  AOI22_X1 U23047 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20108), .B1(
        n20460), .B2(n20107), .ZN(n20090) );
  OAI211_X1 U23048 ( .C1(n20349), .C2(n20147), .A(n20091), .B(n20090), .ZN(
        P1_U3083) );
  OAI22_X1 U23049 ( .A1(n20105), .A2(n20470), .B1(n20403), .B2(n20104), .ZN(
        n20092) );
  INV_X1 U23050 ( .A(n20092), .ZN(n20094) );
  AOI22_X1 U23051 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20108), .B1(
        n20466), .B2(n20107), .ZN(n20093) );
  OAI211_X1 U23052 ( .C1(n9756), .C2(n20147), .A(n20094), .B(n20093), .ZN(
        P1_U3084) );
  OAI22_X1 U23053 ( .A1(n20147), .A2(n20357), .B1(n20408), .B2(n20104), .ZN(
        n20095) );
  INV_X1 U23054 ( .A(n20095), .ZN(n20097) );
  AOI22_X1 U23055 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20108), .B1(
        n20471), .B2(n20107), .ZN(n20096) );
  OAI211_X1 U23056 ( .C1(n20476), .C2(n20105), .A(n20097), .B(n20096), .ZN(
        P1_U3085) );
  OAI22_X1 U23057 ( .A1(n20147), .A2(n20361), .B1(n20413), .B2(n20104), .ZN(
        n20098) );
  INV_X1 U23058 ( .A(n20098), .ZN(n20100) );
  AOI22_X1 U23059 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20108), .B1(
        n20477), .B2(n20107), .ZN(n20099) );
  OAI211_X1 U23060 ( .C1(n20482), .C2(n20105), .A(n20100), .B(n20099), .ZN(
        P1_U3086) );
  OAI22_X1 U23061 ( .A1(n20147), .A2(n20364), .B1(n20418), .B2(n20104), .ZN(
        n20101) );
  INV_X1 U23062 ( .A(n20101), .ZN(n20103) );
  AOI22_X1 U23063 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20108), .B1(
        n20483), .B2(n20107), .ZN(n20102) );
  OAI211_X1 U23064 ( .C1(n9758), .C2(n20105), .A(n20103), .B(n20102), .ZN(
        P1_U3087) );
  OAI22_X1 U23065 ( .A1(n20105), .A2(n20499), .B1(n20425), .B2(n20104), .ZN(
        n20106) );
  INV_X1 U23066 ( .A(n20106), .ZN(n20110) );
  AOI22_X1 U23067 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20108), .B1(
        n20490), .B2(n20107), .ZN(n20109) );
  OAI211_X1 U23068 ( .C1(n20372), .C2(n20147), .A(n20110), .B(n20109), .ZN(
        P1_U3088) );
  NAND2_X1 U23069 ( .A1(n20112), .A2(n20433), .ZN(n20113) );
  NAND2_X1 U23070 ( .A1(n20113), .A2(n20142), .ZN(n20114) );
  NAND2_X1 U23071 ( .A1(n20114), .A2(n20333), .ZN(n20116) );
  NAND2_X1 U23072 ( .A1(n20119), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20115) );
  INV_X1 U23073 ( .A(n20439), .ZN(n20378) );
  OAI22_X1 U23074 ( .A1(n20379), .A2(n20142), .B1(n20141), .B2(n20378), .ZN(
        n20117) );
  INV_X1 U23075 ( .A(n20117), .ZN(n20121) );
  OAI21_X1 U23076 ( .B1(n20119), .B2(n20118), .A(n20447), .ZN(n20144) );
  INV_X1 U23077 ( .A(n20147), .ZN(n20138) );
  INV_X1 U23078 ( .A(n20453), .ZN(n20338) );
  AOI22_X1 U23079 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20144), .B1(
        n20138), .B2(n20338), .ZN(n20120) );
  OAI211_X1 U23080 ( .C1(n20341), .C2(n20187), .A(n20121), .B(n20120), .ZN(
        P1_U3089) );
  OAI22_X1 U23081 ( .A1(n20393), .A2(n20142), .B1(n20141), .B2(n20392), .ZN(
        n20122) );
  INV_X1 U23082 ( .A(n20122), .ZN(n20124) );
  AOI22_X1 U23083 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20144), .B1(
        n20138), .B2(n20342), .ZN(n20123) );
  OAI211_X1 U23084 ( .C1(n20345), .C2(n20187), .A(n20124), .B(n20123), .ZN(
        P1_U3090) );
  OAI22_X1 U23085 ( .A1(n20398), .A2(n20142), .B1(n20141), .B2(n20397), .ZN(
        n20125) );
  INV_X1 U23086 ( .A(n20125), .ZN(n20127) );
  INV_X1 U23087 ( .A(n20465), .ZN(n20346) );
  AOI22_X1 U23088 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20144), .B1(
        n20138), .B2(n20346), .ZN(n20126) );
  OAI211_X1 U23089 ( .C1(n20349), .C2(n20187), .A(n20127), .B(n20126), .ZN(
        P1_U3091) );
  OAI22_X1 U23090 ( .A1(n20403), .A2(n20142), .B1(n20141), .B2(n20402), .ZN(
        n20128) );
  INV_X1 U23091 ( .A(n20128), .ZN(n20130) );
  AOI22_X1 U23092 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20144), .B1(
        n20178), .B2(n9755), .ZN(n20129) );
  OAI211_X1 U23093 ( .C1(n20470), .C2(n20147), .A(n20130), .B(n20129), .ZN(
        P1_U3092) );
  OAI22_X1 U23094 ( .A1(n20408), .A2(n20142), .B1(n20141), .B2(n20407), .ZN(
        n20131) );
  INV_X1 U23095 ( .A(n20131), .ZN(n20133) );
  INV_X1 U23096 ( .A(n20357), .ZN(n20473) );
  AOI22_X1 U23097 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20144), .B1(
        n20178), .B2(n20473), .ZN(n20132) );
  OAI211_X1 U23098 ( .C1(n20476), .C2(n20147), .A(n20133), .B(n20132), .ZN(
        P1_U3093) );
  OAI22_X1 U23099 ( .A1(n20413), .A2(n20142), .B1(n20141), .B2(n20412), .ZN(
        n20134) );
  INV_X1 U23100 ( .A(n20134), .ZN(n20136) );
  AOI22_X1 U23101 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20144), .B1(
        n20178), .B2(n20479), .ZN(n20135) );
  OAI211_X1 U23102 ( .C1(n20482), .C2(n20147), .A(n20136), .B(n20135), .ZN(
        P1_U3094) );
  OAI22_X1 U23103 ( .A1(n20418), .A2(n20142), .B1(n20141), .B2(n20417), .ZN(
        n20137) );
  INV_X1 U23104 ( .A(n20137), .ZN(n20140) );
  AOI22_X1 U23105 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20144), .B1(
        n20138), .B2(n9757), .ZN(n20139) );
  OAI211_X1 U23106 ( .C1(n20364), .C2(n20187), .A(n20140), .B(n20139), .ZN(
        P1_U3095) );
  OAI22_X1 U23107 ( .A1(n20425), .A2(n20142), .B1(n20141), .B2(n20422), .ZN(
        n20143) );
  INV_X1 U23108 ( .A(n20143), .ZN(n20146) );
  AOI22_X1 U23109 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20144), .B1(
        n20178), .B2(n20493), .ZN(n20145) );
  OAI211_X1 U23110 ( .C1(n20499), .C2(n20147), .A(n20146), .B(n20145), .ZN(
        P1_U3096) );
  NAND2_X1 U23111 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20148), .ZN(
        n20253) );
  OR2_X1 U23112 ( .A1(n20286), .A2(n20253), .ZN(n20182) );
  NAND2_X1 U23113 ( .A1(n13201), .A2(n13187), .ZN(n20216) );
  INV_X1 U23114 ( .A(n20149), .ZN(n20150) );
  OR2_X1 U23115 ( .A1(n20216), .A2(n20150), .ZN(n20155) );
  NAND2_X1 U23116 ( .A1(n20151), .A2(n20218), .ZN(n20297) );
  INV_X1 U23117 ( .A(n20297), .ZN(n20153) );
  INV_X1 U23118 ( .A(n20222), .ZN(n20152) );
  NAND2_X1 U23119 ( .A1(n20153), .A2(n20152), .ZN(n20154) );
  AND2_X1 U23120 ( .A1(n20155), .A2(n20154), .ZN(n20181) );
  OAI22_X1 U23121 ( .A1(n20379), .A2(n20182), .B1(n20181), .B2(n20378), .ZN(
        n20156) );
  INV_X1 U23122 ( .A(n20156), .ZN(n20161) );
  INV_X1 U23123 ( .A(n20182), .ZN(n20159) );
  OAI21_X1 U23124 ( .B1(n20204), .B2(n20178), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20157) );
  OAI21_X1 U23125 ( .B1(n9622), .B2(n20216), .A(n20157), .ZN(n20158) );
  AOI22_X1 U23126 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20184), .B1(
        n20204), .B2(n20450), .ZN(n20160) );
  OAI211_X1 U23127 ( .C1(n20453), .C2(n20187), .A(n20161), .B(n20160), .ZN(
        P1_U3097) );
  OAI22_X1 U23128 ( .A1(n20393), .A2(n20182), .B1(n20181), .B2(n20392), .ZN(
        n20162) );
  INV_X1 U23129 ( .A(n20162), .ZN(n20164) );
  AOI22_X1 U23130 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20184), .B1(
        n20178), .B2(n20342), .ZN(n20163) );
  OAI211_X1 U23131 ( .C1(n20345), .C2(n20213), .A(n20164), .B(n20163), .ZN(
        P1_U3098) );
  OAI22_X1 U23132 ( .A1(n20398), .A2(n20182), .B1(n20181), .B2(n20397), .ZN(
        n20165) );
  INV_X1 U23133 ( .A(n20165), .ZN(n20167) );
  AOI22_X1 U23134 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20184), .B1(
        n20204), .B2(n20462), .ZN(n20166) );
  OAI211_X1 U23135 ( .C1(n20465), .C2(n20187), .A(n20167), .B(n20166), .ZN(
        P1_U3099) );
  OAI22_X1 U23136 ( .A1(n20403), .A2(n20182), .B1(n20181), .B2(n20402), .ZN(
        n20168) );
  INV_X1 U23137 ( .A(n20168), .ZN(n20170) );
  AOI22_X1 U23138 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20184), .B1(
        n20178), .B2(n20350), .ZN(n20169) );
  OAI211_X1 U23139 ( .C1(n9756), .C2(n20213), .A(n20170), .B(n20169), .ZN(
        P1_U3100) );
  OAI22_X1 U23140 ( .A1(n20408), .A2(n20182), .B1(n20181), .B2(n20407), .ZN(
        n20171) );
  INV_X1 U23141 ( .A(n20171), .ZN(n20173) );
  AOI22_X1 U23142 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20184), .B1(
        n20178), .B2(n20354), .ZN(n20172) );
  OAI211_X1 U23143 ( .C1(n20357), .C2(n20213), .A(n20173), .B(n20172), .ZN(
        P1_U3101) );
  OAI22_X1 U23144 ( .A1(n20413), .A2(n20182), .B1(n20181), .B2(n20412), .ZN(
        n20174) );
  INV_X1 U23145 ( .A(n20174), .ZN(n20176) );
  AOI22_X1 U23146 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20184), .B1(
        n20204), .B2(n20479), .ZN(n20175) );
  OAI211_X1 U23147 ( .C1(n20482), .C2(n20187), .A(n20176), .B(n20175), .ZN(
        P1_U3102) );
  OAI22_X1 U23148 ( .A1(n20418), .A2(n20182), .B1(n20181), .B2(n20417), .ZN(
        n20177) );
  INV_X1 U23149 ( .A(n20177), .ZN(n20180) );
  AOI22_X1 U23150 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20184), .B1(
        n20178), .B2(n9757), .ZN(n20179) );
  OAI211_X1 U23151 ( .C1(n20364), .C2(n20213), .A(n20180), .B(n20179), .ZN(
        P1_U3103) );
  OAI22_X1 U23152 ( .A1(n20425), .A2(n20182), .B1(n20181), .B2(n20422), .ZN(
        n20183) );
  INV_X1 U23153 ( .A(n20183), .ZN(n20186) );
  AOI22_X1 U23154 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20184), .B1(
        n20204), .B2(n20493), .ZN(n20185) );
  OAI211_X1 U23155 ( .C1(n20499), .C2(n20187), .A(n20186), .B(n20185), .ZN(
        P1_U3104) );
  NOR3_X2 U23156 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20639), .A3(
        n20253), .ZN(n20208) );
  INV_X1 U23157 ( .A(n20216), .ZN(n20254) );
  AOI21_X1 U23158 ( .B1(n20254), .B2(n20330), .A(n20208), .ZN(n20189) );
  INV_X1 U23159 ( .A(n20253), .ZN(n20255) );
  NAND2_X1 U23160 ( .A1(n20255), .A2(n20436), .ZN(n20188) );
  OAI22_X1 U23161 ( .A1(n20189), .A2(n20442), .B1(n20188), .B2(n20437), .ZN(
        n20207) );
  AOI22_X1 U23162 ( .A1(n20440), .A2(n20208), .B1(n20207), .B2(n20439), .ZN(
        n20193) );
  INV_X1 U23163 ( .A(n20188), .ZN(n20191) );
  OAI211_X1 U23164 ( .C1(n20257), .C2(n20334), .A(n20333), .B(n20189), .ZN(
        n20190) );
  OAI211_X1 U23165 ( .C1(n20288), .C2(n20191), .A(n20447), .B(n20190), .ZN(
        n20210) );
  INV_X1 U23166 ( .A(n20246), .ZN(n20209) );
  AOI22_X1 U23167 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20210), .B1(
        n20209), .B2(n20450), .ZN(n20192) );
  OAI211_X1 U23168 ( .C1(n20453), .C2(n20213), .A(n20193), .B(n20192), .ZN(
        P1_U3105) );
  AOI22_X1 U23169 ( .A1(n20455), .A2(n20208), .B1(n20207), .B2(n20454), .ZN(
        n20195) );
  AOI22_X1 U23170 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20210), .B1(
        n20204), .B2(n20342), .ZN(n20194) );
  OAI211_X1 U23171 ( .C1(n20345), .C2(n20246), .A(n20195), .B(n20194), .ZN(
        P1_U3106) );
  AOI22_X1 U23172 ( .A1(n20461), .A2(n20208), .B1(n20207), .B2(n20460), .ZN(
        n20197) );
  AOI22_X1 U23173 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20210), .B1(
        n20209), .B2(n20462), .ZN(n20196) );
  OAI211_X1 U23174 ( .C1(n20465), .C2(n20213), .A(n20197), .B(n20196), .ZN(
        P1_U3107) );
  AOI22_X1 U23175 ( .A1(n20467), .A2(n20208), .B1(n20207), .B2(n20466), .ZN(
        n20199) );
  AOI22_X1 U23176 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20210), .B1(
        n20204), .B2(n20350), .ZN(n20198) );
  OAI211_X1 U23177 ( .C1(n9756), .C2(n20246), .A(n20199), .B(n20198), .ZN(
        P1_U3108) );
  AOI22_X1 U23178 ( .A1(n20472), .A2(n20208), .B1(n20207), .B2(n20471), .ZN(
        n20201) );
  AOI22_X1 U23179 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20210), .B1(
        n20204), .B2(n20354), .ZN(n20200) );
  OAI211_X1 U23180 ( .C1(n20357), .C2(n20246), .A(n20201), .B(n20200), .ZN(
        P1_U3109) );
  AOI22_X1 U23181 ( .A1(n20478), .A2(n20208), .B1(n20207), .B2(n20477), .ZN(
        n20203) );
  AOI22_X1 U23182 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20210), .B1(
        n20209), .B2(n20479), .ZN(n20202) );
  OAI211_X1 U23183 ( .C1(n20482), .C2(n20213), .A(n20203), .B(n20202), .ZN(
        P1_U3110) );
  AOI22_X1 U23184 ( .A1(n20484), .A2(n20208), .B1(n20207), .B2(n20483), .ZN(
        n20206) );
  AOI22_X1 U23185 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20210), .B1(
        n20204), .B2(n9757), .ZN(n20205) );
  OAI211_X1 U23186 ( .C1(n20364), .C2(n20246), .A(n20206), .B(n20205), .ZN(
        P1_U3111) );
  AOI22_X1 U23187 ( .A1(n20492), .A2(n20208), .B1(n20207), .B2(n20490), .ZN(
        n20212) );
  AOI22_X1 U23188 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20210), .B1(
        n20209), .B2(n20493), .ZN(n20211) );
  OAI211_X1 U23189 ( .C1(n20499), .C2(n20213), .A(n20212), .B(n20211), .ZN(
        P1_U3112) );
  OR3_X1 U23190 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20436), .A3(
        n20253), .ZN(n20245) );
  OAI22_X1 U23191 ( .A1(n20284), .A2(n20341), .B1(n20379), .B2(n20245), .ZN(
        n20214) );
  INV_X1 U23192 ( .A(n20214), .ZN(n20226) );
  NAND3_X1 U23193 ( .A1(n20284), .A2(n20246), .A3(n20288), .ZN(n20215) );
  NAND2_X1 U23194 ( .A1(n20215), .A2(n20289), .ZN(n20221) );
  OR2_X1 U23195 ( .A1(n20216), .A2(n20292), .ZN(n20223) );
  AOI22_X1 U23196 ( .A1(n20221), .A2(n20223), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20245), .ZN(n20219) );
  OR2_X1 U23197 ( .A1(n20218), .A2(n20217), .ZN(n20373) );
  NAND2_X1 U23198 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20373), .ZN(n20386) );
  NAND3_X1 U23199 ( .A1(n20220), .A2(n20219), .A3(n20386), .ZN(n20249) );
  INV_X1 U23200 ( .A(n20221), .ZN(n20224) );
  OAI22_X1 U23201 ( .A1(n20224), .A2(n20223), .B1(n20222), .B2(n20373), .ZN(
        n20248) );
  AOI22_X1 U23202 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20249), .B1(
        n20439), .B2(n20248), .ZN(n20225) );
  OAI211_X1 U23203 ( .C1(n20453), .C2(n20246), .A(n20226), .B(n20225), .ZN(
        P1_U3113) );
  OAI22_X1 U23204 ( .A1(n20284), .A2(n20345), .B1(n20393), .B2(n20245), .ZN(
        n20227) );
  INV_X1 U23205 ( .A(n20227), .ZN(n20229) );
  AOI22_X1 U23206 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20249), .B1(
        n20454), .B2(n20248), .ZN(n20228) );
  OAI211_X1 U23207 ( .C1(n20459), .C2(n20246), .A(n20229), .B(n20228), .ZN(
        P1_U3114) );
  OAI22_X1 U23208 ( .A1(n20284), .A2(n20349), .B1(n20398), .B2(n20245), .ZN(
        n20230) );
  INV_X1 U23209 ( .A(n20230), .ZN(n20232) );
  AOI22_X1 U23210 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20249), .B1(
        n20460), .B2(n20248), .ZN(n20231) );
  OAI211_X1 U23211 ( .C1(n20465), .C2(n20246), .A(n20232), .B(n20231), .ZN(
        P1_U3115) );
  OAI22_X1 U23212 ( .A1(n20284), .A2(n9756), .B1(n20403), .B2(n20245), .ZN(
        n20233) );
  INV_X1 U23213 ( .A(n20233), .ZN(n20235) );
  AOI22_X1 U23214 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20249), .B1(
        n20466), .B2(n20248), .ZN(n20234) );
  OAI211_X1 U23215 ( .C1(n20470), .C2(n20246), .A(n20235), .B(n20234), .ZN(
        P1_U3116) );
  OAI22_X1 U23216 ( .A1(n20284), .A2(n20357), .B1(n20408), .B2(n20245), .ZN(
        n20236) );
  INV_X1 U23217 ( .A(n20236), .ZN(n20238) );
  AOI22_X1 U23218 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20249), .B1(
        n20471), .B2(n20248), .ZN(n20237) );
  OAI211_X1 U23219 ( .C1(n20476), .C2(n20246), .A(n20238), .B(n20237), .ZN(
        P1_U3117) );
  OAI22_X1 U23220 ( .A1(n20284), .A2(n20361), .B1(n20413), .B2(n20245), .ZN(
        n20239) );
  INV_X1 U23221 ( .A(n20239), .ZN(n20241) );
  AOI22_X1 U23222 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20249), .B1(
        n20477), .B2(n20248), .ZN(n20240) );
  OAI211_X1 U23223 ( .C1(n20482), .C2(n20246), .A(n20241), .B(n20240), .ZN(
        P1_U3118) );
  OAI22_X1 U23224 ( .A1(n20246), .A2(n9758), .B1(n20418), .B2(n20245), .ZN(
        n20242) );
  INV_X1 U23225 ( .A(n20242), .ZN(n20244) );
  AOI22_X1 U23226 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20249), .B1(
        n20483), .B2(n20248), .ZN(n20243) );
  OAI211_X1 U23227 ( .C1(n20364), .C2(n20284), .A(n20244), .B(n20243), .ZN(
        P1_U3119) );
  OAI22_X1 U23228 ( .A1(n20246), .A2(n20499), .B1(n20425), .B2(n20245), .ZN(
        n20247) );
  INV_X1 U23229 ( .A(n20247), .ZN(n20251) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20249), .B1(
        n20490), .B2(n20248), .ZN(n20250) );
  OAI211_X1 U23231 ( .C1(n20372), .C2(n20284), .A(n20251), .B(n20250), .ZN(
        P1_U3120) );
  NOR2_X1 U23232 ( .A1(n20432), .A2(n20253), .ZN(n20279) );
  AOI21_X1 U23233 ( .B1(n20254), .B2(n20433), .A(n20279), .ZN(n20259) );
  NAND2_X1 U23234 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20255), .ZN(
        n20256) );
  OAI22_X1 U23235 ( .A1(n20259), .A2(n20442), .B1(n20256), .B2(n20437), .ZN(
        n20278) );
  AOI22_X1 U23236 ( .A1(n20440), .A2(n20279), .B1(n20278), .B2(n20439), .ZN(
        n20264) );
  INV_X1 U23237 ( .A(n20256), .ZN(n20262) );
  INV_X1 U23238 ( .A(n20257), .ZN(n20258) );
  OAI21_X1 U23239 ( .B1(n20258), .B2(n20442), .A(n20441), .ZN(n20260) );
  NAND2_X1 U23240 ( .A1(n20260), .A2(n20259), .ZN(n20261) );
  OAI211_X1 U23241 ( .C1(n20288), .C2(n20262), .A(n20447), .B(n20261), .ZN(
        n20281) );
  INV_X1 U23242 ( .A(n20284), .ZN(n20269) );
  AOI22_X1 U23243 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20281), .B1(
        n20269), .B2(n20338), .ZN(n20263) );
  OAI211_X1 U23244 ( .C1(n20341), .C2(n20327), .A(n20264), .B(n20263), .ZN(
        P1_U3121) );
  AOI22_X1 U23245 ( .A1(n20455), .A2(n20279), .B1(n20278), .B2(n20454), .ZN(
        n20266) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20281), .B1(
        n20269), .B2(n20342), .ZN(n20265) );
  OAI211_X1 U23247 ( .C1(n20345), .C2(n20327), .A(n20266), .B(n20265), .ZN(
        P1_U3122) );
  AOI22_X1 U23248 ( .A1(n20461), .A2(n20279), .B1(n20278), .B2(n20460), .ZN(
        n20268) );
  INV_X1 U23249 ( .A(n20327), .ZN(n20280) );
  AOI22_X1 U23250 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20281), .B1(
        n20280), .B2(n20462), .ZN(n20267) );
  OAI211_X1 U23251 ( .C1(n20465), .C2(n20284), .A(n20268), .B(n20267), .ZN(
        P1_U3123) );
  AOI22_X1 U23252 ( .A1(n20467), .A2(n20279), .B1(n20278), .B2(n20466), .ZN(
        n20271) );
  AOI22_X1 U23253 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20281), .B1(
        n20269), .B2(n20350), .ZN(n20270) );
  OAI211_X1 U23254 ( .C1(n9756), .C2(n20327), .A(n20271), .B(n20270), .ZN(
        P1_U3124) );
  AOI22_X1 U23255 ( .A1(n20472), .A2(n20279), .B1(n20278), .B2(n20471), .ZN(
        n20273) );
  AOI22_X1 U23256 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20281), .B1(
        n20280), .B2(n20473), .ZN(n20272) );
  OAI211_X1 U23257 ( .C1(n20476), .C2(n20284), .A(n20273), .B(n20272), .ZN(
        P1_U3125) );
  AOI22_X1 U23258 ( .A1(n20478), .A2(n20279), .B1(n20278), .B2(n20477), .ZN(
        n20275) );
  AOI22_X1 U23259 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20281), .B1(
        n20280), .B2(n20479), .ZN(n20274) );
  OAI211_X1 U23260 ( .C1(n20482), .C2(n20284), .A(n20275), .B(n20274), .ZN(
        P1_U3126) );
  AOI22_X1 U23261 ( .A1(n20484), .A2(n20279), .B1(n20278), .B2(n20483), .ZN(
        n20277) );
  AOI22_X1 U23262 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20281), .B1(
        n20280), .B2(n20485), .ZN(n20276) );
  OAI211_X1 U23263 ( .C1(n9758), .C2(n20284), .A(n20277), .B(n20276), .ZN(
        P1_U3127) );
  AOI22_X1 U23264 ( .A1(n20492), .A2(n20279), .B1(n20278), .B2(n20490), .ZN(
        n20283) );
  AOI22_X1 U23265 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20281), .B1(
        n20280), .B2(n20493), .ZN(n20282) );
  OAI211_X1 U23266 ( .C1(n20499), .C2(n20284), .A(n20283), .B(n20282), .ZN(
        P1_U3128) );
  NAND2_X1 U23267 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20435) );
  OR2_X1 U23268 ( .A1(n20286), .A2(n20435), .ZN(n20321) );
  OAI22_X1 U23269 ( .A1(n20337), .A2(n20341), .B1(n20379), .B2(n20321), .ZN(
        n20287) );
  INV_X1 U23270 ( .A(n20287), .ZN(n20302) );
  INV_X1 U23271 ( .A(n20321), .ZN(n20295) );
  NAND3_X1 U23272 ( .A1(n20327), .A2(n20288), .A3(n20337), .ZN(n20290) );
  NAND2_X1 U23273 ( .A1(n20290), .A2(n20289), .ZN(n20296) );
  NOR2_X1 U23274 ( .A1(n13187), .A2(n20291), .ZN(n20434) );
  NAND2_X1 U23275 ( .A1(n20434), .A2(n20292), .ZN(n20299) );
  AOI22_X1 U23276 ( .A1(n20296), .A2(n20299), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20297), .ZN(n20293) );
  OAI211_X1 U23277 ( .C1(n20295), .C2(n20294), .A(n20387), .B(n20293), .ZN(
        n20324) );
  INV_X1 U23278 ( .A(n20296), .ZN(n20300) );
  OAI22_X1 U23279 ( .A1(n20300), .A2(n20299), .B1(n20298), .B2(n20297), .ZN(
        n20323) );
  AOI22_X1 U23280 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20324), .B1(
        n20439), .B2(n20323), .ZN(n20301) );
  OAI211_X1 U23281 ( .C1(n20453), .C2(n20327), .A(n20302), .B(n20301), .ZN(
        P1_U3129) );
  OAI22_X1 U23282 ( .A1(n20337), .A2(n20345), .B1(n20393), .B2(n20321), .ZN(
        n20303) );
  INV_X1 U23283 ( .A(n20303), .ZN(n20305) );
  AOI22_X1 U23284 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20324), .B1(
        n20454), .B2(n20323), .ZN(n20304) );
  OAI211_X1 U23285 ( .C1(n20459), .C2(n20327), .A(n20305), .B(n20304), .ZN(
        P1_U3130) );
  OAI22_X1 U23286 ( .A1(n20337), .A2(n20349), .B1(n20398), .B2(n20321), .ZN(
        n20306) );
  INV_X1 U23287 ( .A(n20306), .ZN(n20308) );
  AOI22_X1 U23288 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20324), .B1(
        n20460), .B2(n20323), .ZN(n20307) );
  OAI211_X1 U23289 ( .C1(n20465), .C2(n20327), .A(n20308), .B(n20307), .ZN(
        P1_U3131) );
  OAI22_X1 U23290 ( .A1(n20337), .A2(n9756), .B1(n20403), .B2(n20321), .ZN(
        n20309) );
  INV_X1 U23291 ( .A(n20309), .ZN(n20311) );
  AOI22_X1 U23292 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20324), .B1(
        n20466), .B2(n20323), .ZN(n20310) );
  OAI211_X1 U23293 ( .C1(n20470), .C2(n20327), .A(n20311), .B(n20310), .ZN(
        P1_U3132) );
  OAI22_X1 U23294 ( .A1(n20337), .A2(n20357), .B1(n20408), .B2(n20321), .ZN(
        n20312) );
  INV_X1 U23295 ( .A(n20312), .ZN(n20314) );
  AOI22_X1 U23296 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20324), .B1(
        n20471), .B2(n20323), .ZN(n20313) );
  OAI211_X1 U23297 ( .C1(n20476), .C2(n20327), .A(n20314), .B(n20313), .ZN(
        P1_U3133) );
  OAI22_X1 U23298 ( .A1(n20337), .A2(n20361), .B1(n20413), .B2(n20321), .ZN(
        n20315) );
  INV_X1 U23299 ( .A(n20315), .ZN(n20317) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20324), .B1(
        n20477), .B2(n20323), .ZN(n20316) );
  OAI211_X1 U23301 ( .C1(n20482), .C2(n20327), .A(n20317), .B(n20316), .ZN(
        P1_U3134) );
  OAI22_X1 U23302 ( .A1(n20337), .A2(n20364), .B1(n20418), .B2(n20321), .ZN(
        n20318) );
  INV_X1 U23303 ( .A(n20318), .ZN(n20320) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20324), .B1(
        n20483), .B2(n20323), .ZN(n20319) );
  OAI211_X1 U23305 ( .C1(n9758), .C2(n20327), .A(n20320), .B(n20319), .ZN(
        P1_U3135) );
  OAI22_X1 U23306 ( .A1(n20337), .A2(n20372), .B1(n20425), .B2(n20321), .ZN(
        n20322) );
  INV_X1 U23307 ( .A(n20322), .ZN(n20326) );
  AOI22_X1 U23308 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20324), .B1(
        n20490), .B2(n20323), .ZN(n20325) );
  OAI211_X1 U23309 ( .C1(n20499), .C2(n20327), .A(n20326), .B(n20325), .ZN(
        P1_U3136) );
  INV_X1 U23310 ( .A(n20382), .ZN(n20443) );
  INV_X1 U23311 ( .A(n20328), .ZN(n20329) );
  NOR3_X2 U23312 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20639), .A3(
        n20435), .ZN(n20366) );
  AOI21_X1 U23313 ( .B1(n20434), .B2(n20330), .A(n20366), .ZN(n20332) );
  NOR2_X1 U23314 ( .A1(n20435), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20336) );
  INV_X1 U23315 ( .A(n20336), .ZN(n20331) );
  OAI22_X1 U23316 ( .A1(n20332), .A2(n20442), .B1(n20331), .B2(n20437), .ZN(
        n20365) );
  AOI22_X1 U23317 ( .A1(n20440), .A2(n20366), .B1(n20439), .B2(n20365), .ZN(
        n20340) );
  OAI211_X1 U23318 ( .C1(n20382), .C2(n20334), .A(n20333), .B(n20332), .ZN(
        n20335) );
  OAI211_X1 U23319 ( .C1(n20288), .C2(n20336), .A(n20447), .B(n20335), .ZN(
        n20369) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20369), .B1(
        n20368), .B2(n20338), .ZN(n20339) );
  OAI211_X1 U23321 ( .C1(n20341), .C2(n20431), .A(n20340), .B(n20339), .ZN(
        P1_U3137) );
  AOI22_X1 U23322 ( .A1(n20455), .A2(n20366), .B1(n20454), .B2(n20365), .ZN(
        n20344) );
  AOI22_X1 U23323 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20369), .B1(
        n20368), .B2(n20342), .ZN(n20343) );
  OAI211_X1 U23324 ( .C1(n20345), .C2(n20431), .A(n20344), .B(n20343), .ZN(
        P1_U3138) );
  AOI22_X1 U23325 ( .A1(n20461), .A2(n20366), .B1(n20460), .B2(n20365), .ZN(
        n20348) );
  AOI22_X1 U23326 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20369), .B1(
        n20368), .B2(n20346), .ZN(n20347) );
  OAI211_X1 U23327 ( .C1(n20349), .C2(n20431), .A(n20348), .B(n20347), .ZN(
        P1_U3139) );
  AOI22_X1 U23328 ( .A1(n20467), .A2(n20366), .B1(n20466), .B2(n20365), .ZN(
        n20352) );
  AOI22_X1 U23329 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20369), .B1(
        n20368), .B2(n20350), .ZN(n20351) );
  OAI211_X1 U23330 ( .C1(n9756), .C2(n20431), .A(n20352), .B(n20351), .ZN(
        P1_U3140) );
  AOI22_X1 U23331 ( .A1(n20472), .A2(n20366), .B1(n20471), .B2(n20365), .ZN(
        n20356) );
  AOI22_X1 U23332 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20369), .B1(
        n20368), .B2(n20354), .ZN(n20355) );
  OAI211_X1 U23333 ( .C1(n20357), .C2(n20431), .A(n20356), .B(n20355), .ZN(
        P1_U3141) );
  AOI22_X1 U23334 ( .A1(n20478), .A2(n20366), .B1(n20477), .B2(n20365), .ZN(
        n20360) );
  AOI22_X1 U23335 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20369), .B1(
        n20368), .B2(n20358), .ZN(n20359) );
  OAI211_X1 U23336 ( .C1(n20361), .C2(n20431), .A(n20360), .B(n20359), .ZN(
        P1_U3142) );
  AOI22_X1 U23337 ( .A1(n20484), .A2(n20366), .B1(n20483), .B2(n20365), .ZN(
        n20363) );
  AOI22_X1 U23338 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20369), .B1(
        n20368), .B2(n9757), .ZN(n20362) );
  OAI211_X1 U23339 ( .C1(n20364), .C2(n20431), .A(n20363), .B(n20362), .ZN(
        P1_U3143) );
  AOI22_X1 U23340 ( .A1(n20492), .A2(n20366), .B1(n20490), .B2(n20365), .ZN(
        n20371) );
  AOI22_X1 U23341 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20369), .B1(
        n20368), .B2(n20367), .ZN(n20370) );
  OAI211_X1 U23342 ( .C1(n20372), .C2(n20431), .A(n20371), .B(n20370), .ZN(
        P1_U3144) );
  NOR3_X1 U23343 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20436), .A3(
        n20435), .ZN(n20389) );
  INV_X1 U23344 ( .A(n20389), .ZN(n20424) );
  NAND2_X1 U23345 ( .A1(n20434), .A2(n9622), .ZN(n20384) );
  OR2_X1 U23346 ( .A1(n20384), .A2(n20442), .ZN(n20377) );
  INV_X1 U23347 ( .A(n20373), .ZN(n20374) );
  NAND2_X1 U23348 ( .A1(n20375), .A2(n20374), .ZN(n20376) );
  OAI22_X1 U23349 ( .A1(n20379), .A2(n20424), .B1(n20423), .B2(n20378), .ZN(
        n20380) );
  INV_X1 U23350 ( .A(n20380), .ZN(n20391) );
  INV_X1 U23351 ( .A(n20431), .ZN(n20383) );
  OAI21_X1 U23352 ( .B1(n20383), .B2(n20427), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20385) );
  AOI21_X1 U23353 ( .B1(n20385), .B2(n20384), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20388) );
  AOI22_X1 U23354 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20450), .ZN(n20390) );
  OAI211_X1 U23355 ( .C1(n20453), .C2(n20431), .A(n20391), .B(n20390), .ZN(
        P1_U3145) );
  OAI22_X1 U23356 ( .A1(n20393), .A2(n20424), .B1(n20423), .B2(n20392), .ZN(
        n20394) );
  INV_X1 U23357 ( .A(n20394), .ZN(n20396) );
  AOI22_X1 U23358 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20456), .ZN(n20395) );
  OAI211_X1 U23359 ( .C1(n20459), .C2(n20431), .A(n20396), .B(n20395), .ZN(
        P1_U3146) );
  OAI22_X1 U23360 ( .A1(n20398), .A2(n20424), .B1(n20423), .B2(n20397), .ZN(
        n20399) );
  INV_X1 U23361 ( .A(n20399), .ZN(n20401) );
  AOI22_X1 U23362 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20462), .ZN(n20400) );
  OAI211_X1 U23363 ( .C1(n20465), .C2(n20431), .A(n20401), .B(n20400), .ZN(
        P1_U3147) );
  OAI22_X1 U23364 ( .A1(n20403), .A2(n20424), .B1(n20423), .B2(n20402), .ZN(
        n20404) );
  INV_X1 U23365 ( .A(n20404), .ZN(n20406) );
  AOI22_X1 U23366 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n9755), .ZN(n20405) );
  OAI211_X1 U23367 ( .C1(n20470), .C2(n20431), .A(n20406), .B(n20405), .ZN(
        P1_U3148) );
  OAI22_X1 U23368 ( .A1(n20408), .A2(n20424), .B1(n20423), .B2(n20407), .ZN(
        n20409) );
  INV_X1 U23369 ( .A(n20409), .ZN(n20411) );
  AOI22_X1 U23370 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20473), .ZN(n20410) );
  OAI211_X1 U23371 ( .C1(n20476), .C2(n20431), .A(n20411), .B(n20410), .ZN(
        P1_U3149) );
  OAI22_X1 U23372 ( .A1(n20413), .A2(n20424), .B1(n20423), .B2(n20412), .ZN(
        n20414) );
  INV_X1 U23373 ( .A(n20414), .ZN(n20416) );
  AOI22_X1 U23374 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20479), .ZN(n20415) );
  OAI211_X1 U23375 ( .C1(n20482), .C2(n20431), .A(n20416), .B(n20415), .ZN(
        P1_U3150) );
  OAI22_X1 U23376 ( .A1(n20418), .A2(n20424), .B1(n20423), .B2(n20417), .ZN(
        n20419) );
  INV_X1 U23377 ( .A(n20419), .ZN(n20421) );
  AOI22_X1 U23378 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20485), .ZN(n20420) );
  OAI211_X1 U23379 ( .C1(n9758), .C2(n20431), .A(n20421), .B(n20420), .ZN(
        P1_U3151) );
  OAI22_X1 U23380 ( .A1(n20425), .A2(n20424), .B1(n20423), .B2(n20422), .ZN(
        n20426) );
  INV_X1 U23381 ( .A(n20426), .ZN(n20430) );
  AOI22_X1 U23382 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20493), .ZN(n20429) );
  OAI211_X1 U23383 ( .C1(n20499), .C2(n20431), .A(n20430), .B(n20429), .ZN(
        P1_U3152) );
  NOR2_X1 U23384 ( .A1(n20432), .A2(n20435), .ZN(n20491) );
  AOI21_X1 U23385 ( .B1(n20434), .B2(n20433), .A(n20491), .ZN(n20444) );
  NOR2_X1 U23386 ( .A1(n20436), .A2(n20435), .ZN(n20448) );
  INV_X1 U23387 ( .A(n20448), .ZN(n20438) );
  OAI22_X1 U23388 ( .A1(n20444), .A2(n20442), .B1(n20438), .B2(n20437), .ZN(
        n20489) );
  AOI22_X1 U23389 ( .A1(n20440), .A2(n20491), .B1(n20439), .B2(n20489), .ZN(
        n20452) );
  OAI21_X1 U23390 ( .B1(n20443), .B2(n20442), .A(n20441), .ZN(n20445) );
  NAND2_X1 U23391 ( .A1(n20445), .A2(n20444), .ZN(n20446) );
  OAI211_X1 U23392 ( .C1(n20333), .C2(n20448), .A(n20447), .B(n20446), .ZN(
        n20495) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20495), .B1(
        n20494), .B2(n20450), .ZN(n20451) );
  OAI211_X1 U23394 ( .C1(n20453), .C2(n20498), .A(n20452), .B(n20451), .ZN(
        P1_U3153) );
  AOI22_X1 U23395 ( .A1(n20455), .A2(n20491), .B1(n20454), .B2(n20489), .ZN(
        n20458) );
  AOI22_X1 U23396 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20495), .B1(
        n20494), .B2(n20456), .ZN(n20457) );
  OAI211_X1 U23397 ( .C1(n20459), .C2(n20498), .A(n20458), .B(n20457), .ZN(
        P1_U3154) );
  AOI22_X1 U23398 ( .A1(n20461), .A2(n20491), .B1(n20460), .B2(n20489), .ZN(
        n20464) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20495), .B1(
        n20494), .B2(n20462), .ZN(n20463) );
  OAI211_X1 U23400 ( .C1(n20465), .C2(n20498), .A(n20464), .B(n20463), .ZN(
        P1_U3155) );
  AOI22_X1 U23401 ( .A1(n20467), .A2(n20491), .B1(n20466), .B2(n20489), .ZN(
        n20469) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20495), .B1(
        n20494), .B2(n9755), .ZN(n20468) );
  OAI211_X1 U23403 ( .C1(n20470), .C2(n20498), .A(n20469), .B(n20468), .ZN(
        P1_U3156) );
  AOI22_X1 U23404 ( .A1(n20472), .A2(n20491), .B1(n20471), .B2(n20489), .ZN(
        n20475) );
  AOI22_X1 U23405 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20495), .B1(
        n20494), .B2(n20473), .ZN(n20474) );
  OAI211_X1 U23406 ( .C1(n20476), .C2(n20498), .A(n20475), .B(n20474), .ZN(
        P1_U3157) );
  AOI22_X1 U23407 ( .A1(n20478), .A2(n20491), .B1(n20477), .B2(n20489), .ZN(
        n20481) );
  AOI22_X1 U23408 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20495), .B1(
        n20494), .B2(n20479), .ZN(n20480) );
  OAI211_X1 U23409 ( .C1(n20482), .C2(n20498), .A(n20481), .B(n20480), .ZN(
        P1_U3158) );
  AOI22_X1 U23410 ( .A1(n20484), .A2(n20491), .B1(n20483), .B2(n20489), .ZN(
        n20487) );
  AOI22_X1 U23411 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20495), .B1(
        n20494), .B2(n20485), .ZN(n20486) );
  OAI211_X1 U23412 ( .C1(n9758), .C2(n20498), .A(n20487), .B(n20486), .ZN(
        P1_U3159) );
  AOI22_X1 U23413 ( .A1(n20492), .A2(n20491), .B1(n20490), .B2(n20489), .ZN(
        n20497) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20495), .B1(
        n20494), .B2(n20493), .ZN(n20496) );
  OAI211_X1 U23415 ( .C1(n20499), .C2(n20498), .A(n20497), .B(n20496), .ZN(
        P1_U3160) );
  OR2_X1 U23416 ( .A1(n20501), .A2(n20500), .ZN(P1_U3163) );
  AND2_X1 U23417 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20583), .ZN(
        P1_U3164) );
  AND2_X1 U23418 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20583), .ZN(
        P1_U3165) );
  AND2_X1 U23419 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20583), .ZN(
        P1_U3166) );
  AND2_X1 U23420 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20583), .ZN(
        P1_U3167) );
  AND2_X1 U23421 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20583), .ZN(
        P1_U3168) );
  AND2_X1 U23422 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20583), .ZN(
        P1_U3169) );
  AND2_X1 U23423 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20583), .ZN(
        P1_U3170) );
  AND2_X1 U23424 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20583), .ZN(
        P1_U3171) );
  AND2_X1 U23425 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20583), .ZN(
        P1_U3172) );
  AND2_X1 U23426 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20583), .ZN(
        P1_U3173) );
  AND2_X1 U23427 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20583), .ZN(
        P1_U3174) );
  INV_X1 U23428 ( .A(P1_DATAWIDTH_REG_20__SCAN_IN), .ZN(n20648) );
  NOR2_X1 U23429 ( .A1(n20587), .A2(n20648), .ZN(P1_U3175) );
  AND2_X1 U23430 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20583), .ZN(
        P1_U3176) );
  AND2_X1 U23431 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20583), .ZN(
        P1_U3177) );
  AND2_X1 U23432 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20583), .ZN(
        P1_U3178) );
  AND2_X1 U23433 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20583), .ZN(
        P1_U3179) );
  AND2_X1 U23434 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20583), .ZN(
        P1_U3180) );
  AND2_X1 U23435 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20583), .ZN(
        P1_U3181) );
  AND2_X1 U23436 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20583), .ZN(
        P1_U3182) );
  AND2_X1 U23437 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20583), .ZN(
        P1_U3183) );
  AND2_X1 U23438 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20583), .ZN(
        P1_U3184) );
  AND2_X1 U23439 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20583), .ZN(
        P1_U3185) );
  AND2_X1 U23440 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20583), .ZN(P1_U3186) );
  AND2_X1 U23441 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20583), .ZN(P1_U3187) );
  AND2_X1 U23442 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20583), .ZN(P1_U3188) );
  AND2_X1 U23443 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20583), .ZN(P1_U3189) );
  AND2_X1 U23444 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20583), .ZN(P1_U3190) );
  AND2_X1 U23445 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20583), .ZN(P1_U3191) );
  AND2_X1 U23446 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20583), .ZN(P1_U3192) );
  AND2_X1 U23447 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20583), .ZN(P1_U3193) );
  AOI21_X1 U23448 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20507), .A(n20504), 
        .ZN(n20515) );
  NOR2_X1 U23449 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20502) );
  NOR2_X1 U23450 ( .A1(n20502), .A2(n20782), .ZN(n20503) );
  AOI211_X1 U23451 ( .C1(NA), .C2(n20504), .A(n20503), .B(n20508), .ZN(n20505)
         );
  OAI22_X1 U23452 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20515), .B1(n20630), 
        .B2(n20505), .ZN(P1_U3194) );
  AOI21_X1 U23453 ( .B1(n20507), .B2(n20513), .A(n20506), .ZN(n20517) );
  OAI211_X1 U23454 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20508), .A(
        P1_STATE_REG_0__SCAN_IN), .B(HOLD), .ZN(n20516) );
  NOR2_X1 U23455 ( .A1(n20510), .A2(n20509), .ZN(n20511) );
  AOI221_X1 U23456 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20513), .C1(n20512), 
        .C2(n20513), .A(n20511), .ZN(n20514) );
  OAI22_X1 U23457 ( .A1(n20517), .A2(n20516), .B1(n20515), .B2(n20514), .ZN(
        P1_U3196) );
  NAND2_X1 U23458 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20630), .ZN(n20571) );
  NOR2_X1 U23459 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20617), .ZN(n20569) );
  AOI22_X1 U23460 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n20617), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20569), .ZN(n20518) );
  OAI21_X1 U23461 ( .B1(n20609), .B2(n20571), .A(n20518), .ZN(P1_U3197) );
  AOI22_X1 U23462 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20617), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n20569), .ZN(n20519) );
  OAI21_X1 U23463 ( .B1(n19706), .B2(n20571), .A(n20519), .ZN(P1_U3198) );
  INV_X1 U23464 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20521) );
  INV_X1 U23465 ( .A(n20569), .ZN(n20575) );
  OAI222_X1 U23466 ( .A1(n20571), .A2(n20521), .B1(n20520), .B2(n20630), .C1(
        n20522), .C2(n20575), .ZN(P1_U3199) );
  INV_X1 U23467 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20523) );
  OAI222_X1 U23468 ( .A1(n20575), .A2(n20525), .B1(n20523), .B2(n20630), .C1(
        n20522), .C2(n20571), .ZN(P1_U3200) );
  INV_X1 U23469 ( .A(n20571), .ZN(n20573) );
  INV_X1 U23470 ( .A(n20573), .ZN(n20566) );
  INV_X1 U23471 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20524) );
  OAI222_X1 U23472 ( .A1(n20566), .A2(n20525), .B1(n20524), .B2(n20630), .C1(
        n20527), .C2(n20575), .ZN(P1_U3201) );
  INV_X1 U23473 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20526) );
  OAI222_X1 U23474 ( .A1(n20566), .A2(n20527), .B1(n20526), .B2(n20630), .C1(
        n20529), .C2(n20575), .ZN(P1_U3202) );
  INV_X1 U23475 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20528) );
  OAI222_X1 U23476 ( .A1(n20566), .A2(n20529), .B1(n20528), .B2(n20630), .C1(
        n20530), .C2(n20575), .ZN(P1_U3203) );
  INV_X1 U23477 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20531) );
  OAI222_X1 U23478 ( .A1(n20575), .A2(n13588), .B1(n20531), .B2(n20630), .C1(
        n20530), .C2(n20571), .ZN(P1_U3204) );
  INV_X1 U23479 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20532) );
  OAI222_X1 U23480 ( .A1(n20566), .A2(n13588), .B1(n20532), .B2(n20630), .C1(
        n20534), .C2(n20575), .ZN(P1_U3205) );
  INV_X1 U23481 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20533) );
  OAI222_X1 U23482 ( .A1(n20566), .A2(n20534), .B1(n20533), .B2(n20630), .C1(
        n20536), .C2(n20575), .ZN(P1_U3206) );
  INV_X1 U23483 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20535) );
  OAI222_X1 U23484 ( .A1(n20566), .A2(n20536), .B1(n20535), .B2(n20630), .C1(
        n20538), .C2(n20575), .ZN(P1_U3207) );
  AOI22_X1 U23485 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20617), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(n20569), .ZN(n20537) );
  OAI21_X1 U23486 ( .B1(n20538), .B2(n20571), .A(n20537), .ZN(P1_U3208) );
  AOI22_X1 U23487 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20617), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(n20573), .ZN(n20539) );
  OAI21_X1 U23488 ( .B1(n20540), .B2(n20575), .A(n20539), .ZN(P1_U3209) );
  INV_X1 U23489 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20541) );
  OAI222_X1 U23490 ( .A1(n20575), .A2(n20542), .B1(n20541), .B2(n20630), .C1(
        n20540), .C2(n20571), .ZN(P1_U3210) );
  INV_X1 U23491 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20543) );
  OAI222_X1 U23492 ( .A1(n20575), .A2(n20545), .B1(n20543), .B2(n20630), .C1(
        n20542), .C2(n20571), .ZN(P1_U3211) );
  AOI22_X1 U23493 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20617), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20569), .ZN(n20544) );
  OAI21_X1 U23494 ( .B1(n20545), .B2(n20571), .A(n20544), .ZN(P1_U3212) );
  INV_X1 U23495 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20548) );
  AOI22_X1 U23496 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20617), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20573), .ZN(n20546) );
  OAI21_X1 U23497 ( .B1(n20548), .B2(n20575), .A(n20546), .ZN(P1_U3213) );
  AOI22_X1 U23498 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20617), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20569), .ZN(n20547) );
  OAI21_X1 U23499 ( .B1(n20548), .B2(n20571), .A(n20547), .ZN(P1_U3214) );
  AOI22_X1 U23500 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20617), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20573), .ZN(n20549) );
  OAI21_X1 U23501 ( .B1(n20550), .B2(n20575), .A(n20549), .ZN(P1_U3215) );
  INV_X1 U23502 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20551) );
  OAI222_X1 U23503 ( .A1(n20575), .A2(n20553), .B1(n20551), .B2(n20630), .C1(
        n20550), .C2(n20571), .ZN(P1_U3216) );
  INV_X1 U23504 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20552) );
  OAI222_X1 U23505 ( .A1(n20566), .A2(n20553), .B1(n20552), .B2(n20630), .C1(
        n20555), .C2(n20575), .ZN(P1_U3217) );
  INV_X1 U23506 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20554) );
  OAI222_X1 U23507 ( .A1(n20566), .A2(n20555), .B1(n20554), .B2(n20630), .C1(
        n20557), .C2(n20575), .ZN(P1_U3218) );
  INV_X1 U23508 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20556) );
  OAI222_X1 U23509 ( .A1(n20566), .A2(n20557), .B1(n20556), .B2(n20630), .C1(
        n20558), .C2(n20575), .ZN(P1_U3219) );
  INV_X1 U23510 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20559) );
  OAI222_X1 U23511 ( .A1(n20575), .A2(n20561), .B1(n20559), .B2(n20630), .C1(
        n20558), .C2(n20571), .ZN(P1_U3220) );
  INV_X1 U23512 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20560) );
  OAI222_X1 U23513 ( .A1(n20566), .A2(n20561), .B1(n20560), .B2(n20630), .C1(
        n20563), .C2(n20575), .ZN(P1_U3221) );
  INV_X1 U23514 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20562) );
  OAI222_X1 U23515 ( .A1(n20566), .A2(n20563), .B1(n20562), .B2(n20630), .C1(
        n20565), .C2(n20575), .ZN(P1_U3222) );
  INV_X1 U23516 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20564) );
  OAI222_X1 U23517 ( .A1(n20566), .A2(n20565), .B1(n20564), .B2(n20630), .C1(
        n20568), .C2(n20575), .ZN(P1_U3223) );
  INV_X1 U23518 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20567) );
  OAI222_X1 U23519 ( .A1(n20571), .A2(n20568), .B1(n20567), .B2(n20630), .C1(
        n20572), .C2(n20575), .ZN(P1_U3224) );
  AOI22_X1 U23520 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20569), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20617), .ZN(n20570) );
  OAI21_X1 U23521 ( .B1(n20572), .B2(n20571), .A(n20570), .ZN(P1_U3225) );
  AOI22_X1 U23522 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20573), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20617), .ZN(n20574) );
  OAI21_X1 U23523 ( .B1(n20576), .B2(n20575), .A(n20574), .ZN(P1_U3226) );
  INV_X1 U23524 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20775) );
  AOI22_X1 U23525 ( .A1(n20630), .A2(n20577), .B1(n20775), .B2(n20617), .ZN(
        P1_U3458) );
  INV_X1 U23526 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20612) );
  INV_X1 U23527 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20578) );
  AOI22_X1 U23528 ( .A1(n20630), .A2(n20612), .B1(n20578), .B2(n20617), .ZN(
        P1_U3459) );
  INV_X1 U23529 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20579) );
  AOI22_X1 U23530 ( .A1(n20630), .A2(n20580), .B1(n20579), .B2(n20617), .ZN(
        P1_U3460) );
  INV_X1 U23531 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20615) );
  INV_X1 U23532 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20581) );
  AOI22_X1 U23533 ( .A1(n20630), .A2(n20615), .B1(n20581), .B2(n20617), .ZN(
        P1_U3461) );
  INV_X1 U23534 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20584) );
  INV_X1 U23535 ( .A(n20585), .ZN(n20582) );
  AOI21_X1 U23536 ( .B1(n20584), .B2(n20583), .A(n20582), .ZN(P1_U3464) );
  OAI21_X1 U23537 ( .B1(n20587), .B2(n20586), .A(n20585), .ZN(P1_U3465) );
  INV_X1 U23538 ( .A(n20588), .ZN(n20592) );
  INV_X1 U23539 ( .A(n20589), .ZN(n20590) );
  OAI22_X1 U23540 ( .A1(n20592), .A2(n20591), .B1(n20590), .B2(n20597), .ZN(
        n20593) );
  MUX2_X1 U23541 ( .A(n20593), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n20605), .Z(P1_U3469) );
  INV_X1 U23542 ( .A(n20594), .ZN(n20603) );
  NAND2_X1 U23543 ( .A1(n20596), .A2(n20595), .ZN(n20602) );
  INV_X1 U23544 ( .A(n20597), .ZN(n20598) );
  NAND3_X1 U23545 ( .A1(n20600), .A2(n20599), .A3(n20598), .ZN(n20601) );
  OAI211_X1 U23546 ( .C1(n20604), .C2(n20603), .A(n20602), .B(n20601), .ZN(
        n20606) );
  OAI22_X1 U23547 ( .A1(n20607), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n20606), .B2(n20605), .ZN(n20608) );
  INV_X1 U23548 ( .A(n20608), .ZN(P1_U3473) );
  AOI21_X1 U23549 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20610) );
  AOI22_X1 U23550 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20610), .B2(n20609), .ZN(n20613) );
  AOI22_X1 U23551 ( .A1(n20616), .A2(n20613), .B1(n20612), .B2(n20611), .ZN(
        P1_U3481) );
  OAI21_X1 U23552 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20616), .ZN(n20614) );
  OAI21_X1 U23553 ( .B1(n20616), .B2(n20615), .A(n20614), .ZN(P1_U3482) );
  AOI22_X1 U23554 ( .A1(n20630), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20618), 
        .B2(n20617), .ZN(P1_U3483) );
  OAI21_X1 U23555 ( .B1(n20619), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20622) );
  OAI21_X1 U23556 ( .B1(n20622), .B2(n20621), .A(n20620), .ZN(n20629) );
  AOI211_X1 U23557 ( .C1(n20626), .C2(n20625), .A(n20624), .B(n20623), .ZN(
        n20628) );
  NAND2_X1 U23558 ( .A1(n20628), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20627) );
  OAI21_X1 U23559 ( .B1(n20629), .B2(n20628), .A(n20627), .ZN(P1_U3485) );
  MUX2_X1 U23560 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20630), .Z(P1_U3486) );
  AOI22_X1 U23561 ( .A1(n20633), .A2(keyinput124), .B1(keyinput106), .B2(
        n20632), .ZN(n20631) );
  OAI221_X1 U23562 ( .B1(n20633), .B2(keyinput124), .C1(n20632), .C2(
        keyinput106), .A(n20631), .ZN(n20643) );
  INV_X1 U23563 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n20781) );
  AOI22_X1 U23564 ( .A1(n20781), .A2(keyinput127), .B1(keyinput117), .B2(
        n20635), .ZN(n20634) );
  OAI221_X1 U23565 ( .B1(n20781), .B2(keyinput127), .C1(n20635), .C2(
        keyinput117), .A(n20634), .ZN(n20642) );
  INV_X1 U23566 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n20637) );
  AOI22_X1 U23567 ( .A1(n20637), .A2(keyinput99), .B1(keyinput89), .B2(n20762), 
        .ZN(n20636) );
  OAI221_X1 U23568 ( .B1(n20637), .B2(keyinput99), .C1(n20762), .C2(keyinput89), .A(n20636), .ZN(n20641) );
  AOI22_X1 U23569 ( .A1(n20639), .A2(keyinput123), .B1(keyinput88), .B2(n20811), .ZN(n20638) );
  OAI221_X1 U23570 ( .B1(n20639), .B2(keyinput123), .C1(n20811), .C2(
        keyinput88), .A(n20638), .ZN(n20640) );
  NOR4_X1 U23571 ( .A1(n20643), .A2(n20642), .A3(n20641), .A4(n20640), .ZN(
        n20682) );
  AOI22_X1 U23572 ( .A1(n14341), .A2(keyinput83), .B1(keyinput114), .B2(n20791), .ZN(n20644) );
  OAI221_X1 U23573 ( .B1(n14341), .B2(keyinput83), .C1(n20791), .C2(
        keyinput114), .A(n20644), .ZN(n20654) );
  AOI22_X1 U23574 ( .A1(n20646), .A2(keyinput68), .B1(n11072), .B2(keyinput93), 
        .ZN(n20645) );
  OAI221_X1 U23575 ( .B1(n20646), .B2(keyinput68), .C1(n11072), .C2(keyinput93), .A(n20645), .ZN(n20653) );
  AOI22_X1 U23576 ( .A1(n20648), .A2(keyinput74), .B1(n20756), .B2(keyinput122), .ZN(n20647) );
  OAI221_X1 U23577 ( .B1(n20648), .B2(keyinput74), .C1(n20756), .C2(
        keyinput122), .A(n20647), .ZN(n20652) );
  AOI22_X1 U23578 ( .A1(n20809), .A2(keyinput73), .B1(keyinput95), .B2(n20650), 
        .ZN(n20649) );
  OAI221_X1 U23579 ( .B1(n20809), .B2(keyinput73), .C1(n20650), .C2(keyinput95), .A(n20649), .ZN(n20651) );
  NOR4_X1 U23580 ( .A1(n20654), .A2(n20653), .A3(n20652), .A4(n20651), .ZN(
        n20681) );
  INV_X1 U23581 ( .A(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n20656) );
  AOI22_X1 U23582 ( .A1(n20656), .A2(keyinput86), .B1(keyinput100), .B2(n20792), .ZN(n20655) );
  OAI221_X1 U23583 ( .B1(n20656), .B2(keyinput86), .C1(n20792), .C2(
        keyinput100), .A(n20655), .ZN(n20667) );
  AOI22_X1 U23584 ( .A1(n20788), .A2(keyinput101), .B1(n11961), .B2(keyinput65), .ZN(n20657) );
  OAI221_X1 U23585 ( .B1(n20788), .B2(keyinput101), .C1(n11961), .C2(
        keyinput65), .A(n20657), .ZN(n20666) );
  AOI22_X1 U23586 ( .A1(n20660), .A2(keyinput71), .B1(keyinput118), .B2(n20659), .ZN(n20658) );
  OAI221_X1 U23587 ( .B1(n20660), .B2(keyinput71), .C1(n20659), .C2(
        keyinput118), .A(n20658), .ZN(n20665) );
  XOR2_X1 U23588 ( .A(n20661), .B(keyinput72), .Z(n20663) );
  XNOR2_X1 U23589 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B(keyinput98), .ZN(
        n20662) );
  NAND2_X1 U23590 ( .A1(n20663), .A2(n20662), .ZN(n20664) );
  NOR4_X1 U23591 ( .A1(n20667), .A2(n20666), .A3(n20665), .A4(n20664), .ZN(
        n20680) );
  AOI22_X1 U23592 ( .A1(n10395), .A2(keyinput70), .B1(keyinput77), .B2(n20775), 
        .ZN(n20668) );
  OAI221_X1 U23593 ( .B1(n10395), .B2(keyinput70), .C1(n20775), .C2(keyinput77), .A(n20668), .ZN(n20678) );
  AOI22_X1 U23594 ( .A1(n20776), .A2(keyinput126), .B1(keyinput109), .B2(
        n20670), .ZN(n20669) );
  OAI221_X1 U23595 ( .B1(n20776), .B2(keyinput126), .C1(n20670), .C2(
        keyinput109), .A(n20669), .ZN(n20677) );
  INV_X1 U23596 ( .A(DATAI_3_), .ZN(n20672) );
  AOI22_X1 U23597 ( .A1(n20672), .A2(keyinput90), .B1(n10885), .B2(keyinput87), 
        .ZN(n20671) );
  OAI221_X1 U23598 ( .B1(n20672), .B2(keyinput90), .C1(n10885), .C2(keyinput87), .A(n20671), .ZN(n20676) );
  XNOR2_X1 U23599 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(keyinput94), 
        .ZN(n20674) );
  XNOR2_X1 U23600 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B(keyinput112), 
        .ZN(n20673) );
  NAND2_X1 U23601 ( .A1(n20674), .A2(n20673), .ZN(n20675) );
  NOR4_X1 U23602 ( .A1(n20678), .A2(n20677), .A3(n20676), .A4(n20675), .ZN(
        n20679) );
  NAND4_X1 U23603 ( .A1(n20682), .A2(n20681), .A3(n20680), .A4(n20679), .ZN(
        n20824) );
  AOI22_X1 U23604 ( .A1(HOLD), .A2(keyinput121), .B1(
        P3_INSTQUEUE_REG_6__5__SCAN_IN), .B2(keyinput96), .ZN(n20683) );
  OAI221_X1 U23605 ( .B1(HOLD), .B2(keyinput121), .C1(
        P3_INSTQUEUE_REG_6__5__SCAN_IN), .C2(keyinput96), .A(n20683), .ZN(
        n20690) );
  AOI22_X1 U23606 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(keyinput80), 
        .B1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B2(keyinput82), .ZN(n20684) );
  OAI221_X1 U23607 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(keyinput80), 
        .C1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .C2(keyinput82), .A(n20684), .ZN(
        n20689) );
  AOI22_X1 U23608 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(keyinput105), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(keyinput110), .ZN(n20685) );
  OAI221_X1 U23609 ( .B1(P1_DATAO_REG_19__SCAN_IN), .B2(keyinput105), .C1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(keyinput110), .A(n20685), .ZN(
        n20688) );
  AOI22_X1 U23610 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(keyinput113), .B1(
        P2_INSTQUEUE_REG_15__4__SCAN_IN), .B2(keyinput81), .ZN(n20686) );
  OAI221_X1 U23611 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(keyinput113), .C1(
        P2_INSTQUEUE_REG_15__4__SCAN_IN), .C2(keyinput81), .A(n20686), .ZN(
        n20687) );
  NOR4_X1 U23612 ( .A1(n20690), .A2(n20689), .A3(n20688), .A4(n20687), .ZN(
        n20718) );
  AOI22_X1 U23613 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(keyinput84), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(keyinput67), .ZN(n20691) );
  OAI221_X1 U23614 ( .B1(P3_REIP_REG_30__SCAN_IN), .B2(keyinput84), .C1(
        P2_REIP_REG_27__SCAN_IN), .C2(keyinput67), .A(n20691), .ZN(n20698) );
  AOI22_X1 U23615 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(keyinput119), .B1(
        P2_INSTQUEUE_REG_12__4__SCAN_IN), .B2(keyinput91), .ZN(n20692) );
  OAI221_X1 U23616 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(keyinput119), .C1(
        P2_INSTQUEUE_REG_12__4__SCAN_IN), .C2(keyinput91), .A(n20692), .ZN(
        n20697) );
  AOI22_X1 U23617 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(keyinput104), .B1(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(keyinput103), .ZN(n20693) );
  OAI221_X1 U23618 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(keyinput104), .C1(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(keyinput103), .A(n20693), 
        .ZN(n20696) );
  AOI22_X1 U23619 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(keyinput69), 
        .B1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B2(keyinput111), .ZN(n20694) );
  OAI221_X1 U23620 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput69), 
        .C1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .C2(keyinput111), .A(n20694), 
        .ZN(n20695) );
  NOR4_X1 U23621 ( .A1(n20698), .A2(n20697), .A3(n20696), .A4(n20695), .ZN(
        n20717) );
  AOI22_X1 U23622 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(keyinput92), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(keyinput64), .ZN(n20699) );
  OAI221_X1 U23623 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(keyinput92), .C1(
        P2_REIP_REG_4__SCAN_IN), .C2(keyinput64), .A(n20699), .ZN(n20706) );
  AOI22_X1 U23624 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(keyinput66), .B1(
        P1_INSTQUEUE_REG_12__1__SCAN_IN), .B2(keyinput116), .ZN(n20700) );
  OAI221_X1 U23625 ( .B1(P2_DATAO_REG_3__SCAN_IN), .B2(keyinput66), .C1(
        P1_INSTQUEUE_REG_12__1__SCAN_IN), .C2(keyinput116), .A(n20700), .ZN(
        n20705) );
  AOI22_X1 U23626 ( .A1(keyinput120), .A2(BUF1_REG_26__SCAN_IN), .B1(n20812), 
        .B2(keyinput125), .ZN(n20701) );
  OAI221_X1 U23627 ( .B1(keyinput120), .B2(BUF1_REG_26__SCAN_IN), .C1(n20812), 
        .C2(keyinput125), .A(n20701), .ZN(n20704) );
  AOI22_X1 U23628 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(keyinput115), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(keyinput107), .ZN(n20702) );
  OAI221_X1 U23629 ( .B1(P3_EAX_REG_22__SCAN_IN), .B2(keyinput115), .C1(
        P2_BE_N_REG_0__SCAN_IN), .C2(keyinput107), .A(n20702), .ZN(n20703) );
  NOR4_X1 U23630 ( .A1(n20706), .A2(n20705), .A3(n20704), .A4(n20703), .ZN(
        n20716) );
  AOI22_X1 U23631 ( .A1(BUF2_REG_21__SCAN_IN), .A2(keyinput78), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(keyinput75), .ZN(n20707) );
  OAI221_X1 U23632 ( .B1(BUF2_REG_21__SCAN_IN), .B2(keyinput78), .C1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .C2(keyinput75), .A(n20707), .ZN(
        n20714) );
  AOI22_X1 U23633 ( .A1(P3_LWORD_REG_13__SCAN_IN), .A2(keyinput76), .B1(
        P3_EBX_REG_28__SCAN_IN), .B2(keyinput108), .ZN(n20708) );
  OAI221_X1 U23634 ( .B1(P3_LWORD_REG_13__SCAN_IN), .B2(keyinput76), .C1(
        P3_EBX_REG_28__SCAN_IN), .C2(keyinput108), .A(n20708), .ZN(n20713) );
  AOI22_X1 U23635 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(keyinput79), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(keyinput85), .ZN(n20709) );
  OAI221_X1 U23636 ( .B1(P1_UWORD_REG_10__SCAN_IN), .B2(keyinput79), .C1(
        P1_REIP_REG_12__SCAN_IN), .C2(keyinput85), .A(n20709), .ZN(n20712) );
  AOI22_X1 U23637 ( .A1(P3_LWORD_REG_10__SCAN_IN), .A2(keyinput97), .B1(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(keyinput102), .ZN(n20710) );
  OAI221_X1 U23638 ( .B1(P3_LWORD_REG_10__SCAN_IN), .B2(keyinput97), .C1(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(keyinput102), .A(n20710), 
        .ZN(n20711) );
  NOR4_X1 U23639 ( .A1(n20714), .A2(n20713), .A3(n20712), .A4(n20711), .ZN(
        n20715) );
  NAND4_X1 U23640 ( .A1(n20718), .A2(n20717), .A3(n20716), .A4(n20715), .ZN(
        n20823) );
  OAI22_X1 U23641 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(keyinput30), 
        .B1(keyinput44), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n20719) );
  AOI221_X1 U23642 ( .B1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(keyinput30), 
        .C1(P3_EBX_REG_28__SCAN_IN), .C2(keyinput44), .A(n20719), .ZN(n20726)
         );
  OAI22_X1 U23643 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(keyinput2), .B1(
        keyinput51), .B2(P3_EAX_REG_22__SCAN_IN), .ZN(n20720) );
  AOI221_X1 U23644 ( .B1(P2_DATAO_REG_3__SCAN_IN), .B2(keyinput2), .C1(
        P3_EAX_REG_22__SCAN_IN), .C2(keyinput51), .A(n20720), .ZN(n20725) );
  OAI22_X1 U23645 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(keyinput60), 
        .B1(P1_UWORD_REG_10__SCAN_IN), .B2(keyinput15), .ZN(n20721) );
  AOI221_X1 U23646 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(keyinput60), 
        .C1(keyinput15), .C2(P1_UWORD_REG_10__SCAN_IN), .A(n20721), .ZN(n20724) );
  OAI22_X1 U23647 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(keyinput29), .B1(
        keyinput52), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n20722) );
  AOI221_X1 U23648 ( .B1(P2_REIP_REG_5__SCAN_IN), .B2(keyinput29), .C1(
        P1_INSTQUEUE_REG_12__1__SCAN_IN), .C2(keyinput52), .A(n20722), .ZN(
        n20723) );
  NAND4_X1 U23649 ( .A1(n20726), .A2(n20725), .A3(n20724), .A4(n20723), .ZN(
        n20754) );
  OAI22_X1 U23650 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(keyinput40), .B1(
        P2_EBX_REG_27__SCAN_IN), .B2(keyinput7), .ZN(n20727) );
  AOI221_X1 U23651 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(keyinput40), .C1(
        keyinput7), .C2(P2_EBX_REG_27__SCAN_IN), .A(n20727), .ZN(n20734) );
  OAI22_X1 U23652 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(keyinput17), 
        .B1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B2(keyinput22), .ZN(n20728) );
  AOI221_X1 U23653 ( .B1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B2(keyinput17), 
        .C1(keyinput22), .C2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A(n20728), 
        .ZN(n20733) );
  OAI22_X1 U23654 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(keyinput34), .B1(
        keyinput42), .B2(P1_LWORD_REG_9__SCAN_IN), .ZN(n20729) );
  AOI221_X1 U23655 ( .B1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(keyinput34), 
        .C1(P1_LWORD_REG_9__SCAN_IN), .C2(keyinput42), .A(n20729), .ZN(n20732)
         );
  OAI22_X1 U23656 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(keyinput59), 
        .B1(P1_DATAO_REG_25__SCAN_IN), .B2(keyinput54), .ZN(n20730) );
  AOI221_X1 U23657 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(keyinput59), 
        .C1(keyinput54), .C2(P1_DATAO_REG_25__SCAN_IN), .A(n20730), .ZN(n20731) );
  NAND4_X1 U23658 ( .A1(n20734), .A2(n20733), .A3(n20732), .A4(n20731), .ZN(
        n20753) );
  OAI22_X1 U23659 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(keyinput49), .B1(
        P1_DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput10), .ZN(n20735) );
  AOI221_X1 U23660 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(keyinput49), .C1(
        keyinput10), .C2(P1_DATAWIDTH_REG_20__SCAN_IN), .A(n20735), .ZN(n20742) );
  OAI22_X1 U23661 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(keyinput31), 
        .B1(keyinput4), .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n20736) );
  AOI221_X1 U23662 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput31), 
        .C1(P2_DATAO_REG_11__SCAN_IN), .C2(keyinput4), .A(n20736), .ZN(n20741)
         );
  OAI22_X1 U23663 ( .A1(BUF1_REG_26__SCAN_IN), .A2(keyinput56), .B1(DATAI_3_), 
        .B2(keyinput26), .ZN(n20737) );
  AOI221_X1 U23664 ( .B1(BUF1_REG_26__SCAN_IN), .B2(keyinput56), .C1(
        keyinput26), .C2(DATAI_3_), .A(n20737), .ZN(n20740) );
  OAI22_X1 U23665 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(keyinput21), .B1(
        keyinput45), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n20738) );
  AOI221_X1 U23666 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(keyinput21), .C1(
        P3_INSTQUEUE_REG_1__5__SCAN_IN), .C2(keyinput45), .A(n20738), .ZN(
        n20739) );
  NAND4_X1 U23667 ( .A1(n20742), .A2(n20741), .A3(n20740), .A4(n20739), .ZN(
        n20752) );
  OAI22_X1 U23668 ( .A1(P2_EAX_REG_4__SCAN_IN), .A2(keyinput23), .B1(keyinput8), .B2(P1_EBX_REG_5__SCAN_IN), .ZN(n20743) );
  AOI221_X1 U23669 ( .B1(P2_EAX_REG_4__SCAN_IN), .B2(keyinput23), .C1(
        P1_EBX_REG_5__SCAN_IN), .C2(keyinput8), .A(n20743), .ZN(n20750) );
  OAI22_X1 U23670 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(keyinput6), .B1(
        P1_INSTQUEUE_REG_5__2__SCAN_IN), .B2(keyinput35), .ZN(n20744) );
  AOI221_X1 U23671 ( .B1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B2(keyinput6), .C1(
        keyinput35), .C2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A(n20744), .ZN(
        n20749) );
  OAI22_X1 U23672 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(keyinput55), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(keyinput53), .ZN(n20745) );
  AOI221_X1 U23673 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(keyinput55), .C1(
        keyinput53), .C2(P1_DATAO_REG_31__SCAN_IN), .A(n20745), .ZN(n20748) );
  OAI22_X1 U23674 ( .A1(n13674), .A2(keyinput14), .B1(keyinput19), .B2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n20746) );
  AOI221_X1 U23675 ( .B1(n13674), .B2(keyinput14), .C1(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(keyinput19), .A(n20746), .ZN(
        n20747) );
  NAND4_X1 U23676 ( .A1(n20750), .A2(n20749), .A3(n20748), .A4(n20747), .ZN(
        n20751) );
  NOR4_X1 U23677 ( .A1(n20754), .A2(n20753), .A3(n20752), .A4(n20751), .ZN(
        n20822) );
  AOI22_X1 U23678 ( .A1(n20757), .A2(keyinput12), .B1(n20756), .B2(keyinput58), 
        .ZN(n20755) );
  OAI221_X1 U23679 ( .B1(n20757), .B2(keyinput12), .C1(n20756), .C2(keyinput58), .A(n20755), .ZN(n20770) );
  AOI22_X1 U23680 ( .A1(n20760), .A2(keyinput18), .B1(keyinput38), .B2(n20759), 
        .ZN(n20758) );
  OAI221_X1 U23681 ( .B1(n20760), .B2(keyinput18), .C1(n20759), .C2(keyinput38), .A(n20758), .ZN(n20769) );
  AOI22_X1 U23682 ( .A1(n20763), .A2(keyinput3), .B1(keyinput25), .B2(n20762), 
        .ZN(n20761) );
  OAI221_X1 U23683 ( .B1(n20763), .B2(keyinput3), .C1(n20762), .C2(keyinput25), 
        .A(n20761), .ZN(n20768) );
  INV_X1 U23684 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n20764) );
  XOR2_X1 U23685 ( .A(keyinput5), .B(n20764), .Z(n20766) );
  XNOR2_X1 U23686 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B(keyinput27), .ZN(
        n20765) );
  NAND2_X1 U23687 ( .A1(n20766), .A2(n20765), .ZN(n20767) );
  NOR4_X1 U23688 ( .A1(n20770), .A2(n20769), .A3(n20768), .A4(n20767), .ZN(
        n20820) );
  INV_X1 U23689 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n20773) );
  INV_X1 U23690 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n20772) );
  AOI22_X1 U23691 ( .A1(n20773), .A2(keyinput47), .B1(keyinput32), .B2(n20772), 
        .ZN(n20771) );
  OAI221_X1 U23692 ( .B1(n20773), .B2(keyinput47), .C1(n20772), .C2(keyinput32), .A(n20771), .ZN(n20786) );
  AOI22_X1 U23693 ( .A1(n20776), .A2(keyinput62), .B1(keyinput13), .B2(n20775), 
        .ZN(n20774) );
  OAI221_X1 U23694 ( .B1(n20776), .B2(keyinput62), .C1(n20775), .C2(keyinput13), .A(n20774), .ZN(n20785) );
  INV_X1 U23695 ( .A(P3_LWORD_REG_10__SCAN_IN), .ZN(n20779) );
  AOI22_X1 U23696 ( .A1(n20779), .A2(keyinput33), .B1(n20778), .B2(keyinput11), 
        .ZN(n20777) );
  OAI221_X1 U23697 ( .B1(n20779), .B2(keyinput33), .C1(n20778), .C2(keyinput11), .A(n20777), .ZN(n20784) );
  AOI22_X1 U23698 ( .A1(n20782), .A2(keyinput57), .B1(n20781), .B2(keyinput63), 
        .ZN(n20780) );
  OAI221_X1 U23699 ( .B1(n20782), .B2(keyinput57), .C1(n20781), .C2(keyinput63), .A(n20780), .ZN(n20783) );
  NOR4_X1 U23700 ( .A1(n20786), .A2(n20785), .A3(n20784), .A4(n20783), .ZN(
        n20819) );
  AOI22_X1 U23701 ( .A1(n20789), .A2(keyinput41), .B1(n20788), .B2(keyinput37), 
        .ZN(n20787) );
  OAI221_X1 U23702 ( .B1(n20789), .B2(keyinput41), .C1(n20788), .C2(keyinput37), .A(n20787), .ZN(n20801) );
  AOI22_X1 U23703 ( .A1(n20792), .A2(keyinput36), .B1(n20791), .B2(keyinput50), 
        .ZN(n20790) );
  OAI221_X1 U23704 ( .B1(n20792), .B2(keyinput36), .C1(n20791), .C2(keyinput50), .A(n20790), .ZN(n20800) );
  INV_X1 U23705 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20795) );
  AOI22_X1 U23706 ( .A1(n20795), .A2(keyinput48), .B1(keyinput46), .B2(n20794), 
        .ZN(n20793) );
  OAI221_X1 U23707 ( .B1(n20795), .B2(keyinput48), .C1(n20794), .C2(keyinput46), .A(n20793), .ZN(n20799) );
  AOI22_X1 U23708 ( .A1(n20797), .A2(keyinput28), .B1(n11066), .B2(keyinput0), 
        .ZN(n20796) );
  OAI221_X1 U23709 ( .B1(n20797), .B2(keyinput28), .C1(n11066), .C2(keyinput0), 
        .A(n20796), .ZN(n20798) );
  NOR4_X1 U23710 ( .A1(n20801), .A2(n20800), .A3(n20799), .A4(n20798), .ZN(
        n20818) );
  AOI22_X1 U23711 ( .A1(n20804), .A2(keyinput20), .B1(n20803), .B2(keyinput16), 
        .ZN(n20802) );
  OAI221_X1 U23712 ( .B1(n20804), .B2(keyinput20), .C1(n20803), .C2(keyinput16), .A(n20802), .ZN(n20816) );
  AOI22_X1 U23713 ( .A1(n20806), .A2(keyinput43), .B1(n11961), .B2(keyinput1), 
        .ZN(n20805) );
  OAI221_X1 U23714 ( .B1(n20806), .B2(keyinput43), .C1(n11961), .C2(keyinput1), 
        .A(n20805), .ZN(n20815) );
  AOI22_X1 U23715 ( .A1(n20809), .A2(keyinput9), .B1(keyinput39), .B2(n20808), 
        .ZN(n20807) );
  OAI221_X1 U23716 ( .B1(n20809), .B2(keyinput9), .C1(n20808), .C2(keyinput39), 
        .A(n20807), .ZN(n20814) );
  AOI22_X1 U23717 ( .A1(n20812), .A2(keyinput61), .B1(n20811), .B2(keyinput24), 
        .ZN(n20810) );
  OAI221_X1 U23718 ( .B1(n20812), .B2(keyinput61), .C1(n20811), .C2(keyinput24), .A(n20810), .ZN(n20813) );
  NOR4_X1 U23719 ( .A1(n20816), .A2(n20815), .A3(n20814), .A4(n20813), .ZN(
        n20817) );
  AND4_X1 U23720 ( .A1(n20820), .A2(n20819), .A3(n20818), .A4(n20817), .ZN(
        n20821) );
  OAI211_X1 U23721 ( .C1(n20824), .C2(n20823), .A(n20822), .B(n20821), .ZN(
        n20837) );
  AOI22_X1 U23722 ( .A1(n20828), .A2(n20827), .B1(n20826), .B2(n20825), .ZN(
        n20833) );
  AOI22_X1 U23723 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20831), .B1(
        n20830), .B2(n20829), .ZN(n20832) );
  OAI211_X1 U23724 ( .C1(n20835), .C2(n20834), .A(n20833), .B(n20832), .ZN(
        n20836) );
  XNOR2_X1 U23725 ( .A(n20837), .B(n20836), .ZN(P2_U3069) );
  OR2_X1 U14581 ( .A1(n11649), .A2(n11648), .ZN(n19868) );
  INV_X1 U11072 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18583) );
  BUF_X2 U12336 ( .A(n15264), .Z(n13753) );
  AND2_X1 U11331 ( .A1(n10247), .A2(n10527), .ZN(n11584) );
  CLKBUF_X3 U11174 ( .A(n9676), .Z(n9615) );
  CLKBUF_X1 U11070 ( .A(n11699), .Z(n12378) );
  CLKBUF_X1 U11083 ( .A(n11668), .Z(n12254) );
  CLKBUF_X2 U11092 ( .A(n10182), .Z(n10369) );
  INV_X1 U11094 ( .A(n9782), .ZN(n10783) );
  NOR2_X1 U11106 ( .A1(n17993), .A2(n17997), .ZN(n15151) );
  CLKBUF_X1 U11113 ( .A(n13064), .Z(n12466) );
  AND2_X1 U11149 ( .A1(n10130), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14986) );
  CLKBUF_X1 U11156 ( .A(n9767), .Z(n9622) );
  NAND2_X1 U11161 ( .A1(n10364), .A2(n9954), .ZN(n19397) );
  CLKBUF_X1 U11184 ( .A(n15102), .Z(n15224) );
  CLKBUF_X3 U11192 ( .A(n13732), .Z(n16909) );
  CLKBUF_X1 U11196 ( .A(n13770), .Z(n16936) );
  NAND2_X1 U11361 ( .A1(n13689), .A2(n18591), .ZN(n16689) );
  AND4_X1 U11457 ( .A1(n11727), .A2(n11726), .A3(n11725), .A4(n11724), .ZN(
        n11728) );
  CLKBUF_X1 U11480 ( .A(n13224), .Z(n9635) );
  CLKBUF_X1 U12322 ( .A(n16293), .Z(n16291) );
  OR2_X1 U12650 ( .A1(n15288), .A2(n15287), .ZN(n20838) );
  INV_X2 U12879 ( .A(n11181), .ZN(n18933) );
endmodule

