

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput63,
         keyinput62, keyinput61, keyinput60, keyinput59, keyinput58,
         keyinput57, keyinput56, keyinput55, keyinput54, keyinput53,
         keyinput52, keyinput51, keyinput50, keyinput49, keyinput48,
         keyinput47, keyinput46, keyinput45, keyinput44, keyinput43,
         keyinput42, keyinput41, keyinput40, keyinput39, keyinput38,
         keyinput37, keyinput36, keyinput35, keyinput34, keyinput33,
         keyinput32, keyinput31, keyinput30, keyinput29, keyinput28,
         keyinput27, keyinput26, keyinput25, keyinput24, keyinput23,
         keyinput22, keyinput21, keyinput20, keyinput19, keyinput18,
         keyinput17, keyinput16, keyinput15, keyinput14, keyinput13,
         keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7,
         keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1,
         keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6439, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250;

  AND2_X1 U7187 ( .A1(n13887), .A2(n13886), .ZN(n14011) );
  XNOR2_X1 U7188 ( .A(n14361), .B(n7217), .ZN(n14402) );
  XNOR2_X1 U7189 ( .A(n14351), .B(n7212), .ZN(n14395) );
  INV_X1 U7190 ( .A(n6859), .ZN(n14351) );
  NAND2_X1 U7191 ( .A1(n10455), .A2(n10454), .ZN(n10453) );
  NOR2_X1 U7192 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14346), .ZN(n14290) );
  INV_X1 U7193 ( .A(n13262), .ZN(n8927) );
  INV_X1 U7194 ( .A(n6452), .ZN(n11217) );
  NAND2_X1 U7195 ( .A1(n12326), .A2(n12331), .ZN(n9979) );
  AND4_X1 U7196 ( .A1(n9868), .A2(n9867), .A3(n9866), .A4(n9865), .ZN(n11410)
         );
  INV_X2 U7197 ( .A(n8904), .ZN(n8207) );
  BUF_X4 U7198 ( .A(n9733), .Z(n11599) );
  NAND2_X1 U7199 ( .A1(n6698), .A2(n6610), .ZN(n8664) );
  NAND2_X1 U7200 ( .A1(n8183), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8185) );
  INV_X1 U7201 ( .A(n7687), .ZN(n7949) );
  NAND2_X1 U7203 ( .A1(n7679), .A2(n6589), .ZN(n13146) );
  AND3_X1 U7204 ( .A1(n7663), .A2(n7664), .A3(n7666), .ZN(n6588) );
  INV_X1 U7205 ( .A(n14860), .ZN(n11880) );
  INV_X1 U7206 ( .A(n11881), .ZN(n6617) );
  INV_X1 U7207 ( .A(n7508), .ZN(n8101) );
  AND2_X1 U7209 ( .A1(n13315), .A2(n7102), .ZN(n7101) );
  AND2_X1 U7210 ( .A1(n7097), .A2(n7103), .ZN(n7096) );
  OR2_X1 U7211 ( .A1(n8584), .A2(n11270), .ZN(n7035) );
  OR2_X1 U7212 ( .A1(n13313), .A2(n8147), .ZN(n13294) );
  NAND2_X1 U7213 ( .A1(n7662), .A2(n9679), .ZN(n7687) );
  INV_X1 U7214 ( .A(n7662), .ZN(n7948) );
  CLKBUF_X2 U7215 ( .A(n10361), .Z(n11801) );
  INV_X1 U7216 ( .A(n11399), .ZN(n7375) );
  INV_X2 U7217 ( .A(n8245), .ZN(n10393) );
  OR2_X1 U7218 ( .A1(n14957), .A2(n14956), .ZN(n14954) );
  AND2_X1 U7219 ( .A1(n12509), .A2(n12508), .ZN(n12510) );
  INV_X1 U7220 ( .A(n7644), .ZN(n7650) );
  BUF_X1 U7221 ( .A(n12043), .Z(n6442) );
  INV_X1 U7222 ( .A(n8927), .ZN(n13465) );
  INV_X1 U7223 ( .A(n11655), .ZN(n11502) );
  INV_X1 U7225 ( .A(n11545), .ZN(n11501) );
  XOR2_X1 U7226 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n14328), .Z(n14365) );
  NOR2_X2 U7227 ( .A1(n8666), .A2(n14892), .ZN(n12330) );
  CLKBUF_X2 U7228 ( .A(n12045), .Z(n6614) );
  AND2_X1 U7229 ( .A1(n7119), .A2(n6654), .ZN(n13420) );
  NAND2_X1 U7230 ( .A1(n7859), .A2(n7858), .ZN(n13645) );
  OR2_X1 U7231 ( .A1(n7640), .A2(n7869), .ZN(n7642) );
  NAND2_X1 U7232 ( .A1(n9197), .A2(n9163), .ZN(n9202) );
  INV_X1 U7233 ( .A(n8188), .ZN(n11738) );
  NAND2_X1 U7234 ( .A1(n9587), .A2(n7293), .ZN(n11375) );
  AND2_X1 U7235 ( .A1(n14039), .A2(n13901), .ZN(n6439) );
  NOR2_X2 U7236 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7463) );
  NOR2_X4 U7237 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9197) );
  OR2_X2 U7238 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14303), .ZN(n14326) );
  NAND2_X2 U7239 ( .A1(n9804), .A2(n7441), .ZN(n9805) );
  AOI21_X2 U7240 ( .B1(n8675), .B2(n6468), .A(n6449), .ZN(n10770) );
  NOR2_X2 U7241 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7462) );
  OAI21_X2 U7242 ( .B1(n9893), .B2(n6491), .A(n6596), .ZN(n7177) );
  NOR2_X2 U7243 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7461) );
  NAND2_X2 U7244 ( .A1(n11391), .A2(n11383), .ZN(n11675) );
  AOI21_X2 U7245 ( .B1(n10548), .B2(n10549), .A(n6531), .ZN(n10669) );
  OR2_X1 U7246 ( .A1(n11654), .A2(n9858), .ZN(n9861) );
  XNOR2_X2 U7247 ( .A(n8185), .B(n8184), .ZN(n8187) );
  NAND2_X2 U7248 ( .A1(n11857), .A2(n11856), .ZN(n13675) );
  XNOR2_X1 U7250 ( .A(n8231), .B(n8789), .ZN(n12305) );
  NAND2_X2 U7252 ( .A1(n14249), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9615) );
  XNOR2_X2 U7253 ( .A(n7800), .B(n7799), .ZN(n10739) );
  NAND2_X2 U7254 ( .A1(n6972), .A2(n7555), .ZN(n7800) );
  XNOR2_X2 U7255 ( .A(n14353), .B(n13148), .ZN(n15244) );
  NAND2_X2 U7256 ( .A1(n7211), .A2(n14352), .ZN(n14353) );
  XNOR2_X2 U7257 ( .A(n8016), .B(n8015), .ZN(n14273) );
  OAI21_X2 U7258 ( .B1(n8292), .B2(n8291), .A(n8293), .ZN(n8307) );
  NAND2_X2 U7259 ( .A1(n8279), .A2(n8278), .ZN(n8292) );
  NAND2_X2 U7260 ( .A1(n8611), .A2(n8610), .ZN(n8625) );
  NAND2_X2 U7261 ( .A1(n7174), .A2(n13882), .ZN(n14072) );
  XNOR2_X2 U7262 ( .A(n14357), .B(n14358), .ZN(n14401) );
  NAND2_X2 U7263 ( .A1(n14355), .A2(n14356), .ZN(n14357) );
  NAND2_X2 U7264 ( .A1(n13652), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7639) );
  AND2_X2 U7267 ( .A1(n12106), .A2(n8119), .ZN(n7109) );
  XNOR2_X2 U7268 ( .A(n13492), .B(n13139), .ZN(n12106) );
  XNOR2_X2 U7269 ( .A(n7214), .B(P1_ADDR_REG_1__SCAN_IN), .ZN(n14335) );
  INV_X4 U7270 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n7214) );
  XNOR2_X2 U7271 ( .A(n14364), .B(n7215), .ZN(n14403) );
  NAND2_X2 U7272 ( .A1(n7216), .A2(n14363), .ZN(n14364) );
  AND2_X1 U7273 ( .A1(n6481), .A2(n6818), .ZN(n9106) );
  NOR2_X1 U7274 ( .A1(n12642), .A2(n8711), .ZN(n8765) );
  OR2_X1 U7275 ( .A1(n9082), .A2(n9081), .ZN(n11734) );
  AOI21_X1 U7276 ( .B1(n12797), .B2(n7041), .A(n7039), .ZN(n7038) );
  NAND2_X1 U7277 ( .A1(n11180), .A2(n11690), .ZN(n11291) );
  AND2_X1 U7278 ( .A1(n10336), .A2(n10334), .ZN(n7376) );
  CLKBUF_X2 U7279 ( .A(P2_U3947), .Z(n6445) );
  NAND2_X2 U7280 ( .A1(n13811), .A2(n10171), .ZN(n11396) );
  INV_X1 U7281 ( .A(n13808), .ZN(n10478) );
  INV_X1 U7282 ( .A(n14744), .ZN(n10926) );
  INV_X1 U7283 ( .A(n13143), .ZN(n10586) );
  INV_X1 U7284 ( .A(n15068), .ZN(n10027) );
  INV_X1 U7285 ( .A(n12499), .ZN(n8231) );
  CLKBUF_X2 U7286 ( .A(n10135), .Z(n6635) );
  INV_X1 U7287 ( .A(n10042), .ZN(n8783) );
  AND4_X1 U7288 ( .A1(n9623), .A2(n9622), .A3(n9621), .A4(n9620), .ZN(n9731)
         );
  NAND4_X1 U7289 ( .A1(n8242), .A2(n8241), .A3(n8240), .A4(n8239), .ZN(n12498)
         );
  AND3_X1 U7290 ( .A1(n7657), .A2(n7656), .A3(n7655), .ZN(n6613) );
  BUF_X2 U7291 ( .A(n9899), .Z(n11614) );
  OR2_X1 U7292 ( .A1(n12045), .A2(n10274), .ZN(n7664) );
  OR2_X1 U7293 ( .A1(n12045), .A2(n9527), .ZN(n7656) );
  CLKBUF_X2 U7294 ( .A(n7687), .Z(n12061) );
  CLKBUF_X2 U7295 ( .A(n10112), .Z(n11646) );
  INV_X4 U7296 ( .A(n11422), .ZN(n6443) );
  BUF_X2 U7297 ( .A(n8267), .Z(n6448) );
  CLKBUF_X2 U7298 ( .A(n8267), .Z(n6447) );
  NAND2_X2 U7299 ( .A1(n7662), .A2(n11542), .ZN(n8033) );
  XNOR2_X1 U7300 ( .A(n7630), .B(n7629), .ZN(n8158) );
  INV_X1 U7301 ( .A(n8187), .ZN(n8189) );
  NAND2_X1 U7302 ( .A1(n7521), .A2(n7520), .ZN(n7524) );
  INV_X1 U7303 ( .A(n7529), .ZN(n7530) );
  AND2_X1 U7304 ( .A1(n14136), .A2(n14135), .ZN(n6629) );
  NOR2_X1 U7305 ( .A1(n13943), .A2(n6644), .ZN(n14146) );
  NAND2_X1 U7306 ( .A1(n13891), .A2(n7365), .ZN(n13942) );
  NOR2_X1 U7307 ( .A1(n6649), .A2(n6648), .ZN(n13507) );
  AND2_X1 U7308 ( .A1(n6763), .A2(n6762), .ZN(n11717) );
  NAND2_X1 U7309 ( .A1(n7349), .A2(n7352), .ZN(n7348) );
  CLKBUF_X1 U7310 ( .A(n14013), .Z(n6608) );
  NAND2_X1 U7311 ( .A1(n13234), .A2(n13233), .ZN(n13232) );
  NAND2_X1 U7312 ( .A1(n14011), .A2(n7351), .ZN(n14010) );
  NOR2_X1 U7313 ( .A1(n8698), .A2(n12661), .ZN(n6647) );
  AND2_X1 U7314 ( .A1(n11734), .A2(n9083), .ZN(n12990) );
  AOI21_X1 U7315 ( .B1(n7196), .B2(n13954), .A(n7195), .ZN(n7194) );
  INV_X1 U7316 ( .A(n13506), .ZN(n6648) );
  INV_X1 U7317 ( .A(n13893), .ZN(n7195) );
  NAND2_X1 U7318 ( .A1(n6609), .A2(n12735), .ZN(n12728) );
  OR2_X1 U7319 ( .A1(n12186), .A2(n6836), .ZN(n8845) );
  NAND2_X1 U7320 ( .A1(n13759), .A2(n13758), .ZN(n13757) );
  OAI21_X1 U7321 ( .B1(n7036), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n7035), .ZN(
        n8609) );
  NAND2_X1 U7322 ( .A1(n13068), .A2(n13069), .ZN(n13067) );
  NAND2_X1 U7323 ( .A1(n8574), .A2(n8573), .ZN(n12706) );
  NAND2_X1 U7324 ( .A1(n13047), .A2(n13048), .ZN(n13046) );
  NAND2_X1 U7325 ( .A1(n8035), .A2(n8034), .ZN(n13529) );
  NAND2_X1 U7326 ( .A1(n8003), .A2(n8002), .ZN(n13626) );
  NOR2_X1 U7327 ( .A1(n13804), .A2(n11181), .ZN(n11286) );
  NAND2_X1 U7328 ( .A1(n11934), .A2(n11933), .ZN(n11937) );
  NAND2_X1 U7329 ( .A1(n6626), .A2(n7604), .ZN(n8014) );
  NAND2_X1 U7330 ( .A1(n8406), .A2(n12392), .ZN(n12836) );
  NAND2_X1 U7331 ( .A1(n10970), .A2(n8124), .ZN(n11159) );
  NAND2_X1 U7332 ( .A1(n14367), .A2(n14366), .ZN(n14596) );
  CLKBUF_X1 U7333 ( .A(n14538), .Z(n6612) );
  NAND2_X1 U7334 ( .A1(n7589), .A2(n7406), .ZN(n7947) );
  NOR2_X1 U7335 ( .A1(n10713), .A2(n8335), .ZN(n10986) );
  XNOR2_X1 U7336 ( .A(n7150), .B(n10727), .ZN(n10713) );
  NAND2_X1 U7337 ( .A1(n7037), .A2(n12359), .ZN(n10903) );
  OR2_X1 U7338 ( .A1(n7586), .A2(n9751), .ZN(n7589) );
  NAND2_X1 U7339 ( .A1(n6793), .A2(n7151), .ZN(n10712) );
  NAND2_X1 U7340 ( .A1(n7804), .A2(n7803), .ZN(n13479) );
  OAI22_X1 U7341 ( .A1(n10333), .A2(n10332), .B1(n10331), .B2(n14727), .ZN(
        n14678) );
  NAND2_X1 U7342 ( .A1(n10111), .A2(n10110), .ZN(n10333) );
  NAND2_X2 U7343 ( .A1(n10313), .A2(n10312), .ZN(n11435) );
  NAND2_X1 U7344 ( .A1(n7773), .A2(n7772), .ZN(n11923) );
  NOR2_X1 U7345 ( .A1(n9069), .A2(n9065), .ZN(n13116) );
  OR2_X1 U7346 ( .A1(n8394), .A2(n8393), .ZN(n8408) );
  OAI21_X1 U7347 ( .B1(n7766), .B2(n6729), .A(n6727), .ZN(n7830) );
  INV_X2 U7348 ( .A(n14775), .ZN(n6444) );
  AND2_X1 U7349 ( .A1(n12359), .A2(n12349), .ZN(n12346) );
  NAND2_X1 U7350 ( .A1(n7737), .A2(n6965), .ZN(n6962) );
  NAND2_X1 U7351 ( .A1(n7544), .A2(n7543), .ZN(n7737) );
  NAND2_X1 U7352 ( .A1(n8781), .A2(n8780), .ZN(n8788) );
  INV_X1 U7353 ( .A(n11410), .ZN(n6446) );
  INV_X1 U7354 ( .A(n9731), .ZN(n9693) );
  NAND4_X1 U7355 ( .A1(n7709), .A2(n7708), .A3(n7707), .A4(n7706), .ZN(n13144)
         );
  INV_X1 U7356 ( .A(n11867), .ZN(n10361) );
  OAI21_X1 U7357 ( .B1(n8513), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n6840) );
  OAI211_X1 U7358 ( .C1(n7662), .C2(n9525), .A(n7689), .B(n7688), .ZN(n11890)
         );
  NAND2_X1 U7359 ( .A1(n6791), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9932) );
  OR2_X1 U7360 ( .A1(n8033), .A2(n9680), .ZN(n7675) );
  INV_X1 U7361 ( .A(n9685), .ZN(n9677) );
  INV_X2 U7362 ( .A(n11654), .ZN(n11641) );
  CLKBUF_X1 U7363 ( .A(n8033), .Z(n6636) );
  AOI21_X1 U7364 ( .B1(n6965), .B2(n6967), .A(n6523), .ZN(n6963) );
  CLKBUF_X3 U7365 ( .A(n7678), .Z(n12049) );
  CLKBUF_X3 U7366 ( .A(n9859), .Z(n11655) );
  INV_X4 U7367 ( .A(n9773), .ZN(n12602) );
  CLKBUF_X1 U7368 ( .A(n10393), .Z(n9092) );
  CLKBUF_X1 U7369 ( .A(n12085), .Z(n6595) );
  NAND2_X1 U7370 ( .A1(n9272), .A2(n9189), .ZN(n9685) );
  INV_X1 U7371 ( .A(n9618), .ZN(n14258) );
  XNOR2_X1 U7372 ( .A(n9177), .B(P1_IR_REG_25__SCAN_IN), .ZN(n9272) );
  CLKBUF_X1 U7373 ( .A(n8158), .Z(n9481) );
  CLKBUF_X1 U7374 ( .A(n9306), .Z(n14262) );
  XNOR2_X1 U7375 ( .A(n9617), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9618) );
  NAND2_X1 U7376 ( .A1(n9181), .A2(n9180), .ZN(n9273) );
  NAND2_X1 U7377 ( .A1(n9180), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9177) );
  XNOR2_X1 U7378 ( .A(n7492), .B(n7491), .ZN(n7508) );
  MUX2_X1 U7379 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9179), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9181) );
  NAND2_X1 U7380 ( .A1(n9176), .A2(n9183), .ZN(n9180) );
  OR2_X1 U7381 ( .A1(n12984), .A2(n12985), .ZN(n8182) );
  XNOR2_X1 U7382 ( .A(n7524), .B(n9256), .ZN(n7668) );
  INV_X2 U7383 ( .A(n14272), .ZN(n14270) );
  NAND2_X2 U7384 ( .A1(n9679), .A2(P2_U3088), .ZN(n13671) );
  XNOR2_X1 U7385 ( .A(n9253), .B(n9252), .ZN(n9307) );
  NAND2_X1 U7386 ( .A1(n7490), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7492) );
  OAI21_X1 U7387 ( .B1(n9588), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9586) );
  AOI22_X1 U7388 ( .A1(n7935), .A2(n7501), .B1(n7500), .B2(n7499), .ZN(n7502)
         );
  OR2_X1 U7389 ( .A1(n9251), .A2(n9235), .ZN(n9253) );
  OR2_X1 U7390 ( .A1(n14282), .A2(n7210), .ZN(n6864) );
  XNOR2_X1 U7391 ( .A(n9247), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14279) );
  AND2_X1 U7392 ( .A1(n6464), .A2(n8184), .ZN(n6936) );
  INV_X4 U7393 ( .A(n7530), .ZN(n11542) );
  INV_X2 U7394 ( .A(n7530), .ZN(n11363) );
  NOR2_X1 U7395 ( .A1(n6830), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n6828) );
  INV_X1 U7396 ( .A(n7173), .ZN(n9761) );
  NAND2_X1 U7397 ( .A1(n7460), .A2(n7459), .ZN(n7698) );
  AND4_X1 U7398 ( .A1(n6715), .A2(n6714), .A3(n8443), .A4(n6843), .ZN(n8178)
         );
  NAND4_X1 U7399 ( .A1(n9216), .A2(n9160), .A3(n9161), .A4(n9159), .ZN(n9162)
         );
  AND3_X1 U7400 ( .A1(n7259), .A2(n7258), .A3(n7257), .ZN(n9164) );
  AND3_X1 U7401 ( .A1(n8176), .A2(n8174), .A3(n8175), .ZN(n8396) );
  AND2_X1 U7402 ( .A1(n8172), .A2(n8179), .ZN(n7431) );
  INV_X1 U7403 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7259) );
  INV_X1 U7404 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7683) );
  INV_X1 U7405 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8180) );
  INV_X4 U7406 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7407 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n9245) );
  INV_X1 U7408 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9216) );
  INV_X1 U7409 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8172) );
  INV_X1 U7410 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9160) );
  INV_X1 U7411 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9161) );
  INV_X1 U7412 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9159) );
  INV_X1 U7413 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8443) );
  INV_X1 U7414 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7491) );
  NOR2_X1 U7415 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n8175) );
  NOR2_X1 U7416 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8174) );
  NOR2_X1 U7417 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n8176) );
  INV_X1 U7418 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n7258) );
  INV_X1 U7419 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7257) );
  NOR2_X1 U7420 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n6715) );
  NOR2_X1 U7421 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n6714) );
  NOR2_X1 U7422 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8171) );
  OR2_X1 U7423 ( .A1(n10285), .A2(n11890), .ZN(n10286) );
  OAI22_X2 U7424 ( .A1(n14349), .A2(n14294), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14293), .ZN(n14295) );
  OAI21_X2 U7425 ( .B1(n11732), .B2(n13603), .A(n6587), .ZN(n8771) );
  AND2_X1 U7426 ( .A1(n11729), .A2(n11726), .ZN(n6587) );
  AND2_X1 U7427 ( .A1(n7644), .A2(n11324), .ZN(n12043) );
  NAND2_X2 U7428 ( .A1(n9609), .A2(n11375), .ZN(n9684) );
  OAI21_X2 U7429 ( .B1(n7947), .B2(n7946), .A(n7592), .ZN(n7593) );
  NAND2_X2 U7430 ( .A1(n11738), .A2(n8187), .ZN(n8238) );
  XNOR2_X2 U7431 ( .A(n10478), .B(n11435), .ZN(n11682) );
  NAND2_X1 U7432 ( .A1(n11738), .A2(n8189), .ZN(n8267) );
  AND2_X1 U7433 ( .A1(n9140), .A2(n9112), .ZN(n9114) );
  OR2_X1 U7434 ( .A1(n12150), .A2(n10227), .ZN(n12456) );
  INV_X1 U7435 ( .A(n7023), .ZN(n7022) );
  NAND2_X1 U7436 ( .A1(n12119), .A2(n8146), .ZN(n7102) );
  INV_X1 U7437 ( .A(n6490), .ZN(n6830) );
  AOI21_X1 U7438 ( .B1(n7352), .B2(n7351), .A(n6515), .ZN(n7350) );
  NAND2_X1 U7439 ( .A1(n6987), .A2(n6986), .ZN(n6984) );
  NOR2_X1 U7440 ( .A1(n7394), .A2(n6971), .ZN(n6970) );
  INV_X1 U7441 ( .A(n7555), .ZN(n6971) );
  AND2_X1 U7442 ( .A1(n6478), .A2(n7302), .ZN(n7301) );
  INV_X1 U7443 ( .A(n7305), .ZN(n7302) );
  AND2_X1 U7444 ( .A1(n6974), .A2(n6973), .ZN(n7232) );
  INV_X1 U7445 ( .A(n12052), .ZN(n6974) );
  AND2_X1 U7446 ( .A1(n12058), .A2(n12081), .ZN(n6973) );
  NOR2_X1 U7447 ( .A1(n13447), .A2(n7123), .ZN(n7122) );
  INV_X1 U7448 ( .A(n7883), .ZN(n7123) );
  NAND2_X1 U7449 ( .A1(n12241), .A2(n8846), .ZN(n8850) );
  OAI21_X1 U7450 ( .B1(n12223), .B2(n8840), .A(n8844), .ZN(n6835) );
  NAND2_X1 U7451 ( .A1(n10514), .A2(n7145), .ZN(n6787) );
  INV_X1 U7452 ( .A(n10199), .ZN(n7146) );
  NAND2_X1 U7453 ( .A1(n6624), .A2(n6623), .ZN(n6903) );
  INV_X1 U7454 ( .A(n14986), .ZN(n6623) );
  NAND2_X1 U7455 ( .A1(n12550), .A2(n12551), .ZN(n12552) );
  NOR2_X1 U7456 ( .A1(n12573), .A2(n6892), .ZN(n12590) );
  NOR2_X1 U7457 ( .A1(n12555), .A2(n12554), .ZN(n6892) );
  NAND2_X1 U7458 ( .A1(n7059), .A2(n12449), .ZN(n7058) );
  INV_X1 U7459 ( .A(n12450), .ZN(n7059) );
  OR2_X1 U7460 ( .A1(n12747), .A2(n12733), .ZN(n12322) );
  INV_X1 U7461 ( .A(n8686), .ZN(n6709) );
  AND2_X1 U7462 ( .A1(n8687), .A2(n6707), .ZN(n6706) );
  NAND2_X1 U7463 ( .A1(n6708), .A2(n8686), .ZN(n6707) );
  INV_X1 U7464 ( .A(n8685), .ZN(n6708) );
  OR2_X1 U7465 ( .A1(n12976), .A2(n12842), .ZN(n12407) );
  OR2_X1 U7466 ( .A1(n11335), .A2(n14477), .ZN(n6697) );
  NOR2_X1 U7467 ( .A1(n7438), .A2(n8212), .ZN(n8214) );
  OR2_X1 U7468 ( .A1(n8258), .A2(n9256), .ZN(n8213) );
  XNOR2_X1 U7469 ( .A(n8198), .B(n8199), .ZN(n8663) );
  NAND2_X1 U7470 ( .A1(n8722), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8198) );
  INV_X1 U7471 ( .A(n9049), .ZN(n6677) );
  INV_X1 U7472 ( .A(n8928), .ZN(n9052) );
  NOR2_X1 U7473 ( .A1(n13512), .A2(n13514), .ZN(n6923) );
  NAND2_X1 U7474 ( .A1(n13323), .A2(n8012), .ZN(n7090) );
  AND2_X1 U7475 ( .A1(n8149), .A2(n8041), .ZN(n12121) );
  AND2_X1 U7476 ( .A1(n7133), .A2(n6535), .ZN(n7131) );
  NOR2_X1 U7477 ( .A1(n13589), .A2(n6927), .ZN(n6926) );
  INV_X1 U7478 ( .A(n6928), .ZN(n6927) );
  NOR2_X1 U7479 ( .A1(n7828), .A2(n7117), .ZN(n7116) );
  INV_X1 U7480 ( .A(n7813), .ZN(n7117) );
  XNOR2_X1 U7481 ( .A(n13104), .B(n13142), .ZN(n12102) );
  NAND2_X1 U7482 ( .A1(n8101), .A2(n12091), .ZN(n12085) );
  NAND2_X1 U7483 ( .A1(n8057), .A2(n8056), .ZN(n13270) );
  OR2_X1 U7484 ( .A1(n13284), .A2(n8055), .ZN(n8057) );
  NOR2_X1 U7485 ( .A1(n7884), .A2(n7126), .ZN(n7125) );
  INV_X1 U7486 ( .A(n7128), .ZN(n7126) );
  AND2_X1 U7487 ( .A1(n7475), .A2(n6477), .ZN(n7627) );
  NAND2_X1 U7488 ( .A1(n7833), .A2(n7464), .ZN(n7071) );
  NOR3_X1 U7489 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .A3(
        P2_IR_REG_4__SCAN_IN), .ZN(n7464) );
  NOR2_X1 U7490 ( .A1(n7488), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n7509) );
  INV_X1 U7491 ( .A(n10167), .ZN(n7266) );
  INV_X1 U7492 ( .A(n9799), .ZN(n11863) );
  NAND2_X1 U7493 ( .A1(n7364), .A2(n7368), .ZN(n6724) );
  NAND2_X1 U7494 ( .A1(n14132), .A2(n14120), .ZN(n7368) );
  NAND2_X1 U7495 ( .A1(n7367), .A2(n7365), .ZN(n7364) );
  NOR2_X1 U7496 ( .A1(n13997), .A2(n7189), .ZN(n7188) );
  INV_X1 U7497 ( .A(n13889), .ZN(n7189) );
  OR2_X1 U7498 ( .A1(n14214), .A2(n14202), .ZN(n13897) );
  INV_X1 U7499 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9183) );
  INV_X1 U7500 ( .A(n10257), .ZN(n9172) );
  AND2_X1 U7501 ( .A1(n7402), .A2(n7579), .ZN(n7401) );
  OR2_X1 U7502 ( .A1(n6487), .A2(n7403), .ZN(n7402) );
  NAND2_X1 U7503 ( .A1(n7832), .A2(n7567), .ZN(n7854) );
  AOI21_X1 U7504 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n14300), .A(n14299), .ZN(
        n14359) );
  OR2_X1 U7505 ( .A1(n8519), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8532) );
  NAND2_X1 U7506 ( .A1(n9139), .A2(n9113), .ZN(n9123) );
  INV_X1 U7507 ( .A(n12668), .ZN(n8887) );
  NAND2_X1 U7508 ( .A1(n8852), .A2(n12705), .ZN(n9137) );
  OR2_X1 U7509 ( .A1(n12201), .A2(n12204), .ZN(n12202) );
  NAND2_X1 U7510 ( .A1(n9934), .A2(n6792), .ZN(n14908) );
  OR2_X1 U7511 ( .A1(n7140), .A2(n14906), .ZN(n6792) );
  NAND2_X1 U7512 ( .A1(n7140), .A2(n14906), .ZN(n9934) );
  NOR2_X1 U7513 ( .A1(n14939), .A2(n8296), .ZN(n14938) );
  OR2_X1 U7514 ( .A1(n10995), .A2(n10996), .ZN(n6889) );
  NAND2_X1 U7515 ( .A1(n10712), .A2(n10711), .ZN(n7150) );
  NAND2_X1 U7516 ( .A1(n6889), .A2(n6888), .ZN(n14958) );
  INV_X1 U7517 ( .A(n14960), .ZN(n6888) );
  AND2_X1 U7518 ( .A1(n6899), .A2(n6898), .ZN(n12516) );
  INV_X1 U7519 ( .A(n11072), .ZN(n6898) );
  NAND2_X1 U7520 ( .A1(n6878), .A2(n6877), .ZN(n12502) );
  INV_X1 U7521 ( .A(n11069), .ZN(n6877) );
  XNOR2_X1 U7522 ( .A(n12504), .B(n14980), .ZN(n14982) );
  NAND2_X1 U7523 ( .A1(n12502), .A2(n12501), .ZN(n12504) );
  OR2_X1 U7524 ( .A1(n14982), .A2(n14983), .ZN(n6883) );
  NAND2_X1 U7525 ( .A1(n7158), .A2(n7157), .ZN(n12550) );
  INV_X1 U7526 ( .A(n12520), .ZN(n7157) );
  NAND2_X1 U7527 ( .A1(n7031), .A2(n6637), .ZN(n9088) );
  AND2_X1 U7528 ( .A1(n7029), .A2(n6507), .ZN(n6637) );
  INV_X1 U7529 ( .A(n8901), .ZN(n7030) );
  AND2_X1 U7530 ( .A1(n12456), .A2(n9078), .ZN(n12461) );
  NAND2_X1 U7531 ( .A1(n7031), .A2(n6507), .ZN(n8706) );
  NAND2_X1 U7532 ( .A1(n6831), .A2(n12423), .ZN(n12746) );
  NAND2_X1 U7533 ( .A1(n7038), .A2(n12424), .ZN(n6831) );
  NAND2_X1 U7534 ( .A1(n6954), .A2(n6953), .ZN(n8682) );
  AND2_X1 U7535 ( .A1(n7449), .A2(n8680), .ZN(n6953) );
  AOI21_X1 U7536 ( .B1(n7048), .B2(n7050), .A(n7047), .ZN(n7046) );
  INV_X1 U7537 ( .A(n12381), .ZN(n7047) );
  INV_X1 U7538 ( .A(n7053), .ZN(n7048) );
  INV_X1 U7539 ( .A(n8352), .ZN(n8351) );
  NAND2_X2 U7540 ( .A1(n9753), .A2(n9679), .ZN(n12281) );
  INV_X1 U7541 ( .A(n12860), .ZN(n12844) );
  NAND2_X1 U7542 ( .A1(n8614), .A2(n8613), .ZN(n9148) );
  OR2_X1 U7543 ( .A1(n8258), .A2(n11320), .ZN(n8613) );
  OR2_X1 U7544 ( .A1(n11321), .A2(n12281), .ZN(n8614) );
  INV_X1 U7545 ( .A(n12281), .ZN(n12277) );
  INV_X1 U7546 ( .A(n8258), .ZN(n8516) );
  INV_X1 U7547 ( .A(n9753), .ZN(n8515) );
  INV_X1 U7548 ( .A(n12862), .ZN(n12841) );
  NAND2_X1 U7549 ( .A1(n8724), .A2(n8740), .ZN(n9285) );
  OR2_X1 U7550 ( .A1(n6700), .A2(n6699), .ZN(n6611) );
  NAND2_X1 U7551 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), 
        .ZN(n6699) );
  INV_X1 U7552 ( .A(n8663), .ZN(n9773) );
  INV_X1 U7553 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n6712) );
  INV_X1 U7554 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n6711) );
  AOI21_X1 U7555 ( .B1(n7344), .B2(n6685), .A(n6684), .ZN(n6683) );
  INV_X1 U7556 ( .A(n10383), .ZN(n6685) );
  INV_X1 U7557 ( .A(n8965), .ZN(n6684) );
  AND2_X1 U7558 ( .A1(n6673), .A2(n6671), .ZN(n6667) );
  INV_X1 U7559 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7465) );
  NAND2_X1 U7560 ( .A1(n13270), .A2(n12123), .ZN(n8071) );
  AND2_X1 U7561 ( .A1(n13294), .A2(n8148), .ZN(n13315) );
  INV_X1 U7562 ( .A(n7083), .ZN(n7082) );
  NAND2_X1 U7563 ( .A1(n8125), .A2(n7139), .ZN(n7138) );
  OR2_X1 U7564 ( .A1(n7478), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n7480) );
  NAND2_X1 U7565 ( .A1(n10923), .A2(n7286), .ZN(n7285) );
  INV_X1 U7566 ( .A(n10920), .ZN(n7286) );
  NOR2_X1 U7567 ( .A1(n14523), .A2(n7277), .ZN(n7276) );
  INV_X1 U7568 ( .A(n11742), .ZN(n7277) );
  INV_X1 U7569 ( .A(n6724), .ZN(n7363) );
  NAND2_X1 U7570 ( .A1(n13970), .A2(n13890), .ZN(n13944) );
  NOR2_X1 U7571 ( .A1(n7347), .A2(n13979), .ZN(n7346) );
  INV_X1 U7572 ( .A(n7350), .ZN(n7347) );
  BUF_X1 U7573 ( .A(n9856), .Z(n11654) );
  AND2_X1 U7574 ( .A1(n7372), .A2(n11691), .ZN(n7369) );
  NAND2_X1 U7575 ( .A1(n10480), .A2(n11685), .ZN(n10762) );
  NAND2_X1 U7576 ( .A1(n11545), .A2(n9679), .ZN(n9856) );
  NAND2_X1 U7577 ( .A1(n11545), .A2(n11542), .ZN(n9859) );
  NAND2_X1 U7578 ( .A1(n11360), .A2(n11359), .ZN(n11653) );
  NAND2_X1 U7579 ( .A1(n11357), .A2(n11356), .ZN(n11360) );
  NAND2_X1 U7580 ( .A1(n7634), .A2(SI_27_), .ZN(n8077) );
  NAND2_X1 U7581 ( .A1(n7613), .A2(n7612), .ZN(n8032) );
  INV_X1 U7582 ( .A(n8029), .ZN(n7612) );
  NAND2_X1 U7583 ( .A1(n7589), .A2(n7587), .ZN(n7932) );
  INV_X1 U7584 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6863) );
  INV_X1 U7585 ( .A(n6876), .ZN(n14361) );
  OAI21_X1 U7586 ( .B1(n14401), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6497), .ZN(
        n6876) );
  NOR2_X1 U7587 ( .A1(n9101), .A2(n9100), .ZN(n9102) );
  XNOR2_X1 U7588 ( .A(n8099), .B(n8155), .ZN(n11732) );
  NAND2_X1 U7589 ( .A1(n7201), .A2(n7202), .ZN(n7206) );
  INV_X1 U7590 ( .A(n14376), .ZN(n7202) );
  NAND2_X1 U7591 ( .A1(n11881), .A2(n11880), .ZN(n6584) );
  INV_X1 U7592 ( .A(n11919), .ZN(n7251) );
  INV_X1 U7593 ( .A(n11925), .ZN(n7246) );
  AND2_X1 U7594 ( .A1(n12094), .A2(n7248), .ZN(n7247) );
  NAND2_X1 U7595 ( .A1(n11919), .A2(n7249), .ZN(n7248) );
  NAND2_X1 U7596 ( .A1(n11418), .A2(n11421), .ZN(n6986) );
  INV_X1 U7597 ( .A(n6986), .ZN(n6757) );
  NAND2_X1 U7598 ( .A1(n11416), .A2(n11415), .ZN(n11419) );
  AND2_X1 U7599 ( .A1(n6988), .A2(n11420), .ZN(n6987) );
  INV_X1 U7600 ( .A(n11418), .ZN(n6988) );
  INV_X1 U7601 ( .A(n11436), .ZN(n7001) );
  NOR2_X1 U7602 ( .A1(n11439), .A2(n11436), .ZN(n7002) );
  NAND2_X1 U7603 ( .A1(n6993), .A2(n11449), .ZN(n6992) );
  NOR2_X1 U7604 ( .A1(n11449), .A2(n6993), .ZN(n6994) );
  NAND2_X1 U7605 ( .A1(n11980), .A2(n11982), .ZN(n7236) );
  NAND2_X1 U7606 ( .A1(n6760), .A2(n6758), .ZN(n11461) );
  NAND2_X1 U7607 ( .A1(n11457), .A2(n6759), .ZN(n6758) );
  AOI21_X1 U7608 ( .B1(n6983), .B2(n11689), .A(n6982), .ZN(n6981) );
  INV_X1 U7609 ( .A(n11473), .ZN(n6982) );
  NAND2_X1 U7610 ( .A1(n13882), .A2(n11499), .ZN(n6772) );
  NOR2_X1 U7611 ( .A1(n13881), .A2(n11499), .ZN(n6773) );
  NAND2_X1 U7612 ( .A1(n11991), .A2(n11993), .ZN(n7239) );
  INV_X1 U7613 ( .A(n11999), .ZN(n7220) );
  NAND2_X1 U7614 ( .A1(n12009), .A2(n12011), .ZN(n7233) );
  OAI22_X1 U7615 ( .A1(n11587), .A2(n11585), .B1(n11573), .B2(n7000), .ZN(
        n6999) );
  INV_X1 U7616 ( .A(n11572), .ZN(n7000) );
  INV_X1 U7617 ( .A(n8110), .ZN(n7080) );
  NAND2_X1 U7618 ( .A1(n8630), .A2(n7024), .ZN(n12455) );
  NOR2_X1 U7619 ( .A1(n7026), .A2(n7025), .ZN(n7024) );
  INV_X1 U7620 ( .A(n8629), .ZN(n7025) );
  NOR2_X1 U7621 ( .A1(n13022), .A2(n7314), .ZN(n7313) );
  INV_X1 U7622 ( .A(n9021), .ZN(n7314) );
  NOR2_X1 U7623 ( .A1(n7925), .A2(n7924), .ZN(n7923) );
  AOI21_X1 U7624 ( .B1(n6749), .B2(n6748), .A(n6747), .ZN(n6746) );
  INV_X1 U7625 ( .A(n7599), .ZN(n6747) );
  INV_X1 U7626 ( .A(n6975), .ZN(n6748) );
  NAND2_X1 U7627 ( .A1(n7572), .A2(n9348), .ZN(n7579) );
  INV_X1 U7628 ( .A(n7577), .ZN(n7403) );
  NOR2_X1 U7629 ( .A1(n6969), .A2(n6731), .ZN(n6730) );
  INV_X1 U7630 ( .A(n7552), .ZN(n6731) );
  INV_X1 U7631 ( .A(n7393), .ZN(n7392) );
  OAI21_X1 U7632 ( .B1(n7394), .B2(n7556), .A(n7563), .ZN(n7393) );
  NAND2_X1 U7633 ( .A1(n6970), .A2(n7782), .ZN(n6968) );
  NAND2_X1 U7634 ( .A1(n6730), .A2(n7765), .ZN(n6728) );
  NAND2_X1 U7635 ( .A1(n7560), .A2(n7559), .ZN(n7563) );
  INV_X1 U7636 ( .A(SI_11_), .ZN(n7559) );
  INV_X1 U7637 ( .A(n7209), .ZN(n14285) );
  OAI21_X1 U7638 ( .B1(n14342), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6529), .ZN(
        n7209) );
  INV_X1 U7639 ( .A(n6864), .ZN(n14284) );
  NAND2_X1 U7640 ( .A1(n11228), .A2(n8811), .ZN(n8813) );
  OR2_X1 U7641 ( .A1(n9110), .A2(n9132), .ZN(n9140) );
  INV_X1 U7642 ( .A(n12329), .ZN(n12323) );
  AOI21_X1 U7643 ( .B1(n8816), .B2(n6856), .A(n6579), .ZN(n6854) );
  AOI21_X1 U7644 ( .B1(n6851), .B2(n6850), .A(n6849), .ZN(n6848) );
  INV_X1 U7645 ( .A(n6853), .ZN(n6850) );
  INV_X1 U7646 ( .A(n12158), .ZN(n6849) );
  NAND2_X1 U7647 ( .A1(n9930), .A2(n7141), .ZN(n7140) );
  OR2_X1 U7648 ( .A1(n9931), .A2(n10308), .ZN(n7141) );
  AND2_X1 U7649 ( .A1(n10536), .A2(n10535), .ZN(n10538) );
  AND2_X1 U7650 ( .A1(n10999), .A2(n11076), .ZN(n7162) );
  NAND2_X1 U7651 ( .A1(n12541), .A2(n12540), .ZN(n12542) );
  AOI21_X1 U7652 ( .B1(n12586), .B2(n12585), .A(n12584), .ZN(n12607) );
  INV_X1 U7653 ( .A(n12458), .ZN(n6827) );
  NAND2_X1 U7654 ( .A1(n7056), .A2(n6824), .ZN(n6823) );
  INV_X1 U7655 ( .A(n6825), .ZN(n6824) );
  NAND2_X1 U7656 ( .A1(n8616), .A2(n8615), .ZN(n8631) );
  OR2_X1 U7657 ( .A1(n12182), .A2(n12745), .ZN(n12433) );
  INV_X1 U7658 ( .A(n12397), .ZN(n6807) );
  INV_X1 U7659 ( .A(n12407), .ZN(n6805) );
  AOI21_X1 U7660 ( .B1(n7046), .B2(n7049), .A(n7045), .ZN(n7044) );
  INV_X1 U7661 ( .A(n12382), .ZN(n7045) );
  INV_X1 U7662 ( .A(n7046), .ZN(n6813) );
  NOR2_X1 U7663 ( .A1(n8366), .A2(n7051), .ZN(n7050) );
  INV_X1 U7664 ( .A(n12376), .ZN(n7051) );
  INV_X1 U7665 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n10723) );
  NAND2_X1 U7666 ( .A1(n12342), .A2(n12345), .ZN(n6716) );
  NAND2_X1 U7667 ( .A1(n10245), .A2(n10042), .ZN(n12326) );
  NAND2_X1 U7668 ( .A1(n12484), .A2(n12323), .ZN(n12457) );
  NOR2_X1 U7669 ( .A1(n7435), .A2(P3_IR_REG_26__SCAN_IN), .ZN(n7434) );
  NAND2_X1 U7670 ( .A1(n8181), .A2(n7436), .ZN(n7435) );
  INV_X1 U7671 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7436) );
  INV_X1 U7672 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8181) );
  INV_X1 U7673 ( .A(n7020), .ZN(n7019) );
  OAI21_X1 U7674 ( .B1(n8454), .B2(n7021), .A(n8471), .ZN(n7020) );
  INV_X1 U7675 ( .A(n8456), .ZN(n7021) );
  NAND2_X1 U7676 ( .A1(n8408), .A2(n8407), .ZN(n8409) );
  INV_X1 U7677 ( .A(n7013), .ZN(n7012) );
  OAI21_X1 U7678 ( .B1(n8326), .B2(n7014), .A(n8345), .ZN(n7013) );
  INV_X1 U7679 ( .A(n8328), .ZN(n7014) );
  NOR2_X1 U7680 ( .A1(n8398), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8319) );
  INV_X1 U7681 ( .A(n9054), .ZN(n6671) );
  NOR2_X1 U7682 ( .A1(n6489), .A2(n7323), .ZN(n7320) );
  NAND2_X1 U7683 ( .A1(n8989), .A2(n8990), .ZN(n7316) );
  INV_X1 U7684 ( .A(n11245), .ZN(n7317) );
  NAND2_X1 U7685 ( .A1(n6478), .A2(n7307), .ZN(n7303) );
  INV_X1 U7686 ( .A(n7313), .ZN(n7306) );
  INV_X1 U7687 ( .A(n9026), .ZN(n7310) );
  NOR2_X1 U7688 ( .A1(n9027), .A2(n7310), .ZN(n7308) );
  INV_X1 U7689 ( .A(n7229), .ZN(n7226) );
  NAND2_X1 U7690 ( .A1(n6532), .A2(n7232), .ZN(n7227) );
  OAI21_X1 U7691 ( .B1(n12074), .B2(n7231), .A(n7230), .ZN(n7229) );
  NAND2_X1 U7692 ( .A1(n7232), .A2(n7225), .ZN(n7224) );
  INV_X1 U7693 ( .A(n12035), .ZN(n7225) );
  AND2_X1 U7694 ( .A1(n7232), .A2(n12028), .ZN(n7228) );
  NAND2_X1 U7695 ( .A1(n7644), .A2(n7645), .ZN(n7678) );
  INV_X1 U7696 ( .A(n11324), .ZN(n7645) );
  NOR2_X1 U7697 ( .A1(n13626), .A2(n6917), .ZN(n6915) );
  NOR2_X1 U7698 ( .A1(n12107), .A2(n7115), .ZN(n7111) );
  INV_X1 U7699 ( .A(n7827), .ZN(n7115) );
  INV_X1 U7700 ( .A(n7116), .ZN(n7114) );
  INV_X1 U7701 ( .A(n7101), .ZN(n7099) );
  AND2_X1 U7702 ( .A1(n12121), .A2(n13294), .ZN(n7103) );
  INV_X1 U7703 ( .A(n8146), .ZN(n7098) );
  INV_X1 U7704 ( .A(n7065), .ZN(n7064) );
  NAND2_X1 U7705 ( .A1(n8117), .A2(n8116), .ZN(n10506) );
  NOR2_X1 U7706 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n7345) );
  AND3_X1 U7707 ( .A1(n7468), .A2(n7467), .A3(n7466), .ZN(n7474) );
  INV_X1 U7708 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n7510) );
  NAND2_X1 U7709 ( .A1(n11369), .A2(n11370), .ZN(n11663) );
  NAND2_X1 U7710 ( .A1(n11622), .A2(n11625), .ZN(n6995) );
  NOR2_X1 U7711 ( .A1(n11625), .A2(n11622), .ZN(n6996) );
  XNOR2_X1 U7712 ( .A(n14118), .B(n13912), .ZN(n11697) );
  INV_X1 U7713 ( .A(n13885), .ZN(n7182) );
  OAI21_X1 U7714 ( .B1(n7183), .B2(n7182), .A(n13902), .ZN(n7181) );
  AND2_X1 U7715 ( .A1(n13884), .A2(n13883), .ZN(n7183) );
  AND2_X1 U7716 ( .A1(n6459), .A2(n6952), .ZN(n6951) );
  OR2_X1 U7717 ( .A1(n11767), .A2(n14421), .ZN(n11468) );
  OR2_X1 U7718 ( .A1(n11703), .A2(n14279), .ZN(n11369) );
  NAND2_X1 U7719 ( .A1(n14279), .A2(n11703), .ZN(n11370) );
  NOR2_X1 U7720 ( .A1(n7618), .A2(SI_26_), .ZN(n6977) );
  INV_X1 U7721 ( .A(n7617), .ZN(n6740) );
  INV_X1 U7722 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9252) );
  INV_X1 U7723 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7374) );
  NAND2_X1 U7724 ( .A1(n7594), .A2(SI_20_), .ZN(n6975) );
  INV_X1 U7725 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7292) );
  NAND2_X1 U7726 ( .A1(n6735), .A2(n6734), .ZN(n7587) );
  NOR2_X1 U7727 ( .A1(n6736), .A2(SI_18_), .ZN(n6734) );
  OR2_X1 U7728 ( .A1(n9420), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9421) );
  INV_X1 U7729 ( .A(n7799), .ZN(n7556) );
  XNOR2_X1 U7730 ( .A(n7557), .B(SI_10_), .ZN(n7799) );
  NAND2_X1 U7731 ( .A1(n8806), .A2(n11114), .ZN(n8807) );
  NAND2_X1 U7732 ( .A1(n8231), .A2(n8791), .ZN(n8792) );
  INV_X1 U7733 ( .A(n8790), .ZN(n8791) );
  INV_X1 U7734 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10533) );
  AND2_X1 U7735 ( .A1(n12330), .A2(n12326), .ZN(n8785) );
  INV_X1 U7736 ( .A(n8788), .ZN(n12139) );
  INV_X1 U7737 ( .A(n8550), .ZN(n8549) );
  AOI21_X1 U7738 ( .B1(n6848), .B2(n6852), .A(n7416), .ZN(n6846) );
  INV_X1 U7739 ( .A(n6483), .ZN(n7417) );
  NAND2_X1 U7740 ( .A1(n12168), .A2(n12212), .ZN(n6832) );
  NAND2_X1 U7741 ( .A1(n8804), .A2(n8803), .ZN(n11098) );
  NOR2_X1 U7742 ( .A1(n6835), .A2(n12702), .ZN(n6834) );
  NAND2_X1 U7743 ( .A1(n6839), .A2(n6838), .ZN(n7448) );
  INV_X1 U7744 ( .A(n8812), .ZN(n6838) );
  INV_X1 U7745 ( .A(n8813), .ZN(n6839) );
  NAND2_X1 U7746 ( .A1(n8430), .A2(n12159), .ZN(n8447) );
  INV_X1 U7747 ( .A(n8431), .ZN(n8430) );
  AND2_X1 U7748 ( .A1(n12320), .A2(n12467), .ZN(n6592) );
  NOR2_X1 U7749 ( .A1(n12931), .A2(n12624), .ZN(n12470) );
  INV_X1 U7750 ( .A(n6448), .ZN(n8592) );
  INV_X1 U7751 ( .A(n14908), .ZN(n6791) );
  OR2_X1 U7752 ( .A1(n6493), .A2(n10205), .ZN(n14927) );
  NAND2_X1 U7753 ( .A1(n10528), .A2(n10529), .ZN(n14943) );
  XNOR2_X1 U7754 ( .A(n10538), .B(n7145), .ZN(n14937) );
  NAND2_X1 U7755 ( .A1(n6880), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7172) );
  INV_X1 U7756 ( .A(n14937), .ZN(n6880) );
  NAND2_X1 U7757 ( .A1(n6782), .A2(n6781), .ZN(n14939) );
  AOI21_X1 U7758 ( .B1(n7147), .B2(n6785), .A(n6783), .ZN(n6781) );
  INV_X1 U7759 ( .A(n6787), .ZN(n6784) );
  NAND2_X1 U7760 ( .A1(n10531), .A2(n10532), .ZN(n10719) );
  NAND2_X1 U7761 ( .A1(n7172), .A2(n7171), .ZN(n7170) );
  INV_X1 U7762 ( .A(n10539), .ZN(n7171) );
  AND2_X1 U7763 ( .A1(n7147), .A2(n7146), .ZN(n10516) );
  NAND2_X1 U7764 ( .A1(n12516), .A2(n12517), .ZN(n12518) );
  NAND2_X1 U7765 ( .A1(n7156), .A2(n7155), .ZN(n12509) );
  INV_X1 U7766 ( .A(n12506), .ZN(n7155) );
  INV_X1 U7767 ( .A(n6903), .ZN(n14984) );
  XNOR2_X1 U7768 ( .A(n12552), .B(n14457), .ZN(n14459) );
  INV_X1 U7769 ( .A(n12532), .ZN(n7148) );
  OR2_X1 U7770 ( .A1(n12574), .A2(n12575), .ZN(n7167) );
  OR2_X1 U7771 ( .A1(n12574), .A2(n6582), .ZN(n7165) );
  NAND2_X1 U7772 ( .A1(n12593), .A2(n7164), .ZN(n7163) );
  INV_X1 U7773 ( .A(n12595), .ZN(n7164) );
  OR2_X1 U7774 ( .A1(n9148), .A2(n8887), .ZN(n12450) );
  AND2_X1 U7775 ( .A1(n8699), .A2(n12679), .ZN(n12663) );
  NAND2_X1 U7776 ( .A1(n8596), .A2(n12440), .ZN(n12689) );
  OR2_X1 U7777 ( .A1(n12211), .A2(n12705), .ZN(n8596) );
  OR2_X1 U7778 ( .A1(n8575), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8590) );
  NAND2_X1 U7779 ( .A1(n8694), .A2(n8693), .ZN(n12730) );
  OAI21_X1 U7780 ( .B1(n12746), .B2(n12743), .A(n12322), .ZN(n12736) );
  NAND2_X1 U7781 ( .A1(n7040), .A2(n12415), .ZN(n7039) );
  NAND2_X1 U7782 ( .A1(n7041), .A2(n8687), .ZN(n7040) );
  AND2_X1 U7783 ( .A1(n8506), .A2(n7042), .ZN(n7041) );
  OAI21_X1 U7784 ( .B1(n6639), .B2(n6709), .A(n6706), .ZN(n8689) );
  AND2_X1 U7785 ( .A1(n6542), .A2(n6704), .ZN(n6703) );
  NAND2_X1 U7786 ( .A1(n6706), .A2(n6709), .ZN(n6704) );
  AND2_X1 U7787 ( .A1(n12415), .A2(n12418), .ZN(n12772) );
  OR2_X1 U7788 ( .A1(n8482), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8500) );
  NAND2_X1 U7790 ( .A1(n12854), .A2(n12855), .ZN(n8406) );
  INV_X1 U7791 ( .A(n6697), .ZN(n6694) );
  NAND2_X1 U7792 ( .A1(n6693), .A2(n6697), .ZN(n12840) );
  NAND2_X1 U7793 ( .A1(n8682), .A2(n6695), .ZN(n6693) );
  AND2_X1 U7794 ( .A1(n12392), .A2(n12391), .ZN(n12855) );
  INV_X1 U7795 ( .A(n12843), .ZN(n11335) );
  INV_X1 U7796 ( .A(n7050), .ZN(n7049) );
  NOR2_X1 U7797 ( .A1(n8349), .A2(n7054), .ZN(n7053) );
  NOR2_X1 U7798 ( .A1(n12369), .A2(n6934), .ZN(n6933) );
  INV_X1 U7799 ( .A(n8677), .ZN(n6934) );
  AOI21_X1 U7800 ( .B1(n6800), .B2(n6802), .A(n6798), .ZN(n6797) );
  INV_X1 U7801 ( .A(n12366), .ZN(n6798) );
  NAND2_X1 U7802 ( .A1(n8298), .A2(n8297), .ZN(n8333) );
  INV_X1 U7803 ( .A(n8299), .ZN(n8298) );
  OR2_X1 U7804 ( .A1(n8283), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8299) );
  NAND2_X1 U7805 ( .A1(n10300), .A2(n12305), .ZN(n6815) );
  NAND2_X1 U7806 ( .A1(n8882), .A2(n12460), .ZN(n12862) );
  NAND2_X1 U7807 ( .A1(n10247), .A2(n8669), .ZN(n10302) );
  OR2_X1 U7808 ( .A1(n12281), .A2(n9227), .ZN(n8229) );
  INV_X1 U7809 ( .A(n12612), .ZN(n8710) );
  INV_X1 U7810 ( .A(n9756), .ZN(n8868) );
  OAI211_X1 U7811 ( .C1(n8258), .C2(SI_12_), .A(n8404), .B(n8403), .ZN(n14477)
         );
  INV_X1 U7812 ( .A(n12457), .ZN(n12460) );
  NAND2_X1 U7813 ( .A1(n8651), .A2(n12329), .ZN(n15044) );
  INV_X1 U7814 ( .A(n9285), .ZN(n8736) );
  OAI21_X1 U7815 ( .B1(n9285), .B2(P3_D_REG_0__SCAN_IN), .A(n8727), .ZN(n8778)
         );
  OAI21_X1 U7816 ( .B1(n8625), .B2(n8624), .A(n8626), .ZN(n8895) );
  AND2_X1 U7817 ( .A1(n8723), .A2(n8722), .ZN(n8740) );
  INV_X1 U7818 ( .A(n6700), .ZN(n8720) );
  NAND2_X1 U7819 ( .A1(n8558), .A2(n8557), .ZN(n8571) );
  INV_X1 U7820 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8179) );
  XNOR2_X1 U7821 ( .A(n8644), .B(P3_IR_REG_20__SCAN_IN), .ZN(n8757) );
  OR2_X1 U7822 ( .A1(n8528), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8541) );
  NAND2_X1 U7823 ( .A1(n8511), .A2(n8510), .ZN(n8526) );
  NAND2_X1 U7824 ( .A1(n8476), .A2(n8475), .ZN(n8489) );
  AND2_X1 U7825 ( .A1(n8440), .A2(n8425), .ZN(n8438) );
  OR2_X1 U7826 ( .A1(n8409), .A2(n15111), .ZN(n7034) );
  NAND2_X1 U7827 ( .A1(n8409), .A2(n15111), .ZN(n8423) );
  XNOR2_X1 U7828 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8345) );
  XNOR2_X1 U7829 ( .A(n9263), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n8325) );
  CLKBUF_X1 U7830 ( .A(n8327), .Z(n6603) );
  OR2_X1 U7831 ( .A1(n8274), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8398) );
  NAND2_X1 U7832 ( .A1(n8173), .A2(n8172), .ZN(n8274) );
  NAND2_X1 U7833 ( .A1(n6795), .A2(n6794), .ZN(n7173) );
  INV_X1 U7834 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6795) );
  INV_X1 U7835 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6794) );
  AOI21_X1 U7836 ( .B1(n6675), .B2(n6674), .A(n6524), .ZN(n6673) );
  INV_X1 U7837 ( .A(n7342), .ZN(n6674) );
  NAND2_X1 U7838 ( .A1(n6673), .A2(n6670), .ZN(n6669) );
  NAND2_X1 U7839 ( .A1(n6676), .A2(n6671), .ZN(n6670) );
  AND2_X1 U7840 ( .A1(n9033), .A2(n7326), .ZN(n7325) );
  INV_X1 U7841 ( .A(n13063), .ZN(n7326) );
  XNOR2_X1 U7842 ( .A(n8928), .B(n11902), .ZN(n8938) );
  AND2_X1 U7843 ( .A1(n8964), .A2(n10382), .ZN(n7344) );
  AND2_X1 U7844 ( .A1(n6683), .A2(n6681), .ZN(n6680) );
  INV_X1 U7845 ( .A(n10677), .ZN(n6681) );
  INV_X1 U7846 ( .A(n7344), .ZN(n6686) );
  NAND2_X1 U7847 ( .A1(n13030), .A2(n13029), .ZN(n7343) );
  NAND2_X1 U7848 ( .A1(n7650), .A2(n11324), .ZN(n12045) );
  AND2_X1 U7849 ( .A1(n7465), .A2(n7495), .ZN(n7255) );
  NOR2_X2 U7850 ( .A1(n13304), .A2(n13529), .ZN(n13293) );
  AOI21_X1 U7851 ( .B1(n7088), .B2(n7087), .A(n6511), .ZN(n7086) );
  INV_X1 U7852 ( .A(n8012), .ZN(n7087) );
  INV_X1 U7853 ( .A(n12121), .ZN(n13295) );
  NAND2_X1 U7854 ( .A1(n7095), .A2(n7101), .ZN(n13307) );
  XNOR2_X1 U7855 ( .A(n13626), .B(n8011), .ZN(n12119) );
  NAND2_X1 U7856 ( .A1(n7085), .A2(n13384), .ZN(n13382) );
  INV_X1 U7857 ( .A(n13379), .ZN(n7085) );
  OR2_X1 U7858 ( .A1(n13441), .A2(n13440), .ZN(n8128) );
  NOR2_X1 U7859 ( .A1(n6503), .A2(n6458), .ZN(n6654) );
  AOI21_X1 U7860 ( .B1(n7136), .B2(n7134), .A(n6514), .ZN(n7133) );
  INV_X1 U7861 ( .A(n7139), .ZN(n7134) );
  OR2_X1 U7862 ( .A1(n13645), .A2(n13135), .ZN(n7128) );
  NAND2_X1 U7863 ( .A1(n7851), .A2(n6560), .ZN(n7127) );
  AND2_X1 U7864 ( .A1(n9451), .A2(n8159), .ZN(n13426) );
  OR2_X1 U7865 ( .A1(n10972), .A2(n12111), .ZN(n10970) );
  NAND2_X1 U7866 ( .A1(n10506), .A2(n12094), .ZN(n10505) );
  XNOR2_X1 U7867 ( .A(n8102), .B(n6595), .ZN(n6687) );
  NAND2_X1 U7868 ( .A1(n12065), .A2(n8157), .ZN(n13421) );
  NAND2_X1 U7869 ( .A1(n6617), .A2(n14860), .ZN(n11883) );
  INV_X1 U7870 ( .A(n13421), .ZN(n13459) );
  AND2_X1 U7871 ( .A1(n11881), .A2(n14860), .ZN(n10266) );
  NAND2_X1 U7872 ( .A1(n7873), .A2(n7872), .ZN(n13589) );
  AND2_X1 U7873 ( .A1(n9056), .A2(n7503), .ZN(n8770) );
  AND2_X1 U7874 ( .A1(n11882), .A2(n7508), .ZN(n14859) );
  AOI21_X1 U7875 ( .B1(n13665), .B2(n7484), .A(n13663), .ZN(n14846) );
  NOR2_X1 U7876 ( .A1(n7069), .A2(n7071), .ZN(n7070) );
  NOR2_X1 U7877 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n7068) );
  NAND2_X1 U7878 ( .A1(n7469), .A2(n7491), .ZN(n7488) );
  INV_X1 U7879 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n15080) );
  NAND2_X1 U7880 ( .A1(n7837), .A2(n7252), .ZN(n7935) );
  AND2_X1 U7881 ( .A1(n7253), .A2(n7496), .ZN(n7252) );
  INV_X1 U7882 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7496) );
  INV_X1 U7883 ( .A(n10164), .ZN(n10165) );
  INV_X1 U7884 ( .A(n10163), .ZN(n10166) );
  NAND2_X1 U7885 ( .A1(n13793), .A2(n11777), .ZN(n7279) );
  INV_X1 U7886 ( .A(n7270), .ZN(n7269) );
  OAI21_X1 U7887 ( .B1(n13768), .B2(n7271), .A(n13683), .ZN(n7270) );
  INV_X1 U7888 ( .A(n11827), .ZN(n7271) );
  INV_X1 U7889 ( .A(n14622), .ZN(n7262) );
  NOR2_X1 U7890 ( .A1(n7266), .A2(n10368), .ZN(n7261) );
  INV_X1 U7891 ( .A(n7440), .ZN(n7265) );
  INV_X1 U7892 ( .A(n7284), .ZN(n7283) );
  OAI21_X1 U7893 ( .B1(n7285), .B2(n10701), .A(n7287), .ZN(n7284) );
  NAND2_X1 U7894 ( .A1(n11213), .A2(n11212), .ZN(n7287) );
  NAND2_X1 U7895 ( .A1(n10641), .A2(n10642), .ZN(n7298) );
  NAND2_X1 U7896 ( .A1(n11668), .A2(n11669), .ZN(n6765) );
  NAND2_X1 U7897 ( .A1(n11368), .A2(n11367), .ZN(n13867) );
  NAND2_X1 U7898 ( .A1(n13947), .A2(n6956), .ZN(n13874) );
  NOR2_X1 U7899 ( .A1(n13866), .A2(n6957), .ZN(n6956) );
  NAND2_X1 U7900 ( .A1(n14132), .A2(n14123), .ZN(n6957) );
  NAND2_X1 U7901 ( .A1(n13942), .A2(n13892), .ZN(n13933) );
  NAND2_X1 U7902 ( .A1(n13942), .A2(n7196), .ZN(n14130) );
  NAND2_X1 U7903 ( .A1(n13947), .A2(n14132), .ZN(n13931) );
  AOI21_X1 U7904 ( .B1(n7187), .B2(n7185), .A(n6508), .ZN(n7184) );
  INV_X1 U7905 ( .A(n7187), .ZN(n7186) );
  NAND2_X1 U7906 ( .A1(n6941), .A2(n13987), .ZN(n7190) );
  NAND2_X1 U7907 ( .A1(n6628), .A2(n7188), .ZN(n7191) );
  INV_X1 U7908 ( .A(n13997), .ZN(n7353) );
  NAND2_X1 U7909 ( .A1(n6608), .A2(n14012), .ZN(n7354) );
  CLKBUF_X1 U7910 ( .A(n14010), .Z(n6628) );
  NAND2_X1 U7911 ( .A1(n14057), .A2(n7183), .ZN(n14051) );
  NAND2_X1 U7912 ( .A1(n14192), .A2(n13900), .ZN(n14040) );
  AND2_X1 U7913 ( .A1(n13897), .A2(n11674), .ZN(n14099) );
  AND2_X1 U7914 ( .A1(n11306), .A2(n14221), .ZN(n14086) );
  AOI21_X1 U7915 ( .B1(n11690), .B2(n6454), .A(n6509), .ZN(n7372) );
  OR2_X1 U7916 ( .A1(n13804), .A2(n14501), .ZN(n11471) );
  NAND2_X1 U7917 ( .A1(n11172), .A2(n11468), .ZN(n11177) );
  NAND2_X1 U7918 ( .A1(n11177), .A2(n11179), .ZN(n11272) );
  NAND2_X1 U7919 ( .A1(n10829), .A2(n10828), .ZN(n14538) );
  NAND2_X1 U7920 ( .A1(n10477), .A2(n10476), .ZN(n11440) );
  OR2_X1 U7921 ( .A1(n14685), .A2(n11435), .ZN(n10490) );
  NAND2_X1 U7922 ( .A1(n6446), .A2(n11411), .ZN(n7176) );
  NAND2_X1 U7923 ( .A1(n10144), .A2(n10171), .ZN(n10143) );
  NAND2_X1 U7924 ( .A1(n13937), .A2(n14767), .ZN(n14133) );
  XNOR2_X1 U7925 ( .A(n11653), .B(n11652), .ZN(n12060) );
  OAI21_X1 U7926 ( .B1(n8032), .B2(n6572), .A(n6738), .ZN(n8075) );
  INV_X1 U7927 ( .A(n6739), .ZN(n6738) );
  OAI21_X1 U7928 ( .B1(n6742), .B2(n6572), .A(n6976), .ZN(n6739) );
  NAND2_X1 U7929 ( .A1(n7618), .A2(SI_26_), .ZN(n6976) );
  XNOR2_X1 U7930 ( .A(n8075), .B(n8073), .ZN(n7634) );
  AND2_X1 U7931 ( .A1(n6776), .A2(n9165), .ZN(n9186) );
  AND2_X1 U7932 ( .A1(n9840), .A2(n7373), .ZN(n6776) );
  NOR2_X1 U7933 ( .A1(n9185), .A2(n9184), .ZN(n7444) );
  INV_X1 U7934 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9182) );
  XNOR2_X1 U7935 ( .A(n8060), .B(n8059), .ZN(n13661) );
  NAND2_X1 U7936 ( .A1(n6741), .A2(n7617), .ZN(n8060) );
  NAND2_X1 U7937 ( .A1(n8032), .A2(n6742), .ZN(n6741) );
  NAND4_X1 U7938 ( .A1(n7373), .A2(n9165), .A3(n6775), .A4(n6774), .ZN(n10257)
         );
  NOR2_X1 U7939 ( .A1(n9162), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n6775) );
  NAND2_X1 U7940 ( .A1(n7293), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9242) );
  AND2_X1 U7941 ( .A1(n7599), .A2(n7598), .ZN(n7983) );
  INV_X1 U7942 ( .A(n7964), .ZN(n7594) );
  NAND2_X1 U7943 ( .A1(n7593), .A2(n10033), .ZN(n7396) );
  OR2_X1 U7944 ( .A1(n7593), .A2(n10033), .ZN(n7595) );
  NAND2_X1 U7945 ( .A1(n7587), .A2(n7588), .ZN(n7406) );
  INV_X1 U7946 ( .A(n7931), .ZN(n7588) );
  INV_X1 U7947 ( .A(n6736), .ZN(n6733) );
  NAND2_X1 U7948 ( .A1(n7585), .A2(n7584), .ZN(n7919) );
  NAND2_X1 U7949 ( .A1(n7856), .A2(n6487), .ZN(n7400) );
  OR2_X1 U7950 ( .A1(n9202), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n9206) );
  XOR2_X1 U7951 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), .Z(
        n14333) );
  XNOR2_X1 U7952 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14295), .ZN(n14354) );
  NAND2_X1 U7953 ( .A1(n14402), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7216) );
  NAND2_X1 U7954 ( .A1(n10667), .A2(n8799), .ZN(n10809) );
  NAND2_X1 U7955 ( .A1(n8899), .A2(n8898), .ZN(n12150) );
  NAND2_X1 U7956 ( .A1(n10443), .A2(n6833), .ZN(n10548) );
  OR2_X1 U7957 ( .A1(n8794), .A2(n12353), .ZN(n6833) );
  NAND2_X1 U7958 ( .A1(n7420), .A2(n7421), .ZN(n11100) );
  INV_X1 U7959 ( .A(n7422), .ZN(n7421) );
  NAND2_X1 U7960 ( .A1(n10809), .A2(n6495), .ZN(n7420) );
  OAI21_X1 U7961 ( .B1(n8800), .B2(n7423), .A(n8802), .ZN(n7422) );
  AOI21_X1 U7962 ( .B1(n7427), .B2(n7425), .A(n6559), .ZN(n7424) );
  INV_X1 U7963 ( .A(n7427), .ZN(n7426) );
  INV_X1 U7964 ( .A(n12492), .ZN(n11352) );
  NAND2_X1 U7965 ( .A1(n10078), .A2(n10080), .ZN(n10079) );
  NAND2_X1 U7966 ( .A1(n10669), .A2(n10668), .ZN(n10667) );
  NAND4_X1 U7967 ( .A1(n8436), .A2(n8435), .A3(n8434), .A4(n8433), .ZN(n12842)
         );
  AND4_X1 U7968 ( .A1(n8370), .A2(n8369), .A3(n8368), .A4(n8367), .ZN(n12859)
         );
  XNOR2_X1 U7969 ( .A(n6902), .B(n9778), .ZN(n9813) );
  AOI21_X1 U7970 ( .B1(n14898), .B2(n9813), .A(n6900), .ZN(n9919) );
  NOR2_X1 U7971 ( .A1(n6901), .A2(n9778), .ZN(n6900) );
  INV_X1 U7972 ( .A(n6902), .ZN(n6901) );
  INV_X1 U7973 ( .A(n10520), .ZN(n7151) );
  OR2_X1 U7974 ( .A1(n11065), .A2(n6879), .ZN(n6878) );
  NOR2_X1 U7975 ( .A1(n6510), .A2(n11076), .ZN(n6879) );
  NAND2_X1 U7976 ( .A1(n6883), .A2(n6492), .ZN(n7158) );
  INV_X1 U7977 ( .A(n12504), .ZN(n12503) );
  INV_X1 U7978 ( .A(n7149), .ZN(n12533) );
  INV_X1 U7979 ( .A(n12550), .ZN(n12549) );
  INV_X1 U7980 ( .A(n7142), .ZN(n14453) );
  NAND2_X1 U7981 ( .A1(n6789), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7142) );
  AND2_X1 U7982 ( .A1(n7168), .A2(n6479), .ZN(n12557) );
  NAND2_X1 U7983 ( .A1(n6604), .A2(n8909), .ZN(n8910) );
  XNOR2_X1 U7984 ( .A(n8900), .B(n12461), .ZN(n12639) );
  NAND2_X1 U7985 ( .A1(n8893), .A2(n9077), .ZN(n8900) );
  OAI21_X1 U7986 ( .B1(n8708), .B2(n12858), .A(n8709), .ZN(n12642) );
  OAI21_X1 U7987 ( .B1(n6722), .B2(n12858), .A(n6719), .ZN(n12874) );
  NOR2_X1 U7988 ( .A1(n6721), .A2(n6720), .ZN(n6719) );
  XNOR2_X1 U7989 ( .A(n12652), .B(n12655), .ZN(n6722) );
  NOR2_X1 U7990 ( .A1(n12653), .A2(n12860), .ZN(n6720) );
  NAND2_X1 U7991 ( .A1(n8462), .A2(n8461), .ZN(n12914) );
  AND2_X1 U7992 ( .A1(n9085), .A2(n9084), .ZN(n12631) );
  NAND2_X1 U7993 ( .A1(n12633), .A2(n15049), .ZN(n6818) );
  INV_X1 U7994 ( .A(n12150), .ZN(n12637) );
  INV_X1 U7995 ( .A(n9148), .ZN(n12935) );
  NOR2_X1 U7996 ( .A1(n12874), .A2(n6718), .ZN(n12932) );
  AND2_X1 U7997 ( .A1(n12875), .A2(n15049), .ZN(n6718) );
  OR2_X1 U7998 ( .A1(n15050), .A2(n15044), .ZN(n12979) );
  AND2_X1 U7999 ( .A1(n6611), .A2(n8205), .ZN(n6610) );
  NAND2_X1 U8000 ( .A1(n7507), .A2(n7506), .ZN(n9455) );
  OAI21_X1 U8001 ( .B1(n10086), .B2(n7332), .A(n7330), .ZN(n10217) );
  INV_X1 U8002 ( .A(n7331), .ZN(n7330) );
  OAI21_X1 U8003 ( .B1(n6484), .B2(n7332), .A(n10218), .ZN(n7331) );
  INV_X1 U8004 ( .A(n8949), .ZN(n7332) );
  NAND2_X1 U8005 ( .A1(n7819), .A2(n7818), .ZN(n13600) );
  NAND2_X1 U8006 ( .A1(n10096), .A2(n10097), .ZN(n10095) );
  NAND2_X1 U8007 ( .A1(n7939), .A2(n7938), .ZN(n13562) );
  NAND2_X1 U8008 ( .A1(n10086), .A2(n6484), .ZN(n13099) );
  NOR2_X1 U8009 ( .A1(n13258), .A2(n7105), .ZN(n7104) );
  INV_X1 U8010 ( .A(n8070), .ZN(n7105) );
  NAND2_X1 U8011 ( .A1(n7969), .A2(n7968), .ZN(n13553) );
  NAND2_X1 U8012 ( .A1(n12042), .A2(n12041), .ZN(n13501) );
  NAND2_X1 U8013 ( .A1(n13500), .A2(n13502), .ZN(n13604) );
  NAND2_X1 U8014 ( .A1(n14261), .A2(n12059), .ZN(n6961) );
  INV_X1 U8015 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13649) );
  INV_X1 U8016 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n15202) );
  INV_X1 U8017 ( .A(n7460), .ZN(n7696) );
  AND2_X1 U8018 ( .A1(n10702), .A2(n10701), .ZN(n10921) );
  NAND2_X1 U8019 ( .A1(n6725), .A2(n11613), .ZN(n14142) );
  NAND2_X1 U8020 ( .A1(n6726), .A2(n11641), .ZN(n6725) );
  INV_X1 U8021 ( .A(n13659), .ZN(n6726) );
  NAND2_X1 U8022 ( .A1(n11571), .A2(n11570), .ZN(n14175) );
  NAND2_X1 U8023 ( .A1(n11530), .A2(n11529), .ZN(n14187) );
  OR2_X1 U8024 ( .A1(n11581), .A2(n11654), .ZN(n11584) );
  NAND2_X1 U8025 ( .A1(n11030), .A2(n11029), .ZN(n14570) );
  AND2_X1 U8026 ( .A1(n7274), .A2(n11754), .ZN(n7272) );
  INV_X1 U8027 ( .A(n14620), .ZN(n14527) );
  INV_X1 U8028 ( .A(n14004), .ZN(n14166) );
  AND2_X1 U8029 ( .A1(n14618), .A2(n14767), .ZN(n14525) );
  NOR3_X1 U8030 ( .A1(n11717), .A2(n11713), .A3(n11714), .ZN(n11715) );
  NAND2_X1 U8031 ( .A1(n7367), .A2(n13908), .ZN(n7362) );
  OAI21_X1 U8032 ( .B1(n13908), .B2(n7363), .A(n7359), .ZN(n7358) );
  AND2_X1 U8033 ( .A1(n11509), .A2(n11508), .ZN(n14211) );
  AND2_X1 U8034 ( .A1(n11498), .A2(n11497), .ZN(n14097) );
  NAND2_X1 U8035 ( .A1(n14339), .A2(n14340), .ZN(n14391) );
  NAND2_X1 U8036 ( .A1(n7206), .A2(n7203), .ZN(n6862) );
  INV_X1 U8037 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7203) );
  NOR2_X1 U8038 ( .A1(n14606), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7205) );
  AND2_X1 U8039 ( .A1(n11921), .A2(n7251), .ZN(n7250) );
  AND2_X1 U8040 ( .A1(n6443), .A2(n13812), .ZN(n11398) );
  AND2_X1 U8041 ( .A1(n9872), .A2(n11422), .ZN(n11397) );
  NAND2_X1 U8042 ( .A1(n6766), .A2(n11395), .ZN(n11386) );
  NAND2_X1 U8043 ( .A1(n11398), .A2(n11399), .ZN(n6766) );
  INV_X1 U8044 ( .A(n11386), .ZN(n11393) );
  OR2_X1 U8045 ( .A1(n11390), .A2(n11389), .ZN(n11394) );
  NAND2_X1 U8046 ( .A1(n11941), .A2(n11943), .ZN(n7243) );
  NAND2_X1 U8047 ( .A1(n11426), .A2(n6755), .ZN(n11429) );
  OAI21_X1 U8048 ( .B1(n11419), .B2(n6987), .A(n6756), .ZN(n6755) );
  NOR2_X1 U8049 ( .A1(n6757), .A2(n11425), .ZN(n6756) );
  NAND2_X1 U8050 ( .A1(n11969), .A2(n11971), .ZN(n7221) );
  OR2_X1 U8051 ( .A1(n11454), .A2(n11455), .ZN(n6761) );
  AOI21_X1 U8052 ( .B1(n6994), .B2(n6992), .A(n6990), .ZN(n6989) );
  NOR2_X1 U8053 ( .A1(n11474), .A2(n6457), .ZN(n6980) );
  INV_X1 U8054 ( .A(n6773), .ZN(n6770) );
  INV_X1 U8055 ( .A(n6768), .ZN(n6767) );
  OAI21_X1 U8056 ( .B1(n6979), .B2(n6773), .A(n6526), .ZN(n6768) );
  NOR2_X1 U8057 ( .A1(n6467), .A2(n6517), .ZN(n6979) );
  OR2_X1 U8058 ( .A1(n12000), .A2(n7220), .ZN(n6642) );
  NAND2_X1 U8059 ( .A1(n12000), .A2(n7220), .ZN(n7219) );
  INV_X1 U8060 ( .A(n11538), .ZN(n7003) );
  NOR2_X1 U8061 ( .A1(n11541), .A2(n11538), .ZN(n7004) );
  MUX2_X1 U8062 ( .A(n14180), .B(n14047), .S(n11422), .Z(n11557) );
  NAND2_X1 U8063 ( .A1(n6960), .A2(n6959), .ZN(n12038) );
  NAND2_X1 U8064 ( .A1(n13244), .A2(n12031), .ZN(n6959) );
  NAND2_X1 U8065 ( .A1(n13512), .A2(n12077), .ZN(n6960) );
  NAND2_X1 U8066 ( .A1(n7407), .A2(n7408), .ZN(n11597) );
  NAND2_X1 U8067 ( .A1(n11585), .A2(n11587), .ZN(n7408) );
  INV_X1 U8068 ( .A(n6999), .ZN(n6998) );
  INV_X1 U8069 ( .A(n11596), .ZN(n6754) );
  NAND2_X1 U8070 ( .A1(n7395), .A2(n7558), .ZN(n7394) );
  INV_X1 U8071 ( .A(n7814), .ZN(n7395) );
  OR2_X1 U8072 ( .A1(n8835), .A2(n8836), .ZN(n8841) );
  INV_X1 U8073 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8199) );
  NAND2_X1 U8074 ( .A1(n7312), .A2(n9026), .ZN(n9028) );
  NAND2_X1 U8075 ( .A1(n13067), .A2(n7313), .ZN(n7312) );
  INV_X1 U8076 ( .A(n12080), .ZN(n7230) );
  INV_X1 U8077 ( .A(n12081), .ZN(n7231) );
  NOR2_X1 U8078 ( .A1(n7791), .A2(n7790), .ZN(n7789) );
  OAI21_X1 U8079 ( .B1(n7107), .B2(n7066), .A(n10782), .ZN(n7065) );
  NOR2_X1 U8080 ( .A1(n10454), .A2(n7073), .ZN(n7072) );
  INV_X1 U8081 ( .A(n8114), .ZN(n7073) );
  NOR2_X1 U8082 ( .A1(n7080), .A2(n7077), .ZN(n7076) );
  INV_X1 U8083 ( .A(n8109), .ZN(n7077) );
  NAND2_X1 U8084 ( .A1(n10291), .A2(n8108), .ZN(n10021) );
  INV_X1 U8085 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7517) );
  INV_X1 U8086 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7518) );
  OAI21_X1 U8087 ( .B1(n6753), .B2(n6752), .A(n7386), .ZN(n11623) );
  NAND2_X1 U8088 ( .A1(n11610), .A2(n7387), .ZN(n7386) );
  AOI21_X1 U8089 ( .B1(n11597), .B2(n11598), .A(n6754), .ZN(n6753) );
  OAI21_X1 U8090 ( .B1(n11597), .B2(n11598), .A(n6522), .ZN(n6752) );
  NOR2_X1 U8091 ( .A1(n7403), .A2(n7399), .ZN(n7398) );
  INV_X1 U8092 ( .A(n7853), .ZN(n7399) );
  NAND2_X1 U8093 ( .A1(n7856), .A2(n7571), .ZN(n7867) );
  OAI21_X1 U8094 ( .B1(n11542), .B2(P2_DATAO_REG_11__SCAN_IN), .A(n6627), .ZN(
        n7560) );
  NAND2_X1 U8095 ( .A1(n11542), .A2(n9346), .ZN(n6627) );
  INV_X1 U8096 ( .A(n6966), .ZN(n6965) );
  OAI21_X1 U8097 ( .B1(n7545), .B2(n6967), .A(n7548), .ZN(n6966) );
  INV_X1 U8098 ( .A(n7547), .ZN(n6967) );
  OAI21_X1 U8099 ( .B1(n11542), .B2(n7532), .A(n7531), .ZN(n7534) );
  NAND2_X1 U8100 ( .A1(n11542), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7531) );
  INV_X1 U8101 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14286) );
  AOI21_X1 U8102 ( .B1(n14302), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n14301), .ZN(
        n14303) );
  AND2_X1 U8103 ( .A1(n14360), .A2(n14359), .ZN(n14301) );
  OR2_X1 U8104 ( .A1(n10197), .A2(n6779), .ZN(n6778) );
  AND2_X1 U8105 ( .A1(n10202), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6779) );
  AND2_X1 U8106 ( .A1(n6778), .A2(n14922), .ZN(n10198) );
  NAND2_X1 U8107 ( .A1(n10537), .A2(n10515), .ZN(n6786) );
  OAI211_X1 U8108 ( .C1(n14937), .C2(n6882), .A(n6881), .B(n10725), .ZN(n10992) );
  OR2_X1 U8109 ( .A1(n10540), .A2(n8301), .ZN(n6882) );
  NAND2_X1 U8110 ( .A1(n10539), .A2(n7169), .ZN(n6881) );
  NAND2_X1 U8111 ( .A1(n6622), .A2(n6621), .ZN(n6899) );
  INV_X1 U8112 ( .A(n11014), .ZN(n6621) );
  OR2_X1 U8113 ( .A1(n11077), .A2(n11078), .ZN(n7156) );
  NAND2_X1 U8114 ( .A1(n14462), .A2(n14461), .ZN(n6625) );
  OR2_X1 U8115 ( .A1(n12542), .A2(n14457), .ZN(n6619) );
  NOR2_X1 U8116 ( .A1(n7060), .A2(n6826), .ZN(n6825) );
  INV_X1 U8117 ( .A(n12445), .ZN(n6826) );
  INV_X1 U8118 ( .A(n12449), .ZN(n7060) );
  INV_X1 U8119 ( .A(n8704), .ZN(n7027) );
  OR2_X1 U8120 ( .A1(n8601), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8617) );
  NAND2_X1 U8121 ( .A1(n12788), .A2(n7043), .ZN(n7042) );
  NOR2_X1 U8122 ( .A1(n12855), .A2(n6696), .ZN(n6695) );
  INV_X1 U8123 ( .A(n8681), .ZN(n6696) );
  INV_X1 U8124 ( .A(n6801), .ZN(n6800) );
  OAI21_X1 U8125 ( .B1(n12300), .B2(n6802), .A(n12363), .ZN(n6801) );
  INV_X1 U8126 ( .A(n12361), .ZN(n6802) );
  AND2_X1 U8127 ( .A1(n10905), .A2(n10909), .ZN(n10906) );
  INV_X1 U8128 ( .A(n8258), .ZN(n8227) );
  AND2_X1 U8129 ( .A1(n7434), .A2(n6490), .ZN(n6904) );
  NAND2_X1 U8130 ( .A1(n8583), .A2(n8582), .ZN(n8584) );
  NAND2_X1 U8131 ( .A1(n8581), .A2(n8580), .ZN(n8583) );
  NAND2_X1 U8132 ( .A1(n8526), .A2(n8525), .ZN(n8527) );
  NAND2_X1 U8133 ( .A1(n8527), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8540) );
  AND2_X1 U8134 ( .A1(n8426), .A2(n8443), .ZN(n8459) );
  INV_X1 U8135 ( .A(n7432), .ZN(n8177) );
  INV_X1 U8136 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8377) );
  NOR2_X1 U8137 ( .A1(n13087), .A2(n7341), .ZN(n7340) );
  INV_X1 U8138 ( .A(n9004), .ZN(n7341) );
  AND2_X1 U8139 ( .A1(n7923), .A2(n7646), .ZN(n7955) );
  INV_X1 U8140 ( .A(n7340), .ZN(n7335) );
  AND2_X1 U8141 ( .A1(n9048), .A2(n9042), .ZN(n7342) );
  OAI21_X1 U8142 ( .B1(n13384), .B2(n7084), .A(n12115), .ZN(n7083) );
  NOR2_X1 U8143 ( .A1(n7877), .A2(n7876), .ZN(n7875) );
  AND2_X1 U8144 ( .A1(n7122), .A2(n6476), .ZN(n7121) );
  INV_X1 U8145 ( .A(n7125), .ZN(n7120) );
  OR2_X1 U8146 ( .A1(n11944), .A2(n11128), .ZN(n7139) );
  NOR2_X1 U8147 ( .A1(n13645), .A2(n11944), .ZN(n6928) );
  OR2_X1 U8148 ( .A1(n7860), .A2(n11127), .ZN(n7877) );
  AND2_X1 U8149 ( .A1(n7789), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7805) );
  NAND2_X1 U8150 ( .A1(n8043), .A2(n8042), .ZN(n13284) );
  XNOR2_X1 U8151 ( .A(n13145), .B(n10027), .ZN(n12098) );
  NAND2_X1 U8152 ( .A1(n6920), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7630) );
  AND2_X1 U8153 ( .A1(n7474), .A2(n7465), .ZN(n6690) );
  OR2_X1 U8154 ( .A1(n7801), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n7816) );
  NOR2_X2 U8155 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7670) );
  NOR2_X1 U8156 ( .A1(n9287), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9342) );
  NAND2_X1 U8157 ( .A1(n13893), .A2(n11698), .ZN(n13932) );
  OR2_X1 U8158 ( .A1(n13937), .A2(n14120), .ZN(n11698) );
  INV_X1 U8159 ( .A(n7188), .ZN(n7185) );
  INV_X1 U8160 ( .A(n11589), .ZN(n11588) );
  NAND2_X1 U8161 ( .A1(n14033), .A2(n13903), .ZN(n14013) );
  NOR2_X1 U8162 ( .A1(n11278), .A2(n11277), .ZN(n11308) );
  OR2_X1 U8163 ( .A1(n11183), .A2(n11182), .ZN(n11278) );
  NAND2_X1 U8164 ( .A1(n11044), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11183) );
  OR2_X1 U8165 ( .A1(n10490), .A2(n11440), .ZN(n6932) );
  INV_X1 U8166 ( .A(n7176), .ZN(n6597) );
  NAND2_X1 U8167 ( .A1(n11334), .A2(n14109), .ZN(n11383) );
  OAI21_X1 U8168 ( .B1(n8075), .B2(n7625), .A(n7624), .ZN(n11357) );
  AND2_X1 U8169 ( .A1(n7614), .A2(n6743), .ZN(n6742) );
  INV_X1 U8170 ( .A(n8044), .ZN(n6743) );
  AOI21_X1 U8171 ( .B1(n6450), .B2(n6750), .A(n6568), .ZN(n6745) );
  OAI21_X1 U8172 ( .B1(n7593), .B2(n6750), .A(n6746), .ZN(n7999) );
  NOR2_X1 U8173 ( .A1(n7917), .A2(n15122), .ZN(n6736) );
  NAND2_X1 U8174 ( .A1(n7917), .A2(n15122), .ZN(n6737) );
  NAND2_X1 U8175 ( .A1(n7581), .A2(n7580), .ZN(n7584) );
  INV_X1 U8176 ( .A(SI_16_), .ZN(n7580) );
  NOR2_X1 U8177 ( .A1(n7885), .A2(n7576), .ZN(n7577) );
  INV_X1 U8178 ( .A(n7571), .ZN(n7404) );
  INV_X1 U8179 ( .A(n6730), .ZN(n6729) );
  AND2_X1 U8180 ( .A1(n6728), .A2(n6549), .ZN(n6727) );
  AND2_X1 U8181 ( .A1(n7567), .A2(n7566), .ZN(n7829) );
  OR2_X1 U8182 ( .A1(n9282), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9287) );
  AND2_X1 U8183 ( .A1(n14283), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7210) );
  NOR2_X1 U8184 ( .A1(n14298), .A2(n14297), .ZN(n14330) );
  NOR2_X1 U8185 ( .A1(n14354), .A2(n14296), .ZN(n14297) );
  AOI21_X1 U8186 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14306), .A(n14305), .ZN(
        n14369) );
  NOR2_X1 U8187 ( .A1(n14325), .A2(n14324), .ZN(n14305) );
  OAI22_X1 U8188 ( .A1(n14977), .A2(P1_ADDR_REG_13__SCAN_IN), .B1(n14323), 
        .B2(n14310), .ZN(n14374) );
  AND2_X1 U8189 ( .A1(n6856), .A2(n6855), .ZN(n6853) );
  NAND2_X1 U8190 ( .A1(n7409), .A2(n10079), .ZN(n7411) );
  NOR2_X1 U8191 ( .A1(n10357), .A2(n7410), .ZN(n7409) );
  INV_X1 U8192 ( .A(n8792), .ZN(n7410) );
  OR2_X1 U8193 ( .A1(n9116), .A2(n9141), .ZN(n9121) );
  OR2_X1 U8194 ( .A1(n8778), .A2(n12477), .ZN(n8781) );
  AND2_X1 U8195 ( .A1(n12474), .A2(n8779), .ZN(n8780) );
  AND2_X1 U8196 ( .A1(n9132), .A2(n8857), .ZN(n9115) );
  NOR2_X1 U8197 ( .A1(n8822), .A2(n7419), .ZN(n7418) );
  INV_X1 U8198 ( .A(n8819), .ZN(n7419) );
  AND2_X1 U8199 ( .A1(n9137), .A2(n8854), .ZN(n12213) );
  OR2_X1 U8200 ( .A1(n11104), .A2(n8801), .ZN(n8802) );
  AND2_X1 U8201 ( .A1(n12176), .A2(n7428), .ZN(n7427) );
  NAND2_X1 U8202 ( .A1(n12250), .A2(n8829), .ZN(n7428) );
  INV_X1 U8203 ( .A(n8829), .ZN(n7425) );
  OR3_X1 U8204 ( .A1(n8383), .A2(P3_REG3_REG_11__SCAN_IN), .A3(
        P3_REG3_REG_12__SCAN_IN), .ZN(n8416) );
  OR2_X1 U8205 ( .A1(n11336), .A2(n11335), .ZN(n6856) );
  OR2_X1 U8206 ( .A1(n6485), .A2(n6837), .ZN(n6836) );
  NAND2_X1 U8207 ( .A1(n8835), .A2(n8836), .ZN(n6837) );
  INV_X1 U8208 ( .A(n6835), .ZN(n8846) );
  INV_X1 U8209 ( .A(n12498), .ZN(n10082) );
  INV_X1 U8210 ( .A(n8500), .ZN(n8499) );
  INV_X1 U8211 ( .A(n12497), .ZN(n8797) );
  OR2_X1 U8212 ( .A1(n8818), .A2(n12842), .ZN(n8819) );
  OAI21_X1 U8213 ( .B1(n11338), .B2(n6852), .A(n6848), .ZN(n8820) );
  AND2_X1 U8214 ( .A1(n10399), .A2(n10398), .ZN(n12280) );
  OR2_X1 U8215 ( .A1(n9763), .A2(n10254), .ZN(n9815) );
  AND2_X1 U8216 ( .A1(n9820), .A2(n9819), .ZN(n9822) );
  NAND2_X1 U8217 ( .A1(n9816), .A2(n9817), .ZN(n9930) );
  NOR2_X1 U8218 ( .A1(n15055), .A2(n14910), .ZN(n14909) );
  INV_X1 U8219 ( .A(n11325), .ZN(n14906) );
  OR2_X1 U8220 ( .A1(n10198), .A2(n6777), .ZN(n14925) );
  NOR2_X1 U8221 ( .A1(n6778), .A2(n14922), .ZN(n6777) );
  INV_X1 U8222 ( .A(n6887), .ZN(n6886) );
  NAND2_X1 U8223 ( .A1(n10195), .A2(n10196), .ZN(n10528) );
  NAND2_X1 U8224 ( .A1(n10719), .A2(n10720), .ZN(n11008) );
  AND2_X1 U8225 ( .A1(n14954), .A2(n10990), .ZN(n11075) );
  NAND2_X1 U8226 ( .A1(n7161), .A2(n11000), .ZN(n7160) );
  INV_X1 U8227 ( .A(n10999), .ZN(n7161) );
  INV_X1 U8228 ( .A(n6899), .ZN(n11071) );
  INV_X1 U8229 ( .A(n7156), .ZN(n12507) );
  NAND2_X1 U8230 ( .A1(n6790), .A2(n6482), .ZN(n7149) );
  NAND2_X1 U8231 ( .A1(n6903), .A2(n6575), .ZN(n12541) );
  AND2_X1 U8232 ( .A1(n6619), .A2(n6618), .ZN(n14462) );
  NAND2_X1 U8233 ( .A1(n12542), .A2(n14457), .ZN(n6618) );
  INV_X1 U8234 ( .A(n7168), .ZN(n14458) );
  INV_X1 U8235 ( .A(n6625), .ZN(n14464) );
  NAND2_X1 U8236 ( .A1(n6890), .A2(n6891), .ZN(n12573) );
  OR2_X1 U8237 ( .A1(n6479), .A2(n12556), .ZN(n6890) );
  NAND2_X1 U8238 ( .A1(n6893), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7168) );
  OAI21_X1 U8239 ( .B1(n12568), .B2(n6453), .A(n12567), .ZN(n12570) );
  NAND2_X1 U8240 ( .A1(n6844), .A2(n6843), .ZN(n8494) );
  INV_X1 U8241 ( .A(n8478), .ZN(n6844) );
  OR2_X1 U8242 ( .A1(n12565), .A2(n12784), .ZN(n7154) );
  OR2_X1 U8243 ( .A1(n12565), .A2(n6583), .ZN(n7152) );
  OR2_X1 U8244 ( .A1(n6475), .A2(n12582), .ZN(n7153) );
  INV_X1 U8245 ( .A(n12609), .ZN(n6620) );
  NAND2_X1 U8246 ( .A1(n6821), .A2(n6819), .ZN(n12271) );
  AOI21_X1 U8247 ( .B1(n6462), .B2(n7057), .A(n6820), .ZN(n6819) );
  INV_X1 U8248 ( .A(n12456), .ZN(n6820) );
  NAND2_X1 U8249 ( .A1(n9117), .A2(n7026), .ZN(n9077) );
  NOR2_X1 U8250 ( .A1(n7026), .A2(n12862), .ZN(n6721) );
  NOR2_X1 U8251 ( .A1(n12663), .A2(n12672), .ZN(n8700) );
  INV_X1 U8252 ( .A(n12665), .ZN(n12672) );
  NAND2_X1 U8253 ( .A1(n8562), .A2(n8561), .ZN(n8575) );
  AND4_X1 U8254 ( .A1(n8538), .A2(n8537), .A3(n8536), .A4(n8535), .ZN(n12733)
         );
  INV_X1 U8255 ( .A(n12730), .ZN(n6609) );
  INV_X1 U8256 ( .A(n12490), .ZN(n12745) );
  AND2_X1 U8257 ( .A1(n12765), .A2(n8691), .ZN(n12754) );
  NAND2_X1 U8258 ( .A1(n12754), .A2(n7446), .ZN(n12753) );
  NAND2_X1 U8259 ( .A1(n12797), .A2(n12406), .ZN(n12787) );
  NAND2_X1 U8260 ( .A1(n12787), .A2(n12788), .ZN(n12786) );
  NAND2_X1 U8261 ( .A1(n8463), .A2(n12195), .ZN(n8482) );
  AND2_X1 U8262 ( .A1(n12409), .A2(n12406), .ZN(n12798) );
  AOI21_X1 U8263 ( .B1(n6806), .B2(n6810), .A(n6805), .ZN(n6804) );
  AOI21_X1 U8264 ( .B1(n6455), .B2(n6694), .A(n6562), .ZN(n6692) );
  NAND2_X1 U8265 ( .A1(n12819), .A2(n12824), .ZN(n12818) );
  AOI21_X1 U8266 ( .B1(n7044), .B2(n6813), .A(n6812), .ZN(n6811) );
  INV_X1 U8267 ( .A(n7044), .ZN(n6814) );
  INV_X1 U8268 ( .A(n12387), .ZN(n6812) );
  OR2_X1 U8269 ( .A1(n8333), .A2(n8332), .ZN(n8352) );
  NAND2_X1 U8270 ( .A1(n10948), .A2(n8678), .ZN(n10949) );
  NAND2_X1 U8271 ( .A1(n6935), .A2(n8677), .ZN(n10933) );
  NAND2_X1 U8272 ( .A1(n8675), .A2(n8674), .ZN(n10656) );
  NAND2_X1 U8273 ( .A1(n8671), .A2(n6716), .ZN(n10558) );
  INV_X1 U8274 ( .A(n8785), .ZN(n6816) );
  INV_X1 U8275 ( .A(n12305), .ZN(n10299) );
  INV_X1 U8276 ( .A(n8668), .ZN(n10245) );
  NAND2_X1 U8277 ( .A1(n12285), .A2(n12284), .ZN(n14474) );
  NAND2_X1 U8278 ( .A1(n8600), .A2(n8599), .ZN(n8866) );
  NAND2_X1 U8279 ( .A1(n8587), .A2(n8586), .ZN(n12211) );
  NAND2_X1 U8280 ( .A1(n8547), .A2(n8546), .ZN(n12182) );
  OR2_X1 U8281 ( .A1(n10162), .A2(n12281), .ZN(n8547) );
  NAND2_X1 U8282 ( .A1(n11734), .A2(n11733), .ZN(n11737) );
  OAI22_X1 U8283 ( .A1(n9080), .A2(n9079), .B1(P1_DATAO_REG_28__SCAN_IN), .B2(
        n14264), .ZN(n9082) );
  NAND2_X1 U8284 ( .A1(n7433), .A2(n6905), .ZN(n7061) );
  INV_X1 U8285 ( .A(n7435), .ZN(n7433) );
  XNOR2_X1 U8286 ( .A(n8741), .B(n6905), .ZN(n9754) );
  NAND2_X1 U8287 ( .A1(n8541), .A2(n8540), .ZN(n8544) );
  NAND2_X1 U8288 ( .A1(n8544), .A2(n8543), .ZN(n8558) );
  OAI21_X1 U8289 ( .B1(n8527), .B2(P1_DATAO_REG_20__SCAN_IN), .A(n8540), .ZN(
        n8528) );
  NAND2_X1 U8290 ( .A1(n8508), .A2(n8507), .ZN(n8511) );
  AND2_X1 U8291 ( .A1(n8525), .A2(n8509), .ZN(n8510) );
  NAND2_X1 U8292 ( .A1(n6842), .A2(n6841), .ZN(n8513) );
  INV_X1 U8293 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n6841) );
  INV_X1 U8294 ( .A(n8494), .ZN(n6842) );
  AND2_X1 U8295 ( .A1(n8507), .A2(n8490), .ZN(n8491) );
  NAND2_X1 U8296 ( .A1(n8492), .A2(n8491), .ZN(n8508) );
  NAND2_X1 U8297 ( .A1(n7017), .A2(n7015), .ZN(n8476) );
  AOI21_X1 U8298 ( .B1(n7019), .B2(n7021), .A(n7016), .ZN(n7015) );
  INV_X1 U8299 ( .A(n8473), .ZN(n7016) );
  AND2_X1 U8300 ( .A1(n8488), .A2(n8474), .ZN(n8475) );
  NOR2_X1 U8301 ( .A1(n8274), .A2(n8177), .ZN(n8426) );
  AND2_X1 U8302 ( .A1(n9344), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8389) );
  AND2_X1 U8303 ( .A1(n8402), .A2(n8410), .ZN(n12514) );
  NAND2_X1 U8304 ( .A1(n7010), .A2(n7009), .ZN(n8361) );
  AOI21_X1 U8305 ( .B1(n7012), .B2(n7014), .A(n6530), .ZN(n7009) );
  NAND2_X1 U8306 ( .A1(n8327), .A2(n7012), .ZN(n7010) );
  AND2_X1 U8307 ( .A1(n8319), .A2(n8318), .ZN(n8323) );
  AND2_X1 U8308 ( .A1(n9220), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8291) );
  XNOR2_X1 U8309 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8306) );
  XNOR2_X1 U8310 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8276) );
  NAND2_X1 U8311 ( .A1(n9213), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8235) );
  XNOR2_X1 U8312 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8254) );
  NAND2_X1 U8313 ( .A1(n8225), .A2(n8224), .ZN(n8234) );
  XNOR2_X1 U8314 ( .A(n7511), .B(n7510), .ZN(n12090) );
  NOR2_X1 U8315 ( .A1(n13017), .A2(n7338), .ZN(n7337) );
  INV_X1 U8316 ( .A(n9009), .ZN(n7338) );
  NAND2_X1 U8317 ( .A1(n13046), .A2(n7340), .ZN(n7339) );
  NOR2_X1 U8318 ( .A1(n6664), .A2(n7318), .ZN(n6659) );
  NAND2_X1 U8319 ( .A1(n7321), .A2(n11245), .ZN(n7318) );
  NAND2_X1 U8320 ( .A1(n7322), .A2(n7324), .ZN(n7321) );
  AND2_X1 U8321 ( .A1(n7315), .A2(n6661), .ZN(n6660) );
  NAND2_X1 U8322 ( .A1(n6663), .A2(n6662), .ZN(n6661) );
  OAI21_X1 U8323 ( .B1(n7320), .B2(n7317), .A(n7316), .ZN(n7315) );
  NAND2_X1 U8324 ( .A1(n6655), .A2(n9032), .ZN(n9033) );
  NAND2_X1 U8325 ( .A1(n13008), .A2(n13007), .ZN(n13006) );
  NAND2_X1 U8326 ( .A1(n10384), .A2(n10383), .ZN(n8958) );
  OAI21_X1 U8327 ( .B1(n13046), .B2(n7336), .A(n7333), .ZN(n13068) );
  AOI21_X1 U8328 ( .B1(n7337), .B2(n7335), .A(n7334), .ZN(n7333) );
  INV_X1 U8329 ( .A(n7337), .ZN(n7336) );
  INV_X1 U8330 ( .A(n9015), .ZN(n7334) );
  NOR2_X1 U8331 ( .A1(n7311), .A2(n7306), .ZN(n7305) );
  NAND2_X1 U8332 ( .A1(n9027), .A2(n7310), .ZN(n7309) );
  NAND2_X1 U8333 ( .A1(n7308), .A2(n7306), .ZN(n7304) );
  INV_X1 U8334 ( .A(n7308), .ZN(n7307) );
  XNOR2_X1 U8335 ( .A(n8928), .B(n6635), .ZN(n8921) );
  NAND2_X1 U8336 ( .A1(n7343), .A2(n7342), .ZN(n13110) );
  NAND2_X1 U8337 ( .A1(n6665), .A2(n6663), .ZN(n11089) );
  OAI21_X1 U8338 ( .B1(n12036), .B2(n7224), .A(n6527), .ZN(n6646) );
  INV_X1 U8339 ( .A(n6614), .ZN(n8022) );
  OR2_X1 U8340 ( .A1(n7678), .A2(n9424), .ZN(n7663) );
  AND2_X1 U8341 ( .A1(n7255), .A2(n7254), .ZN(n7253) );
  INV_X1 U8342 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7254) );
  NOR2_X1 U8343 ( .A1(n6922), .A2(n12037), .ZN(n6921) );
  INV_X1 U8344 ( .A(n6923), .ZN(n6922) );
  NAND2_X1 U8345 ( .A1(n13261), .A2(n6923), .ZN(n13238) );
  AND2_X1 U8346 ( .A1(n13261), .A2(n13253), .ZN(n13250) );
  INV_X1 U8347 ( .A(n13247), .ZN(n13261) );
  AOI21_X1 U8348 ( .B1(n7096), .B2(n7099), .A(n7093), .ZN(n7092) );
  INV_X1 U8349 ( .A(n8149), .ZN(n7093) );
  INV_X1 U8350 ( .A(n8020), .ZN(n8036) );
  NAND2_X1 U8351 ( .A1(n13358), .A2(n6466), .ZN(n13304) );
  OR2_X1 U8352 ( .A1(n13324), .A2(n13323), .ZN(n13326) );
  NAND2_X1 U8353 ( .A1(n13358), .A2(n6915), .ZN(n13328) );
  NAND2_X1 U8354 ( .A1(n13358), .A2(n8103), .ZN(n13359) );
  OR2_X1 U8355 ( .A1(n13562), .A2(n13404), .ZN(n13394) );
  OR2_X1 U8356 ( .A1(n7910), .A2(n7909), .ZN(n7925) );
  NAND2_X1 U8357 ( .A1(n7130), .A2(n7129), .ZN(n13441) );
  AOI21_X1 U8358 ( .B1(n7131), .B2(n7137), .A(n6498), .ZN(n7129) );
  NOR2_X1 U8359 ( .A1(n13580), .A2(n6925), .ZN(n6924) );
  INV_X1 U8360 ( .A(n6926), .ZN(n6925) );
  NAND2_X1 U8361 ( .A1(n7135), .A2(n7139), .ZN(n11146) );
  OR2_X1 U8362 ( .A1(n11159), .A2(n8125), .ZN(n7135) );
  AND2_X1 U8363 ( .A1(n9451), .A2(n9481), .ZN(n13427) );
  NAND2_X1 U8364 ( .A1(n11167), .A2(n14493), .ZN(n11166) );
  NAND2_X1 U8365 ( .A1(n11167), .A2(n6928), .ZN(n13466) );
  AOI21_X1 U8366 ( .B1(n7114), .B2(n7827), .A(n11944), .ZN(n7113) );
  OR2_X1 U8367 ( .A1(n7844), .A2(n7843), .ZN(n7860) );
  AND2_X1 U8368 ( .A1(n10976), .A2(n10975), .ZN(n11167) );
  OAI21_X1 U8369 ( .B1(n10506), .B2(n7108), .A(n7106), .ZN(n10893) );
  AOI21_X1 U8370 ( .B1(n7109), .B2(n7107), .A(n6500), .ZN(n7106) );
  INV_X1 U8371 ( .A(n7109), .ZN(n7108) );
  NOR2_X1 U8372 ( .A1(n10890), .A2(n13479), .ZN(n10976) );
  OR2_X1 U8373 ( .A1(n10779), .A2(n13492), .ZN(n10890) );
  NAND2_X1 U8374 ( .A1(n7067), .A2(n7107), .ZN(n10499) );
  NOR2_X1 U8375 ( .A1(n10456), .A2(n11918), .ZN(n10502) );
  NAND2_X1 U8376 ( .A1(n6911), .A2(n6910), .ZN(n10456) );
  INV_X1 U8377 ( .A(n10429), .ZN(n6911) );
  NAND2_X1 U8378 ( .A1(n10584), .A2(n8110), .ZN(n10434) );
  NAND2_X1 U8379 ( .A1(n6913), .A2(n6912), .ZN(n10429) );
  NOR2_X1 U8380 ( .A1(n10286), .A2(n15068), .ZN(n10592) );
  NAND2_X1 U8381 ( .A1(n11898), .A2(n10585), .ZN(n10584) );
  NAND2_X1 U8382 ( .A1(n10019), .A2(n8109), .ZN(n10585) );
  NAND2_X1 U8383 ( .A1(n7091), .A2(n7096), .ZN(n13298) );
  OR2_X1 U8384 ( .A1(n13319), .A2(n7099), .ZN(n7091) );
  NAND2_X1 U8385 ( .A1(n7124), .A2(n7883), .ZN(n13448) );
  NAND2_X1 U8386 ( .A1(n7127), .A2(n7125), .ZN(n7124) );
  INV_X1 U8387 ( .A(n14864), .ZN(n14873) );
  INV_X1 U8388 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7641) );
  INV_X1 U8389 ( .A(n7476), .ZN(n7482) );
  NOR2_X1 U8390 ( .A1(n7770), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n7784) );
  OR2_X1 U8391 ( .A1(n7767), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n7770) );
  OR2_X1 U8392 ( .A1(n7835), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n7767) );
  CLKBUF_X1 U8393 ( .A(n7670), .Z(n7671) );
  AND2_X1 U8394 ( .A1(n11036), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n11044) );
  INV_X1 U8395 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9877) );
  OR2_X1 U8396 ( .A1(n10315), .A2(n10314), .ZN(n10340) );
  NOR2_X1 U8397 ( .A1(n10844), .A2(n10843), .ZN(n11036) );
  OR2_X1 U8398 ( .A1(n10836), .A2(n10835), .ZN(n10844) );
  AND2_X1 U8399 ( .A1(n7275), .A2(n6537), .ZN(n7274) );
  OR2_X1 U8400 ( .A1(n14523), .A2(n7278), .ZN(n7275) );
  NAND2_X1 U8401 ( .A1(n13767), .A2(n13768), .ZN(n13766) );
  NOR2_X1 U8402 ( .A1(n10340), .A2(n11218), .ZN(n10748) );
  NOR2_X1 U8403 ( .A1(n9878), .A2(n9877), .ZN(n9900) );
  NAND2_X1 U8404 ( .A1(n9899), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9714) );
  NOR2_X1 U8405 ( .A1(n6724), .A2(n13908), .ZN(n7357) );
  NAND2_X1 U8406 ( .A1(n7363), .A2(n7360), .ZN(n7359) );
  NAND2_X1 U8407 ( .A1(n7366), .A2(n7361), .ZN(n7360) );
  INV_X1 U8408 ( .A(n13932), .ZN(n13925) );
  NAND2_X1 U8409 ( .A1(n14029), .A2(n6937), .ZN(n13961) );
  NOR2_X1 U8410 ( .A1(n14150), .A2(n6939), .ZN(n6937) );
  AND2_X1 U8411 ( .A1(n13979), .A2(n7190), .ZN(n7187) );
  NAND2_X1 U8412 ( .A1(n14029), .A2(n6460), .ZN(n13999) );
  NAND2_X1 U8413 ( .A1(n14029), .A2(n14020), .ZN(n14015) );
  OR2_X1 U8414 ( .A1(n14180), .A2(n14047), .ZN(n13886) );
  OAI21_X1 U8415 ( .B1(n14057), .B2(n7182), .A(n7180), .ZN(n13887) );
  INV_X1 U8416 ( .A(n7181), .ZN(n7180) );
  NOR2_X1 U8417 ( .A1(n11531), .A2(n15206), .ZN(n11546) );
  NOR2_X1 U8418 ( .A1(n14069), .A2(n6950), .ZN(n6949) );
  INV_X1 U8419 ( .A(n6951), .ZN(n6950) );
  NAND2_X1 U8420 ( .A1(n6599), .A2(n6598), .ZN(n7174) );
  INV_X1 U8421 ( .A(n13881), .ZN(n6598) );
  NAND2_X1 U8422 ( .A1(n11306), .A2(n6459), .ZN(n14087) );
  AND2_X1 U8423 ( .A1(n11286), .A2(n11289), .ZN(n11306) );
  AND4_X1 U8424 ( .A1(n11041), .A2(n11040), .A3(n11039), .A4(n11038), .ZN(
        n14421) );
  NAND2_X1 U8425 ( .A1(n11042), .A2(n11061), .ZN(n11172) );
  NAND2_X1 U8426 ( .A1(n6948), .A2(n6947), .ZN(n14418) );
  INV_X1 U8427 ( .A(n14570), .ZN(n6947) );
  INV_X1 U8428 ( .A(n6948), .ZN(n14416) );
  OAI21_X1 U8429 ( .B1(n10762), .B2(n7384), .A(n7382), .ZN(n14536) );
  INV_X1 U8430 ( .A(n6932), .ZN(n10855) );
  NAND2_X1 U8431 ( .A1(n14688), .A2(n14687), .ZN(n14685) );
  OR2_X1 U8432 ( .A1(n10114), .A2(n10113), .ZN(n10315) );
  AND2_X1 U8433 ( .A1(n10123), .A2(n10654), .ZN(n14688) );
  NOR2_X1 U8434 ( .A1(n9898), .A2(n11417), .ZN(n10123) );
  NAND2_X1 U8435 ( .A1(n6631), .A2(n6501), .ZN(n9913) );
  OR2_X1 U8436 ( .A1(n10143), .A2(n11411), .ZN(n9898) );
  NAND2_X1 U8437 ( .A1(n9855), .A2(n9854), .ZN(n10142) );
  NAND2_X1 U8438 ( .A1(n9874), .A2(n9873), .ZN(n10140) );
  AND2_X1 U8439 ( .A1(n9740), .A2(n11399), .ZN(n10144) );
  AND2_X1 U8440 ( .A1(n14278), .A2(n11545), .ZN(n14180) );
  OR2_X1 U8441 ( .A1(n11377), .A2(n13816), .ZN(n14420) );
  INV_X1 U8442 ( .A(n14420), .ZN(n14745) );
  OAI21_X1 U8443 ( .B1(n9272), .B2(n9276), .A(n9275), .ZN(n9606) );
  NOR2_X1 U8444 ( .A1(n9592), .A2(n9677), .ZN(n9850) );
  XNOR2_X1 U8445 ( .A(n11357), .B(n11356), .ZN(n11642) );
  XNOR2_X1 U8446 ( .A(n9250), .B(n9249), .ZN(n9306) );
  INV_X1 U8447 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9249) );
  INV_X1 U8448 ( .A(n9178), .ZN(n9176) );
  NAND2_X1 U8449 ( .A1(n7999), .A2(SI_22_), .ZN(n8013) );
  NAND2_X1 U8450 ( .A1(n9172), .A2(n9244), .ZN(n9588) );
  AND2_X1 U8451 ( .A1(n7291), .A2(n9244), .ZN(n7290) );
  AND2_X1 U8452 ( .A1(n9167), .A2(n7292), .ZN(n7291) );
  NAND2_X1 U8453 ( .A1(n7800), .A2(n7556), .ZN(n7391) );
  XNOR2_X1 U8454 ( .A(n7766), .B(n7765), .ZN(n10310) );
  XNOR2_X1 U8455 ( .A(n7752), .B(n7751), .ZN(n10325) );
  NAND2_X1 U8456 ( .A1(n6964), .A2(n7547), .ZN(n7752) );
  NAND2_X1 U8457 ( .A1(n7737), .A2(n7545), .ZN(n6964) );
  AND2_X1 U8458 ( .A1(n9841), .A2(n9216), .ZN(n9261) );
  NOR2_X1 U8459 ( .A1(n9206), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9841) );
  INV_X1 U8460 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9163) );
  NAND2_X1 U8461 ( .A1(n7198), .A2(n14345), .ZN(n14348) );
  XNOR2_X1 U8462 ( .A(n14346), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n14347) );
  NAND2_X1 U8463 ( .A1(n14594), .A2(n6634), .ZN(n14371) );
  OAI21_X1 U8464 ( .B1(n14596), .B2(n14595), .A(P2_ADDR_REG_11__SCAN_IN), .ZN(
        n6634) );
  NOR2_X1 U8465 ( .A1(n14445), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6866) );
  NOR2_X1 U8466 ( .A1(n14445), .A2(n14440), .ZN(n6867) );
  INV_X1 U8467 ( .A(n12494), .ZN(n11104) );
  NAND2_X1 U8468 ( .A1(n10809), .A2(n10808), .ZN(n10807) );
  AND3_X1 U8469 ( .A1(n8313), .A2(n8312), .A3(n8311), .ZN(n10812) );
  NAND2_X1 U8470 ( .A1(n6847), .A2(n6851), .ZN(n12157) );
  NAND2_X1 U8471 ( .A1(n11338), .A2(n6853), .ZN(n6847) );
  AND3_X1 U8472 ( .A1(n8595), .A2(n8594), .A3(n8593), .ZN(n12705) );
  CLKBUF_X1 U8473 ( .A(n12168), .Z(n12169) );
  NAND2_X1 U8474 ( .A1(n11098), .A2(n6512), .ZN(n11228) );
  NAND2_X1 U8475 ( .A1(n11098), .A2(n8807), .ZN(n11227) );
  NAND2_X1 U8476 ( .A1(n10079), .A2(n8792), .ZN(n10356) );
  NAND2_X1 U8477 ( .A1(n10807), .A2(n8800), .ZN(n10881) );
  NAND2_X1 U8478 ( .A1(n10881), .A2(n10880), .ZN(n10879) );
  NAND2_X1 U8479 ( .A1(n7414), .A2(n6483), .ZN(n12194) );
  NAND2_X1 U8480 ( .A1(n8820), .A2(n7418), .ZN(n7414) );
  AOI21_X1 U8481 ( .B1(n7415), .B2(n7417), .A(n6564), .ZN(n7413) );
  NAND2_X1 U8482 ( .A1(n8531), .A2(n8530), .ZN(n12747) );
  OR2_X1 U8483 ( .A1(n10034), .A2(n12281), .ZN(n8531) );
  NAND2_X1 U8484 ( .A1(n8560), .A2(n8559), .ZN(n12722) );
  INV_X1 U8485 ( .A(n8789), .ZN(n8230) );
  OR2_X1 U8486 ( .A1(n12251), .A2(n12250), .ZN(n12252) );
  AND4_X1 U8487 ( .A1(n8305), .A2(n8304), .A3(n8303), .A4(n8302), .ZN(n10884)
         );
  OAI21_X2 U8488 ( .B1(n8863), .B2(n8862), .A(n8861), .ZN(n12216) );
  INV_X1 U8489 ( .A(n12216), .ZN(n14886) );
  NAND2_X1 U8490 ( .A1(n8820), .A2(n8819), .ZN(n12260) );
  INV_X1 U8491 ( .A(n14891), .ZN(n12268) );
  XNOR2_X1 U8492 ( .A(n6591), .B(n12612), .ZN(n12476) );
  AOI21_X1 U8493 ( .B1(n12294), .B2(n12293), .A(n12292), .ZN(n12295) );
  OR2_X1 U8494 ( .A1(n12470), .A2(n12291), .ZN(n12292) );
  AOI21_X1 U8495 ( .B1(n12635), .B2(n8207), .A(n8662), .ZN(n10227) );
  NAND2_X1 U8496 ( .A1(n8623), .A2(n8622), .ZN(n12668) );
  INV_X1 U8497 ( .A(n12653), .ZN(n12686) );
  NAND4_X1 U8498 ( .A1(n8288), .A2(n8287), .A3(n8286), .A4(n8285), .ZN(n12496)
         );
  NAND4_X1 U8499 ( .A1(n8250), .A2(n8249), .A3(n8248), .A4(n8247), .ZN(n12353)
         );
  OR2_X1 U8500 ( .A1(n8904), .A2(n8215), .ZN(n8218) );
  OR2_X1 U8501 ( .A1(n8238), .A2(n8206), .ZN(n8209) );
  NAND2_X1 U8502 ( .A1(n8207), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8208) );
  INV_X1 U8503 ( .A(n9932), .ZN(n14907) );
  INV_X1 U8504 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14935) );
  INV_X1 U8505 ( .A(n7172), .ZN(n14936) );
  NAND2_X1 U8506 ( .A1(n7170), .A2(n7169), .ZN(n10726) );
  INV_X1 U8507 ( .A(n7170), .ZN(n10541) );
  NOR2_X1 U8508 ( .A1(n10516), .A2(n10515), .ZN(n10517) );
  INV_X1 U8509 ( .A(n6889), .ZN(n14961) );
  INV_X1 U8510 ( .A(n7150), .ZN(n10985) );
  XNOR2_X1 U8511 ( .A(n11075), .B(n11076), .ZN(n10991) );
  NOR2_X1 U8512 ( .A1(n10991), .A2(n11004), .ZN(n11077) );
  OR2_X1 U8513 ( .A1(n14976), .A2(n12849), .ZN(n6790) );
  INV_X1 U8514 ( .A(n6883), .ZN(n14981) );
  AND2_X1 U8515 ( .A1(n12587), .A2(n12588), .ZN(n6909) );
  NAND2_X1 U8516 ( .A1(n7153), .A2(n7152), .ZN(n12600) );
  NAND2_X1 U8517 ( .A1(n7165), .A2(n7163), .ZN(n12614) );
  XNOR2_X1 U8518 ( .A(n12615), .B(n12616), .ZN(n6897) );
  AND3_X1 U8519 ( .A1(n7165), .A2(n7163), .A3(n12613), .ZN(n12615) );
  AND3_X1 U8520 ( .A1(n7153), .A2(n7152), .A3(n12599), .ZN(n12601) );
  XNOR2_X1 U8521 ( .A(n12271), .B(n12317), .ZN(n12633) );
  NAND2_X1 U8522 ( .A1(n8893), .A2(n8639), .ZN(n12648) );
  NAND2_X1 U8523 ( .A1(n7055), .A2(n12449), .ZN(n8638) );
  INV_X1 U8524 ( .A(n7038), .ZN(n12758) );
  NAND2_X1 U8525 ( .A1(n8689), .A2(n8688), .ZN(n12767) );
  NAND2_X1 U8526 ( .A1(n8481), .A2(n8480), .ZN(n12910) );
  NAND2_X1 U8527 ( .A1(n6639), .A2(n8685), .ZN(n6705) );
  NAND2_X1 U8528 ( .A1(n6808), .A2(n12397), .ZN(n12825) );
  NAND2_X1 U8529 ( .A1(n6809), .A2(n12396), .ZN(n6808) );
  INV_X1 U8530 ( .A(n12836), .ZN(n6809) );
  OAI21_X1 U8531 ( .B1(n8682), .B2(n6694), .A(n6455), .ZN(n12838) );
  NAND2_X1 U8532 ( .A1(n8682), .A2(n8681), .ZN(n12856) );
  NAND2_X1 U8533 ( .A1(n6954), .A2(n8680), .ZN(n11236) );
  OAI21_X1 U8534 ( .B1(n8331), .B2(n7049), .A(n7046), .ZN(n11238) );
  NAND2_X1 U8535 ( .A1(n7052), .A2(n12376), .ZN(n11115) );
  NAND2_X1 U8536 ( .A1(n8331), .A2(n7053), .ZN(n7052) );
  INV_X1 U8537 ( .A(n10812), .ZN(n15027) );
  NAND2_X1 U8538 ( .A1(n6799), .A2(n12361), .ZN(n10769) );
  NAND2_X1 U8539 ( .A1(n10903), .A2(n12300), .ZN(n6799) );
  NOR2_X1 U8540 ( .A1(n12868), .A2(n10244), .ZN(n12647) );
  NAND2_X1 U8541 ( .A1(n8518), .A2(n8517), .ZN(n12962) );
  NAND2_X1 U8542 ( .A1(n8429), .A2(n8428), .ZN(n12976) );
  AND2_X1 U8543 ( .A1(n8726), .A2(n8725), .ZN(n10055) );
  AND2_X1 U8544 ( .A1(n9754), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12981) );
  XNOR2_X1 U8545 ( .A(n8895), .B(n8628), .ZN(n12155) );
  NAND2_X1 U8546 ( .A1(n8716), .A2(n8715), .ZN(n10818) );
  AND2_X1 U8547 ( .A1(n8643), .A2(n8642), .ZN(n12484) );
  XNOR2_X1 U8548 ( .A(n8647), .B(n6829), .ZN(n12329) );
  INV_X1 U8549 ( .A(n8757), .ZN(n10032) );
  INV_X1 U8550 ( .A(SI_19_), .ZN(n15087) );
  INV_X1 U8551 ( .A(SI_17_), .ZN(n15122) );
  NAND2_X1 U8552 ( .A1(n7018), .A2(n8456), .ZN(n8472) );
  NAND2_X1 U8553 ( .A1(n8455), .A2(n8454), .ZN(n7018) );
  INV_X1 U8554 ( .A(SI_14_), .ZN(n9302) );
  INV_X1 U8555 ( .A(SI_13_), .ZN(n9299) );
  NAND2_X1 U8556 ( .A1(n7034), .A2(n8423), .ZN(n8422) );
  INV_X1 U8557 ( .A(SI_12_), .ZN(n9268) );
  XNOR2_X1 U8558 ( .A(n8358), .B(P3_IR_REG_10__SCAN_IN), .ZN(n14967) );
  NAND2_X1 U8559 ( .A1(n7011), .A2(n8328), .ZN(n8346) );
  NAND2_X1 U8560 ( .A1(n6603), .A2(n8326), .ZN(n7011) );
  XNOR2_X1 U8561 ( .A(n8290), .B(n8289), .ZN(n10525) );
  INV_X1 U8562 ( .A(n8173), .ZN(n8251) );
  NAND2_X1 U8563 ( .A1(n7173), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8220) );
  NAND2_X1 U8564 ( .A1(n6486), .A2(P3_IR_REG_1__SCAN_IN), .ZN(n7144) );
  AND2_X1 U8565 ( .A1(n12090), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9155) );
  NAND2_X1 U8566 ( .A1(n13110), .A2(n9049), .ZN(n12999) );
  NAND2_X1 U8567 ( .A1(n6682), .A2(n6683), .ZN(n10678) );
  OR2_X1 U8568 ( .A1(n10384), .A2(n6686), .ZN(n6682) );
  NAND2_X1 U8569 ( .A1(n7951), .A2(n7950), .ZN(n13559) );
  OAI211_X1 U8570 ( .C1(n7343), .C2(n6672), .A(n6668), .B(n6666), .ZN(n9062)
         );
  NAND2_X1 U8571 ( .A1(n6675), .A2(n9054), .ZN(n6672) );
  OAI21_X1 U8572 ( .B1(n6673), .B2(n9054), .A(n6669), .ZN(n6668) );
  NOR2_X1 U8573 ( .A1(n13512), .A2(n13122), .ZN(n9063) );
  NAND2_X1 U8574 ( .A1(n13067), .A2(n9021), .ZN(n13023) );
  NAND2_X1 U8575 ( .A1(n7908), .A2(n7907), .ZN(n13577) );
  NAND2_X1 U8576 ( .A1(n13006), .A2(n9033), .ZN(n13062) );
  INV_X1 U8577 ( .A(n10067), .ZN(n8935) );
  XNOR2_X1 U8578 ( .A(n8938), .B(n8937), .ZN(n10067) );
  NAND2_X1 U8579 ( .A1(n8958), .A2(n10382), .ZN(n10617) );
  OAI211_X1 U8580 ( .C1(n13067), .C2(n7307), .A(n7299), .B(n6478), .ZN(n13078)
         );
  NAND2_X1 U8581 ( .A1(n13067), .A2(n7305), .ZN(n7299) );
  NAND2_X1 U8582 ( .A1(n6680), .A2(n6686), .ZN(n6678) );
  NAND2_X1 U8583 ( .A1(n13046), .A2(n9004), .ZN(n13088) );
  AND2_X1 U8584 ( .A1(n10086), .A2(n8943), .ZN(n13101) );
  NAND2_X1 U8585 ( .A1(n7343), .A2(n9042), .ZN(n13113) );
  NAND2_X1 U8586 ( .A1(n9961), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13118) );
  AND2_X1 U8587 ( .A1(n7681), .A2(n6544), .ZN(n6589) );
  OR2_X1 U8588 ( .A1(n8094), .A2(n10268), .ZN(n7658) );
  AND2_X1 U8589 ( .A1(n7837), .A2(n7465), .ZN(n7870) );
  NAND2_X1 U8590 ( .A1(n7837), .A2(n7255), .ZN(n7892) );
  AOI21_X1 U8591 ( .B1(n8166), .B2(n13421), .A(n8165), .ZN(n11729) );
  NAND2_X1 U8592 ( .A1(n13256), .A2(n6465), .ZN(n13230) );
  NAND2_X1 U8593 ( .A1(n8071), .A2(n8070), .ZN(n13257) );
  NAND2_X1 U8594 ( .A1(n8062), .A2(n8061), .ZN(n13520) );
  NAND2_X1 U8595 ( .A1(n8047), .A2(n8046), .ZN(n13525) );
  NAND2_X1 U8596 ( .A1(n7100), .A2(n8146), .ZN(n13308) );
  OR2_X1 U8597 ( .A1(n13319), .A2(n12119), .ZN(n7100) );
  NAND2_X1 U8598 ( .A1(n8018), .A2(n8017), .ZN(n13313) );
  NAND2_X1 U8599 ( .A1(n13382), .A2(n7945), .ZN(n13365) );
  NAND2_X1 U8600 ( .A1(n7132), .A2(n7133), .ZN(n13458) );
  OR2_X1 U8601 ( .A1(n11159), .A2(n7137), .ZN(n7132) );
  NAND2_X1 U8602 ( .A1(n7127), .A2(n7128), .ZN(n13456) );
  NAND2_X1 U8603 ( .A1(n7118), .A2(n7813), .ZN(n10969) );
  NAND2_X1 U8604 ( .A1(n10505), .A2(n8119), .ZN(n10781) );
  NAND2_X1 U8605 ( .A1(n7074), .A2(n8114), .ZN(n10457) );
  NAND2_X1 U8606 ( .A1(n13490), .A2(n10570), .ZN(n13474) );
  AND2_X1 U8607 ( .A1(n13490), .A2(n15069), .ZN(n13493) );
  INV_X1 U8608 ( .A(n13410), .ZN(n14833) );
  INV_X1 U8609 ( .A(n13501), .ZN(n13607) );
  NAND2_X1 U8610 ( .A1(n12063), .A2(n12062), .ZN(n13610) );
  OR2_X1 U8611 ( .A1(n11268), .A2(n6636), .ZN(n8003) );
  NAND2_X1 U8612 ( .A1(n7922), .A2(n7921), .ZN(n13634) );
  AND2_X1 U8613 ( .A1(n9455), .A2(n9155), .ZN(n14854) );
  XNOR2_X1 U8614 ( .A(n7062), .B(n7628), .ZN(n13658) );
  NAND2_X1 U8615 ( .A1(n7631), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7062) );
  NAND2_X1 U8616 ( .A1(n7481), .A2(n7480), .ZN(n11271) );
  INV_X1 U8617 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11269) );
  NAND2_X1 U8618 ( .A1(n7488), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7489) );
  INV_X1 U8619 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10077) );
  INV_X1 U8620 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9990) );
  INV_X1 U8621 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9846) );
  INV_X1 U8622 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9676) );
  INV_X1 U8623 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9346) );
  INV_X1 U8624 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9220) );
  INV_X1 U8625 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9204) );
  INV_X1 U8626 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9214) );
  INV_X1 U8627 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9212) );
  CLKBUF_X1 U8628 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n13673) );
  NAND2_X1 U8629 ( .A1(n13766), .A2(n11827), .ZN(n13684) );
  NAND2_X1 U8630 ( .A1(n10739), .A2(n11641), .ZN(n10742) );
  NAND2_X1 U8631 ( .A1(n10168), .A2(n10167), .ZN(n14621) );
  AND3_X1 U8632 ( .A1(n11312), .A2(n11311), .A3(n11310), .ZN(n14202) );
  NOR2_X1 U8633 ( .A1(n13691), .A2(n7281), .ZN(n7280) );
  INV_X1 U8634 ( .A(n11799), .ZN(n7281) );
  NAND2_X1 U8635 ( .A1(n7282), .A2(n11799), .ZN(n13692) );
  OR2_X1 U8636 ( .A1(n10921), .A2(n7285), .ZN(n11214) );
  NOR2_X1 U8637 ( .A1(n10921), .A2(n10920), .ZN(n10922) );
  NAND2_X1 U8638 ( .A1(n13757), .A2(n11812), .ZN(n13702) );
  NAND2_X1 U8639 ( .A1(n7273), .A2(n7274), .ZN(n13710) );
  NAND2_X1 U8640 ( .A1(n11276), .A2(n11275), .ZN(n14227) );
  AND2_X1 U8641 ( .A1(n11300), .A2(n11299), .ZN(n14221) );
  AOI21_X1 U8642 ( .B1(n7269), .B2(n7271), .A(n6513), .ZN(n7267) );
  XNOR2_X1 U8643 ( .A(n11837), .B(n11838), .ZN(n13750) );
  NAND2_X1 U8644 ( .A1(n7265), .A2(n10368), .ZN(n7264) );
  AND2_X1 U8645 ( .A1(n14513), .A2(n14511), .ZN(n11762) );
  INV_X1 U8646 ( .A(n14097), .ZN(n14214) );
  AND2_X1 U8647 ( .A1(n7298), .A2(n10646), .ZN(n7295) );
  AND2_X1 U8648 ( .A1(n7294), .A2(n7298), .ZN(n10647) );
  NAND2_X1 U8649 ( .A1(n6764), .A2(n6461), .ZN(n6762) );
  INV_X1 U8650 ( .A(n13867), .ZN(n14115) );
  INV_X1 U8651 ( .A(n13874), .ZN(n13873) );
  AOI21_X1 U8652 ( .B1(n12060), .B2(n11641), .A(n11656), .ZN(n14118) );
  INV_X1 U8653 ( .A(n14155), .ZN(n14139) );
  AND2_X1 U8654 ( .A1(n13944), .A2(n13954), .ZN(n6644) );
  NAND2_X1 U8655 ( .A1(n7191), .A2(n7190), .ZN(n13993) );
  NAND2_X1 U8656 ( .A1(n7191), .A2(n7187), .ZN(n14160) );
  NAND2_X1 U8657 ( .A1(n7348), .A2(n7350), .ZN(n13978) );
  AND2_X1 U8658 ( .A1(n7354), .A2(n7355), .ZN(n13998) );
  NAND2_X1 U8659 ( .A1(n7354), .A2(n7352), .ZN(n14164) );
  NAND2_X1 U8660 ( .A1(n6628), .A2(n13889), .ZN(n13996) );
  NAND2_X1 U8661 ( .A1(n14051), .A2(n13885), .ZN(n14026) );
  INV_X1 U8662 ( .A(n14187), .ZN(n14049) );
  NOR2_X1 U8663 ( .A1(n7381), .A2(n14058), .ZN(n7380) );
  INV_X1 U8664 ( .A(n13898), .ZN(n7381) );
  NAND2_X1 U8665 ( .A1(n14079), .A2(n13898), .ZN(n14059) );
  NAND2_X1 U8666 ( .A1(n7370), .A2(n7372), .ZN(n11304) );
  NAND2_X1 U8667 ( .A1(n11272), .A2(n11471), .ZN(n11302) );
  NAND2_X1 U8668 ( .A1(n11176), .A2(n11175), .ZN(n13804) );
  INV_X1 U8669 ( .A(n14558), .ZN(n14504) );
  NAND2_X1 U8670 ( .A1(n11035), .A2(n11034), .ZN(n11767) );
  NAND2_X1 U8671 ( .A1(n11060), .A2(n11059), .ZN(n11062) );
  NOR2_X1 U8672 ( .A1(n11061), .A2(n7179), .ZN(n7178) );
  INV_X1 U8673 ( .A(n11059), .ZN(n7179) );
  NOR2_X1 U8674 ( .A1(n11379), .A2(n11703), .ZN(n7288) );
  NAND2_X1 U8675 ( .A1(n10834), .A2(n10833), .ZN(n13712) );
  NAND2_X1 U8676 ( .A1(n7385), .A2(n10762), .ZN(n14762) );
  AND2_X1 U8677 ( .A1(n10762), .A2(n10761), .ZN(n10764) );
  AND2_X1 U8678 ( .A1(n7377), .A2(n10334), .ZN(n10337) );
  NAND2_X1 U8679 ( .A1(n7377), .A2(n7376), .ZN(n10479) );
  NAND2_X1 U8680 ( .A1(n7378), .A2(n7379), .ZN(n7377) );
  INV_X1 U8681 ( .A(n7175), .ZN(n10102) );
  AOI21_X1 U8682 ( .B1(n9893), .B2(n7176), .A(n6491), .ZN(n7175) );
  INV_X1 U8683 ( .A(n14700), .ZN(n14544) );
  INV_X1 U8684 ( .A(n14096), .ZN(n14683) );
  INV_X1 U8685 ( .A(n14066), .ZN(n14690) );
  NAND2_X1 U8686 ( .A1(n9851), .A2(n14706), .ZN(n14437) );
  INV_X2 U8687 ( .A(n14787), .ZN(n14790) );
  INV_X1 U8688 ( .A(n14124), .ZN(n14127) );
  AND2_X1 U8689 ( .A1(n14134), .A2(n14133), .ZN(n14135) );
  OR2_X1 U8690 ( .A1(n9722), .A2(n9847), .ZN(n14775) );
  XNOR2_X1 U8691 ( .A(n11366), .B(n11365), .ZN(n14254) );
  OAI21_X1 U8692 ( .B1(n11653), .B2(n11651), .A(n11362), .ZN(n11366) );
  INV_X1 U8693 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9614) );
  XNOR2_X1 U8694 ( .A(n8080), .B(n8079), .ZN(n14261) );
  NAND2_X1 U8695 ( .A1(n8077), .A2(n8076), .ZN(n8080) );
  NAND2_X1 U8696 ( .A1(n8077), .A2(n7637), .ZN(n13659) );
  CLKBUF_X1 U8697 ( .A(n9307), .Z(n14631) );
  NAND2_X1 U8698 ( .A1(n9186), .A2(n7444), .ZN(n9248) );
  NAND2_X1 U8699 ( .A1(n8014), .A2(n8013), .ZN(n8016) );
  XNOR2_X1 U8700 ( .A(n11544), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14278) );
  NAND2_X1 U8701 ( .A1(n6626), .A2(n9679), .ZN(n11544) );
  OAI21_X1 U8702 ( .B1(n10257), .B2(n9246), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9247) );
  NAND2_X1 U8703 ( .A1(n6751), .A2(n6749), .ZN(n7982) );
  NAND2_X1 U8704 ( .A1(n7595), .A2(n7396), .ZN(n7965) );
  INV_X1 U8705 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10259) );
  NAND2_X1 U8706 ( .A1(n7405), .A2(n7589), .ZN(n7934) );
  INV_X1 U8707 ( .A(n7406), .ZN(n7405) );
  INV_X1 U8708 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9995) );
  INV_X1 U8709 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9844) );
  INV_X1 U8710 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9948) );
  INV_X1 U8711 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9423) );
  INV_X1 U8712 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9292) );
  INV_X1 U8713 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n15155) );
  INV_X1 U8714 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9263) );
  INV_X1 U8715 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9237) );
  INV_X1 U8716 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9218) );
  INV_X1 U8717 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7532) );
  INV_X1 U8718 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14337) );
  AOI21_X1 U8719 ( .B1(n14392), .B2(n14341), .A(n14389), .ZN(n15246) );
  XNOR2_X1 U8720 ( .A(n14332), .B(n7199), .ZN(n15240) );
  INV_X1 U8721 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7199) );
  XNOR2_X1 U8722 ( .A(n14347), .B(n14348), .ZN(n15241) );
  INV_X1 U8723 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7212) );
  INV_X1 U8724 ( .A(n14362), .ZN(n7217) );
  INV_X1 U8725 ( .A(n14365), .ZN(n7215) );
  XNOR2_X1 U8726 ( .A(n14371), .B(n14370), .ZN(n14598) );
  NAND2_X1 U8727 ( .A1(n7200), .A2(n6858), .ZN(n14372) );
  INV_X1 U8728 ( .A(n14599), .ZN(n6858) );
  NAND2_X1 U8729 ( .A1(n6862), .A2(n6860), .ZN(n14380) );
  NOR2_X1 U8730 ( .A1(n14603), .A2(n6861), .ZN(n6860) );
  INV_X1 U8731 ( .A(n14606), .ZN(n6861) );
  INV_X1 U8732 ( .A(n6878), .ZN(n11070) );
  INV_X1 U8733 ( .A(n7158), .ZN(n12505) );
  INV_X1 U8734 ( .A(n6789), .ZN(n14454) );
  AND2_X1 U8735 ( .A1(n7142), .A2(n6496), .ZN(n12538) );
  INV_X1 U8736 ( .A(n8910), .ZN(n12641) );
  AND2_X1 U8737 ( .A1(n9108), .A2(n7033), .ZN(n7032) );
  OR2_X1 U8738 ( .A1(n15066), .A2(n9107), .ZN(n7033) );
  OR2_X1 U8739 ( .A1(n12631), .A2(n12928), .ZN(n9108) );
  NOR2_X1 U8740 ( .A1(n6606), .A2(n6502), .ZN(n6605) );
  NOR2_X1 U8741 ( .A1(n15066), .A2(n8911), .ZN(n6606) );
  OR2_X1 U8742 ( .A1(n15066), .A2(n8766), .ZN(n6955) );
  NAND2_X1 U8743 ( .A1(n6717), .A2(n6471), .ZN(n12877) );
  NAND2_X1 U8744 ( .A1(n12932), .A2(n15066), .ZN(n6717) );
  AND2_X1 U8745 ( .A1(n9105), .A2(n6578), .ZN(n6817) );
  OR2_X1 U8746 ( .A1(n12631), .A2(n12979), .ZN(n9105) );
  OAI21_X1 U8747 ( .B1(n8765), .B2(n15050), .A(n6470), .ZN(P3_U3454) );
  NAND2_X1 U8748 ( .A1(n13099), .A2(n8949), .ZN(n10219) );
  AND2_X1 U8749 ( .A1(n10095), .A2(n8926), .ZN(n10039) );
  NAND2_X1 U8750 ( .A1(n6931), .A2(n6930), .ZN(P2_U3530) );
  AOI21_X1 U8751 ( .B1(n13501), .B2(n13596), .A(n6573), .ZN(n6930) );
  NAND2_X1 U8752 ( .A1(n13604), .A2(n14885), .ZN(n6931) );
  INV_X1 U8753 ( .A(n6653), .ZN(n6652) );
  OAI21_X1 U8754 ( .B1(n8774), .B2(n8170), .A(n8168), .ZN(n6653) );
  AND2_X1 U8755 ( .A1(n13512), .A2(n13596), .ZN(n6615) );
  NAND2_X1 U8756 ( .A1(n6651), .A2(n6650), .ZN(P2_U3495) );
  AOI22_X1 U8757 ( .A1(n13512), .A2(n13646), .B1(P2_REG0_REG_28__SCAN_IN), 
        .B2(n14879), .ZN(n6650) );
  NAND2_X1 U8758 ( .A1(n13612), .A2(n14880), .ZN(n6651) );
  OAI21_X1 U8759 ( .B1(n14257), .B2(n13666), .A(n7327), .ZN(P2_U3297) );
  NOR2_X1 U8760 ( .A1(n7329), .A2(n7328), .ZN(n7327) );
  AOI21_X1 U8761 ( .B1(n11743), .B2(n11742), .A(n7442), .ZN(n14524) );
  INV_X1 U8762 ( .A(n7206), .ZN(n14602) );
  AND2_X1 U8763 ( .A1(n6862), .A2(n7207), .ZN(n14607) );
  OAI21_X1 U8764 ( .B1(n14444), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6872), .ZN(
        n7208) );
  INV_X2 U8765 ( .A(n11926), .ZN(n12030) );
  MUX2_X2 U8766 ( .A(n6978), .B(n11379), .S(n11663), .Z(n11422) );
  NOR2_X1 U8767 ( .A1(n8676), .A2(n10906), .ZN(n6449) );
  AND2_X1 U8768 ( .A1(n6746), .A2(n6561), .ZN(n6450) );
  OR2_X1 U8769 ( .A1(n7594), .A2(SI_20_), .ZN(n6451) );
  AND2_X1 U8770 ( .A1(n9684), .A2(n9610), .ZN(n6452) );
  INV_X1 U8771 ( .A(n12094), .ZN(n7107) );
  INV_X1 U8772 ( .A(n13954), .ZN(n7365) );
  AND2_X1 U8773 ( .A1(n6625), .A2(n6619), .ZN(n6453) );
  INV_X1 U8774 ( .A(n14012), .ZN(n7351) );
  AND2_X1 U8775 ( .A1(n11471), .A2(n11692), .ZN(n6454) );
  INV_X1 U8776 ( .A(n6689), .ZN(n6688) );
  INV_X2 U8777 ( .A(n12077), .ZN(n12031) );
  AND2_X1 U8778 ( .A1(n12839), .A2(n6505), .ZN(n6455) );
  AND2_X1 U8779 ( .A1(n14142), .A2(n14147), .ZN(n6456) );
  NOR3_X1 U8780 ( .A1(n11480), .A2(n11479), .A3(n11485), .ZN(n6457) );
  INV_X1 U8781 ( .A(n6852), .ZN(n6851) );
  NOR2_X1 U8782 ( .A1(n6854), .A2(n12231), .ZN(n6852) );
  INV_X1 U8783 ( .A(n12489), .ZN(n7026) );
  NOR2_X1 U8784 ( .A1(n13580), .A2(n13425), .ZN(n6458) );
  INV_X1 U8785 ( .A(n7323), .ZN(n7322) );
  INV_X1 U8786 ( .A(n7137), .ZN(n7136) );
  NAND2_X1 U8787 ( .A1(n8126), .A2(n7138), .ZN(n7137) );
  AND2_X1 U8788 ( .A1(n14097), .A2(n14221), .ZN(n6459) );
  INV_X1 U8789 ( .A(n14445), .ZN(n6873) );
  AND2_X1 U8790 ( .A1(n14020), .A2(n6941), .ZN(n6460) );
  OR2_X1 U8791 ( .A1(n11672), .A2(n11671), .ZN(n6461) );
  AND2_X1 U8792 ( .A1(n6823), .A2(n6827), .ZN(n6462) );
  NOR2_X1 U8793 ( .A1(n11435), .A2(n10478), .ZN(n6463) );
  OAI21_X1 U8794 ( .B1(n7999), .B2(SI_22_), .A(n8013), .ZN(n11543) );
  INV_X1 U8795 ( .A(n11543), .ZN(n6626) );
  NAND2_X1 U8796 ( .A1(n8845), .A2(n8846), .ZN(n12240) );
  AND2_X1 U8797 ( .A1(n7434), .A2(n6518), .ZN(n6464) );
  AND2_X1 U8798 ( .A1(n13233), .A2(n8072), .ZN(n6465) );
  INV_X1 U8799 ( .A(n8990), .ZN(n7324) );
  NAND2_X1 U8800 ( .A1(n11608), .A2(n11607), .ZN(n14150) );
  AND2_X1 U8801 ( .A1(n6915), .A2(n6914), .ZN(n6466) );
  NOR2_X1 U8802 ( .A1(n6981), .A2(n6457), .ZN(n6467) );
  INV_X1 U8803 ( .A(n14132), .ZN(n13937) );
  AND2_X1 U8804 ( .A1(n11634), .A2(n11633), .ZN(n14132) );
  INV_X1 U8805 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7459) );
  NAND2_X1 U8806 ( .A1(n7986), .A2(n7985), .ZN(n13549) );
  INV_X1 U8807 ( .A(n13549), .ZN(n6918) );
  AND2_X1 U8808 ( .A1(n6528), .A2(n8674), .ZN(n6468) );
  NOR3_X1 U8809 ( .A1(n6558), .A2(n14073), .A3(n14572), .ZN(n6469) );
  NAND2_X1 U8810 ( .A1(n7339), .A2(n9009), .ZN(n13016) );
  INV_X1 U8811 ( .A(n13512), .ZN(n13613) );
  NAND2_X1 U8812 ( .A1(n6961), .A2(n8081), .ZN(n13512) );
  NAND2_X1 U8813 ( .A1(n11167), .A2(n6926), .ZN(n6929) );
  AND2_X1 U8814 ( .A1(n8752), .A2(n6574), .ZN(n6470) );
  NAND2_X1 U8815 ( .A1(n10499), .A2(n7781), .ZN(n10778) );
  INV_X1 U8816 ( .A(n9609), .ZN(n6978) );
  INV_X1 U8817 ( .A(n11908), .ZN(n6912) );
  OR2_X1 U8818 ( .A1(n15066), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n6471) );
  NOR2_X1 U8819 ( .A1(n12537), .A2(n14455), .ZN(n6472) );
  NOR2_X1 U8820 ( .A1(n12556), .A2(n14460), .ZN(n6473) );
  AND3_X1 U8821 ( .A1(n8218), .A2(n8217), .A3(n8216), .ZN(n6474) );
  INV_X1 U8822 ( .A(n11858), .ZN(n10169) );
  OR2_X1 U8823 ( .A1(n12591), .A2(n12580), .ZN(n6475) );
  INV_X1 U8824 ( .A(n14078), .ZN(n6771) );
  NAND2_X1 U8825 ( .A1(n13645), .A2(n13135), .ZN(n6476) );
  AND4_X1 U8826 ( .A1(n7474), .A2(n7473), .A3(n7472), .A4(n7471), .ZN(n6477)
         );
  INV_X1 U8827 ( .A(n9027), .ZN(n7311) );
  NAND2_X1 U8828 ( .A1(n6701), .A2(n8697), .ZN(n12661) );
  AND2_X1 U8829 ( .A1(n7304), .A2(n7309), .ZN(n6478) );
  NAND2_X1 U8830 ( .A1(n14457), .A2(n12552), .ZN(n6479) );
  NAND2_X1 U8831 ( .A1(n8187), .A2(n8188), .ZN(n8245) );
  NOR2_X1 U8832 ( .A1(n12223), .A2(n12224), .ZN(n6480) );
  AND2_X1 U8833 ( .A1(n9103), .A2(n9102), .ZN(n6481) );
  OR2_X1 U8834 ( .A1(n12511), .A2(n12510), .ZN(n6482) );
  OR2_X1 U8835 ( .A1(n8821), .A2(n12160), .ZN(n6483) );
  AND2_X1 U8836 ( .A1(n13100), .A2(n8943), .ZN(n6484) );
  NAND4_X1 U8837 ( .A1(n8194), .A2(n8193), .A3(n8192), .A4(n8191), .ZN(n8666)
         );
  OR2_X1 U8838 ( .A1(n12998), .A2(n6677), .ZN(n6676) );
  NAND2_X1 U8839 ( .A1(n6477), .A2(n7070), .ZN(n7631) );
  NOR2_X1 U8840 ( .A1(n8833), .A2(n12183), .ZN(n6485) );
  NAND2_X1 U8841 ( .A1(n8219), .A2(n6474), .ZN(n12499) );
  INV_X1 U8842 ( .A(n7200), .ZN(n14600) );
  AND2_X1 U8843 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n6486) );
  NAND2_X1 U8844 ( .A1(n6822), .A2(n7056), .ZN(n8893) );
  XNOR2_X1 U8845 ( .A(n13775), .B(n14047), .ZN(n13902) );
  INV_X1 U8846 ( .A(n13902), .ZN(n6630) );
  NAND2_X1 U8847 ( .A1(n7268), .A2(n7267), .ZN(n13749) );
  NAND2_X1 U8848 ( .A1(n12252), .A2(n8829), .ZN(n12175) );
  NOR2_X1 U8849 ( .A1(n7578), .A2(n7404), .ZN(n6487) );
  INV_X1 U8850 ( .A(n13908), .ZN(n7361) );
  NAND2_X1 U8851 ( .A1(n7841), .A2(n7840), .ZN(n11944) );
  NAND2_X1 U8852 ( .A1(n8981), .A2(n8980), .ZN(n6488) );
  AND2_X1 U8853 ( .A1(n8989), .A2(n7324), .ZN(n6489) );
  INV_X1 U8854 ( .A(n14922), .ZN(n10203) );
  NAND2_X1 U8855 ( .A1(n6705), .A2(n8686), .ZN(n12780) );
  AND2_X1 U8856 ( .A1(n8180), .A2(n6905), .ZN(n6490) );
  INV_X1 U8857 ( .A(n13967), .ZN(n14147) );
  NAND2_X1 U8858 ( .A1(n13326), .A2(n8012), .ZN(n13314) );
  AND2_X1 U8859 ( .A1(n11410), .A2(n11409), .ZN(n6491) );
  INV_X1 U8860 ( .A(n11703), .ZN(n14022) );
  OR2_X1 U8861 ( .A1(n12511), .A2(n12503), .ZN(n6492) );
  INV_X1 U8862 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14918) );
  AND3_X2 U8863 ( .A1(n7676), .A2(n7675), .A3(n7674), .ZN(n10135) );
  INV_X1 U8864 ( .A(n10135), .ZN(n11885) );
  INV_X1 U8865 ( .A(n11692), .ZN(n11301) );
  NAND2_X1 U8866 ( .A1(n14057), .A2(n13883), .ZN(n14050) );
  XNOR2_X1 U8867 ( .A(n14142), .B(n13967), .ZN(n13954) );
  AND2_X1 U8868 ( .A1(n10204), .A2(n10203), .ZN(n6493) );
  NAND2_X1 U8869 ( .A1(n7400), .A2(n7577), .ZN(n7890) );
  INV_X1 U8870 ( .A(n10880), .ZN(n7423) );
  OR3_X1 U8871 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        P3_IR_REG_1__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U8872 ( .A1(n8851), .A2(n12212), .ZN(n12167) );
  AND2_X1 U8873 ( .A1(n10880), .A2(n10808), .ZN(n6495) );
  NAND2_X1 U8874 ( .A1(n14457), .A2(n12535), .ZN(n6496) );
  INV_X1 U8875 ( .A(n11611), .ZN(n7387) );
  OR2_X1 U8876 ( .A1(n14358), .A2(n14357), .ZN(n6497) );
  NAND2_X1 U8877 ( .A1(n11644), .A2(n11643), .ZN(n13909) );
  AND2_X1 U8878 ( .A1(n13589), .A2(n12093), .ZN(n6498) );
  MUX2_X1 U8879 ( .A(n14142), .B(n13967), .S(n6443), .Z(n11624) );
  OR2_X1 U8880 ( .A1(n14371), .A2(n14370), .ZN(n6499) );
  XNOR2_X1 U8881 ( .A(n13514), .B(n13126), .ZN(n13258) );
  INV_X1 U8882 ( .A(n11409), .ZN(n11411) );
  NAND2_X1 U8883 ( .A1(n7895), .A2(n7894), .ZN(n13580) );
  AND2_X1 U8884 ( .A1(n11516), .A2(n11515), .ZN(n14197) );
  INV_X1 U8885 ( .A(n13514), .ZN(n13253) );
  OAI21_X2 U8886 ( .B1(n13659), .B2(n6636), .A(n7638), .ZN(n13514) );
  AND2_X1 U8887 ( .A1(n13492), .A2(n8120), .ZN(n6500) );
  OR2_X1 U8888 ( .A1(n11410), .A2(n11411), .ZN(n6501) );
  INV_X1 U8889 ( .A(n11455), .ZN(n6990) );
  NOR2_X1 U8890 ( .A1(n7353), .A2(n13904), .ZN(n7352) );
  NOR2_X1 U8891 ( .A1(n12637), .A2(n12928), .ZN(n6502) );
  AND2_X1 U8892 ( .A1(n7122), .A2(n7120), .ZN(n6503) );
  AND2_X1 U8893 ( .A1(n12597), .A2(n6906), .ZN(n6504) );
  OR2_X1 U8894 ( .A1(n6695), .A2(n6694), .ZN(n6505) );
  NAND2_X1 U8895 ( .A1(n14029), .A2(n6938), .ZN(n6942) );
  AND2_X1 U8896 ( .A1(n8235), .A2(n8224), .ZN(n6506) );
  INV_X1 U8897 ( .A(n7057), .ZN(n7056) );
  NAND2_X1 U8898 ( .A1(n12452), .A2(n7058), .ZN(n7057) );
  NAND2_X1 U8899 ( .A1(n7028), .A2(n7027), .ZN(n6507) );
  NAND2_X1 U8900 ( .A1(n13358), .A2(n6916), .ZN(n6919) );
  AND2_X1 U8901 ( .A1(n13983), .A2(n14004), .ZN(n6508) );
  AND2_X1 U8902 ( .A1(n14227), .A2(n13802), .ZN(n6509) );
  AND2_X1 U8903 ( .A1(n14958), .A2(n10999), .ZN(n6510) );
  INV_X1 U8904 ( .A(n11451), .ZN(n6993) );
  AND2_X1 U8905 ( .A1(n13313), .A2(n13129), .ZN(n6511) );
  NAND2_X1 U8906 ( .A1(n7633), .A2(n7632), .ZN(n12037) );
  INV_X1 U8907 ( .A(n12396), .ZN(n6810) );
  AND2_X1 U8908 ( .A1(n8808), .A2(n8807), .ZN(n6512) );
  AND2_X1 U8909 ( .A1(n11833), .A2(n11832), .ZN(n6513) );
  INV_X1 U8910 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n6905) );
  INV_X1 U8911 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7629) );
  INV_X1 U8912 ( .A(n11474), .ZN(n6983) );
  NOR2_X1 U8913 ( .A1(n13645), .A2(n13463), .ZN(n6514) );
  NOR2_X1 U8914 ( .A1(n14170), .A2(n13987), .ZN(n6515) );
  INV_X1 U8915 ( .A(n11689), .ZN(n11061) );
  NAND2_X1 U8916 ( .A1(n8845), .A2(n6834), .ZN(n12241) );
  XOR2_X1 U8917 ( .A(n14452), .B(n14451), .Z(n6516) );
  NAND2_X1 U8918 ( .A1(n11495), .A2(n11494), .ZN(n6517) );
  NOR2_X1 U8919 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n6518) );
  NOR2_X1 U8920 ( .A1(n14132), .A2(n14120), .ZN(n6519) );
  INV_X1 U8921 ( .A(n10540), .ZN(n7169) );
  INV_X1 U8922 ( .A(n11690), .ZN(n11179) );
  OR2_X1 U8923 ( .A1(n6463), .A2(n10335), .ZN(n6520) );
  AND4_X1 U8924 ( .A1(n7432), .A2(n7430), .A3(n8173), .A4(n6828), .ZN(n8712)
         );
  OR2_X1 U8925 ( .A1(n7429), .A2(n8177), .ZN(n6521) );
  OR2_X1 U8926 ( .A1(n7387), .A2(n11610), .ZN(n6522) );
  INV_X1 U8927 ( .A(n6917), .ZN(n6916) );
  NAND2_X1 U8928 ( .A1(n8103), .A2(n6918), .ZN(n6917) );
  INV_X1 U8929 ( .A(n6939), .ZN(n6938) );
  NAND2_X1 U8930 ( .A1(n6460), .A2(n6940), .ZN(n6939) );
  AND2_X1 U8931 ( .A1(n7549), .A2(SI_7_), .ZN(n6523) );
  NOR2_X1 U8932 ( .A1(n9051), .A2(n9050), .ZN(n6524) );
  INV_X1 U8933 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7626) );
  OR2_X1 U8934 ( .A1(n7265), .A2(n10368), .ZN(n6525) );
  AND2_X1 U8935 ( .A1(n6772), .A2(n6771), .ZN(n6526) );
  AND2_X1 U8936 ( .A1(n7227), .A2(n7226), .ZN(n6527) );
  NOR2_X1 U8937 ( .A1(n12346), .A2(n8676), .ZN(n6528) );
  INV_X1 U8938 ( .A(n7197), .ZN(n7196) );
  NAND2_X1 U8939 ( .A1(n13925), .A2(n13892), .ZN(n7197) );
  OR2_X1 U8940 ( .A1(n14284), .A2(n14918), .ZN(n6529) );
  AND2_X1 U8941 ( .A1(n15155), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n6530) );
  INV_X1 U8942 ( .A(n7416), .ZN(n7415) );
  OAI21_X1 U8943 ( .B1(n7418), .B2(n7417), .A(n12193), .ZN(n7416) );
  INV_X1 U8944 ( .A(n7367), .ZN(n7366) );
  NOR2_X1 U8945 ( .A1(n6456), .A2(n6519), .ZN(n7367) );
  INV_X1 U8946 ( .A(n7089), .ZN(n7088) );
  NAND2_X1 U8947 ( .A1(n7090), .A2(n8028), .ZN(n7089) );
  OAI22_X1 U8948 ( .A1(n11667), .A2(n11670), .B1(n11668), .B2(n11669), .ZN(
        n6764) );
  AND2_X1 U8949 ( .A1(n8796), .A2(n8797), .ZN(n6531) );
  OAI21_X1 U8950 ( .B1(n6787), .B2(n7146), .A(n6786), .ZN(n6783) );
  INV_X1 U8951 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9344) );
  NAND2_X1 U8952 ( .A1(n8092), .A2(n8091), .ZN(n13233) );
  INV_X1 U8953 ( .A(n6958), .ZN(n13910) );
  NOR2_X1 U8954 ( .A1(n13931), .A2(n13909), .ZN(n6958) );
  INV_X1 U8955 ( .A(n6676), .ZN(n6675) );
  NAND2_X1 U8956 ( .A1(n12034), .A2(n12057), .ZN(n6532) );
  AND3_X1 U8957 ( .A1(n12130), .A2(n7508), .A3(n12131), .ZN(n6533) );
  NOR2_X1 U8958 ( .A1(n11542), .A2(n9257), .ZN(n6534) );
  OR2_X1 U8959 ( .A1(n13589), .A2(n12093), .ZN(n6535) );
  OR2_X1 U8960 ( .A1(n14348), .A2(n14347), .ZN(n6536) );
  OR2_X1 U8961 ( .A1(n11749), .A2(n11748), .ZN(n6537) );
  AND3_X1 U8962 ( .A1(n6713), .A2(n6712), .A3(n6711), .ZN(n6538) );
  AND2_X1 U8963 ( .A1(n14144), .A2(n14145), .ZN(n6539) );
  INV_X1 U8964 ( .A(n14281), .ZN(n14336) );
  NAND2_X1 U8965 ( .A1(n6863), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14281) );
  INV_X1 U8966 ( .A(n7028), .ZN(n12452) );
  NAND2_X1 U8967 ( .A1(n7022), .A2(n12455), .ZN(n7028) );
  NAND2_X1 U8968 ( .A1(n8637), .A2(n8636), .ZN(n12489) );
  AND2_X1 U8969 ( .A1(n7345), .A2(n7629), .ZN(n6540) );
  INV_X1 U8970 ( .A(n7781), .ZN(n7066) );
  AND2_X1 U8971 ( .A1(n11780), .A2(n11782), .ZN(n6541) );
  AND2_X1 U8972 ( .A1(n8690), .A2(n8688), .ZN(n6542) );
  NOR2_X1 U8973 ( .A1(n12824), .A2(n6807), .ZN(n6806) );
  INV_X1 U8974 ( .A(n7945), .ZN(n7084) );
  AND2_X1 U8975 ( .A1(n8201), .A2(n8203), .ZN(n6543) );
  AND2_X1 U8976 ( .A1(n7680), .A2(n7682), .ZN(n6544) );
  AND2_X1 U8977 ( .A1(n11814), .A2(n11812), .ZN(n6545) );
  OR2_X1 U8978 ( .A1(n11574), .A2(n11572), .ZN(n6546) );
  INV_X1 U8979 ( .A(n11921), .ZN(n7249) );
  AND2_X1 U8980 ( .A1(n7167), .A2(n7166), .ZN(n6547) );
  OR2_X1 U8981 ( .A1(n11941), .A2(n11943), .ZN(n6548) );
  AND2_X1 U8982 ( .A1(n7392), .A2(n6968), .ZN(n6549) );
  AND2_X1 U8983 ( .A1(n7154), .A2(n6475), .ZN(n6550) );
  AND2_X1 U8984 ( .A1(n6690), .A2(n15123), .ZN(n6551) );
  INV_X1 U8985 ( .A(n13884), .ZN(n14053) );
  AND2_X1 U8986 ( .A1(n13885), .A2(n11673), .ZN(n13884) );
  NAND2_X1 U8987 ( .A1(n12010), .A2(n7235), .ZN(n6552) );
  NAND2_X1 U8988 ( .A1(n11981), .A2(n7238), .ZN(n6553) );
  NAND2_X1 U8989 ( .A1(n11992), .A2(n7241), .ZN(n6554) );
  INV_X1 U8990 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8184) );
  INV_X1 U8991 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n6843) );
  AND2_X1 U8992 ( .A1(n6751), .A2(n6451), .ZN(n6555) );
  INV_X1 U8993 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9166) );
  INV_X1 U8994 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9187) );
  NAND2_X1 U8995 ( .A1(n11970), .A2(n7223), .ZN(n6556) );
  INV_X1 U8996 ( .A(n6664), .ZN(n6663) );
  NAND2_X1 U8997 ( .A1(n11090), .A2(n6488), .ZN(n6664) );
  NAND2_X1 U8998 ( .A1(n12498), .A2(n8793), .ZN(n6557) );
  NAND2_X2 U8999 ( .A1(n14859), .A2(n12091), .ZN(n13262) );
  INV_X1 U9000 ( .A(n11000), .ZN(n11076) );
  INV_X1 U9001 ( .A(n13313), .ZN(n6914) );
  INV_X1 U9002 ( .A(n10537), .ZN(n7145) );
  NAND4_X1 U9003 ( .A1(n8339), .A2(n8338), .A3(n8337), .A4(n8336), .ZN(n12493)
         );
  CLKBUF_X3 U9004 ( .A(n7475), .Z(n7837) );
  INV_X1 U9005 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n6713) );
  NAND2_X1 U9006 ( .A1(n11595), .A2(n11594), .ZN(n13983) );
  INV_X1 U9007 ( .A(n13983), .ZN(n6940) );
  NAND2_X1 U9008 ( .A1(n8630), .A2(n8629), .ZN(n9117) );
  INV_X1 U9009 ( .A(n6750), .ZN(n6749) );
  NAND2_X1 U9010 ( .A1(n6451), .A2(n7983), .ZN(n6750) );
  INV_X1 U9011 ( .A(n14138), .ZN(n14120) );
  NAND2_X1 U9012 ( .A1(n7273), .A2(n7272), .ZN(n13708) );
  AND2_X1 U9013 ( .A1(n11306), .A2(n6951), .ZN(n6558) );
  NAND2_X1 U9014 ( .A1(n7193), .A2(n11296), .ZN(n13878) );
  INV_X1 U9015 ( .A(n12406), .ZN(n7043) );
  NAND2_X1 U9016 ( .A1(n11584), .A2(n11583), .ZN(n14170) );
  INV_X1 U9017 ( .A(n14170), .ZN(n6941) );
  INV_X1 U9018 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n6829) );
  NAND2_X1 U9019 ( .A1(n7279), .A2(n11780), .ZN(n13726) );
  NOR2_X1 U9020 ( .A1(n6945), .A2(n9162), .ZN(n9840) );
  INV_X1 U9021 ( .A(n11458), .ZN(n6759) );
  AND2_X1 U9022 ( .A1(n6665), .A2(n6488), .ZN(n11088) );
  AND2_X1 U9023 ( .A1(n8830), .A2(n12491), .ZN(n6559) );
  AND2_X1 U9024 ( .A1(n7852), .A2(n6476), .ZN(n6560) );
  OR2_X1 U9025 ( .A1(n8000), .A2(n15215), .ZN(n6561) );
  AND2_X1 U9026 ( .A1(n12847), .A2(n12821), .ZN(n6562) );
  NAND2_X1 U9027 ( .A1(n14221), .A2(n14210), .ZN(n6563) );
  AND2_X1 U9028 ( .A1(n8824), .A2(n12805), .ZN(n6564) );
  INV_X1 U9029 ( .A(n12231), .ZN(n6855) );
  AND2_X1 U9030 ( .A1(n7339), .A2(n7337), .ZN(n6565) );
  INV_X1 U9031 ( .A(n9778), .ZN(n9812) );
  NOR2_X1 U9032 ( .A1(n14205), .A2(n14193), .ZN(n6566) );
  NAND2_X1 U9033 ( .A1(n7837), .A2(n7253), .ZN(n6567) );
  OR2_X1 U9034 ( .A1(n8015), .A2(n7605), .ZN(n6568) );
  INV_X1 U9035 ( .A(n6946), .ZN(n11181) );
  NOR2_X1 U9036 ( .A1(n14418), .A2(n11767), .ZN(n6946) );
  AND2_X1 U9037 ( .A1(n7584), .A2(n6737), .ZN(n6569) );
  AND2_X1 U9038 ( .A1(n8768), .A2(n6955), .ZN(n6570) );
  OR2_X1 U9039 ( .A1(n6759), .A2(n11457), .ZN(n6571) );
  INV_X1 U9040 ( .A(n13904), .ZN(n7355) );
  NAND2_X1 U9041 ( .A1(n7502), .A2(n7493), .ZN(n13312) );
  INV_X1 U9042 ( .A(n13312), .ZN(n6689) );
  OR2_X1 U9043 ( .A1(n9609), .A2(n14279), .ZN(n9687) );
  INV_X1 U9044 ( .A(n9687), .ZN(n7289) );
  OR2_X1 U9045 ( .A1(n6740), .A2(n6977), .ZN(n6572) );
  NAND2_X1 U9046 ( .A1(n11504), .A2(n11503), .ZN(n14205) );
  INV_X1 U9047 ( .A(n14205), .ZN(n6952) );
  AND2_X2 U9048 ( .A1(n8770), .A2(n10263), .ZN(n14880) );
  AND2_X1 U9049 ( .A1(n14883), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6573) );
  AND2_X2 U9050 ( .A1(n8770), .A2(n7514), .ZN(n14885) );
  OR2_X1 U9051 ( .A1(n15052), .A2(n8750), .ZN(n6574) );
  OR2_X1 U9052 ( .A1(n14768), .A2(n10743), .ZN(n14531) );
  INV_X1 U9053 ( .A(n14531), .ZN(n7384) );
  NOR2_X1 U9054 ( .A1(n12522), .A2(n12521), .ZN(n6575) );
  AND2_X1 U9055 ( .A1(n10505), .A2(n7109), .ZN(n6576) );
  AND2_X1 U9056 ( .A1(n8958), .A2(n7344), .ZN(n6577) );
  OR2_X1 U9057 ( .A1(n15052), .A2(n9104), .ZN(n6578) );
  AND2_X1 U9058 ( .A1(n11665), .A2(n11370), .ZN(n14574) );
  NAND2_X1 U9059 ( .A1(n6687), .A2(n6688), .ZN(n8915) );
  NAND4_X1 U9060 ( .A1(n8211), .A2(n8210), .A3(n8209), .A4(n8208), .ZN(n10042)
         );
  INV_X1 U9061 ( .A(n13104), .ZN(n6910) );
  XNOR2_X1 U9062 ( .A(n7489), .B(n15080), .ZN(n11882) );
  AND2_X2 U9063 ( .A1(n10057), .A2(n8764), .ZN(n15066) );
  INV_X2 U9064 ( .A(n15050), .ZN(n15052) );
  NAND2_X1 U9065 ( .A1(n12612), .A2(n10032), .ZN(n12474) );
  INV_X1 U9066 ( .A(n7147), .ZN(n6780) );
  AND2_X1 U9067 ( .A1(n8817), .A2(n12861), .ZN(n6579) );
  NAND2_X1 U9068 ( .A1(n11902), .A2(n10592), .ZN(n10593) );
  INV_X1 U9069 ( .A(n10593), .ZN(n6913) );
  NOR2_X1 U9070 ( .A1(n14926), .A2(n10205), .ZN(n6580) );
  AND2_X1 U9071 ( .A1(n11390), .A2(n11391), .ZN(n6581) );
  INV_X1 U9072 ( .A(n14945), .ZN(n14987) );
  AND2_X1 U9073 ( .A1(P3_U3897), .A2(n8664), .ZN(n14945) );
  OR2_X1 U9074 ( .A1(n12595), .A2(n12575), .ZN(n6582) );
  OR2_X1 U9075 ( .A1(n12582), .A2(n12784), .ZN(n6583) );
  AND2_X1 U9076 ( .A1(n8712), .A2(n6936), .ZN(n12984) );
  NAND2_X1 U9077 ( .A1(n7289), .A2(n7288), .ZN(n14419) );
  NAND2_X1 U9078 ( .A1(n11960), .A2(n11959), .ZN(n11963) );
  NAND2_X1 U9079 ( .A1(n12027), .A2(n12026), .ZN(n12036) );
  INV_X1 U9080 ( .A(n12084), .ZN(n12092) );
  AOI21_X1 U9081 ( .B1(n7247), .B2(n7250), .A(n7246), .ZN(n7245) );
  XNOR2_X1 U9082 ( .A(n11926), .B(n6584), .ZN(n7218) );
  NAND2_X1 U9083 ( .A1(n10235), .A2(n12102), .ZN(n7074) );
  OAI21_X2 U9084 ( .B1(n13385), .B2(n8136), .A(n8135), .ZN(n13367) );
  NAND2_X1 U9085 ( .A1(n13422), .A2(n8130), .ZN(n13412) );
  NAND2_X1 U9086 ( .A1(n8106), .A2(n12096), .ZN(n9832) );
  OAI21_X1 U9087 ( .B1(n13351), .B2(n13337), .A(n8142), .ZN(n8144) );
  NAND2_X1 U9088 ( .A1(n10895), .A2(n12107), .ZN(n10894) );
  NAND2_X1 U9089 ( .A1(n7092), .A2(n7094), .ZN(n13278) );
  NAND2_X1 U9090 ( .A1(n6886), .A2(n6884), .ZN(n10536) );
  NOR2_X1 U9091 ( .A1(n11001), .A2(n11003), .ZN(n11065) );
  NAND2_X1 U9092 ( .A1(n14958), .A2(n7162), .ZN(n7159) );
  NOR2_X1 U9093 ( .A1(n10728), .A2(n15062), .ZN(n10995) );
  NAND2_X1 U9094 ( .A1(n6897), .A2(n14896), .ZN(n6896) );
  OAI21_X1 U9095 ( .B1(P3_IR_REG_31__SCAN_IN), .B2(P3_IR_REG_1__SCAN_IN), .A(
        n7144), .ZN(n7143) );
  XNOR2_X2 U9096 ( .A(n7639), .B(n13649), .ZN(n7644) );
  NAND3_X1 U9097 ( .A1(n6586), .A2(n6585), .A3(n7219), .ZN(n6600) );
  NAND2_X1 U9098 ( .A1(n11998), .A2(n11997), .ZN(n6585) );
  NAND2_X1 U9099 ( .A1(n6590), .A2(n11994), .ZN(n6586) );
  NAND2_X2 U9100 ( .A1(n6613), .A2(n7658), .ZN(n11881) );
  OAI21_X2 U9101 ( .B1(n13324), .B2(n7089), .A(n7086), .ZN(n13290) );
  NAND2_X2 U9102 ( .A1(n7998), .A2(n7997), .ZN(n13324) );
  XNOR2_X2 U9103 ( .A(n11885), .B(n8917), .ZN(n12096) );
  NAND2_X2 U9104 ( .A1(n7665), .A2(n6588), .ZN(n8917) );
  OR2_X1 U9105 ( .A1(n7678), .A2(n9526), .ZN(n7655) );
  XNOR2_X2 U9106 ( .A(n13146), .B(n11890), .ZN(n12095) );
  NAND2_X1 U9107 ( .A1(n11884), .A2(n7218), .ZN(n11889) );
  NAND2_X1 U9108 ( .A1(n7244), .A2(n7245), .ZN(n11929) );
  NAND2_X1 U9109 ( .A1(n11995), .A2(n11996), .ZN(n6590) );
  NAND3_X1 U9110 ( .A1(n12319), .A2(n12472), .A3(n6592), .ZN(n6591) );
  NAND2_X1 U9111 ( .A1(n8441), .A2(n8440), .ZN(n8455) );
  INV_X1 U9112 ( .A(n12290), .ZN(n12931) );
  OAI211_X1 U9113 ( .C1(n12476), .C2(n12477), .A(n6594), .B(n6593), .ZN(n12478) );
  OR2_X1 U9114 ( .A1(n12473), .A2(n12475), .ZN(n6593) );
  NAND2_X1 U9115 ( .A1(n12473), .A2(n8652), .ZN(n6594) );
  NAND2_X1 U9116 ( .A1(n12279), .A2(n12278), .ZN(n12290) );
  XNOR2_X1 U9117 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8233) );
  NAND2_X1 U9118 ( .A1(n8309), .A2(n8308), .ZN(n8327) );
  NAND2_X1 U9119 ( .A1(n9088), .A2(n9087), .ZN(n9090) );
  OAI21_X1 U9120 ( .B1(n9106), .B2(n15050), .A(n6817), .ZN(P3_U3456) );
  OAI21_X1 U9121 ( .B1(n9106), .B2(n15064), .A(n7032), .ZN(P3_U3488) );
  NAND2_X1 U9122 ( .A1(n11060), .A2(n7178), .ZN(n14566) );
  NAND2_X1 U9123 ( .A1(n13972), .A2(n13971), .ZN(n13970) );
  INV_X1 U9124 ( .A(n13944), .ZN(n13891) );
  NAND2_X1 U9125 ( .A1(n10330), .A2(n10329), .ZN(n10471) );
  INV_X1 U9126 ( .A(n14085), .ZN(n6599) );
  NAND2_X2 U9127 ( .A1(n9306), .A2(n9307), .ZN(n11545) );
  NAND2_X1 U9128 ( .A1(n9730), .A2(n11677), .ZN(n9855) );
  NOR2_X1 U9129 ( .A1(n11679), .A2(n6597), .ZN(n6596) );
  NAND2_X2 U9130 ( .A1(n10141), .A2(n9862), .ZN(n9893) );
  NAND2_X1 U9131 ( .A1(n9779), .A2(n11675), .ZN(n9781) );
  NAND2_X1 U9132 ( .A1(n14432), .A2(n14433), .ZN(n11060) );
  NAND2_X1 U9133 ( .A1(n11295), .A2(n11301), .ZN(n7193) );
  NAND2_X2 U9134 ( .A1(n7437), .A2(n14058), .ZN(n14057) );
  NAND2_X1 U9135 ( .A1(n6600), .A2(n6642), .ZN(n12003) );
  BUF_X1 U9136 ( .A(n6441), .Z(n6601) );
  NAND2_X1 U9137 ( .A1(n10018), .A2(n12098), .ZN(n10017) );
  NAND2_X1 U9138 ( .A1(n10428), .A2(n10433), .ZN(n10427) );
  NAND2_X1 U9139 ( .A1(n13420), .A2(n13419), .ZN(n13418) );
  OR2_X2 U9140 ( .A1(n10266), .A2(n12096), .ZN(n9831) );
  NAND3_X1 U9141 ( .A1(n6602), .A2(n6869), .A3(n6865), .ZN(n14444) );
  NAND3_X1 U9142 ( .A1(n6870), .A2(n6875), .A3(n14445), .ZN(n6602) );
  NAND2_X1 U9143 ( .A1(n14395), .A2(n14394), .ZN(n7211) );
  NAND2_X1 U9144 ( .A1(n7206), .A2(n7205), .ZN(n7204) );
  NOR2_X1 U9145 ( .A1(n14331), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n14287) );
  XNOR2_X1 U9146 ( .A(n7208), .B(n6516), .ZN(SUB_1596_U4) );
  OAI22_X1 U9147 ( .A1(n14335), .A2(n14281), .B1(P1_ADDR_REG_1__SCAN_IN), .B2(
        n7214), .ZN(n7213) );
  NAND2_X1 U9148 ( .A1(n8439), .A2(n8438), .ZN(n8441) );
  NAND2_X1 U9149 ( .A1(n12029), .A2(n7228), .ZN(n6632) );
  NAND2_X1 U9150 ( .A1(n8195), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8221) );
  NAND3_X1 U9151 ( .A1(n8903), .A2(n9088), .A3(n12837), .ZN(n6604) );
  NAND2_X1 U9152 ( .A1(n6607), .A2(n6605), .ZN(P3_U3487) );
  OR2_X1 U9153 ( .A1(n8913), .A2(n15064), .ZN(n6607) );
  AOI21_X1 U9154 ( .B1(n13955), .B2(n13954), .A(n6456), .ZN(n13926) );
  NAND2_X1 U9155 ( .A1(n11025), .A2(n11024), .ZN(n14431) );
  NAND2_X1 U9156 ( .A1(n13896), .A2(n13895), .ZN(n14100) );
  NAND2_X1 U9157 ( .A1(n7391), .A2(n7558), .ZN(n7815) );
  NAND2_X4 U9158 ( .A1(n8664), .A2(n8663), .ZN(n9753) );
  NAND2_X1 U9159 ( .A1(n6732), .A2(n7552), .ZN(n7783) );
  NAND2_X1 U9160 ( .A1(n13976), .A2(n13905), .ZN(n13959) );
  NAND2_X1 U9161 ( .A1(n12802), .A2(n8684), .ZN(n12791) );
  NAND2_X1 U9162 ( .A1(n12717), .A2(n8696), .ZN(n6701) );
  OAI21_X1 U9163 ( .B1(n7385), .B2(n7384), .A(n14532), .ZN(n7383) );
  NAND2_X1 U9164 ( .A1(n6645), .A2(n6632), .ZN(n12084) );
  NAND2_X1 U9165 ( .A1(n11907), .A2(n11906), .ZN(n11913) );
  NAND2_X1 U9166 ( .A1(n11952), .A2(n11951), .ZN(n11955) );
  NAND2_X1 U9167 ( .A1(n12019), .A2(n12018), .ZN(n12022) );
  NAND2_X1 U9168 ( .A1(n11913), .A2(n11912), .ZN(n11910) );
  AND2_X2 U9169 ( .A1(n7670), .A2(n7683), .ZN(n7460) );
  OR2_X1 U9170 ( .A1(n13511), .A2(n6615), .ZN(P2_U3527) );
  NAND2_X1 U9171 ( .A1(n10232), .A2(n10234), .ZN(n10231) );
  NAND2_X1 U9172 ( .A1(n13231), .A2(n13230), .ZN(n13508) );
  NAND2_X1 U9173 ( .A1(n6616), .A2(n11886), .ZN(n11887) );
  NAND2_X1 U9174 ( .A1(n11889), .A2(n11888), .ZN(n6616) );
  INV_X1 U9175 ( .A(n14985), .ZN(n6624) );
  NOR2_X1 U9176 ( .A1(n12570), .A2(n12569), .ZN(n12584) );
  INV_X1 U9177 ( .A(n11013), .ZN(n6622) );
  NOR2_X1 U9178 ( .A1(n14965), .A2(n14966), .ZN(n14964) );
  OAI22_X1 U9179 ( .A1(n10192), .A2(n10191), .B1(n10190), .B2(n10202), .ZN(
        n14921) );
  XNOR2_X1 U9180 ( .A(n12608), .B(n6620), .ZN(n12618) );
  OAI22_X1 U9181 ( .A1(n9919), .A2(n9918), .B1(n9917), .B2(n9916), .ZN(n14905)
         );
  AND2_X2 U9182 ( .A1(n14566), .A2(n11178), .ZN(n11180) );
  AND2_X1 U9183 ( .A1(n6896), .A2(n6895), .ZN(n6894) );
  INV_X1 U9184 ( .A(n6710), .ZN(n8640) );
  AND2_X2 U9185 ( .A1(n11395), .A2(n11396), .ZN(n11404) );
  AOI21_X2 U9186 ( .B1(n14072), .B2(n14078), .A(n6566), .ZN(n7437) );
  NAND2_X1 U9187 ( .A1(n10581), .A2(n7718), .ZN(n10428) );
  NAND2_X1 U9188 ( .A1(n13229), .A2(n13228), .ZN(n13231) );
  INV_X1 U9189 ( .A(n12096), .ZN(n6638) );
  NAND2_X1 U9190 ( .A1(n10889), .A2(n8121), .ZN(n7118) );
  NAND2_X1 U9191 ( .A1(n7118), .A2(n7116), .ZN(n7112) );
  NAND2_X1 U9192 ( .A1(n7101), .A2(n7098), .ZN(n7097) );
  INV_X1 U9193 ( .A(n6970), .ZN(n6969) );
  AOI21_X2 U9194 ( .B1(n13243), .B2(n13258), .A(n8154), .ZN(n13234) );
  AND2_X2 U9195 ( .A1(n7627), .A2(n6540), .ZN(n7640) );
  NAND2_X2 U9196 ( .A1(n8144), .A2(n8143), .ZN(n13319) );
  OAI21_X1 U9197 ( .B1(n11898), .B2(n7080), .A(n8111), .ZN(n7079) );
  INV_X1 U9198 ( .A(n7079), .ZN(n7078) );
  NAND2_X1 U9199 ( .A1(n10738), .A2(n10737), .ZN(n10859) );
  NAND2_X1 U9200 ( .A1(n11291), .A2(n11290), .ZN(n11295) );
  NAND2_X1 U9201 ( .A1(n9733), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9630) );
  NAND2_X1 U9202 ( .A1(n7348), .A2(n7346), .ZN(n13976) );
  NAND2_X1 U9203 ( .A1(n7371), .A2(n6454), .ZN(n7370) );
  NAND2_X1 U9204 ( .A1(n6439), .A2(n6630), .ZN(n14033) );
  XNOR2_X1 U9205 ( .A(n13894), .B(n13908), .ZN(n14128) );
  INV_X1 U9206 ( .A(n7383), .ZN(n7382) );
  INV_X1 U9207 ( .A(n6945), .ZN(n6774) );
  INV_X1 U9208 ( .A(n9911), .ZN(n6631) );
  NAND2_X1 U9209 ( .A1(n14137), .A2(n6629), .ZN(n14236) );
  NAND2_X1 U9210 ( .A1(n14536), .A2(n10830), .ZN(n10842) );
  NAND2_X2 U9211 ( .A1(n14531), .A2(n10744), .ZN(n11684) );
  NAND2_X1 U9212 ( .A1(n12092), .A2(n12091), .ZN(n6633) );
  NAND2_X1 U9213 ( .A1(n6633), .A2(n6533), .ZN(n12136) );
  INV_X1 U9214 ( .A(n14441), .ZN(n6868) );
  INV_X1 U9215 ( .A(n7213), .ZN(n14334) );
  XNOR2_X2 U9216 ( .A(n14285), .B(n14286), .ZN(n14331) );
  OAI21_X1 U9217 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(n15241), .A(n6536), .ZN(
        n6859) );
  NAND2_X1 U9218 ( .A1(n15240), .A2(n15239), .ZN(n7198) );
  XNOR2_X1 U9219 ( .A(n14335), .B(n14281), .ZN(n14338) );
  OR2_X2 U9220 ( .A1(n11158), .A2(n14493), .ZN(n7851) );
  NAND2_X1 U9221 ( .A1(n11112), .A2(n12304), .ZN(n6954) );
  NAND2_X1 U9222 ( .A1(n6700), .A2(n6543), .ZN(n6698) );
  NAND2_X1 U9223 ( .A1(n10770), .A2(n10768), .ZN(n6935) );
  NOR2_X1 U9224 ( .A1(n8700), .A2(n6647), .ZN(n12664) );
  NAND2_X1 U9225 ( .A1(n8169), .A2(n6652), .ZN(P2_U3528) );
  NAND2_X1 U9226 ( .A1(n14040), .A2(n14053), .ZN(n14039) );
  NAND2_X1 U9227 ( .A1(n7783), .A2(n7553), .ZN(n6972) );
  OAI21_X1 U9228 ( .B1(n14146), .B2(n14755), .A(n6539), .ZN(n14237) );
  NAND2_X1 U9229 ( .A1(n7370), .A2(n7369), .ZN(n13896) );
  NAND3_X1 U9230 ( .A1(n6641), .A2(n6640), .A3(n6548), .ZN(n7242) );
  NAND2_X1 U9231 ( .A1(n11940), .A2(n11939), .ZN(n6640) );
  NAND2_X1 U9232 ( .A1(n11936), .A2(n11935), .ZN(n6641) );
  NAND2_X1 U9233 ( .A1(n7240), .A2(n7239), .ZN(n11995) );
  NAND2_X1 U9234 ( .A1(n7222), .A2(n7221), .ZN(n11974) );
  NAND2_X1 U9235 ( .A1(n7234), .A2(n7233), .ZN(n12014) );
  NAND2_X1 U9236 ( .A1(n7237), .A2(n7236), .ZN(n11985) );
  NAND2_X1 U9237 ( .A1(n7476), .A2(n7345), .ZN(n6920) );
  NAND2_X1 U9238 ( .A1(n8424), .A2(n8423), .ZN(n8439) );
  INV_X1 U9239 ( .A(n8585), .ZN(n7036) );
  NAND2_X1 U9240 ( .A1(n8379), .A2(n8378), .ZN(n8390) );
  NAND2_X1 U9241 ( .A1(n8363), .A2(n8362), .ZN(n8376) );
  NAND2_X1 U9242 ( .A1(n8235), .A2(n7006), .ZN(n7005) );
  OAI21_X2 U9243 ( .B1(n8895), .B2(n8894), .A(n8896), .ZN(n9080) );
  NOR2_X1 U9244 ( .A1(n14619), .A2(n7440), .ZN(n10367) );
  XNOR2_X1 U9245 ( .A(n6643), .B(n11217), .ZN(n10163) );
  NAND2_X1 U9246 ( .A1(n9800), .A2(n9801), .ZN(n6643) );
  OR2_X2 U9247 ( .A1(n11254), .A2(n11253), .ZN(n11255) );
  NAND2_X1 U9248 ( .A1(n13777), .A2(n13776), .ZN(n7282) );
  OAI21_X2 U9249 ( .B1(n10702), .B2(n7285), .A(n7283), .ZN(n11251) );
  NAND3_X1 U9250 ( .A1(n10370), .A2(n10371), .A3(n7297), .ZN(n7296) );
  AND3_X1 U9251 ( .A1(n7373), .A2(n6943), .A3(n6774), .ZN(n6944) );
  INV_X1 U9252 ( .A(n6646), .ZN(n6645) );
  NAND2_X1 U9253 ( .A1(n7177), .A2(n10103), .ZN(n10322) );
  NAND3_X1 U9254 ( .A1(n7034), .A2(n8423), .A3(P1_DATAO_REG_13__SCAN_IN), .ZN(
        n8424) );
  NAND2_X1 U9255 ( .A1(n8307), .A2(n8306), .ZN(n8309) );
  NAND2_X1 U9256 ( .A1(n8361), .A2(n8360), .ZN(n8363) );
  NAND2_X1 U9257 ( .A1(n8376), .A2(n8375), .ZN(n8379) );
  NAND2_X1 U9258 ( .A1(n8257), .A2(n8256), .ZN(n8277) );
  NAND2_X1 U9259 ( .A1(n13237), .A2(n13236), .ZN(n6649) );
  NAND2_X2 U9260 ( .A1(n6962), .A2(n6963), .ZN(n7766) );
  OAI21_X1 U9261 ( .B1(n12619), .B2(n14995), .A(n6894), .ZN(P3_U3201) );
  NOR2_X1 U9262 ( .A1(n14964), .A2(n11012), .ZN(n11013) );
  AOI21_X1 U9263 ( .B1(n12618), .B2(n14945), .A(n12617), .ZN(n6895) );
  NAND2_X1 U9264 ( .A1(n7112), .A2(n7827), .ZN(n11158) );
  INV_X1 U9265 ( .A(n9031), .ZN(n6655) );
  NAND2_X1 U9266 ( .A1(n9029), .A2(n9030), .ZN(n9031) );
  NAND2_X1 U9267 ( .A1(n6658), .A2(n6656), .ZN(n13037) );
  NAND2_X1 U9268 ( .A1(n6657), .A2(n6660), .ZN(n6656) );
  OR2_X1 U9269 ( .A1(n8983), .A2(n6664), .ZN(n6657) );
  NAND2_X1 U9270 ( .A1(n6665), .A2(n6659), .ZN(n6658) );
  NAND2_X1 U9271 ( .A1(n8983), .A2(n8982), .ZN(n6665) );
  INV_X1 U9272 ( .A(n8982), .ZN(n6662) );
  NAND2_X1 U9273 ( .A1(n7343), .A2(n6667), .ZN(n6666) );
  NAND2_X1 U9274 ( .A1(n10384), .A2(n6680), .ZN(n6679) );
  NAND3_X1 U9275 ( .A1(n6679), .A2(n6678), .A3(n8970), .ZN(n10819) );
  OAI21_X2 U9276 ( .B1(n11882), .B2(n6689), .A(n6595), .ZN(n8928) );
  INV_X1 U9277 ( .A(n11882), .ZN(n8102) );
  NAND2_X1 U9278 ( .A1(n7837), .A2(n6690), .ZN(n7493) );
  NAND2_X1 U9279 ( .A1(n7837), .A2(n6551), .ZN(n7490) );
  NAND2_X4 U9280 ( .A1(n9753), .A2(n11542), .ZN(n8258) );
  NAND2_X1 U9281 ( .A1(n8682), .A2(n6455), .ZN(n6691) );
  NAND2_X1 U9282 ( .A1(n6691), .A2(n6692), .ZN(n12819) );
  NOR2_X2 U9283 ( .A1(n8642), .A2(n7061), .ZN(n6700) );
  NAND2_X1 U9284 ( .A1(n12791), .A2(n6706), .ZN(n6702) );
  NAND2_X1 U9285 ( .A1(n6702), .A2(n6703), .ZN(n12765) );
  NAND4_X1 U9286 ( .A1(n7430), .A2(n7432), .A3(n8173), .A4(n6829), .ZN(n6710)
         );
  AND2_X2 U9287 ( .A1(n9761), .A2(n8171), .ZN(n8173) );
  AND2_X2 U9288 ( .A1(n8396), .A2(n6538), .ZN(n7432) );
  AND2_X2 U9289 ( .A1(n8178), .A2(n7431), .ZN(n7430) );
  NAND2_X1 U9290 ( .A1(n10558), .A2(n8672), .ZN(n10687) );
  INV_X1 U9291 ( .A(n6716), .ZN(n12298) );
  OAI21_X2 U9292 ( .B1(n7686), .B2(n7685), .A(n7528), .ZN(n6723) );
  NAND2_X1 U9293 ( .A1(n6723), .A2(n7533), .ZN(n7536) );
  XNOR2_X1 U9294 ( .A(n6723), .B(n7700), .ZN(n9857) );
  NAND2_X1 U9295 ( .A1(n7766), .A2(n7550), .ZN(n6732) );
  NAND2_X1 U9296 ( .A1(n7830), .A2(n7829), .ZN(n7832) );
  NAND2_X1 U9297 ( .A1(n7585), .A2(n6569), .ZN(n6735) );
  AND2_X1 U9298 ( .A1(n6735), .A2(n6733), .ZN(n7586) );
  NAND2_X1 U9299 ( .A1(n8032), .A2(n7614), .ZN(n8045) );
  NAND2_X1 U9300 ( .A1(n6744), .A2(n6745), .ZN(n7607) );
  NAND2_X1 U9301 ( .A1(n7593), .A2(n6450), .ZN(n6744) );
  NAND2_X1 U9302 ( .A1(n7593), .A2(n6975), .ZN(n6751) );
  NAND3_X1 U9303 ( .A1(n11456), .A2(n6761), .A3(n6571), .ZN(n6760) );
  NAND4_X1 U9304 ( .A1(n11640), .A2(n6461), .A3(n11639), .A4(n6765), .ZN(n6763) );
  NAND4_X1 U9305 ( .A1(n11466), .A2(n11465), .A3(n6770), .A4(n6980), .ZN(n6769) );
  NAND2_X1 U9306 ( .A1(n6769), .A2(n6767), .ZN(n11513) );
  NAND2_X1 U9307 ( .A1(n6780), .A2(n6784), .ZN(n6782) );
  AND2_X1 U9308 ( .A1(n10537), .A2(n7146), .ZN(n6785) );
  XNOR2_X1 U9309 ( .A(n12535), .B(n12553), .ZN(n6789) );
  NAND2_X1 U9310 ( .A1(n6789), .A2(n6472), .ZN(n6788) );
  OAI21_X1 U9311 ( .B1(n6496), .B2(n12537), .A(n6788), .ZN(n12564) );
  INV_X1 U9312 ( .A(n6790), .ZN(n14975) );
  NAND2_X1 U9313 ( .A1(n7149), .A2(n7148), .ZN(n12534) );
  XNOR2_X1 U9314 ( .A(n12510), .B(n12511), .ZN(n14976) );
  INV_X1 U9315 ( .A(n10521), .ZN(n6793) );
  NAND2_X1 U9316 ( .A1(n10903), .A2(n6800), .ZN(n6796) );
  NAND2_X1 U9317 ( .A1(n6796), .A2(n6797), .ZN(n10931) );
  NAND2_X1 U9318 ( .A1(n12836), .A2(n6806), .ZN(n6803) );
  NAND2_X1 U9319 ( .A1(n6803), .A2(n6804), .ZN(n12809) );
  OAI21_X1 U9320 ( .B1(n8331), .B2(n6814), .A(n6811), .ZN(n12854) );
  NAND2_X1 U9321 ( .A1(n6815), .A2(n12340), .ZN(n10557) );
  NAND2_X1 U9322 ( .A1(n6816), .A2(n12331), .ZN(n10300) );
  NAND2_X1 U9323 ( .A1(n12671), .A2(n6462), .ZN(n6821) );
  NAND2_X1 U9324 ( .A1(n12671), .A2(n6825), .ZN(n6822) );
  NAND2_X1 U9325 ( .A1(n12671), .A2(n12445), .ZN(n12654) );
  NAND3_X1 U9326 ( .A1(n7432), .A2(n7430), .A3(n8173), .ZN(n8646) );
  NAND3_X1 U9327 ( .A1(n8851), .A2(n12212), .A3(n12719), .ZN(n12168) );
  NAND2_X2 U9328 ( .A1(n6832), .A2(n12213), .ZN(n9139) );
  XNOR2_X2 U9329 ( .A(n6840), .B(n8514), .ZN(n12612) );
  NAND2_X1 U9330 ( .A1(n11338), .A2(n6848), .ZN(n6845) );
  NAND2_X1 U9331 ( .A1(n6845), .A2(n6846), .ZN(n7412) );
  OAI21_X1 U9332 ( .B1(n11338), .B2(n8816), .A(n6856), .ZN(n12233) );
  AND2_X1 U9333 ( .A1(n14372), .A2(n6857), .ZN(n14601) );
  NAND2_X1 U9334 ( .A1(n14600), .A2(n14599), .ZN(n6857) );
  INV_X1 U9335 ( .A(n7207), .ZN(n14603) );
  NAND2_X1 U9336 ( .A1(n14377), .A2(n14376), .ZN(n7207) );
  XNOR2_X2 U9337 ( .A(n6864), .B(P3_ADDR_REG_3__SCAN_IN), .ZN(n14342) );
  NAND2_X1 U9338 ( .A1(n6868), .A2(n6871), .ZN(n6875) );
  NAND2_X1 U9339 ( .A1(n14386), .A2(n6866), .ZN(n6865) );
  NAND2_X1 U9340 ( .A1(n14386), .A2(n14442), .ZN(n6870) );
  NAND2_X1 U9341 ( .A1(n6868), .A2(n6867), .ZN(n6869) );
  NAND2_X1 U9342 ( .A1(n6870), .A2(n6875), .ZN(n6874) );
  INV_X1 U9343 ( .A(n6875), .ZN(n14439) );
  INV_X1 U9344 ( .A(n14440), .ZN(n6871) );
  NAND2_X1 U9345 ( .A1(n6874), .A2(n6873), .ZN(n6872) );
  NAND2_X1 U9346 ( .A1(n14927), .A2(n6885), .ZN(n6884) );
  INV_X1 U9347 ( .A(n10205), .ZN(n6885) );
  OAI21_X1 U9348 ( .B1(n10205), .B2(P3_REG1_REG_5__SCAN_IN), .A(n10206), .ZN(
        n6887) );
  NOR2_X1 U9349 ( .A1(n14927), .A2(n8268), .ZN(n14926) );
  NAND2_X1 U9350 ( .A1(n6893), .A2(n6473), .ZN(n6891) );
  INV_X1 U9351 ( .A(n14459), .ZN(n6893) );
  MUX2_X1 U9352 ( .A(n9774), .B(n10254), .S(n9773), .Z(n6902) );
  NAND2_X1 U9353 ( .A1(n8640), .A2(n6904), .ZN(n8722) );
  NAND2_X1 U9354 ( .A1(n8640), .A2(n8180), .ZN(n8642) );
  OAI21_X1 U9355 ( .B1(n12598), .B2(n14995), .A(n6504), .ZN(P3_U3200) );
  AND2_X1 U9356 ( .A1(n6908), .A2(n6907), .ZN(n6906) );
  AOI21_X1 U9357 ( .B1(n14944), .B2(n12606), .A(n12589), .ZN(n6907) );
  OAI21_X1 U9358 ( .B1(n12605), .B2(n6909), .A(n14945), .ZN(n6908) );
  INV_X1 U9359 ( .A(n6919), .ZN(n13342) );
  NAND2_X1 U9360 ( .A1(n13261), .A2(n6921), .ZN(n13221) );
  NAND2_X1 U9361 ( .A1(n11167), .A2(n6924), .ZN(n13450) );
  INV_X1 U9362 ( .A(n6929), .ZN(n13449) );
  NOR2_X2 U9363 ( .A1(n6932), .A2(n14768), .ZN(n14542) );
  NAND2_X1 U9364 ( .A1(n6935), .A2(n6933), .ZN(n10948) );
  NAND2_X1 U9365 ( .A1(n8712), .A2(n6464), .ZN(n8183) );
  INV_X1 U9366 ( .A(n6942), .ZN(n13982) );
  NAND3_X1 U9367 ( .A1(n9174), .A2(n9245), .A3(n9173), .ZN(n9185) );
  NOR2_X1 U9368 ( .A1(n9162), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n6943) );
  AND3_X2 U9369 ( .A1(n6944), .A2(n9165), .A3(n7444), .ZN(n9251) );
  NAND4_X1 U9370 ( .A1(n9158), .A2(n9157), .A3(n9288), .A4(n9260), .ZN(n6945)
         );
  AND2_X2 U9371 ( .A1(n9871), .A2(n9870), .ZN(n11409) );
  NOR2_X2 U9372 ( .A1(n14541), .A2(n13712), .ZN(n6948) );
  NAND2_X1 U9373 ( .A1(n11306), .A2(n6949), .ZN(n14065) );
  OAI21_X1 U9374 ( .B1(n8765), .B2(n15064), .A(n6570), .ZN(P3_U3486) );
  NAND2_X2 U9375 ( .A1(n12664), .A2(n8705), .ZN(n7031) );
  XNOR2_X2 U9376 ( .A(n7527), .B(SI_2_), .ZN(n7686) );
  NAND2_X2 U9377 ( .A1(n7526), .A2(n7525), .ZN(n7527) );
  NAND3_X1 U9378 ( .A1(n7595), .A2(n7594), .A3(n7396), .ZN(n7967) );
  NAND2_X1 U9379 ( .A1(n11419), .A2(n6986), .ZN(n6985) );
  NAND3_X1 U9380 ( .A1(n6985), .A2(n6984), .A3(n11425), .ZN(n11424) );
  OAI21_X1 U9381 ( .B1(n11450), .B2(n6994), .A(n6992), .ZN(n11454) );
  NAND2_X1 U9382 ( .A1(n6991), .A2(n6989), .ZN(n11453) );
  NAND2_X1 U9383 ( .A1(n11450), .A2(n6992), .ZN(n6991) );
  OAI21_X1 U9384 ( .B1(n11623), .B2(n6996), .A(n6995), .ZN(n11637) );
  NAND2_X1 U9385 ( .A1(n6997), .A2(n6998), .ZN(n7407) );
  NAND3_X1 U9386 ( .A1(n11561), .A2(n11560), .A3(n6546), .ZN(n6997) );
  OAI22_X1 U9387 ( .A1(n11437), .A2(n7002), .B1(n11438), .B2(n7001), .ZN(
        n11443) );
  NAND2_X1 U9388 ( .A1(n11443), .A2(n11444), .ZN(n11442) );
  OAI22_X1 U9389 ( .A1(n11539), .A2(n7004), .B1(n11540), .B2(n7003), .ZN(
        n11556) );
  INV_X1 U9390 ( .A(n11556), .ZN(n11559) );
  INV_X1 U9391 ( .A(n11461), .ZN(n11464) );
  NAND2_X1 U9392 ( .A1(n8225), .A2(n6506), .ZN(n7007) );
  INV_X1 U9393 ( .A(n8233), .ZN(n7006) );
  NAND3_X1 U9394 ( .A1(n7007), .A2(n7005), .A3(n8254), .ZN(n8257) );
  NAND2_X1 U9395 ( .A1(n7008), .A2(n8235), .ZN(n8255) );
  NAND2_X1 U9396 ( .A1(n8234), .A2(n8233), .ZN(n7008) );
  NAND2_X1 U9397 ( .A1(n8455), .A2(n7019), .ZN(n7017) );
  AOI21_X1 U9398 ( .B1(n8630), .B2(n8629), .A(n12489), .ZN(n7023) );
  NOR2_X1 U9399 ( .A1(n12461), .A2(n7030), .ZN(n7029) );
  NAND3_X1 U9400 ( .A1(n6507), .A2(n7031), .A3(n8901), .ZN(n8902) );
  OAI21_X2 U9401 ( .B1(n8571), .B2(n8570), .A(n8572), .ZN(n8581) );
  OAI21_X2 U9402 ( .B1(n8390), .B2(n8389), .A(n8391), .ZN(n8394) );
  NAND2_X1 U9403 ( .A1(n7035), .A2(n8585), .ZN(n8597) );
  NAND2_X1 U9404 ( .A1(n10657), .A2(n12346), .ZN(n7037) );
  NAND2_X1 U9405 ( .A1(n8262), .A2(n8261), .ZN(n10657) );
  NAND2_X1 U9406 ( .A1(n8331), .A2(n12372), .ZN(n10946) );
  INV_X1 U9407 ( .A(n12372), .ZN(n7054) );
  NAND2_X1 U9408 ( .A1(n12654), .A2(n12450), .ZN(n7055) );
  NAND2_X1 U9409 ( .A1(n12708), .A2(n12707), .ZN(n12709) );
  NAND2_X1 U9410 ( .A1(n8556), .A2(n12433), .ZN(n12721) );
  NAND2_X1 U9411 ( .A1(n8243), .A2(n12342), .ZN(n10685) );
  NAND2_X1 U9412 ( .A1(n12808), .A2(n12405), .ZN(n12799) );
  XNOR2_X1 U9413 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n8223) );
  NAND2_X2 U9414 ( .A1(n8158), .A2(n13658), .ZN(n7662) );
  INV_X1 U9415 ( .A(n10501), .ZN(n7067) );
  NAND2_X1 U9416 ( .A1(n7063), .A2(n7064), .ZN(n7798) );
  NAND2_X1 U9417 ( .A1(n10501), .A2(n7781), .ZN(n7063) );
  NAND2_X1 U9418 ( .A1(n7460), .A2(n7068), .ZN(n7069) );
  NOR2_X2 U9419 ( .A1(n7698), .A2(n7071), .ZN(n7475) );
  NAND2_X1 U9420 ( .A1(n7074), .A2(n7072), .ZN(n8117) );
  NAND2_X1 U9421 ( .A1(n7078), .A2(n7075), .ZN(n8113) );
  NAND2_X1 U9422 ( .A1(n10019), .A2(n7076), .ZN(n7075) );
  NAND2_X1 U9423 ( .A1(n7081), .A2(n7082), .ZN(n7963) );
  NAND2_X1 U9424 ( .A1(n13379), .A2(n7945), .ZN(n7081) );
  NAND2_X1 U9425 ( .A1(n13319), .A2(n7096), .ZN(n7094) );
  NAND2_X1 U9426 ( .A1(n13319), .A2(n8146), .ZN(n7095) );
  NAND2_X1 U9427 ( .A1(n13256), .A2(n8072), .ZN(n13229) );
  NAND2_X2 U9428 ( .A1(n8071), .A2(n7104), .ZN(n13256) );
  NAND2_X1 U9429 ( .A1(n10889), .A2(n7111), .ZN(n7110) );
  NAND2_X1 U9430 ( .A1(n7110), .A2(n7113), .ZN(n7850) );
  NAND3_X1 U9431 ( .A1(n7851), .A2(n7852), .A3(n7121), .ZN(n7119) );
  NAND2_X1 U9432 ( .A1(n7851), .A2(n7852), .ZN(n11155) );
  NAND2_X1 U9433 ( .A1(n11159), .A2(n7131), .ZN(n7130) );
  OAI21_X1 U9434 ( .B1(n9778), .B2(n9762), .A(n9814), .ZN(n9763) );
  OR2_X2 U9435 ( .A1(n7143), .A2(n9761), .ZN(n9778) );
  OR2_X1 U9436 ( .A1(n14923), .A2(n10198), .ZN(n7147) );
  INV_X1 U9437 ( .A(n7154), .ZN(n12581) );
  OAI211_X1 U9438 ( .C1(n14958), .C2(n11076), .A(n7159), .B(n7160), .ZN(n11001) );
  NOR2_X1 U9439 ( .A1(n10204), .A2(n10203), .ZN(n10205) );
  INV_X1 U9440 ( .A(n7167), .ZN(n12592) );
  INV_X1 U9441 ( .A(n12593), .ZN(n7166) );
  INV_X1 U9442 ( .A(n14109), .ZN(n9708) );
  INV_X1 U9443 ( .A(n11334), .ZN(n13813) );
  OR2_X2 U9444 ( .A1(n11334), .A2(n14109), .ZN(n11391) );
  AND4_X4 U9445 ( .A1(n9631), .A2(n9630), .A3(n9629), .A4(n9632), .ZN(n11334)
         );
  INV_X1 U9446 ( .A(n9202), .ZN(n9165) );
  OAI21_X2 U9447 ( .B1(n14010), .B2(n7186), .A(n7184), .ZN(n13972) );
  NAND2_X1 U9448 ( .A1(n7193), .A2(n7192), .ZN(n13880) );
  AND2_X1 U9449 ( .A1(n6563), .A2(n11296), .ZN(n7192) );
  OAI21_X2 U9450 ( .B1(n13891), .B2(n7197), .A(n7194), .ZN(n13894) );
  XNOR2_X2 U9451 ( .A(n14289), .B(n14935), .ZN(n14346) );
  NOR2_X2 U9452 ( .A1(n14287), .A2(n14288), .ZN(n14289) );
  OAI21_X2 U9453 ( .B1(n14598), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n6499), .ZN(
        n7200) );
  INV_X1 U9454 ( .A(n14377), .ZN(n7201) );
  OAI21_X1 U9455 ( .B1(n7207), .B2(n14606), .A(n7204), .ZN(n14605) );
  INV_X2 U9456 ( .A(n12030), .ZN(n12032) );
  NAND3_X1 U9457 ( .A1(n11968), .A2(n11967), .A3(n6556), .ZN(n7222) );
  INV_X1 U9458 ( .A(n11969), .ZN(n7223) );
  NAND3_X1 U9459 ( .A1(n12008), .A2(n12007), .A3(n6552), .ZN(n7234) );
  INV_X1 U9460 ( .A(n12009), .ZN(n7235) );
  NAND3_X1 U9461 ( .A1(n11979), .A2(n11978), .A3(n6553), .ZN(n7237) );
  INV_X1 U9462 ( .A(n11980), .ZN(n7238) );
  NAND3_X1 U9463 ( .A1(n11990), .A2(n11989), .A3(n6554), .ZN(n7240) );
  INV_X1 U9464 ( .A(n11991), .ZN(n7241) );
  NAND2_X1 U9465 ( .A1(n7242), .A2(n7243), .ZN(n11947) );
  NAND2_X1 U9466 ( .A1(n11920), .A2(n7247), .ZN(n7244) );
  OAI21_X1 U9467 ( .B1(n9699), .B2(n7256), .A(n9804), .ZN(n9720) );
  NAND2_X1 U9468 ( .A1(n9699), .A2(n7256), .ZN(n9804) );
  XNOR2_X1 U9469 ( .A(n9690), .B(n9803), .ZN(n7256) );
  NOR2_X1 U9470 ( .A1(n14622), .A2(n7266), .ZN(n7260) );
  AND2_X2 U9471 ( .A1(n7260), .A2(n10168), .ZN(n14619) );
  NAND3_X1 U9472 ( .A1(n7262), .A2(n10168), .A3(n7261), .ZN(n7263) );
  OAI211_X2 U9473 ( .C1(n14619), .C2(n7264), .A(n6525), .B(n7263), .ZN(n10177)
         );
  NAND2_X1 U9474 ( .A1(n13767), .A2(n7269), .ZN(n7268) );
  NAND2_X1 U9475 ( .A1(n11743), .A2(n7276), .ZN(n7273) );
  INV_X1 U9476 ( .A(n7442), .ZN(n7278) );
  NAND2_X1 U9477 ( .A1(n7279), .A2(n6541), .ZN(n13727) );
  NAND2_X1 U9478 ( .A1(n7282), .A2(n7280), .ZN(n13693) );
  NAND2_X1 U9479 ( .A1(n13757), .A2(n6545), .ZN(n13700) );
  NOR2_X2 U9480 ( .A1(n9687), .A2(n11379), .ZN(n14686) );
  NAND2_X2 U9481 ( .A1(n14419), .A2(n11858), .ZN(n9799) );
  OR2_X1 U9482 ( .A1(n11334), .A2(n9799), .ZN(n9689) );
  NAND2_X1 U9483 ( .A1(n9172), .A2(n7290), .ZN(n7293) );
  NAND2_X1 U9484 ( .A1(n7296), .A2(n7295), .ZN(n10698) );
  CLKBUF_X1 U9485 ( .A(n7296), .Z(n7294) );
  NAND2_X1 U9486 ( .A1(n10371), .A2(n10370), .ZN(n10372) );
  INV_X1 U9487 ( .A(n7294), .ZN(n10640) );
  INV_X1 U9488 ( .A(n10373), .ZN(n7297) );
  NAND2_X1 U9489 ( .A1(n13067), .A2(n7301), .ZN(n7300) );
  OAI211_X1 U9490 ( .C1(n13067), .C2(n7303), .A(n7300), .B(n13079), .ZN(n9030)
         );
  OAI211_X1 U9491 ( .C1(n11089), .C2(n7324), .A(n7322), .B(n7319), .ZN(n11244)
         );
  NAND2_X1 U9492 ( .A1(n11089), .A2(n6489), .ZN(n7319) );
  NOR2_X1 U9493 ( .A1(n8989), .A2(n7324), .ZN(n7323) );
  NAND2_X1 U9494 ( .A1(n13006), .A2(n7325), .ZN(n13060) );
  NOR2_X1 U9495 ( .A1(n7644), .A2(P2_U3088), .ZN(n7328) );
  NOR2_X1 U9496 ( .A1(n13671), .A2(n12138), .ZN(n7329) );
  NAND2_X1 U9497 ( .A1(n10037), .A2(n8934), .ZN(n10066) );
  NAND3_X1 U9498 ( .A1(n10038), .A2(n8926), .A3(n10095), .ZN(n10037) );
  INV_X1 U9499 ( .A(n14013), .ZN(n7349) );
  NAND2_X1 U9500 ( .A1(n13955), .A2(n7357), .ZN(n7356) );
  OAI211_X1 U9501 ( .C1(n13955), .C2(n7362), .A(n7358), .B(n7356), .ZN(n14125)
         );
  INV_X1 U9502 ( .A(n11177), .ZN(n7371) );
  AND2_X1 U9503 ( .A1(n9164), .A2(n7374), .ZN(n7373) );
  NAND3_X1 U9504 ( .A1(n9165), .A2(n9840), .A3(n9164), .ZN(n9991) );
  NAND3_X1 U9505 ( .A1(n11390), .A2(n11391), .A3(n9732), .ZN(n9874) );
  XNOR2_X2 U9506 ( .A(n7375), .B(n13812), .ZN(n9732) );
  INV_X1 U9507 ( .A(n9732), .ZN(n11677) );
  OAI22_X1 U9508 ( .A1(n14678), .A2(n6520), .B1(n7376), .B2(n6463), .ZN(n10480) );
  INV_X1 U9509 ( .A(n14678), .ZN(n7378) );
  INV_X1 U9510 ( .A(n10335), .ZN(n7379) );
  NAND2_X2 U9511 ( .A1(n14079), .A2(n7380), .ZN(n14192) );
  NAND2_X2 U9512 ( .A1(n14080), .A2(n6771), .ZN(n14079) );
  AND2_X1 U9513 ( .A1(n10763), .A2(n10761), .ZN(n7385) );
  INV_X1 U9514 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7389) );
  AND2_X2 U9515 ( .A1(n7390), .A2(n7388), .ZN(n7529) );
  NAND4_X1 U9516 ( .A1(n7518), .A2(n7389), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7388) );
  NAND4_X1 U9517 ( .A1(n7517), .A2(n7516), .A3(n7515), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7390) );
  INV_X1 U9518 ( .A(n7529), .ZN(n7519) );
  NAND2_X1 U9519 ( .A1(n7854), .A2(n7853), .ZN(n7856) );
  NAND2_X1 U9520 ( .A1(n7397), .A2(n7401), .ZN(n7904) );
  NAND2_X1 U9521 ( .A1(n7854), .A2(n7398), .ZN(n7397) );
  AND2_X1 U9522 ( .A1(n7411), .A2(n6557), .ZN(n10444) );
  INV_X1 U9523 ( .A(n7411), .ZN(n10355) );
  NAND2_X1 U9524 ( .A1(n7412), .A2(n7413), .ZN(n12201) );
  OAI21_X1 U9525 ( .B1(n12251), .B2(n7426), .A(n7424), .ZN(n12223) );
  NAND3_X1 U9526 ( .A1(n8173), .A2(n8178), .A3(n8172), .ZN(n7429) );
  NAND2_X1 U9527 ( .A1(n8712), .A2(n8181), .ZN(n8715) );
  NOR2_X2 U9528 ( .A1(n14142), .A2(n13961), .ZN(n13947) );
  NAND2_X1 U9529 ( .A1(n13510), .A2(n13509), .ZN(n13511) );
  AND2_X1 U9530 ( .A1(n12648), .A2(n15036), .ZN(n8711) );
  NAND2_X1 U9531 ( .A1(n13612), .A2(n14885), .ZN(n13510) );
  NAND2_X1 U9532 ( .A1(n12272), .A2(n12468), .ZN(n12294) );
  AND2_X1 U9533 ( .A1(n7906), .A2(n7935), .ZN(n10628) );
  NAND2_X1 U9534 ( .A1(n8919), .A2(n8918), .ZN(n10129) );
  NAND2_X1 U9535 ( .A1(n8997), .A2(n8996), .ZN(n13038) );
  NAND2_X1 U9536 ( .A1(n13215), .A2(n13214), .ZN(n13222) );
  INV_X1 U9537 ( .A(n13221), .ZN(n13215) );
  INV_X1 U9538 ( .A(n14686), .ZN(n14572) );
  NAND2_X1 U9539 ( .A1(n12092), .A2(n12087), .ZN(n12088) );
  NOR2_X1 U9540 ( .A1(n13465), .A2(n13312), .ZN(n9060) );
  NAND2_X1 U9541 ( .A1(n8783), .A2(n8668), .ZN(n12331) );
  XNOR2_X1 U9542 ( .A(n8921), .B(n8920), .ZN(n10132) );
  OR2_X1 U9543 ( .A1(n9616), .A2(n9235), .ZN(n9617) );
  INV_X1 U9544 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7516) );
  AOI21_X1 U9545 ( .B1(n9062), .B2(n13098), .A(n13120), .ZN(n9076) );
  INV_X1 U9546 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7515) );
  INV_X1 U9547 ( .A(n14180), .ZN(n13775) );
  NOR2_X2 U9548 ( .A1(n14180), .A2(n14041), .ZN(n14029) );
  NAND2_X1 U9549 ( .A1(n7608), .A2(SI_24_), .ZN(n7614) );
  NAND2_X1 U9550 ( .A1(n9613), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9250) );
  NAND2_X1 U9551 ( .A1(n6442), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7666) );
  INV_X1 U9552 ( .A(n6442), .ZN(n8082) );
  NAND2_X1 U9553 ( .A1(n8214), .A2(n8213), .ZN(n8668) );
  XNOR2_X1 U9554 ( .A(n10245), .B(n8788), .ZN(n8782) );
  NAND2_X1 U9555 ( .A1(n10393), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8193) );
  AND2_X1 U9556 ( .A1(n9059), .A2(n9058), .ZN(n13098) );
  AND2_X1 U9557 ( .A1(n14885), .A2(n14873), .ZN(n13596) );
  INV_X1 U9558 ( .A(n9117), .ZN(n12645) );
  AND2_X1 U9559 ( .A1(n9753), .A2(n6534), .ZN(n7438) );
  OR2_X1 U9560 ( .A1(n12637), .A2(n12979), .ZN(n7439) );
  AND2_X1 U9561 ( .A1(n10174), .A2(n10173), .ZN(n7440) );
  OR2_X1 U9562 ( .A1(n9802), .A2(n9803), .ZN(n7441) );
  AND2_X1 U9563 ( .A1(n11741), .A2(n11740), .ZN(n7442) );
  OR2_X1 U9564 ( .A1(n10697), .A2(n10696), .ZN(n7443) );
  INV_X1 U9565 ( .A(n12833), .ZN(n12863) );
  INV_X1 U9566 ( .A(n12858), .ZN(n12837) );
  INV_X1 U9567 ( .A(n12060), .ZN(n14257) );
  INV_X1 U9568 ( .A(n8837), .ZN(n8835) );
  INV_X1 U9569 ( .A(SI_20_), .ZN(n10033) );
  OR2_X1 U9570 ( .A1(n13213), .A2(n13212), .ZN(P2_U3233) );
  NAND2_X1 U9571 ( .A1(n12423), .A2(n12424), .ZN(n7446) );
  INV_X1 U9572 ( .A(n14767), .ZN(n14748) );
  XOR2_X1 U9573 ( .A(n11703), .B(n11702), .Z(n7447) );
  OR2_X1 U9574 ( .A1(n12859), .A2(n14481), .ZN(n7449) );
  MUX2_X1 U9575 ( .A(n13145), .B(n15068), .S(n12032), .Z(n11896) );
  MUX2_X1 U9576 ( .A(n13143), .B(n11908), .S(n12032), .Z(n11909) );
  INV_X1 U9577 ( .A(n14221), .ZN(n11492) );
  NAND2_X1 U9578 ( .A1(n11493), .A2(n11492), .ZN(n11494) );
  MUX2_X1 U9579 ( .A(n13428), .B(n13634), .S(n12031), .Z(n11980) );
  MUX2_X1 U9580 ( .A(n13131), .B(n13553), .S(n12031), .Z(n11996) );
  MUX2_X1 U9581 ( .A(n13129), .B(n13313), .S(n12031), .Z(n12009) );
  MUX2_X1 U9582 ( .A(n13128), .B(n13529), .S(n12031), .Z(n12015) );
  AND3_X1 U9583 ( .A1(n15080), .A2(n15123), .A3(n7491), .ZN(n7473) );
  INV_X1 U9584 ( .A(n8849), .ZN(n8847) );
  INV_X1 U9585 ( .A(n10992), .ZN(n10993) );
  INV_X1 U9586 ( .A(n12772), .ZN(n8690) );
  INV_X1 U9587 ( .A(n12032), .ZN(n12077) );
  OR2_X1 U9588 ( .A1(n11352), .A2(n8810), .ZN(n8811) );
  AND2_X1 U9589 ( .A1(n12290), .A2(n12318), .ZN(n12291) );
  INV_X1 U9590 ( .A(n8563), .ZN(n8562) );
  INV_X1 U9591 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12159) );
  INV_X1 U9592 ( .A(n12317), .ZN(n9089) );
  INV_X1 U9593 ( .A(n8464), .ZN(n8463) );
  INV_X1 U9594 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n9936) );
  NAND2_X1 U9595 ( .A1(n10302), .A2(n10299), .ZN(n10301) );
  INV_X1 U9596 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8200) );
  INV_X1 U9597 ( .A(n13040), .ZN(n8996) );
  AND2_X1 U9598 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7705) );
  NAND2_X1 U9599 ( .A1(n11308), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11517) );
  OAI21_X1 U9600 ( .B1(n10140), .B2(n9875), .A(n11396), .ZN(n9911) );
  INV_X1 U9601 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9167) );
  NAND2_X1 U9602 ( .A1(n7568), .A2(n9299), .ZN(n7571) );
  INV_X1 U9603 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9260) );
  INV_X1 U9604 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14283) );
  INV_X1 U9605 ( .A(n9120), .ZN(n9118) );
  OR2_X1 U9606 ( .A1(n8532), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8550) );
  INV_X1 U9607 ( .A(n8590), .ZN(n8589) );
  OR2_X1 U9608 ( .A1(n8631), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8657) );
  OR2_X1 U9609 ( .A1(n8447), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8464) );
  INV_X1 U9610 ( .A(n9941), .ZN(n10202) );
  XNOR2_X1 U9611 ( .A(n10992), .B(n10727), .ZN(n10728) );
  NOR2_X1 U9612 ( .A1(n10227), .A2(n12860), .ZN(n9100) );
  AND2_X1 U9613 ( .A1(n12433), .A2(n12432), .ZN(n12731) );
  NAND2_X1 U9614 ( .A1(n8499), .A2(n8498), .ZN(n8519) );
  NAND2_X1 U9615 ( .A1(n8415), .A2(n8414), .ZN(n8431) );
  NAND2_X1 U9616 ( .A1(n15006), .A2(n10082), .ZN(n12342) );
  NAND2_X1 U9617 ( .A1(n10949), .A2(n8679), .ZN(n11112) );
  AND2_X1 U9618 ( .A1(n8710), .A2(n12484), .ZN(n8743) );
  INV_X1 U9619 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8203) );
  INV_X1 U9620 ( .A(n13112), .ZN(n9048) );
  AND2_X1 U9621 ( .A1(n9479), .A2(n9478), .ZN(n9648) );
  NOR2_X1 U9622 ( .A1(n8048), .A2(n7647), .ZN(n8065) );
  NAND2_X1 U9623 ( .A1(n8036), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8048) );
  OR2_X1 U9624 ( .A1(n7775), .A2(n7774), .ZN(n7791) );
  XNOR2_X1 U9625 ( .A(n13144), .B(n14872), .ZN(n11898) );
  NAND2_X1 U9626 ( .A1(n10166), .A2(n10165), .ZN(n10167) );
  NOR2_X1 U9627 ( .A1(n10918), .A2(n10919), .ZN(n10920) );
  INV_X1 U9628 ( .A(n13729), .ZN(n11782) );
  NAND2_X1 U9629 ( .A1(n10361), .A2(n9693), .ZN(n9695) );
  AND2_X1 U9630 ( .A1(n13916), .A2(n11628), .ZN(n11874) );
  OR3_X1 U9631 ( .A1(n11517), .A2(n13760), .A3(n13695), .ZN(n11531) );
  INV_X1 U9632 ( .A(n14118), .ZN(n13866) );
  INV_X1 U9633 ( .A(n11682), .ZN(n10336) );
  INV_X1 U9634 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9244) );
  AND2_X1 U9635 ( .A1(n7571), .A2(n7570), .ZN(n7853) );
  INV_X1 U9636 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9288) );
  NOR2_X1 U9637 ( .A1(n14330), .A2(n14329), .ZN(n14299) );
  NAND2_X1 U9638 ( .A1(n9191), .A2(n12981), .ZN(n9756) );
  INV_X1 U9639 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n8297) );
  NAND2_X1 U9640 ( .A1(n8549), .A2(n8548), .ZN(n8563) );
  INV_X1 U9641 ( .A(n12820), .ZN(n12160) );
  NAND2_X1 U9642 ( .A1(n8589), .A2(n8588), .ZN(n8601) );
  NAND2_X1 U9643 ( .A1(n8885), .A2(n8881), .ZN(n12261) );
  OR2_X1 U9644 ( .A1(n8872), .A2(n9756), .ZN(n8863) );
  OR2_X1 U9645 ( .A1(n8638), .A2(n12452), .ZN(n8639) );
  INV_X1 U9646 ( .A(n8687), .ZN(n12788) );
  NAND2_X1 U9647 ( .A1(n12809), .A2(n12810), .ZN(n12808) );
  OR2_X1 U9648 ( .A1(n8882), .A2(n12457), .ZN(n12860) );
  INV_X1 U9649 ( .A(n10909), .ZN(n12300) );
  INV_X1 U9650 ( .A(n12484), .ZN(n8651) );
  NAND2_X1 U9651 ( .A1(n8609), .A2(n8608), .ZN(n8611) );
  NAND2_X1 U9652 ( .A1(n8489), .A2(n8488), .ZN(n8492) );
  OR2_X1 U9653 ( .A1(n7987), .A2(n13024), .ZN(n8004) );
  NAND2_X1 U9654 ( .A1(n8936), .A2(n8935), .ZN(n10064) );
  OR2_X1 U9655 ( .A1(n14850), .A2(n10261), .ZN(n9069) );
  NOR2_X1 U9656 ( .A1(n8004), .A2(n13081), .ZN(n8019) );
  INV_X1 U9657 ( .A(n13610), .ZN(n13214) );
  INV_X1 U9658 ( .A(n8164), .ZN(n8165) );
  INV_X1 U9659 ( .A(n13358), .ZN(n13370) );
  INV_X1 U9660 ( .A(n13493), .ZN(n14839) );
  NAND2_X1 U9661 ( .A1(n14883), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n13509) );
  INV_X1 U9662 ( .A(n12123), .ZN(n13269) );
  INV_X1 U9663 ( .A(n11944), .ZN(n14493) );
  XNOR2_X1 U9664 ( .A(n11923), .B(n13140), .ZN(n12094) );
  AND2_X1 U9665 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n7501) );
  INV_X1 U9666 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7869) );
  INV_X1 U9667 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10843) );
  OR2_X1 U9668 ( .A1(n13917), .A2(n13915), .ZN(n13733) );
  NOR2_X1 U9669 ( .A1(n10178), .A2(n9592), .ZN(n11720) );
  AND2_X1 U9670 ( .A1(n11627), .A2(n11617), .ZN(n13948) );
  AND2_X1 U9671 ( .A1(n11546), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11562) );
  INV_X1 U9672 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11218) );
  INV_X1 U9673 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10835) );
  INV_X1 U9674 ( .A(n11375), .ZN(n11379) );
  OR2_X1 U9675 ( .A1(n9712), .A2(n9711), .ZN(n13917) );
  NOR2_X1 U9676 ( .A1(n11655), .A2(n15172), .ZN(n11656) );
  AND2_X1 U9677 ( .A1(n9713), .A2(n13816), .ZN(n14766) );
  NAND2_X1 U9678 ( .A1(n14019), .A2(n9700), .ZN(n14767) );
  AND2_X1 U9679 ( .A1(n7584), .A2(n7583), .ZN(n7903) );
  NAND2_X1 U9680 ( .A1(n8351), .A2(n8350), .ZN(n8383) );
  NAND2_X1 U9681 ( .A1(n8814), .A2(n7448), .ZN(n11338) );
  AND2_X1 U9682 ( .A1(n8885), .A2(n8884), .ZN(n12264) );
  NAND2_X1 U9683 ( .A1(n8879), .A2(n8878), .ZN(n12243) );
  INV_X1 U9684 ( .A(n12280), .ZN(n12624) );
  AND2_X1 U9685 ( .A1(n8607), .A2(n8606), .ZN(n12653) );
  AND4_X1 U9686 ( .A1(n8421), .A2(n8420), .A3(n8419), .A4(n8418), .ZN(n12861)
         );
  OR2_X1 U9687 ( .A1(n8245), .A2(n10308), .ZN(n8219) );
  NOR2_X1 U9688 ( .A1(n10987), .A2(n10986), .ZN(n14957) );
  INV_X1 U9689 ( .A(n14979), .ZN(n14944) );
  INV_X1 U9690 ( .A(n12872), .ZN(n12831) );
  INV_X1 U9691 ( .A(n12828), .ZN(n12864) );
  INV_X1 U9692 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10564) );
  AND2_X1 U9693 ( .A1(n8868), .A2(n8867), .ZN(n12828) );
  AND2_X1 U9694 ( .A1(n8755), .A2(n8754), .ZN(n10057) );
  INV_X1 U9695 ( .A(n15044), .ZN(n15007) );
  OR2_X1 U9696 ( .A1(n11117), .A2(n15036), .ZN(n15049) );
  INV_X1 U9697 ( .A(n15039), .ZN(n15036) );
  NAND2_X1 U9698 ( .A1(n9964), .A2(n8916), .ZN(n10131) );
  NAND2_X1 U9699 ( .A1(n9061), .A2(n13487), .ZN(n13120) );
  OR2_X1 U9700 ( .A1(n14808), .A2(n14807), .ZN(n14809) );
  INV_X1 U9701 ( .A(n14806), .ZN(n14824) );
  INV_X1 U9702 ( .A(n12124), .ZN(n8155) );
  INV_X1 U9703 ( .A(n13474), .ZN(n14842) );
  AND2_X1 U9704 ( .A1(n14876), .A2(n8915), .ZN(n13603) );
  INV_X1 U9705 ( .A(n13603), .ZN(n13584) );
  AND3_X1 U9706 ( .A1(n14850), .A2(n14854), .A3(n8769), .ZN(n10263) );
  INV_X1 U9707 ( .A(n13733), .ZN(n14625) );
  INV_X1 U9708 ( .A(n14628), .ZN(n13798) );
  AND4_X1 U9709 ( .A1(n11632), .A2(n11631), .A3(n11630), .A4(n11629), .ZN(
        n14138) );
  AND3_X1 U9710 ( .A1(n11521), .A2(n11520), .A3(n11519), .ZN(n14203) );
  AND4_X1 U9711 ( .A1(n11049), .A2(n11048), .A3(n11047), .A4(n11046), .ZN(
        n14501) );
  INV_X1 U9712 ( .A(n14668), .ZN(n14652) );
  INV_X1 U9713 ( .A(n14666), .ZN(n14643) );
  XOR2_X1 U9714 ( .A(n13928), .B(n13909), .Z(n13908) );
  INV_X1 U9715 ( .A(n14574), .ZN(n14763) );
  INV_X1 U9716 ( .A(n14197), .ZN(n14069) );
  AND2_X1 U9717 ( .A1(n14437), .A2(n14763), .ZN(n14434) );
  INV_X1 U9718 ( .A(n9847), .ZN(n13915) );
  AND2_X1 U9719 ( .A1(n9853), .A2(n14730), .ZN(n14755) );
  INV_X1 U9720 ( .A(n14755), .ZN(n14774) );
  AND2_X1 U9721 ( .A1(n9608), .A2(n9607), .ZN(n9847) );
  NAND2_X1 U9722 ( .A1(n9254), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9592) );
  AND2_X1 U9723 ( .A1(n9290), .A2(n9293), .ZN(n10475) );
  NAND2_X1 U9724 ( .A1(n8740), .A2(n8739), .ZN(n9191) );
  INV_X1 U9725 ( .A(n8890), .ZN(n8891) );
  AND2_X1 U9726 ( .A1(n10399), .A2(n9097), .ZN(n12289) );
  INV_X1 U9727 ( .A(n12705), .ZN(n12667) );
  OR2_X1 U9728 ( .A1(n9765), .A2(n9773), .ZN(n14989) );
  OR2_X1 U9729 ( .A1(n9765), .A2(n9764), .ZN(n14995) );
  INV_X1 U9730 ( .A(n12863), .ZN(n12868) );
  OR2_X1 U9731 ( .A1(n12833), .A2(n11118), .ZN(n12872) );
  AND2_X1 U9732 ( .A1(n10059), .A2(n12864), .ZN(n12833) );
  INV_X1 U9733 ( .A(n12647), .ZN(n10957) );
  NAND2_X1 U9734 ( .A1(n9117), .A2(n8767), .ZN(n8768) );
  INV_X1 U9735 ( .A(n15066), .ZN(n15064) );
  NAND2_X1 U9736 ( .A1(n15066), .A2(n15007), .ZN(n12928) );
  AND2_X1 U9737 ( .A1(n8749), .A2(n8748), .ZN(n15050) );
  NAND2_X1 U9738 ( .A1(n9285), .A2(n12981), .ZN(n9286) );
  INV_X1 U9739 ( .A(n8740), .ZN(n11322) );
  INV_X1 U9740 ( .A(SI_15_), .ZN(n9348) );
  INV_X1 U9741 ( .A(n14397), .ZN(n12997) );
  AND2_X1 U9742 ( .A1(n9073), .A2(n9072), .ZN(n9074) );
  INV_X1 U9743 ( .A(n13120), .ZN(n13077) );
  INV_X1 U9744 ( .A(n13098), .ZN(n13122) );
  INV_X1 U9745 ( .A(n14822), .ZN(n10637) );
  OR2_X1 U9746 ( .A1(n10264), .A2(n6689), .ZN(n13410) );
  INV_X1 U9747 ( .A(n13490), .ZN(n15079) );
  AND2_X1 U9748 ( .A1(n13392), .A2(n13391), .ZN(n13568) );
  INV_X1 U9749 ( .A(n14885), .ZN(n14883) );
  NAND2_X1 U9750 ( .A1(n14880), .A2(n14873), .ZN(n13640) );
  INV_X1 U9751 ( .A(n14880), .ZN(n14879) );
  NOR2_X1 U9752 ( .A1(n14851), .A2(n14846), .ZN(n14847) );
  INV_X1 U9753 ( .A(n14847), .ZN(n14848) );
  INV_X1 U9754 ( .A(n14854), .ZN(n14851) );
  XNOR2_X1 U9755 ( .A(n7483), .B(n7626), .ZN(n13663) );
  INV_X1 U9756 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9419) );
  AND2_X1 U9757 ( .A1(n10182), .A2(n14274), .ZN(n14628) );
  NAND2_X1 U9758 ( .A1(n9706), .A2(n9705), .ZN(n14620) );
  OR2_X1 U9759 ( .A1(n14635), .A2(n11719), .ZN(n14668) );
  OR2_X1 U9760 ( .A1(n14635), .A2(n13816), .ZN(n14670) );
  NAND2_X1 U9761 ( .A1(n14437), .A2(n14009), .ZN(n14700) );
  NAND2_X1 U9762 ( .A1(n9850), .A2(n9849), .ZN(n14706) );
  OR2_X1 U9763 ( .A1(n9722), .A2(n13915), .ZN(n14787) );
  NAND2_X1 U9764 ( .A1(n9850), .A2(n9606), .ZN(n14708) );
  INV_X1 U9765 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10075) );
  INV_X1 U9766 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n15111) );
  NOR2_X2 U9767 ( .A1(n9191), .A2(n9190), .ZN(P3_U3897) );
  NOR2_X1 U9768 ( .A1(n9455), .A2(n9156), .ZN(P2_U3947) );
  INV_X1 U9769 ( .A(n13817), .ZN(P1_U4016) );
  NOR4_X1 U9770 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n7458) );
  OR4_X1 U9771 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n7455) );
  NOR4_X1 U9772 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n7453) );
  NOR4_X1 U9773 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n7452) );
  NOR4_X1 U9774 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n7451) );
  NOR4_X1 U9775 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n7450) );
  NAND4_X1 U9776 ( .A1(n7453), .A2(n7452), .A3(n7451), .A4(n7450), .ZN(n7454)
         );
  NOR4_X1 U9777 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        n7455), .A4(n7454), .ZN(n7457) );
  NOR4_X1 U9778 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n7456) );
  NAND3_X1 U9779 ( .A1(n7458), .A2(n7457), .A3(n7456), .ZN(n7485) );
  AND3_X2 U9780 ( .A1(n7463), .A2(n7462), .A3(n7461), .ZN(n7833) );
  NOR2_X1 U9781 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7468) );
  NOR2_X1 U9782 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7467) );
  NOR2_X1 U9783 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n7466) );
  INV_X1 U9784 ( .A(n7490), .ZN(n7469) );
  NAND2_X1 U9785 ( .A1(n7509), .A2(n7510), .ZN(n7478) );
  NAND2_X1 U9786 ( .A1(n7480), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7470) );
  MUX2_X1 U9787 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7470), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n7477) );
  INV_X2 U9788 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n15123) );
  NOR2_X1 U9789 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n7472) );
  NOR2_X1 U9790 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n7471) );
  NAND2_X1 U9791 ( .A1(n7477), .A2(n7482), .ZN(n13665) );
  NAND2_X1 U9792 ( .A1(n7478), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7479) );
  MUX2_X1 U9793 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7479), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n7481) );
  INV_X1 U9794 ( .A(P2_B_REG_SCAN_IN), .ZN(n8162) );
  XOR2_X1 U9795 ( .A(n11271), .B(n8162), .Z(n7484) );
  NAND2_X1 U9796 ( .A1(n7482), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7483) );
  NAND2_X1 U9797 ( .A1(n7485), .A2(n14846), .ZN(n9056) );
  INV_X1 U9798 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14852) );
  NAND2_X1 U9799 ( .A1(n14846), .A2(n14852), .ZN(n7487) );
  NAND2_X1 U9800 ( .A1(n13665), .A2(n13663), .ZN(n7486) );
  NAND2_X1 U9801 ( .A1(n7487), .A2(n7486), .ZN(n14853) );
  NAND2_X1 U9802 ( .A1(n7493), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7494) );
  XNOR2_X2 U9803 ( .A(n7494), .B(n15123), .ZN(n12091) );
  INV_X1 U9804 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7495) );
  INV_X1 U9805 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7498) );
  INV_X1 U9806 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7497) );
  NAND3_X1 U9807 ( .A1(n7498), .A2(n7497), .A3(P2_IR_REG_19__SCAN_IN), .ZN(
        n7500) );
  XNOR2_X1 U9808 ( .A(P2_IR_REG_31__SCAN_IN), .B(P2_IR_REG_19__SCAN_IN), .ZN(
        n7499) );
  INV_X1 U9809 ( .A(n9060), .ZN(n9068) );
  AND2_X1 U9810 ( .A1(n14853), .A2(n9068), .ZN(n7503) );
  INV_X1 U9811 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14849) );
  NAND2_X1 U9812 ( .A1(n14846), .A2(n14849), .ZN(n7505) );
  NAND2_X1 U9813 ( .A1(n11271), .A2(n13663), .ZN(n7504) );
  NAND2_X1 U9814 ( .A1(n7505), .A2(n7504), .ZN(n14850) );
  INV_X1 U9815 ( .A(n13665), .ZN(n7507) );
  NOR2_X1 U9816 ( .A1(n11271), .A2(n13663), .ZN(n7506) );
  NAND2_X1 U9817 ( .A1(n13312), .A2(n12091), .ZN(n12064) );
  NAND2_X1 U9818 ( .A1(n8102), .A2(n8101), .ZN(n9057) );
  INV_X1 U9819 ( .A(n9057), .ZN(n9451) );
  NAND2_X1 U9820 ( .A1(n12064), .A2(n9451), .ZN(n8769) );
  OR2_X1 U9821 ( .A1(n7509), .A2(n7869), .ZN(n7511) );
  AND2_X1 U9822 ( .A1(n8769), .A2(n12090), .ZN(n7512) );
  AND2_X1 U9823 ( .A1(n9455), .A2(n7512), .ZN(n9070) );
  NAND2_X1 U9824 ( .A1(n9070), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7513) );
  NOR2_X1 U9825 ( .A1(n14850), .A2(n7513), .ZN(n7514) );
  NAND2_X1 U9826 ( .A1(n12064), .A2(n14859), .ZN(n14864) );
  INV_X1 U9827 ( .A(n13596), .ZN(n8170) );
  NAND2_X1 U9828 ( .A1(n7519), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7521) );
  NAND2_X1 U9829 ( .A1(n7529), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7520) );
  INV_X1 U9830 ( .A(SI_1_), .ZN(n9256) );
  AND2_X1 U9831 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7522) );
  NAND2_X1 U9832 ( .A1(n7530), .A2(n7522), .ZN(n9627) );
  AND2_X1 U9833 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7523) );
  NAND2_X1 U9834 ( .A1(n7529), .A2(n7523), .ZN(n7660) );
  NAND2_X1 U9835 ( .A1(n9627), .A2(n7660), .ZN(n7667) );
  NAND2_X1 U9836 ( .A1(n7668), .A2(n7667), .ZN(n7526) );
  NAND2_X1 U9837 ( .A1(n7524), .A2(SI_1_), .ZN(n7525) );
  INV_X1 U9838 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9725) );
  INV_X1 U9839 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9213) );
  MUX2_X1 U9840 ( .A(n9725), .B(n9213), .S(n11363), .Z(n7685) );
  NAND2_X1 U9841 ( .A1(n7527), .A2(SI_2_), .ZN(n7528) );
  XNOR2_X1 U9842 ( .A(n7534), .B(SI_3_), .ZN(n7700) );
  INV_X1 U9843 ( .A(n7700), .ZN(n7533) );
  NAND2_X1 U9844 ( .A1(n7534), .A2(SI_3_), .ZN(n7535) );
  NAND2_X1 U9845 ( .A1(n7536), .A2(n7535), .ZN(n7711) );
  MUX2_X1 U9846 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n11542), .Z(n7538) );
  XNOR2_X1 U9847 ( .A(n7538), .B(SI_4_), .ZN(n7710) );
  INV_X1 U9848 ( .A(n7710), .ZN(n7537) );
  NAND2_X1 U9849 ( .A1(n7711), .A2(n7537), .ZN(n7540) );
  NAND2_X1 U9850 ( .A1(n7538), .A2(SI_4_), .ZN(n7539) );
  NAND2_X1 U9851 ( .A1(n7540), .A2(n7539), .ZN(n7719) );
  MUX2_X1 U9852 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n11542), .Z(n7542) );
  XNOR2_X1 U9853 ( .A(n7542), .B(SI_5_), .ZN(n7720) );
  INV_X1 U9854 ( .A(n7720), .ZN(n7541) );
  NAND2_X1 U9855 ( .A1(n7719), .A2(n7541), .ZN(n7544) );
  NAND2_X1 U9856 ( .A1(n7542), .A2(SI_5_), .ZN(n7543) );
  MUX2_X1 U9857 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n11542), .Z(n7546) );
  XNOR2_X1 U9858 ( .A(n7546), .B(SI_6_), .ZN(n7738) );
  INV_X1 U9859 ( .A(n7738), .ZN(n7545) );
  NAND2_X1 U9860 ( .A1(n7546), .A2(SI_6_), .ZN(n7547) );
  MUX2_X1 U9861 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n11542), .Z(n7549) );
  XNOR2_X1 U9862 ( .A(n7549), .B(SI_7_), .ZN(n7751) );
  INV_X1 U9863 ( .A(n7751), .ZN(n7548) );
  MUX2_X1 U9864 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n11542), .Z(n7551) );
  XNOR2_X1 U9865 ( .A(n7551), .B(SI_8_), .ZN(n7765) );
  INV_X1 U9866 ( .A(n7765), .ZN(n7550) );
  NAND2_X1 U9867 ( .A1(n7551), .A2(SI_8_), .ZN(n7552) );
  MUX2_X1 U9868 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n11542), .Z(n7554) );
  XNOR2_X1 U9869 ( .A(n7554), .B(SI_9_), .ZN(n7782) );
  INV_X1 U9870 ( .A(n7782), .ZN(n7553) );
  NAND2_X1 U9871 ( .A1(n7554), .A2(SI_9_), .ZN(n7555) );
  MUX2_X1 U9872 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n11542), .Z(n7557) );
  NAND2_X1 U9873 ( .A1(n7557), .A2(SI_10_), .ZN(n7558) );
  INV_X1 U9874 ( .A(n7560), .ZN(n7561) );
  NAND2_X1 U9875 ( .A1(n7561), .A2(SI_11_), .ZN(n7562) );
  NAND2_X1 U9876 ( .A1(n7563), .A2(n7562), .ZN(n7814) );
  MUX2_X1 U9877 ( .A(n9423), .B(n9419), .S(n11542), .Z(n7564) );
  NAND2_X1 U9878 ( .A1(n7564), .A2(n9268), .ZN(n7567) );
  INV_X1 U9879 ( .A(n7564), .ZN(n7565) );
  NAND2_X1 U9880 ( .A1(n7565), .A2(SI_12_), .ZN(n7566) );
  MUX2_X1 U9881 ( .A(n15111), .B(n9676), .S(n11542), .Z(n7568) );
  INV_X1 U9882 ( .A(n7568), .ZN(n7569) );
  NAND2_X1 U9883 ( .A1(n7569), .A2(SI_13_), .ZN(n7570) );
  MUX2_X1 U9884 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n11542), .Z(n7888) );
  NOR2_X1 U9885 ( .A1(n7888), .A2(SI_14_), .ZN(n7578) );
  MUX2_X1 U9886 ( .A(n9844), .B(n9846), .S(n11542), .Z(n7572) );
  INV_X1 U9887 ( .A(n7572), .ZN(n7573) );
  NAND2_X1 U9888 ( .A1(n7573), .A2(SI_15_), .ZN(n7574) );
  NAND2_X1 U9889 ( .A1(n7579), .A2(n7574), .ZN(n7885) );
  INV_X1 U9890 ( .A(n7888), .ZN(n7575) );
  NOR2_X1 U9891 ( .A1(n7575), .A2(n9302), .ZN(n7576) );
  MUX2_X1 U9892 ( .A(n9995), .B(n9990), .S(n11542), .Z(n7581) );
  INV_X1 U9893 ( .A(n7581), .ZN(n7582) );
  NAND2_X1 U9894 ( .A1(n7582), .A2(SI_16_), .ZN(n7583) );
  NAND2_X1 U9895 ( .A1(n7904), .A2(n7903), .ZN(n7585) );
  MUX2_X1 U9896 ( .A(n10075), .B(n10077), .S(n11542), .Z(n7917) );
  INV_X1 U9897 ( .A(SI_18_), .ZN(n9751) );
  MUX2_X1 U9898 ( .A(n10259), .B(n15202), .S(n11363), .Z(n7931) );
  MUX2_X1 U9899 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n11363), .Z(n7590) );
  XNOR2_X1 U9900 ( .A(n7590), .B(SI_19_), .ZN(n7946) );
  INV_X1 U9901 ( .A(n7590), .ZN(n7591) );
  NAND2_X1 U9902 ( .A1(n7591), .A2(n15087), .ZN(n7592) );
  INV_X1 U9903 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n15142) );
  INV_X1 U9904 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10866) );
  MUX2_X1 U9905 ( .A(n15142), .B(n10866), .S(n11363), .Z(n7964) );
  MUX2_X1 U9906 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n11363), .Z(n7596) );
  NAND2_X1 U9907 ( .A1(n7596), .A2(SI_21_), .ZN(n7599) );
  INV_X1 U9908 ( .A(n7596), .ZN(n7597) );
  INV_X1 U9909 ( .A(SI_21_), .ZN(n15192) );
  NAND2_X1 U9910 ( .A1(n7597), .A2(n15192), .ZN(n7598) );
  INV_X1 U9911 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7600) );
  MUX2_X1 U9912 ( .A(n7600), .B(n11269), .S(n11363), .Z(n8000) );
  INV_X1 U9913 ( .A(SI_22_), .ZN(n15215) );
  MUX2_X1 U9914 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n11363), .Z(n7601) );
  NAND2_X1 U9915 ( .A1(n7601), .A2(SI_23_), .ZN(n7606) );
  INV_X1 U9916 ( .A(n7601), .ZN(n7602) );
  INV_X1 U9917 ( .A(SI_23_), .ZN(n10470) );
  NAND2_X1 U9918 ( .A1(n7602), .A2(n10470), .ZN(n7603) );
  NAND2_X1 U9919 ( .A1(n7606), .A2(n7603), .ZN(n8015) );
  INV_X1 U9920 ( .A(n8000), .ZN(n7604) );
  NOR2_X1 U9921 ( .A1(n7604), .A2(SI_22_), .ZN(n7605) );
  NAND2_X1 U9922 ( .A1(n7607), .A2(n7606), .ZN(n7608) );
  INV_X1 U9923 ( .A(n7608), .ZN(n7610) );
  INV_X1 U9924 ( .A(SI_24_), .ZN(n7609) );
  NAND2_X1 U9925 ( .A1(n7610), .A2(n7609), .ZN(n7611) );
  NAND2_X1 U9926 ( .A1(n7614), .A2(n7611), .ZN(n8030) );
  INV_X1 U9927 ( .A(n8030), .ZN(n7613) );
  INV_X1 U9928 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11582) );
  INV_X1 U9929 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11270) );
  MUX2_X1 U9930 ( .A(n11582), .B(n11270), .S(n11363), .Z(n8029) );
  MUX2_X1 U9931 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n11542), .Z(n7615) );
  XNOR2_X1 U9932 ( .A(n7615), .B(SI_25_), .ZN(n8044) );
  INV_X1 U9933 ( .A(n7615), .ZN(n7616) );
  INV_X1 U9934 ( .A(SI_25_), .ZN(n10943) );
  NAND2_X1 U9935 ( .A1(n7616), .A2(n10943), .ZN(n7617) );
  INV_X1 U9936 ( .A(SI_26_), .ZN(n11320) );
  INV_X1 U9937 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14265) );
  INV_X1 U9938 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13662) );
  MUX2_X1 U9939 ( .A(n14265), .B(n13662), .S(n11363), .Z(n8058) );
  INV_X1 U9940 ( .A(n8058), .ZN(n7618) );
  INV_X1 U9941 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n11612) );
  INV_X1 U9942 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13660) );
  MUX2_X1 U9943 ( .A(n11612), .B(n13660), .S(n11363), .Z(n8073) );
  MUX2_X1 U9944 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n11363), .Z(n8078) );
  NAND2_X1 U9945 ( .A1(n8078), .A2(SI_28_), .ZN(n7619) );
  OAI21_X1 U9946 ( .B1(n8073), .B2(n7635), .A(n7619), .ZN(n7625) );
  NAND2_X1 U9947 ( .A1(n8073), .A2(n7635), .ZN(n7620) );
  NAND2_X1 U9948 ( .A1(n7620), .A2(SI_28_), .ZN(n7623) );
  INV_X1 U9949 ( .A(n8078), .ZN(n7622) );
  NOR2_X1 U9950 ( .A1(SI_27_), .A2(SI_28_), .ZN(n7621) );
  AOI22_X1 U9951 ( .A1(n7623), .A2(n7622), .B1(n7621), .B2(n8073), .ZN(n7624)
         );
  INV_X1 U9952 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14260) );
  INV_X1 U9953 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n11323) );
  MUX2_X1 U9954 ( .A(n14260), .B(n11323), .S(n11363), .Z(n11358) );
  XNOR2_X1 U9955 ( .A(n11358), .B(SI_29_), .ZN(n11356) );
  INV_X1 U9956 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7628) );
  INV_X4 U9957 ( .A(n8033), .ZN(n12059) );
  NAND2_X1 U9958 ( .A1(n11642), .A2(n12059), .ZN(n7633) );
  INV_X1 U9959 ( .A(n11363), .ZN(n9679) );
  OR2_X1 U9960 ( .A1(n12061), .A2(n11323), .ZN(n7632) );
  INV_X1 U9961 ( .A(n7634), .ZN(n7636) );
  INV_X1 U9962 ( .A(SI_27_), .ZN(n7635) );
  NAND2_X1 U9963 ( .A1(n7636), .A2(n7635), .ZN(n7637) );
  OR2_X1 U9964 ( .A1(n12061), .A2(n13660), .ZN(n7638) );
  NAND2_X1 U9965 ( .A1(n7640), .A2(n7641), .ZN(n13652) );
  NAND2_X1 U9966 ( .A1(n8093), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n7654) );
  INV_X1 U9967 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n7643) );
  OR2_X1 U9968 ( .A1(n8082), .A2(n7643), .ZN(n7653) );
  NAND2_X4 U9969 ( .A1(n7650), .A2(n7645), .ZN(n8094) );
  NAND2_X1 U9970 ( .A1(n7705), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7744) );
  INV_X1 U9971 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7743) );
  NOR2_X1 U9972 ( .A1(n7744), .A2(n7743), .ZN(n7742) );
  NAND2_X1 U9973 ( .A1(n7742), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7775) );
  INV_X1 U9974 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7774) );
  INV_X1 U9975 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7790) );
  NAND2_X1 U9976 ( .A1(n7805), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7844) );
  INV_X1 U9977 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7843) );
  INV_X1 U9978 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11127) );
  INV_X1 U9979 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7876) );
  NAND2_X1 U9980 ( .A1(n7875), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7910) );
  INV_X1 U9981 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7909) );
  INV_X1 U9982 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7924) );
  AND2_X1 U9983 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n7646) );
  NAND2_X1 U9984 ( .A1(n7955), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7987) );
  INV_X1 U9985 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13024) );
  INV_X1 U9986 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13081) );
  NAND2_X1 U9987 ( .A1(n8019), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8020) );
  INV_X1 U9988 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n7647) );
  NAND2_X1 U9989 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(n8065), .ZN(n8064) );
  INV_X1 U9990 ( .A(n8064), .ZN(n7648) );
  NAND2_X1 U9991 ( .A1(n7648), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8085) );
  INV_X1 U9992 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13000) );
  NAND2_X1 U9993 ( .A1(n8064), .A2(n13000), .ZN(n7649) );
  NAND2_X1 U9994 ( .A1(n8085), .A2(n7649), .ZN(n13251) );
  OR2_X1 U9995 ( .A1(n8094), .A2(n13251), .ZN(n7652) );
  INV_X1 U9996 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13252) );
  OR2_X1 U9997 ( .A1(n6614), .A2(n13252), .ZN(n7651) );
  NAND4_X1 U9998 ( .A1(n7654), .A2(n7653), .A3(n7652), .A4(n7651), .ZN(n13126)
         );
  INV_X1 U9999 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10268) );
  NAND2_X1 U10000 ( .A1(n6442), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7657) );
  INV_X1 U10001 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9527) );
  INV_X1 U10002 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9526) );
  NAND2_X1 U10003 ( .A1(n11542), .A2(SI_0_), .ZN(n7659) );
  INV_X1 U10004 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8195) );
  NAND2_X1 U10005 ( .A1(n7659), .A2(n8195), .ZN(n7661) );
  AND2_X1 U10006 ( .A1(n7661), .A2(n7660), .ZN(n13674) );
  MUX2_X1 U10007 ( .A(n13673), .B(n13674), .S(n7662), .Z(n14860) );
  INV_X1 U10008 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10275) );
  OR2_X1 U10009 ( .A1(n8094), .A2(n10275), .ZN(n7665) );
  INV_X1 U10010 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10274) );
  INV_X1 U10011 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9424) );
  OR2_X1 U10012 ( .A1(n7687), .A2(n9212), .ZN(n7676) );
  XNOR2_X1 U10013 ( .A(n7668), .B(n7667), .ZN(n9680) );
  NAND2_X1 U10014 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n13673), .ZN(n7669) );
  MUX2_X1 U10015 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7669), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n7673) );
  INV_X1 U10016 ( .A(n7671), .ZN(n7672) );
  NAND2_X1 U10017 ( .A1(n7673), .A2(n7672), .ZN(n9546) );
  OR2_X1 U10018 ( .A1(n7662), .A2(n9546), .ZN(n7674) );
  INV_X1 U10019 ( .A(n8917), .ZN(n10293) );
  NAND2_X1 U10020 ( .A1(n10293), .A2(n6635), .ZN(n7677) );
  NAND2_X1 U10021 ( .A1(n9831), .A2(n7677), .ZN(n10281) );
  NAND2_X1 U10022 ( .A1(n6441), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7682) );
  INV_X1 U10023 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10288) );
  OR2_X1 U10024 ( .A1(n8094), .A2(n10288), .ZN(n7681) );
  INV_X1 U10025 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n15082) );
  OR2_X1 U10026 ( .A1(n12045), .A2(n15082), .ZN(n7680) );
  INV_X1 U10027 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9427) );
  OR2_X1 U10028 ( .A1(n12049), .A2(n9427), .ZN(n7679) );
  OR2_X1 U10029 ( .A1(n7671), .A2(n7869), .ZN(n7684) );
  XNOR2_X1 U10030 ( .A(n7684), .B(n7683), .ZN(n9525) );
  XNOR2_X1 U10031 ( .A(n7686), .B(n7685), .ZN(n9724) );
  OR2_X1 U10032 ( .A1(n8033), .A2(n9724), .ZN(n7689) );
  OR2_X1 U10033 ( .A1(n7687), .A2(n9213), .ZN(n7688) );
  INV_X1 U10034 ( .A(n12095), .ZN(n7690) );
  NAND2_X1 U10035 ( .A1(n10281), .A2(n7690), .ZN(n10283) );
  INV_X1 U10036 ( .A(n13146), .ZN(n10133) );
  INV_X1 U10037 ( .A(n11890), .ZN(n14865) );
  NAND2_X1 U10038 ( .A1(n10133), .A2(n14865), .ZN(n7691) );
  NAND2_X1 U10039 ( .A1(n10283), .A2(n7691), .ZN(n10018) );
  NAND2_X1 U10040 ( .A1(n6442), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7695) );
  OR2_X1 U10041 ( .A1(n8094), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7694) );
  INV_X1 U10042 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9461) );
  OR2_X1 U10043 ( .A1(n12045), .A2(n9461), .ZN(n7693) );
  INV_X1 U10044 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9430) );
  OR2_X1 U10045 ( .A1(n12049), .A2(n9430), .ZN(n7692) );
  NAND4_X1 U10046 ( .A1(n7695), .A2(n7694), .A3(n7693), .A4(n7692), .ZN(n13145) );
  NAND2_X1 U10047 ( .A1(n7696), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7697) );
  MUX2_X1 U10048 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7697), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n7699) );
  NAND2_X1 U10049 ( .A1(n7699), .A2(n7698), .ZN(n9512) );
  NAND2_X1 U10050 ( .A1(n9857), .A2(n12059), .ZN(n7702) );
  OR2_X1 U10051 ( .A1(n12061), .A2(n9214), .ZN(n7701) );
  OAI211_X2 U10052 ( .C1(n7662), .C2(n9512), .A(n7702), .B(n7701), .ZN(n15068)
         );
  INV_X1 U10053 ( .A(n13145), .ZN(n10587) );
  NAND2_X1 U10054 ( .A1(n10587), .A2(n10027), .ZN(n7703) );
  NAND2_X1 U10055 ( .A1(n10017), .A2(n7703), .ZN(n10582) );
  NAND2_X1 U10056 ( .A1(n8093), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7709) );
  INV_X1 U10057 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7704) );
  OR2_X1 U10058 ( .A1(n8082), .A2(n7704), .ZN(n7708) );
  INV_X1 U10059 ( .A(n7705), .ZN(n7730) );
  OAI21_X1 U10060 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n7730), .ZN(n10595) );
  OR2_X1 U10061 ( .A1(n8094), .A2(n10595), .ZN(n7707) );
  INV_X1 U10062 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10591) );
  OR2_X1 U10063 ( .A1(n6614), .A2(n10591), .ZN(n7706) );
  XNOR2_X1 U10064 ( .A(n7711), .B(n7710), .ZN(n9869) );
  NAND2_X1 U10065 ( .A1(n9869), .A2(n12059), .ZN(n7717) );
  NAND2_X1 U10066 ( .A1(n7698), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7712) );
  MUX2_X1 U10067 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7712), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n7715) );
  INV_X1 U10068 ( .A(n7698), .ZN(n7714) );
  INV_X1 U10069 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7713) );
  NAND2_X1 U10070 ( .A1(n7714), .A2(n7713), .ZN(n7722) );
  NAND2_X1 U10071 ( .A1(n7715), .A2(n7722), .ZN(n9558) );
  INV_X1 U10072 ( .A(n9558), .ZN(n9465) );
  AOI22_X1 U10073 ( .A1(n7949), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7948), .B2(
        n9465), .ZN(n7716) );
  NAND2_X1 U10074 ( .A1(n7717), .A2(n7716), .ZN(n14872) );
  INV_X1 U10075 ( .A(n11898), .ZN(n12099) );
  NAND2_X1 U10076 ( .A1(n10582), .A2(n12099), .ZN(n10581) );
  INV_X1 U10077 ( .A(n13144), .ZN(n10432) );
  INV_X1 U10078 ( .A(n14872), .ZN(n11902) );
  NAND2_X1 U10079 ( .A1(n10432), .A2(n11902), .ZN(n7718) );
  XNOR2_X1 U10080 ( .A(n7719), .B(n7720), .ZN(n9894) );
  NAND2_X1 U10081 ( .A1(n9894), .A2(n12059), .ZN(n7727) );
  NAND2_X1 U10082 ( .A1(n7722), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7721) );
  MUX2_X1 U10083 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7721), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n7725) );
  INV_X1 U10084 ( .A(n7722), .ZN(n7724) );
  INV_X1 U10085 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7723) );
  NAND2_X1 U10086 ( .A1(n7724), .A2(n7723), .ZN(n7835) );
  AND2_X1 U10087 ( .A1(n7725), .A2(n7835), .ZN(n9563) );
  AOI22_X1 U10088 ( .A1(n7949), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7948), .B2(
        n9563), .ZN(n7726) );
  NAND2_X1 U10089 ( .A1(n7727), .A2(n7726), .ZN(n11908) );
  NAND2_X1 U10090 ( .A1(n8093), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7735) );
  INV_X1 U10091 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7728) );
  OR2_X1 U10092 ( .A1(n8082), .A2(n7728), .ZN(n7734) );
  INV_X1 U10093 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7729) );
  NAND2_X1 U10094 ( .A1(n7730), .A2(n7729), .ZN(n7731) );
  NAND2_X1 U10095 ( .A1(n7744), .A2(n7731), .ZN(n10602) );
  OR2_X1 U10096 ( .A1(n8094), .A2(n10602), .ZN(n7733) );
  INV_X1 U10097 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10601) );
  OR2_X1 U10098 ( .A1(n6614), .A2(n10601), .ZN(n7732) );
  NAND4_X1 U10099 ( .A1(n7735), .A2(n7734), .A3(n7733), .A4(n7732), .ZN(n13143) );
  XNOR2_X1 U10100 ( .A(n11908), .B(n13143), .ZN(n12101) );
  INV_X1 U10101 ( .A(n12101), .ZN(n10433) );
  OR2_X1 U10102 ( .A1(n11908), .A2(n13143), .ZN(n7736) );
  NAND2_X1 U10103 ( .A1(n10427), .A2(n7736), .ZN(n10232) );
  XNOR2_X1 U10104 ( .A(n7737), .B(n7738), .ZN(n10104) );
  NAND2_X1 U10105 ( .A1(n10104), .A2(n12059), .ZN(n7741) );
  NAND2_X1 U10106 ( .A1(n7835), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7739) );
  XNOR2_X1 U10107 ( .A(n7739), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9468) );
  AOI22_X1 U10108 ( .A1(n7949), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7948), .B2(
        n9468), .ZN(n7740) );
  NAND2_X1 U10109 ( .A1(n7741), .A2(n7740), .ZN(n13104) );
  NAND2_X1 U10110 ( .A1(n6601), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7749) );
  INV_X1 U10111 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9440) );
  OR2_X1 U10112 ( .A1(n12049), .A2(n9440), .ZN(n7748) );
  INV_X1 U10113 ( .A(n7742), .ZN(n7758) );
  NAND2_X1 U10114 ( .A1(n7744), .A2(n7743), .ZN(n7745) );
  NAND2_X1 U10115 ( .A1(n7758), .A2(n7745), .ZN(n13105) );
  OR2_X1 U10116 ( .A1(n8094), .A2(n13105), .ZN(n7747) );
  INV_X1 U10117 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10611) );
  OR2_X1 U10118 ( .A1(n6614), .A2(n10611), .ZN(n7746) );
  NAND4_X1 U10119 ( .A1(n7749), .A2(n7748), .A3(n7747), .A4(n7746), .ZN(n13142) );
  INV_X1 U10120 ( .A(n12102), .ZN(n10234) );
  OR2_X1 U10121 ( .A1(n13104), .A2(n13142), .ZN(n7750) );
  NAND2_X1 U10122 ( .A1(n10231), .A2(n7750), .ZN(n10455) );
  NAND2_X1 U10123 ( .A1(n10325), .A2(n12059), .ZN(n7755) );
  NAND2_X1 U10124 ( .A1(n7767), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7753) );
  XNOR2_X1 U10125 ( .A(n7753), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13153) );
  AOI22_X1 U10126 ( .A1(n7949), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7948), .B2(
        n13153), .ZN(n7754) );
  NAND2_X1 U10127 ( .A1(n7755), .A2(n7754), .ZN(n11918) );
  NAND2_X1 U10128 ( .A1(n8093), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7763) );
  INV_X1 U10129 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7756) );
  OR2_X1 U10130 ( .A1(n8082), .A2(n7756), .ZN(n7762) );
  INV_X1 U10131 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7757) );
  NAND2_X1 U10132 ( .A1(n7758), .A2(n7757), .ZN(n7759) );
  NAND2_X1 U10133 ( .A1(n7775), .A2(n7759), .ZN(n14835) );
  OR2_X1 U10134 ( .A1(n8094), .A2(n14835), .ZN(n7761) );
  INV_X1 U10135 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9469) );
  OR2_X1 U10136 ( .A1(n6614), .A2(n9469), .ZN(n7760) );
  NAND4_X1 U10137 ( .A1(n7763), .A2(n7762), .A3(n7761), .A4(n7760), .ZN(n13141) );
  XNOR2_X1 U10138 ( .A(n11918), .B(n13141), .ZN(n12104) );
  INV_X1 U10139 ( .A(n12104), .ZN(n10454) );
  OR2_X1 U10140 ( .A1(n11918), .A2(n13141), .ZN(n7764) );
  NAND2_X1 U10141 ( .A1(n10310), .A2(n12059), .ZN(n7773) );
  NAND2_X1 U10142 ( .A1(n7770), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7768) );
  MUX2_X1 U10143 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7768), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n7769) );
  INV_X1 U10144 ( .A(n7769), .ZN(n7771) );
  NOR2_X1 U10145 ( .A1(n7771), .A2(n7784), .ZN(n13168) );
  AOI22_X1 U10146 ( .A1(n7949), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7948), .B2(
        n13168), .ZN(n7772) );
  NAND2_X1 U10147 ( .A1(n6441), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7780) );
  INV_X1 U10148 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10576) );
  OR2_X1 U10149 ( .A1(n6614), .A2(n10576), .ZN(n7779) );
  NAND2_X1 U10150 ( .A1(n7775), .A2(n7774), .ZN(n7776) );
  NAND2_X1 U10151 ( .A1(n7791), .A2(n7776), .ZN(n10571) );
  OR2_X1 U10152 ( .A1(n8094), .A2(n10571), .ZN(n7778) );
  INV_X1 U10153 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9444) );
  OR2_X1 U10154 ( .A1(n12049), .A2(n9444), .ZN(n7777) );
  NAND4_X1 U10155 ( .A1(n7780), .A2(n7779), .A3(n7778), .A4(n7777), .ZN(n13140) );
  NAND2_X1 U10156 ( .A1(n11923), .A2(n13140), .ZN(n7781) );
  XNOR2_X1 U10157 ( .A(n7783), .B(n7782), .ZN(n10474) );
  NAND2_X1 U10158 ( .A1(n10474), .A2(n12059), .ZN(n7787) );
  INV_X1 U10159 ( .A(n7784), .ZN(n7801) );
  NAND2_X1 U10160 ( .A1(n7801), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7785) );
  XNOR2_X1 U10161 ( .A(n7785), .B(P2_IR_REG_9__SCAN_IN), .ZN(n13186) );
  AOI22_X1 U10162 ( .A1(n7949), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7948), .B2(
        n13186), .ZN(n7786) );
  NAND2_X2 U10163 ( .A1(n7787), .A2(n7786), .ZN(n13492) );
  NAND2_X1 U10164 ( .A1(n8093), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7796) );
  INV_X1 U10165 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7788) );
  OR2_X1 U10166 ( .A1(n8082), .A2(n7788), .ZN(n7795) );
  INV_X1 U10167 ( .A(n7789), .ZN(n7807) );
  NAND2_X1 U10168 ( .A1(n7791), .A2(n7790), .ZN(n7792) );
  NAND2_X1 U10169 ( .A1(n7807), .A2(n7792), .ZN(n13488) );
  OR2_X1 U10170 ( .A1(n8094), .A2(n13488), .ZN(n7794) );
  INV_X1 U10171 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n13489) );
  OR2_X1 U10172 ( .A1(n6614), .A2(n13489), .ZN(n7793) );
  NAND4_X1 U10173 ( .A1(n7796), .A2(n7795), .A3(n7794), .A4(n7793), .ZN(n13139) );
  INV_X1 U10174 ( .A(n12106), .ZN(n10782) );
  NAND2_X1 U10175 ( .A1(n13492), .A2(n13139), .ZN(n7797) );
  NAND2_X1 U10176 ( .A1(n7798), .A2(n7797), .ZN(n10889) );
  NAND2_X1 U10177 ( .A1(n10739), .A2(n12059), .ZN(n7804) );
  NAND2_X1 U10178 ( .A1(n7816), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7802) );
  XNOR2_X1 U10179 ( .A(n7802), .B(P2_IR_REG_10__SCAN_IN), .ZN(n9476) );
  AOI22_X1 U10180 ( .A1(n7949), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n9476), 
        .B2(n7948), .ZN(n7803) );
  NAND2_X1 U10181 ( .A1(n6601), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7812) );
  INV_X1 U10182 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n13477) );
  OR2_X1 U10183 ( .A1(n6614), .A2(n13477), .ZN(n7811) );
  INV_X1 U10184 ( .A(n7805), .ZN(n7820) );
  INV_X1 U10185 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7806) );
  NAND2_X1 U10186 ( .A1(n7807), .A2(n7806), .ZN(n7808) );
  NAND2_X1 U10187 ( .A1(n7820), .A2(n7808), .ZN(n13476) );
  OR2_X1 U10188 ( .A1(n8094), .A2(n13476), .ZN(n7810) );
  INV_X1 U10189 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9450) );
  OR2_X1 U10190 ( .A1(n12049), .A2(n9450), .ZN(n7809) );
  NAND4_X1 U10191 ( .A1(n7812), .A2(n7811), .A3(n7810), .A4(n7809), .ZN(n13138) );
  XNOR2_X1 U10192 ( .A(n13479), .B(n13138), .ZN(n12107) );
  INV_X1 U10193 ( .A(n12107), .ZN(n8121) );
  NAND2_X1 U10194 ( .A1(n13479), .A2(n13138), .ZN(n7813) );
  XNOR2_X1 U10195 ( .A(n7814), .B(n7815), .ZN(n10826) );
  NAND2_X1 U10196 ( .A1(n10826), .A2(n12059), .ZN(n7819) );
  OAI21_X1 U10197 ( .B1(n7816), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7817) );
  XNOR2_X1 U10198 ( .A(n7817), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9645) );
  AOI22_X1 U10199 ( .A1(n9645), .A2(n7948), .B1(n7949), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n7818) );
  NAND2_X1 U10200 ( .A1(n6601), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7826) );
  INV_X1 U10201 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n15175) );
  NAND2_X1 U10202 ( .A1(n7820), .A2(n15175), .ZN(n7821) );
  NAND2_X1 U10203 ( .A1(n7844), .A2(n7821), .ZN(n10978) );
  OR2_X1 U10204 ( .A1(n8094), .A2(n10978), .ZN(n7825) );
  INV_X1 U10205 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10979) );
  OR2_X1 U10206 ( .A1(n6614), .A2(n10979), .ZN(n7824) );
  INV_X1 U10207 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7822) );
  OR2_X1 U10208 ( .A1(n12049), .A2(n7822), .ZN(n7823) );
  NAND4_X1 U10209 ( .A1(n7826), .A2(n7825), .A3(n7824), .A4(n7823), .ZN(n13137) );
  AND2_X1 U10210 ( .A1(n13600), .A2(n13137), .ZN(n7828) );
  OR2_X1 U10211 ( .A1(n13600), .A2(n13137), .ZN(n7827) );
  OR2_X1 U10212 ( .A1(n7830), .A2(n7829), .ZN(n7831) );
  NAND2_X1 U10213 ( .A1(n7832), .A2(n7831), .ZN(n10831) );
  NAND2_X1 U10214 ( .A1(n10831), .A2(n12059), .ZN(n7841) );
  INV_X1 U10215 ( .A(n7833), .ZN(n7834) );
  OAI21_X1 U10216 ( .B1(n7835), .B2(n7834), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7836) );
  MUX2_X1 U10217 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7836), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n7839) );
  INV_X1 U10218 ( .A(n7837), .ZN(n7838) );
  AND2_X1 U10219 ( .A1(n7839), .A2(n7838), .ZN(n9954) );
  AOI22_X1 U10220 ( .A1(n7949), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7948), 
        .B2(n9954), .ZN(n7840) );
  NAND2_X1 U10221 ( .A1(n8093), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7849) );
  INV_X1 U10222 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7842) );
  OR2_X1 U10223 ( .A1(n8082), .A2(n7842), .ZN(n7848) );
  NAND2_X1 U10224 ( .A1(n7844), .A2(n7843), .ZN(n7845) );
  NAND2_X1 U10225 ( .A1(n7860), .A2(n7845), .ZN(n11164) );
  OR2_X1 U10226 ( .A1(n8094), .A2(n11164), .ZN(n7847) );
  INV_X1 U10227 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11165) );
  OR2_X1 U10228 ( .A1(n6614), .A2(n11165), .ZN(n7846) );
  NAND4_X1 U10229 ( .A1(n7849), .A2(n7848), .A3(n7847), .A4(n7846), .ZN(n13136) );
  NAND2_X1 U10230 ( .A1(n7850), .A2(n13136), .ZN(n7852) );
  OR2_X1 U10231 ( .A1(n7854), .A2(n7853), .ZN(n7855) );
  NAND2_X1 U10232 ( .A1(n7856), .A2(n7855), .ZN(n11026) );
  NAND2_X1 U10233 ( .A1(n11026), .A2(n12059), .ZN(n7859) );
  OR2_X1 U10234 ( .A1(n7837), .A2(n7869), .ZN(n7857) );
  XNOR2_X1 U10235 ( .A(n7857), .B(P2_IR_REG_13__SCAN_IN), .ZN(n14805) );
  AOI22_X1 U10236 ( .A1(n7949), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7948), 
        .B2(n14805), .ZN(n7858) );
  NAND2_X1 U10237 ( .A1(n6601), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7866) );
  INV_X1 U10238 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11151) );
  OR2_X1 U10239 ( .A1(n6614), .A2(n11151), .ZN(n7865) );
  NAND2_X1 U10240 ( .A1(n7860), .A2(n11127), .ZN(n7861) );
  NAND2_X1 U10241 ( .A1(n7877), .A2(n7861), .ZN(n11150) );
  OR2_X1 U10242 ( .A1(n8094), .A2(n11150), .ZN(n7864) );
  INV_X1 U10243 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7862) );
  OR2_X1 U10244 ( .A1(n12049), .A2(n7862), .ZN(n7863) );
  NAND4_X1 U10245 ( .A1(n7866), .A2(n7865), .A3(n7864), .A4(n7863), .ZN(n13135) );
  NAND2_X1 U10246 ( .A1(n7867), .A2(n9302), .ZN(n7886) );
  OR2_X1 U10247 ( .A1(n7867), .A2(n9302), .ZN(n7868) );
  NAND2_X1 U10248 ( .A1(n7886), .A2(n7868), .ZN(n7889) );
  XNOR2_X1 U10249 ( .A(n7889), .B(n7888), .ZN(n11032) );
  NAND2_X1 U10250 ( .A1(n11032), .A2(n12059), .ZN(n7873) );
  OR2_X1 U10251 ( .A1(n7870), .A2(n7869), .ZN(n7871) );
  XNOR2_X1 U10252 ( .A(n7871), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10402) );
  AOI22_X1 U10253 ( .A1(n7949), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7948), 
        .B2(n10402), .ZN(n7872) );
  NAND2_X1 U10254 ( .A1(n8022), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7882) );
  INV_X1 U10255 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7874) );
  OR2_X1 U10256 ( .A1(n8082), .A2(n7874), .ZN(n7881) );
  INV_X1 U10257 ( .A(n7875), .ZN(n7897) );
  NAND2_X1 U10258 ( .A1(n7877), .A2(n7876), .ZN(n7878) );
  NAND2_X1 U10259 ( .A1(n7897), .A2(n7878), .ZN(n13467) );
  OR2_X1 U10260 ( .A1(n8094), .A2(n13467), .ZN(n7880) );
  INV_X1 U10261 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10415) );
  OR2_X1 U10262 ( .A1(n12049), .A2(n10415), .ZN(n7879) );
  NAND4_X1 U10263 ( .A1(n7882), .A2(n7881), .A3(n7880), .A4(n7879), .ZN(n13134) );
  NOR2_X1 U10264 ( .A1(n13589), .A2(n13134), .ZN(n7884) );
  NAND2_X1 U10265 ( .A1(n13589), .A2(n13134), .ZN(n7883) );
  AND2_X1 U10266 ( .A1(n7886), .A2(n7885), .ZN(n7887) );
  OAI21_X1 U10267 ( .B1(n7889), .B2(n7888), .A(n7887), .ZN(n7891) );
  NAND2_X1 U10268 ( .A1(n7891), .A2(n7890), .ZN(n11173) );
  NAND2_X1 U10269 ( .A1(n11173), .A2(n12059), .ZN(n7895) );
  NAND2_X1 U10270 ( .A1(n7892), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7893) );
  XNOR2_X1 U10271 ( .A(n7893), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14821) );
  AOI22_X1 U10272 ( .A1(n7949), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7948), 
        .B2(n14821), .ZN(n7894) );
  INV_X1 U10273 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7896) );
  NAND2_X1 U10274 ( .A1(n7897), .A2(n7896), .ZN(n7898) );
  NAND2_X1 U10275 ( .A1(n7910), .A2(n7898), .ZN(n13444) );
  OR2_X1 U10276 ( .A1(n13444), .A2(n8094), .ZN(n7902) );
  INV_X1 U10277 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n13638) );
  OR2_X1 U10278 ( .A1(n8082), .A2(n13638), .ZN(n7901) );
  INV_X1 U10279 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n13585) );
  OR2_X1 U10280 ( .A1(n12049), .A2(n13585), .ZN(n7900) );
  INV_X1 U10281 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n13445) );
  OR2_X1 U10282 ( .A1(n6614), .A2(n13445), .ZN(n7899) );
  NAND4_X1 U10283 ( .A1(n7902), .A2(n7901), .A3(n7900), .A4(n7899), .ZN(n13425) );
  INV_X1 U10284 ( .A(n13425), .ZN(n13461) );
  XNOR2_X1 U10285 ( .A(n13580), .B(n13461), .ZN(n13440) );
  INV_X1 U10286 ( .A(n13440), .ZN(n13447) );
  XNOR2_X1 U10287 ( .A(n7904), .B(n7903), .ZN(n11273) );
  NAND2_X1 U10288 ( .A1(n11273), .A2(n12059), .ZN(n7908) );
  NAND2_X1 U10289 ( .A1(n6567), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7905) );
  MUX2_X1 U10290 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7905), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n7906) );
  AOI22_X1 U10291 ( .A1(n7949), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7948), 
        .B2(n10628), .ZN(n7907) );
  NAND2_X1 U10292 ( .A1(n7910), .A2(n7909), .ZN(n7911) );
  NAND2_X1 U10293 ( .A1(n7925), .A2(n7911), .ZN(n13431) );
  NAND2_X1 U10294 ( .A1(n6601), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7913) );
  NAND2_X1 U10295 ( .A1(n8022), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7912) );
  AND2_X1 U10296 ( .A1(n7913), .A2(n7912), .ZN(n7915) );
  NAND2_X1 U10297 ( .A1(n8093), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7914) );
  OAI211_X1 U10298 ( .C1(n13431), .C2(n8094), .A(n7915), .B(n7914), .ZN(n13133) );
  INV_X1 U10299 ( .A(n13133), .ZN(n8129) );
  XNOR2_X1 U10300 ( .A(n13577), .B(n8129), .ZN(n13419) );
  NAND2_X1 U10301 ( .A1(n13577), .A2(n13133), .ZN(n7916) );
  NAND2_X1 U10302 ( .A1(n13418), .A2(n7916), .ZN(n13403) );
  XNOR2_X1 U10303 ( .A(n7917), .B(SI_17_), .ZN(n7918) );
  XNOR2_X1 U10304 ( .A(n7919), .B(n7918), .ZN(n11297) );
  NAND2_X1 U10305 ( .A1(n11297), .A2(n12059), .ZN(n7922) );
  NAND2_X1 U10306 ( .A1(n7935), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7920) );
  XNOR2_X1 U10307 ( .A(n7920), .B(P2_IR_REG_17__SCAN_IN), .ZN(n10631) );
  AOI22_X1 U10308 ( .A1(n7949), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7948), 
        .B2(n10631), .ZN(n7921) );
  INV_X1 U10309 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13407) );
  INV_X1 U10310 ( .A(n7923), .ZN(n7954) );
  NAND2_X1 U10311 ( .A1(n7925), .A2(n7924), .ZN(n7926) );
  NAND2_X1 U10312 ( .A1(n7954), .A2(n7926), .ZN(n13406) );
  OR2_X1 U10313 ( .A1(n13406), .A2(n8094), .ZN(n7928) );
  AOI22_X1 U10314 ( .A1(n8093), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n6601), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n7927) );
  OAI211_X1 U10315 ( .C1(n6614), .C2(n13407), .A(n7928), .B(n7927), .ZN(n13428) );
  INV_X1 U10316 ( .A(n13428), .ZN(n13388) );
  XNOR2_X1 U10317 ( .A(n13634), .B(n13388), .ZN(n13411) );
  NAND2_X1 U10318 ( .A1(n13403), .A2(n13411), .ZN(n7930) );
  NAND2_X1 U10319 ( .A1(n13634), .A2(n13428), .ZN(n7929) );
  NAND2_X1 U10320 ( .A1(n7930), .A2(n7929), .ZN(n13379) );
  NAND2_X1 U10321 ( .A1(n7932), .A2(n7931), .ZN(n7933) );
  NAND2_X1 U10322 ( .A1(n7934), .A2(n7933), .ZN(n11496) );
  OR2_X1 U10323 ( .A1(n11496), .A2(n6636), .ZN(n7939) );
  OR2_X1 U10324 ( .A1(n7935), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U10325 ( .A1(n7936), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7937) );
  XNOR2_X1 U10326 ( .A(n7937), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13199) );
  AOI22_X1 U10327 ( .A1(n13199), .A2(n7948), .B1(n7949), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n7938) );
  XNOR2_X1 U10328 ( .A(n7954), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n13396) );
  INV_X1 U10329 ( .A(n8094), .ZN(n7989) );
  NAND2_X1 U10330 ( .A1(n13396), .A2(n7989), .ZN(n7944) );
  INV_X1 U10331 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13197) );
  NAND2_X1 U10332 ( .A1(n6601), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7941) );
  NAND2_X1 U10333 ( .A1(n8022), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7940) );
  OAI211_X1 U10334 ( .C1(n12049), .C2(n13197), .A(n7941), .B(n7940), .ZN(n7942) );
  INV_X1 U10335 ( .A(n7942), .ZN(n7943) );
  NAND2_X1 U10336 ( .A1(n7944), .A2(n7943), .ZN(n13132) );
  INV_X1 U10337 ( .A(n13132), .ZN(n8134) );
  XNOR2_X1 U10338 ( .A(n13562), .B(n8134), .ZN(n13384) );
  INV_X1 U10339 ( .A(n13384), .ZN(n13380) );
  OR2_X1 U10340 ( .A1(n13562), .A2(n13132), .ZN(n7945) );
  XNOR2_X1 U10341 ( .A(n7947), .B(n7946), .ZN(n11500) );
  NAND2_X1 U10342 ( .A1(n11500), .A2(n12059), .ZN(n7951) );
  AOI22_X1 U10343 ( .A1(n7949), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6689), 
        .B2(n7948), .ZN(n7950) );
  INV_X1 U10344 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7953) );
  INV_X1 U10345 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7952) );
  OAI21_X1 U10346 ( .B1(n7954), .B2(n7953), .A(n7952), .ZN(n7956) );
  INV_X1 U10347 ( .A(n7955), .ZN(n7971) );
  AND2_X1 U10348 ( .A1(n7956), .A2(n7971), .ZN(n13372) );
  NAND2_X1 U10349 ( .A1(n13372), .A2(n7989), .ZN(n7962) );
  INV_X1 U10350 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n7959) );
  NAND2_X1 U10351 ( .A1(n8022), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n7958) );
  NAND2_X1 U10352 ( .A1(n6601), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n7957) );
  OAI211_X1 U10353 ( .C1(n12049), .C2(n7959), .A(n7958), .B(n7957), .ZN(n7960)
         );
  INV_X1 U10354 ( .A(n7960), .ZN(n7961) );
  NAND2_X1 U10355 ( .A1(n7962), .A2(n7961), .ZN(n13386) );
  NAND2_X1 U10356 ( .A1(n13559), .A2(n13386), .ZN(n12115) );
  OR2_X1 U10357 ( .A1(n13559), .A2(n13386), .ZN(n12116) );
  NAND2_X1 U10358 ( .A1(n7963), .A2(n12116), .ZN(n13348) );
  NAND2_X1 U10359 ( .A1(n7965), .A2(n7964), .ZN(n7966) );
  NAND2_X1 U10360 ( .A1(n7967), .A2(n7966), .ZN(n11514) );
  OR2_X1 U10361 ( .A1(n11514), .A2(n6636), .ZN(n7969) );
  OR2_X1 U10362 ( .A1(n12061), .A2(n10866), .ZN(n7968) );
  INV_X1 U10363 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7970) );
  NAND2_X1 U10364 ( .A1(n7971), .A2(n7970), .ZN(n7972) );
  NAND2_X1 U10365 ( .A1(n7987), .A2(n7972), .ZN(n13355) );
  OR2_X1 U10366 ( .A1(n13355), .A2(n8094), .ZN(n7978) );
  INV_X1 U10367 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n7975) );
  NAND2_X1 U10368 ( .A1(n6601), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n7974) );
  NAND2_X1 U10369 ( .A1(n8022), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n7973) );
  OAI211_X1 U10370 ( .C1(n7975), .C2(n12049), .A(n7974), .B(n7973), .ZN(n7976)
         );
  INV_X1 U10371 ( .A(n7976), .ZN(n7977) );
  NAND2_X1 U10372 ( .A1(n7978), .A2(n7977), .ZN(n13131) );
  NAND2_X1 U10373 ( .A1(n13553), .A2(n13131), .ZN(n7979) );
  NAND2_X1 U10374 ( .A1(n13348), .A2(n7979), .ZN(n7981) );
  OR2_X1 U10375 ( .A1(n13553), .A2(n13131), .ZN(n7980) );
  NAND2_X1 U10376 ( .A1(n7981), .A2(n7980), .ZN(n13336) );
  OR2_X1 U10377 ( .A1(n6555), .A2(n7983), .ZN(n7984) );
  NAND2_X1 U10378 ( .A1(n7982), .A2(n7984), .ZN(n11527) );
  OR2_X1 U10379 ( .A1(n11527), .A2(n6636), .ZN(n7986) );
  INV_X1 U10380 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11111) );
  OR2_X1 U10381 ( .A1(n12061), .A2(n11111), .ZN(n7985) );
  NAND2_X1 U10382 ( .A1(n7987), .A2(n13024), .ZN(n7988) );
  AND2_X1 U10383 ( .A1(n8004), .A2(n7988), .ZN(n13343) );
  NAND2_X1 U10384 ( .A1(n13343), .A2(n7989), .ZN(n7995) );
  INV_X1 U10385 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n7992) );
  NAND2_X1 U10386 ( .A1(n6601), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7991) );
  NAND2_X1 U10387 ( .A1(n8022), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7990) );
  OAI211_X1 U10388 ( .C1(n12049), .C2(n7992), .A(n7991), .B(n7990), .ZN(n7993)
         );
  INV_X1 U10389 ( .A(n7993), .ZN(n7994) );
  NAND2_X1 U10390 ( .A1(n7995), .A2(n7994), .ZN(n13353) );
  XNOR2_X1 U10391 ( .A(n13549), .B(n13353), .ZN(n13338) );
  INV_X1 U10392 ( .A(n13338), .ZN(n7996) );
  NAND2_X1 U10393 ( .A1(n13336), .A2(n7996), .ZN(n7998) );
  INV_X1 U10394 ( .A(n13353), .ZN(n13071) );
  NAND2_X1 U10395 ( .A1(n6918), .A2(n13071), .ZN(n7997) );
  NAND2_X1 U10396 ( .A1(n11543), .A2(n8000), .ZN(n8001) );
  NAND2_X1 U10397 ( .A1(n8014), .A2(n8001), .ZN(n11268) );
  OR2_X1 U10398 ( .A1(n12061), .A2(n11269), .ZN(n8002) );
  AND2_X1 U10399 ( .A1(n8004), .A2(n13081), .ZN(n8005) );
  OR2_X1 U10400 ( .A1(n8005), .A2(n8019), .ZN(n13329) );
  INV_X1 U10401 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8008) );
  NAND2_X1 U10402 ( .A1(n6601), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8007) );
  NAND2_X1 U10403 ( .A1(n8022), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8006) );
  OAI211_X1 U10404 ( .C1(n12049), .C2(n8008), .A(n8007), .B(n8006), .ZN(n8009)
         );
  INV_X1 U10405 ( .A(n8009), .ZN(n8010) );
  OAI21_X1 U10406 ( .B1(n13329), .B2(n8094), .A(n8010), .ZN(n13130) );
  INV_X1 U10407 ( .A(n13130), .ZN(n8011) );
  INV_X1 U10408 ( .A(n12119), .ZN(n13323) );
  NAND2_X1 U10409 ( .A1(n13626), .A2(n13130), .ZN(n8012) );
  NAND2_X1 U10410 ( .A1(n14273), .A2(n12059), .ZN(n8018) );
  INV_X1 U10411 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n13672) );
  OR2_X1 U10412 ( .A1(n12061), .A2(n13672), .ZN(n8017) );
  OR2_X1 U10413 ( .A1(n8019), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8021) );
  NAND2_X1 U10414 ( .A1(n8021), .A2(n8020), .ZN(n13306) );
  OR2_X1 U10415 ( .A1(n13306), .A2(n8094), .ZN(n8027) );
  INV_X1 U10416 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n13540) );
  NAND2_X1 U10417 ( .A1(n6601), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8024) );
  NAND2_X1 U10418 ( .A1(n8022), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8023) );
  OAI211_X1 U10419 ( .C1(n12049), .C2(n13540), .A(n8024), .B(n8023), .ZN(n8025) );
  INV_X1 U10420 ( .A(n8025), .ZN(n8026) );
  NAND2_X1 U10421 ( .A1(n8027), .A2(n8026), .ZN(n13129) );
  OR2_X1 U10422 ( .A1(n13313), .A2(n13129), .ZN(n8028) );
  NAND2_X1 U10423 ( .A1(n8030), .A2(n8029), .ZN(n8031) );
  NAND2_X1 U10424 ( .A1(n8032), .A2(n8031), .ZN(n11581) );
  OR2_X1 U10425 ( .A1(n11581), .A2(n6636), .ZN(n8035) );
  OR2_X1 U10426 ( .A1(n12061), .A2(n11270), .ZN(n8034) );
  NAND2_X1 U10427 ( .A1(n6601), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8040) );
  INV_X1 U10428 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n13535) );
  OR2_X1 U10429 ( .A1(n12049), .A2(n13535), .ZN(n8039) );
  OAI21_X1 U10430 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n8036), .A(n8048), .ZN(
        n13291) );
  OR2_X1 U10431 ( .A1(n8094), .A2(n13291), .ZN(n8038) );
  INV_X1 U10432 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13292) );
  OR2_X1 U10433 ( .A1(n6614), .A2(n13292), .ZN(n8037) );
  NAND4_X1 U10434 ( .A1(n8040), .A2(n8039), .A3(n8038), .A4(n8037), .ZN(n13128) );
  INV_X1 U10435 ( .A(n13128), .ZN(n13032) );
  NAND2_X1 U10436 ( .A1(n13529), .A2(n13032), .ZN(n8149) );
  OR2_X1 U10437 ( .A1(n13529), .A2(n13032), .ZN(n8041) );
  NAND2_X1 U10438 ( .A1(n13290), .A2(n13295), .ZN(n8043) );
  NAND2_X1 U10439 ( .A1(n13529), .A2(n13128), .ZN(n8042) );
  XNOR2_X1 U10440 ( .A(n8045), .B(n8044), .ZN(n13664) );
  NAND2_X1 U10441 ( .A1(n13664), .A2(n12059), .ZN(n8047) );
  INV_X1 U10442 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13667) );
  OR2_X1 U10443 ( .A1(n12061), .A2(n13667), .ZN(n8046) );
  NAND2_X1 U10444 ( .A1(n6601), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8054) );
  INV_X1 U10445 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n15221) );
  OR2_X1 U10446 ( .A1(n12049), .A2(n15221), .ZN(n8053) );
  INV_X1 U10447 ( .A(n8048), .ZN(n8050) );
  INV_X1 U10448 ( .A(n8065), .ZN(n8049) );
  OAI21_X1 U10449 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n8050), .A(n8049), .ZN(
        n13282) );
  OR2_X1 U10450 ( .A1(n8094), .A2(n13282), .ZN(n8052) );
  INV_X1 U10451 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13283) );
  OR2_X1 U10452 ( .A1(n6614), .A2(n13283), .ZN(n8051) );
  NAND4_X1 U10453 ( .A1(n8054), .A2(n8053), .A3(n8052), .A4(n8051), .ZN(n13127) );
  AND2_X1 U10454 ( .A1(n13525), .A2(n13127), .ZN(n8055) );
  OR2_X1 U10455 ( .A1(n13525), .A2(n13127), .ZN(n8056) );
  XNOR2_X1 U10456 ( .A(n8058), .B(SI_26_), .ZN(n8059) );
  NAND2_X1 U10457 ( .A1(n13661), .A2(n12059), .ZN(n8062) );
  OR2_X1 U10458 ( .A1(n12061), .A2(n13662), .ZN(n8061) );
  NAND2_X1 U10459 ( .A1(n6601), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8069) );
  INV_X1 U10460 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8063) );
  OR2_X1 U10461 ( .A1(n12049), .A2(n8063), .ZN(n8068) );
  OAI21_X1 U10462 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(n8065), .A(n8064), .ZN(
        n13267) );
  OR2_X1 U10463 ( .A1(n8094), .A2(n13267), .ZN(n8067) );
  INV_X1 U10464 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13268) );
  OR2_X1 U10465 ( .A1(n6614), .A2(n13268), .ZN(n8066) );
  NAND4_X1 U10466 ( .A1(n8069), .A2(n8068), .A3(n8067), .A4(n8066), .ZN(n13245) );
  INV_X1 U10467 ( .A(n13245), .ZN(n13031) );
  XNOR2_X1 U10468 ( .A(n13520), .B(n13031), .ZN(n12123) );
  OR2_X1 U10469 ( .A1(n13520), .A2(n13245), .ZN(n8070) );
  NAND2_X1 U10470 ( .A1(n13514), .A2(n13126), .ZN(n8072) );
  INV_X1 U10471 ( .A(n8073), .ZN(n8074) );
  NAND2_X1 U10472 ( .A1(n8075), .A2(n8074), .ZN(n8076) );
  XNOR2_X1 U10473 ( .A(n8078), .B(SI_28_), .ZN(n8079) );
  INV_X1 U10474 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13657) );
  OR2_X1 U10475 ( .A1(n12061), .A2(n13657), .ZN(n8081) );
  NAND2_X1 U10476 ( .A1(n8093), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8090) );
  INV_X1 U10477 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n15133) );
  OR2_X1 U10478 ( .A1(n8082), .A2(n15133), .ZN(n8089) );
  INV_X1 U10479 ( .A(n8085), .ZN(n8083) );
  NAND2_X1 U10480 ( .A1(n8083), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n11724) );
  INV_X1 U10481 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8084) );
  NAND2_X1 U10482 ( .A1(n8085), .A2(n8084), .ZN(n8086) );
  NAND2_X1 U10483 ( .A1(n11724), .A2(n8086), .ZN(n13239) );
  OR2_X1 U10484 ( .A1(n8094), .A2(n13239), .ZN(n8088) );
  INV_X1 U10485 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n15186) );
  OR2_X1 U10486 ( .A1(n6614), .A2(n15186), .ZN(n8087) );
  NAND4_X1 U10487 ( .A1(n8090), .A2(n8089), .A3(n8088), .A4(n8087), .ZN(n13244) );
  NAND2_X1 U10488 ( .A1(n13512), .A2(n13244), .ZN(n8092) );
  OR2_X1 U10489 ( .A1(n13512), .A2(n13244), .ZN(n8091) );
  INV_X1 U10490 ( .A(n13233), .ZN(n13228) );
  NAND2_X1 U10491 ( .A1(n13231), .A2(n8092), .ZN(n8099) );
  NAND2_X1 U10492 ( .A1(n8093), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8098) );
  NAND2_X1 U10493 ( .A1(n6601), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8097) );
  OR2_X1 U10494 ( .A1(n8094), .A2(n11724), .ZN(n8096) );
  INV_X1 U10495 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n11725) );
  OR2_X1 U10496 ( .A1(n6614), .A2(n11725), .ZN(n8095) );
  NAND4_X1 U10497 ( .A1(n8098), .A2(n8097), .A3(n8096), .A4(n8095), .ZN(n13125) );
  XNOR2_X1 U10498 ( .A(n12037), .B(n13125), .ZN(n12124) );
  INV_X1 U10499 ( .A(n12091), .ZN(n12097) );
  NOR2_X1 U10500 ( .A1(n13312), .A2(n12097), .ZN(n8100) );
  NAND2_X1 U10501 ( .A1(n8100), .A2(n11882), .ZN(n14876) );
  INV_X1 U10502 ( .A(n13525), .ZN(n8104) );
  INV_X1 U10503 ( .A(n13626), .ZN(n8145) );
  NAND2_X1 U10504 ( .A1(n11880), .A2(n6635), .ZN(n10285) );
  INV_X1 U10505 ( .A(n11923), .ZN(n10572) );
  NAND2_X1 U10506 ( .A1(n10502), .A2(n10572), .ZN(n10779) );
  INV_X1 U10507 ( .A(n13600), .ZN(n10975) );
  NOR2_X1 U10508 ( .A1(n13450), .A2(n13577), .ZN(n13435) );
  INV_X1 U10509 ( .A(n13634), .ZN(n13405) );
  NAND2_X1 U10510 ( .A1(n13435), .A2(n13405), .ZN(n13404) );
  NOR2_X2 U10511 ( .A1(n13394), .A2(n13559), .ZN(n13358) );
  INV_X1 U10512 ( .A(n13553), .ZN(n8103) );
  NAND2_X1 U10513 ( .A1(n8104), .A2(n13293), .ZN(n13275) );
  OR2_X1 U10514 ( .A1(n13275), .A2(n13520), .ZN(n13247) );
  AOI21_X1 U10515 ( .B1(n13238), .B2(n12037), .A(n13465), .ZN(n8105) );
  INV_X1 U10516 ( .A(n12037), .ZN(n8774) );
  NAND2_X1 U10517 ( .A1(n8105), .A2(n13221), .ZN(n11726) );
  INV_X1 U10518 ( .A(n13244), .ZN(n13001) );
  INV_X1 U10519 ( .A(n11883), .ZN(n8106) );
  NAND2_X1 U10520 ( .A1(n10293), .A2(n11885), .ZN(n8107) );
  NAND2_X1 U10521 ( .A1(n9832), .A2(n8107), .ZN(n10292) );
  NAND2_X1 U10522 ( .A1(n10292), .A2(n12095), .ZN(n10291) );
  NAND2_X1 U10523 ( .A1(n10133), .A2(n11890), .ZN(n8108) );
  INV_X1 U10524 ( .A(n12098), .ZN(n10020) );
  NAND2_X1 U10525 ( .A1(n10021), .A2(n10020), .ZN(n10019) );
  NAND2_X1 U10526 ( .A1(n10587), .A2(n15068), .ZN(n8109) );
  NAND2_X1 U10527 ( .A1(n10432), .A2(n14872), .ZN(n8110) );
  OR2_X1 U10528 ( .A1(n10586), .A2(n11908), .ZN(n8111) );
  NAND2_X1 U10529 ( .A1(n11908), .A2(n10586), .ZN(n8112) );
  NAND2_X1 U10530 ( .A1(n8113), .A2(n8112), .ZN(n10235) );
  INV_X1 U10531 ( .A(n13142), .ZN(n10431) );
  NAND2_X1 U10532 ( .A1(n13104), .A2(n10431), .ZN(n8114) );
  INV_X1 U10533 ( .A(n13141), .ZN(n8115) );
  OR2_X1 U10534 ( .A1(n11918), .A2(n8115), .ZN(n8116) );
  INV_X1 U10535 ( .A(n13140), .ZN(n8118) );
  OR2_X1 U10536 ( .A1(n11923), .A2(n8118), .ZN(n8119) );
  INV_X1 U10537 ( .A(n13139), .ZN(n8120) );
  INV_X1 U10538 ( .A(n13138), .ZN(n8122) );
  OR2_X1 U10539 ( .A1(n13479), .A2(n8122), .ZN(n8123) );
  NAND2_X1 U10540 ( .A1(n10894), .A2(n8123), .ZN(n10972) );
  INV_X1 U10541 ( .A(n13137), .ZN(n11160) );
  XNOR2_X1 U10542 ( .A(n13600), .B(n11160), .ZN(n12111) );
  NAND2_X1 U10543 ( .A1(n13600), .A2(n11160), .ZN(n8124) );
  INV_X1 U10544 ( .A(n13136), .ZN(n11128) );
  AND2_X1 U10545 ( .A1(n11944), .A2(n11128), .ZN(n8125) );
  INV_X1 U10546 ( .A(n13135), .ZN(n13463) );
  XNOR2_X1 U10547 ( .A(n13645), .B(n13463), .ZN(n12112) );
  INV_X1 U10548 ( .A(n12112), .ZN(n8126) );
  INV_X1 U10549 ( .A(n13134), .ZN(n12093) );
  OR2_X1 U10550 ( .A1(n13580), .A2(n13461), .ZN(n8127) );
  NAND2_X1 U10551 ( .A1(n8128), .A2(n8127), .ZN(n13423) );
  INV_X1 U10552 ( .A(n13419), .ZN(n13424) );
  NAND2_X1 U10553 ( .A1(n13423), .A2(n13424), .ZN(n13422) );
  OR2_X1 U10554 ( .A1(n13577), .A2(n8129), .ZN(n8130) );
  NAND2_X1 U10555 ( .A1(n13634), .A2(n13388), .ZN(n8131) );
  NAND2_X1 U10556 ( .A1(n13412), .A2(n8131), .ZN(n8133) );
  OR2_X1 U10557 ( .A1(n13634), .A2(n13388), .ZN(n8132) );
  NAND2_X1 U10558 ( .A1(n8133), .A2(n8132), .ZN(n13385) );
  NOR2_X1 U10559 ( .A1(n13562), .A2(n8134), .ZN(n8136) );
  NAND2_X1 U10560 ( .A1(n13562), .A2(n8134), .ZN(n8135) );
  INV_X1 U10561 ( .A(n13386), .ZN(n13094) );
  OR2_X1 U10562 ( .A1(n13559), .A2(n13094), .ZN(n8137) );
  NAND2_X1 U10563 ( .A1(n13367), .A2(n8137), .ZN(n8139) );
  NAND2_X1 U10564 ( .A1(n13559), .A2(n13094), .ZN(n8138) );
  NAND2_X1 U10565 ( .A1(n8139), .A2(n8138), .ZN(n13351) );
  INV_X1 U10566 ( .A(n13131), .ZN(n8140) );
  AND2_X1 U10567 ( .A1(n13553), .A2(n8140), .ZN(n13337) );
  OAI22_X1 U10568 ( .A1(n13549), .A2(n13071), .B1(n8140), .B2(n13553), .ZN(
        n8141) );
  INV_X1 U10569 ( .A(n8141), .ZN(n8142) );
  NAND2_X1 U10570 ( .A1(n13549), .A2(n13071), .ZN(n8143) );
  NAND2_X1 U10571 ( .A1(n8145), .A2(n13130), .ZN(n8146) );
  INV_X1 U10572 ( .A(n13129), .ZN(n8147) );
  NAND2_X1 U10573 ( .A1(n13313), .A2(n8147), .ZN(n8148) );
  XNOR2_X1 U10574 ( .A(n13525), .B(n13127), .ZN(n13285) );
  NAND2_X1 U10575 ( .A1(n13278), .A2(n13285), .ZN(n8151) );
  INV_X1 U10576 ( .A(n13127), .ZN(n13115) );
  NAND2_X1 U10577 ( .A1(n13525), .A2(n13115), .ZN(n8150) );
  NAND2_X1 U10578 ( .A1(n8151), .A2(n8150), .ZN(n13263) );
  NAND2_X1 U10579 ( .A1(n13263), .A2(n13269), .ZN(n8153) );
  NAND2_X1 U10580 ( .A1(n13520), .A2(n13031), .ZN(n8152) );
  NAND2_X1 U10581 ( .A1(n8153), .A2(n8152), .ZN(n13243) );
  INV_X1 U10582 ( .A(n13126), .ZN(n13114) );
  AND2_X1 U10583 ( .A1(n13514), .A2(n13114), .ZN(n8154) );
  OAI21_X1 U10584 ( .B1(n13001), .B2(n13512), .A(n13232), .ZN(n8156) );
  XNOR2_X1 U10585 ( .A(n8156), .B(n8155), .ZN(n8166) );
  OR2_X1 U10586 ( .A1(n11882), .A2(n13312), .ZN(n12065) );
  OR2_X1 U10587 ( .A1(n7508), .A2(n12091), .ZN(n8157) );
  INV_X1 U10588 ( .A(n9481), .ZN(n8159) );
  INV_X1 U10589 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n15189) );
  INV_X1 U10590 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n13224) );
  OR2_X1 U10591 ( .A1(n6614), .A2(n13224), .ZN(n8161) );
  NAND2_X1 U10592 ( .A1(n6601), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8160) );
  OAI211_X1 U10593 ( .C1(n12049), .C2(n15189), .A(n8161), .B(n8160), .ZN(
        n13124) );
  OR2_X1 U10594 ( .A1(n13658), .A2(n8162), .ZN(n8163) );
  AND2_X1 U10595 ( .A1(n13427), .A2(n8163), .ZN(n13217) );
  AOI22_X1 U10596 ( .A1(n13426), .A2(n13244), .B1(n13124), .B2(n13217), .ZN(
        n8164) );
  NAND2_X1 U10597 ( .A1(n8771), .A2(n14885), .ZN(n8169) );
  INV_X1 U10598 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8167) );
  OR2_X1 U10599 ( .A1(n14885), .A2(n8167), .ZN(n8168) );
  INV_X1 U10600 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n8750) );
  XNOR2_X2 U10601 ( .A(n8182), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8188) );
  INV_X1 U10602 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n8186) );
  OR2_X1 U10603 ( .A1(n6447), .A2(n8186), .ZN(n8194) );
  NAND2_X4 U10604 ( .A1(n8189), .A2(n8188), .ZN(n8904) );
  INV_X1 U10605 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n8190) );
  OR2_X1 U10606 ( .A1(n8904), .A2(n8190), .ZN(n8192) );
  NAND2_X1 U10607 ( .A1(n8659), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8191) );
  INV_X1 U10608 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9624) );
  NAND2_X1 U10609 ( .A1(n9624), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8196) );
  AND2_X1 U10610 ( .A1(n8221), .A2(n8196), .ZN(n8197) );
  INV_X1 U10611 ( .A(SI_0_), .ZN(n9625) );
  MUX2_X1 U10612 ( .A(n8197), .B(n9625), .S(n11542), .Z(n9193) );
  NAND2_X1 U10613 ( .A1(n8200), .A2(n8199), .ZN(n8204) );
  INV_X1 U10614 ( .A(n8204), .ZN(n8201) );
  XNOR2_X1 U10615 ( .A(P3_IR_REG_31__SCAN_IN), .B(P3_IR_REG_28__SCAN_IN), .ZN(
        n8202) );
  OAI21_X1 U10616 ( .B1(n8204), .B2(n8203), .A(n8202), .ZN(n8205) );
  MUX2_X1 U10617 ( .A(n15107), .B(n9193), .S(n9753), .Z(n14892) );
  NAND2_X1 U10618 ( .A1(n10393), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8211) );
  INV_X1 U10619 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n9774) );
  OR2_X1 U10620 ( .A1(n8267), .A2(n9774), .ZN(n8210) );
  INV_X1 U10621 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8206) );
  XNOR2_X1 U10622 ( .A(n8221), .B(n8223), .ZN(n9257) );
  NOR2_X1 U10623 ( .A1(n9753), .A2(n9778), .ZN(n8212) );
  INV_X1 U10624 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10308) );
  INV_X1 U10625 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n8215) );
  NAND2_X1 U10626 ( .A1(n8659), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8217) );
  INV_X1 U10627 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9923) );
  OR2_X1 U10628 ( .A1(n6448), .A2(n9923), .ZN(n8216) );
  XNOR2_X2 U10629 ( .A(n8220), .B(P3_IR_REG_2__SCAN_IN), .ZN(n9931) );
  INV_X1 U10630 ( .A(n8221), .ZN(n8222) );
  NAND2_X1 U10631 ( .A1(n8223), .A2(n8222), .ZN(n8225) );
  NAND2_X1 U10632 ( .A1(n9212), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8224) );
  XNOR2_X1 U10633 ( .A(n8233), .B(n8234), .ZN(n9227) );
  INV_X1 U10634 ( .A(SI_2_), .ZN(n8226) );
  NAND2_X1 U10635 ( .A1(n8227), .A2(n8226), .ZN(n8228) );
  OAI211_X1 U10636 ( .C1(n9931), .C2(n9753), .A(n8229), .B(n8228), .ZN(n8789)
         );
  NAND2_X1 U10637 ( .A1(n8231), .A2(n8230), .ZN(n12340) );
  NAND2_X1 U10638 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6494), .ZN(n8232) );
  XNOR2_X1 U10639 ( .A(n8232), .B(P3_IR_REG_3__SCAN_IN), .ZN(n11325) );
  XNOR2_X1 U10640 ( .A(n8255), .B(n8254), .ZN(n11326) );
  OR2_X1 U10641 ( .A1(n12281), .A2(n11326), .ZN(n8237) );
  OR2_X1 U10642 ( .A1(n8258), .A2(SI_3_), .ZN(n8236) );
  OAI211_X1 U10643 ( .C1(n11325), .C2(n9753), .A(n8237), .B(n8236), .ZN(n10354) );
  INV_X1 U10644 ( .A(n10354), .ZN(n15006) );
  INV_X4 U10645 ( .A(n8238), .ZN(n8659) );
  NAND2_X1 U10646 ( .A1(n8659), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8242) );
  NAND2_X1 U10647 ( .A1(n8592), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8241) );
  INV_X1 U10648 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10563) );
  OR2_X1 U10649 ( .A1(n8245), .A2(n10563), .ZN(n8240) );
  OR2_X1 U10650 ( .A1(n8904), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8239) );
  NAND2_X1 U10651 ( .A1(n12498), .A2(n10354), .ZN(n12345) );
  NAND2_X1 U10652 ( .A1(n10557), .A2(n12298), .ZN(n8243) );
  NAND2_X1 U10653 ( .A1(n8659), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8250) );
  NAND2_X1 U10654 ( .A1(n8592), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8249) );
  NAND2_X1 U10655 ( .A1(n10564), .A2(n9936), .ZN(n8265) );
  NAND2_X1 U10656 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8244) );
  AND2_X1 U10657 ( .A1(n8265), .A2(n8244), .ZN(n10686) );
  OR2_X1 U10658 ( .A1(n8904), .A2(n10686), .ZN(n8248) );
  INV_X1 U10659 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n8246) );
  OR2_X1 U10660 ( .A1(n8245), .A2(n8246), .ZN(n8247) );
  NAND2_X1 U10661 ( .A1(n8251), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8252) );
  MUX2_X1 U10662 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8252), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8253) );
  AND2_X1 U10663 ( .A1(n8253), .A2(n8274), .ZN(n9941) );
  NAND2_X1 U10664 ( .A1(n9214), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8256) );
  XNOR2_X1 U10665 ( .A(n8277), .B(n8276), .ZN(n9229) );
  OR2_X1 U10666 ( .A1(n12281), .A2(n9229), .ZN(n8260) );
  OR2_X1 U10667 ( .A1(n8258), .A2(SI_4_), .ZN(n8259) );
  OAI211_X1 U10668 ( .C1(n9941), .C2(n9753), .A(n8260), .B(n8259), .ZN(n15012)
         );
  XNOR2_X1 U10669 ( .A(n12353), .B(n15012), .ZN(n10684) );
  INV_X1 U10670 ( .A(n10684), .ZN(n12344) );
  NAND2_X1 U10671 ( .A1(n10685), .A2(n12344), .ZN(n8262) );
  INV_X1 U10672 ( .A(n12353), .ZN(n12350) );
  INV_X1 U10673 ( .A(n15012), .ZN(n8673) );
  NAND2_X1 U10674 ( .A1(n12350), .A2(n8673), .ZN(n8261) );
  NAND2_X1 U10675 ( .A1(n10393), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8272) );
  NAND2_X1 U10676 ( .A1(n8659), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8271) );
  INV_X1 U10677 ( .A(n8265), .ZN(n8264) );
  INV_X1 U10678 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U10679 ( .A1(n8264), .A2(n8263), .ZN(n8283) );
  NAND2_X1 U10680 ( .A1(n8265), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8266) );
  AND2_X1 U10681 ( .A1(n8283), .A2(n8266), .ZN(n10550) );
  OR2_X1 U10682 ( .A1(n8904), .A2(n10550), .ZN(n8270) );
  INV_X1 U10683 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n8268) );
  OR2_X1 U10684 ( .A1(n6448), .A2(n8268), .ZN(n8269) );
  NAND4_X1 U10685 ( .A1(n8272), .A2(n8271), .A3(n8270), .A4(n8269), .ZN(n12497) );
  NAND2_X1 U10686 ( .A1(n8274), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8273) );
  MUX2_X1 U10687 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8273), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8275) );
  NAND2_X1 U10688 ( .A1(n8275), .A2(n8398), .ZN(n14922) );
  NAND2_X1 U10689 ( .A1(n8277), .A2(n8276), .ZN(n8279) );
  NAND2_X1 U10690 ( .A1(n9204), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8278) );
  XNOR2_X1 U10691 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8280) );
  XNOR2_X1 U10692 ( .A(n8292), .B(n8280), .ZN(n9231) );
  OR2_X1 U10693 ( .A1(n12281), .A2(n9231), .ZN(n8282) );
  OR2_X1 U10694 ( .A1(n8258), .A2(SI_5_), .ZN(n8281) );
  OAI211_X1 U10695 ( .C1(n10203), .C2(n9753), .A(n8282), .B(n8281), .ZN(n15017) );
  INV_X1 U10696 ( .A(n15017), .ZN(n10662) );
  NAND2_X1 U10697 ( .A1(n8797), .A2(n10662), .ZN(n12359) );
  NAND2_X1 U10698 ( .A1(n12497), .A2(n15017), .ZN(n12349) );
  NAND2_X1 U10699 ( .A1(n10393), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8288) );
  NAND2_X1 U10700 ( .A1(n8659), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8287) );
  NAND2_X1 U10701 ( .A1(n8283), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8284) );
  AND2_X1 U10702 ( .A1(n8299), .A2(n8284), .ZN(n10904) );
  OR2_X1 U10703 ( .A1(n8904), .A2(n10904), .ZN(n8286) );
  INV_X1 U10704 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10188) );
  OR2_X1 U10705 ( .A1(n6447), .A2(n10188), .ZN(n8285) );
  INV_X1 U10706 ( .A(n12496), .ZN(n10771) );
  NAND2_X1 U10707 ( .A1(n8398), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8290) );
  INV_X1 U10708 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8289) );
  INV_X1 U10709 ( .A(SI_6_), .ZN(n9258) );
  OR2_X1 U10710 ( .A1(n8258), .A2(n9258), .ZN(n8295) );
  NAND2_X1 U10711 ( .A1(n9218), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8293) );
  XNOR2_X1 U10712 ( .A(n8307), .B(n8306), .ZN(n9259) );
  OR2_X1 U10713 ( .A1(n12281), .A2(n9259), .ZN(n8294) );
  OAI211_X1 U10714 ( .C1(n9753), .C2(n10525), .A(n8295), .B(n8294), .ZN(n10674) );
  NAND2_X1 U10715 ( .A1(n10771), .A2(n10674), .ZN(n12361) );
  INV_X1 U10716 ( .A(n10674), .ZN(n15022) );
  NAND2_X1 U10717 ( .A1(n12496), .A2(n15022), .ZN(n12360) );
  NAND2_X1 U10718 ( .A1(n12361), .A2(n12360), .ZN(n10909) );
  NAND2_X1 U10719 ( .A1(n8659), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8305) );
  INV_X1 U10720 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n8296) );
  OR2_X1 U10721 ( .A1(n8245), .A2(n8296), .ZN(n8304) );
  NAND2_X1 U10722 ( .A1(n8299), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8300) );
  AND2_X1 U10723 ( .A1(n8333), .A2(n8300), .ZN(n10815) );
  OR2_X1 U10724 ( .A1(n8904), .A2(n10815), .ZN(n8303) );
  INV_X1 U10725 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n8301) );
  OR2_X1 U10726 ( .A1(n6447), .A2(n8301), .ZN(n8302) );
  OR2_X1 U10727 ( .A1(n8258), .A2(SI_7_), .ZN(n8313) );
  NAND2_X1 U10728 ( .A1(n9237), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8308) );
  XNOR2_X1 U10729 ( .A(n6603), .B(n8325), .ZN(n9233) );
  OR2_X1 U10730 ( .A1(n12281), .A2(n9233), .ZN(n8312) );
  INV_X1 U10731 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n12985) );
  NOR2_X1 U10732 ( .A1(n8319), .A2(n12985), .ZN(n8310) );
  XNOR2_X1 U10733 ( .A(n8310), .B(P3_IR_REG_7__SCAN_IN), .ZN(n10537) );
  OR2_X1 U10734 ( .A1(n9753), .A2(n7145), .ZN(n8311) );
  NAND2_X1 U10735 ( .A1(n10884), .A2(n10812), .ZN(n12366) );
  INV_X1 U10736 ( .A(n10884), .ZN(n12495) );
  NAND2_X1 U10737 ( .A1(n12495), .A2(n15027), .ZN(n12367) );
  NAND2_X1 U10738 ( .A1(n12366), .A2(n12367), .ZN(n10768) );
  INV_X1 U10739 ( .A(n10768), .ZN(n12363) );
  NAND2_X1 U10740 ( .A1(n8659), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8317) );
  NAND2_X1 U10741 ( .A1(n9092), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8316) );
  XNOR2_X1 U10742 ( .A(n8333), .B(n10533), .ZN(n10937) );
  OR2_X1 U10743 ( .A1(n8904), .A2(n10937), .ZN(n8315) );
  INV_X1 U10744 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n10522) );
  OR2_X1 U10745 ( .A1(n6448), .A2(n10522), .ZN(n8314) );
  NAND4_X1 U10746 ( .A1(n8317), .A2(n8316), .A3(n8315), .A4(n8314), .ZN(n12494) );
  INV_X1 U10747 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8318) );
  INV_X1 U10748 ( .A(n8323), .ZN(n8320) );
  NAND2_X1 U10749 ( .A1(n8320), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8321) );
  INV_X1 U10750 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8322) );
  MUX2_X1 U10751 ( .A(n8321), .B(P3_IR_REG_31__SCAN_IN), .S(n8322), .Z(n8324)
         );
  NAND2_X1 U10752 ( .A1(n8323), .A2(n8322), .ZN(n8341) );
  NAND2_X1 U10753 ( .A1(n8324), .A2(n8341), .ZN(n10716) );
  INV_X1 U10754 ( .A(n8325), .ZN(n8326) );
  NAND2_X1 U10755 ( .A1(n9263), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8328) );
  XNOR2_X1 U10756 ( .A(n8346), .B(n8345), .ZN(n9269) );
  OR2_X1 U10757 ( .A1(n12281), .A2(n9269), .ZN(n8330) );
  INV_X1 U10758 ( .A(SI_8_), .ZN(n9270) );
  OR2_X1 U10759 ( .A1(n8258), .A2(n9270), .ZN(n8329) );
  OAI211_X1 U10760 ( .C1(n9753), .C2(n10716), .A(n8330), .B(n8329), .ZN(n10886) );
  XNOR2_X1 U10761 ( .A(n12494), .B(n10886), .ZN(n12369) );
  NAND2_X1 U10762 ( .A1(n10931), .A2(n12369), .ZN(n8331) );
  NAND2_X1 U10763 ( .A1(n11104), .A2(n10886), .ZN(n12372) );
  NAND2_X1 U10764 ( .A1(n8659), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8339) );
  NAND2_X1 U10765 ( .A1(n8592), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8338) );
  OAI21_X1 U10766 ( .B1(n8333), .B2(P3_REG3_REG_8__SCAN_IN), .A(
        P3_REG3_REG_9__SCAN_IN), .ZN(n8334) );
  NAND2_X1 U10767 ( .A1(n10533), .A2(n10723), .ZN(n8332) );
  AND2_X1 U10768 ( .A1(n8334), .A2(n8352), .ZN(n11105) );
  OR2_X1 U10769 ( .A1(n8904), .A2(n11105), .ZN(n8337) );
  INV_X1 U10770 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n8335) );
  OR2_X1 U10771 ( .A1(n8245), .A2(n8335), .ZN(n8336) );
  INV_X1 U10772 ( .A(n12493), .ZN(n11114) );
  NAND2_X1 U10773 ( .A1(n8341), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8340) );
  MUX2_X1 U10774 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8340), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n8344) );
  INV_X1 U10775 ( .A(n8341), .ZN(n8343) );
  INV_X1 U10776 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8342) );
  NAND2_X1 U10777 ( .A1(n8343), .A2(n8342), .ZN(n8371) );
  NAND2_X1 U10778 ( .A1(n8344), .A2(n8371), .ZN(n10727) );
  INV_X1 U10779 ( .A(n10727), .ZN(n10994) );
  OR2_X1 U10780 ( .A1(n8258), .A2(SI_9_), .ZN(n8348) );
  XNOR2_X1 U10781 ( .A(n9292), .B(P1_DATAO_REG_9__SCAN_IN), .ZN(n8359) );
  XNOR2_X1 U10782 ( .A(n8361), .B(n8359), .ZN(n9221) );
  OR2_X1 U10783 ( .A1(n12281), .A2(n9221), .ZN(n8347) );
  OAI211_X1 U10784 ( .C1(n10994), .C2(n9753), .A(n8348), .B(n8347), .ZN(n15038) );
  INV_X1 U10785 ( .A(n15038), .ZN(n11108) );
  NAND2_X1 U10786 ( .A1(n11114), .A2(n11108), .ZN(n12377) );
  INV_X1 U10787 ( .A(n12377), .ZN(n8349) );
  NAND2_X1 U10788 ( .A1(n12493), .A2(n15038), .ZN(n12376) );
  NAND2_X1 U10789 ( .A1(n8659), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8357) );
  NAND2_X1 U10790 ( .A1(n10393), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8356) );
  INV_X1 U10791 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n8350) );
  NAND2_X1 U10792 ( .A1(n8352), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8353) );
  AND2_X1 U10793 ( .A1(n8383), .A2(n8353), .ZN(n11235) );
  OR2_X1 U10794 ( .A1(n8904), .A2(n11235), .ZN(n8355) );
  INV_X1 U10795 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n10997) );
  OR2_X1 U10796 ( .A1(n6447), .A2(n10997), .ZN(n8354) );
  NAND4_X1 U10797 ( .A1(n8357), .A2(n8356), .A3(n8355), .A4(n8354), .ZN(n12492) );
  NAND2_X1 U10798 ( .A1(n8371), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8358) );
  OR2_X1 U10799 ( .A1(n8258), .A2(SI_10_), .ZN(n8365) );
  INV_X1 U10800 ( .A(n8359), .ZN(n8360) );
  NAND2_X1 U10801 ( .A1(n9292), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8362) );
  XNOR2_X1 U10802 ( .A(n8377), .B(P1_DATAO_REG_10__SCAN_IN), .ZN(n8374) );
  XNOR2_X1 U10803 ( .A(n8376), .B(n8374), .ZN(n9225) );
  OR2_X1 U10804 ( .A1(n12281), .A2(n9225), .ZN(n8364) );
  OAI211_X1 U10805 ( .C1(n14967), .C2(n9753), .A(n8365), .B(n8364), .ZN(n15045) );
  NAND2_X1 U10806 ( .A1(n12492), .A2(n15045), .ZN(n12380) );
  INV_X1 U10807 ( .A(n12380), .ZN(n8366) );
  INV_X1 U10808 ( .A(n15045), .ZN(n11232) );
  NAND2_X1 U10809 ( .A1(n11352), .A2(n11232), .ZN(n12381) );
  NAND2_X1 U10810 ( .A1(n8659), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8370) );
  INV_X1 U10811 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11004) );
  OR2_X1 U10812 ( .A1(n8245), .A2(n11004), .ZN(n8369) );
  INV_X1 U10813 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11015) );
  XNOR2_X1 U10814 ( .A(n8383), .B(n11015), .ZN(n11239) );
  OR2_X1 U10815 ( .A1(n8904), .A2(n11239), .ZN(n8368) );
  INV_X1 U10816 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n11003) );
  OR2_X1 U10817 ( .A1(n6448), .A2(n11003), .ZN(n8367) );
  OAI21_X1 U10818 ( .B1(n8371), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8373) );
  INV_X1 U10819 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8372) );
  XNOR2_X1 U10820 ( .A(n8373), .B(n8372), .ZN(n11000) );
  OR2_X1 U10821 ( .A1(n8258), .A2(SI_11_), .ZN(n8382) );
  INV_X1 U10822 ( .A(n8374), .ZN(n8375) );
  NAND2_X1 U10823 ( .A1(n8377), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8378) );
  XNOR2_X1 U10824 ( .A(n9346), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n8380) );
  XNOR2_X1 U10825 ( .A(n8390), .B(n8380), .ZN(n9223) );
  OR2_X1 U10826 ( .A1(n12281), .A2(n9223), .ZN(n8381) );
  OAI211_X1 U10827 ( .C1(n11076), .C2(n9753), .A(n8382), .B(n8381), .ZN(n14481) );
  XNOR2_X1 U10828 ( .A(n12859), .B(n14481), .ZN(n12382) );
  INV_X1 U10829 ( .A(n14481), .ZN(n12388) );
  NAND2_X1 U10830 ( .A1(n12859), .A2(n12388), .ZN(n12387) );
  NAND2_X1 U10831 ( .A1(n8659), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8388) );
  NAND2_X1 U10832 ( .A1(n10393), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8387) );
  OAI21_X1 U10833 ( .B1(n8383), .B2(P3_REG3_REG_11__SCAN_IN), .A(
        P3_REG3_REG_12__SCAN_IN), .ZN(n8384) );
  AND2_X1 U10834 ( .A1(n8384), .A2(n8416), .ZN(n12865) );
  OR2_X1 U10835 ( .A1(n8904), .A2(n12865), .ZN(n8386) );
  INV_X1 U10836 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n11066) );
  OR2_X1 U10837 ( .A1(n6447), .A2(n11066), .ZN(n8385) );
  NAND4_X1 U10838 ( .A1(n8388), .A2(n8387), .A3(n8386), .A4(n8385), .ZN(n12843) );
  NAND2_X1 U10839 ( .A1(n9346), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8391) );
  NAND2_X1 U10840 ( .A1(n9423), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8407) );
  NAND2_X1 U10841 ( .A1(n9419), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8392) );
  NAND2_X1 U10842 ( .A1(n8407), .A2(n8392), .ZN(n8393) );
  NAND2_X1 U10843 ( .A1(n8394), .A2(n8393), .ZN(n8395) );
  NAND2_X1 U10844 ( .A1(n8408), .A2(n8395), .ZN(n9267) );
  NAND2_X1 U10845 ( .A1(n9267), .A2(n12277), .ZN(n8404) );
  INV_X1 U10846 ( .A(n8396), .ZN(n8397) );
  NOR2_X1 U10847 ( .A1(n8398), .A2(n8397), .ZN(n8401) );
  INV_X1 U10848 ( .A(n8401), .ZN(n8399) );
  NAND2_X1 U10849 ( .A1(n8399), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8400) );
  MUX2_X1 U10850 ( .A(n8400), .B(P3_IR_REG_31__SCAN_IN), .S(n6713), .Z(n8402)
         );
  NAND2_X1 U10851 ( .A1(n8401), .A2(n6713), .ZN(n8410) );
  OR2_X1 U10852 ( .A1(n9753), .A2(n12514), .ZN(n8403) );
  INV_X1 U10853 ( .A(n14477), .ZN(n8405) );
  NAND2_X1 U10854 ( .A1(n11335), .A2(n8405), .ZN(n12392) );
  NAND2_X1 U10855 ( .A1(n12843), .A2(n14477), .ZN(n12391) );
  XNOR2_X1 U10856 ( .A(n8422), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9297) );
  NAND2_X1 U10857 ( .A1(n9297), .A2(n12277), .ZN(n8413) );
  NAND2_X1 U10858 ( .A1(n8410), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8411) );
  XNOR2_X1 U10859 ( .A(n8411), .B(P3_IR_REG_13__SCAN_IN), .ZN(n12511) );
  AOI22_X1 U10860 ( .A1(n8516), .A2(SI_13_), .B1(n8515), .B2(n12511), .ZN(
        n8412) );
  NAND2_X1 U10861 ( .A1(n8413), .A2(n8412), .ZN(n12847) );
  INV_X1 U10862 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12849) );
  OR2_X1 U10863 ( .A1(n8245), .A2(n12849), .ZN(n8421) );
  INV_X1 U10864 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n15159) );
  OR2_X1 U10865 ( .A1(n8238), .A2(n15159), .ZN(n8420) );
  INV_X1 U10866 ( .A(n8416), .ZN(n8415) );
  INV_X1 U10867 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8414) );
  NAND2_X1 U10868 ( .A1(n8416), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8417) );
  AND2_X1 U10869 ( .A1(n8431), .A2(n8417), .ZN(n12848) );
  OR2_X1 U10870 ( .A1(n8904), .A2(n12848), .ZN(n8419) );
  INV_X1 U10871 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14983) );
  OR2_X1 U10872 ( .A1(n6447), .A2(n14983), .ZN(n8418) );
  NAND2_X1 U10873 ( .A1(n12847), .A2(n12861), .ZN(n12396) );
  OR2_X1 U10874 ( .A1(n12847), .A2(n12861), .ZN(n12397) );
  NAND2_X1 U10875 ( .A1(n9948), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8440) );
  INV_X1 U10876 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9949) );
  NAND2_X1 U10877 ( .A1(n9949), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8425) );
  XNOR2_X1 U10878 ( .A(n8439), .B(n8438), .ZN(n9303) );
  NAND2_X1 U10879 ( .A1(n9303), .A2(n12277), .ZN(n8429) );
  OR2_X1 U10880 ( .A1(n8426), .A2(n12985), .ZN(n8427) );
  XNOR2_X1 U10881 ( .A(n8427), .B(n8443), .ZN(n12527) );
  AOI22_X1 U10882 ( .A1(n8516), .A2(n9302), .B1(n8515), .B2(n12527), .ZN(n8428) );
  NAND2_X1 U10883 ( .A1(n10393), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8436) );
  NAND2_X1 U10884 ( .A1(n8659), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8435) );
  NAND2_X1 U10885 ( .A1(n8431), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8432) );
  AND2_X1 U10886 ( .A1(n8447), .A2(n8432), .ZN(n12826) );
  OR2_X1 U10887 ( .A1(n8904), .A2(n12826), .ZN(n8434) );
  INV_X1 U10888 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12923) );
  OR2_X1 U10889 ( .A1(n6448), .A2(n12923), .ZN(n8433) );
  NAND2_X1 U10890 ( .A1(n12976), .A2(n12842), .ZN(n12401) );
  NAND2_X1 U10891 ( .A1(n12407), .A2(n12401), .ZN(n12824) );
  INV_X1 U10892 ( .A(n12824), .ZN(n8437) );
  NAND2_X1 U10893 ( .A1(n9844), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8456) );
  NAND2_X1 U10894 ( .A1(n9846), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8442) );
  NAND2_X1 U10895 ( .A1(n8456), .A2(n8442), .ZN(n8453) );
  XNOR2_X1 U10896 ( .A(n8455), .B(n8453), .ZN(n9347) );
  NAND2_X1 U10897 ( .A1(n9347), .A2(n12277), .ZN(n8446) );
  OR2_X1 U10898 ( .A1(n8459), .A2(n12985), .ZN(n8444) );
  XNOR2_X1 U10899 ( .A(n8444), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U10900 ( .A1(n8516), .A2(SI_15_), .B1(n8515), .B2(n12553), .ZN(
        n8445) );
  NAND2_X1 U10901 ( .A1(n8446), .A2(n8445), .ZN(n12811) );
  NAND2_X1 U10902 ( .A1(n10393), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U10903 ( .A1(n8659), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8451) );
  NAND2_X1 U10904 ( .A1(n8447), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8448) );
  AND2_X1 U10905 ( .A1(n8464), .A2(n8448), .ZN(n12812) );
  OR2_X1 U10906 ( .A1(n8904), .A2(n12812), .ZN(n8450) );
  INV_X1 U10907 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14460) );
  OR2_X1 U10908 ( .A1(n6447), .A2(n14460), .ZN(n8449) );
  NAND4_X1 U10909 ( .A1(n8452), .A2(n8451), .A3(n8450), .A4(n8449), .ZN(n12820) );
  OR2_X1 U10910 ( .A1(n12811), .A2(n12160), .ZN(n12400) );
  NAND2_X1 U10911 ( .A1(n12811), .A2(n12160), .ZN(n12405) );
  NAND2_X1 U10912 ( .A1(n12400), .A2(n12405), .ZN(n12803) );
  INV_X1 U10913 ( .A(n12803), .ZN(n12810) );
  INV_X1 U10914 ( .A(n8453), .ZN(n8454) );
  NAND2_X1 U10915 ( .A1(n9995), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8473) );
  NAND2_X1 U10916 ( .A1(n9990), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U10917 ( .A1(n8473), .A2(n8457), .ZN(n8470) );
  XNOR2_X1 U10918 ( .A(n8472), .B(n8470), .ZN(n14398) );
  NAND2_X1 U10919 ( .A1(n14398), .A2(n12277), .ZN(n8462) );
  INV_X1 U10920 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8458) );
  NAND2_X1 U10921 ( .A1(n8459), .A2(n8458), .ZN(n8478) );
  NAND2_X1 U10922 ( .A1(n8478), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8460) );
  XNOR2_X1 U10923 ( .A(n8460), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U10924 ( .A1(n8516), .A2(SI_16_), .B1(n8515), .B2(n12555), .ZN(
        n8461) );
  NAND2_X1 U10925 ( .A1(n9092), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8469) );
  NAND2_X1 U10926 ( .A1(n8659), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8468) );
  INV_X1 U10927 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n12195) );
  NAND2_X1 U10928 ( .A1(n8464), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8465) );
  AND2_X1 U10929 ( .A1(n8482), .A2(n8465), .ZN(n12794) );
  OR2_X1 U10930 ( .A1(n8904), .A2(n12794), .ZN(n8467) );
  INV_X1 U10931 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12554) );
  OR2_X1 U10932 ( .A1(n6448), .A2(n12554), .ZN(n8466) );
  NAND4_X1 U10933 ( .A1(n8469), .A2(n8468), .A3(n8467), .A4(n8466), .ZN(n12805) );
  INV_X1 U10934 ( .A(n12805), .ZN(n12262) );
  OR2_X1 U10935 ( .A1(n12914), .A2(n12262), .ZN(n12409) );
  NAND2_X1 U10936 ( .A1(n12914), .A2(n12262), .ZN(n12406) );
  NAND2_X1 U10937 ( .A1(n12799), .A2(n12798), .ZN(n12797) );
  INV_X1 U10938 ( .A(n8470), .ZN(n8471) );
  NAND2_X1 U10939 ( .A1(n10075), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U10940 ( .A1(n10077), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8474) );
  OR2_X1 U10941 ( .A1(n8476), .A2(n8475), .ZN(n8477) );
  NAND2_X1 U10942 ( .A1(n8489), .A2(n8477), .ZN(n9637) );
  OR2_X1 U10943 ( .A1(n9637), .A2(n12281), .ZN(n8481) );
  NAND2_X1 U10944 ( .A1(n8494), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8479) );
  XNOR2_X1 U10945 ( .A(n8479), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U10946 ( .A1(n8516), .A2(SI_17_), .B1(n8515), .B2(n12591), .ZN(
        n8480) );
  NAND2_X1 U10947 ( .A1(n8659), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8487) );
  INV_X1 U10948 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12784) );
  OR2_X1 U10949 ( .A1(n8245), .A2(n12784), .ZN(n8486) );
  NAND2_X1 U10950 ( .A1(n8482), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8483) );
  AND2_X1 U10951 ( .A1(n8500), .A2(n8483), .ZN(n12783) );
  OR2_X1 U10952 ( .A1(n8904), .A2(n12783), .ZN(n8485) );
  INV_X1 U10953 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12575) );
  OR2_X1 U10954 ( .A1(n6447), .A2(n12575), .ZN(n8484) );
  NAND4_X1 U10955 ( .A1(n8487), .A2(n8486), .A3(n8485), .A4(n8484), .ZN(n12792) );
  INV_X1 U10956 ( .A(n12792), .ZN(n12769) );
  OR2_X1 U10957 ( .A1(n12910), .A2(n12769), .ZN(n12412) );
  NAND2_X1 U10958 ( .A1(n12910), .A2(n12769), .ZN(n12771) );
  NAND2_X1 U10959 ( .A1(n12412), .A2(n12771), .ZN(n8687) );
  NAND2_X1 U10960 ( .A1(n10259), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8507) );
  NAND2_X1 U10961 ( .A1(n15202), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8490) );
  OR2_X1 U10962 ( .A1(n8492), .A2(n8491), .ZN(n8493) );
  NAND2_X1 U10963 ( .A1(n8508), .A2(n8493), .ZN(n9750) );
  OR2_X1 U10964 ( .A1(n9750), .A2(n12281), .ZN(n8497) );
  NAND2_X1 U10965 ( .A1(n8513), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8495) );
  XNOR2_X1 U10966 ( .A(n8495), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12606) );
  AOI22_X1 U10967 ( .A1(n8516), .A2(SI_18_), .B1(n8515), .B2(n12606), .ZN(
        n8496) );
  NAND2_X1 U10968 ( .A1(n8497), .A2(n8496), .ZN(n12249) );
  NAND2_X1 U10969 ( .A1(n8659), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8505) );
  NAND2_X1 U10970 ( .A1(n10393), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8504) );
  INV_X1 U10971 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n8498) );
  NAND2_X1 U10972 ( .A1(n8500), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8501) );
  AND2_X1 U10973 ( .A1(n8519), .A2(n8501), .ZN(n12774) );
  OR2_X1 U10974 ( .A1(n8904), .A2(n12774), .ZN(n8503) );
  INV_X1 U10975 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12908) );
  OR2_X1 U10976 ( .A1(n6448), .A2(n12908), .ZN(n8502) );
  NAND4_X1 U10977 ( .A1(n8505), .A2(n8504), .A3(n8503), .A4(n8502), .ZN(n12781) );
  INV_X1 U10978 ( .A(n12781), .ZN(n12205) );
  OR2_X1 U10979 ( .A1(n12249), .A2(n12205), .ZN(n12415) );
  NAND2_X1 U10980 ( .A1(n12249), .A2(n12205), .ZN(n12418) );
  INV_X1 U10981 ( .A(n12771), .ZN(n12416) );
  NOR2_X1 U10982 ( .A1(n8690), .A2(n12416), .ZN(n8506) );
  INV_X1 U10983 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10467) );
  NAND2_X1 U10984 ( .A1(n10467), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8525) );
  INV_X1 U10985 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10465) );
  NAND2_X1 U10986 ( .A1(n10465), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8509) );
  OR2_X1 U10987 ( .A1(n8511), .A2(n8510), .ZN(n8512) );
  NAND2_X1 U10988 ( .A1(n8526), .A2(n8512), .ZN(n9811) );
  NAND2_X1 U10989 ( .A1(n9811), .A2(n12277), .ZN(n8518) );
  INV_X1 U10990 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8514) );
  AOI22_X1 U10991 ( .A1(n8516), .A2(n15087), .B1(n8515), .B2(n12612), .ZN(
        n8517) );
  NAND2_X1 U10992 ( .A1(n8659), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8524) );
  NAND2_X1 U10993 ( .A1(n8592), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U10994 ( .A1(n8519), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8520) );
  AND2_X1 U10995 ( .A1(n8532), .A2(n8520), .ZN(n12759) );
  OR2_X1 U10996 ( .A1(n8904), .A2(n12759), .ZN(n8522) );
  INV_X1 U10997 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12760) );
  OR2_X1 U10998 ( .A1(n8245), .A2(n12760), .ZN(n8521) );
  NAND4_X1 U10999 ( .A1(n8524), .A2(n8523), .A3(n8522), .A4(n8521), .ZN(n12491) );
  NAND2_X1 U11000 ( .A1(n12962), .A2(n12491), .ZN(n12424) );
  OR2_X1 U11001 ( .A1(n12962), .A2(n12491), .ZN(n12423) );
  NAND2_X1 U11002 ( .A1(n8528), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8529) );
  NAND2_X1 U11003 ( .A1(n8541), .A2(n8529), .ZN(n10034) );
  OR2_X1 U11004 ( .A1(n8258), .A2(n10033), .ZN(n8530) );
  NAND2_X1 U11005 ( .A1(n8532), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U11006 ( .A1(n8550), .A2(n8533), .ZN(n12748) );
  NAND2_X1 U11007 ( .A1(n8207), .A2(n12748), .ZN(n8538) );
  INV_X1 U11008 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n8534) );
  OR2_X1 U11009 ( .A1(n8245), .A2(n8534), .ZN(n8537) );
  INV_X1 U11010 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12956) );
  OR2_X1 U11011 ( .A1(n8238), .A2(n12956), .ZN(n8536) );
  INV_X1 U11012 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12900) );
  OR2_X1 U11013 ( .A1(n6447), .A2(n12900), .ZN(n8535) );
  NAND2_X1 U11014 ( .A1(n12747), .A2(n12733), .ZN(n12321) );
  NAND2_X1 U11015 ( .A1(n12322), .A2(n12321), .ZN(n12743) );
  INV_X1 U11016 ( .A(n12743), .ZN(n8539) );
  INV_X1 U11017 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11528) );
  NAND2_X1 U11018 ( .A1(n11528), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U11019 ( .A1(n11111), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8542) );
  AND2_X1 U11020 ( .A1(n8557), .A2(n8542), .ZN(n8543) );
  OR2_X1 U11021 ( .A1(n8544), .A2(n8543), .ZN(n8545) );
  NAND2_X1 U11022 ( .A1(n8558), .A2(n8545), .ZN(n10162) );
  OR2_X1 U11023 ( .A1(n8258), .A2(n15192), .ZN(n8546) );
  NAND2_X1 U11024 ( .A1(n10393), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8555) );
  INV_X1 U11025 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U11026 ( .A1(n8550), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8551) );
  NAND2_X1 U11027 ( .A1(n8563), .A2(n8551), .ZN(n12737) );
  NAND2_X1 U11028 ( .A1(n8207), .A2(n12737), .ZN(n8554) );
  INV_X1 U11029 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n15207) );
  OR2_X1 U11030 ( .A1(n8238), .A2(n15207), .ZN(n8553) );
  INV_X1 U11031 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12896) );
  OR2_X1 U11032 ( .A1(n6448), .A2(n12896), .ZN(n8552) );
  NAND4_X1 U11033 ( .A1(n8555), .A2(n8554), .A3(n8553), .A4(n8552), .ZN(n12490) );
  NAND2_X1 U11034 ( .A1(n12182), .A2(n12745), .ZN(n12432) );
  NAND2_X1 U11035 ( .A1(n12736), .A2(n12432), .ZN(n8556) );
  XNOR2_X1 U11036 ( .A(n11269), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8570) );
  XNOR2_X1 U11037 ( .A(n8571), .B(n8570), .ZN(n10228) );
  NAND2_X1 U11038 ( .A1(n10228), .A2(n12277), .ZN(n8560) );
  OR2_X1 U11039 ( .A1(n8258), .A2(n15215), .ZN(n8559) );
  INV_X1 U11040 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U11041 ( .A1(n8563), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8564) );
  NAND2_X1 U11042 ( .A1(n8575), .A2(n8564), .ZN(n12723) );
  NAND2_X1 U11043 ( .A1(n12723), .A2(n8207), .ZN(n8568) );
  NAND2_X1 U11044 ( .A1(n9092), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U11045 ( .A1(n8659), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U11046 ( .A1(n8592), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8565) );
  NAND4_X1 U11047 ( .A1(n8568), .A2(n8567), .A3(n8566), .A4(n8565), .ZN(n12702) );
  INV_X1 U11048 ( .A(n12702), .ZN(n12734) );
  NAND2_X1 U11049 ( .A1(n12722), .A2(n12734), .ZN(n12431) );
  NAND2_X1 U11050 ( .A1(n12721), .A2(n12431), .ZN(n8569) );
  OR2_X1 U11051 ( .A1(n12722), .A2(n12734), .ZN(n12430) );
  NAND2_X1 U11052 ( .A1(n8569), .A2(n12430), .ZN(n12708) );
  NAND2_X1 U11053 ( .A1(n11269), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8572) );
  XNOR2_X1 U11054 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8580) );
  XNOR2_X1 U11055 ( .A(n8581), .B(n8580), .ZN(n10468) );
  NAND2_X1 U11056 ( .A1(n10468), .A2(n12277), .ZN(n8574) );
  OR2_X1 U11057 ( .A1(n8258), .A2(n10470), .ZN(n8573) );
  INV_X1 U11058 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12888) );
  NAND2_X1 U11059 ( .A1(n8575), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U11060 ( .A1(n8590), .A2(n8576), .ZN(n12711) );
  NAND2_X1 U11061 ( .A1(n12711), .A2(n8207), .ZN(n8578) );
  AOI22_X1 U11062 ( .A1(n9092), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n8659), .B2(
        P3_REG0_REG_23__SCAN_IN), .ZN(n8577) );
  OAI211_X1 U11063 ( .C1(n6448), .C2(n12888), .A(n8578), .B(n8577), .ZN(n12685) );
  NAND2_X1 U11064 ( .A1(n12706), .A2(n12685), .ZN(n12681) );
  OR2_X1 U11065 ( .A1(n12706), .A2(n12685), .ZN(n8579) );
  NAND2_X1 U11066 ( .A1(n12681), .A2(n8579), .ZN(n12707) );
  NAND2_X1 U11067 ( .A1(n13672), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8582) );
  NAND2_X1 U11068 ( .A1(n8584), .A2(n11270), .ZN(n8585) );
  XNOR2_X1 U11069 ( .A(n8597), .B(n11582), .ZN(n10816) );
  NAND2_X1 U11070 ( .A1(n10816), .A2(n12277), .ZN(n8587) );
  OR2_X1 U11071 ( .A1(n8258), .A2(n7609), .ZN(n8586) );
  INV_X1 U11072 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U11073 ( .A1(n8590), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8591) );
  NAND2_X1 U11074 ( .A1(n8601), .A2(n8591), .ZN(n12694) );
  NAND2_X1 U11075 ( .A1(n12694), .A2(n8207), .ZN(n8595) );
  AOI22_X1 U11076 ( .A1(n8592), .A2(P3_REG1_REG_24__SCAN_IN), .B1(n8659), .B2(
        P3_REG0_REG_24__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U11077 ( .A1(n10393), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8593) );
  NAND2_X1 U11078 ( .A1(n12211), .A2(n12705), .ZN(n12440) );
  INV_X1 U11079 ( .A(n12685), .ZN(n12719) );
  NOR2_X1 U11080 ( .A1(n12706), .A2(n12719), .ZN(n12690) );
  NOR2_X1 U11081 ( .A1(n12689), .A2(n12690), .ZN(n12442) );
  NAND2_X1 U11082 ( .A1(n12709), .A2(n12442), .ZN(n12692) );
  NAND2_X1 U11083 ( .A1(n12692), .A2(n12440), .ZN(n12673) );
  XNOR2_X1 U11084 ( .A(n13667), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8598) );
  XNOR2_X1 U11085 ( .A(n8609), .B(n8598), .ZN(n10942) );
  NAND2_X1 U11086 ( .A1(n10942), .A2(n12277), .ZN(n8600) );
  OR2_X1 U11087 ( .A1(n8258), .A2(n10943), .ZN(n8599) );
  NAND2_X1 U11088 ( .A1(n8601), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8602) );
  NAND2_X1 U11089 ( .A1(n8617), .A2(n8602), .ZN(n12674) );
  NAND2_X1 U11090 ( .A1(n12674), .A2(n8207), .ZN(n8607) );
  INV_X1 U11091 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12880) );
  NAND2_X1 U11092 ( .A1(n10393), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U11093 ( .A1(n8659), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8603) );
  OAI211_X1 U11094 ( .C1(n12880), .C2(n6447), .A(n8604), .B(n8603), .ZN(n8605)
         );
  INV_X1 U11095 ( .A(n8605), .ZN(n8606) );
  OR2_X1 U11096 ( .A1(n8866), .A2(n12653), .ZN(n12446) );
  NAND2_X1 U11097 ( .A1(n8866), .A2(n12653), .ZN(n12445) );
  NAND2_X1 U11098 ( .A1(n12446), .A2(n12445), .ZN(n12665) );
  NAND2_X1 U11099 ( .A1(n12673), .A2(n12672), .ZN(n12671) );
  NAND2_X1 U11100 ( .A1(n13667), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8608) );
  INV_X1 U11101 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14271) );
  NAND2_X1 U11102 ( .A1(n14271), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8610) );
  AOI22_X1 U11103 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n13662), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n14265), .ZN(n8612) );
  XNOR2_X1 U11104 ( .A(n8625), .B(n8612), .ZN(n11321) );
  INV_X1 U11105 ( .A(n8617), .ZN(n8616) );
  INV_X1 U11106 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U11107 ( .A1(n8617), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U11108 ( .A1(n8631), .A2(n8618), .ZN(n12656) );
  NAND2_X1 U11109 ( .A1(n12656), .A2(n8207), .ZN(n8623) );
  INV_X1 U11110 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12876) );
  NAND2_X1 U11111 ( .A1(n9092), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8620) );
  NAND2_X1 U11112 ( .A1(n8659), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8619) );
  OAI211_X1 U11113 ( .C1(n12876), .C2(n6448), .A(n8620), .B(n8619), .ZN(n8621)
         );
  INV_X1 U11114 ( .A(n8621), .ZN(n8622) );
  NAND2_X1 U11115 ( .A1(n9148), .A2(n8887), .ZN(n12449) );
  NOR2_X1 U11116 ( .A1(n13662), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8624) );
  NAND2_X1 U11117 ( .A1(n13662), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8626) );
  AOI22_X1 U11118 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n13660), .B2(n11612), .ZN(n8627) );
  INV_X1 U11119 ( .A(n8627), .ZN(n8628) );
  NAND2_X1 U11120 ( .A1(n12155), .A2(n12277), .ZN(n8630) );
  OR2_X1 U11121 ( .A1(n8258), .A2(n7635), .ZN(n8629) );
  NAND2_X1 U11122 ( .A1(n8631), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8632) );
  NAND2_X1 U11123 ( .A1(n8657), .A2(n8632), .ZN(n12643) );
  NAND2_X1 U11124 ( .A1(n12643), .A2(n8207), .ZN(n8637) );
  INV_X1 U11125 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n8766) );
  NAND2_X1 U11126 ( .A1(n8659), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U11127 ( .A1(n9092), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8633) );
  OAI211_X1 U11128 ( .C1(n8766), .C2(n6447), .A(n8634), .B(n8633), .ZN(n8635)
         );
  INV_X1 U11129 ( .A(n8635), .ZN(n8636) );
  NAND2_X1 U11130 ( .A1(n6710), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8641) );
  MUX2_X1 U11131 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8641), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n8643) );
  NAND2_X1 U11132 ( .A1(n6521), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8644) );
  NAND2_X1 U11133 ( .A1(n12484), .A2(n10032), .ZN(n8645) );
  NAND2_X1 U11134 ( .A1(n8710), .A2(n8645), .ZN(n8648) );
  NAND2_X1 U11135 ( .A1(n8646), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8647) );
  NAND2_X1 U11136 ( .A1(n8648), .A2(n12329), .ZN(n8650) );
  OAI21_X1 U11137 ( .B1(n8757), .B2(n12323), .A(n8651), .ZN(n8649) );
  NAND2_X1 U11138 ( .A1(n8650), .A2(n8649), .ZN(n8871) );
  INV_X1 U11139 ( .A(n12474), .ZN(n8652) );
  NAND3_X1 U11140 ( .A1(n8871), .A2(n8652), .A3(n15044), .ZN(n8654) );
  AND2_X1 U11141 ( .A1(n12484), .A2(n8757), .ZN(n8653) );
  NAND2_X1 U11142 ( .A1(n12612), .A2(n8653), .ZN(n8759) );
  NAND2_X1 U11143 ( .A1(n8654), .A2(n8759), .ZN(n11117) );
  INV_X1 U11144 ( .A(n8657), .ZN(n8656) );
  INV_X1 U11145 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8655) );
  NAND2_X1 U11146 ( .A1(n8656), .A2(n8655), .ZN(n12620) );
  NAND2_X1 U11147 ( .A1(n8657), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U11148 ( .A1(n12620), .A2(n8658), .ZN(n12635) );
  INV_X1 U11149 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n8911) );
  NAND2_X1 U11150 ( .A1(n8659), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8661) );
  NAND2_X1 U11151 ( .A1(n10393), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8660) );
  OAI211_X1 U11152 ( .C1(n6448), .C2(n8911), .A(n8661), .B(n8660), .ZN(n8662)
         );
  INV_X1 U11153 ( .A(n8664), .ZN(n12481) );
  NAND2_X1 U11154 ( .A1(n9773), .A2(n12481), .ZN(n9764) );
  NAND2_X1 U11155 ( .A1(n9753), .A2(n9764), .ZN(n8882) );
  OAI22_X1 U11156 ( .A1(n10227), .A2(n12862), .B1(n8887), .B2(n12860), .ZN(
        n8665) );
  AOI21_X1 U11157 ( .B1(n12648), .B2(n11117), .A(n8665), .ZN(n8709) );
  INV_X1 U11158 ( .A(n14892), .ZN(n8667) );
  NAND2_X1 U11159 ( .A1(n8666), .A2(n8667), .ZN(n10248) );
  NAND2_X1 U11160 ( .A1(n9979), .A2(n10248), .ZN(n10247) );
  NAND2_X1 U11161 ( .A1(n8783), .A2(n10245), .ZN(n8669) );
  NAND2_X1 U11162 ( .A1(n8231), .A2(n8789), .ZN(n8670) );
  NAND2_X1 U11163 ( .A1(n10301), .A2(n8670), .ZN(n10560) );
  INV_X1 U11164 ( .A(n10560), .ZN(n8671) );
  NAND2_X1 U11165 ( .A1(n12498), .A2(n15006), .ZN(n8672) );
  NAND2_X1 U11166 ( .A1(n10687), .A2(n10684), .ZN(n8675) );
  NAND2_X1 U11167 ( .A1(n12353), .A2(n8673), .ZN(n8674) );
  AND2_X1 U11168 ( .A1(n12496), .A2(n10674), .ZN(n8676) );
  NAND2_X1 U11169 ( .A1(n8797), .A2(n15017), .ZN(n10905) );
  OR2_X1 U11170 ( .A1(n10884), .A2(n15027), .ZN(n8677) );
  NAND2_X1 U11171 ( .A1(n12377), .A2(n12376), .ZN(n12301) );
  INV_X1 U11172 ( .A(n10886), .ZN(n15032) );
  NAND2_X1 U11173 ( .A1(n11104), .A2(n15032), .ZN(n10947) );
  AND2_X1 U11174 ( .A1(n12301), .A2(n10947), .ZN(n8678) );
  NAND2_X1 U11175 ( .A1(n12493), .A2(n11108), .ZN(n8679) );
  NAND2_X1 U11176 ( .A1(n12381), .A2(n12380), .ZN(n12304) );
  NAND2_X1 U11177 ( .A1(n12492), .A2(n11232), .ZN(n8680) );
  NAND2_X1 U11178 ( .A1(n12859), .A2(n14481), .ZN(n8681) );
  NAND2_X1 U11179 ( .A1(n12397), .A2(n12396), .ZN(n12839) );
  INV_X1 U11180 ( .A(n12861), .ZN(n12821) );
  INV_X1 U11181 ( .A(n12842), .ZN(n12234) );
  OR2_X1 U11182 ( .A1(n12976), .A2(n12234), .ZN(n8683) );
  NAND2_X1 U11183 ( .A1(n12818), .A2(n8683), .ZN(n12804) );
  NAND2_X1 U11184 ( .A1(n12804), .A2(n12803), .ZN(n12802) );
  NAND2_X1 U11185 ( .A1(n12811), .A2(n12820), .ZN(n8684) );
  OR2_X1 U11186 ( .A1(n12914), .A2(n12805), .ZN(n8685) );
  NAND2_X1 U11187 ( .A1(n12914), .A2(n12805), .ZN(n8686) );
  NAND2_X1 U11188 ( .A1(n12910), .A2(n12792), .ZN(n8688) );
  OR2_X1 U11189 ( .A1(n12249), .A2(n12781), .ZN(n8691) );
  INV_X1 U11190 ( .A(n12491), .ZN(n12770) );
  OR2_X1 U11191 ( .A1(n12962), .A2(n12770), .ZN(n8692) );
  NAND2_X1 U11192 ( .A1(n12753), .A2(n8692), .ZN(n12742) );
  NAND2_X1 U11193 ( .A1(n12742), .A2(n12743), .ZN(n8694) );
  INV_X1 U11194 ( .A(n12733), .ZN(n12755) );
  NAND2_X1 U11195 ( .A1(n12747), .A2(n12755), .ZN(n8693) );
  OR2_X1 U11196 ( .A1(n12182), .A2(n12490), .ZN(n8695) );
  NAND2_X1 U11197 ( .A1(n12728), .A2(n8695), .ZN(n12717) );
  NAND2_X1 U11198 ( .A1(n12722), .A2(n12702), .ZN(n8696) );
  OR2_X1 U11199 ( .A1(n12722), .A2(n12702), .ZN(n8697) );
  INV_X1 U11200 ( .A(n12689), .ZN(n12682) );
  OR2_X1 U11201 ( .A1(n12707), .A2(n12682), .ZN(n12662) );
  OR2_X1 U11202 ( .A1(n12662), .A2(n12672), .ZN(n8698) );
  NAND2_X1 U11203 ( .A1(n12211), .A2(n12667), .ZN(n8699) );
  OR2_X1 U11204 ( .A1(n12682), .A2(n12681), .ZN(n12679) );
  NAND2_X1 U11205 ( .A1(n8866), .A2(n12686), .ZN(n12651) );
  NAND2_X1 U11206 ( .A1(n9148), .A2(n12668), .ZN(n8701) );
  AND2_X1 U11207 ( .A1(n12651), .A2(n8701), .ZN(n8703) );
  NAND2_X1 U11208 ( .A1(n12664), .A2(n8703), .ZN(n8702) );
  OR2_X1 U11209 ( .A1(n9148), .A2(n12668), .ZN(n8704) );
  AND2_X1 U11210 ( .A1(n8702), .A2(n8704), .ZN(n8707) );
  AND2_X1 U11211 ( .A1(n8703), .A2(n7028), .ZN(n8705) );
  AOI21_X1 U11212 ( .B1(n12452), .B2(n8707), .A(n8706), .ZN(n8708) );
  NOR2_X1 U11213 ( .A1(n12329), .A2(n10032), .ZN(n12479) );
  NOR2_X2 U11214 ( .A1(n8743), .A2(n12479), .ZN(n12858) );
  NAND2_X1 U11215 ( .A1(n8710), .A2(n10032), .ZN(n12475) );
  OR2_X1 U11216 ( .A1(n12475), .A2(n12484), .ZN(n15039) );
  INV_X1 U11217 ( .A(n8712), .ZN(n8713) );
  NAND2_X1 U11218 ( .A1(n8713), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8714) );
  MUX2_X1 U11219 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8714), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8716) );
  XNOR2_X1 U11220 ( .A(n10818), .B(P3_B_REG_SCAN_IN), .ZN(n8719) );
  NAND2_X1 U11221 ( .A1(n8715), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8717) );
  MUX2_X1 U11222 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8717), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8718) );
  NAND2_X1 U11223 ( .A1(n8718), .A2(n8720), .ZN(n10945) );
  NAND2_X1 U11224 ( .A1(n8719), .A2(n10945), .ZN(n8724) );
  NAND2_X1 U11225 ( .A1(n8720), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8721) );
  MUX2_X1 U11226 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8721), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n8723) );
  INV_X1 U11227 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n15222) );
  NAND2_X1 U11228 ( .A1(n8736), .A2(n15222), .ZN(n8726) );
  NAND2_X1 U11229 ( .A1(n11322), .A2(n10945), .ZN(n8725) );
  NAND2_X1 U11230 ( .A1(n11322), .A2(n10818), .ZN(n8727) );
  INV_X1 U11231 ( .A(n8778), .ZN(n12982) );
  NOR2_X1 U11232 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .ZN(
        n8731) );
  NOR4_X1 U11233 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_6__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n8730) );
  NOR4_X1 U11234 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_29__SCAN_IN), .ZN(n8729) );
  NOR4_X1 U11235 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_D_REG_25__SCAN_IN), .A3(
        P3_D_REG_20__SCAN_IN), .A4(P3_D_REG_19__SCAN_IN), .ZN(n8728) );
  NAND4_X1 U11236 ( .A1(n8731), .A2(n8730), .A3(n8729), .A4(n8728), .ZN(n8738)
         );
  NOR4_X1 U11237 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n8735) );
  NOR4_X1 U11238 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_21__SCAN_IN), .ZN(n8734) );
  NOR4_X1 U11239 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8733) );
  NOR4_X1 U11240 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n8732) );
  NAND4_X1 U11241 ( .A1(n8735), .A2(n8734), .A3(n8733), .A4(n8732), .ZN(n8737)
         );
  OAI21_X1 U11242 ( .B1(n8738), .B2(n8737), .A(n8736), .ZN(n8753) );
  NAND3_X1 U11243 ( .A1(n10055), .A2(n12982), .A3(n8753), .ZN(n8872) );
  NOR2_X1 U11244 ( .A1(n10945), .A2(n10818), .ZN(n8739) );
  NAND2_X1 U11245 ( .A1(n8642), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8741) );
  INV_X1 U11246 ( .A(n8863), .ZN(n8869) );
  NAND2_X1 U11247 ( .A1(n12329), .A2(n8757), .ZN(n12477) );
  INV_X1 U11248 ( .A(n12477), .ZN(n8742) );
  AND2_X1 U11249 ( .A1(n8743), .A2(n8742), .ZN(n8870) );
  NAND2_X1 U11250 ( .A1(n8869), .A2(n8870), .ZN(n8749) );
  NOR2_X1 U11251 ( .A1(n12474), .A2(n12457), .ZN(n8744) );
  NAND2_X1 U11252 ( .A1(n8868), .A2(n8744), .ZN(n8883) );
  INV_X1 U11253 ( .A(n10055), .ZN(n8745) );
  NAND3_X1 U11254 ( .A1(n8778), .A2(n8745), .A3(n8753), .ZN(n8877) );
  NAND2_X1 U11255 ( .A1(n8868), .A2(n8871), .ZN(n8746) );
  OAI22_X1 U11256 ( .A1(n8872), .A2(n8883), .B1(n8877), .B2(n8746), .ZN(n8747)
         );
  INV_X1 U11257 ( .A(n8747), .ZN(n8748) );
  INV_X1 U11258 ( .A(n12979), .ZN(n8751) );
  NAND2_X1 U11259 ( .A1(n9117), .A2(n8751), .ZN(n8752) );
  XNOR2_X1 U11260 ( .A(n10055), .B(n8778), .ZN(n8755) );
  AND2_X1 U11261 ( .A1(n8868), .A2(n8753), .ZN(n8754) );
  NAND2_X1 U11262 ( .A1(n12612), .A2(n12484), .ZN(n8756) );
  OAI21_X1 U11263 ( .B1(n8757), .B2(n15044), .A(n8756), .ZN(n8758) );
  AOI21_X1 U11264 ( .B1(n8758), .B2(n12474), .A(n12460), .ZN(n8762) );
  NAND2_X1 U11265 ( .A1(n12474), .A2(n12460), .ZN(n10051) );
  NAND2_X1 U11266 ( .A1(n8759), .A2(n12457), .ZN(n10053) );
  NAND2_X1 U11267 ( .A1(n10051), .A2(n10053), .ZN(n8760) );
  NAND2_X1 U11268 ( .A1(n10055), .A2(n8760), .ZN(n8761) );
  OAI21_X1 U11269 ( .B1(n10055), .B2(n8762), .A(n8761), .ZN(n8763) );
  INV_X1 U11270 ( .A(n8763), .ZN(n8764) );
  INV_X1 U11271 ( .A(n12928), .ZN(n8767) );
  NAND2_X1 U11272 ( .A1(n8771), .A2(n14880), .ZN(n8777) );
  INV_X1 U11273 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8772) );
  OR2_X1 U11274 ( .A1(n14880), .A2(n8772), .ZN(n8773) );
  OAI21_X1 U11275 ( .B1(n8774), .B2(n13640), .A(n8773), .ZN(n8775) );
  INV_X1 U11276 ( .A(n8775), .ZN(n8776) );
  NAND2_X1 U11277 ( .A1(n8777), .A2(n8776), .ZN(P2_U3496) );
  INV_X2 U11278 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NAND2_X1 U11279 ( .A1(n12323), .A2(n10032), .ZN(n8779) );
  INV_X4 U11280 ( .A(n12139), .ZN(n9980) );
  XNOR2_X1 U11281 ( .A(n12910), .B(n9980), .ZN(n8825) );
  INV_X1 U11282 ( .A(n8825), .ZN(n8826) );
  XNOR2_X1 U11283 ( .A(n15012), .B(n9980), .ZN(n8794) );
  NOR2_X1 U11284 ( .A1(n8782), .A2(n10042), .ZN(n8786) );
  NOR3_X1 U11285 ( .A1(n8783), .A2(n10245), .A3(n8788), .ZN(n8784) );
  NOR2_X1 U11286 ( .A1(n8786), .A2(n8784), .ZN(n9984) );
  OAI211_X1 U11287 ( .C1(n8785), .C2(n12139), .A(n9984), .B(n10248), .ZN(n9983) );
  INV_X1 U11288 ( .A(n8786), .ZN(n8787) );
  NAND2_X1 U11289 ( .A1(n9983), .A2(n8787), .ZN(n10078) );
  XNOR2_X1 U11290 ( .A(n8789), .B(n8788), .ZN(n8790) );
  XOR2_X1 U11291 ( .A(n12499), .B(n8790), .Z(n10080) );
  XNOR2_X1 U11292 ( .A(n10354), .B(n8788), .ZN(n8793) );
  XNOR2_X1 U11293 ( .A(n8793), .B(n12498), .ZN(n10357) );
  XOR2_X1 U11294 ( .A(n12353), .B(n8794), .Z(n10445) );
  NAND2_X1 U11295 ( .A1(n10444), .A2(n10445), .ZN(n10443) );
  XNOR2_X1 U11296 ( .A(n15017), .B(n9980), .ZN(n8795) );
  XOR2_X1 U11297 ( .A(n12497), .B(n8795), .Z(n10549) );
  INV_X1 U11298 ( .A(n8795), .ZN(n8796) );
  XNOR2_X1 U11299 ( .A(n10674), .B(n9980), .ZN(n8798) );
  XNOR2_X1 U11300 ( .A(n8798), .B(n12496), .ZN(n10668) );
  OR2_X1 U11301 ( .A1(n10771), .A2(n8798), .ZN(n8799) );
  XNOR2_X1 U11302 ( .A(n10768), .B(n12139), .ZN(n10808) );
  OR2_X1 U11303 ( .A1(n10808), .A2(n10884), .ZN(n8800) );
  XNOR2_X1 U11304 ( .A(n9980), .B(n10886), .ZN(n8801) );
  XNOR2_X1 U11305 ( .A(n8801), .B(n12494), .ZN(n10880) );
  INV_X1 U11306 ( .A(n11100), .ZN(n8804) );
  XNOR2_X1 U11307 ( .A(n9980), .B(n15038), .ZN(n8805) );
  XNOR2_X1 U11308 ( .A(n12493), .B(n8805), .ZN(n11101) );
  INV_X1 U11309 ( .A(n11101), .ZN(n8803) );
  INV_X1 U11310 ( .A(n8805), .ZN(n8806) );
  XNOR2_X1 U11311 ( .A(n15045), .B(n9980), .ZN(n8809) );
  XNOR2_X1 U11312 ( .A(n8809), .B(n12492), .ZN(n11226) );
  INV_X1 U11313 ( .A(n11226), .ZN(n8808) );
  INV_X1 U11314 ( .A(n8809), .ZN(n8810) );
  XNOR2_X1 U11315 ( .A(n14481), .B(n9980), .ZN(n8812) );
  NAND2_X1 U11316 ( .A1(n8813), .A2(n8812), .ZN(n11346) );
  NAND2_X1 U11317 ( .A1(n11346), .A2(n12859), .ZN(n8814) );
  XOR2_X1 U11318 ( .A(n9980), .B(n14477), .Z(n11336) );
  INV_X1 U11319 ( .A(n11336), .ZN(n8815) );
  NOR2_X1 U11320 ( .A1(n8815), .A2(n12843), .ZN(n8816) );
  XNOR2_X1 U11321 ( .A(n12847), .B(n9980), .ZN(n8817) );
  NOR2_X1 U11322 ( .A1(n8817), .A2(n12861), .ZN(n12231) );
  XNOR2_X1 U11323 ( .A(n12976), .B(n9980), .ZN(n8818) );
  XOR2_X1 U11324 ( .A(n12842), .B(n8818), .Z(n12158) );
  XNOR2_X1 U11325 ( .A(n12811), .B(n12139), .ZN(n12258) );
  NOR2_X1 U11326 ( .A1(n12258), .A2(n12820), .ZN(n8822) );
  INV_X1 U11327 ( .A(n12258), .ZN(n8821) );
  XNOR2_X1 U11328 ( .A(n12914), .B(n9980), .ZN(n8823) );
  XNOR2_X1 U11329 ( .A(n8823), .B(n12805), .ZN(n12193) );
  INV_X1 U11330 ( .A(n8823), .ZN(n8824) );
  XOR2_X1 U11331 ( .A(n12792), .B(n8825), .Z(n12204) );
  OAI21_X1 U11332 ( .B1(n8826), .B2(n12792), .A(n12202), .ZN(n12251) );
  XNOR2_X1 U11333 ( .A(n12249), .B(n9980), .ZN(n8827) );
  XOR2_X1 U11334 ( .A(n12781), .B(n8827), .Z(n12250) );
  INV_X1 U11335 ( .A(n8827), .ZN(n8828) );
  NAND2_X1 U11336 ( .A1(n8828), .A2(n12781), .ZN(n8829) );
  XNOR2_X1 U11337 ( .A(n12962), .B(n9980), .ZN(n8830) );
  XOR2_X1 U11338 ( .A(n12491), .B(n8830), .Z(n12176) );
  XNOR2_X1 U11339 ( .A(n12747), .B(n9980), .ZN(n8831) );
  NAND2_X1 U11340 ( .A1(n8831), .A2(n12733), .ZN(n12183) );
  OAI21_X1 U11341 ( .B1(n8831), .B2(n12733), .A(n12183), .ZN(n12224) );
  XNOR2_X1 U11342 ( .A(n12182), .B(n9980), .ZN(n8834) );
  XNOR2_X1 U11343 ( .A(n8834), .B(n12490), .ZN(n12184) );
  INV_X1 U11344 ( .A(n12184), .ZN(n8833) );
  OR2_X1 U11345 ( .A1(n12224), .A2(n8833), .ZN(n8832) );
  NOR2_X1 U11346 ( .A1(n12223), .A2(n8832), .ZN(n12186) );
  NAND2_X1 U11347 ( .A1(n8834), .A2(n12745), .ZN(n8836) );
  XNOR2_X1 U11348 ( .A(n12722), .B(n9980), .ZN(n8837) );
  INV_X1 U11349 ( .A(n8841), .ZN(n8839) );
  AND2_X1 U11350 ( .A1(n12184), .A2(n8837), .ZN(n8838) );
  NOR2_X1 U11351 ( .A1(n8839), .A2(n8838), .ZN(n8843) );
  OR2_X1 U11352 ( .A1(n12224), .A2(n8843), .ZN(n8840) );
  AND2_X1 U11353 ( .A1(n12183), .A2(n8841), .ZN(n8842) );
  OR2_X1 U11354 ( .A1(n8843), .A2(n8842), .ZN(n8844) );
  INV_X1 U11355 ( .A(n8850), .ZN(n8848) );
  XNOR2_X1 U11356 ( .A(n12706), .B(n9980), .ZN(n8849) );
  NAND2_X1 U11357 ( .A1(n8848), .A2(n8847), .ZN(n8851) );
  NAND2_X2 U11358 ( .A1(n8850), .A2(n8849), .ZN(n12212) );
  XNOR2_X1 U11359 ( .A(n12211), .B(n9980), .ZN(n8852) );
  INV_X1 U11360 ( .A(n8852), .ZN(n8853) );
  NAND2_X1 U11361 ( .A1(n8853), .A2(n12667), .ZN(n8854) );
  INV_X1 U11362 ( .A(n9139), .ZN(n12217) );
  INV_X1 U11363 ( .A(n9137), .ZN(n8858) );
  XNOR2_X1 U11364 ( .A(n8866), .B(n9980), .ZN(n8855) );
  NAND2_X1 U11365 ( .A1(n8855), .A2(n12653), .ZN(n9132) );
  INV_X1 U11366 ( .A(n8855), .ZN(n8856) );
  NAND2_X1 U11367 ( .A1(n8856), .A2(n12686), .ZN(n8857) );
  NOR3_X1 U11368 ( .A1(n12217), .A2(n8858), .A3(n9115), .ZN(n8865) );
  NAND2_X1 U11369 ( .A1(n9139), .A2(n9137), .ZN(n8859) );
  NAND2_X1 U11370 ( .A1(n8859), .A2(n9115), .ZN(n9136) );
  INV_X1 U11371 ( .A(n9136), .ZN(n8864) );
  NAND2_X1 U11372 ( .A1(n8871), .A2(n15044), .ZN(n8862) );
  NAND2_X1 U11373 ( .A1(n8868), .A2(n8870), .ZN(n8860) );
  OR2_X1 U11374 ( .A1(n8877), .A2(n8860), .ZN(n8861) );
  OAI21_X1 U11375 ( .B1(n8865), .B2(n8864), .A(n12216), .ZN(n8892) );
  INV_X1 U11376 ( .A(n8866), .ZN(n12939) );
  NOR2_X1 U11377 ( .A1(n12475), .A2(n15044), .ZN(n8867) );
  AOI21_X2 U11378 ( .B1(n8869), .B2(n15007), .A(n12828), .ZN(n14891) );
  INV_X1 U11379 ( .A(n8877), .ZN(n8885) );
  INV_X1 U11380 ( .A(n8870), .ZN(n8875) );
  NAND2_X1 U11381 ( .A1(n8872), .A2(n8871), .ZN(n8874) );
  AND3_X1 U11382 ( .A1(n9191), .A2(n9754), .A3(n10051), .ZN(n8873) );
  OAI211_X1 U11383 ( .C1(n8885), .C2(n8875), .A(n8874), .B(n8873), .ZN(n8876)
         );
  NAND2_X1 U11384 ( .A1(n8876), .A2(P3_STATE_REG_SCAN_IN), .ZN(n8879) );
  INV_X1 U11385 ( .A(n8883), .ZN(n12482) );
  NAND2_X1 U11386 ( .A1(n8877), .A2(n12482), .ZN(n8878) );
  INV_X1 U11387 ( .A(n8882), .ZN(n8880) );
  NOR2_X1 U11388 ( .A1(n8883), .A2(n8880), .ZN(n8881) );
  NOR2_X1 U11389 ( .A1(n8883), .A2(n8882), .ZN(n8884) );
  AOI22_X1 U11390 ( .A1(n12667), .A2(n12264), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n8886) );
  OAI21_X1 U11391 ( .B1(n8887), .B2(n12261), .A(n8886), .ZN(n8888) );
  AOI21_X1 U11392 ( .B1(n12674), .B2(n12243), .A(n8888), .ZN(n8889) );
  OAI21_X1 U11393 ( .B1(n12939), .B2(n14891), .A(n8889), .ZN(n8890) );
  NAND2_X1 U11394 ( .A1(n8892), .A2(n8891), .ZN(P3_U3165) );
  NOR2_X1 U11395 ( .A1(n11612), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8894) );
  NAND2_X1 U11396 ( .A1(n11612), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8896) );
  INV_X1 U11397 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14264) );
  AOI22_X1 U11398 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(
        P1_DATAO_REG_28__SCAN_IN), .B1(n13657), .B2(n14264), .ZN(n8897) );
  XNOR2_X1 U11399 ( .A(n9080), .B(n8897), .ZN(n12993) );
  NAND2_X1 U11400 ( .A1(n12993), .A2(n12277), .ZN(n8899) );
  INV_X1 U11401 ( .A(SI_28_), .ZN(n12994) );
  OR2_X1 U11402 ( .A1(n8258), .A2(n12994), .ZN(n8898) );
  NAND2_X1 U11403 ( .A1(n12150), .A2(n10227), .ZN(n9078) );
  OR2_X1 U11404 ( .A1(n9117), .A2(n12489), .ZN(n8901) );
  NAND2_X1 U11405 ( .A1(n8902), .A2(n12461), .ZN(n8903) );
  OR2_X1 U11406 ( .A1(n12620), .A2(n8904), .ZN(n10399) );
  INV_X1 U11407 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9107) );
  NAND2_X1 U11408 ( .A1(n10393), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8906) );
  INV_X1 U11409 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9104) );
  OR2_X1 U11410 ( .A1(n8238), .A2(n9104), .ZN(n8905) );
  OAI211_X1 U11411 ( .C1(n6447), .C2(n9107), .A(n8906), .B(n8905), .ZN(n8907)
         );
  INV_X1 U11412 ( .A(n8907), .ZN(n8908) );
  NAND2_X1 U11413 ( .A1(n10399), .A2(n8908), .ZN(n12488) );
  AOI22_X1 U11414 ( .A1(n12488), .A2(n12841), .B1(n12844), .B2(n12489), .ZN(
        n8909) );
  AOI21_X1 U11415 ( .B1(n12639), .B2(n15049), .A(n8910), .ZN(n8913) );
  INV_X1 U11416 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n8912) );
  MUX2_X1 U11417 ( .A(n8913), .B(n8912), .S(n15050), .Z(n8914) );
  NAND2_X1 U11418 ( .A1(n8914), .A2(n7439), .ZN(P3_U3455) );
  NAND2_X1 U11419 ( .A1(n10266), .A2(n13262), .ZN(n9964) );
  OR2_X1 U11420 ( .A1(n8928), .A2(n14860), .ZN(n8916) );
  INV_X1 U11421 ( .A(n10131), .ZN(n8919) );
  NAND2_X1 U11422 ( .A1(n8917), .A2(n13262), .ZN(n8920) );
  INV_X1 U11423 ( .A(n10132), .ZN(n8918) );
  NAND2_X1 U11424 ( .A1(n8921), .A2(n8920), .ZN(n8922) );
  NAND2_X1 U11425 ( .A1(n10129), .A2(n8922), .ZN(n10096) );
  NAND2_X1 U11426 ( .A1(n13146), .A2(n13262), .ZN(n8925) );
  XNOR2_X1 U11427 ( .A(n8928), .B(n11890), .ZN(n8923) );
  XNOR2_X1 U11428 ( .A(n8925), .B(n8923), .ZN(n10097) );
  INV_X1 U11429 ( .A(n8923), .ZN(n8924) );
  NAND2_X1 U11430 ( .A1(n8925), .A2(n8924), .ZN(n8926) );
  AND2_X1 U11431 ( .A1(n13145), .A2(n13262), .ZN(n8930) );
  XNOR2_X1 U11432 ( .A(n15068), .B(n8928), .ZN(n8929) );
  NAND2_X1 U11433 ( .A1(n8930), .A2(n8929), .ZN(n8934) );
  INV_X1 U11434 ( .A(n8929), .ZN(n8932) );
  INV_X1 U11435 ( .A(n8930), .ZN(n8931) );
  NAND2_X1 U11436 ( .A1(n8932), .A2(n8931), .ZN(n8933) );
  AND2_X1 U11437 ( .A1(n8934), .A2(n8933), .ZN(n10038) );
  INV_X1 U11438 ( .A(n10066), .ZN(n8936) );
  NAND2_X1 U11439 ( .A1(n13144), .A2(n13262), .ZN(n8937) );
  NAND2_X1 U11440 ( .A1(n8938), .A2(n8937), .ZN(n8939) );
  NAND2_X1 U11441 ( .A1(n10064), .A2(n8939), .ZN(n10087) );
  XNOR2_X1 U11442 ( .A(n11908), .B(n8928), .ZN(n8940) );
  NAND2_X1 U11443 ( .A1(n13143), .A2(n13262), .ZN(n8941) );
  XNOR2_X1 U11444 ( .A(n8940), .B(n8941), .ZN(n10088) );
  NAND2_X1 U11445 ( .A1(n10087), .A2(n10088), .ZN(n10086) );
  INV_X1 U11446 ( .A(n8940), .ZN(n8942) );
  NAND2_X1 U11447 ( .A1(n8942), .A2(n8941), .ZN(n8943) );
  XNOR2_X1 U11448 ( .A(n13104), .B(n8928), .ZN(n8944) );
  AND2_X1 U11449 ( .A1(n13142), .A2(n13465), .ZN(n8945) );
  NAND2_X1 U11450 ( .A1(n8944), .A2(n8945), .ZN(n8949) );
  INV_X1 U11451 ( .A(n8944), .ZN(n8947) );
  INV_X1 U11452 ( .A(n8945), .ZN(n8946) );
  NAND2_X1 U11453 ( .A1(n8947), .A2(n8946), .ZN(n8948) );
  AND2_X1 U11454 ( .A1(n8949), .A2(n8948), .ZN(n13100) );
  XNOR2_X1 U11455 ( .A(n11918), .B(n8928), .ZN(n8952) );
  NAND2_X1 U11456 ( .A1(n13141), .A2(n13262), .ZN(n8950) );
  XNOR2_X1 U11457 ( .A(n8952), .B(n8950), .ZN(n10218) );
  INV_X1 U11458 ( .A(n8950), .ZN(n8951) );
  NAND2_X1 U11459 ( .A1(n8952), .A2(n8951), .ZN(n8953) );
  NAND2_X1 U11460 ( .A1(n10217), .A2(n8953), .ZN(n10384) );
  XNOR2_X1 U11461 ( .A(n11923), .B(n9052), .ZN(n8954) );
  NAND2_X1 U11462 ( .A1(n13140), .A2(n13262), .ZN(n8955) );
  NAND2_X1 U11463 ( .A1(n8954), .A2(n8955), .ZN(n10383) );
  INV_X1 U11464 ( .A(n8954), .ZN(n8957) );
  INV_X1 U11465 ( .A(n8955), .ZN(n8956) );
  NAND2_X1 U11466 ( .A1(n8957), .A2(n8956), .ZN(n10382) );
  XNOR2_X1 U11467 ( .A(n13492), .B(n9052), .ZN(n8959) );
  NAND2_X1 U11468 ( .A1(n13139), .A2(n13262), .ZN(n8960) );
  NAND2_X1 U11469 ( .A1(n8959), .A2(n8960), .ZN(n8965) );
  INV_X1 U11470 ( .A(n8959), .ZN(n8962) );
  INV_X1 U11471 ( .A(n8960), .ZN(n8961) );
  NAND2_X1 U11472 ( .A1(n8962), .A2(n8961), .ZN(n8963) );
  NAND2_X1 U11473 ( .A1(n8965), .A2(n8963), .ZN(n10618) );
  INV_X1 U11474 ( .A(n10618), .ZN(n8964) );
  XNOR2_X1 U11475 ( .A(n13479), .B(n9052), .ZN(n8966) );
  NAND2_X1 U11476 ( .A1(n13138), .A2(n13262), .ZN(n8967) );
  XNOR2_X1 U11477 ( .A(n8966), .B(n8967), .ZN(n10677) );
  INV_X1 U11478 ( .A(n8966), .ZN(n8969) );
  INV_X1 U11479 ( .A(n8967), .ZN(n8968) );
  NAND2_X1 U11480 ( .A1(n8969), .A2(n8968), .ZN(n8970) );
  XNOR2_X1 U11481 ( .A(n13600), .B(n8928), .ZN(n8973) );
  NAND2_X1 U11482 ( .A1(n13137), .A2(n13262), .ZN(n8971) );
  XNOR2_X1 U11483 ( .A(n8973), .B(n8971), .ZN(n10820) );
  NAND2_X1 U11484 ( .A1(n10819), .A2(n10820), .ZN(n10958) );
  XNOR2_X1 U11485 ( .A(n11944), .B(n8928), .ZN(n8975) );
  AND2_X1 U11486 ( .A1(n13136), .A2(n13262), .ZN(n8976) );
  NAND2_X1 U11487 ( .A1(n8975), .A2(n8976), .ZN(n10960) );
  INV_X1 U11488 ( .A(n8971), .ZN(n8972) );
  NAND2_X1 U11489 ( .A1(n8973), .A2(n8972), .ZN(n10959) );
  AND2_X1 U11490 ( .A1(n10960), .A2(n10959), .ZN(n8974) );
  NAND2_X1 U11491 ( .A1(n10958), .A2(n8974), .ZN(n8983) );
  XNOR2_X1 U11492 ( .A(n13645), .B(n8928), .ZN(n8981) );
  NAND2_X1 U11493 ( .A1(n13135), .A2(n13262), .ZN(n8979) );
  XNOR2_X1 U11494 ( .A(n8981), .B(n8979), .ZN(n11125) );
  INV_X1 U11495 ( .A(n8975), .ZN(n8978) );
  INV_X1 U11496 ( .A(n8976), .ZN(n8977) );
  NAND2_X1 U11497 ( .A1(n8978), .A2(n8977), .ZN(n11123) );
  AND2_X1 U11498 ( .A1(n11125), .A2(n11123), .ZN(n8982) );
  INV_X1 U11499 ( .A(n8979), .ZN(n8980) );
  XNOR2_X1 U11500 ( .A(n13589), .B(n9052), .ZN(n8984) );
  NAND2_X1 U11501 ( .A1(n13134), .A2(n13262), .ZN(n8985) );
  NAND2_X1 U11502 ( .A1(n8984), .A2(n8985), .ZN(n8989) );
  INV_X1 U11503 ( .A(n8984), .ZN(n8987) );
  INV_X1 U11504 ( .A(n8985), .ZN(n8986) );
  NAND2_X1 U11505 ( .A1(n8987), .A2(n8986), .ZN(n8988) );
  AND2_X1 U11506 ( .A1(n8989), .A2(n8988), .ZN(n11090) );
  XNOR2_X1 U11507 ( .A(n13580), .B(n8928), .ZN(n8990) );
  AND2_X1 U11508 ( .A1(n13425), .A2(n13262), .ZN(n11245) );
  INV_X1 U11509 ( .A(n13037), .ZN(n8997) );
  XNOR2_X1 U11510 ( .A(n13577), .B(n9052), .ZN(n8991) );
  NAND2_X1 U11511 ( .A1(n13133), .A2(n13262), .ZN(n8992) );
  NAND2_X1 U11512 ( .A1(n8991), .A2(n8992), .ZN(n8998) );
  INV_X1 U11513 ( .A(n8991), .ZN(n8994) );
  INV_X1 U11514 ( .A(n8992), .ZN(n8993) );
  NAND2_X1 U11515 ( .A1(n8994), .A2(n8993), .ZN(n8995) );
  NAND2_X1 U11516 ( .A1(n8998), .A2(n8995), .ZN(n13040) );
  NAND2_X1 U11517 ( .A1(n13038), .A2(n8998), .ZN(n13047) );
  XNOR2_X1 U11518 ( .A(n13634), .B(n9052), .ZN(n8999) );
  NAND2_X1 U11519 ( .A1(n13428), .A2(n13262), .ZN(n9000) );
  NAND2_X1 U11520 ( .A1(n8999), .A2(n9000), .ZN(n9004) );
  INV_X1 U11521 ( .A(n8999), .ZN(n9002) );
  INV_X1 U11522 ( .A(n9000), .ZN(n9001) );
  NAND2_X1 U11523 ( .A1(n9002), .A2(n9001), .ZN(n9003) );
  AND2_X1 U11524 ( .A1(n9004), .A2(n9003), .ZN(n13048) );
  XNOR2_X1 U11525 ( .A(n13562), .B(n9052), .ZN(n9005) );
  NAND2_X1 U11526 ( .A1(n13132), .A2(n13262), .ZN(n9006) );
  XNOR2_X1 U11527 ( .A(n9005), .B(n9006), .ZN(n13087) );
  INV_X1 U11528 ( .A(n9005), .ZN(n9008) );
  INV_X1 U11529 ( .A(n9006), .ZN(n9007) );
  NAND2_X1 U11530 ( .A1(n9008), .A2(n9007), .ZN(n9009) );
  XNOR2_X1 U11531 ( .A(n13559), .B(n9052), .ZN(n9010) );
  NAND2_X1 U11532 ( .A1(n13386), .A2(n13465), .ZN(n9011) );
  NAND2_X1 U11533 ( .A1(n9010), .A2(n9011), .ZN(n9015) );
  INV_X1 U11534 ( .A(n9010), .ZN(n9013) );
  INV_X1 U11535 ( .A(n9011), .ZN(n9012) );
  NAND2_X1 U11536 ( .A1(n9013), .A2(n9012), .ZN(n9014) );
  NAND2_X1 U11537 ( .A1(n9015), .A2(n9014), .ZN(n13017) );
  XNOR2_X1 U11538 ( .A(n13553), .B(n9052), .ZN(n9016) );
  NAND2_X1 U11539 ( .A1(n13131), .A2(n13262), .ZN(n9017) );
  NAND2_X1 U11540 ( .A1(n9016), .A2(n9017), .ZN(n9021) );
  INV_X1 U11541 ( .A(n9016), .ZN(n9019) );
  INV_X1 U11542 ( .A(n9017), .ZN(n9018) );
  NAND2_X1 U11543 ( .A1(n9019), .A2(n9018), .ZN(n9020) );
  AND2_X1 U11544 ( .A1(n9021), .A2(n9020), .ZN(n13069) );
  XNOR2_X1 U11545 ( .A(n13549), .B(n9052), .ZN(n9022) );
  NAND2_X1 U11546 ( .A1(n13353), .A2(n13465), .ZN(n9023) );
  XNOR2_X1 U11547 ( .A(n9022), .B(n9023), .ZN(n13022) );
  INV_X1 U11548 ( .A(n9022), .ZN(n9025) );
  INV_X1 U11549 ( .A(n9023), .ZN(n9024) );
  NAND2_X1 U11550 ( .A1(n9025), .A2(n9024), .ZN(n9026) );
  XNOR2_X1 U11551 ( .A(n13626), .B(n9052), .ZN(n9027) );
  AND2_X1 U11552 ( .A1(n13130), .A2(n13262), .ZN(n13079) );
  NAND2_X1 U11553 ( .A1(n9028), .A2(n7311), .ZN(n9029) );
  XNOR2_X1 U11554 ( .A(n13313), .B(n9052), .ZN(n9032) );
  XNOR2_X1 U11555 ( .A(n9031), .B(n9032), .ZN(n13008) );
  NAND2_X1 U11556 ( .A1(n13129), .A2(n13262), .ZN(n13007) );
  XNOR2_X1 U11557 ( .A(n13529), .B(n9052), .ZN(n9034) );
  NAND2_X1 U11558 ( .A1(n13128), .A2(n13262), .ZN(n9035) );
  XNOR2_X1 U11559 ( .A(n9034), .B(n9035), .ZN(n13063) );
  INV_X1 U11560 ( .A(n9034), .ZN(n9037) );
  INV_X1 U11561 ( .A(n9035), .ZN(n9036) );
  NAND2_X1 U11562 ( .A1(n9037), .A2(n9036), .ZN(n9038) );
  NAND2_X1 U11563 ( .A1(n13060), .A2(n9038), .ZN(n13030) );
  XNOR2_X1 U11564 ( .A(n13525), .B(n8928), .ZN(n9041) );
  NAND2_X1 U11565 ( .A1(n13127), .A2(n13262), .ZN(n9039) );
  XNOR2_X1 U11566 ( .A(n9041), .B(n9039), .ZN(n13029) );
  INV_X1 U11567 ( .A(n9039), .ZN(n9040) );
  NAND2_X1 U11568 ( .A1(n9041), .A2(n9040), .ZN(n9042) );
  XNOR2_X1 U11569 ( .A(n13520), .B(n9052), .ZN(n9043) );
  NAND2_X1 U11570 ( .A1(n13245), .A2(n13262), .ZN(n9044) );
  NAND2_X1 U11571 ( .A1(n9043), .A2(n9044), .ZN(n9049) );
  INV_X1 U11572 ( .A(n9043), .ZN(n9046) );
  INV_X1 U11573 ( .A(n9044), .ZN(n9045) );
  NAND2_X1 U11574 ( .A1(n9046), .A2(n9045), .ZN(n9047) );
  NAND2_X1 U11575 ( .A1(n9049), .A2(n9047), .ZN(n13112) );
  XNOR2_X1 U11576 ( .A(n13514), .B(n9052), .ZN(n9051) );
  NAND2_X1 U11577 ( .A1(n13126), .A2(n13262), .ZN(n9050) );
  XNOR2_X1 U11578 ( .A(n9051), .B(n9050), .ZN(n12998) );
  NAND2_X1 U11579 ( .A1(n13244), .A2(n13262), .ZN(n9053) );
  XNOR2_X1 U11580 ( .A(n9053), .B(n9052), .ZN(n9054) );
  INV_X1 U11581 ( .A(n14853), .ZN(n9055) );
  NAND2_X1 U11582 ( .A1(n9056), .A2(n9055), .ZN(n10261) );
  NOR2_X1 U11583 ( .A1(n9069), .A2(n14851), .ZN(n9059) );
  AND2_X1 U11584 ( .A1(n14864), .A2(n9057), .ZN(n9058) );
  AND2_X1 U11585 ( .A1(n14859), .A2(n12097), .ZN(n15069) );
  NAND2_X1 U11586 ( .A1(n9059), .A2(n15069), .ZN(n9061) );
  NAND2_X2 U11587 ( .A1(n14854), .A2(n9060), .ZN(n13487) );
  INV_X1 U11588 ( .A(n9062), .ZN(n9064) );
  NAND2_X1 U11589 ( .A1(n9064), .A2(n9063), .ZN(n9075) );
  INV_X1 U11590 ( .A(n12064), .ZN(n12132) );
  NAND2_X1 U11591 ( .A1(n14854), .A2(n12132), .ZN(n9065) );
  NAND2_X1 U11592 ( .A1(n13125), .A2(n13427), .ZN(n9067) );
  NAND2_X1 U11593 ( .A1(n13126), .A2(n13426), .ZN(n9066) );
  NAND2_X1 U11594 ( .A1(n9067), .A2(n9066), .ZN(n13235) );
  AOI22_X1 U11595 ( .A1(n13116), .A2(n13235), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9073) );
  NAND2_X1 U11596 ( .A1(n9069), .A2(n9068), .ZN(n9071) );
  NAND2_X1 U11597 ( .A1(n9071), .A2(n9070), .ZN(n9961) );
  OR2_X1 U11598 ( .A1(n13239), .A2(n13118), .ZN(n9072) );
  OAI211_X1 U11599 ( .C1(n9076), .C2(n13613), .A(n9075), .B(n9074), .ZN(
        P2_U3192) );
  NAND2_X1 U11600 ( .A1(n9078), .A2(n9077), .ZN(n12458) );
  NOR2_X1 U11601 ( .A1(n13657), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9079) );
  XNOR2_X1 U11602 ( .A(n14260), .B(P1_DATAO_REG_29__SCAN_IN), .ZN(n9081) );
  NAND2_X1 U11603 ( .A1(n9082), .A2(n9081), .ZN(n9083) );
  NAND2_X1 U11604 ( .A1(n12990), .A2(n12277), .ZN(n9085) );
  INV_X1 U11605 ( .A(SI_29_), .ZN(n12992) );
  OR2_X1 U11606 ( .A1(n8258), .A2(n12992), .ZN(n9084) );
  NAND2_X1 U11607 ( .A1(n12631), .A2(n12488), .ZN(n12468) );
  INV_X1 U11608 ( .A(n12631), .ZN(n9086) );
  INV_X1 U11609 ( .A(n12488), .ZN(n12145) );
  NAND2_X1 U11610 ( .A1(n9086), .A2(n12145), .ZN(n12464) );
  NAND2_X1 U11611 ( .A1(n12468), .A2(n12464), .ZN(n12317) );
  OR2_X1 U11612 ( .A1(n10227), .A2(n12637), .ZN(n9087) );
  XNOR2_X1 U11613 ( .A(n9090), .B(n9089), .ZN(n9091) );
  NAND2_X1 U11614 ( .A1(n9091), .A2(n12837), .ZN(n9103) );
  INV_X1 U11615 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n9095) );
  NAND2_X1 U11616 ( .A1(n9092), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9094) );
  INV_X1 U11617 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14485) );
  OR2_X1 U11618 ( .A1(n8238), .A2(n14485), .ZN(n9093) );
  OAI211_X1 U11619 ( .C1(n9095), .C2(n6447), .A(n9094), .B(n9093), .ZN(n9096)
         );
  INV_X1 U11620 ( .A(n9096), .ZN(n9097) );
  INV_X1 U11621 ( .A(P3_B_REG_SCAN_IN), .ZN(n9098) );
  NOR2_X1 U11622 ( .A1(n8664), .A2(n9098), .ZN(n9099) );
  OR2_X1 U11623 ( .A1(n12862), .A2(n9099), .ZN(n12622) );
  NOR2_X1 U11624 ( .A1(n12289), .A2(n12622), .ZN(n9101) );
  XNOR2_X1 U11625 ( .A(n9148), .B(n12139), .ZN(n9109) );
  NOR2_X1 U11626 ( .A1(n9109), .A2(n12668), .ZN(n9111) );
  AOI21_X1 U11627 ( .B1(n9109), .B2(n12668), .A(n9111), .ZN(n9134) );
  INV_X1 U11628 ( .A(n9134), .ZN(n9110) );
  INV_X1 U11629 ( .A(n9111), .ZN(n9112) );
  AND2_X1 U11630 ( .A1(n9137), .A2(n9114), .ZN(n9113) );
  INV_X1 U11631 ( .A(n9114), .ZN(n9116) );
  AND2_X1 U11632 ( .A1(n9115), .A2(n9134), .ZN(n9141) );
  NAND2_X1 U11633 ( .A1(n9123), .A2(n9121), .ZN(n9119) );
  XNOR2_X1 U11634 ( .A(n9117), .B(n12139), .ZN(n12146) );
  NOR2_X1 U11635 ( .A1(n12146), .A2(n12489), .ZN(n12141) );
  AOI21_X1 U11636 ( .B1(n12146), .B2(n12489), .A(n12141), .ZN(n9120) );
  NAND2_X1 U11637 ( .A1(n9119), .A2(n9118), .ZN(n9124) );
  AND2_X1 U11638 ( .A1(n9121), .A2(n9120), .ZN(n9122) );
  NAND2_X1 U11639 ( .A1(n9123), .A2(n9122), .ZN(n12153) );
  NAND2_X1 U11640 ( .A1(n9124), .A2(n12153), .ZN(n9125) );
  NAND2_X1 U11641 ( .A1(n9125), .A2(n12216), .ZN(n9131) );
  AOI22_X1 U11642 ( .A1(n12668), .A2(n12264), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9126) );
  OAI21_X1 U11643 ( .B1(n10227), .B2(n12261), .A(n9126), .ZN(n9127) );
  AOI21_X1 U11644 ( .B1(n12643), .B2(n12243), .A(n9127), .ZN(n9128) );
  OAI21_X1 U11645 ( .B1(n12645), .B2(n14891), .A(n9128), .ZN(n9129) );
  INV_X1 U11646 ( .A(n9129), .ZN(n9130) );
  NAND2_X1 U11647 ( .A1(n9131), .A2(n9130), .ZN(P3_U3154) );
  INV_X1 U11648 ( .A(n9132), .ZN(n9133) );
  NOR2_X1 U11649 ( .A1(n9134), .A2(n9133), .ZN(n9135) );
  NAND2_X1 U11650 ( .A1(n9136), .A2(n9135), .ZN(n9146) );
  AND2_X1 U11651 ( .A1(n9137), .A2(n9140), .ZN(n9138) );
  NAND2_X1 U11652 ( .A1(n9139), .A2(n9138), .ZN(n9144) );
  INV_X1 U11653 ( .A(n9140), .ZN(n9142) );
  OR2_X1 U11654 ( .A1(n9142), .A2(n9141), .ZN(n9143) );
  NAND2_X1 U11655 ( .A1(n9144), .A2(n9143), .ZN(n9145) );
  NAND2_X1 U11656 ( .A1(n9146), .A2(n9145), .ZN(n9147) );
  NAND2_X1 U11657 ( .A1(n9147), .A2(n12216), .ZN(n9154) );
  AOI22_X1 U11658 ( .A1(n12686), .A2(n12264), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9149) );
  OAI21_X1 U11659 ( .B1(n7026), .B2(n12261), .A(n9149), .ZN(n9150) );
  AOI21_X1 U11660 ( .B1(n12656), .B2(n12243), .A(n9150), .ZN(n9151) );
  OAI21_X1 U11661 ( .B1(n12935), .B2(n14891), .A(n9151), .ZN(n9152) );
  INV_X1 U11662 ( .A(n9152), .ZN(n9153) );
  NAND2_X1 U11663 ( .A1(n9154), .A2(n9153), .ZN(P3_U3180) );
  INV_X1 U11664 ( .A(n9155), .ZN(n9156) );
  NOR2_X1 U11665 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n9158) );
  NOR2_X2 U11666 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), 
        .ZN(n9157) );
  INV_X1 U11667 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9243) );
  INV_X1 U11668 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9168) );
  NAND2_X1 U11669 ( .A1(n9243), .A2(n9168), .ZN(n9169) );
  OAI21_X1 U11670 ( .B1(n7293), .B2(n9169), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9171) );
  INV_X1 U11671 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9170) );
  XNOR2_X1 U11672 ( .A(n9171), .B(n9170), .ZN(n9254) );
  NOR2_X1 U11673 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n9174) );
  NOR2_X1 U11674 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n9173) );
  INV_X1 U11675 ( .A(n9185), .ZN(n9175) );
  NAND2_X1 U11676 ( .A1(n9172), .A2(n9175), .ZN(n9178) );
  NAND2_X1 U11677 ( .A1(n9178), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9179) );
  NAND3_X1 U11678 ( .A1(n9183), .A2(n9182), .A3(n9166), .ZN(n9184) );
  NAND2_X1 U11679 ( .A1(n9248), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9188) );
  XNOR2_X1 U11680 ( .A(n9188), .B(n9187), .ZN(n14267) );
  NOR2_X1 U11681 ( .A1(n9273), .A2(n14267), .ZN(n9189) );
  OR2_X2 U11682 ( .A1(n9592), .A2(n9685), .ZN(n13817) );
  INV_X2 U11683 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U11684 ( .A(n12981), .ZN(n9190) );
  NAND2_X1 U11685 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_STATE_REG_SCAN_IN), .ZN(
        n9192) );
  OAI21_X1 U11686 ( .B1(n9193), .B2(P3_STATE_REG_SCAN_IN), .A(n9192), .ZN(
        P3_U3295) );
  NAND2_X1 U11687 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9194) );
  MUX2_X1 U11688 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9194), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9196) );
  INV_X1 U11689 ( .A(n9197), .ZN(n9195) );
  NAND2_X1 U11690 ( .A1(n9196), .A2(n9195), .ZN(n9683) );
  AND2_X1 U11691 ( .A1(n11542), .A2(P1_U3086), .ZN(n9295) );
  INV_X2 U11692 ( .A(n9295), .ZN(n14276) );
  INV_X1 U11693 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9678) );
  NOR2_X1 U11694 ( .A1(n11542), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14272) );
  OAI222_X1 U11695 ( .A1(P1_U3086), .A2(n9683), .B1(n14276), .B2(n9678), .C1(
        n14270), .C2(n9680), .ZN(P1_U3354) );
  INV_X1 U11696 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9235) );
  NOR2_X1 U11697 ( .A1(n9197), .A2(n9235), .ZN(n9198) );
  MUX2_X1 U11698 ( .A(n9235), .B(n9198), .S(P1_IR_REG_2__SCAN_IN), .Z(n9199)
         );
  INV_X1 U11699 ( .A(n9199), .ZN(n9200) );
  NAND2_X1 U11700 ( .A1(n9200), .A2(n9202), .ZN(n9726) );
  OAI222_X1 U11701 ( .A1(n14276), .A2(n9725), .B1(n14270), .B2(n9724), .C1(
        P1_U3086), .C2(n9726), .ZN(P1_U3353) );
  NAND2_X1 U11702 ( .A1(n9202), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9201) );
  MUX2_X1 U11703 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9201), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9203) );
  NAND2_X1 U11704 ( .A1(n9203), .A2(n9206), .ZN(n13833) );
  OAI222_X1 U11705 ( .A1(n14276), .A2(n7532), .B1(n14270), .B2(n9858), .C1(
        P1_U3086), .C2(n13833), .ZN(P1_U3352) );
  AND2_X1 U11706 ( .A1(n11542), .A2(P2_U3088), .ZN(n13668) );
  INV_X2 U11707 ( .A(n13668), .ZN(n13666) );
  INV_X1 U11708 ( .A(n9869), .ZN(n9210) );
  OAI222_X1 U11709 ( .A1(n13671), .A2(n9204), .B1(n13666), .B2(n9210), .C1(
        P2_U3088), .C2(n9558), .ZN(P2_U3323) );
  INV_X1 U11710 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9211) );
  NAND2_X1 U11711 ( .A1(n9206), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9205) );
  MUX2_X1 U11712 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9205), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n9208) );
  INV_X1 U11713 ( .A(n9841), .ZN(n9207) );
  AND2_X1 U11714 ( .A1(n9208), .A2(n9207), .ZN(n14658) );
  INV_X1 U11715 ( .A(n14658), .ZN(n9209) );
  OAI222_X1 U11716 ( .A1(n14276), .A2(n9211), .B1(n14270), .B2(n9210), .C1(
        P1_U3086), .C2(n9209), .ZN(P1_U3351) );
  OAI222_X1 U11717 ( .A1(P2_U3088), .A2(n9546), .B1(n13671), .B2(n9212), .C1(
        n13666), .C2(n9680), .ZN(P2_U3326) );
  OAI222_X1 U11718 ( .A1(n13671), .A2(n9213), .B1(n13666), .B2(n9724), .C1(
        P2_U3088), .C2(n9525), .ZN(P2_U3325) );
  OAI222_X1 U11719 ( .A1(n13671), .A2(n9214), .B1(n13666), .B2(n9858), .C1(
        P2_U3088), .C2(n9512), .ZN(P2_U3324) );
  INV_X1 U11720 ( .A(n9894), .ZN(n9219) );
  NOR2_X1 U11721 ( .A1(n9841), .A2(n9235), .ZN(n9215) );
  MUX2_X1 U11722 ( .A(n9235), .B(n9215), .S(P1_IR_REG_5__SCAN_IN), .Z(n9217)
         );
  OR2_X1 U11723 ( .A1(n9217), .A2(n9261), .ZN(n9330) );
  OAI222_X1 U11724 ( .A1(n14276), .A2(n9218), .B1(n14270), .B2(n9219), .C1(
        P1_U3086), .C2(n9330), .ZN(P1_U3350) );
  INV_X1 U11725 ( .A(n9563), .ZN(n9572) );
  OAI222_X1 U11726 ( .A1(n13671), .A2(n9220), .B1(n13666), .B2(n9219), .C1(
        P2_U3088), .C2(n9572), .ZN(P2_U3322) );
  NOR2_X2 U11727 ( .A1(n11542), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14397) );
  NAND2_X1 U11728 ( .A1(n11542), .A2(P3_U3151), .ZN(n12995) );
  INV_X1 U11729 ( .A(n12995), .ZN(n14396) );
  AOI222_X1 U11730 ( .A1(n9221), .A2(n14397), .B1(SI_9_), .B2(n14396), .C1(
        n10994), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9222) );
  INV_X1 U11731 ( .A(n9222), .ZN(P3_U3286) );
  AOI222_X1 U11732 ( .A1(n9223), .A2(n14397), .B1(SI_11_), .B2(n14396), .C1(
        n11076), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9224) );
  INV_X1 U11733 ( .A(n9224), .ZN(P3_U3284) );
  AOI222_X1 U11734 ( .A1(n9225), .A2(n14397), .B1(SI_10_), .B2(n14396), .C1(
        n14967), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9226) );
  INV_X1 U11735 ( .A(n9226), .ZN(P3_U3285) );
  AOI222_X1 U11736 ( .A1(n9227), .A2(n14397), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9931), .C1(SI_2_), .C2(n14396), .ZN(n9228) );
  INV_X1 U11737 ( .A(n9228), .ZN(P3_U3293) );
  AOI222_X1 U11738 ( .A1(n9229), .A2(n14397), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9941), .C1(SI_4_), .C2(n14396), .ZN(n9230) );
  INV_X1 U11739 ( .A(n9230), .ZN(P3_U3291) );
  AOI222_X1 U11740 ( .A1(n9231), .A2(n14397), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10203), .C1(SI_5_), .C2(n14396), .ZN(n9232) );
  INV_X1 U11741 ( .A(n9232), .ZN(P3_U3290) );
  AOI222_X1 U11742 ( .A1(n9233), .A2(n14397), .B1(n7145), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_7_), .C2(n14396), .ZN(n9234) );
  INV_X1 U11743 ( .A(n9234), .ZN(P3_U3288) );
  INV_X1 U11744 ( .A(n10104), .ZN(n9238) );
  OR2_X1 U11745 ( .A1(n9261), .A2(n9235), .ZN(n9236) );
  XNOR2_X1 U11746 ( .A(n9236), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10105) );
  INV_X1 U11747 ( .A(n10105), .ZN(n9350) );
  OAI222_X1 U11748 ( .A1(n14276), .A2(n9237), .B1(n14270), .B2(n9238), .C1(
        P1_U3086), .C2(n9350), .ZN(P1_U3349) );
  INV_X1 U11749 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9239) );
  INV_X1 U11750 ( .A(n9468), .ZN(n14792) );
  OAI222_X1 U11751 ( .A1(n13671), .A2(n9239), .B1(n13666), .B2(n9238), .C1(
        P2_U3088), .C2(n14792), .ZN(P2_U3321) );
  INV_X1 U11752 ( .A(n9254), .ZN(n9240) );
  NAND2_X1 U11753 ( .A1(n9240), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14274) );
  INV_X1 U11754 ( .A(n14274), .ZN(n9241) );
  OR2_X1 U11755 ( .A1(n9850), .A2(n9241), .ZN(n9305) );
  XNOR2_X1 U11756 ( .A(n9242), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9609) );
  NAND3_X1 U11757 ( .A1(n9245), .A2(n9244), .A3(n9243), .ZN(n9246) );
  NAND2_X1 U11758 ( .A1(n9609), .A2(n14279), .ZN(n11377) );
  INV_X1 U11759 ( .A(n11377), .ZN(n9713) );
  NAND2_X1 U11760 ( .A1(n9251), .A2(n9252), .ZN(n9613) );
  AOI21_X1 U11761 ( .B1(n9713), .B2(n9254), .A(n11501), .ZN(n9304) );
  INV_X1 U11762 ( .A(n9304), .ZN(n9255) );
  AND2_X1 U11763 ( .A1(n9305), .A2(n9255), .ZN(n14633) );
  NOR2_X1 U11764 ( .A1(n14633), .A2(P1_U4016), .ZN(P1_U3085) );
  OAI222_X1 U11765 ( .A1(n12997), .A2(n9257), .B1(n12995), .B2(n9256), .C1(
        P3_U3151), .C2(n9778), .ZN(P3_U3294) );
  OAI222_X1 U11766 ( .A1(n12997), .A2(n9259), .B1(n12995), .B2(n9258), .C1(
        P3_U3151), .C2(n10525), .ZN(P3_U3289) );
  INV_X1 U11767 ( .A(n10325), .ZN(n9265) );
  NAND2_X1 U11768 ( .A1(n9261), .A2(n9260), .ZN(n9282) );
  NAND2_X1 U11769 ( .A1(n9282), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9262) );
  XNOR2_X1 U11770 ( .A(n9262), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10326) );
  INV_X1 U11771 ( .A(n10326), .ZN(n9356) );
  OAI222_X1 U11772 ( .A1(n14276), .A2(n9263), .B1(n14270), .B2(n9265), .C1(
        P1_U3086), .C2(n9356), .ZN(P1_U3348) );
  INV_X1 U11773 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9266) );
  INV_X1 U11774 ( .A(n13153), .ZN(n9264) );
  OAI222_X1 U11775 ( .A1(n13671), .A2(n9266), .B1(n13666), .B2(n9265), .C1(
        P2_U3088), .C2(n9264), .ZN(P2_U3320) );
  INV_X1 U11776 ( .A(n12514), .ZN(n11083) );
  OAI222_X1 U11777 ( .A1(P3_U3151), .A2(n11083), .B1(n12995), .B2(n9268), .C1(
        n12997), .C2(n9267), .ZN(P3_U3283) );
  OAI222_X1 U11778 ( .A1(P3_U3151), .A2(n10716), .B1(n12995), .B2(n9270), .C1(
        n12997), .C2(n9269), .ZN(P3_U3287) );
  NAND2_X1 U11779 ( .A1(n10055), .A2(n12981), .ZN(n9271) );
  OAI21_X1 U11780 ( .B1(n15222), .B2(n12981), .A(n9271), .ZN(P3_U3377) );
  NAND2_X1 U11781 ( .A1(n9273), .A2(P1_B_REG_SCAN_IN), .ZN(n9276) );
  INV_X1 U11782 ( .A(n14267), .ZN(n9278) );
  OAI21_X1 U11783 ( .B1(n9273), .B2(P1_B_REG_SCAN_IN), .A(n9278), .ZN(n9274)
         );
  INV_X1 U11784 ( .A(n9274), .ZN(n9275) );
  INV_X1 U11785 ( .A(n14708), .ZN(n14707) );
  NAND2_X1 U11786 ( .A1(n9273), .A2(n14267), .ZN(n9607) );
  OAI22_X1 U11787 ( .A1(n14707), .A2(P1_D_REG_0__SCAN_IN), .B1(n9592), .B2(
        n9607), .ZN(n9277) );
  INV_X1 U11788 ( .A(n9277), .ZN(P1_U3445) );
  OR2_X1 U11789 ( .A1(n9272), .A2(n9278), .ZN(n9603) );
  OAI22_X1 U11790 ( .A1(n14707), .A2(P1_D_REG_1__SCAN_IN), .B1(n9592), .B2(
        n9603), .ZN(n9279) );
  INV_X1 U11791 ( .A(n9279), .ZN(P1_U3446) );
  INV_X1 U11792 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9281) );
  INV_X1 U11793 ( .A(n10310), .ZN(n9284) );
  INV_X1 U11794 ( .A(n13168), .ZN(n9280) );
  OAI222_X1 U11795 ( .A1(n13671), .A2(n9281), .B1(n13666), .B2(n9284), .C1(
        P2_U3088), .C2(n9280), .ZN(P2_U3319) );
  NAND2_X1 U11796 ( .A1(n9287), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9283) );
  XNOR2_X1 U11797 ( .A(n9283), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10311) );
  INV_X1 U11798 ( .A(n10311), .ZN(n9408) );
  OAI222_X1 U11799 ( .A1(n14276), .A2(n15155), .B1(n14270), .B2(n9284), .C1(
        P1_U3086), .C2(n9408), .ZN(P1_U3347) );
  AND2_X1 U11800 ( .A1(n9286), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U11801 ( .A1(n9286), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U11802 ( .A1(n9286), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U11803 ( .A1(n9286), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U11804 ( .A1(n9286), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U11805 ( .A1(n9286), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U11806 ( .A1(n9286), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U11807 ( .A1(n9286), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U11808 ( .A1(n9286), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U11809 ( .A1(n9286), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U11810 ( .A1(n9286), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U11811 ( .A1(n9286), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U11812 ( .A1(n9286), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U11813 ( .A1(n9286), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U11814 ( .A1(n9286), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U11815 ( .A1(n9286), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U11816 ( .A1(n9286), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U11817 ( .A1(n9286), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U11818 ( .A1(n9286), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U11819 ( .A1(n9286), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U11820 ( .A1(n9286), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U11821 ( .A1(n9286), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U11822 ( .A1(n9286), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U11823 ( .A1(n9286), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U11824 ( .A1(n9286), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U11825 ( .A1(n9286), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U11826 ( .A1(n9286), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U11827 ( .A1(n9286), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U11828 ( .A1(n9286), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U11829 ( .A1(n9286), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  INV_X1 U11830 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n15190) );
  INV_X1 U11831 ( .A(n10474), .ZN(n9291) );
  INV_X1 U11832 ( .A(n13186), .ZN(n9449) );
  OAI222_X1 U11833 ( .A1(n13671), .A2(n15190), .B1(n13666), .B2(n9291), .C1(
        P2_U3088), .C2(n9449), .ZN(P2_U3318) );
  OR2_X1 U11834 ( .A1(n9342), .A2(n9235), .ZN(n9289) );
  OR2_X1 U11835 ( .A1(n9289), .A2(n9288), .ZN(n9290) );
  NAND2_X1 U11836 ( .A1(n9289), .A2(n9288), .ZN(n9293) );
  INV_X1 U11837 ( .A(n10475), .ZN(n9398) );
  OAI222_X1 U11838 ( .A1(n14276), .A2(n9292), .B1(n14270), .B2(n9291), .C1(
        P1_U3086), .C2(n9398), .ZN(P1_U3346) );
  INV_X1 U11839 ( .A(n10739), .ZN(n9300) );
  NAND2_X1 U11840 ( .A1(n9293), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9294) );
  XNOR2_X1 U11841 ( .A(n9294), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10740) );
  AOI22_X1 U11842 ( .A1(n10740), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9295), .ZN(n9296) );
  OAI21_X1 U11843 ( .B1(n9300), .B2(n14270), .A(n9296), .ZN(P1_U3345) );
  INV_X1 U11844 ( .A(n12511), .ZN(n14980) );
  INV_X1 U11845 ( .A(n9297), .ZN(n9298) );
  OAI222_X1 U11846 ( .A1(P3_U3151), .A2(n14980), .B1(n12995), .B2(n9299), .C1(
        n12997), .C2(n9298), .ZN(P3_U3282) );
  INV_X1 U11847 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9301) );
  INV_X1 U11848 ( .A(n9476), .ZN(n9500) );
  OAI222_X1 U11849 ( .A1(n13671), .A2(n9301), .B1(n13666), .B2(n9300), .C1(
        P2_U3088), .C2(n9500), .ZN(P2_U3317) );
  OAI222_X1 U11850 ( .A1(n12527), .A2(P3_U3151), .B1(n12997), .B2(n9303), .C1(
        n9302), .C2(n12995), .ZN(P3_U3281) );
  NAND2_X1 U11851 ( .A1(n9305), .A2(n9304), .ZN(n14635) );
  INV_X1 U11852 ( .A(n14262), .ZN(n13816) );
  INV_X1 U11853 ( .A(n14631), .ZN(n11719) );
  INV_X1 U11854 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9308) );
  MUX2_X1 U11855 ( .A(n9308), .B(P1_REG1_REG_5__SCAN_IN), .S(n9330), .Z(n9313)
         );
  INV_X1 U11856 ( .A(n9683), .ZN(n9315) );
  INV_X1 U11857 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9795) );
  MUX2_X1 U11858 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9795), .S(n9683), .Z(n9368)
         );
  NAND2_X1 U11859 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9369) );
  NOR2_X1 U11860 ( .A1(n9368), .A2(n9369), .ZN(n9367) );
  AOI21_X1 U11861 ( .B1(n9315), .B2(P1_REG1_REG_1__SCAN_IN), .A(n9367), .ZN(
        n13825) );
  INV_X1 U11862 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9746) );
  MUX2_X1 U11863 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9746), .S(n9726), .Z(n13824) );
  NOR2_X1 U11864 ( .A1(n13825), .A2(n13824), .ZN(n13837) );
  NOR2_X1 U11865 ( .A1(n9726), .A2(n9746), .ZN(n13832) );
  INV_X1 U11866 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9309) );
  MUX2_X1 U11867 ( .A(n9309), .B(P1_REG1_REG_3__SCAN_IN), .S(n13833), .Z(n9310) );
  OAI21_X1 U11868 ( .B1(n13837), .B2(n13832), .A(n9310), .ZN(n14649) );
  INV_X1 U11869 ( .A(n13833), .ZN(n9311) );
  NAND2_X1 U11870 ( .A1(n9311), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n14648) );
  INV_X1 U11871 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14778) );
  MUX2_X1 U11872 ( .A(n14778), .B(P1_REG1_REG_4__SCAN_IN), .S(n14658), .Z(
        n14647) );
  AOI21_X1 U11873 ( .B1(n14649), .B2(n14648), .A(n14647), .ZN(n14646) );
  AOI21_X1 U11874 ( .B1(n14658), .B2(P1_REG1_REG_4__SCAN_IN), .A(n14646), .ZN(
        n9312) );
  NAND2_X1 U11875 ( .A1(n9312), .A2(n9313), .ZN(n9326) );
  OAI21_X1 U11876 ( .B1(n9313), .B2(n9312), .A(n9326), .ZN(n9322) );
  OR3_X1 U11877 ( .A1(n14635), .A2(n14631), .A3(n14262), .ZN(n14666) );
  INV_X1 U11878 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9314) );
  MUX2_X1 U11879 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9314), .S(n9683), .Z(n9371)
         );
  NAND2_X1 U11880 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n13815) );
  NOR2_X1 U11881 ( .A1(n9371), .A2(n13815), .ZN(n9370) );
  AOI21_X1 U11882 ( .B1(n9315), .B2(P1_REG2_REG_1__SCAN_IN), .A(n9370), .ZN(
        n13823) );
  INV_X1 U11883 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10154) );
  MUX2_X1 U11884 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10154), .S(n9726), .Z(
        n13822) );
  OR2_X1 U11885 ( .A1(n13823), .A2(n13822), .ZN(n13840) );
  INV_X1 U11886 ( .A(n9726), .ZN(n13828) );
  NAND2_X1 U11887 ( .A1(n13828), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13839) );
  INV_X1 U11888 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9316) );
  MUX2_X1 U11889 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9316), .S(n13833), .Z(
        n13838) );
  AOI21_X1 U11890 ( .B1(n13840), .B2(n13839), .A(n13838), .ZN(n14645) );
  NOR2_X1 U11891 ( .A1(n13833), .A2(n9316), .ZN(n14639) );
  INV_X1 U11892 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9887) );
  MUX2_X1 U11893 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9887), .S(n14658), .Z(n9317) );
  OAI21_X1 U11894 ( .B1(n14645), .B2(n14639), .A(n9317), .ZN(n14642) );
  NAND2_X1 U11895 ( .A1(n14658), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9319) );
  INV_X1 U11896 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9329) );
  MUX2_X1 U11897 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9329), .S(n9330), .Z(n9318)
         );
  AOI21_X1 U11898 ( .B1(n14642), .B2(n9319), .A(n9318), .ZN(n9333) );
  AND3_X1 U11899 ( .A1(n14642), .A2(n9319), .A3(n9318), .ZN(n9320) );
  NOR3_X1 U11900 ( .A1(n14666), .A2(n9333), .A3(n9320), .ZN(n9321) );
  AOI21_X1 U11901 ( .B1(n14652), .B2(n9322), .A(n9321), .ZN(n9325) );
  NAND2_X1 U11902 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10374) );
  INV_X1 U11903 ( .A(n10374), .ZN(n9323) );
  AOI21_X1 U11904 ( .B1(n14633), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n9323), .ZN(
        n9324) );
  OAI211_X1 U11905 ( .C1(n9330), .C2(n14670), .A(n9325), .B(n9324), .ZN(
        P1_U3248) );
  INV_X1 U11906 ( .A(n9330), .ZN(n9895) );
  OAI21_X1 U11907 ( .B1(n9895), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9326), .ZN(
        n9328) );
  INV_X1 U11908 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14780) );
  MUX2_X1 U11909 ( .A(n14780), .B(P1_REG1_REG_6__SCAN_IN), .S(n10105), .Z(
        n9327) );
  NOR2_X1 U11910 ( .A1(n9328), .A2(n9327), .ZN(n9385) );
  AOI211_X1 U11911 ( .C1(n9328), .C2(n9327), .A(n14668), .B(n9385), .ZN(n9337)
         );
  NOR2_X1 U11912 ( .A1(n9330), .A2(n9329), .ZN(n9332) );
  INV_X1 U11913 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10122) );
  MUX2_X1 U11914 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10122), .S(n10105), .Z(
        n9331) );
  OAI21_X1 U11915 ( .B1(n9333), .B2(n9332), .A(n9331), .ZN(n9378) );
  INV_X1 U11916 ( .A(n9378), .ZN(n9335) );
  NOR3_X1 U11917 ( .A1(n9333), .A2(n9332), .A3(n9331), .ZN(n9334) );
  NOR3_X1 U11918 ( .A1(n14666), .A2(n9335), .A3(n9334), .ZN(n9336) );
  NOR2_X1 U11919 ( .A1(n9337), .A2(n9336), .ZN(n9340) );
  INV_X1 U11920 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9338) );
  NOR2_X1 U11921 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9338), .ZN(n10650) );
  AOI21_X1 U11922 ( .B1(n14633), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10650), .ZN(
        n9339) );
  OAI211_X1 U11923 ( .C1(n9350), .C2(n14670), .A(n9340), .B(n9339), .ZN(
        P1_U3249) );
  INV_X1 U11924 ( .A(n10826), .ZN(n9345) );
  NOR2_X1 U11925 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9341) );
  NAND2_X1 U11926 ( .A1(n9342), .A2(n9341), .ZN(n9420) );
  NAND2_X1 U11927 ( .A1(n9420), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9343) );
  XNOR2_X1 U11928 ( .A(n9343), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10827) );
  INV_X1 U11929 ( .A(n10827), .ZN(n9660) );
  OAI222_X1 U11930 ( .A1(n14276), .A2(n9344), .B1(n14270), .B2(n9345), .C1(
        P1_U3086), .C2(n9660), .ZN(P1_U3344) );
  INV_X1 U11931 ( .A(n9645), .ZN(n9484) );
  OAI222_X1 U11932 ( .A1(n13671), .A2(n9346), .B1(n13666), .B2(n9345), .C1(
        P2_U3088), .C2(n9484), .ZN(P2_U3316) );
  INV_X1 U11933 ( .A(n12553), .ZN(n14457) );
  INV_X1 U11934 ( .A(n9347), .ZN(n9349) );
  OAI222_X1 U11935 ( .A1(n14457), .A2(P3_U3151), .B1(n12997), .B2(n9349), .C1(
        n9348), .C2(n12995), .ZN(P3_U3280) );
  INV_X1 U11936 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n14782) );
  NOR2_X1 U11937 ( .A1(n9350), .A2(n14780), .ZN(n9380) );
  MUX2_X1 U11938 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n14782), .S(n10326), .Z(
        n9351) );
  OAI21_X1 U11939 ( .B1(n9385), .B2(n9380), .A(n9351), .ZN(n9383) );
  OAI21_X1 U11940 ( .B1(n14782), .B2(n9356), .A(n9383), .ZN(n9406) );
  INV_X1 U11941 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9352) );
  MUX2_X1 U11942 ( .A(n9352), .B(P1_REG1_REG_8__SCAN_IN), .S(n10311), .Z(n9407) );
  NOR2_X1 U11943 ( .A1(n9406), .A2(n9407), .ZN(n9405) );
  NOR2_X1 U11944 ( .A1(n10311), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9394) );
  INV_X1 U11945 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n14785) );
  MUX2_X1 U11946 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n14785), .S(n10475), .Z(
        n9395) );
  OAI21_X1 U11947 ( .B1(n9405), .B2(n9394), .A(n9395), .ZN(n9393) );
  OAI21_X1 U11948 ( .B1(n10475), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9393), .ZN(
        n9354) );
  INV_X1 U11949 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14788) );
  MUX2_X1 U11950 ( .A(n14788), .B(P1_REG1_REG_10__SCAN_IN), .S(n10740), .Z(
        n9353) );
  NOR2_X1 U11951 ( .A1(n9354), .A2(n9353), .ZN(n9578) );
  AOI211_X1 U11952 ( .C1(n9354), .C2(n9353), .A(n14668), .B(n9578), .ZN(n9366)
         );
  NAND2_X1 U11953 ( .A1(n10105), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9377) );
  INV_X1 U11954 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9355) );
  MUX2_X1 U11955 ( .A(n9355), .B(P1_REG2_REG_7__SCAN_IN), .S(n10326), .Z(n9376) );
  AOI21_X1 U11956 ( .B1(n9378), .B2(n9377), .A(n9376), .ZN(n9415) );
  NOR2_X1 U11957 ( .A1(n9356), .A2(n9355), .ZN(n9410) );
  INV_X1 U11958 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10338) );
  MUX2_X1 U11959 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10338), .S(n10311), .Z(
        n9357) );
  OAI21_X1 U11960 ( .B1(n9415), .B2(n9410), .A(n9357), .ZN(n9413) );
  NAND2_X1 U11961 ( .A1(n10311), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9391) );
  INV_X1 U11962 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n15094) );
  MUX2_X1 U11963 ( .A(n15094), .B(P1_REG2_REG_9__SCAN_IN), .S(n10475), .Z(
        n9390) );
  AOI21_X1 U11964 ( .B1(n9413), .B2(n9391), .A(n9390), .ZN(n9404) );
  NOR2_X1 U11965 ( .A1(n9398), .A2(n15094), .ZN(n9359) );
  INV_X1 U11966 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10757) );
  MUX2_X1 U11967 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10757), .S(n10740), .Z(
        n9358) );
  OAI21_X1 U11968 ( .B1(n9404), .B2(n9359), .A(n9358), .ZN(n9576) );
  INV_X1 U11969 ( .A(n9576), .ZN(n9361) );
  NOR3_X1 U11970 ( .A1(n9404), .A2(n9359), .A3(n9358), .ZN(n9360) );
  NOR3_X1 U11971 ( .A1(n9361), .A2(n9360), .A3(n14666), .ZN(n9365) );
  INV_X1 U11972 ( .A(n10740), .ZN(n9363) );
  NAND2_X1 U11973 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11262)
         );
  NAND2_X1 U11974 ( .A1(n14633), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n9362) );
  OAI211_X1 U11975 ( .C1(n14670), .C2(n9363), .A(n11262), .B(n9362), .ZN(n9364) );
  OR3_X1 U11976 ( .A1(n9366), .A2(n9365), .A3(n9364), .ZN(P1_U3253) );
  AOI211_X1 U11977 ( .C1(n9369), .C2(n9368), .A(n9367), .B(n14668), .ZN(n9373)
         );
  AOI211_X1 U11978 ( .C1(n13815), .C2(n9371), .A(n9370), .B(n14666), .ZN(n9372) );
  NOR2_X1 U11979 ( .A1(n9373), .A2(n9372), .ZN(n9375) );
  AOI22_X1 U11980 ( .A1(n14633), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9374) );
  OAI211_X1 U11981 ( .C1(n9683), .C2(n14670), .A(n9375), .B(n9374), .ZN(
        P1_U3244) );
  NAND3_X1 U11982 ( .A1(n9378), .A2(n9377), .A3(n9376), .ZN(n9379) );
  NAND2_X1 U11983 ( .A1(n14643), .A2(n9379), .ZN(n9389) );
  INV_X1 U11984 ( .A(n9380), .ZN(n9382) );
  MUX2_X1 U11985 ( .A(n14782), .B(P1_REG1_REG_7__SCAN_IN), .S(n10326), .Z(
        n9381) );
  NAND2_X1 U11986 ( .A1(n9382), .A2(n9381), .ZN(n9384) );
  OAI211_X1 U11987 ( .C1(n9385), .C2(n9384), .A(n9383), .B(n14652), .ZN(n9388)
         );
  INV_X1 U11988 ( .A(n14670), .ZN(n14657) );
  INV_X1 U11989 ( .A(n14633), .ZN(n14674) );
  INV_X1 U11990 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14296) );
  NAND2_X1 U11991 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10705) );
  OAI21_X1 U11992 ( .B1(n14674), .B2(n14296), .A(n10705), .ZN(n9386) );
  AOI21_X1 U11993 ( .B1(n10326), .B2(n14657), .A(n9386), .ZN(n9387) );
  OAI211_X1 U11994 ( .C1(n9415), .C2(n9389), .A(n9388), .B(n9387), .ZN(
        P1_U3250) );
  NAND3_X1 U11995 ( .A1(n9413), .A2(n9391), .A3(n9390), .ZN(n9392) );
  NAND2_X1 U11996 ( .A1(n9392), .A2(n14643), .ZN(n9403) );
  INV_X1 U11997 ( .A(n9393), .ZN(n9397) );
  NOR3_X1 U11998 ( .A1(n9405), .A2(n9395), .A3(n9394), .ZN(n9396) );
  OAI21_X1 U11999 ( .B1(n9397), .B2(n9396), .A(n14652), .ZN(n9402) );
  NOR2_X1 U12000 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11218), .ZN(n9400) );
  NOR2_X1 U12001 ( .A1(n14670), .A2(n9398), .ZN(n9399) );
  AOI211_X1 U12002 ( .C1(n14633), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n9400), .B(
        n9399), .ZN(n9401) );
  OAI211_X1 U12003 ( .C1(n9404), .C2(n9403), .A(n9402), .B(n9401), .ZN(
        P1_U3252) );
  AOI21_X1 U12004 ( .B1(n9407), .B2(n9406), .A(n9405), .ZN(n9418) );
  AND2_X1 U12005 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10928) );
  NOR2_X1 U12006 ( .A1(n14670), .A2(n9408), .ZN(n9409) );
  AOI211_X1 U12007 ( .C1(n14633), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10928), .B(
        n9409), .ZN(n9417) );
  INV_X1 U12008 ( .A(n9410), .ZN(n9412) );
  MUX2_X1 U12009 ( .A(n10338), .B(P1_REG2_REG_8__SCAN_IN), .S(n10311), .Z(
        n9411) );
  NAND2_X1 U12010 ( .A1(n9412), .A2(n9411), .ZN(n9414) );
  OAI211_X1 U12011 ( .C1(n9415), .C2(n9414), .A(n9413), .B(n14643), .ZN(n9416)
         );
  OAI211_X1 U12012 ( .C1(n9418), .C2(n14668), .A(n9417), .B(n9416), .ZN(
        P1_U3251) );
  INV_X1 U12013 ( .A(n10831), .ZN(n9422) );
  INV_X1 U12014 ( .A(n9954), .ZN(n9644) );
  OAI222_X1 U12015 ( .A1(n13671), .A2(n9419), .B1(n13666), .B2(n9422), .C1(
        P2_U3088), .C2(n9644), .ZN(P2_U3315) );
  NAND2_X1 U12016 ( .A1(n9421), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9672) );
  XNOR2_X1 U12017 ( .A(n9672), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10832) );
  INV_X1 U12018 ( .A(n10832), .ZN(n9969) );
  OAI222_X1 U12019 ( .A1(n14276), .A2(n9423), .B1(n14270), .B2(n9422), .C1(
        P1_U3086), .C2(n9969), .ZN(P1_U3343) );
  INV_X1 U12020 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n13178) );
  MUX2_X1 U12021 ( .A(n9424), .B(P2_REG1_REG_1__SCAN_IN), .S(n9546), .Z(n9426)
         );
  AND2_X1 U12022 ( .A1(n13673), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9425) );
  NAND2_X1 U12023 ( .A1(n9426), .A2(n9425), .ZN(n9536) );
  INV_X1 U12024 ( .A(n9546), .ZN(n9457) );
  NAND2_X1 U12025 ( .A1(n9457), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9514) );
  NAND2_X1 U12026 ( .A1(n9536), .A2(n9514), .ZN(n9429) );
  MUX2_X1 U12027 ( .A(n9427), .B(P2_REG1_REG_2__SCAN_IN), .S(n9525), .Z(n9428)
         );
  NAND2_X1 U12028 ( .A1(n9429), .A2(n9428), .ZN(n9516) );
  INV_X1 U12029 ( .A(n9525), .ZN(n9460) );
  NAND2_X1 U12030 ( .A1(n9460), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9502) );
  NAND2_X1 U12031 ( .A1(n9516), .A2(n9502), .ZN(n9432) );
  MUX2_X1 U12032 ( .A(n9430), .B(P2_REG1_REG_3__SCAN_IN), .S(n9512), .Z(n9431)
         );
  NAND2_X1 U12033 ( .A1(n9432), .A2(n9431), .ZN(n9553) );
  OR2_X1 U12034 ( .A1(n9512), .A2(n9430), .ZN(n9552) );
  NAND2_X1 U12035 ( .A1(n9553), .A2(n9552), .ZN(n9435) );
  INV_X1 U12036 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9433) );
  MUX2_X1 U12037 ( .A(n9433), .B(P2_REG1_REG_4__SCAN_IN), .S(n9558), .Z(n9434)
         );
  NAND2_X1 U12038 ( .A1(n9435), .A2(n9434), .ZN(n9566) );
  NAND2_X1 U12039 ( .A1(n9465), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9565) );
  NAND2_X1 U12040 ( .A1(n9566), .A2(n9565), .ZN(n9438) );
  INV_X1 U12041 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9436) );
  MUX2_X1 U12042 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9436), .S(n9563), .Z(n9437)
         );
  NAND2_X1 U12043 ( .A1(n9438), .A2(n9437), .ZN(n9568) );
  NAND2_X1 U12044 ( .A1(n9563), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9439) );
  NAND2_X1 U12045 ( .A1(n9568), .A2(n9439), .ZN(n14800) );
  MUX2_X1 U12046 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9440), .S(n9468), .Z(n14799) );
  NAND2_X1 U12047 ( .A1(n14800), .A2(n14799), .ZN(n14798) );
  NAND2_X1 U12048 ( .A1(n9468), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n13151) );
  NAND2_X1 U12049 ( .A1(n14798), .A2(n13151), .ZN(n9443) );
  INV_X1 U12050 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9441) );
  MUX2_X1 U12051 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9441), .S(n13153), .Z(n9442) );
  NAND2_X1 U12052 ( .A1(n9443), .A2(n9442), .ZN(n13171) );
  NAND2_X1 U12053 ( .A1(n13153), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n13170) );
  NAND2_X1 U12054 ( .A1(n13171), .A2(n13170), .ZN(n9446) );
  MUX2_X1 U12055 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9444), .S(n13168), .Z(n9445) );
  NAND2_X1 U12056 ( .A1(n9446), .A2(n9445), .ZN(n13173) );
  NAND2_X1 U12057 ( .A1(n13168), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9447) );
  NAND2_X1 U12058 ( .A1(n13173), .A2(n9447), .ZN(n13177) );
  MUX2_X1 U12059 ( .A(n13178), .B(P2_REG1_REG_9__SCAN_IN), .S(n13186), .Z(
        n9448) );
  NOR2_X1 U12060 ( .A1(n13177), .A2(n9448), .ZN(n13189) );
  AOI21_X1 U12061 ( .B1(n13178), .B2(n9449), .A(n13189), .ZN(n9495) );
  MUX2_X1 U12062 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9450), .S(n9476), .Z(n9494) );
  NAND2_X1 U12063 ( .A1(n9495), .A2(n9494), .ZN(n9493) );
  OAI21_X1 U12064 ( .B1(n9450), .B2(n9500), .A(n9493), .ZN(n9640) );
  XOR2_X1 U12065 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9645), .Z(n9639) );
  XNOR2_X1 U12066 ( .A(n9640), .B(n9639), .ZN(n9488) );
  INV_X1 U12067 ( .A(n12090), .ZN(n9454) );
  NAND2_X1 U12068 ( .A1(n12090), .A2(n9451), .ZN(n9452) );
  NAND2_X1 U12069 ( .A1(n9452), .A2(n7662), .ZN(n9453) );
  OAI21_X1 U12070 ( .B1(n9455), .B2(n9454), .A(n9453), .ZN(n9482) );
  OR2_X1 U12071 ( .A1(n9481), .A2(P2_U3088), .ZN(n13655) );
  INV_X1 U12072 ( .A(n13658), .ZN(n12133) );
  NOR2_X1 U12073 ( .A1(n13655), .A2(n12133), .ZN(n9456) );
  NAND2_X1 U12074 ( .A1(n9482), .A2(n9456), .ZN(n14812) );
  MUX2_X1 U12075 ( .A(n10274), .B(P2_REG2_REG_1__SCAN_IN), .S(n9546), .Z(n9540) );
  AND2_X1 U12076 ( .A1(n13673), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9541) );
  NAND2_X1 U12077 ( .A1(n9540), .A2(n9541), .ZN(n9539) );
  NAND2_X1 U12078 ( .A1(n9457), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9519) );
  NAND2_X1 U12079 ( .A1(n9539), .A2(n9519), .ZN(n9459) );
  MUX2_X1 U12080 ( .A(n15082), .B(P2_REG2_REG_2__SCAN_IN), .S(n9525), .Z(n9458) );
  NAND2_X1 U12081 ( .A1(n9459), .A2(n9458), .ZN(n9521) );
  NAND2_X1 U12082 ( .A1(n9460), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9506) );
  NAND2_X1 U12083 ( .A1(n9521), .A2(n9506), .ZN(n9463) );
  MUX2_X1 U12084 ( .A(n9461), .B(P2_REG2_REG_3__SCAN_IN), .S(n9512), .Z(n9462)
         );
  NAND2_X1 U12085 ( .A1(n9463), .A2(n9462), .ZN(n9508) );
  OR2_X1 U12086 ( .A1(n9512), .A2(n9461), .ZN(n9464) );
  NAND2_X1 U12087 ( .A1(n9508), .A2(n9464), .ZN(n9549) );
  MUX2_X1 U12088 ( .A(n10591), .B(P2_REG2_REG_4__SCAN_IN), .S(n9558), .Z(n9548) );
  NAND2_X1 U12089 ( .A1(n9549), .A2(n9548), .ZN(n9547) );
  NAND2_X1 U12090 ( .A1(n9465), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9466) );
  NAND2_X1 U12091 ( .A1(n9547), .A2(n9466), .ZN(n9561) );
  MUX2_X1 U12092 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10601), .S(n9563), .Z(n9560) );
  NAND2_X1 U12093 ( .A1(n9561), .A2(n9560), .ZN(n9559) );
  NAND2_X1 U12094 ( .A1(n9563), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9467) );
  NAND2_X1 U12095 ( .A1(n9559), .A2(n9467), .ZN(n14797) );
  MUX2_X1 U12096 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10611), .S(n9468), .Z(
        n14796) );
  NAND2_X1 U12097 ( .A1(n14797), .A2(n14796), .ZN(n14795) );
  NAND2_X1 U12098 ( .A1(n9468), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n13155) );
  NAND2_X1 U12099 ( .A1(n14795), .A2(n13155), .ZN(n9471) );
  MUX2_X1 U12100 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9469), .S(n13153), .Z(n9470) );
  NAND2_X1 U12101 ( .A1(n9471), .A2(n9470), .ZN(n13165) );
  NAND2_X1 U12102 ( .A1(n13153), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n13164) );
  NAND2_X1 U12103 ( .A1(n13165), .A2(n13164), .ZN(n9473) );
  MUX2_X1 U12104 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10576), .S(n13168), .Z(
        n9472) );
  NAND2_X1 U12105 ( .A1(n9473), .A2(n9472), .ZN(n13167) );
  NAND2_X1 U12106 ( .A1(n13168), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9474) );
  AND2_X1 U12107 ( .A1(n13167), .A2(n9474), .ZN(n13183) );
  MUX2_X1 U12108 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n13489), .S(n13186), .Z(
        n9475) );
  NAND2_X1 U12109 ( .A1(n13183), .A2(n9475), .ZN(n13181) );
  OR2_X1 U12110 ( .A1(n13186), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n13182) );
  NAND2_X1 U12111 ( .A1(n13181), .A2(n13182), .ZN(n9491) );
  MUX2_X1 U12112 ( .A(n13477), .B(P2_REG2_REG_10__SCAN_IN), .S(n9476), .Z(
        n9490) );
  NOR2_X1 U12113 ( .A1(n9491), .A2(n9490), .ZN(n9489) );
  AOI21_X1 U12114 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n9476), .A(n9489), .ZN(
        n9479) );
  MUX2_X1 U12115 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10979), .S(n9645), .Z(
        n9478) );
  INV_X1 U12116 ( .A(n9648), .ZN(n9477) );
  OAI21_X1 U12117 ( .B1(n9479), .B2(n9478), .A(n9477), .ZN(n9486) );
  NOR2_X1 U12118 ( .A1(n13655), .A2(n13658), .ZN(n9480) );
  NAND2_X1 U12119 ( .A1(n9482), .A2(n9480), .ZN(n14806) );
  AND2_X1 U12120 ( .A1(n9481), .A2(n9482), .ZN(n14791) );
  AND2_X1 U12121 ( .A1(n14791), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14822) );
  NAND2_X1 U12122 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10821)
         );
  OR2_X1 U12123 ( .A1(n9482), .A2(P2_U3088), .ZN(n13211) );
  INV_X1 U12124 ( .A(n13211), .ZN(n14820) );
  NAND2_X1 U12125 ( .A1(n14820), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n9483) );
  OAI211_X1 U12126 ( .C1(n10637), .C2(n9484), .A(n10821), .B(n9483), .ZN(n9485) );
  AOI21_X1 U12127 ( .B1(n9486), .B2(n14824), .A(n9485), .ZN(n9487) );
  OAI21_X1 U12128 ( .B1(n9488), .B2(n14812), .A(n9487), .ZN(P2_U3225) );
  AOI211_X1 U12129 ( .C1(n9491), .C2(n9490), .A(n14806), .B(n9489), .ZN(n9492)
         );
  INV_X1 U12130 ( .A(n9492), .ZN(n9499) );
  NAND2_X1 U12131 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n10679)
         );
  INV_X1 U12132 ( .A(n14812), .ZN(n14827) );
  OAI211_X1 U12133 ( .C1(n9495), .C2(n9494), .A(n14827), .B(n9493), .ZN(n9496)
         );
  NAND2_X1 U12134 ( .A1(n10679), .A2(n9496), .ZN(n9497) );
  AOI21_X1 U12135 ( .B1(n14820), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n9497), .ZN(
        n9498) );
  OAI211_X1 U12136 ( .C1(n10637), .C2(n9500), .A(n9499), .B(n9498), .ZN(
        P2_U3224) );
  MUX2_X1 U12137 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9430), .S(n9512), .Z(n9501)
         );
  NAND3_X1 U12138 ( .A1(n9516), .A2(n9502), .A3(n9501), .ZN(n9503) );
  NAND2_X1 U12139 ( .A1(n9553), .A2(n9503), .ZN(n9504) );
  INV_X1 U12140 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n15070) );
  OAI22_X1 U12141 ( .A1(n14812), .A2(n9504), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15070), .ZN(n9510) );
  MUX2_X1 U12142 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n9461), .S(n9512), .Z(n9505)
         );
  NAND3_X1 U12143 ( .A1(n9521), .A2(n9506), .A3(n9505), .ZN(n9507) );
  AND3_X1 U12144 ( .A1(n14824), .A2(n9508), .A3(n9507), .ZN(n9509) );
  AOI211_X1 U12145 ( .C1(n14820), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n9510), .B(
        n9509), .ZN(n9511) );
  OAI21_X1 U12146 ( .B1(n9512), .B2(n10637), .A(n9511), .ZN(P2_U3217) );
  MUX2_X1 U12147 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9427), .S(n9525), .Z(n9513)
         );
  NAND3_X1 U12148 ( .A1(n9536), .A2(n9514), .A3(n9513), .ZN(n9515) );
  NAND2_X1 U12149 ( .A1(n9516), .A2(n9515), .ZN(n9517) );
  OAI22_X1 U12150 ( .A1(n14812), .A2(n9517), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10288), .ZN(n9523) );
  MUX2_X1 U12151 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n15082), .S(n9525), .Z(n9518) );
  NAND3_X1 U12152 ( .A1(n9539), .A2(n9519), .A3(n9518), .ZN(n9520) );
  AND3_X1 U12153 ( .A1(n14824), .A2(n9521), .A3(n9520), .ZN(n9522) );
  AOI211_X1 U12154 ( .C1(n14820), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n9523), .B(
        n9522), .ZN(n9524) );
  OAI21_X1 U12155 ( .B1(n9525), .B2(n10637), .A(n9524), .ZN(P2_U3216) );
  OAI22_X1 U12156 ( .A1(n9527), .A2(n14806), .B1(n14812), .B2(n9526), .ZN(
        n9530) );
  NAND2_X1 U12157 ( .A1(n14827), .A2(n9526), .ZN(n9528) );
  OAI211_X1 U12158 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n14806), .A(n10637), .B(
        n9528), .ZN(n9529) );
  MUX2_X1 U12159 ( .A(n9530), .B(n9529), .S(n13673), .Z(n9533) );
  INV_X1 U12160 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9531) );
  OAI22_X1 U12161 ( .A1(n13211), .A2(n9531), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10268), .ZN(n9532) );
  OR2_X1 U12162 ( .A1(n9533), .A2(n9532), .ZN(P2_U3214) );
  INV_X1 U12163 ( .A(n13673), .ZN(n9535) );
  MUX2_X1 U12164 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9424), .S(n9546), .Z(n9534)
         );
  OAI21_X1 U12165 ( .B1(n9526), .B2(n9535), .A(n9534), .ZN(n9537) );
  NAND2_X1 U12166 ( .A1(n9537), .A2(n9536), .ZN(n9538) );
  OAI22_X1 U12167 ( .A1(n14812), .A2(n9538), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10275), .ZN(n9544) );
  OAI211_X1 U12168 ( .C1(n9541), .C2(n9540), .A(n14824), .B(n9539), .ZN(n9542)
         );
  INV_X1 U12169 ( .A(n9542), .ZN(n9543) );
  AOI211_X1 U12170 ( .C1(n14820), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n9544), .B(
        n9543), .ZN(n9545) );
  OAI21_X1 U12171 ( .B1(n9546), .B2(n10637), .A(n9545), .ZN(P2_U3215) );
  NAND2_X1 U12172 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10068) );
  OAI211_X1 U12173 ( .C1(n9549), .C2(n9548), .A(n14824), .B(n9547), .ZN(n9550)
         );
  NAND2_X1 U12174 ( .A1(n10068), .A2(n9550), .ZN(n9556) );
  MUX2_X1 U12175 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9433), .S(n9558), .Z(n9551)
         );
  NAND3_X1 U12176 ( .A1(n9553), .A2(n9552), .A3(n9551), .ZN(n9554) );
  AND3_X1 U12177 ( .A1(n14827), .A2(n9566), .A3(n9554), .ZN(n9555) );
  AOI211_X1 U12178 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n14820), .A(n9556), .B(
        n9555), .ZN(n9557) );
  OAI21_X1 U12179 ( .B1(n9558), .B2(n10637), .A(n9557), .ZN(P2_U3218) );
  NAND2_X1 U12180 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10090) );
  OAI211_X1 U12181 ( .C1(n9561), .C2(n9560), .A(n14824), .B(n9559), .ZN(n9562)
         );
  NAND2_X1 U12182 ( .A1(n10090), .A2(n9562), .ZN(n9570) );
  MUX2_X1 U12183 ( .A(n9436), .B(P2_REG1_REG_5__SCAN_IN), .S(n9563), .Z(n9564)
         );
  NAND3_X1 U12184 ( .A1(n9566), .A2(n9565), .A3(n9564), .ZN(n9567) );
  AND3_X1 U12185 ( .A1(n14827), .A2(n9568), .A3(n9567), .ZN(n9569) );
  AOI211_X1 U12186 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n14820), .A(n9570), .B(
        n9569), .ZN(n9571) );
  OAI21_X1 U12187 ( .B1(n9572), .B2(n10637), .A(n9571), .ZN(P2_U3219) );
  NAND2_X1 U12188 ( .A1(n10740), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9575) );
  INV_X1 U12189 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9573) );
  MUX2_X1 U12190 ( .A(n9573), .B(P1_REG2_REG_11__SCAN_IN), .S(n10827), .Z(
        n9574) );
  AOI21_X1 U12191 ( .B1(n9576), .B2(n9575), .A(n9574), .ZN(n9655) );
  NAND3_X1 U12192 ( .A1(n9576), .A2(n9575), .A3(n9574), .ZN(n9577) );
  NAND2_X1 U12193 ( .A1(n9577), .A2(n14643), .ZN(n9585) );
  INV_X1 U12194 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14585) );
  MUX2_X1 U12195 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n14585), .S(n10827), .Z(
        n9580) );
  AOI21_X1 U12196 ( .B1(n10740), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9578), .ZN(
        n9579) );
  NAND2_X1 U12197 ( .A1(n9579), .A2(n9580), .ZN(n9664) );
  OAI21_X1 U12198 ( .B1(n9580), .B2(n9579), .A(n9664), .ZN(n9581) );
  NAND2_X1 U12199 ( .A1(n9581), .A2(n14652), .ZN(n9584) );
  INV_X1 U12200 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n15218) );
  NAND2_X1 U12201 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14528)
         );
  OAI21_X1 U12202 ( .B1(n14674), .B2(n15218), .A(n14528), .ZN(n9582) );
  AOI21_X1 U12203 ( .B1(n10827), .B2(n14657), .A(n9582), .ZN(n9583) );
  OAI211_X1 U12204 ( .C1(n9655), .C2(n9585), .A(n9584), .B(n9583), .ZN(
        P1_U3254) );
  MUX2_X1 U12205 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9586), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n9587) );
  NAND2_X1 U12206 ( .A1(n9588), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9589) );
  XNOR2_X2 U12207 ( .A(n9589), .B(P1_IR_REG_19__SCAN_IN), .ZN(n11703) );
  AND2_X1 U12208 ( .A1(n11375), .A2(n14022), .ZN(n9590) );
  OR2_X1 U12209 ( .A1(n11377), .A2(n9590), .ZN(n9591) );
  NAND2_X1 U12210 ( .A1(n9591), .A2(n9685), .ZN(n10178) );
  NOR4_X1 U12211 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n9601) );
  NOR4_X1 U12212 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n9600) );
  OR4_X1 U12213 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n9598) );
  NOR4_X1 U12214 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9596) );
  NOR4_X1 U12215 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n9595) );
  NOR4_X1 U12216 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9594) );
  NOR4_X1 U12217 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9593) );
  NAND4_X1 U12218 ( .A1(n9596), .A2(n9595), .A3(n9594), .A4(n9593), .ZN(n9597)
         );
  NOR4_X1 U12219 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9598), .A4(n9597), .ZN(n9599) );
  AND3_X1 U12220 ( .A1(n9601), .A2(n9600), .A3(n9599), .ZN(n9602) );
  OR2_X1 U12221 ( .A1(n9606), .A2(n9602), .ZN(n9703) );
  NAND2_X1 U12222 ( .A1(n11720), .A2(n9703), .ZN(n9712) );
  OR2_X1 U12223 ( .A1(n9606), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9604) );
  AND2_X1 U12224 ( .A1(n9604), .A2(n9603), .ZN(n9704) );
  INV_X1 U12225 ( .A(n9704), .ZN(n9711) );
  NAND2_X1 U12226 ( .A1(n11375), .A2(n11703), .ZN(n9852) );
  INV_X1 U12227 ( .A(n9852), .ZN(n14697) );
  NAND2_X1 U12228 ( .A1(n7289), .A2(n14697), .ZN(n9848) );
  NAND2_X1 U12229 ( .A1(n9711), .A2(n9848), .ZN(n9605) );
  OR2_X1 U12230 ( .A1(n9712), .A2(n9605), .ZN(n9722) );
  OR2_X1 U12231 ( .A1(n9606), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9608) );
  INV_X1 U12232 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9635) );
  NAND2_X1 U12233 ( .A1(n14022), .A2(n14279), .ZN(n9610) );
  INV_X1 U12234 ( .A(n11369), .ZN(n9611) );
  OR2_X1 U12235 ( .A1(n9684), .A2(n9611), .ZN(n9612) );
  NAND2_X1 U12236 ( .A1(n11217), .A2(n9612), .ZN(n9853) );
  OR2_X1 U12237 ( .A1(n9852), .A2(n14279), .ZN(n14730) );
  NAND2_X1 U12238 ( .A1(n9609), .A2(n11379), .ZN(n11665) );
  NOR2_X2 U12239 ( .A1(n9613), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n9616) );
  NAND2_X1 U12240 ( .A1(n9616), .A2(n9614), .ZN(n14249) );
  XNOR2_X2 U12241 ( .A(n9615), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9619) );
  INV_X1 U12242 ( .A(n9619), .ZN(n14256) );
  AND2_X2 U12243 ( .A1(n14256), .A2(n14258), .ZN(n9733) );
  NAND2_X1 U12244 ( .A1(n9733), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9623) );
  AND2_X2 U12245 ( .A1(n14256), .A2(n9618), .ZN(n9899) );
  NAND2_X1 U12246 ( .A1(n9899), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9622) );
  AND2_X2 U12247 ( .A1(n9619), .A2(n14258), .ZN(n9734) );
  NAND2_X1 U12248 ( .A1(n9734), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9621) );
  AND2_X2 U12249 ( .A1(n9619), .A2(n9618), .ZN(n10112) );
  NAND2_X1 U12250 ( .A1(n10112), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9620) );
  OAI21_X1 U12251 ( .B1(n11542), .B2(n9625), .A(n9624), .ZN(n9626) );
  AND2_X1 U12252 ( .A1(n9627), .A2(n9626), .ZN(n14280) );
  MUX2_X1 U12253 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14280), .S(n11545), .Z(n11331) );
  INV_X1 U12254 ( .A(n11331), .ZN(n11388) );
  NAND2_X1 U12255 ( .A1(n9693), .A2(n11331), .ZN(n9779) );
  INV_X1 U12256 ( .A(n9779), .ZN(n9628) );
  AOI21_X1 U12257 ( .B1(n9731), .B2(n11388), .A(n9628), .ZN(n14698) );
  OAI21_X1 U12258 ( .B1(n14774), .B2(n14763), .A(n14698), .ZN(n9633) );
  NAND2_X1 U12259 ( .A1(n11331), .A2(n7289), .ZN(n14696) );
  NAND2_X1 U12260 ( .A1(n10112), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9632) );
  NAND2_X1 U12261 ( .A1(n9899), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9631) );
  NAND2_X1 U12262 ( .A1(n9734), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9629) );
  NAND2_X1 U12263 ( .A1(n13813), .A2(n14745), .ZN(n14695) );
  NAND3_X1 U12264 ( .A1(n9633), .A2(n14696), .A3(n14695), .ZN(n14232) );
  NAND2_X1 U12265 ( .A1(n14232), .A2(n6444), .ZN(n9634) );
  OAI21_X1 U12266 ( .B1(n6444), .B2(n9635), .A(n9634), .ZN(P1_U3459) );
  INV_X2 U12267 ( .A(P3_U3897), .ZN(n12500) );
  NAND2_X1 U12268 ( .A1(n12500), .A2(P3_DATAO_REG_11__SCAN_IN), .ZN(n9636) );
  OAI21_X1 U12269 ( .B1(n12859), .B2(n12500), .A(n9636), .ZN(P3_U3502) );
  INV_X1 U12270 ( .A(n12591), .ZN(n12585) );
  OAI222_X1 U12271 ( .A1(P3_U3151), .A2(n12585), .B1(n12995), .B2(n15122), 
        .C1(n12997), .C2(n9637), .ZN(P3_U3278) );
  INV_X1 U12272 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n15201) );
  NAND2_X1 U12273 ( .A1(n12792), .A2(P3_U3897), .ZN(n9638) );
  OAI21_X1 U12274 ( .B1(P3_U3897), .B2(n15201), .A(n9638), .ZN(P3_U3508) );
  AOI22_X1 U12275 ( .A1(n9640), .A2(n9639), .B1(P2_REG1_REG_11__SCAN_IN), .B2(
        n9645), .ZN(n9642) );
  INV_X1 U12276 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n15112) );
  MUX2_X1 U12277 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n15112), .S(n9954), .Z(
        n9641) );
  NAND2_X1 U12278 ( .A1(n9642), .A2(n9641), .ZN(n9953) );
  OAI21_X1 U12279 ( .B1(n9642), .B2(n9641), .A(n9953), .ZN(n9652) );
  AND2_X1 U12280 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n10965) );
  AOI21_X1 U12281 ( .B1(n14820), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n10965), 
        .ZN(n9643) );
  OAI21_X1 U12282 ( .B1(n10637), .B2(n9644), .A(n9643), .ZN(n9651) );
  NOR2_X1 U12283 ( .A1(n9645), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9646) );
  MUX2_X1 U12284 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11165), .S(n9954), .Z(
        n9647) );
  OAI21_X1 U12285 ( .B1(n9648), .B2(n9646), .A(n9647), .ZN(n9951) );
  OR3_X1 U12286 ( .A1(n9648), .A2(n9647), .A3(n9646), .ZN(n9649) );
  AOI21_X1 U12287 ( .B1(n9951), .B2(n9649), .A(n14806), .ZN(n9650) );
  AOI211_X1 U12288 ( .C1(n14827), .C2(n9652), .A(n9651), .B(n9650), .ZN(n9653)
         );
  INV_X1 U12289 ( .A(n9653), .ZN(P2_U3226) );
  INV_X1 U12290 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n15177) );
  NAND2_X1 U12291 ( .A1(n12353), .A2(P3_U3897), .ZN(n9654) );
  OAI21_X1 U12292 ( .B1(P3_U3897), .B2(n15177), .A(n9654), .ZN(P3_U3495) );
  INV_X1 U12293 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9970) );
  MUX2_X1 U12294 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n9970), .S(n10832), .Z(
        n9656) );
  INV_X1 U12295 ( .A(n9656), .ZN(n9659) );
  AOI21_X1 U12296 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n10827), .A(n9655), .ZN(
        n9657) );
  INV_X1 U12297 ( .A(n9657), .ZN(n9658) );
  AND2_X1 U12298 ( .A1(n9657), .A2(n9656), .ZN(n9968) );
  AOI21_X1 U12299 ( .B1(n9659), .B2(n9658), .A(n9968), .ZN(n9670) );
  NAND2_X1 U12300 ( .A1(n9660), .A2(n14585), .ZN(n9662) );
  INV_X1 U12301 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9661) );
  MUX2_X1 U12302 ( .A(n9661), .B(P1_REG1_REG_12__SCAN_IN), .S(n10832), .Z(
        n9663) );
  AOI21_X1 U12303 ( .B1(n9664), .B2(n9662), .A(n9663), .ZN(n9967) );
  AND3_X1 U12304 ( .A1(n9664), .A2(n9663), .A3(n9662), .ZN(n9665) );
  OAI21_X1 U12305 ( .B1(n9967), .B2(n9665), .A(n14652), .ZN(n9669) );
  NOR2_X1 U12306 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10835), .ZN(n9667) );
  NOR2_X1 U12307 ( .A1(n14670), .A2(n9969), .ZN(n9666) );
  AOI211_X1 U12308 ( .C1(n14633), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n9667), .B(
        n9666), .ZN(n9668) );
  OAI211_X1 U12309 ( .C1(n9670), .C2(n14666), .A(n9669), .B(n9668), .ZN(
        P1_U3255) );
  INV_X1 U12310 ( .A(n11026), .ZN(n9675) );
  INV_X1 U12311 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9671) );
  NAND2_X1 U12312 ( .A1(n9672), .A2(n9671), .ZN(n9673) );
  NAND2_X1 U12313 ( .A1(n9673), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9945) );
  INV_X1 U12314 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9944) );
  XNOR2_X1 U12315 ( .A(n9945), .B(n9944), .ZN(n11027) );
  OAI222_X1 U12316 ( .A1(n14276), .A2(n15111), .B1(n14270), .B2(n9675), .C1(
        P1_U3086), .C2(n11027), .ZN(P1_U3342) );
  INV_X1 U12317 ( .A(n14805), .ZN(n9674) );
  OAI222_X1 U12318 ( .A1(n13671), .A2(n9676), .B1(n13666), .B2(n9675), .C1(
        P2_U3088), .C2(n9674), .ZN(P2_U3314) );
  OR2_X4 U12319 ( .A1(n9684), .A2(n9677), .ZN(n11867) );
  OR2_X1 U12320 ( .A1(n9859), .A2(n9678), .ZN(n9682) );
  OR2_X1 U12321 ( .A1(n9856), .A2(n9680), .ZN(n9681) );
  OAI211_X2 U12322 ( .C1(n11545), .C2(n9683), .A(n9682), .B(n9681), .ZN(n14109) );
  AND2_X4 U12323 ( .A1(n9685), .A2(n9684), .ZN(n11858) );
  OAI22_X1 U12324 ( .A1(n11334), .A2(n11867), .B1(n9708), .B2(n10169), .ZN(
        n9686) );
  XNOR2_X1 U12325 ( .A(n9686), .B(n11217), .ZN(n9803) );
  NAND2_X1 U12326 ( .A1(n10361), .A2(n14109), .ZN(n9688) );
  NAND2_X1 U12327 ( .A1(n9689), .A2(n9688), .ZN(n9802) );
  INV_X1 U12328 ( .A(n9802), .ZN(n9690) );
  OR2_X1 U12329 ( .A1(n9731), .A2(n9799), .ZN(n9692) );
  AOI22_X1 U12330 ( .A1(n10361), .A2(n11331), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n9677), .ZN(n9691) );
  AND2_X1 U12331 ( .A1(n9692), .A2(n9691), .ZN(n11329) );
  AOI22_X1 U12332 ( .A1(n11331), .A2(n11858), .B1(n9677), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9694) );
  AND2_X1 U12333 ( .A1(n9695), .A2(n9694), .ZN(n11328) );
  INV_X1 U12334 ( .A(n11328), .ZN(n9696) );
  NAND2_X1 U12335 ( .A1(n11329), .A2(n9696), .ZN(n9698) );
  NAND2_X1 U12336 ( .A1(n11328), .A2(n11217), .ZN(n9697) );
  NAND2_X1 U12337 ( .A1(n9698), .A2(n9697), .ZN(n9699) );
  NAND2_X1 U12338 ( .A1(n7289), .A2(n11379), .ZN(n14019) );
  NAND2_X1 U12339 ( .A1(n7289), .A2(n11703), .ZN(n9700) );
  INV_X1 U12340 ( .A(n9850), .ZN(n9701) );
  OR2_X1 U12341 ( .A1(n9701), .A2(n9713), .ZN(n9702) );
  NOR2_X1 U12342 ( .A1(n14767), .A2(n9702), .ZN(n9706) );
  NAND3_X1 U12343 ( .A1(n9847), .A2(n9704), .A3(n9703), .ZN(n9707) );
  INV_X1 U12344 ( .A(n9707), .ZN(n9705) );
  NAND2_X1 U12345 ( .A1(n9707), .A2(n9848), .ZN(n10180) );
  AND2_X1 U12346 ( .A1(n10180), .A2(n9850), .ZN(n14618) );
  INV_X1 U12347 ( .A(n14525), .ZN(n14500) );
  NAND2_X1 U12348 ( .A1(n10180), .A2(n11720), .ZN(n11330) );
  INV_X1 U12349 ( .A(n11330), .ZN(n9710) );
  INV_X1 U12350 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9709) );
  OAI22_X1 U12351 ( .A1(n14500), .A2(n9708), .B1(n9710), .B2(n9709), .ZN(n9719) );
  NAND2_X1 U12352 ( .A1(n14625), .A2(n14766), .ZN(n14503) );
  NAND2_X1 U12353 ( .A1(n14625), .A2(n14745), .ZN(n14502) );
  NAND2_X1 U12354 ( .A1(n10112), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9717) );
  NAND2_X1 U12355 ( .A1(n9733), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9716) );
  NAND2_X1 U12356 ( .A1(n9734), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9715) );
  NAND4_X4 U12357 ( .A1(n9717), .A2(n9716), .A3(n9715), .A4(n9714), .ZN(n13812) );
  INV_X1 U12358 ( .A(n13812), .ZN(n9872) );
  OAI22_X1 U12359 ( .A1(n9731), .A2(n14503), .B1(n14502), .B2(n9872), .ZN(
        n9718) );
  AOI211_X1 U12360 ( .C1(n9720), .C2(n14527), .A(n9719), .B(n9718), .ZN(n9721)
         );
  INV_X1 U12361 ( .A(n9721), .ZN(P1_U3222) );
  NAND2_X1 U12362 ( .A1(n11334), .A2(n9708), .ZN(n9723) );
  NAND2_X1 U12363 ( .A1(n9781), .A2(n9723), .ZN(n9730) );
  OR2_X1 U12364 ( .A1(n9856), .A2(n9724), .ZN(n9729) );
  OR2_X1 U12365 ( .A1(n9859), .A2(n9725), .ZN(n9728) );
  OR2_X1 U12366 ( .A1(n11545), .A2(n9726), .ZN(n9727) );
  AND3_X2 U12367 ( .A1(n9729), .A2(n9728), .A3(n9727), .ZN(n11399) );
  OAI21_X1 U12368 ( .B1(n9730), .B2(n11677), .A(n9855), .ZN(n10158) );
  INV_X1 U12369 ( .A(n10158), .ZN(n9744) );
  NAND2_X1 U12370 ( .A1(n9731), .A2(n11331), .ZN(n11381) );
  NAND2_X1 U12371 ( .A1(n11383), .A2(n11381), .ZN(n11390) );
  OAI21_X1 U12372 ( .B1(n6581), .B2(n9732), .A(n9874), .ZN(n9739) );
  INV_X1 U12373 ( .A(n14766), .ZN(n14209) );
  INV_X1 U12374 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10145) );
  NAND2_X1 U12375 ( .A1(n10112), .A2(n10145), .ZN(n9738) );
  NAND2_X1 U12376 ( .A1(n11599), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9737) );
  NAND2_X1 U12377 ( .A1(n9734), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9736) );
  NAND2_X1 U12378 ( .A1(n9899), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9735) );
  AND4_X2 U12379 ( .A1(n9738), .A2(n9737), .A3(n9736), .A4(n9735), .ZN(n10172)
         );
  OAI22_X1 U12380 ( .A1(n11334), .A2(n14209), .B1(n10172), .B2(n14420), .ZN(
        n9808) );
  AOI21_X1 U12381 ( .B1(n9739), .B2(n14763), .A(n9808), .ZN(n10161) );
  OR2_X1 U12382 ( .A1(n14109), .A2(n11331), .ZN(n9783) );
  INV_X1 U12383 ( .A(n9783), .ZN(n9740) );
  NAND2_X1 U12384 ( .A1(n7375), .A2(n9783), .ZN(n9741) );
  NAND2_X1 U12385 ( .A1(n9741), .A2(n14686), .ZN(n9742) );
  NOR2_X1 U12386 ( .A1(n10144), .A2(n9742), .ZN(n10157) );
  AOI21_X1 U12387 ( .B1(n7375), .B2(n14767), .A(n10157), .ZN(n9743) );
  OAI211_X1 U12388 ( .C1(n9744), .C2(n14755), .A(n10161), .B(n9743), .ZN(n9747) );
  NAND2_X1 U12389 ( .A1(n9747), .A2(n14790), .ZN(n9745) );
  OAI21_X1 U12390 ( .B1(n14790), .B2(n9746), .A(n9745), .ZN(P1_U3530) );
  INV_X1 U12391 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9749) );
  NAND2_X1 U12392 ( .A1(n9747), .A2(n6444), .ZN(n9748) );
  OAI21_X1 U12393 ( .B1(n6444), .B2(n9749), .A(n9748), .ZN(P1_U3465) );
  INV_X1 U12394 ( .A(n12606), .ZN(n12594) );
  OAI222_X1 U12395 ( .A1(P3_U3151), .A2(n12594), .B1(n12995), .B2(n9751), .C1(
        n12997), .C2(n9750), .ZN(P3_U3277) );
  NAND2_X1 U12396 ( .A1(n12460), .A2(n9754), .ZN(n9752) );
  AND2_X1 U12397 ( .A1(n9753), .A2(n9752), .ZN(n9767) );
  INV_X1 U12398 ( .A(n9754), .ZN(n9755) );
  NAND2_X1 U12399 ( .A1(n9755), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12486) );
  NAND2_X1 U12400 ( .A1(n9756), .A2(n12486), .ZN(n9768) );
  NAND2_X1 U12401 ( .A1(n9767), .A2(n9768), .ZN(n9765) );
  MUX2_X1 U12402 ( .A(n9765), .B(n12500), .S(n12481), .Z(n14979) );
  INV_X1 U12403 ( .A(n14989), .ZN(n14896) );
  NAND2_X1 U12404 ( .A1(n15107), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9757) );
  NAND2_X1 U12405 ( .A1(n9812), .A2(n9757), .ZN(n9820) );
  OR3_X1 U12406 ( .A1(n8186), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        P3_IR_REG_1__SCAN_IN), .ZN(n9758) );
  AOI21_X1 U12407 ( .B1(n9820), .B2(n9758), .A(n9774), .ZN(n9760) );
  NAND2_X1 U12408 ( .A1(n9774), .A2(n9758), .ZN(n9819) );
  INV_X1 U12409 ( .A(n9819), .ZN(n9759) );
  OAI22_X1 U12410 ( .A1(n9760), .A2(n9759), .B1(n9820), .B2(
        P3_REG1_REG_1__SCAN_IN), .ZN(n9772) );
  INV_X1 U12411 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n15107) );
  AND2_X1 U12412 ( .A1(P3_REG2_REG_0__SCAN_IN), .A2(n15107), .ZN(n9762) );
  NAND2_X1 U12413 ( .A1(P3_REG2_REG_0__SCAN_IN), .A2(n9761), .ZN(n9814) );
  INV_X1 U12414 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10254) );
  NAND2_X1 U12415 ( .A1(n9763), .A2(n10254), .ZN(n9766) );
  AOI21_X1 U12416 ( .B1(n9815), .B2(n9766), .A(n14995), .ZN(n9771) );
  INV_X1 U12417 ( .A(n9767), .ZN(n9769) );
  AND2_X1 U12418 ( .A1(n9769), .A2(n9768), .ZN(n14972) );
  INV_X1 U12419 ( .A(n14972), .ZN(n14978) );
  INV_X1 U12420 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10246) );
  OAI22_X1 U12421 ( .A1(n14978), .A2(n7214), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10246), .ZN(n9770) );
  AOI211_X1 U12422 ( .C1(n14896), .C2(n9772), .A(n9771), .B(n9770), .ZN(n9777)
         );
  MUX2_X1 U12423 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n12602), .Z(n14899) );
  NOR2_X1 U12424 ( .A1(n14899), .A2(n15107), .ZN(n14898) );
  XNOR2_X1 U12425 ( .A(n9813), .B(n14898), .ZN(n9775) );
  NAND2_X1 U12426 ( .A1(n9775), .A2(n14945), .ZN(n9776) );
  OAI211_X1 U12427 ( .C1(n14979), .C2(n9778), .A(n9777), .B(n9776), .ZN(
        P3_U3183) );
  OR2_X1 U12428 ( .A1(n9779), .A2(n11675), .ZN(n9780) );
  NAND2_X1 U12429 ( .A1(n9781), .A2(n9780), .ZN(n14108) );
  INV_X1 U12430 ( .A(n14108), .ZN(n9793) );
  INV_X1 U12431 ( .A(n9853), .ZN(n14733) );
  NAND2_X1 U12432 ( .A1(n14108), .A2(n14733), .ZN(n9788) );
  NAND2_X1 U12433 ( .A1(n14109), .A2(n11331), .ZN(n9782) );
  AND2_X1 U12434 ( .A1(n9783), .A2(n9782), .ZN(n9789) );
  XNOR2_X1 U12435 ( .A(n11334), .B(n9789), .ZN(n9784) );
  MUX2_X1 U12436 ( .A(n9784), .B(n11675), .S(n9693), .Z(n9785) );
  NAND2_X1 U12437 ( .A1(n9785), .A2(n14763), .ZN(n9787) );
  AOI22_X1 U12438 ( .A1(n9693), .A2(n14766), .B1(n14745), .B2(n13812), .ZN(
        n9786) );
  NAND3_X1 U12439 ( .A1(n9788), .A2(n9787), .A3(n9786), .ZN(n14104) );
  INV_X1 U12440 ( .A(n14104), .ZN(n9792) );
  INV_X1 U12441 ( .A(n9789), .ZN(n9790) );
  NOR2_X1 U12442 ( .A1(n9790), .A2(n14572), .ZN(n14110) );
  AOI21_X1 U12443 ( .B1(n14109), .B2(n14767), .A(n14110), .ZN(n9791) );
  OAI211_X1 U12444 ( .C1(n9793), .C2(n14730), .A(n9792), .B(n9791), .ZN(n9796)
         );
  NAND2_X1 U12445 ( .A1(n9796), .A2(n14790), .ZN(n9794) );
  OAI21_X1 U12446 ( .B1(n14790), .B2(n9795), .A(n9794), .ZN(P1_U3529) );
  INV_X1 U12447 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9798) );
  NAND2_X1 U12448 ( .A1(n9796), .A2(n6444), .ZN(n9797) );
  OAI21_X1 U12449 ( .B1(n6444), .B2(n9798), .A(n9797), .ZN(P1_U3462) );
  OAI22_X1 U12450 ( .A1(n9872), .A2(n9799), .B1(n11399), .B2(n11867), .ZN(
        n10164) );
  NAND2_X1 U12451 ( .A1(n13812), .A2(n10361), .ZN(n9801) );
  OR2_X1 U12452 ( .A1(n11399), .A2(n10169), .ZN(n9800) );
  XOR2_X1 U12453 ( .A(n10164), .B(n10163), .Z(n9806) );
  NAND2_X1 U12454 ( .A1(n9805), .A2(n9806), .ZN(n10168) );
  OAI21_X1 U12455 ( .B1(n9806), .B2(n9805), .A(n10168), .ZN(n9807) );
  NAND2_X1 U12456 ( .A1(n9807), .A2(n14527), .ZN(n9810) );
  AOI22_X1 U12457 ( .A1(n14625), .A2(n9808), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n11330), .ZN(n9809) );
  OAI211_X1 U12458 ( .C1(n11399), .C2(n14500), .A(n9810), .B(n9809), .ZN(
        P1_U3237) );
  OAI222_X1 U12459 ( .A1(n12997), .A2(n9811), .B1(P3_U3151), .B2(n12612), .C1(
        n12995), .C2(n15087), .ZN(P3_U3276) );
  MUX2_X1 U12460 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12602), .Z(n9917) );
  XOR2_X1 U12461 ( .A(n9931), .B(n9917), .Z(n9918) );
  XOR2_X1 U12462 ( .A(n9918), .B(n9919), .Z(n9829) );
  AOI22_X1 U12463 ( .A1(n14972), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n9826) );
  INV_X1 U12464 ( .A(n14995), .ZN(n14897) );
  XNOR2_X1 U12465 ( .A(n9931), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n9817) );
  NAND2_X1 U12466 ( .A1(n9815), .A2(n9814), .ZN(n9816) );
  OAI21_X1 U12467 ( .B1(n9817), .B2(n9816), .A(n9930), .ZN(n9818) );
  NAND2_X1 U12468 ( .A1(n14897), .A2(n9818), .ZN(n9825) );
  XNOR2_X1 U12469 ( .A(n9931), .B(P3_REG1_REG_2__SCAN_IN), .ZN(n9821) );
  NAND2_X1 U12470 ( .A1(n9821), .A2(n9822), .ZN(n9922) );
  OAI21_X1 U12471 ( .B1(n9822), .B2(n9821), .A(n9922), .ZN(n9823) );
  NAND2_X1 U12472 ( .A1(n14896), .A2(n9823), .ZN(n9824) );
  NAND3_X1 U12473 ( .A1(n9826), .A2(n9825), .A3(n9824), .ZN(n9827) );
  AOI21_X1 U12474 ( .B1(n9931), .B2(n14944), .A(n9827), .ZN(n9828) );
  OAI21_X1 U12475 ( .B1(n9829), .B2(n14987), .A(n9828), .ZN(P3_U3184) );
  NAND2_X1 U12476 ( .A1(n12096), .A2(n10266), .ZN(n9830) );
  NAND2_X1 U12477 ( .A1(n9831), .A2(n9830), .ZN(n9836) );
  INV_X1 U12478 ( .A(n9836), .ZN(n10280) );
  INV_X1 U12479 ( .A(n8915), .ZN(n13383) );
  INV_X1 U12480 ( .A(n13426), .ZN(n13464) );
  INV_X1 U12481 ( .A(n13427), .ZN(n13462) );
  OAI22_X1 U12482 ( .A1(n6617), .A2(n13464), .B1(n10133), .B2(n13462), .ZN(
        n9835) );
  NAND2_X1 U12483 ( .A1(n6638), .A2(n11883), .ZN(n9833) );
  AOI21_X1 U12484 ( .B1(n9833), .B2(n9832), .A(n13459), .ZN(n9834) );
  AOI211_X1 U12485 ( .C1(n13383), .C2(n9836), .A(n9835), .B(n9834), .ZN(n10273) );
  OAI211_X1 U12486 ( .C1(n11880), .C2(n6635), .A(n8927), .B(n10285), .ZN(
        n10276) );
  OAI211_X1 U12487 ( .C1(n10280), .C2(n14876), .A(n10273), .B(n10276), .ZN(
        n10049) );
  INV_X1 U12488 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9837) );
  OAI22_X1 U12489 ( .A1(n13640), .A2(n6635), .B1(n14880), .B2(n9837), .ZN(
        n9838) );
  AOI21_X1 U12490 ( .B1(n10049), .B2(n14880), .A(n9838), .ZN(n9839) );
  INV_X1 U12491 ( .A(n9839), .ZN(P2_U3433) );
  INV_X1 U12492 ( .A(n11173), .ZN(n9845) );
  NAND2_X1 U12493 ( .A1(n9841), .A2(n9840), .ZN(n9842) );
  NAND2_X1 U12494 ( .A1(n9842), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9843) );
  XNOR2_X1 U12495 ( .A(n9843), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11174) );
  INV_X1 U12496 ( .A(n11174), .ZN(n14669) );
  OAI222_X1 U12497 ( .A1(n14276), .A2(n9844), .B1(n14270), .B2(n9845), .C1(
        P1_U3086), .C2(n14669), .ZN(P1_U3340) );
  INV_X1 U12498 ( .A(n14821), .ZN(n10419) );
  OAI222_X1 U12499 ( .A1(n13671), .A2(n9846), .B1(n13666), .B2(n9845), .C1(
        P2_U3088), .C2(n10419), .ZN(P2_U3312) );
  OR2_X1 U12500 ( .A1(n13917), .A2(n9847), .ZN(n9851) );
  INV_X1 U12501 ( .A(n9848), .ZN(n9849) );
  OR2_X1 U12502 ( .A1(n9852), .A2(n6978), .ZN(n14106) );
  NAND2_X1 U12503 ( .A1(n9853), .A2(n14106), .ZN(n14009) );
  NAND2_X1 U12504 ( .A1(n9872), .A2(n11399), .ZN(n9854) );
  INV_X1 U12505 ( .A(n9857), .ZN(n9858) );
  OR2_X1 U12506 ( .A1(n11655), .A2(n7532), .ZN(n9860) );
  OAI211_X1 U12507 ( .C1(n11545), .C2(n13833), .A(n9861), .B(n9860), .ZN(
        n14615) );
  NAND2_X1 U12508 ( .A1(n10172), .A2(n14615), .ZN(n11395) );
  INV_X1 U12509 ( .A(n10172), .ZN(n13811) );
  INV_X2 U12510 ( .A(n14615), .ZN(n10171) );
  INV_X1 U12511 ( .A(n11404), .ZN(n11676) );
  NAND2_X1 U12512 ( .A1(n10142), .A2(n11676), .ZN(n10141) );
  NAND2_X1 U12513 ( .A1(n10172), .A2(n10171), .ZN(n9862) );
  NAND2_X1 U12514 ( .A1(n11614), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9868) );
  NAND2_X1 U12515 ( .A1(n11599), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9867) );
  INV_X1 U12516 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9863) );
  NAND2_X1 U12517 ( .A1(n10145), .A2(n9863), .ZN(n9864) );
  NAND2_X1 U12518 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9878) );
  AND2_X1 U12519 ( .A1(n9864), .A2(n9878), .ZN(n9889) );
  NAND2_X1 U12520 ( .A1(n10112), .A2(n9889), .ZN(n9866) );
  NAND2_X1 U12521 ( .A1(n9734), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9865) );
  AOI22_X1 U12522 ( .A1(n11502), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n11501), 
        .B2(n14658), .ZN(n9871) );
  NAND2_X1 U12523 ( .A1(n9869), .A2(n11641), .ZN(n9870) );
  XNOR2_X1 U12524 ( .A(n6446), .B(n11411), .ZN(n11678) );
  XNOR2_X1 U12525 ( .A(n9893), .B(n11678), .ZN(n14717) );
  NAND2_X1 U12526 ( .A1(n9872), .A2(n7375), .ZN(n9873) );
  INV_X1 U12527 ( .A(n11395), .ZN(n9875) );
  XNOR2_X1 U12528 ( .A(n9911), .B(n11678), .ZN(n9876) );
  NOR2_X1 U12529 ( .A1(n9876), .A2(n14574), .ZN(n14721) );
  OR2_X1 U12530 ( .A1(n10172), .A2(n14209), .ZN(n9885) );
  NAND2_X1 U12531 ( .A1(n9899), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9883) );
  NAND2_X1 U12532 ( .A1(n9733), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9882) );
  AND2_X1 U12533 ( .A1(n9878), .A2(n9877), .ZN(n9879) );
  NOR2_X1 U12534 ( .A1(n9900), .A2(n9879), .ZN(n10379) );
  NAND2_X1 U12535 ( .A1(n10112), .A2(n10379), .ZN(n9881) );
  NAND2_X1 U12536 ( .A1(n9734), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9880) );
  NAND4_X1 U12537 ( .A1(n9883), .A2(n9882), .A3(n9881), .A4(n9880), .ZN(n13810) );
  NAND2_X1 U12538 ( .A1(n13810), .A2(n14745), .ZN(n9884) );
  NAND2_X1 U12539 ( .A1(n9885), .A2(n9884), .ZN(n14718) );
  NOR2_X1 U12540 ( .A1(n14721), .A2(n14718), .ZN(n9886) );
  MUX2_X1 U12541 ( .A(n9887), .B(n9886), .S(n14437), .Z(n9892) );
  INV_X1 U12542 ( .A(n9898), .ZN(n9888) );
  AOI211_X1 U12543 ( .C1(n11411), .C2(n10143), .A(n14572), .B(n9888), .ZN(
        n14719) );
  NAND2_X1 U12544 ( .A1(n14437), .A2(n14022), .ZN(n14066) );
  INV_X1 U12545 ( .A(n14019), .ZN(n14426) );
  NAND2_X1 U12546 ( .A1(n14437), .A2(n14426), .ZN(n14096) );
  INV_X1 U12547 ( .A(n9889), .ZN(n10184) );
  OAI22_X1 U12548 ( .A1(n14096), .A2(n11409), .B1(n10184), .B2(n14706), .ZN(
        n9890) );
  AOI21_X1 U12549 ( .B1(n14719), .B2(n14690), .A(n9890), .ZN(n9891) );
  OAI211_X1 U12550 ( .C1(n14700), .C2(n14717), .A(n9892), .B(n9891), .ZN(
        P1_U3289) );
  NAND2_X1 U12551 ( .A1(n9894), .A2(n11641), .ZN(n9897) );
  AOI22_X1 U12552 ( .A1(n11502), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11501), 
        .B2(n9895), .ZN(n9896) );
  NAND2_X1 U12553 ( .A1(n9897), .A2(n9896), .ZN(n11417) );
  XNOR2_X1 U12554 ( .A(n11417), .B(n13810), .ZN(n11679) );
  XNOR2_X1 U12555 ( .A(n10102), .B(n11679), .ZN(n10014) );
  AOI211_X1 U12556 ( .C1(n11417), .C2(n9898), .A(n14572), .B(n10123), .ZN(
        n10010) );
  INV_X1 U12557 ( .A(n11417), .ZN(n10376) );
  OR2_X1 U12558 ( .A1(n11410), .A2(n14209), .ZN(n9907) );
  NAND2_X1 U12559 ( .A1(n11614), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9905) );
  NAND2_X1 U12560 ( .A1(n11599), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9904) );
  NAND2_X1 U12561 ( .A1(n9900), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10114) );
  OR2_X1 U12562 ( .A1(n9900), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9901) );
  AND2_X1 U12563 ( .A1(n10114), .A2(n9901), .ZN(n10651) );
  NAND2_X1 U12564 ( .A1(n11646), .A2(n10651), .ZN(n9903) );
  NAND2_X1 U12565 ( .A1(n9734), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9902) );
  NAND4_X1 U12566 ( .A1(n9905), .A2(n9904), .A3(n9903), .A4(n9902), .ZN(n13809) );
  NAND2_X1 U12567 ( .A1(n13809), .A2(n14745), .ZN(n9906) );
  AND2_X1 U12568 ( .A1(n9907), .A2(n9906), .ZN(n10375) );
  MUX2_X1 U12569 ( .A(n9329), .B(n10375), .S(n14437), .Z(n9909) );
  INV_X1 U12570 ( .A(n14706), .ZN(n14682) );
  NAND2_X1 U12571 ( .A1(n14682), .A2(n10379), .ZN(n9908) );
  OAI211_X1 U12572 ( .C1(n10376), .C2(n14096), .A(n9909), .B(n9908), .ZN(n9910) );
  AOI21_X1 U12573 ( .B1(n10010), .B2(n14690), .A(n9910), .ZN(n9915) );
  NAND2_X1 U12574 ( .A1(n11410), .A2(n11411), .ZN(n9912) );
  NAND2_X1 U12575 ( .A1(n9913), .A2(n9912), .ZN(n10108) );
  XNOR2_X1 U12576 ( .A(n10108), .B(n11679), .ZN(n10012) );
  NAND2_X1 U12577 ( .A1(n10012), .A2(n14434), .ZN(n9914) );
  OAI211_X1 U12578 ( .C1(n10014), .C2(n14700), .A(n9915), .B(n9914), .ZN(
        P1_U3288) );
  MUX2_X1 U12579 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12602), .Z(n10190) );
  XOR2_X1 U12580 ( .A(n9941), .B(n10190), .Z(n10191) );
  INV_X1 U12581 ( .A(n9931), .ZN(n9916) );
  MUX2_X1 U12582 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12602), .Z(n9920) );
  XNOR2_X1 U12583 ( .A(n9920), .B(n11325), .ZN(n14904) );
  INV_X1 U12584 ( .A(n9920), .ZN(n9921) );
  AOI22_X1 U12585 ( .A1(n14905), .A2(n14904), .B1(n11325), .B2(n9921), .ZN(
        n10192) );
  XOR2_X1 U12586 ( .A(n10191), .B(n10192), .Z(n9943) );
  OAI21_X1 U12587 ( .B1(n9931), .B2(n9923), .A(n9922), .ZN(n9924) );
  NAND2_X1 U12588 ( .A1(n9924), .A2(n14906), .ZN(n9928) );
  INV_X1 U12589 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15055) );
  OAI21_X1 U12590 ( .B1(n9924), .B2(n14906), .A(n9928), .ZN(n14910) );
  INV_X1 U12591 ( .A(n14909), .ZN(n9926) );
  INV_X1 U12592 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n9925) );
  XNOR2_X1 U12593 ( .A(n9941), .B(n9925), .ZN(n9927) );
  AOI21_X1 U12594 ( .B1(n9928), .B2(n9926), .A(n9927), .ZN(n10201) );
  AND3_X1 U12595 ( .A1(n9928), .A2(n9927), .A3(n9926), .ZN(n9929) );
  NOR2_X1 U12596 ( .A1(n10201), .A2(n9929), .ZN(n9939) );
  XNOR2_X1 U12597 ( .A(n10202), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n9933) );
  AOI21_X1 U12598 ( .B1(n9934), .B2(n9932), .A(n9933), .ZN(n10197) );
  AND3_X1 U12599 ( .A1(n9934), .A2(n9933), .A3(n9932), .ZN(n9935) );
  OAI21_X1 U12600 ( .B1(n10197), .B2(n9935), .A(n14897), .ZN(n9938) );
  NOR2_X1 U12601 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9936), .ZN(n10446) );
  AOI21_X1 U12602 ( .B1(n14972), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10446), .ZN(
        n9937) );
  OAI211_X1 U12603 ( .C1(n9939), .C2(n14989), .A(n9938), .B(n9937), .ZN(n9940)
         );
  AOI21_X1 U12604 ( .B1(n9941), .B2(n14944), .A(n9940), .ZN(n9942) );
  OAI21_X1 U12605 ( .B1(n9943), .B2(n14987), .A(n9942), .ZN(P3_U3186) );
  INV_X1 U12606 ( .A(n11032), .ZN(n9950) );
  NAND2_X1 U12607 ( .A1(n9945), .A2(n9944), .ZN(n9946) );
  NAND2_X1 U12608 ( .A1(n9946), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9947) );
  XNOR2_X1 U12609 ( .A(n9947), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11033) );
  INV_X1 U12610 ( .A(n11033), .ZN(n10798) );
  OAI222_X1 U12611 ( .A1(n14276), .A2(n9948), .B1(n14270), .B2(n9950), .C1(
        n10798), .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U12612 ( .A(n10402), .ZN(n10416) );
  OAI222_X1 U12613 ( .A1(P2_U3088), .A2(n10416), .B1(n13666), .B2(n9950), .C1(
        n9949), .C2(n13671), .ZN(P2_U3313) );
  NAND2_X1 U12614 ( .A1(n14805), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9952) );
  OAI21_X1 U12615 ( .B1(n9954), .B2(P2_REG2_REG_12__SCAN_IN), .A(n9951), .ZN(
        n14808) );
  MUX2_X1 U12616 ( .A(n11151), .B(P2_REG2_REG_13__SCAN_IN), .S(n14805), .Z(
        n14807) );
  NAND2_X1 U12617 ( .A1(n9952), .A2(n14809), .ZN(n10401) );
  XNOR2_X1 U12618 ( .A(n10401), .B(n10402), .ZN(n10403) );
  XOR2_X1 U12619 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n10403), .Z(n9960) );
  NAND2_X1 U12620 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n11092)
         );
  OAI21_X1 U12621 ( .B1(n9954), .B2(P2_REG1_REG_12__SCAN_IN), .A(n9953), .ZN(
        n14813) );
  XNOR2_X1 U12622 ( .A(n14805), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n14814) );
  NOR2_X1 U12623 ( .A1(n14813), .A2(n14814), .ZN(n14811) );
  AOI21_X1 U12624 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n14805), .A(n14811), 
        .ZN(n10418) );
  XNOR2_X1 U12625 ( .A(n10402), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n10417) );
  XOR2_X1 U12626 ( .A(n10418), .B(n10417), .Z(n9955) );
  NAND2_X1 U12627 ( .A1(n14827), .A2(n9955), .ZN(n9956) );
  NAND2_X1 U12628 ( .A1(n11092), .A2(n9956), .ZN(n9957) );
  AOI21_X1 U12629 ( .B1(n14820), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n9957), .ZN(
        n9959) );
  NAND2_X1 U12630 ( .A1(n14822), .A2(n10402), .ZN(n9958) );
  OAI211_X1 U12631 ( .C1(n9960), .C2(n14806), .A(n9959), .B(n9958), .ZN(
        P2_U3228) );
  NAND2_X1 U12632 ( .A1(n13116), .A2(n13427), .ZN(n13093) );
  NOR2_X1 U12633 ( .A1(n9961), .A2(P2_U3088), .ZN(n10134) );
  INV_X1 U12634 ( .A(n10134), .ZN(n9962) );
  AOI22_X1 U12635 ( .A1(n9962), .A2(P2_REG3_REG_0__SCAN_IN), .B1(n14860), .B2(
        n13120), .ZN(n9966) );
  OAI21_X1 U12636 ( .B1(n6617), .B2(n8927), .A(n11880), .ZN(n9963) );
  NAND3_X1 U12637 ( .A1(n13098), .A2(n9964), .A3(n9963), .ZN(n9965) );
  OAI211_X1 U12638 ( .C1(n10293), .C2(n13093), .A(n9966), .B(n9965), .ZN(
        P2_U3204) );
  INV_X1 U12639 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n14579) );
  MUX2_X1 U12640 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n14579), .S(n11027), .Z(
        n9996) );
  AOI21_X1 U12641 ( .B1(n9661), .B2(n9969), .A(n9967), .ZN(n9998) );
  XOR2_X1 U12642 ( .A(n9996), .B(n9998), .Z(n9978) );
  NOR2_X1 U12643 ( .A1(n14670), .A2(n11027), .ZN(n9976) );
  NAND2_X1 U12644 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14516)
         );
  AOI21_X1 U12645 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(n9973) );
  INV_X1 U12646 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9971) );
  MUX2_X1 U12647 ( .A(n9971), .B(P1_REG2_REG_13__SCAN_IN), .S(n11027), .Z(
        n9972) );
  NAND2_X1 U12648 ( .A1(n9973), .A2(n9972), .ZN(n10002) );
  OAI211_X1 U12649 ( .C1(n9973), .C2(n9972), .A(n10002), .B(n14643), .ZN(n9974) );
  NAND2_X1 U12650 ( .A1(n14516), .A2(n9974), .ZN(n9975) );
  AOI211_X1 U12651 ( .C1(n14633), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n9976), .B(
        n9975), .ZN(n9977) );
  OAI21_X1 U12652 ( .B1(n9978), .B2(n14668), .A(n9977), .ZN(P1_U3256) );
  INV_X1 U12653 ( .A(n12330), .ZN(n9981) );
  NAND3_X1 U12654 ( .A1(n9981), .A2(n9979), .A3(n9980), .ZN(n9982) );
  OAI211_X1 U12655 ( .C1(n9984), .C2(n10248), .A(n9983), .B(n9982), .ZN(n9988)
         );
  INV_X1 U12656 ( .A(n12261), .ZN(n14888) );
  AOI22_X1 U12657 ( .A1(n14888), .A2(n12499), .B1(n12264), .B2(n8666), .ZN(
        n9985) );
  OAI21_X1 U12658 ( .B1(n14891), .B2(n10245), .A(n9985), .ZN(n9987) );
  NOR2_X1 U12659 ( .A1(n12243), .A2(P3_U3151), .ZN(n14895) );
  NOR2_X1 U12660 ( .A1(n14895), .A2(n10246), .ZN(n9986) );
  AOI211_X1 U12661 ( .C1(n9988), .C2(n12216), .A(n9987), .B(n9986), .ZN(n9989)
         );
  INV_X1 U12662 ( .A(n9989), .ZN(P3_U3162) );
  INV_X1 U12663 ( .A(n10628), .ZN(n10624) );
  INV_X1 U12664 ( .A(n11273), .ZN(n9994) );
  OAI222_X1 U12665 ( .A1(P2_U3088), .A2(n10624), .B1(n13666), .B2(n9994), .C1(
        n9990), .C2(n13671), .ZN(P2_U3311) );
  NAND2_X1 U12666 ( .A1(n9991), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9992) );
  MUX2_X1 U12667 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9992), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n9993) );
  INV_X1 U12668 ( .A(n9186), .ZN(n10073) );
  AND2_X1 U12669 ( .A1(n9993), .A2(n10073), .ZN(n11274) );
  INV_X1 U12670 ( .A(n11274), .ZN(n10806) );
  OAI222_X1 U12671 ( .A1(n14276), .A2(n9995), .B1(n14270), .B2(n9994), .C1(
        n10806), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U12672 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14568) );
  AOI22_X1 U12673 ( .A1(n11033), .A2(n14568), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n10798), .ZN(n10001) );
  INV_X1 U12674 ( .A(n9996), .ZN(n9997) );
  NAND2_X1 U12675 ( .A1(n9998), .A2(n9997), .ZN(n9999) );
  OAI21_X1 U12676 ( .B1(n11027), .B2(n14579), .A(n9999), .ZN(n10000) );
  NOR2_X1 U12677 ( .A1(n10001), .A2(n10000), .ZN(n10797) );
  AOI21_X1 U12678 ( .B1(n10001), .B2(n10000), .A(n10797), .ZN(n10009) );
  INV_X1 U12679 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n15216) );
  AOI22_X1 U12680 ( .A1(n11033), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n15216), 
        .B2(n10798), .ZN(n10004) );
  OAI21_X1 U12681 ( .B1(n11027), .B2(n9971), .A(n10002), .ZN(n10003) );
  NAND2_X1 U12682 ( .A1(n10004), .A2(n10003), .ZN(n10790) );
  OAI211_X1 U12683 ( .C1(n10004), .C2(n10003), .A(n14643), .B(n10790), .ZN(
        n10008) );
  NAND2_X1 U12684 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14508)
         );
  NAND2_X1 U12685 ( .A1(n14633), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n10005) );
  OAI211_X1 U12686 ( .C1(n14670), .C2(n10798), .A(n14508), .B(n10005), .ZN(
        n10006) );
  INV_X1 U12687 ( .A(n10006), .ZN(n10007) );
  OAI211_X1 U12688 ( .C1(n10009), .C2(n14668), .A(n10008), .B(n10007), .ZN(
        P1_U3257) );
  INV_X1 U12689 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10016) );
  OAI21_X1 U12690 ( .B1(n10376), .B2(n14748), .A(n10375), .ZN(n10011) );
  AOI211_X1 U12691 ( .C1(n10012), .C2(n14763), .A(n10011), .B(n10010), .ZN(
        n10013) );
  OAI21_X1 U12692 ( .B1(n14755), .B2(n10014), .A(n10013), .ZN(n14231) );
  NAND2_X1 U12693 ( .A1(n14231), .A2(n6444), .ZN(n10015) );
  OAI21_X1 U12694 ( .B1(n6444), .B2(n10016), .A(n10015), .ZN(P1_U3474) );
  INV_X1 U12695 ( .A(n14876), .ZN(n14869) );
  OAI21_X1 U12696 ( .B1(n10018), .B2(n12098), .A(n10017), .ZN(n15076) );
  AOI211_X1 U12697 ( .C1(n15068), .C2(n10286), .A(n13262), .B(n10592), .ZN(
        n15067) );
  INV_X1 U12698 ( .A(n15076), .ZN(n10025) );
  OAI21_X1 U12699 ( .B1(n10021), .B2(n10020), .A(n10019), .ZN(n10023) );
  OAI22_X1 U12700 ( .A1(n10133), .A2(n13464), .B1(n10432), .B2(n13462), .ZN(
        n10022) );
  AOI21_X1 U12701 ( .B1(n10023), .B2(n13421), .A(n10022), .ZN(n10024) );
  OAI21_X1 U12702 ( .B1(n10025), .B2(n8915), .A(n10024), .ZN(n15074) );
  AOI211_X1 U12703 ( .C1(n14869), .C2(n15076), .A(n15067), .B(n15074), .ZN(
        n10031) );
  INV_X1 U12704 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10026) );
  OAI22_X1 U12705 ( .A1(n13640), .A2(n10027), .B1(n14880), .B2(n10026), .ZN(
        n10028) );
  INV_X1 U12706 ( .A(n10028), .ZN(n10029) );
  OAI21_X1 U12707 ( .B1(n10031), .B2(n14879), .A(n10029), .ZN(P2_U3439) );
  AOI22_X1 U12708 ( .A1(n13596), .A2(n15068), .B1(n14883), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n10030) );
  OAI21_X1 U12709 ( .B1(n10031), .B2(n14883), .A(n10030), .ZN(P2_U3502) );
  OAI222_X1 U12710 ( .A1(n12997), .A2(n10034), .B1(n12995), .B2(n10033), .C1(
        P3_U3151), .C2(n10032), .ZN(P3_U3275) );
  AOI22_X1 U12711 ( .A1(n13118), .A2(n15070), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_STATE_REG_SCAN_IN), .ZN(n10036) );
  NAND2_X1 U12712 ( .A1(n13116), .A2(n13426), .ZN(n13072) );
  OAI22_X1 U12713 ( .A1(n10133), .A2(n13072), .B1(n13093), .B2(n10432), .ZN(
        n10035) );
  AOI211_X1 U12714 ( .C1(n15068), .C2(n13120), .A(n10036), .B(n10035), .ZN(
        n10041) );
  OAI211_X1 U12715 ( .C1(n10039), .C2(n10038), .A(n10037), .B(n13098), .ZN(
        n10040) );
  NAND2_X1 U12716 ( .A1(n10041), .A2(n10040), .ZN(P2_U3190) );
  INV_X1 U12717 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10045) );
  NAND2_X1 U12718 ( .A1(n8666), .A2(n14892), .ZN(n12325) );
  INV_X1 U12719 ( .A(n12325), .ZN(n10043) );
  NOR2_X1 U12720 ( .A1(n12330), .A2(n10043), .ZN(n14887) );
  NOR3_X1 U12721 ( .A1(n14887), .A2(n15007), .A3(n12460), .ZN(n10044) );
  AOI21_X1 U12722 ( .B1(n12841), .B2(n10042), .A(n10044), .ZN(n10060) );
  MUX2_X1 U12723 ( .A(n10045), .B(n10060), .S(n15052), .Z(n10046) );
  OAI21_X1 U12724 ( .B1(n14892), .B2(n12979), .A(n10046), .ZN(P3_U3390) );
  MUX2_X1 U12725 ( .A(n8186), .B(n10060), .S(n15066), .Z(n10047) );
  OAI21_X1 U12726 ( .B1(n14892), .B2(n12928), .A(n10047), .ZN(P3_U3459) );
  OAI22_X1 U12727 ( .A1(n8170), .A2(n6635), .B1(n14885), .B2(n9424), .ZN(
        n10048) );
  AOI21_X1 U12728 ( .B1(n14885), .B2(n10049), .A(n10048), .ZN(n10050) );
  INV_X1 U12729 ( .A(n10050), .ZN(P2_U3500) );
  INV_X1 U12730 ( .A(n10051), .ZN(n10052) );
  NOR2_X1 U12731 ( .A1(n10055), .A2(n10052), .ZN(n10054) );
  MUX2_X1 U12732 ( .A(n10055), .B(n10054), .S(n10053), .Z(n10056) );
  NAND2_X1 U12733 ( .A1(n10057), .A2(n10056), .ZN(n10059) );
  NAND2_X1 U12734 ( .A1(n12475), .A2(n15007), .ZN(n10058) );
  OR2_X2 U12735 ( .A1(n10059), .A2(n10058), .ZN(n12866) );
  INV_X1 U12736 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10061) );
  MUX2_X1 U12737 ( .A(n10061), .B(n10060), .S(n12863), .Z(n10063) );
  NAND2_X1 U12738 ( .A1(n12828), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10062) );
  OAI211_X1 U12739 ( .C1(n14892), .C2(n12866), .A(n10063), .B(n10062), .ZN(
        P3_U3233) );
  INV_X1 U12740 ( .A(n10064), .ZN(n10065) );
  AOI21_X1 U12741 ( .B1(n10067), .B2(n10066), .A(n10065), .ZN(n10072) );
  OAI21_X1 U12742 ( .B1(n13093), .B2(n10586), .A(n10068), .ZN(n10070) );
  OAI22_X1 U12743 ( .A1(n13072), .A2(n10587), .B1(n13118), .B2(n10595), .ZN(
        n10069) );
  AOI211_X1 U12744 ( .C1(n14872), .C2(n13120), .A(n10070), .B(n10069), .ZN(
        n10071) );
  OAI21_X1 U12745 ( .B1(n10072), .B2(n13122), .A(n10071), .ZN(P2_U3202) );
  INV_X1 U12746 ( .A(n11297), .ZN(n10076) );
  NAND2_X1 U12747 ( .A1(n10073), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10074) );
  XNOR2_X1 U12748 ( .A(n10074), .B(P1_IR_REG_17__SCAN_IN), .ZN(n11298) );
  INV_X1 U12749 ( .A(n11298), .ZN(n11137) );
  OAI222_X1 U12750 ( .A1(n14276), .A2(n10075), .B1(n14270), .B2(n10076), .C1(
        n11137), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U12751 ( .A(n10631), .ZN(n11198) );
  OAI222_X1 U12752 ( .A1(n13671), .A2(n10077), .B1(n13666), .B2(n10076), .C1(
        n11198), .C2(P2_U3088), .ZN(P2_U3310) );
  OAI21_X1 U12753 ( .B1(n10080), .B2(n10078), .A(n10079), .ZN(n10081) );
  NAND2_X1 U12754 ( .A1(n10081), .A2(n12216), .ZN(n10085) );
  INV_X1 U12755 ( .A(n12264), .ZN(n12227) );
  OAI22_X1 U12756 ( .A1(n8783), .A2(n12227), .B1(n10082), .B2(n12261), .ZN(
        n10083) );
  AOI21_X1 U12757 ( .B1(n12268), .B2(n8230), .A(n10083), .ZN(n10084) );
  OAI211_X1 U12758 ( .C1(n8215), .C2(n14895), .A(n10085), .B(n10084), .ZN(
        P3_U3177) );
  OAI21_X1 U12759 ( .B1(n10088), .B2(n10087), .A(n10086), .ZN(n10089) );
  NAND2_X1 U12760 ( .A1(n10089), .A2(n13098), .ZN(n10094) );
  INV_X1 U12761 ( .A(n13093), .ZN(n11095) );
  INV_X1 U12762 ( .A(n10090), .ZN(n10092) );
  OAI22_X1 U12763 ( .A1(n13072), .A2(n10432), .B1(n13118), .B2(n10602), .ZN(
        n10091) );
  AOI211_X1 U12764 ( .C1(n11095), .C2(n13142), .A(n10092), .B(n10091), .ZN(
        n10093) );
  OAI211_X1 U12765 ( .C1(n6912), .C2(n13077), .A(n10094), .B(n10093), .ZN(
        P2_U3199) );
  OAI21_X1 U12766 ( .B1(n10097), .B2(n10096), .A(n10095), .ZN(n10100) );
  OAI22_X1 U12767 ( .A1(n10293), .A2(n13072), .B1(n13093), .B2(n10587), .ZN(
        n10099) );
  OAI22_X1 U12768 ( .A1(n13077), .A2(n14865), .B1(n10134), .B2(n10288), .ZN(
        n10098) );
  AOI211_X1 U12769 ( .C1(n13098), .C2(n10100), .A(n10099), .B(n10098), .ZN(
        n10101) );
  INV_X1 U12770 ( .A(n10101), .ZN(P2_U3209) );
  INV_X1 U12771 ( .A(n13810), .ZN(n10109) );
  NAND2_X1 U12772 ( .A1(n10376), .A2(n10109), .ZN(n10103) );
  NAND2_X1 U12773 ( .A1(n10104), .A2(n11641), .ZN(n10107) );
  AOI22_X1 U12774 ( .A1(n11502), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11501), 
        .B2(n10105), .ZN(n10106) );
  NAND2_X1 U12775 ( .A1(n10107), .A2(n10106), .ZN(n14727) );
  XNOR2_X1 U12776 ( .A(n14727), .B(n13809), .ZN(n11680) );
  XNOR2_X1 U12777 ( .A(n10322), .B(n11680), .ZN(n14729) );
  NAND2_X1 U12778 ( .A1(n10108), .A2(n11679), .ZN(n10111) );
  NAND2_X1 U12779 ( .A1(n10109), .A2(n11417), .ZN(n10110) );
  INV_X1 U12780 ( .A(n11680), .ZN(n10321) );
  XNOR2_X1 U12781 ( .A(n10333), .B(n10321), .ZN(n10120) );
  NAND2_X1 U12782 ( .A1(n11614), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10119) );
  NAND2_X1 U12783 ( .A1(n11599), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10118) );
  INV_X1 U12784 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10113) );
  NAND2_X1 U12785 ( .A1(n10114), .A2(n10113), .ZN(n10115) );
  AND2_X1 U12786 ( .A1(n10315), .A2(n10115), .ZN(n14681) );
  NAND2_X1 U12787 ( .A1(n11646), .A2(n14681), .ZN(n10117) );
  NAND2_X1 U12788 ( .A1(n9734), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10116) );
  NAND4_X1 U12789 ( .A1(n10119), .A2(n10118), .A3(n10117), .A4(n10116), .ZN(
        n14744) );
  AOI22_X1 U12790 ( .A1(n14745), .A2(n14744), .B1(n13810), .B2(n14766), .ZN(
        n10648) );
  OAI21_X1 U12791 ( .B1(n10120), .B2(n14574), .A(n10648), .ZN(n14725) );
  INV_X1 U12792 ( .A(n14725), .ZN(n10121) );
  MUX2_X1 U12793 ( .A(n10122), .B(n10121), .S(n14437), .Z(n10128) );
  INV_X1 U12794 ( .A(n10123), .ZN(n10124) );
  INV_X1 U12795 ( .A(n14727), .ZN(n10654) );
  AOI211_X1 U12796 ( .C1(n14727), .C2(n10124), .A(n14572), .B(n14688), .ZN(
        n14726) );
  INV_X1 U12797 ( .A(n10651), .ZN(n10125) );
  OAI22_X1 U12798 ( .A1(n14096), .A2(n10654), .B1(n10125), .B2(n14706), .ZN(
        n10126) );
  AOI21_X1 U12799 ( .B1(n14726), .B2(n14690), .A(n10126), .ZN(n10127) );
  OAI211_X1 U12800 ( .C1(n14700), .C2(n14729), .A(n10128), .B(n10127), .ZN(
        P1_U3287) );
  INV_X1 U12801 ( .A(n10129), .ZN(n10130) );
  AOI21_X1 U12802 ( .B1(n10132), .B2(n10131), .A(n10130), .ZN(n10139) );
  INV_X1 U12803 ( .A(n13072), .ZN(n13090) );
  NOR2_X1 U12804 ( .A1(n13093), .A2(n10133), .ZN(n10137) );
  OAI22_X1 U12805 ( .A1(n13077), .A2(n6635), .B1(n10134), .B2(n10275), .ZN(
        n10136) );
  AOI211_X1 U12806 ( .C1(n13090), .C2(n11881), .A(n10137), .B(n10136), .ZN(
        n10138) );
  OAI21_X1 U12807 ( .B1(n10139), .B2(n13122), .A(n10138), .ZN(P2_U3194) );
  INV_X1 U12808 ( .A(n14434), .ZN(n14701) );
  XNOR2_X1 U12809 ( .A(n10140), .B(n11404), .ZN(n14715) );
  INV_X1 U12810 ( .A(n14715), .ZN(n10152) );
  OAI21_X1 U12811 ( .B1(n10142), .B2(n11676), .A(n10141), .ZN(n14709) );
  OAI211_X1 U12812 ( .C1(n10144), .C2(n10171), .A(n14686), .B(n10143), .ZN(
        n14711) );
  AOI22_X1 U12813 ( .A1(n14683), .A2(n14615), .B1(n14682), .B2(n10145), .ZN(
        n10149) );
  OR2_X1 U12814 ( .A1(n11410), .A2(n14420), .ZN(n10147) );
  NAND2_X1 U12815 ( .A1(n13812), .A2(n14766), .ZN(n10146) );
  NAND2_X1 U12816 ( .A1(n10147), .A2(n10146), .ZN(n14624) );
  INV_X1 U12817 ( .A(n14624), .ZN(n14712) );
  MUX2_X1 U12818 ( .A(n9316), .B(n14712), .S(n14437), .Z(n10148) );
  OAI211_X1 U12819 ( .C1(n14711), .C2(n14066), .A(n10149), .B(n10148), .ZN(
        n10150) );
  AOI21_X1 U12820 ( .B1(n14544), .B2(n14709), .A(n10150), .ZN(n10151) );
  OAI21_X1 U12821 ( .B1(n14701), .B2(n10152), .A(n10151), .ZN(P1_U3290) );
  INV_X2 U12822 ( .A(n14437), .ZN(n14704) );
  INV_X1 U12823 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10153) );
  OAI22_X1 U12824 ( .A1(n14437), .A2(n10154), .B1(n10153), .B2(n14706), .ZN(
        n10156) );
  NOR2_X1 U12825 ( .A1(n14096), .A2(n11399), .ZN(n10155) );
  AOI211_X1 U12826 ( .C1(n10157), .C2(n14690), .A(n10156), .B(n10155), .ZN(
        n10160) );
  NAND2_X1 U12827 ( .A1(n14544), .A2(n10158), .ZN(n10159) );
  OAI211_X1 U12828 ( .C1(n14704), .C2(n10161), .A(n10160), .B(n10159), .ZN(
        P1_U3291) );
  OAI222_X1 U12829 ( .A1(n12997), .A2(n10162), .B1(n12995), .B2(n15192), .C1(
        P3_U3151), .C2(n12329), .ZN(P3_U3274) );
  OAI22_X1 U12830 ( .A1(n10172), .A2(n11867), .B1(n10171), .B2(n10169), .ZN(
        n10170) );
  XNOR2_X1 U12831 ( .A(n10170), .B(n11217), .ZN(n10174) );
  OAI22_X1 U12832 ( .A1(n10172), .A2(n9799), .B1(n10171), .B2(n11867), .ZN(
        n10173) );
  XNOR2_X1 U12833 ( .A(n10174), .B(n10173), .ZN(n14622) );
  OAI22_X1 U12834 ( .A1(n11410), .A2(n9799), .B1(n11409), .B2(n11867), .ZN(
        n10368) );
  OAI22_X1 U12835 ( .A1(n11410), .A2(n11867), .B1(n11409), .B2(n10169), .ZN(
        n10175) );
  XNOR2_X1 U12836 ( .A(n10175), .B(n11861), .ZN(n10176) );
  NAND2_X1 U12837 ( .A1(n10177), .A2(n10176), .ZN(n10371) );
  OAI211_X1 U12838 ( .C1(n10177), .C2(n10176), .A(n10371), .B(n14527), .ZN(
        n10187) );
  NOR2_X1 U12839 ( .A1(n14748), .A2(n11409), .ZN(n14720) );
  INV_X1 U12840 ( .A(n10178), .ZN(n10179) );
  NAND2_X1 U12841 ( .A1(n10180), .A2(n10179), .ZN(n10181) );
  NAND2_X1 U12842 ( .A1(n10181), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10182) );
  NAND2_X1 U12843 ( .A1(n14625), .A2(n14718), .ZN(n10183) );
  NAND2_X1 U12844 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14637) );
  OAI211_X1 U12845 ( .C1(n14628), .C2(n10184), .A(n10183), .B(n14637), .ZN(
        n10185) );
  AOI21_X1 U12846 ( .B1(n14618), .B2(n14720), .A(n10185), .ZN(n10186) );
  NAND2_X1 U12847 ( .A1(n10187), .A2(n10186), .ZN(P1_U3230) );
  INV_X1 U12848 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10189) );
  MUX2_X1 U12849 ( .A(n10189), .B(n10188), .S(n12602), .Z(n10527) );
  XNOR2_X1 U12850 ( .A(n10527), .B(n10525), .ZN(n10196) );
  MUX2_X1 U12851 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12602), .Z(n10193) );
  OR2_X1 U12852 ( .A1(n10193), .A2(n14922), .ZN(n10194) );
  XNOR2_X1 U12853 ( .A(n10193), .B(n10203), .ZN(n14920) );
  NAND2_X1 U12854 ( .A1(n14921), .A2(n14920), .ZN(n14919) );
  NAND2_X1 U12855 ( .A1(n10194), .A2(n14919), .ZN(n10195) );
  OAI21_X1 U12856 ( .B1(n10196), .B2(n10195), .A(n10528), .ZN(n10215) );
  NOR2_X1 U12857 ( .A1(n14979), .A2(n10525), .ZN(n10214) );
  INV_X1 U12858 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n14924) );
  NOR2_X1 U12859 ( .A1(n14924), .A2(n14925), .ZN(n14923) );
  NAND2_X1 U12860 ( .A1(n10525), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10514) );
  OAI21_X1 U12861 ( .B1(n10525), .B2(P3_REG2_REG_6__SCAN_IN), .A(n10514), .ZN(
        n10199) );
  AOI21_X1 U12862 ( .B1(n6780), .B2(n10199), .A(n10516), .ZN(n10212) );
  INV_X1 U12863 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10200) );
  NOR2_X1 U12864 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10200), .ZN(n10670) );
  AOI21_X1 U12865 ( .B1(n14972), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n10670), .ZN(
        n10211) );
  AOI21_X1 U12866 ( .B1(P3_REG1_REG_4__SCAN_IN), .B2(n10202), .A(n10201), .ZN(
        n10204) );
  NAND2_X1 U12867 ( .A1(n10525), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10535) );
  OAI21_X1 U12868 ( .B1(n10525), .B2(P3_REG1_REG_6__SCAN_IN), .A(n10535), .ZN(
        n10207) );
  INV_X1 U12869 ( .A(n10207), .ZN(n10206) );
  NAND2_X1 U12870 ( .A1(n10207), .A2(n6580), .ZN(n10208) );
  NAND2_X1 U12871 ( .A1(n10536), .A2(n10208), .ZN(n10209) );
  NAND2_X1 U12872 ( .A1(n14896), .A2(n10209), .ZN(n10210) );
  OAI211_X1 U12873 ( .C1(n10212), .C2(n14995), .A(n10211), .B(n10210), .ZN(
        n10213) );
  AOI211_X1 U12874 ( .C1(n14945), .C2(n10215), .A(n10214), .B(n10213), .ZN(
        n10216) );
  INV_X1 U12875 ( .A(n10216), .ZN(P3_U3188) );
  OAI211_X1 U12876 ( .C1(n10219), .C2(n10218), .A(n10217), .B(n13098), .ZN(
        n10225) );
  NAND2_X1 U12877 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n13147) );
  NAND2_X1 U12878 ( .A1(n13142), .A2(n13426), .ZN(n10221) );
  NAND2_X1 U12879 ( .A1(n13140), .A2(n13427), .ZN(n10220) );
  NAND2_X1 U12880 ( .A1(n10221), .A2(n10220), .ZN(n10458) );
  NAND2_X1 U12881 ( .A1(n13116), .A2(n10458), .ZN(n10222) );
  OAI211_X1 U12882 ( .C1(n13118), .C2(n14835), .A(n13147), .B(n10222), .ZN(
        n10223) );
  AOI21_X1 U12883 ( .B1(n11918), .B2(n13120), .A(n10223), .ZN(n10224) );
  NAND2_X1 U12884 ( .A1(n10225), .A2(n10224), .ZN(P2_U3185) );
  NAND2_X1 U12885 ( .A1(n12500), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n10226) );
  OAI21_X1 U12886 ( .B1(n10227), .B2(n12500), .A(n10226), .ZN(P3_U3519) );
  INV_X1 U12887 ( .A(n10228), .ZN(n10230) );
  OAI22_X1 U12888 ( .A1(n12484), .A2(P3_U3151), .B1(SI_22_), .B2(n12995), .ZN(
        n10229) );
  AOI21_X1 U12889 ( .B1(n10230), .B2(n14397), .A(n10229), .ZN(P3_U3273) );
  OAI21_X1 U12890 ( .B1(n10232), .B2(n10234), .A(n10231), .ZN(n10608) );
  INV_X1 U12891 ( .A(n10456), .ZN(n10233) );
  AOI211_X1 U12892 ( .C1(n13104), .C2(n10429), .A(n13465), .B(n10233), .ZN(
        n10613) );
  XNOR2_X1 U12893 ( .A(n10235), .B(n10234), .ZN(n10238) );
  NAND2_X1 U12894 ( .A1(n13143), .A2(n13426), .ZN(n10237) );
  NAND2_X1 U12895 ( .A1(n13141), .A2(n13427), .ZN(n10236) );
  AND2_X1 U12896 ( .A1(n10237), .A2(n10236), .ZN(n13102) );
  OAI21_X1 U12897 ( .B1(n10238), .B2(n13459), .A(n13102), .ZN(n10609) );
  AOI211_X1 U12898 ( .C1(n13584), .C2(n10608), .A(n10613), .B(n10609), .ZN(
        n10243) );
  INV_X1 U12899 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10239) );
  OAI22_X1 U12900 ( .A1(n13640), .A2(n6910), .B1(n14880), .B2(n10239), .ZN(
        n10240) );
  INV_X1 U12901 ( .A(n10240), .ZN(n10241) );
  OAI21_X1 U12902 ( .B1(n10243), .B2(n14879), .A(n10241), .ZN(P2_U3448) );
  AOI22_X1 U12903 ( .A1(n13596), .A2(n13104), .B1(n14883), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n10242) );
  OAI21_X1 U12904 ( .B1(n10243), .B2(n14883), .A(n10242), .ZN(P2_U3505) );
  XNOR2_X1 U12905 ( .A(n9979), .B(n12330), .ZN(n14997) );
  NOR2_X1 U12906 ( .A1(n12475), .A2(n12329), .ZN(n11116) );
  INV_X1 U12907 ( .A(n11116), .ZN(n10244) );
  NOR2_X1 U12908 ( .A1(n10245), .A2(n15044), .ZN(n14999) );
  NOR2_X1 U12909 ( .A1(n12864), .A2(n10246), .ZN(n10252) );
  INV_X1 U12910 ( .A(n11117), .ZN(n10953) );
  AOI22_X1 U12911 ( .A1(n12844), .A2(n8666), .B1(n12499), .B2(n12841), .ZN(
        n10251) );
  OAI21_X1 U12912 ( .B1(n9979), .B2(n10248), .A(n10247), .ZN(n10249) );
  NAND2_X1 U12913 ( .A1(n10249), .A2(n12837), .ZN(n10250) );
  OAI211_X1 U12914 ( .C1(n14997), .C2(n10953), .A(n10251), .B(n10250), .ZN(
        n14998) );
  AOI211_X1 U12915 ( .C1(n14999), .C2(n12475), .A(n10252), .B(n14998), .ZN(
        n10253) );
  MUX2_X1 U12916 ( .A(n10254), .B(n10253), .S(n12863), .Z(n10255) );
  OAI21_X1 U12917 ( .B1(n14997), .B2(n10957), .A(n10255), .ZN(P3_U3232) );
  NAND2_X1 U12918 ( .A1(n12500), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10256) );
  OAI21_X1 U12919 ( .B1(n12289), .B2(n12500), .A(n10256), .ZN(P3_U3521) );
  NAND2_X1 U12920 ( .A1(n10257), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10258) );
  XNOR2_X1 U12921 ( .A(n10258), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13851) );
  INV_X1 U12922 ( .A(n13851), .ZN(n11145) );
  OAI222_X1 U12923 ( .A1(P1_U3086), .A2(n11145), .B1(n14270), .B2(n11496), 
        .C1(n10259), .C2(n14276), .ZN(P1_U3337) );
  INV_X1 U12924 ( .A(n13199), .ZN(n10260) );
  OAI222_X1 U12925 ( .A1(P2_U3088), .A2(n10260), .B1(n13666), .B2(n11496), 
        .C1(n15202), .C2(n13671), .ZN(P2_U3309) );
  INV_X1 U12926 ( .A(n10261), .ZN(n10262) );
  NAND2_X1 U12927 ( .A1(n10263), .A2(n10262), .ZN(n10264) );
  NAND2_X2 U12928 ( .A1(n10264), .A2(n13487), .ZN(n13490) );
  AOI21_X1 U12929 ( .B1(n14833), .B2(n8927), .A(n13493), .ZN(n10272) );
  NOR2_X2 U12930 ( .A1(n12085), .A2(n13312), .ZN(n15077) );
  NAND2_X1 U12931 ( .A1(n13490), .A2(n15077), .ZN(n13393) );
  NOR2_X1 U12932 ( .A1(n11881), .A2(n14860), .ZN(n10265) );
  OR2_X1 U12933 ( .A1(n10266), .A2(n10265), .ZN(n14855) );
  NOR2_X1 U12934 ( .A1(n13393), .A2(n14855), .ZN(n10270) );
  AOI21_X1 U12935 ( .B1(n13459), .B2(n8915), .A(n14855), .ZN(n10267) );
  AOI21_X1 U12936 ( .B1(n13427), .B2(n8917), .A(n10267), .ZN(n14856) );
  OAI22_X1 U12937 ( .A1(n15079), .A2(n14856), .B1(n10268), .B2(n13487), .ZN(
        n10269) );
  AOI211_X1 U12938 ( .C1(n15079), .C2(P2_REG2_REG_0__SCAN_IN), .A(n10270), .B(
        n10269), .ZN(n10271) );
  OAI21_X1 U12939 ( .B1(n10272), .B2(n11880), .A(n10271), .ZN(P2_U3265) );
  MUX2_X1 U12940 ( .A(n10274), .B(n10273), .S(n13490), .Z(n10279) );
  OAI22_X1 U12941 ( .A1(n13410), .A2(n10276), .B1(n10275), .B2(n13487), .ZN(
        n10277) );
  AOI21_X1 U12942 ( .B1(n13493), .B2(n11885), .A(n10277), .ZN(n10278) );
  OAI211_X1 U12943 ( .C1(n10280), .C2(n13393), .A(n10279), .B(n10278), .ZN(
        P2_U3264) );
  INV_X1 U12944 ( .A(n10281), .ZN(n10282) );
  NAND2_X1 U12945 ( .A1(n10282), .A2(n12095), .ZN(n10284) );
  AND2_X1 U12946 ( .A1(n10283), .A2(n10284), .ZN(n14862) );
  NOR2_X1 U12947 ( .A1(n13490), .A2(n15082), .ZN(n10290) );
  AOI21_X1 U12948 ( .B1(n10285), .B2(n11890), .A(n13465), .ZN(n10287) );
  NAND2_X1 U12949 ( .A1(n10287), .A2(n10286), .ZN(n14863) );
  OAI22_X1 U12950 ( .A1(n13410), .A2(n14863), .B1(n10288), .B2(n13487), .ZN(
        n10289) );
  AOI211_X1 U12951 ( .C1(n13493), .C2(n11890), .A(n10290), .B(n10289), .ZN(
        n10298) );
  OAI21_X1 U12952 ( .B1(n10292), .B2(n12095), .A(n10291), .ZN(n10295) );
  OAI22_X1 U12953 ( .A1(n10293), .A2(n13464), .B1(n10587), .B2(n13462), .ZN(
        n10294) );
  AOI21_X1 U12954 ( .B1(n10295), .B2(n13421), .A(n10294), .ZN(n10296) );
  OAI21_X1 U12955 ( .B1(n14862), .B2(n8915), .A(n10296), .ZN(n14866) );
  NAND2_X1 U12956 ( .A1(n14866), .A2(n13490), .ZN(n10297) );
  OAI211_X1 U12957 ( .C1(n14862), .C2(n13393), .A(n10298), .B(n10297), .ZN(
        P2_U3263) );
  XNOR2_X1 U12958 ( .A(n10299), .B(n10300), .ZN(n15001) );
  NOR2_X1 U12959 ( .A1(n8789), .A2(n15044), .ZN(n15003) );
  NOR2_X1 U12960 ( .A1(n12864), .A2(n8215), .ZN(n10306) );
  AOI22_X1 U12961 ( .A1(n12841), .A2(n12498), .B1(n10042), .B2(n12844), .ZN(
        n10305) );
  OAI21_X1 U12962 ( .B1(n10302), .B2(n10299), .A(n10301), .ZN(n10303) );
  NAND2_X1 U12963 ( .A1(n10303), .A2(n12837), .ZN(n10304) );
  OAI211_X1 U12964 ( .C1(n15001), .C2(n10953), .A(n10305), .B(n10304), .ZN(
        n15002) );
  AOI211_X1 U12965 ( .C1(n15003), .C2(n12475), .A(n10306), .B(n15002), .ZN(
        n10307) );
  MUX2_X1 U12966 ( .A(n10308), .B(n10307), .S(n12863), .Z(n10309) );
  OAI21_X1 U12967 ( .B1(n15001), .B2(n10957), .A(n10309), .ZN(P3_U3231) );
  NAND2_X1 U12968 ( .A1(n10310), .A2(n11641), .ZN(n10313) );
  AOI22_X1 U12969 ( .A1(n11502), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11501), 
        .B2(n10311), .ZN(n10312) );
  NAND2_X1 U12970 ( .A1(n11599), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10320) );
  NAND2_X1 U12971 ( .A1(n11614), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10319) );
  INV_X1 U12972 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10314) );
  NAND2_X1 U12973 ( .A1(n10315), .A2(n10314), .ZN(n10316) );
  NAND2_X1 U12974 ( .A1(n10340), .A2(n10316), .ZN(n10925) );
  INV_X1 U12975 ( .A(n10925), .ZN(n10346) );
  NAND2_X1 U12976 ( .A1(n11646), .A2(n10346), .ZN(n10318) );
  NAND2_X1 U12977 ( .A1(n9734), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10317) );
  NAND4_X1 U12978 ( .A1(n10320), .A2(n10319), .A3(n10318), .A4(n10317), .ZN(
        n13808) );
  NAND2_X1 U12979 ( .A1(n10322), .A2(n10321), .ZN(n10324) );
  OR2_X1 U12980 ( .A1(n14727), .A2(n13809), .ZN(n10323) );
  NAND2_X1 U12981 ( .A1(n10324), .A2(n10323), .ZN(n14676) );
  NAND2_X1 U12982 ( .A1(n10325), .A2(n11641), .ZN(n10328) );
  AOI22_X1 U12983 ( .A1(n11502), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11501), 
        .B2(n10326), .ZN(n10327) );
  NAND2_X1 U12984 ( .A1(n10328), .A2(n10327), .ZN(n14684) );
  XNOR2_X1 U12985 ( .A(n14684), .B(n10926), .ZN(n14677) );
  NAND2_X1 U12986 ( .A1(n14676), .A2(n14677), .ZN(n10330) );
  OR2_X1 U12987 ( .A1(n14684), .A2(n14744), .ZN(n10329) );
  XOR2_X1 U12988 ( .A(n10471), .B(n11682), .Z(n14742) );
  INV_X1 U12989 ( .A(n13809), .ZN(n10331) );
  AND2_X1 U12990 ( .A1(n14727), .A2(n10331), .ZN(n10332) );
  NOR2_X1 U12991 ( .A1(n14684), .A2(n10926), .ZN(n10335) );
  NAND2_X1 U12992 ( .A1(n14684), .A2(n10926), .ZN(n10334) );
  OAI211_X1 U12993 ( .C1(n10337), .C2(n10336), .A(n14763), .B(n10479), .ZN(
        n14750) );
  MUX2_X1 U12994 ( .A(n14750), .B(n10338), .S(n14704), .Z(n10351) );
  INV_X1 U12995 ( .A(n14684), .ZN(n14687) );
  AOI21_X1 U12996 ( .B1(n14685), .B2(n11435), .A(n14572), .ZN(n10339) );
  AND2_X1 U12997 ( .A1(n10339), .A2(n10490), .ZN(n14743) );
  NAND2_X1 U12998 ( .A1(n14437), .A2(n14766), .ZN(n14064) );
  AND2_X1 U12999 ( .A1(n14437), .A2(n14745), .ZN(n14061) );
  NAND2_X1 U13000 ( .A1(n11614), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10345) );
  NAND2_X1 U13001 ( .A1(n11599), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10344) );
  AND2_X1 U13002 ( .A1(n10340), .A2(n11218), .ZN(n10341) );
  NOR2_X1 U13003 ( .A1(n10748), .A2(n10341), .ZN(n11221) );
  NAND2_X1 U13004 ( .A1(n11646), .A2(n11221), .ZN(n10343) );
  NAND2_X1 U13005 ( .A1(n11657), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10342) );
  NAND4_X1 U13006 ( .A1(n10345), .A2(n10344), .A3(n10343), .A4(n10342), .ZN(
        n14765) );
  AOI22_X1 U13007 ( .A1(n14061), .A2(n14765), .B1(n10346), .B2(n14682), .ZN(
        n10348) );
  NAND2_X1 U13008 ( .A1(n14683), .A2(n11435), .ZN(n10347) );
  OAI211_X1 U13009 ( .C1(n10926), .C2(n14064), .A(n10348), .B(n10347), .ZN(
        n10349) );
  AOI21_X1 U13010 ( .B1(n14743), .B2(n14690), .A(n10349), .ZN(n10350) );
  OAI211_X1 U13011 ( .C1(n14700), .C2(n14742), .A(n10351), .B(n10350), .ZN(
        P1_U3285) );
  NAND2_X1 U13012 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_U3151), .ZN(n14916) );
  OAI21_X1 U13013 ( .B1(n12350), .B2(n12261), .A(n14916), .ZN(n10352) );
  AOI21_X1 U13014 ( .B1(n12264), .B2(n12499), .A(n10352), .ZN(n10353) );
  OAI21_X1 U13015 ( .B1(n14891), .B2(n10354), .A(n10353), .ZN(n10359) );
  AOI211_X1 U13016 ( .C1(n10357), .C2(n10356), .A(n14886), .B(n10355), .ZN(
        n10358) );
  AOI211_X1 U13017 ( .C1(n10564), .C2(n12243), .A(n10359), .B(n10358), .ZN(
        n10360) );
  INV_X1 U13018 ( .A(n10360), .ZN(P3_U3158) );
  NAND2_X1 U13019 ( .A1(n11417), .A2(n11858), .ZN(n10363) );
  NAND2_X1 U13020 ( .A1(n13810), .A2(n11801), .ZN(n10362) );
  NAND2_X1 U13021 ( .A1(n10363), .A2(n10362), .ZN(n10364) );
  XNOR2_X1 U13022 ( .A(n10364), .B(n11861), .ZN(n10639) );
  NAND2_X1 U13023 ( .A1(n11863), .A2(n13810), .ZN(n10366) );
  NAND2_X1 U13024 ( .A1(n11417), .A2(n11801), .ZN(n10365) );
  NAND2_X1 U13025 ( .A1(n10366), .A2(n10365), .ZN(n10638) );
  XNOR2_X1 U13026 ( .A(n10639), .B(n10638), .ZN(n10373) );
  INV_X1 U13027 ( .A(n10367), .ZN(n10369) );
  NAND2_X1 U13028 ( .A1(n10369), .A2(n10368), .ZN(n10370) );
  AOI21_X1 U13029 ( .B1(n10373), .B2(n10372), .A(n10640), .ZN(n10381) );
  OAI21_X1 U13030 ( .B1(n10375), .B2(n13733), .A(n10374), .ZN(n10378) );
  NOR2_X1 U13031 ( .A1(n14500), .A2(n10376), .ZN(n10377) );
  AOI211_X1 U13032 ( .C1(n10379), .C2(n13798), .A(n10378), .B(n10377), .ZN(
        n10380) );
  OAI21_X1 U13033 ( .B1(n10381), .B2(n14620), .A(n10380), .ZN(P1_U3227) );
  NAND2_X1 U13034 ( .A1(n10383), .A2(n10382), .ZN(n10385) );
  XOR2_X1 U13035 ( .A(n10385), .B(n10384), .Z(n10392) );
  NAND2_X1 U13036 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n13160) );
  NAND2_X1 U13037 ( .A1(n13141), .A2(n13426), .ZN(n10387) );
  NAND2_X1 U13038 ( .A1(n13139), .A2(n13427), .ZN(n10386) );
  AND2_X1 U13039 ( .A1(n10387), .A2(n10386), .ZN(n10507) );
  INV_X1 U13040 ( .A(n10507), .ZN(n10388) );
  NAND2_X1 U13041 ( .A1(n13116), .A2(n10388), .ZN(n10389) );
  OAI211_X1 U13042 ( .C1(n13118), .C2(n10571), .A(n13160), .B(n10389), .ZN(
        n10390) );
  AOI21_X1 U13043 ( .B1(n11923), .B2(n13120), .A(n10390), .ZN(n10391) );
  OAI21_X1 U13044 ( .B1(n10392), .B2(n13122), .A(n10391), .ZN(P2_U3193) );
  INV_X1 U13045 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n15124) );
  INV_X1 U13046 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n10396) );
  NAND2_X1 U13047 ( .A1(n10393), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n10395) );
  INV_X1 U13048 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12929) );
  OR2_X1 U13049 ( .A1(n8238), .A2(n12929), .ZN(n10394) );
  OAI211_X1 U13050 ( .C1(n10396), .C2(n6448), .A(n10395), .B(n10394), .ZN(
        n10397) );
  INV_X1 U13051 ( .A(n10397), .ZN(n10398) );
  NAND2_X1 U13052 ( .A1(n12624), .A2(P3_U3897), .ZN(n10400) );
  OAI21_X1 U13053 ( .B1(P3_U3897), .B2(n15124), .A(n10400), .ZN(P3_U3522) );
  NAND2_X1 U13054 ( .A1(n10402), .A2(n10401), .ZN(n10406) );
  INV_X1 U13055 ( .A(n10403), .ZN(n10404) );
  NAND2_X1 U13056 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n10404), .ZN(n10405) );
  NAND2_X1 U13057 ( .A1(n10406), .A2(n10405), .ZN(n10407) );
  NAND2_X1 U13058 ( .A1(n14821), .A2(n10407), .ZN(n10408) );
  XNOR2_X1 U13059 ( .A(n10419), .B(n10407), .ZN(n14825) );
  NAND2_X1 U13060 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14825), .ZN(n14823) );
  NAND2_X1 U13061 ( .A1(n10408), .A2(n14823), .ZN(n10413) );
  INV_X1 U13062 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10410) );
  NAND2_X1 U13063 ( .A1(n10628), .A2(n10410), .ZN(n10409) );
  OAI21_X1 U13064 ( .B1(n10628), .B2(n10410), .A(n10409), .ZN(n10412) );
  NAND2_X1 U13065 ( .A1(n10624), .A2(n10410), .ZN(n10411) );
  OAI211_X1 U13066 ( .C1(n10410), .C2(n10624), .A(n10413), .B(n10411), .ZN(
        n10623) );
  OAI211_X1 U13067 ( .C1(n10413), .C2(n10412), .A(n10623), .B(n14824), .ZN(
        n10426) );
  NAND2_X1 U13068 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13041)
         );
  INV_X1 U13069 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10414) );
  XNOR2_X1 U13070 ( .A(n10628), .B(n10414), .ZN(n10629) );
  OAI22_X1 U13071 ( .A1(n10418), .A2(n10417), .B1(n10416), .B2(n10415), .ZN(
        n10420) );
  NAND2_X1 U13072 ( .A1(n14821), .A2(n10420), .ZN(n10421) );
  XNOR2_X1 U13073 ( .A(n10420), .B(n10419), .ZN(n14828) );
  NAND2_X1 U13074 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14828), .ZN(n14826) );
  NAND2_X1 U13075 ( .A1(n10421), .A2(n14826), .ZN(n10630) );
  XOR2_X1 U13076 ( .A(n10629), .B(n10630), .Z(n10422) );
  NAND2_X1 U13077 ( .A1(n14827), .A2(n10422), .ZN(n10423) );
  NAND2_X1 U13078 ( .A1(n13041), .A2(n10423), .ZN(n10424) );
  AOI21_X1 U13079 ( .B1(n14820), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n10424), 
        .ZN(n10425) );
  OAI211_X1 U13080 ( .C1(n10637), .C2(n10624), .A(n10426), .B(n10425), .ZN(
        P2_U3230) );
  OAI21_X1 U13081 ( .B1(n10428), .B2(n10433), .A(n10427), .ZN(n10599) );
  AOI21_X1 U13082 ( .B1(n10593), .B2(n11908), .A(n13465), .ZN(n10430) );
  AND2_X1 U13083 ( .A1(n10430), .A2(n10429), .ZN(n10604) );
  OAI22_X1 U13084 ( .A1(n10432), .A2(n13464), .B1(n10431), .B2(n13462), .ZN(
        n10437) );
  XNOR2_X1 U13085 ( .A(n10434), .B(n10433), .ZN(n10435) );
  NOR2_X1 U13086 ( .A1(n10435), .A2(n13459), .ZN(n10436) );
  AOI211_X1 U13087 ( .C1(n13383), .C2(n10599), .A(n10437), .B(n10436), .ZN(
        n10600) );
  INV_X1 U13088 ( .A(n10600), .ZN(n10438) );
  AOI211_X1 U13089 ( .C1(n14869), .C2(n10599), .A(n10604), .B(n10438), .ZN(
        n10442) );
  AOI22_X1 U13090 ( .A1(n13596), .A2(n11908), .B1(n14883), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n10439) );
  OAI21_X1 U13091 ( .B1(n10442), .B2(n14883), .A(n10439), .ZN(P2_U3504) );
  OAI22_X1 U13092 ( .A1(n13640), .A2(n6912), .B1(n14880), .B2(n7728), .ZN(
        n10440) );
  INV_X1 U13093 ( .A(n10440), .ZN(n10441) );
  OAI21_X1 U13094 ( .B1(n10442), .B2(n14879), .A(n10441), .ZN(P2_U3445) );
  OAI21_X1 U13095 ( .B1(n10445), .B2(n10444), .A(n10443), .ZN(n10451) );
  INV_X1 U13096 ( .A(n12243), .ZN(n12266) );
  NOR2_X1 U13097 ( .A1(n12266), .A2(n10686), .ZN(n10450) );
  AOI21_X1 U13098 ( .B1(n14888), .B2(n12497), .A(n10446), .ZN(n10448) );
  NAND2_X1 U13099 ( .A1(n12264), .A2(n12498), .ZN(n10447) );
  OAI211_X1 U13100 ( .C1(n14891), .C2(n15012), .A(n10448), .B(n10447), .ZN(
        n10449) );
  AOI211_X1 U13101 ( .C1(n10451), .C2(n12216), .A(n10450), .B(n10449), .ZN(
        n10452) );
  INV_X1 U13102 ( .A(n10452), .ZN(P3_U3170) );
  OAI21_X1 U13103 ( .B1(n10455), .B2(n10454), .A(n10453), .ZN(n14843) );
  AOI211_X1 U13104 ( .C1(n11918), .C2(n10456), .A(n13262), .B(n10502), .ZN(
        n14834) );
  XNOR2_X1 U13105 ( .A(n10457), .B(n12104), .ZN(n10459) );
  AOI21_X1 U13106 ( .B1(n10459), .B2(n13421), .A(n10458), .ZN(n14845) );
  INV_X1 U13107 ( .A(n14845), .ZN(n10460) );
  AOI211_X1 U13108 ( .C1(n13584), .C2(n14843), .A(n14834), .B(n10460), .ZN(
        n10464) );
  INV_X1 U13109 ( .A(n11918), .ZN(n14840) );
  OAI22_X1 U13110 ( .A1(n13640), .A2(n14840), .B1(n14880), .B2(n7756), .ZN(
        n10461) );
  INV_X1 U13111 ( .A(n10461), .ZN(n10462) );
  OAI21_X1 U13112 ( .B1(n10464), .B2(n14879), .A(n10462), .ZN(P2_U3451) );
  AOI22_X1 U13113 ( .A1(n13596), .A2(n11918), .B1(n14883), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n10463) );
  OAI21_X1 U13114 ( .B1(n10464), .B2(n14883), .A(n10463), .ZN(P2_U3506) );
  INV_X1 U13115 ( .A(n11500), .ZN(n10466) );
  OAI222_X1 U13116 ( .A1(n13671), .A2(n10465), .B1(n13666), .B2(n10466), .C1(
        n13312), .C2(P2_U3088), .ZN(P2_U3308) );
  OAI222_X1 U13117 ( .A1(n14276), .A2(n10467), .B1(n14270), .B2(n10466), .C1(
        P1_U3086), .C2(n14022), .ZN(P1_U3336) );
  NAND2_X1 U13118 ( .A1(n10468), .A2(n14397), .ZN(n10469) );
  OAI211_X1 U13119 ( .C1(n10470), .C2(n12995), .A(n10469), .B(n12486), .ZN(
        P3_U3272) );
  NAND2_X1 U13120 ( .A1(n10471), .A2(n11682), .ZN(n10473) );
  OR2_X1 U13121 ( .A1(n11435), .A2(n13808), .ZN(n10472) );
  NAND2_X1 U13122 ( .A1(n10473), .A2(n10472), .ZN(n10736) );
  NAND2_X1 U13123 ( .A1(n10474), .A2(n11641), .ZN(n10477) );
  AOI22_X1 U13124 ( .A1(n11502), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11501), 
        .B2(n10475), .ZN(n10476) );
  XNOR2_X1 U13125 ( .A(n11440), .B(n14765), .ZN(n11685) );
  XNOR2_X1 U13126 ( .A(n10736), .B(n11685), .ZN(n14756) );
  OAI21_X1 U13127 ( .B1(n10480), .B2(n11685), .A(n10762), .ZN(n10481) );
  NAND2_X1 U13128 ( .A1(n10481), .A2(n14763), .ZN(n10489) );
  NAND2_X1 U13129 ( .A1(n13808), .A2(n14766), .ZN(n10488) );
  NAND2_X1 U13130 ( .A1(n11599), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10486) );
  NAND2_X1 U13131 ( .A1(n11614), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10485) );
  INV_X1 U13132 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10482) );
  XNOR2_X1 U13133 ( .A(n10748), .B(n10482), .ZN(n11261) );
  NAND2_X1 U13134 ( .A1(n11646), .A2(n11261), .ZN(n10484) );
  NAND2_X1 U13135 ( .A1(n11657), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10483) );
  NAND4_X1 U13136 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n14520) );
  NAND2_X1 U13137 ( .A1(n14520), .A2(n14745), .ZN(n10487) );
  AND2_X1 U13138 ( .A1(n10488), .A2(n10487), .ZN(n11219) );
  NAND2_X1 U13139 ( .A1(n10489), .A2(n11219), .ZN(n14759) );
  NAND2_X1 U13140 ( .A1(n14759), .A2(n14437), .ZN(n10498) );
  NAND2_X1 U13141 ( .A1(n10490), .A2(n11440), .ZN(n10491) );
  NAND2_X1 U13142 ( .A1(n10491), .A2(n14686), .ZN(n10492) );
  NOR2_X1 U13143 ( .A1(n10855), .A2(n10492), .ZN(n14757) );
  INV_X1 U13144 ( .A(n11221), .ZN(n10495) );
  NAND2_X1 U13145 ( .A1(n11440), .A2(n14683), .ZN(n10494) );
  NAND2_X1 U13146 ( .A1(n14704), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10493) );
  OAI211_X1 U13147 ( .C1(n14706), .C2(n10495), .A(n10494), .B(n10493), .ZN(
        n10496) );
  AOI21_X1 U13148 ( .B1(n14757), .B2(n14690), .A(n10496), .ZN(n10497) );
  OAI211_X1 U13149 ( .C1(n14756), .C2(n14700), .A(n10498), .B(n10497), .ZN(
        P1_U3284) );
  INV_X1 U13150 ( .A(n10499), .ZN(n10500) );
  AOI21_X1 U13151 ( .B1(n12094), .B2(n10501), .A(n10500), .ZN(n10568) );
  INV_X1 U13152 ( .A(n10502), .ZN(n10504) );
  INV_X1 U13153 ( .A(n10779), .ZN(n10503) );
  AOI211_X1 U13154 ( .C1(n11923), .C2(n10504), .A(n13465), .B(n10503), .ZN(
        n10574) );
  OAI211_X1 U13155 ( .C1(n10506), .C2(n12094), .A(n10505), .B(n13421), .ZN(
        n10508) );
  NAND2_X1 U13156 ( .A1(n10508), .A2(n10507), .ZN(n10575) );
  AOI211_X1 U13157 ( .C1(n10568), .C2(n13584), .A(n10574), .B(n10575), .ZN(
        n10513) );
  INV_X1 U13158 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10509) );
  OAI22_X1 U13159 ( .A1(n13640), .A2(n10572), .B1(n14880), .B2(n10509), .ZN(
        n10510) );
  INV_X1 U13160 ( .A(n10510), .ZN(n10511) );
  OAI21_X1 U13161 ( .B1(n10513), .B2(n14879), .A(n10511), .ZN(P2_U3454) );
  AOI22_X1 U13162 ( .A1(n13596), .A2(n11923), .B1(n14883), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n10512) );
  OAI21_X1 U13163 ( .B1(n10513), .B2(n14883), .A(n10512), .ZN(P2_U3507) );
  INV_X1 U13164 ( .A(n10514), .ZN(n10515) );
  NOR2_X1 U13165 ( .A1(n7145), .A2(n10517), .ZN(n10518) );
  NOR2_X1 U13166 ( .A1(n10518), .A2(n14938), .ZN(n10521) );
  NAND2_X1 U13167 ( .A1(n10716), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n10711) );
  OAI21_X1 U13168 ( .B1(n10716), .B2(P3_REG2_REG_8__SCAN_IN), .A(n10711), .ZN(
        n10520) );
  INV_X1 U13169 ( .A(n10712), .ZN(n10519) );
  AOI21_X1 U13170 ( .B1(n10521), .B2(n10520), .A(n10519), .ZN(n10547) );
  INV_X1 U13171 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10523) );
  MUX2_X1 U13172 ( .A(n10523), .B(n10522), .S(n12602), .Z(n10718) );
  XNOR2_X1 U13173 ( .A(n10718), .B(n10716), .ZN(n10532) );
  MUX2_X1 U13174 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12602), .Z(n10524) );
  OR2_X1 U13175 ( .A1(n10524), .A2(n10537), .ZN(n10530) );
  XNOR2_X1 U13176 ( .A(n10524), .B(n7145), .ZN(n14942) );
  INV_X1 U13177 ( .A(n10525), .ZN(n10526) );
  NAND2_X1 U13178 ( .A1(n10527), .A2(n10526), .ZN(n10529) );
  NAND2_X1 U13179 ( .A1(n14942), .A2(n14943), .ZN(n14941) );
  NAND2_X1 U13180 ( .A1(n10530), .A2(n14941), .ZN(n10531) );
  OAI21_X1 U13181 ( .B1(n10532), .B2(n10531), .A(n10719), .ZN(n10545) );
  NOR2_X1 U13182 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10533), .ZN(n10882) );
  AOI21_X1 U13183 ( .B1(n14972), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n10882), .ZN(
        n10534) );
  OAI21_X1 U13184 ( .B1(n14979), .B2(n10716), .A(n10534), .ZN(n10544) );
  NOR2_X1 U13185 ( .A1(n7145), .A2(n10538), .ZN(n10539) );
  NAND2_X1 U13186 ( .A1(n10716), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n10725) );
  OAI21_X1 U13187 ( .B1(n10716), .B2(P3_REG1_REG_8__SCAN_IN), .A(n10725), .ZN(
        n10540) );
  NAND2_X1 U13188 ( .A1(n10541), .A2(n10540), .ZN(n10542) );
  AOI21_X1 U13189 ( .B1(n10726), .B2(n10542), .A(n14989), .ZN(n10543) );
  AOI211_X1 U13190 ( .C1(n14945), .C2(n10545), .A(n10544), .B(n10543), .ZN(
        n10546) );
  OAI21_X1 U13191 ( .B1(n10547), .B2(n14995), .A(n10546), .ZN(P3_U3190) );
  XOR2_X1 U13192 ( .A(n10549), .B(n10548), .Z(n10556) );
  INV_X1 U13193 ( .A(n10550), .ZN(n10661) );
  NAND2_X1 U13194 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(P3_U3151), .ZN(n14933) );
  INV_X1 U13195 ( .A(n14933), .ZN(n10551) );
  AOI21_X1 U13196 ( .B1(n14888), .B2(n12496), .A(n10551), .ZN(n10553) );
  NAND2_X1 U13197 ( .A1(n12264), .A2(n12353), .ZN(n10552) );
  OAI211_X1 U13198 ( .C1(n14891), .C2(n15017), .A(n10553), .B(n10552), .ZN(
        n10554) );
  AOI21_X1 U13199 ( .B1(n10661), .B2(n12243), .A(n10554), .ZN(n10555) );
  OAI21_X1 U13200 ( .B1(n10556), .B2(n14886), .A(n10555), .ZN(P3_U3167) );
  XNOR2_X1 U13201 ( .A(n10557), .B(n12298), .ZN(n15008) );
  INV_X1 U13202 ( .A(n15008), .ZN(n10567) );
  OAI22_X1 U13203 ( .A1(n12350), .A2(n12862), .B1(n8231), .B2(n12860), .ZN(
        n10562) );
  INV_X1 U13204 ( .A(n10558), .ZN(n10559) );
  AOI211_X1 U13205 ( .C1(n12298), .C2(n10560), .A(n12858), .B(n10559), .ZN(
        n10561) );
  AOI211_X1 U13206 ( .C1(n15008), .C2(n11117), .A(n10562), .B(n10561), .ZN(
        n15010) );
  MUX2_X1 U13207 ( .A(n10563), .B(n15010), .S(n12863), .Z(n10566) );
  INV_X1 U13208 ( .A(n12866), .ZN(n12796) );
  AOI22_X1 U13209 ( .A1(n12796), .A2(n15006), .B1(n12828), .B2(n10564), .ZN(
        n10565) );
  OAI211_X1 U13210 ( .C1(n10567), .C2(n10957), .A(n10566), .B(n10565), .ZN(
        P3_U3230) );
  INV_X1 U13211 ( .A(n10568), .ZN(n10580) );
  INV_X1 U13212 ( .A(n15077), .ZN(n10569) );
  NAND2_X1 U13213 ( .A1(n10569), .A2(n8915), .ZN(n10570) );
  OAI22_X1 U13214 ( .A1(n14839), .A2(n10572), .B1(n13487), .B2(n10571), .ZN(
        n10573) );
  AOI21_X1 U13215 ( .B1(n10574), .B2(n14833), .A(n10573), .ZN(n10579) );
  INV_X1 U13216 ( .A(n10575), .ZN(n10577) );
  MUX2_X1 U13217 ( .A(n10577), .B(n10576), .S(n15079), .Z(n10578) );
  OAI211_X1 U13218 ( .C1(n10580), .C2(n13474), .A(n10579), .B(n10578), .ZN(
        P2_U3257) );
  OAI21_X1 U13219 ( .B1(n10582), .B2(n12099), .A(n10581), .ZN(n10583) );
  INV_X1 U13220 ( .A(n10583), .ZN(n14877) );
  OAI21_X1 U13221 ( .B1(n10585), .B2(n11898), .A(n10584), .ZN(n10590) );
  OAI22_X1 U13222 ( .A1(n10587), .A2(n13464), .B1(n10586), .B2(n13462), .ZN(
        n10589) );
  NOR2_X1 U13223 ( .A1(n14877), .A2(n8915), .ZN(n10588) );
  AOI211_X1 U13224 ( .C1(n13421), .C2(n10590), .A(n10589), .B(n10588), .ZN(
        n14875) );
  MUX2_X1 U13225 ( .A(n10591), .B(n14875), .S(n13490), .Z(n10598) );
  INV_X1 U13226 ( .A(n10592), .ZN(n10594) );
  AOI211_X1 U13227 ( .C1(n14872), .C2(n10594), .A(n13465), .B(n6913), .ZN(
        n14871) );
  OAI22_X1 U13228 ( .A1(n14839), .A2(n11902), .B1(n10595), .B2(n13487), .ZN(
        n10596) );
  AOI21_X1 U13229 ( .B1(n14833), .B2(n14871), .A(n10596), .ZN(n10597) );
  OAI211_X1 U13230 ( .C1(n14877), .C2(n13393), .A(n10598), .B(n10597), .ZN(
        P2_U3261) );
  INV_X1 U13231 ( .A(n10599), .ZN(n10607) );
  MUX2_X1 U13232 ( .A(n10601), .B(n10600), .S(n13490), .Z(n10606) );
  OAI22_X1 U13233 ( .A1(n14839), .A2(n6912), .B1(n13487), .B2(n10602), .ZN(
        n10603) );
  AOI21_X1 U13234 ( .B1(n14833), .B2(n10604), .A(n10603), .ZN(n10605) );
  OAI211_X1 U13235 ( .C1(n10607), .C2(n13393), .A(n10606), .B(n10605), .ZN(
        P2_U3260) );
  INV_X1 U13236 ( .A(n10608), .ZN(n10616) );
  INV_X1 U13237 ( .A(n10609), .ZN(n10610) );
  MUX2_X1 U13238 ( .A(n10611), .B(n10610), .S(n13490), .Z(n10615) );
  OAI22_X1 U13239 ( .A1(n14839), .A2(n6910), .B1(n13487), .B2(n13105), .ZN(
        n10612) );
  AOI21_X1 U13240 ( .B1(n10613), .B2(n14833), .A(n10612), .ZN(n10614) );
  OAI211_X1 U13241 ( .C1(n13474), .C2(n10616), .A(n10615), .B(n10614), .ZN(
        P2_U3259) );
  AOI21_X1 U13242 ( .B1(n10618), .B2(n10617), .A(n6577), .ZN(n10622) );
  NOR2_X1 U13243 ( .A1(n13118), .A2(n13488), .ZN(n10620) );
  INV_X1 U13244 ( .A(n13116), .ZN(n13082) );
  AOI22_X1 U13245 ( .A1(n13426), .A2(n13140), .B1(n13138), .B2(n13427), .ZN(
        n10783) );
  NAND2_X1 U13246 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n13192) );
  OAI21_X1 U13247 ( .B1(n13082), .B2(n10783), .A(n13192), .ZN(n10619) );
  AOI211_X1 U13248 ( .C1(n13492), .C2(n13120), .A(n10620), .B(n10619), .ZN(
        n10621) );
  OAI21_X1 U13249 ( .B1(n10622), .B2(n13122), .A(n10621), .ZN(P2_U3203) );
  OAI21_X1 U13250 ( .B1(n10410), .B2(n10624), .A(n10623), .ZN(n10627) );
  NAND2_X1 U13251 ( .A1(n10631), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11203) );
  INV_X1 U13252 ( .A(n11203), .ZN(n10625) );
  AOI21_X1 U13253 ( .B1(n13407), .B2(n11198), .A(n10625), .ZN(n10626) );
  NAND2_X1 U13254 ( .A1(n10626), .A2(n10627), .ZN(n11202) );
  OAI211_X1 U13255 ( .C1(n10627), .C2(n10626), .A(n14824), .B(n11202), .ZN(
        n10636) );
  NAND2_X1 U13256 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13052)
         );
  AOI22_X1 U13257 ( .A1(n10630), .A2(n10629), .B1(n10628), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n11200) );
  XNOR2_X1 U13258 ( .A(n10631), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n11199) );
  XOR2_X1 U13259 ( .A(n11200), .B(n11199), .Z(n10632) );
  NAND2_X1 U13260 ( .A1(n14827), .A2(n10632), .ZN(n10633) );
  NAND2_X1 U13261 ( .A1(n13052), .A2(n10633), .ZN(n10634) );
  AOI21_X1 U13262 ( .B1(n14820), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n10634), 
        .ZN(n10635) );
  OAI211_X1 U13263 ( .C1(n10637), .C2(n11198), .A(n10636), .B(n10635), .ZN(
        P2_U3231) );
  INV_X1 U13264 ( .A(n10638), .ZN(n10642) );
  INV_X1 U13265 ( .A(n10639), .ZN(n10641) );
  NAND2_X1 U13266 ( .A1(n14727), .A2(n11858), .ZN(n10644) );
  NAND2_X1 U13267 ( .A1(n13809), .A2(n11801), .ZN(n10643) );
  NAND2_X1 U13268 ( .A1(n10644), .A2(n10643), .ZN(n10645) );
  XNOR2_X1 U13269 ( .A(n10645), .B(n11217), .ZN(n10695) );
  AOI22_X1 U13270 ( .A1(n14727), .A2(n11801), .B1(n11863), .B2(n13809), .ZN(
        n10696) );
  XNOR2_X1 U13271 ( .A(n10695), .B(n10696), .ZN(n10646) );
  OAI211_X1 U13272 ( .C1(n10647), .C2(n10646), .A(n10698), .B(n14527), .ZN(
        n10653) );
  NOR2_X1 U13273 ( .A1(n13733), .A2(n10648), .ZN(n10649) );
  AOI211_X1 U13274 ( .C1(n10651), .C2(n13798), .A(n10650), .B(n10649), .ZN(
        n10652) );
  OAI211_X1 U13275 ( .C1(n10654), .C2(n14500), .A(n10653), .B(n10652), .ZN(
        P1_U3239) );
  OR2_X1 U13276 ( .A1(n10656), .A2(n12346), .ZN(n10907) );
  INV_X1 U13277 ( .A(n10907), .ZN(n10655) );
  AOI21_X1 U13278 ( .B1(n12346), .B2(n10656), .A(n10655), .ZN(n10660) );
  AOI22_X1 U13279 ( .A1(n12844), .A2(n12353), .B1(n12496), .B2(n12841), .ZN(
        n10659) );
  XNOR2_X1 U13280 ( .A(n10657), .B(n12346), .ZN(n15020) );
  NAND2_X1 U13281 ( .A1(n15020), .A2(n11117), .ZN(n10658) );
  OAI211_X1 U13282 ( .C1(n10660), .C2(n12858), .A(n10659), .B(n10658), .ZN(
        n15018) );
  INV_X1 U13283 ( .A(n15018), .ZN(n10666) );
  AOI22_X1 U13284 ( .A1(n12796), .A2(n10662), .B1(n12828), .B2(n10661), .ZN(
        n10663) );
  OAI21_X1 U13285 ( .B1(n14924), .B2(n12863), .A(n10663), .ZN(n10664) );
  AOI21_X1 U13286 ( .B1(n15020), .B2(n12647), .A(n10664), .ZN(n10665) );
  OAI21_X1 U13287 ( .B1(n10666), .B2(n12833), .A(n10665), .ZN(P3_U3228) );
  OAI211_X1 U13288 ( .C1(n10669), .C2(n10668), .A(n10667), .B(n12216), .ZN(
        n10676) );
  INV_X1 U13289 ( .A(n10670), .ZN(n10672) );
  NAND2_X1 U13290 ( .A1(n12264), .A2(n12497), .ZN(n10671) );
  OAI211_X1 U13291 ( .C1(n10884), .C2(n12261), .A(n10672), .B(n10671), .ZN(
        n10673) );
  AOI21_X1 U13292 ( .B1(n12268), .B2(n10674), .A(n10673), .ZN(n10675) );
  OAI211_X1 U13293 ( .C1(n10904), .C2(n12266), .A(n10676), .B(n10675), .ZN(
        P3_U3179) );
  XNOR2_X1 U13294 ( .A(n10678), .B(n10677), .ZN(n10683) );
  NOR2_X1 U13295 ( .A1(n13118), .A2(n13476), .ZN(n10681) );
  AOI22_X1 U13296 ( .A1(n13427), .A2(n13137), .B1(n13139), .B2(n13426), .ZN(
        n10896) );
  OAI21_X1 U13297 ( .B1(n13082), .B2(n10896), .A(n10679), .ZN(n10680) );
  AOI211_X1 U13298 ( .C1(n13479), .C2(n13120), .A(n10681), .B(n10680), .ZN(
        n10682) );
  OAI21_X1 U13299 ( .B1(n10683), .B2(n13122), .A(n10682), .ZN(P2_U3189) );
  XNOR2_X1 U13300 ( .A(n10685), .B(n10684), .ZN(n15013) );
  INV_X1 U13301 ( .A(n15013), .ZN(n10693) );
  OAI22_X1 U13302 ( .A1(n12866), .A2(n15012), .B1(n10686), .B2(n12864), .ZN(
        n10692) );
  XNOR2_X1 U13303 ( .A(n10687), .B(n12344), .ZN(n10688) );
  NAND2_X1 U13304 ( .A1(n10688), .A2(n12837), .ZN(n10690) );
  AOI22_X1 U13305 ( .A1(n12844), .A2(n12498), .B1(n12497), .B2(n12841), .ZN(
        n10689) );
  OAI211_X1 U13306 ( .C1(n15013), .C2(n10953), .A(n10690), .B(n10689), .ZN(
        n15015) );
  MUX2_X1 U13307 ( .A(n15015), .B(P3_REG2_REG_4__SCAN_IN), .S(n12833), .Z(
        n10691) );
  AOI211_X1 U13308 ( .C1(n10693), .C2(n12647), .A(n10692), .B(n10691), .ZN(
        n10694) );
  INV_X1 U13309 ( .A(n10694), .ZN(P3_U3229) );
  INV_X1 U13310 ( .A(n10695), .ZN(n10697) );
  NAND2_X1 U13311 ( .A1(n10698), .A2(n7443), .ZN(n10702) );
  AND2_X1 U13312 ( .A1(n11863), .A2(n14744), .ZN(n10699) );
  AOI21_X1 U13313 ( .B1(n14684), .B2(n11801), .A(n10699), .ZN(n10919) );
  AOI22_X1 U13314 ( .A1(n14684), .A2(n11858), .B1(n11801), .B2(n14744), .ZN(
        n10700) );
  XNOR2_X1 U13315 ( .A(n10700), .B(n11217), .ZN(n10918) );
  XOR2_X1 U13316 ( .A(n10919), .B(n10918), .Z(n10701) );
  OAI21_X1 U13317 ( .B1(n10702), .B2(n10701), .A(n14527), .ZN(n10710) );
  NAND2_X1 U13318 ( .A1(n13809), .A2(n14766), .ZN(n10704) );
  NAND2_X1 U13319 ( .A1(n13808), .A2(n14745), .ZN(n10703) );
  AND2_X1 U13320 ( .A1(n10704), .A2(n10703), .ZN(n14736) );
  OAI21_X1 U13321 ( .B1(n13733), .B2(n14736), .A(n10705), .ZN(n10708) );
  NAND2_X1 U13322 ( .A1(n14684), .A2(n14767), .ZN(n14735) );
  INV_X1 U13323 ( .A(n14618), .ZN(n10706) );
  NOR2_X1 U13324 ( .A1(n14735), .A2(n10706), .ZN(n10707) );
  AOI211_X1 U13325 ( .C1(n14681), .C2(n13798), .A(n10708), .B(n10707), .ZN(
        n10709) );
  OAI21_X1 U13326 ( .B1(n10710), .B2(n10921), .A(n10709), .ZN(P1_U3213) );
  AOI21_X1 U13327 ( .B1(n8335), .B2(n10713), .A(n10986), .ZN(n10734) );
  MUX2_X1 U13328 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n12602), .Z(n10714) );
  NOR2_X1 U13329 ( .A1(n10714), .A2(n10727), .ZN(n11007) );
  NAND2_X1 U13330 ( .A1(n10714), .A2(n10727), .ZN(n11009) );
  INV_X1 U13331 ( .A(n11009), .ZN(n10715) );
  OR2_X1 U13332 ( .A1(n11007), .A2(n10715), .ZN(n10722) );
  INV_X1 U13333 ( .A(n10716), .ZN(n10717) );
  NAND2_X1 U13334 ( .A1(n10718), .A2(n10717), .ZN(n10720) );
  INV_X1 U13335 ( .A(n11008), .ZN(n10721) );
  XNOR2_X1 U13336 ( .A(n10722), .B(n10721), .ZN(n10732) );
  NOR2_X1 U13337 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10723), .ZN(n11102) );
  AOI21_X1 U13338 ( .B1(n14972), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11102), .ZN(
        n10724) );
  OAI21_X1 U13339 ( .B1(n14979), .B2(n10727), .A(n10724), .ZN(n10731) );
  INV_X1 U13340 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15062) );
  AOI21_X1 U13341 ( .B1(n15062), .B2(n10728), .A(n10995), .ZN(n10729) );
  NOR2_X1 U13342 ( .A1(n10729), .A2(n14989), .ZN(n10730) );
  AOI211_X1 U13343 ( .C1(n14945), .C2(n10732), .A(n10731), .B(n10730), .ZN(
        n10733) );
  OAI21_X1 U13344 ( .B1(n10734), .B2(n14995), .A(n10733), .ZN(P3_U3191) );
  INV_X1 U13345 ( .A(n11685), .ZN(n10735) );
  NAND2_X1 U13346 ( .A1(n10736), .A2(n10735), .ZN(n10738) );
  OR2_X1 U13347 ( .A1(n11440), .A2(n14765), .ZN(n10737) );
  AOI22_X1 U13348 ( .A1(n11501), .A2(n10740), .B1(n11502), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n10741) );
  NAND2_X2 U13349 ( .A1(n10742), .A2(n10741), .ZN(n14768) );
  INV_X1 U13350 ( .A(n14520), .ZN(n10743) );
  NAND2_X1 U13351 ( .A1(n14768), .A2(n10743), .ZN(n10744) );
  XNOR2_X1 U13352 ( .A(n10859), .B(n11684), .ZN(n14773) );
  XNOR2_X1 U13353 ( .A(n10855), .B(n14768), .ZN(n10755) );
  NAND2_X1 U13354 ( .A1(n10748), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10746) );
  INV_X1 U13355 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10745) );
  NAND2_X1 U13356 ( .A1(n10746), .A2(n10745), .ZN(n10749) );
  AND2_X1 U13357 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n10747) );
  NAND2_X1 U13358 ( .A1(n10748), .A2(n10747), .ZN(n10836) );
  NAND2_X1 U13359 ( .A1(n10749), .A2(n10836), .ZN(n14530) );
  INV_X1 U13360 ( .A(n14530), .ZN(n14537) );
  NAND2_X1 U13361 ( .A1(n11646), .A2(n14537), .ZN(n10753) );
  NAND2_X1 U13362 ( .A1(n11599), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10752) );
  NAND2_X1 U13363 ( .A1(n11657), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10751) );
  NAND2_X1 U13364 ( .A1(n9899), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10750) );
  NAND4_X1 U13365 ( .A1(n10753), .A2(n10752), .A3(n10751), .A4(n10750), .ZN(
        n14404) );
  AND2_X1 U13366 ( .A1(n14404), .A2(n14745), .ZN(n10754) );
  AOI21_X1 U13367 ( .B1(n10755), .B2(n14686), .A(n10754), .ZN(n14770) );
  INV_X1 U13368 ( .A(n14064), .ZN(n14094) );
  INV_X1 U13369 ( .A(n11261), .ZN(n10756) );
  OAI22_X1 U13370 ( .A1(n14437), .A2(n10757), .B1(n10756), .B2(n14706), .ZN(
        n10758) );
  AOI21_X1 U13371 ( .B1(n14094), .B2(n14765), .A(n10758), .ZN(n10760) );
  NAND2_X1 U13372 ( .A1(n14768), .A2(n14683), .ZN(n10759) );
  OAI211_X1 U13373 ( .C1(n14770), .C2(n14066), .A(n10760), .B(n10759), .ZN(
        n10766) );
  INV_X1 U13374 ( .A(n14765), .ZN(n11264) );
  NAND2_X1 U13375 ( .A1(n11440), .A2(n11264), .ZN(n10761) );
  INV_X1 U13376 ( .A(n11684), .ZN(n10763) );
  OR2_X1 U13377 ( .A1(n10764), .A2(n10763), .ZN(n14764) );
  AND3_X1 U13378 ( .A1(n14764), .A2(n14434), .A3(n14762), .ZN(n10765) );
  AOI211_X1 U13379 ( .C1(n14544), .C2(n14773), .A(n10766), .B(n10765), .ZN(
        n10767) );
  INV_X1 U13380 ( .A(n10767), .ZN(P1_U3283) );
  XNOR2_X1 U13381 ( .A(n10769), .B(n10768), .ZN(n15028) );
  XNOR2_X1 U13382 ( .A(n10770), .B(n12363), .ZN(n10773) );
  OAI22_X1 U13383 ( .A1(n11104), .A2(n12862), .B1(n10771), .B2(n12860), .ZN(
        n10772) );
  AOI21_X1 U13384 ( .B1(n10773), .B2(n12837), .A(n10772), .ZN(n10774) );
  OAI21_X1 U13385 ( .B1(n10953), .B2(n15028), .A(n10774), .ZN(n15030) );
  NAND2_X1 U13386 ( .A1(n15030), .A2(n12863), .ZN(n10777) );
  OAI22_X1 U13387 ( .A1(n12866), .A2(n15027), .B1(n10815), .B2(n12864), .ZN(
        n10775) );
  AOI21_X1 U13388 ( .B1(n12833), .B2(P3_REG2_REG_7__SCAN_IN), .A(n10775), .ZN(
        n10776) );
  OAI211_X1 U13389 ( .C1(n15028), .C2(n10957), .A(n10777), .B(n10776), .ZN(
        P3_U3226) );
  XNOR2_X1 U13390 ( .A(n10778), .B(n12106), .ZN(n13494) );
  AOI21_X1 U13391 ( .B1(n10779), .B2(n13492), .A(n13465), .ZN(n10780) );
  AND2_X1 U13392 ( .A1(n10780), .A2(n10890), .ZN(n13495) );
  AOI21_X1 U13393 ( .B1(n10782), .B2(n10781), .A(n6576), .ZN(n10784) );
  OAI21_X1 U13394 ( .B1(n10784), .B2(n13459), .A(n10783), .ZN(n13486) );
  AOI211_X1 U13395 ( .C1(n13584), .C2(n13494), .A(n13495), .B(n13486), .ZN(
        n10789) );
  AOI22_X1 U13396 ( .A1(n13596), .A2(n13492), .B1(n14883), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n10785) );
  OAI21_X1 U13397 ( .B1(n10789), .B2(n14883), .A(n10785), .ZN(P2_U3508) );
  INV_X1 U13398 ( .A(n13492), .ZN(n10786) );
  OAI22_X1 U13399 ( .A1(n13640), .A2(n10786), .B1(n14880), .B2(n7788), .ZN(
        n10787) );
  INV_X1 U13400 ( .A(n10787), .ZN(n10788) );
  OAI21_X1 U13401 ( .B1(n10789), .B2(n14879), .A(n10788), .ZN(P2_U3457) );
  OAI21_X1 U13402 ( .B1(n15216), .B2(n10798), .A(n10790), .ZN(n10791) );
  NOR2_X1 U13403 ( .A1(n11174), .A2(n10791), .ZN(n10792) );
  XNOR2_X1 U13404 ( .A(n11174), .B(n10791), .ZN(n14664) );
  NOR2_X1 U13405 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14664), .ZN(n14663) );
  NOR2_X1 U13406 ( .A1(n10792), .A2(n14663), .ZN(n10795) );
  NOR2_X1 U13407 ( .A1(n11274), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n10793) );
  AOI21_X1 U13408 ( .B1(n11274), .B2(P1_REG2_REG_16__SCAN_IN), .A(n10793), 
        .ZN(n10794) );
  NAND2_X1 U13409 ( .A1(n10794), .A2(n10795), .ZN(n10867) );
  OAI211_X1 U13410 ( .C1(n10795), .C2(n10794), .A(n14643), .B(n10867), .ZN(
        n10805) );
  NAND2_X1 U13411 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13731)
         );
  INV_X1 U13412 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10796) );
  XNOR2_X1 U13413 ( .A(n11274), .B(n10796), .ZN(n10872) );
  AOI21_X1 U13414 ( .B1(n10798), .B2(n14568), .A(n10797), .ZN(n10799) );
  NOR2_X1 U13415 ( .A1(n11174), .A2(n10799), .ZN(n10800) );
  XNOR2_X1 U13416 ( .A(n11174), .B(n10799), .ZN(n14662) );
  NOR2_X1 U13417 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14662), .ZN(n14661) );
  NOR2_X1 U13418 ( .A1(n10800), .A2(n14661), .ZN(n10873) );
  XOR2_X1 U13419 ( .A(n10872), .B(n10873), .Z(n10801) );
  NAND2_X1 U13420 ( .A1(n14652), .A2(n10801), .ZN(n10802) );
  NAND2_X1 U13421 ( .A1(n13731), .A2(n10802), .ZN(n10803) );
  AOI21_X1 U13422 ( .B1(n14633), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10803), 
        .ZN(n10804) );
  OAI211_X1 U13423 ( .C1(n14670), .C2(n10806), .A(n10805), .B(n10804), .ZN(
        P1_U3259) );
  OAI211_X1 U13424 ( .C1(n10809), .C2(n10808), .A(n10807), .B(n12216), .ZN(
        n10814) );
  NAND2_X1 U13425 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(P3_U3151), .ZN(n14951) );
  NAND2_X1 U13426 ( .A1(n12264), .A2(n12496), .ZN(n10810) );
  OAI211_X1 U13427 ( .C1(n11104), .C2(n12261), .A(n14951), .B(n10810), .ZN(
        n10811) );
  AOI21_X1 U13428 ( .B1(n12268), .B2(n10812), .A(n10811), .ZN(n10813) );
  OAI211_X1 U13429 ( .C1(n10815), .C2(n12266), .A(n10814), .B(n10813), .ZN(
        P3_U3153) );
  INV_X1 U13430 ( .A(n10816), .ZN(n10817) );
  OAI222_X1 U13431 ( .A1(n10818), .A2(P3_U3151), .B1(n12997), .B2(n10817), 
        .C1(n7609), .C2(n12995), .ZN(P3_U3271) );
  XNOR2_X1 U13432 ( .A(n10819), .B(n10820), .ZN(n10825) );
  NOR2_X1 U13433 ( .A1(n13118), .A2(n10978), .ZN(n10823) );
  AOI22_X1 U13434 ( .A1(n13427), .A2(n13136), .B1(n13138), .B2(n13426), .ZN(
        n10973) );
  OAI21_X1 U13435 ( .B1(n13082), .B2(n10973), .A(n10821), .ZN(n10822) );
  AOI211_X1 U13436 ( .C1(n13600), .C2(n13120), .A(n10823), .B(n10822), .ZN(
        n10824) );
  OAI21_X1 U13437 ( .B1(n10825), .B2(n13122), .A(n10824), .ZN(P2_U3208) );
  NAND2_X1 U13438 ( .A1(n10826), .A2(n11641), .ZN(n10829) );
  AOI22_X1 U13439 ( .A1(n11502), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n10827), 
        .B2(n11501), .ZN(n10828) );
  XNOR2_X1 U13440 ( .A(n14538), .B(n14404), .ZN(n14532) );
  INV_X1 U13441 ( .A(n14404), .ZN(n10854) );
  OR2_X1 U13442 ( .A1(n6612), .A2(n10854), .ZN(n10830) );
  NAND2_X1 U13443 ( .A1(n10831), .A2(n11641), .ZN(n10834) );
  AOI22_X1 U13444 ( .A1(n10832), .A2(n11501), .B1(n11502), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n10833) );
  NAND2_X1 U13445 ( .A1(n11614), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10841) );
  NAND2_X1 U13446 ( .A1(n11599), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10840) );
  NAND2_X1 U13447 ( .A1(n10836), .A2(n10835), .ZN(n10837) );
  AND2_X1 U13448 ( .A1(n10844), .A2(n10837), .ZN(n13713) );
  NAND2_X1 U13449 ( .A1(n11646), .A2(n13713), .ZN(n10839) );
  NAND2_X1 U13450 ( .A1(n11657), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10838) );
  NAND4_X1 U13451 ( .A1(n10841), .A2(n10840), .A3(n10839), .A4(n10838), .ZN(
        n14519) );
  XNOR2_X1 U13452 ( .A(n13712), .B(n14519), .ZN(n11687) );
  NAND2_X1 U13453 ( .A1(n10842), .A2(n11687), .ZN(n11025) );
  OAI211_X1 U13454 ( .C1(n10842), .C2(n11687), .A(n14763), .B(n11025), .ZN(
        n14410) );
  AOI22_X1 U13455 ( .A1(n14704), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n13713), 
        .B2(n14682), .ZN(n10853) );
  NAND2_X1 U13456 ( .A1(n11599), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n10851) );
  NAND2_X1 U13457 ( .A1(n11614), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10850) );
  NAND2_X1 U13458 ( .A1(n11657), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10849) );
  INV_X1 U13459 ( .A(n11036), .ZN(n10846) );
  NAND2_X1 U13460 ( .A1(n10844), .A2(n10843), .ZN(n10845) );
  NAND2_X1 U13461 ( .A1(n10846), .A2(n10845), .ZN(n14518) );
  INV_X1 U13462 ( .A(n14518), .ZN(n10847) );
  NAND2_X1 U13463 ( .A1(n11646), .A2(n10847), .ZN(n10848) );
  NAND4_X1 U13464 ( .A1(n10851), .A2(n10850), .A3(n10849), .A4(n10848), .ZN(
        n14558) );
  NAND2_X1 U13465 ( .A1(n14061), .A2(n14558), .ZN(n10852) );
  OAI211_X1 U13466 ( .C1(n10854), .C2(n14064), .A(n10853), .B(n10852), .ZN(
        n10858) );
  INV_X1 U13467 ( .A(n6612), .ZN(n14582) );
  NAND2_X1 U13468 ( .A1(n14542), .A2(n14582), .ZN(n14541) );
  AOI21_X1 U13469 ( .B1(n14541), .B2(n13712), .A(n14572), .ZN(n10856) );
  NAND2_X1 U13470 ( .A1(n10856), .A2(n14416), .ZN(n14406) );
  NOR2_X1 U13471 ( .A1(n14406), .A2(n14066), .ZN(n10857) );
  AOI211_X1 U13472 ( .C1(n14683), .C2(n13712), .A(n10858), .B(n10857), .ZN(
        n10865) );
  NAND2_X1 U13473 ( .A1(n10859), .A2(n11684), .ZN(n10861) );
  OR2_X1 U13474 ( .A1(n14768), .A2(n14520), .ZN(n10860) );
  NAND2_X1 U13475 ( .A1(n10861), .A2(n10860), .ZN(n14539) );
  INV_X1 U13476 ( .A(n14532), .ZN(n14540) );
  NAND2_X1 U13477 ( .A1(n14539), .A2(n14540), .ZN(n10863) );
  OR2_X1 U13478 ( .A1(n6612), .A2(n14404), .ZN(n10862) );
  NAND2_X1 U13479 ( .A1(n10863), .A2(n10862), .ZN(n11056) );
  XNOR2_X1 U13480 ( .A(n11056), .B(n11687), .ZN(n14411) );
  INV_X1 U13481 ( .A(n14411), .ZN(n14413) );
  NAND2_X1 U13482 ( .A1(n14413), .A2(n14544), .ZN(n10864) );
  OAI211_X1 U13483 ( .C1(n14410), .C2(n14704), .A(n10865), .B(n10864), .ZN(
        P1_U3281) );
  OAI222_X1 U13484 ( .A1(n14276), .A2(n15142), .B1(n14270), .B2(n11514), .C1(
        n11375), .C2(P1_U3086), .ZN(P1_U3335) );
  OAI222_X1 U13485 ( .A1(n13671), .A2(n10866), .B1(P2_U3088), .B2(n12091), 
        .C1(n13666), .C2(n11514), .ZN(P2_U3307) );
  NAND2_X1 U13486 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n11274), .ZN(n10868) );
  NAND2_X1 U13487 ( .A1(n10868), .A2(n10867), .ZN(n10871) );
  INV_X1 U13488 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U13489 ( .A1(n11298), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10869), 
        .B2(n11137), .ZN(n10870) );
  NAND2_X1 U13490 ( .A1(n10870), .A2(n10871), .ZN(n11133) );
  OAI211_X1 U13491 ( .C1(n10871), .C2(n10870), .A(n14643), .B(n11133), .ZN(
        n10878) );
  NAND2_X1 U13492 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13742)
         );
  AOI22_X1 U13493 ( .A1(n10873), .A2(n10872), .B1(P1_REG1_REG_16__SCAN_IN), 
        .B2(n11274), .ZN(n11139) );
  XNOR2_X1 U13494 ( .A(n11298), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n11138) );
  XOR2_X1 U13495 ( .A(n11139), .B(n11138), .Z(n10874) );
  NAND2_X1 U13496 ( .A1(n14652), .A2(n10874), .ZN(n10875) );
  NAND2_X1 U13497 ( .A1(n13742), .A2(n10875), .ZN(n10876) );
  AOI21_X1 U13498 ( .B1(n14633), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n10876), 
        .ZN(n10877) );
  OAI211_X1 U13499 ( .C1(n14670), .C2(n11137), .A(n10878), .B(n10877), .ZN(
        P1_U3260) );
  OAI211_X1 U13500 ( .C1(n10881), .C2(n10880), .A(n10879), .B(n12216), .ZN(
        n10888) );
  AOI21_X1 U13501 ( .B1(n14888), .B2(n12493), .A(n10882), .ZN(n10883) );
  OAI21_X1 U13502 ( .B1(n10884), .B2(n12227), .A(n10883), .ZN(n10885) );
  AOI21_X1 U13503 ( .B1(n12268), .B2(n10886), .A(n10885), .ZN(n10887) );
  OAI211_X1 U13504 ( .C1(n12266), .C2(n10937), .A(n10888), .B(n10887), .ZN(
        P3_U3161) );
  XNOR2_X1 U13505 ( .A(n10889), .B(n12107), .ZN(n13480) );
  NAND2_X1 U13506 ( .A1(n10890), .A2(n13479), .ZN(n10891) );
  NAND2_X1 U13507 ( .A1(n10891), .A2(n8927), .ZN(n10892) );
  NOR2_X1 U13508 ( .A1(n10976), .A2(n10892), .ZN(n13481) );
  INV_X1 U13509 ( .A(n10893), .ZN(n10895) );
  OAI211_X1 U13510 ( .C1(n10895), .C2(n12107), .A(n13421), .B(n10894), .ZN(
        n10897) );
  NAND2_X1 U13511 ( .A1(n10897), .A2(n10896), .ZN(n13475) );
  AOI211_X1 U13512 ( .C1(n13584), .C2(n13480), .A(n13481), .B(n13475), .ZN(
        n10902) );
  INV_X1 U13513 ( .A(n13640), .ZN(n13646) );
  INV_X1 U13514 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10898) );
  NOR2_X1 U13515 ( .A1(n14880), .A2(n10898), .ZN(n10899) );
  AOI21_X1 U13516 ( .B1(n13646), .B2(n13479), .A(n10899), .ZN(n10900) );
  OAI21_X1 U13517 ( .B1(n10902), .B2(n14879), .A(n10900), .ZN(P2_U3460) );
  AOI22_X1 U13518 ( .A1(n13596), .A2(n13479), .B1(n14883), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n10901) );
  OAI21_X1 U13519 ( .B1(n10902), .B2(n14883), .A(n10901), .ZN(P2_U3509) );
  XNOR2_X1 U13520 ( .A(n10903), .B(n12300), .ZN(n15025) );
  OAI22_X1 U13521 ( .A1(n12866), .A2(n15022), .B1(n10904), .B2(n12864), .ZN(
        n10915) );
  AND2_X1 U13522 ( .A1(n10907), .A2(n10905), .ZN(n10910) );
  NAND2_X1 U13523 ( .A1(n10907), .A2(n10906), .ZN(n10908) );
  OAI211_X1 U13524 ( .C1(n10910), .C2(n10909), .A(n10908), .B(n12837), .ZN(
        n10913) );
  AOI22_X1 U13525 ( .A1(n12495), .A2(n12841), .B1(n12844), .B2(n12497), .ZN(
        n10912) );
  NAND2_X1 U13526 ( .A1(n15025), .A2(n11117), .ZN(n10911) );
  NAND3_X1 U13527 ( .A1(n10913), .A2(n10912), .A3(n10911), .ZN(n15023) );
  MUX2_X1 U13528 ( .A(n15023), .B(P3_REG2_REG_6__SCAN_IN), .S(n12833), .Z(
        n10914) );
  AOI211_X1 U13529 ( .C1(n15025), .C2(n12647), .A(n10915), .B(n10914), .ZN(
        n10916) );
  INV_X1 U13530 ( .A(n10916), .ZN(P3_U3227) );
  INV_X1 U13531 ( .A(n11435), .ZN(n14749) );
  AOI22_X1 U13532 ( .A1(n11435), .A2(n11801), .B1(n11863), .B2(n13808), .ZN(
        n11212) );
  AOI22_X1 U13533 ( .A1(n11435), .A2(n11858), .B1(n11801), .B2(n13808), .ZN(
        n10917) );
  XNOR2_X1 U13534 ( .A(n10917), .B(n11217), .ZN(n11213) );
  XOR2_X1 U13535 ( .A(n11212), .B(n11213), .Z(n10923) );
  OAI21_X1 U13536 ( .B1(n10923), .B2(n10922), .A(n11214), .ZN(n10924) );
  NAND2_X1 U13537 ( .A1(n10924), .A2(n14527), .ZN(n10930) );
  INV_X1 U13538 ( .A(n14502), .ZN(n13746) );
  OAI22_X1 U13539 ( .A1(n14503), .A2(n10926), .B1(n14628), .B2(n10925), .ZN(
        n10927) );
  AOI211_X1 U13540 ( .C1(n13746), .C2(n14765), .A(n10928), .B(n10927), .ZN(
        n10929) );
  OAI211_X1 U13541 ( .C1(n14749), .C2(n14500), .A(n10930), .B(n10929), .ZN(
        P1_U3221) );
  XNOR2_X1 U13542 ( .A(n10931), .B(n12369), .ZN(n15035) );
  INV_X1 U13543 ( .A(n15035), .ZN(n10941) );
  INV_X1 U13544 ( .A(n10948), .ZN(n10932) );
  AOI21_X1 U13545 ( .B1(n12369), .B2(n10933), .A(n10932), .ZN(n10936) );
  AOI22_X1 U13546 ( .A1(n12495), .A2(n12844), .B1(n12841), .B2(n12493), .ZN(
        n10935) );
  NAND2_X1 U13547 ( .A1(n15035), .A2(n11117), .ZN(n10934) );
  OAI211_X1 U13548 ( .C1(n10936), .C2(n12858), .A(n10935), .B(n10934), .ZN(
        n15033) );
  NAND2_X1 U13549 ( .A1(n15033), .A2(n12863), .ZN(n10940) );
  OAI22_X1 U13550 ( .A1(n12866), .A2(n15032), .B1(n10937), .B2(n12864), .ZN(
        n10938) );
  AOI21_X1 U13551 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n12868), .A(n10938), .ZN(
        n10939) );
  OAI211_X1 U13552 ( .C1(n10941), .C2(n10957), .A(n10940), .B(n10939), .ZN(
        P3_U3225) );
  INV_X1 U13553 ( .A(n10942), .ZN(n10944) );
  OAI222_X1 U13554 ( .A1(P3_U3151), .A2(n10945), .B1(n12997), .B2(n10944), 
        .C1(n10943), .C2(n12995), .ZN(P3_U3270) );
  OAI222_X1 U13555 ( .A1(n14276), .A2(n11528), .B1(n14270), .B2(n11527), .C1(
        n6978), .C2(P1_U3086), .ZN(P1_U3334) );
  XNOR2_X1 U13556 ( .A(n10946), .B(n12301), .ZN(n15040) );
  AND2_X1 U13557 ( .A1(n10948), .A2(n10947), .ZN(n10950) );
  OAI211_X1 U13558 ( .C1(n10950), .C2(n12301), .A(n12837), .B(n10949), .ZN(
        n10952) );
  AOI22_X1 U13559 ( .A1(n12844), .A2(n12494), .B1(n12492), .B2(n12841), .ZN(
        n10951) );
  OAI211_X1 U13560 ( .C1(n10953), .C2(n15040), .A(n10952), .B(n10951), .ZN(
        n15042) );
  NAND2_X1 U13561 ( .A1(n15042), .A2(n12863), .ZN(n10956) );
  OAI22_X1 U13562 ( .A1(n12866), .A2(n15038), .B1(n11105), .B2(n12864), .ZN(
        n10954) );
  AOI21_X1 U13563 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n12868), .A(n10954), .ZN(
        n10955) );
  OAI211_X1 U13564 ( .C1(n15040), .C2(n10957), .A(n10956), .B(n10955), .ZN(
        P3_U3224) );
  NAND2_X1 U13565 ( .A1(n10958), .A2(n10959), .ZN(n10963) );
  NAND2_X1 U13566 ( .A1(n11123), .A2(n10960), .ZN(n10962) );
  OR2_X1 U13567 ( .A1(n10963), .A2(n10962), .ZN(n11124) );
  INV_X1 U13568 ( .A(n11124), .ZN(n10961) );
  AOI21_X1 U13569 ( .B1(n10963), .B2(n10962), .A(n10961), .ZN(n10968) );
  OAI22_X1 U13570 ( .A1(n13072), .A2(n11160), .B1(n13118), .B2(n11164), .ZN(
        n10964) );
  AOI211_X1 U13571 ( .C1(n11095), .C2(n13135), .A(n10965), .B(n10964), .ZN(
        n10967) );
  NAND2_X1 U13572 ( .A1(n11944), .A2(n13120), .ZN(n10966) );
  OAI211_X1 U13573 ( .C1(n10968), .C2(n13122), .A(n10967), .B(n10966), .ZN(
        P2_U3196) );
  XNOR2_X1 U13574 ( .A(n10969), .B(n12111), .ZN(n13602) );
  INV_X1 U13575 ( .A(n10970), .ZN(n10971) );
  AOI21_X1 U13576 ( .B1(n12111), .B2(n10972), .A(n10971), .ZN(n10974) );
  OAI21_X1 U13577 ( .B1(n10974), .B2(n13459), .A(n10973), .ZN(n13598) );
  OAI21_X1 U13578 ( .B1(n10976), .B2(n10975), .A(n8927), .ZN(n10977) );
  NOR2_X1 U13579 ( .A1(n10977), .A2(n11167), .ZN(n13599) );
  NAND2_X1 U13580 ( .A1(n13599), .A2(n14833), .ZN(n10982) );
  OAI22_X1 U13581 ( .A1(n13490), .A2(n10979), .B1(n10978), .B2(n13487), .ZN(
        n10980) );
  AOI21_X1 U13582 ( .B1(n13600), .B2(n13493), .A(n10980), .ZN(n10981) );
  NAND2_X1 U13583 ( .A1(n10982), .A2(n10981), .ZN(n10983) );
  AOI21_X1 U13584 ( .B1(n13598), .B2(n13490), .A(n10983), .ZN(n10984) );
  OAI21_X1 U13585 ( .B1(n13602), .B2(n13474), .A(n10984), .ZN(P2_U3254) );
  NOR2_X1 U13586 ( .A1(n10994), .A2(n10985), .ZN(n10987) );
  INV_X1 U13587 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10988) );
  OR2_X1 U13588 ( .A1(n14967), .A2(n10988), .ZN(n10990) );
  NAND2_X1 U13589 ( .A1(n14967), .A2(n10988), .ZN(n10989) );
  NAND2_X1 U13590 ( .A1(n10990), .A2(n10989), .ZN(n14956) );
  AOI21_X1 U13591 ( .B1(n11004), .B2(n10991), .A(n11077), .ZN(n11022) );
  NOR2_X1 U13592 ( .A1(n10994), .A2(n10993), .ZN(n10996) );
  OR2_X1 U13593 ( .A1(n14967), .A2(n10997), .ZN(n10999) );
  NAND2_X1 U13594 ( .A1(n14967), .A2(n10997), .ZN(n10998) );
  NAND2_X1 U13595 ( .A1(n10999), .A2(n10998), .ZN(n14960) );
  AOI21_X1 U13596 ( .B1(n11003), .B2(n11001), .A(n11065), .ZN(n11002) );
  NOR2_X1 U13597 ( .A1(n11002), .A2(n14989), .ZN(n11020) );
  MUX2_X1 U13598 ( .A(n11004), .B(n11003), .S(n12602), .Z(n11005) );
  AND2_X1 U13599 ( .A1(n11005), .A2(n11076), .ZN(n11072) );
  NOR2_X1 U13600 ( .A1(n11005), .A2(n11076), .ZN(n11006) );
  OR2_X1 U13601 ( .A1(n11072), .A2(n11006), .ZN(n11014) );
  MUX2_X1 U13602 ( .A(n10988), .B(n10997), .S(n12602), .Z(n11011) );
  AND2_X1 U13603 ( .A1(n11011), .A2(n14967), .ZN(n11012) );
  AOI21_X1 U13604 ( .B1(n11009), .B2(n11008), .A(n11007), .ZN(n14965) );
  INV_X1 U13605 ( .A(n11012), .ZN(n11010) );
  OAI21_X1 U13606 ( .B1(n14967), .B2(n11011), .A(n11010), .ZN(n14966) );
  AOI21_X1 U13607 ( .B1(n11014), .B2(n11013), .A(n11071), .ZN(n11018) );
  NOR2_X1 U13608 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11015), .ZN(n11349) );
  AOI21_X1 U13609 ( .B1(n14972), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11349), 
        .ZN(n11017) );
  NAND2_X1 U13610 ( .A1(n14944), .A2(n11076), .ZN(n11016) );
  OAI211_X1 U13611 ( .C1(n11018), .C2(n14987), .A(n11017), .B(n11016), .ZN(
        n11019) );
  NOR2_X1 U13612 ( .A1(n11020), .A2(n11019), .ZN(n11021) );
  OAI21_X1 U13613 ( .B1(n11022), .B2(n14995), .A(n11021), .ZN(P3_U3193) );
  INV_X1 U13614 ( .A(n14519), .ZN(n11023) );
  OR2_X1 U13615 ( .A1(n13712), .A2(n11023), .ZN(n11024) );
  NAND2_X1 U13616 ( .A1(n11026), .A2(n11641), .ZN(n11030) );
  OAI22_X1 U13617 ( .A1(n11027), .A2(n11545), .B1(n11655), .B2(n15111), .ZN(
        n11028) );
  INV_X1 U13618 ( .A(n11028), .ZN(n11029) );
  XNOR2_X1 U13619 ( .A(n14570), .B(n14504), .ZN(n14433) );
  INV_X1 U13620 ( .A(n14433), .ZN(n14430) );
  NAND2_X1 U13621 ( .A1(n14431), .A2(n14430), .ZN(n14429) );
  OR2_X1 U13622 ( .A1(n14570), .A2(n14504), .ZN(n11031) );
  NAND2_X1 U13623 ( .A1(n14429), .A2(n11031), .ZN(n11042) );
  NAND2_X1 U13624 ( .A1(n11032), .A2(n11641), .ZN(n11035) );
  AOI22_X1 U13625 ( .A1(n11033), .A2(n11501), .B1(n11502), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11034) );
  NOR2_X1 U13626 ( .A1(n11036), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n11037) );
  OR2_X1 U13627 ( .A1(n11044), .A2(n11037), .ZN(n14510) );
  INV_X1 U13628 ( .A(n14510), .ZN(n11043) );
  NAND2_X1 U13629 ( .A1(n10112), .A2(n11043), .ZN(n11041) );
  NAND2_X1 U13630 ( .A1(n11599), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11040) );
  NAND2_X1 U13631 ( .A1(n11657), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11039) );
  NAND2_X1 U13632 ( .A1(n9899), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11038) );
  NAND2_X1 U13633 ( .A1(n11767), .A2(n14421), .ZN(n11467) );
  NAND2_X1 U13634 ( .A1(n11468), .A2(n11467), .ZN(n11689) );
  OAI211_X1 U13635 ( .C1(n11042), .C2(n11061), .A(n11172), .B(n14763), .ZN(
        n14563) );
  AOI22_X1 U13636 ( .A1(n14704), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n11043), 
        .B2(n14682), .ZN(n11051) );
  NAND2_X1 U13637 ( .A1(n11599), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11049) );
  NAND2_X1 U13638 ( .A1(n11657), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11048) );
  OR2_X1 U13639 ( .A1(n11044), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11045) );
  AND2_X1 U13640 ( .A1(n11183), .A2(n11045), .ZN(n13799) );
  NAND2_X1 U13641 ( .A1(n11646), .A2(n13799), .ZN(n11047) );
  NAND2_X1 U13642 ( .A1(n11614), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11046) );
  INV_X1 U13643 ( .A(n14501), .ZN(n14559) );
  NAND2_X1 U13644 ( .A1(n14061), .A2(n14559), .ZN(n11050) );
  OAI211_X1 U13645 ( .C1(n14504), .C2(n14064), .A(n11051), .B(n11050), .ZN(
        n11054) );
  AOI21_X1 U13646 ( .B1(n11767), .B2(n14418), .A(n14572), .ZN(n11052) );
  NAND2_X1 U13647 ( .A1(n11052), .A2(n11181), .ZN(n14561) );
  NOR2_X1 U13648 ( .A1(n14561), .A2(n14066), .ZN(n11053) );
  AOI211_X1 U13649 ( .C1(n14683), .C2(n11767), .A(n11054), .B(n11053), .ZN(
        n11064) );
  INV_X1 U13650 ( .A(n11687), .ZN(n11055) );
  NAND2_X1 U13651 ( .A1(n11056), .A2(n11055), .ZN(n11058) );
  OR2_X1 U13652 ( .A1(n13712), .A2(n14519), .ZN(n11057) );
  NAND2_X1 U13653 ( .A1(n11058), .A2(n11057), .ZN(n14432) );
  OR2_X1 U13654 ( .A1(n14570), .A2(n14558), .ZN(n11059) );
  NAND2_X1 U13655 ( .A1(n11062), .A2(n11061), .ZN(n14557) );
  NAND3_X1 U13656 ( .A1(n14566), .A2(n14557), .A3(n14544), .ZN(n11063) );
  OAI211_X1 U13657 ( .C1(n14563), .C2(n14704), .A(n11064), .B(n11063), .ZN(
        P1_U3279) );
  NAND2_X1 U13658 ( .A1(n11083), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12501) );
  NAND2_X1 U13659 ( .A1(n12514), .A2(n11066), .ZN(n11067) );
  NAND2_X1 U13660 ( .A1(n12501), .A2(n11067), .ZN(n11069) );
  INV_X1 U13661 ( .A(n12502), .ZN(n11068) );
  AOI21_X1 U13662 ( .B1(n11070), .B2(n11069), .A(n11068), .ZN(n11087) );
  INV_X1 U13663 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11073) );
  MUX2_X1 U13664 ( .A(n11073), .B(n11066), .S(n12602), .Z(n12513) );
  XNOR2_X1 U13665 ( .A(n12513), .B(n12514), .ZN(n12515) );
  XNOR2_X1 U13666 ( .A(n12516), .B(n12515), .ZN(n11085) );
  INV_X1 U13667 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11074) );
  NOR2_X1 U13668 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11074), .ZN(n11339) );
  AOI21_X1 U13669 ( .B1(n14972), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11339), 
        .ZN(n11082) );
  NOR2_X1 U13670 ( .A1(n11076), .A2(n11075), .ZN(n11078) );
  NAND2_X1 U13671 ( .A1(n11083), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12508) );
  NAND2_X1 U13672 ( .A1(n12514), .A2(n11073), .ZN(n11079) );
  NAND2_X1 U13673 ( .A1(n12508), .A2(n11079), .ZN(n12506) );
  XNOR2_X1 U13674 ( .A(n12507), .B(n12506), .ZN(n11080) );
  NAND2_X1 U13675 ( .A1(n14897), .A2(n11080), .ZN(n11081) );
  OAI211_X1 U13676 ( .C1(n14979), .C2(n11083), .A(n11082), .B(n11081), .ZN(
        n11084) );
  AOI21_X1 U13677 ( .B1(n14945), .B2(n11085), .A(n11084), .ZN(n11086) );
  OAI21_X1 U13678 ( .B1(n11087), .B2(n14989), .A(n11086), .ZN(P3_U3194) );
  INV_X1 U13679 ( .A(n13589), .ZN(n13470) );
  OAI21_X1 U13680 ( .B1(n11090), .B2(n11088), .A(n11089), .ZN(n11091) );
  NAND2_X1 U13681 ( .A1(n11091), .A2(n13098), .ZN(n11097) );
  INV_X1 U13682 ( .A(n11092), .ZN(n11094) );
  OAI22_X1 U13683 ( .A1(n13072), .A2(n13463), .B1(n13118), .B2(n13467), .ZN(
        n11093) );
  AOI211_X1 U13684 ( .C1(n11095), .C2(n13425), .A(n11094), .B(n11093), .ZN(
        n11096) );
  OAI211_X1 U13685 ( .C1(n13470), .C2(n13077), .A(n11097), .B(n11096), .ZN(
        P2_U3187) );
  INV_X1 U13686 ( .A(n11098), .ZN(n11099) );
  AOI21_X1 U13687 ( .B1(n11101), .B2(n11100), .A(n11099), .ZN(n11110) );
  AOI21_X1 U13688 ( .B1(n12492), .B2(n14888), .A(n11102), .ZN(n11103) );
  OAI21_X1 U13689 ( .B1(n11104), .B2(n12227), .A(n11103), .ZN(n11107) );
  NOR2_X1 U13690 ( .A1(n12266), .A2(n11105), .ZN(n11106) );
  AOI211_X1 U13691 ( .C1(n11108), .C2(n12268), .A(n11107), .B(n11106), .ZN(
        n11109) );
  OAI21_X1 U13692 ( .B1(n11110), .B2(n14886), .A(n11109), .ZN(P3_U3171) );
  OAI222_X1 U13693 ( .A1(n13671), .A2(n11111), .B1(P2_U3088), .B2(n7508), .C1(
        n13666), .C2(n11527), .ZN(P2_U3306) );
  XNOR2_X1 U13694 ( .A(n11112), .B(n12304), .ZN(n11113) );
  OAI222_X1 U13695 ( .A1(n12862), .A2(n12859), .B1(n12860), .B2(n11114), .C1(
        n11113), .C2(n12858), .ZN(n15046) );
  INV_X1 U13696 ( .A(n15046), .ZN(n11122) );
  XNOR2_X1 U13697 ( .A(n11115), .B(n12304), .ZN(n15048) );
  NOR2_X1 U13698 ( .A1(n11117), .A2(n11116), .ZN(n11118) );
  NOR2_X1 U13699 ( .A1(n12863), .A2(n10988), .ZN(n11120) );
  OAI22_X1 U13700 ( .A1(n12866), .A2(n15045), .B1(n11235), .B2(n12864), .ZN(
        n11119) );
  AOI211_X1 U13701 ( .C1(n15048), .C2(n12831), .A(n11120), .B(n11119), .ZN(
        n11121) );
  OAI21_X1 U13702 ( .B1(n11122), .B2(n12833), .A(n11121), .ZN(P3_U3223) );
  NAND2_X1 U13703 ( .A1(n11124), .A2(n11123), .ZN(n11126) );
  XOR2_X1 U13704 ( .A(n11126), .B(n11125), .Z(n11132) );
  OAI22_X1 U13705 ( .A1(n13093), .A2(n12093), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11127), .ZN(n11130) );
  OAI22_X1 U13706 ( .A1(n13072), .A2(n11128), .B1(n13118), .B2(n11150), .ZN(
        n11129) );
  AOI211_X1 U13707 ( .C1(n13645), .C2(n13120), .A(n11130), .B(n11129), .ZN(
        n11131) );
  OAI21_X1 U13708 ( .B1(n11132), .B2(n13122), .A(n11131), .ZN(P2_U3206) );
  NAND2_X1 U13709 ( .A1(n11298), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11134) );
  NAND2_X1 U13710 ( .A1(n11134), .A2(n11133), .ZN(n13852) );
  XOR2_X1 U13711 ( .A(n13851), .B(n13852), .Z(n11135) );
  NAND2_X1 U13712 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n11135), .ZN(n13854) );
  OAI211_X1 U13713 ( .C1(n11135), .C2(P1_REG2_REG_18__SCAN_IN), .A(n14643), 
        .B(n13854), .ZN(n11144) );
  NAND2_X1 U13714 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13778)
         );
  INV_X1 U13715 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n11136) );
  OAI22_X1 U13716 ( .A1(n11139), .A2(n11138), .B1(n11137), .B2(n11136), .ZN(
        n13846) );
  XOR2_X1 U13717 ( .A(n13851), .B(n13846), .Z(n11140) );
  NAND2_X1 U13718 ( .A1(n11140), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n13848) );
  OAI211_X1 U13719 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n11140), .A(n14652), 
        .B(n13848), .ZN(n11141) );
  NAND2_X1 U13720 ( .A1(n13778), .A2(n11141), .ZN(n11142) );
  AOI21_X1 U13721 ( .B1(n14633), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n11142), 
        .ZN(n11143) );
  OAI211_X1 U13722 ( .C1(n14670), .C2(n11145), .A(n11144), .B(n11143), .ZN(
        P1_U3261) );
  XNOR2_X1 U13723 ( .A(n11146), .B(n12112), .ZN(n11147) );
  NAND2_X1 U13724 ( .A1(n11147), .A2(n13421), .ZN(n11149) );
  AOI22_X1 U13725 ( .A1(n13426), .A2(n13136), .B1(n13134), .B2(n13427), .ZN(
        n11148) );
  AND2_X1 U13726 ( .A1(n11149), .A2(n11148), .ZN(n13593) );
  OAI22_X1 U13727 ( .A1(n13490), .A2(n11151), .B1(n11150), .B2(n13487), .ZN(
        n11154) );
  AOI21_X1 U13728 ( .B1(n11166), .B2(n13645), .A(n13465), .ZN(n11152) );
  NAND2_X1 U13729 ( .A1(n11152), .A2(n13466), .ZN(n13592) );
  NOR2_X1 U13730 ( .A1(n13592), .A2(n13410), .ZN(n11153) );
  AOI211_X1 U13731 ( .C1(n13493), .C2(n13645), .A(n11154), .B(n11153), .ZN(
        n11157) );
  XNOR2_X1 U13732 ( .A(n11155), .B(n12112), .ZN(n13594) );
  OR2_X1 U13733 ( .A1(n13594), .A2(n13474), .ZN(n11156) );
  OAI211_X1 U13734 ( .C1(n13593), .C2(n15079), .A(n11157), .B(n11156), .ZN(
        P2_U3252) );
  XNOR2_X1 U13735 ( .A(n11944), .B(n13136), .ZN(n12109) );
  XNOR2_X1 U13736 ( .A(n11158), .B(n12109), .ZN(n14491) );
  XNOR2_X1 U13737 ( .A(n11159), .B(n12109), .ZN(n11162) );
  OAI22_X1 U13738 ( .A1(n11160), .A2(n13464), .B1(n13463), .B2(n13462), .ZN(
        n11161) );
  AOI21_X1 U13739 ( .B1(n11162), .B2(n13421), .A(n11161), .ZN(n11163) );
  OAI21_X1 U13740 ( .B1(n14491), .B2(n8915), .A(n11163), .ZN(n14494) );
  NAND2_X1 U13741 ( .A1(n14494), .A2(n13490), .ZN(n11171) );
  OAI22_X1 U13742 ( .A1(n13490), .A2(n11165), .B1(n11164), .B2(n13487), .ZN(
        n11169) );
  OAI211_X1 U13743 ( .C1(n11167), .C2(n14493), .A(n8927), .B(n11166), .ZN(
        n14492) );
  NOR2_X1 U13744 ( .A1(n14492), .A2(n13410), .ZN(n11168) );
  AOI211_X1 U13745 ( .C1(n13493), .C2(n11944), .A(n11169), .B(n11168), .ZN(
        n11170) );
  OAI211_X1 U13746 ( .C1(n14491), .C2(n13393), .A(n11171), .B(n11170), .ZN(
        P2_U3253) );
  NAND2_X1 U13747 ( .A1(n11173), .A2(n11641), .ZN(n11176) );
  AOI22_X1 U13748 ( .A1(n11502), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11501), 
        .B2(n11174), .ZN(n11175) );
  NAND2_X1 U13749 ( .A1(n13804), .A2(n14501), .ZN(n11472) );
  NAND2_X1 U13750 ( .A1(n11471), .A2(n11472), .ZN(n11690) );
  OAI21_X1 U13751 ( .B1(n11177), .B2(n11179), .A(n11272), .ZN(n14552) );
  INV_X1 U13752 ( .A(n14421), .ZN(n14548) );
  NAND2_X1 U13753 ( .A1(n11767), .A2(n14548), .ZN(n11178) );
  OAI21_X1 U13754 ( .B1(n11180), .B2(n11690), .A(n11291), .ZN(n14555) );
  INV_X1 U13755 ( .A(n13804), .ZN(n14551) );
  INV_X1 U13756 ( .A(n11286), .ZN(n11287) );
  OAI211_X1 U13757 ( .C1(n14551), .C2(n6946), .A(n11287), .B(n14686), .ZN(
        n14550) );
  NAND2_X1 U13758 ( .A1(n11614), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11188) );
  NAND2_X1 U13759 ( .A1(n11599), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n11187) );
  INV_X1 U13760 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n11182) );
  NAND2_X1 U13761 ( .A1(n11183), .A2(n11182), .ZN(n11184) );
  AND2_X1 U13762 ( .A1(n11278), .A2(n11184), .ZN(n13730) );
  NAND2_X1 U13763 ( .A1(n11646), .A2(n13730), .ZN(n11186) );
  NAND2_X1 U13764 ( .A1(n11657), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11185) );
  NAND4_X1 U13765 ( .A1(n11188), .A2(n11187), .A3(n11186), .A4(n11185), .ZN(
        n14547) );
  INV_X1 U13766 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11190) );
  INV_X1 U13767 ( .A(n13799), .ZN(n11189) );
  OAI22_X1 U13768 ( .A1(n14437), .A2(n11190), .B1(n11189), .B2(n14706), .ZN(
        n11191) );
  AOI21_X1 U13769 ( .B1(n14061), .B2(n14547), .A(n11191), .ZN(n11192) );
  OAI21_X1 U13770 ( .B1(n14421), .B2(n14064), .A(n11192), .ZN(n11193) );
  AOI21_X1 U13771 ( .B1(n13804), .B2(n14683), .A(n11193), .ZN(n11194) );
  OAI21_X1 U13772 ( .B1(n14550), .B2(n14066), .A(n11194), .ZN(n11195) );
  AOI21_X1 U13773 ( .B1(n14555), .B2(n14544), .A(n11195), .ZN(n11196) );
  OAI21_X1 U13774 ( .B1(n14552), .B2(n14701), .A(n11196), .ZN(P1_U3278) );
  INV_X1 U13775 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11197) );
  OAI22_X1 U13776 ( .A1(n11200), .A2(n11199), .B1(n11198), .B2(n11197), .ZN(
        n13200) );
  XNOR2_X1 U13777 ( .A(n13200), .B(n13199), .ZN(n13198) );
  XOR2_X1 U13778 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13198), .Z(n11211) );
  INV_X1 U13779 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n11201) );
  NAND2_X1 U13780 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13091)
         );
  OAI21_X1 U13781 ( .B1(n13211), .B2(n11201), .A(n13091), .ZN(n11209) );
  NAND2_X1 U13782 ( .A1(n11203), .A2(n11202), .ZN(n11204) );
  NOR2_X1 U13783 ( .A1(n11204), .A2(n13199), .ZN(n13195) );
  AOI21_X1 U13784 ( .B1(n11204), .B2(n13199), .A(n13195), .ZN(n11205) );
  INV_X1 U13785 ( .A(n11205), .ZN(n11206) );
  NOR2_X1 U13786 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n11206), .ZN(n13194) );
  AOI21_X1 U13787 ( .B1(n11206), .B2(P2_REG2_REG_18__SCAN_IN), .A(n13194), 
        .ZN(n11207) );
  NOR2_X1 U13788 ( .A1(n11207), .A2(n14806), .ZN(n11208) );
  AOI211_X1 U13789 ( .C1(n14822), .C2(n13199), .A(n11209), .B(n11208), .ZN(
        n11210) );
  OAI21_X1 U13790 ( .B1(n11211), .B2(n14812), .A(n11210), .ZN(P2_U3232) );
  AND2_X1 U13791 ( .A1(n11863), .A2(n14765), .ZN(n11215) );
  AOI21_X1 U13792 ( .B1(n11440), .B2(n11801), .A(n11215), .ZN(n11252) );
  XNOR2_X1 U13793 ( .A(n11251), .B(n11252), .ZN(n11257) );
  AOI22_X1 U13794 ( .A1(n11440), .A2(n11858), .B1(n11801), .B2(n14765), .ZN(
        n11216) );
  XOR2_X1 U13795 ( .A(n11217), .B(n11216), .Z(n11256) );
  XOR2_X1 U13796 ( .A(n11257), .B(n11256), .Z(n11225) );
  OAI22_X1 U13797 ( .A1(n13733), .A2(n11219), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11218), .ZN(n11220) );
  AOI21_X1 U13798 ( .B1(n11221), .B2(n13798), .A(n11220), .ZN(n11224) );
  INV_X1 U13799 ( .A(n11440), .ZN(n11222) );
  NOR2_X1 U13800 ( .A1(n11222), .A2(n14748), .ZN(n14758) );
  NAND2_X1 U13801 ( .A1(n14758), .A2(n14618), .ZN(n11223) );
  OAI211_X1 U13802 ( .C1(n11225), .C2(n14620), .A(n11224), .B(n11223), .ZN(
        P1_U3231) );
  AOI21_X1 U13803 ( .B1(n11227), .B2(n11226), .A(n14886), .ZN(n11229) );
  NAND2_X1 U13804 ( .A1(n11229), .A2(n11228), .ZN(n11234) );
  NAND2_X1 U13805 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n14962)
         );
  NAND2_X1 U13806 ( .A1(n12264), .A2(n12493), .ZN(n11230) );
  OAI211_X1 U13807 ( .C1(n12859), .C2(n12261), .A(n14962), .B(n11230), .ZN(
        n11231) );
  AOI21_X1 U13808 ( .B1(n12268), .B2(n11232), .A(n11231), .ZN(n11233) );
  OAI211_X1 U13809 ( .C1(n11235), .C2(n12266), .A(n11234), .B(n11233), .ZN(
        P3_U3157) );
  XOR2_X1 U13810 ( .A(n12382), .B(n11236), .Z(n11237) );
  OAI222_X1 U13811 ( .A1(n12862), .A2(n11335), .B1(n12860), .B2(n11352), .C1(
        n11237), .C2(n12858), .ZN(n14482) );
  INV_X1 U13812 ( .A(n14482), .ZN(n11243) );
  XNOR2_X1 U13813 ( .A(n11238), .B(n12382), .ZN(n14484) );
  INV_X1 U13814 ( .A(n11239), .ZN(n11348) );
  AOI22_X1 U13815 ( .A1(n12796), .A2(n12388), .B1(n11348), .B2(n12828), .ZN(
        n11240) );
  OAI21_X1 U13816 ( .B1(n11004), .B2(n12863), .A(n11240), .ZN(n11241) );
  AOI21_X1 U13817 ( .B1(n14484), .B2(n12831), .A(n11241), .ZN(n11242) );
  OAI21_X1 U13818 ( .B1(n11243), .B2(n12833), .A(n11242), .ZN(P3_U3222) );
  XNOR2_X1 U13819 ( .A(n11244), .B(n11245), .ZN(n11250) );
  AOI22_X1 U13820 ( .A1(n13133), .A2(n13427), .B1(n13426), .B2(n13134), .ZN(
        n13442) );
  INV_X1 U13821 ( .A(n13442), .ZN(n11246) );
  AOI22_X1 U13822 ( .A1(n13116), .A2(n11246), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11247) );
  OAI21_X1 U13823 ( .B1(n13444), .B2(n13118), .A(n11247), .ZN(n11248) );
  AOI21_X1 U13824 ( .B1(n13580), .B2(n13120), .A(n11248), .ZN(n11249) );
  OAI21_X1 U13825 ( .B1(n11250), .B2(n13122), .A(n11249), .ZN(P2_U3213) );
  INV_X1 U13826 ( .A(n11251), .ZN(n11254) );
  INV_X1 U13827 ( .A(n11252), .ZN(n11253) );
  OAI21_X2 U13828 ( .B1(n11257), .B2(n11256), .A(n11255), .ZN(n11743) );
  NAND2_X1 U13829 ( .A1(n14768), .A2(n11858), .ZN(n11259) );
  NAND2_X1 U13830 ( .A1(n14520), .A2(n11801), .ZN(n11258) );
  NAND2_X1 U13831 ( .A1(n11259), .A2(n11258), .ZN(n11260) );
  XNOR2_X1 U13832 ( .A(n11260), .B(n11861), .ZN(n11739) );
  AOI22_X1 U13833 ( .A1(n14768), .A2(n11801), .B1(n11863), .B2(n14520), .ZN(
        n11740) );
  XNOR2_X1 U13834 ( .A(n11739), .B(n11740), .ZN(n11742) );
  XOR2_X1 U13835 ( .A(n11743), .B(n11742), .Z(n11267) );
  AOI22_X1 U13836 ( .A1(n13746), .A2(n14404), .B1(n11261), .B2(n13798), .ZN(
        n11263) );
  OAI211_X1 U13837 ( .C1(n11264), .C2(n14503), .A(n11263), .B(n11262), .ZN(
        n11265) );
  AOI21_X1 U13838 ( .B1(n14525), .B2(n14768), .A(n11265), .ZN(n11266) );
  OAI21_X1 U13839 ( .B1(n11267), .B2(n14620), .A(n11266), .ZN(P1_U3217) );
  OAI222_X1 U13840 ( .A1(n13671), .A2(n11269), .B1(P2_U3088), .B2(n11882), 
        .C1(n13666), .C2(n11268), .ZN(P2_U3305) );
  OAI222_X1 U13841 ( .A1(P2_U3088), .A2(n11271), .B1(n13666), .B2(n11581), 
        .C1(n11270), .C2(n13671), .ZN(P2_U3303) );
  OAI222_X1 U13842 ( .A1(n9273), .A2(P1_U3086), .B1(n14270), .B2(n11581), .C1(
        n11582), .C2(n14276), .ZN(P1_U3331) );
  NAND2_X1 U13843 ( .A1(n11273), .A2(n11641), .ZN(n11276) );
  AOI22_X1 U13844 ( .A1(n11502), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11501), 
        .B2(n11274), .ZN(n11275) );
  XNOR2_X1 U13845 ( .A(n14227), .B(n14547), .ZN(n11692) );
  XNOR2_X1 U13846 ( .A(n11302), .B(n11301), .ZN(n11285) );
  OR2_X1 U13847 ( .A1(n14501), .A2(n14209), .ZN(n11283) );
  INV_X1 U13848 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11277) );
  AND2_X1 U13849 ( .A1(n11278), .A2(n11277), .ZN(n11279) );
  OR2_X1 U13850 ( .A1(n11279), .A2(n11308), .ZN(n13743) );
  INV_X1 U13851 ( .A(n11646), .ZN(n11553) );
  AOI22_X1 U13852 ( .A1(n11657), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n11599), 
        .B2(P1_REG0_REG_17__SCAN_IN), .ZN(n11281) );
  NAND2_X1 U13853 ( .A1(n11614), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n11280) );
  OAI211_X1 U13854 ( .C1(n13743), .C2(n11553), .A(n11281), .B(n11280), .ZN(
        n14093) );
  NAND2_X1 U13855 ( .A1(n14093), .A2(n14745), .ZN(n11282) );
  AND2_X1 U13856 ( .A1(n11283), .A2(n11282), .ZN(n13734) );
  INV_X1 U13857 ( .A(n13734), .ZN(n11284) );
  AOI21_X1 U13858 ( .B1(n11285), .B2(n14763), .A(n11284), .ZN(n14229) );
  INV_X1 U13859 ( .A(n14227), .ZN(n11289) );
  AOI211_X1 U13860 ( .C1(n14227), .C2(n11287), .A(n14572), .B(n11306), .ZN(
        n14226) );
  AOI22_X1 U13861 ( .A1(n14704), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n13730), 
        .B2(n14682), .ZN(n11288) );
  OAI21_X1 U13862 ( .B1(n11289), .B2(n14096), .A(n11288), .ZN(n11293) );
  OR2_X1 U13863 ( .A1(n13804), .A2(n14559), .ZN(n11290) );
  XNOR2_X1 U13864 ( .A(n11295), .B(n11692), .ZN(n14230) );
  NOR2_X1 U13865 ( .A1(n14230), .A2(n14700), .ZN(n11292) );
  AOI211_X1 U13866 ( .C1(n14226), .C2(n14690), .A(n11293), .B(n11292), .ZN(
        n11294) );
  OAI21_X1 U13867 ( .B1(n14704), .B2(n14229), .A(n11294), .ZN(P1_U3277) );
  OR2_X1 U13868 ( .A1(n14227), .A2(n14547), .ZN(n11296) );
  NAND2_X1 U13869 ( .A1(n11297), .A2(n11641), .ZN(n11300) );
  AOI22_X1 U13870 ( .A1(n11502), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11501), 
        .B2(n11298), .ZN(n11299) );
  XNOR2_X1 U13871 ( .A(n11492), .B(n14093), .ZN(n11691) );
  XNOR2_X1 U13872 ( .A(n13878), .B(n11691), .ZN(n14225) );
  INV_X1 U13873 ( .A(n11691), .ZN(n11305) );
  INV_X1 U13874 ( .A(n14547), .ZN(n13802) );
  INV_X1 U13875 ( .A(n13896), .ZN(n11303) );
  AOI21_X1 U13876 ( .B1(n11305), .B2(n11304), .A(n11303), .ZN(n14223) );
  OAI21_X1 U13877 ( .B1(n11306), .B2(n14221), .A(n14686), .ZN(n11307) );
  OR2_X1 U13878 ( .A1(n14086), .A2(n11307), .ZN(n14220) );
  NOR2_X1 U13879 ( .A1(n14706), .A2(n13743), .ZN(n11314) );
  INV_X1 U13880 ( .A(n14061), .ZN(n14091) );
  OR2_X1 U13881 ( .A1(n11308), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11309) );
  AND2_X1 U13882 ( .A1(n11517), .A2(n11309), .ZN(n14089) );
  NAND2_X1 U13883 ( .A1(n14089), .A2(n11646), .ZN(n11312) );
  AOI22_X1 U13884 ( .A1(n11657), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n11599), 
        .B2(P1_REG0_REG_18__SCAN_IN), .ZN(n11311) );
  NAND2_X1 U13885 ( .A1(n11614), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n11310) );
  NOR2_X1 U13886 ( .A1(n14091), .A2(n14202), .ZN(n11313) );
  AOI211_X1 U13887 ( .C1(n14704), .C2(P1_REG2_REG_17__SCAN_IN), .A(n11314), 
        .B(n11313), .ZN(n11315) );
  OAI21_X1 U13888 ( .B1(n13802), .B2(n14064), .A(n11315), .ZN(n11316) );
  AOI21_X1 U13889 ( .B1(n11492), .B2(n14683), .A(n11316), .ZN(n11317) );
  OAI21_X1 U13890 ( .B1(n14220), .B2(n14066), .A(n11317), .ZN(n11318) );
  AOI21_X1 U13891 ( .B1(n14223), .B2(n14434), .A(n11318), .ZN(n11319) );
  OAI21_X1 U13892 ( .B1(n14700), .B2(n14225), .A(n11319), .ZN(P1_U3276) );
  OAI222_X1 U13893 ( .A1(n11322), .A2(P3_U3151), .B1(n12997), .B2(n11321), 
        .C1(n11320), .C2(n12995), .ZN(P3_U3269) );
  OAI222_X1 U13894 ( .A1(n14276), .A2(n11612), .B1(n14270), .B2(n13659), .C1(
        n14631), .C2(P1_U3086), .ZN(P1_U3328) );
  INV_X1 U13895 ( .A(n11642), .ZN(n14259) );
  OAI222_X1 U13896 ( .A1(n13666), .A2(n14259), .B1(P2_U3088), .B2(n11324), 
        .C1(n11323), .C2(n13671), .ZN(P2_U3298) );
  AOI222_X1 U13897 ( .A1(n11326), .A2(n14397), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11325), .C1(SI_3_), .C2(n14396), .ZN(n11327) );
  INV_X1 U13898 ( .A(n11327), .ZN(P3_U3292) );
  XOR2_X1 U13899 ( .A(n11329), .B(n11328), .Z(n13814) );
  NAND2_X1 U13900 ( .A1(n13814), .A2(n14527), .ZN(n11333) );
  AOI22_X1 U13901 ( .A1(n14525), .A2(n11331), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n11330), .ZN(n11332) );
  OAI211_X1 U13902 ( .C1(n11334), .C2(n14502), .A(n11333), .B(n11332), .ZN(
        P1_U3232) );
  XNOR2_X1 U13903 ( .A(n11336), .B(n11335), .ZN(n11337) );
  XNOR2_X1 U13904 ( .A(n11338), .B(n11337), .ZN(n11345) );
  INV_X1 U13905 ( .A(n12865), .ZN(n11343) );
  AOI21_X1 U13906 ( .B1(n12821), .B2(n14888), .A(n11339), .ZN(n11341) );
  OR2_X1 U13907 ( .A1(n12859), .A2(n12227), .ZN(n11340) );
  OAI211_X1 U13908 ( .C1(n14891), .C2(n14477), .A(n11341), .B(n11340), .ZN(
        n11342) );
  AOI21_X1 U13909 ( .B1(n11343), .B2(n12243), .A(n11342), .ZN(n11344) );
  OAI21_X1 U13910 ( .B1(n11345), .B2(n14886), .A(n11344), .ZN(P3_U3164) );
  NAND2_X1 U13911 ( .A1(n11346), .A2(n7448), .ZN(n11347) );
  XNOR2_X1 U13912 ( .A(n11347), .B(n12859), .ZN(n11355) );
  NAND2_X1 U13913 ( .A1(n12243), .A2(n11348), .ZN(n11351) );
  AOI21_X1 U13914 ( .B1(n14888), .B2(n12843), .A(n11349), .ZN(n11350) );
  OAI211_X1 U13915 ( .C1(n11352), .C2(n12227), .A(n11351), .B(n11350), .ZN(
        n11353) );
  AOI21_X1 U13916 ( .B1(n12388), .B2(n12268), .A(n11353), .ZN(n11354) );
  OAI21_X1 U13917 ( .B1(n11355), .B2(n14886), .A(n11354), .ZN(P3_U3176) );
  NAND2_X1 U13918 ( .A1(n11358), .A2(n12992), .ZN(n11359) );
  MUX2_X1 U13919 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n11363), .Z(n11361) );
  XNOR2_X1 U13920 ( .A(n11361), .B(SI_30_), .ZN(n11651) );
  NAND2_X1 U13921 ( .A1(n11361), .A2(SI_30_), .ZN(n11362) );
  MUX2_X1 U13922 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n11363), .Z(n11364) );
  XNOR2_X1 U13923 ( .A(n11364), .B(SI_31_), .ZN(n11365) );
  NAND2_X1 U13924 ( .A1(n14254), .A2(n11641), .ZN(n11368) );
  INV_X1 U13925 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14251) );
  OR2_X1 U13926 ( .A1(n11655), .A2(n14251), .ZN(n11367) );
  NOR2_X1 U13927 ( .A1(n13867), .A2(n11422), .ZN(n11708) );
  NAND2_X1 U13928 ( .A1(n11614), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n11373) );
  NAND2_X1 U13929 ( .A1(n11657), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n11372) );
  NAND2_X1 U13930 ( .A1(n11599), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n11371) );
  AND3_X1 U13931 ( .A1(n11373), .A2(n11372), .A3(n11371), .ZN(n13870) );
  INV_X1 U13932 ( .A(n13870), .ZN(n13807) );
  INV_X1 U13933 ( .A(n14279), .ZN(n11374) );
  NAND2_X1 U13934 ( .A1(n11375), .A2(n11374), .ZN(n11376) );
  NAND2_X1 U13935 ( .A1(n11377), .A2(n11376), .ZN(n11378) );
  NAND2_X1 U13936 ( .A1(n11378), .A2(n14106), .ZN(n11713) );
  NAND2_X1 U13937 ( .A1(n6978), .A2(n11379), .ZN(n11712) );
  NAND2_X1 U13938 ( .A1(n11713), .A2(n11712), .ZN(n11704) );
  NAND2_X1 U13939 ( .A1(n13867), .A2(n11422), .ZN(n11706) );
  NOR2_X1 U13940 ( .A1(n11706), .A2(n13807), .ZN(n11380) );
  AOI211_X1 U13941 ( .C1(n11708), .C2(n13807), .A(n11704), .B(n11380), .ZN(
        n11718) );
  NAND2_X1 U13942 ( .A1(n11397), .A2(n7375), .ZN(n11385) );
  INV_X1 U13943 ( .A(n11381), .ZN(n11382) );
  NAND2_X1 U13944 ( .A1(n11382), .A2(n11391), .ZN(n11384) );
  NAND4_X1 U13945 ( .A1(n11385), .A2(n11384), .A3(n11422), .A4(n11383), .ZN(
        n11387) );
  OR2_X1 U13946 ( .A1(n11387), .A2(n11386), .ZN(n11408) );
  AOI21_X1 U13947 ( .B1(n9693), .B2(n11388), .A(n9684), .ZN(n11389) );
  AND2_X1 U13948 ( .A1(n11391), .A2(n6443), .ZN(n11392) );
  NAND4_X1 U13949 ( .A1(n11394), .A2(n11393), .A3(n11392), .A4(n11396), .ZN(
        n11407) );
  MUX2_X1 U13950 ( .A(n11396), .B(n11395), .S(n6443), .Z(n11406) );
  OR3_X1 U13951 ( .A1(n11397), .A2(n13812), .A3(n11399), .ZN(n11402) );
  INV_X1 U13952 ( .A(n11398), .ZN(n11400) );
  NAND3_X1 U13953 ( .A1(n11400), .A2(n11399), .A3(n13812), .ZN(n11401) );
  NAND2_X1 U13954 ( .A1(n11402), .A2(n11401), .ZN(n11403) );
  NAND2_X1 U13955 ( .A1(n11404), .A2(n11403), .ZN(n11405) );
  NAND4_X1 U13956 ( .A1(n11408), .A2(n11407), .A3(n11406), .A4(n11405), .ZN(
        n11414) );
  MUX2_X1 U13957 ( .A(n11410), .B(n11409), .S(n11422), .Z(n11413) );
  MUX2_X1 U13958 ( .A(n6446), .B(n11411), .S(n6443), .Z(n11412) );
  OAI21_X1 U13959 ( .B1(n11414), .B2(n11413), .A(n11412), .ZN(n11416) );
  NAND2_X1 U13960 ( .A1(n11414), .A2(n11413), .ZN(n11415) );
  MUX2_X1 U13961 ( .A(n13810), .B(n11417), .S(n6443), .Z(n11420) );
  MUX2_X1 U13963 ( .A(n13810), .B(n11417), .S(n11609), .Z(n11418) );
  INV_X1 U13964 ( .A(n11420), .ZN(n11421) );
  MUX2_X1 U13965 ( .A(n13809), .B(n14727), .S(n11609), .Z(n11425) );
  MUX2_X1 U13966 ( .A(n13809), .B(n14727), .S(n6443), .Z(n11423) );
  NAND2_X1 U13967 ( .A1(n11424), .A2(n11423), .ZN(n11426) );
  MUX2_X1 U13968 ( .A(n14744), .B(n14684), .S(n6443), .Z(n11430) );
  NAND2_X1 U13969 ( .A1(n11429), .A2(n11430), .ZN(n11428) );
  MUX2_X1 U13970 ( .A(n14744), .B(n14684), .S(n11609), .Z(n11427) );
  NAND2_X1 U13971 ( .A1(n11428), .A2(n11427), .ZN(n11434) );
  INV_X1 U13972 ( .A(n11429), .ZN(n11432) );
  INV_X1 U13973 ( .A(n11430), .ZN(n11431) );
  NAND2_X1 U13974 ( .A1(n11432), .A2(n11431), .ZN(n11433) );
  NAND2_X1 U13975 ( .A1(n11434), .A2(n11433), .ZN(n11437) );
  MUX2_X1 U13976 ( .A(n13808), .B(n11435), .S(n11609), .Z(n11438) );
  MUX2_X1 U13977 ( .A(n13808), .B(n11435), .S(n6443), .Z(n11436) );
  INV_X1 U13978 ( .A(n11438), .ZN(n11439) );
  MUX2_X1 U13979 ( .A(n14765), .B(n11440), .S(n6443), .Z(n11444) );
  MUX2_X1 U13980 ( .A(n14765), .B(n11440), .S(n11609), .Z(n11441) );
  NAND2_X1 U13981 ( .A1(n11442), .A2(n11441), .ZN(n11448) );
  INV_X1 U13982 ( .A(n11443), .ZN(n11446) );
  INV_X1 U13983 ( .A(n11444), .ZN(n11445) );
  NAND2_X1 U13984 ( .A1(n11446), .A2(n11445), .ZN(n11447) );
  NAND2_X1 U13985 ( .A1(n11448), .A2(n11447), .ZN(n11450) );
  MUX2_X1 U13986 ( .A(n14520), .B(n14768), .S(n11609), .Z(n11451) );
  MUX2_X1 U13987 ( .A(n14520), .B(n14768), .S(n6443), .Z(n11449) );
  MUX2_X1 U13988 ( .A(n14404), .B(n6612), .S(n6443), .Z(n11455) );
  MUX2_X1 U13989 ( .A(n14404), .B(n6612), .S(n11422), .Z(n11452) );
  NAND2_X1 U13990 ( .A1(n11453), .A2(n11452), .ZN(n11456) );
  MUX2_X1 U13991 ( .A(n14519), .B(n13712), .S(n11609), .Z(n11458) );
  MUX2_X1 U13992 ( .A(n14519), .B(n13712), .S(n6443), .Z(n11457) );
  MUX2_X1 U13993 ( .A(n14558), .B(n14570), .S(n6443), .Z(n11462) );
  NAND2_X1 U13994 ( .A1(n11461), .A2(n11462), .ZN(n11460) );
  MUX2_X1 U13995 ( .A(n14558), .B(n14570), .S(n11422), .Z(n11459) );
  NAND2_X1 U13996 ( .A1(n11460), .A2(n11459), .ZN(n11466) );
  INV_X1 U13997 ( .A(n11462), .ZN(n11463) );
  NAND2_X1 U13998 ( .A1(n11464), .A2(n11463), .ZN(n11465) );
  NAND2_X1 U13999 ( .A1(n11472), .A2(n11467), .ZN(n11470) );
  NAND2_X1 U14000 ( .A1(n11471), .A2(n11468), .ZN(n11469) );
  MUX2_X1 U14001 ( .A(n11470), .B(n11469), .S(n6443), .Z(n11474) );
  MUX2_X1 U14002 ( .A(n11472), .B(n11471), .S(n11609), .Z(n11473) );
  MUX2_X1 U14003 ( .A(n14547), .B(n14227), .S(n6443), .Z(n11490) );
  NAND2_X1 U14004 ( .A1(n11490), .A2(n14093), .ZN(n11475) );
  NAND2_X1 U14005 ( .A1(n13802), .A2(n6443), .ZN(n11487) );
  AOI21_X1 U14006 ( .B1(n11475), .B2(n11487), .A(n14221), .ZN(n11480) );
  INV_X1 U14007 ( .A(n14093), .ZN(n14210) );
  NAND2_X1 U14008 ( .A1(n11490), .A2(n14210), .ZN(n11476) );
  OR2_X1 U14009 ( .A1(n14227), .A2(n6443), .ZN(n11481) );
  AOI21_X1 U14010 ( .B1(n11476), .B2(n11481), .A(n11492), .ZN(n11479) );
  NAND2_X1 U14011 ( .A1(n14093), .A2(n11609), .ZN(n11483) );
  OR2_X1 U14012 ( .A1(n14227), .A2(n11483), .ZN(n11478) );
  NOR2_X1 U14013 ( .A1(n14093), .A2(n11609), .ZN(n11488) );
  NAND2_X1 U14014 ( .A1(n11488), .A2(n13802), .ZN(n11477) );
  NAND2_X1 U14015 ( .A1(n11478), .A2(n11477), .ZN(n11485) );
  INV_X1 U14016 ( .A(n11481), .ZN(n11482) );
  NAND2_X1 U14017 ( .A1(n11490), .A2(n11482), .ZN(n11484) );
  NAND2_X1 U14018 ( .A1(n11484), .A2(n11483), .ZN(n11486) );
  AOI22_X1 U14019 ( .A1(n11486), .A2(n14221), .B1(n11490), .B2(n11485), .ZN(
        n11495) );
  INV_X1 U14020 ( .A(n11487), .ZN(n11489) );
  AOI21_X1 U14021 ( .B1(n11490), .B2(n11489), .A(n11488), .ZN(n11491) );
  INV_X1 U14022 ( .A(n11491), .ZN(n11493) );
  OR2_X1 U14023 ( .A1(n11496), .A2(n11654), .ZN(n11498) );
  AOI22_X1 U14024 ( .A1(n11502), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11501), 
        .B2(n13851), .ZN(n11497) );
  INV_X1 U14025 ( .A(n14202), .ZN(n14218) );
  OR2_X1 U14026 ( .A1(n14214), .A2(n14218), .ZN(n13882) );
  MUX2_X1 U14027 ( .A(n14202), .B(n14097), .S(n11422), .Z(n11499) );
  AND2_X1 U14028 ( .A1(n14214), .A2(n14218), .ZN(n13881) );
  NAND2_X1 U14029 ( .A1(n11500), .A2(n11641), .ZN(n11504) );
  AOI22_X1 U14030 ( .A1(n11502), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n11703), 
        .B2(n11501), .ZN(n11503) );
  XNOR2_X1 U14031 ( .A(n11517), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n14074) );
  NAND2_X1 U14032 ( .A1(n14074), .A2(n11646), .ZN(n11509) );
  INV_X1 U14033 ( .A(n11614), .ZN(n11662) );
  INV_X1 U14034 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13849) );
  NAND2_X1 U14035 ( .A1(n11657), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11506) );
  NAND2_X1 U14036 ( .A1(n11599), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11505) );
  OAI211_X1 U14037 ( .C1(n11662), .C2(n13849), .A(n11506), .B(n11505), .ZN(
        n11507) );
  INV_X1 U14038 ( .A(n11507), .ZN(n11508) );
  XNOR2_X1 U14039 ( .A(n14205), .B(n14211), .ZN(n14078) );
  INV_X1 U14040 ( .A(n14211), .ZN(n14193) );
  NAND2_X1 U14041 ( .A1(n14193), .A2(n6443), .ZN(n11511) );
  OR2_X1 U14042 ( .A1(n14193), .A2(n6443), .ZN(n11510) );
  MUX2_X1 U14043 ( .A(n11511), .B(n11510), .S(n14205), .Z(n11512) );
  NAND2_X1 U14044 ( .A1(n11513), .A2(n11512), .ZN(n11524) );
  OR2_X1 U14045 ( .A1(n11514), .A2(n11654), .ZN(n11516) );
  OR2_X1 U14046 ( .A1(n11655), .A2(n15142), .ZN(n11515) );
  INV_X1 U14047 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n13695) );
  INV_X1 U14048 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13760) );
  OAI21_X1 U14049 ( .B1(n11517), .B2(n13695), .A(n13760), .ZN(n11518) );
  AND2_X1 U14050 ( .A1(n11518), .A2(n11531), .ZN(n14060) );
  NAND2_X1 U14051 ( .A1(n14060), .A2(n11646), .ZN(n11521) );
  AOI22_X1 U14052 ( .A1(n9899), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n11599), 
        .B2(P1_REG0_REG_20__SCAN_IN), .ZN(n11520) );
  NAND2_X1 U14053 ( .A1(n11657), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n11519) );
  MUX2_X1 U14054 ( .A(n14197), .B(n14203), .S(n11422), .Z(n11523) );
  INV_X1 U14055 ( .A(n14203), .ZN(n13899) );
  MUX2_X1 U14056 ( .A(n13899), .B(n14069), .S(n11422), .Z(n11522) );
  OAI21_X1 U14057 ( .B1(n11524), .B2(n11523), .A(n11522), .ZN(n11526) );
  NAND2_X1 U14058 ( .A1(n11524), .A2(n11523), .ZN(n11525) );
  NAND2_X1 U14059 ( .A1(n11526), .A2(n11525), .ZN(n11539) );
  OR2_X1 U14060 ( .A1(n11527), .A2(n11654), .ZN(n11530) );
  OR2_X1 U14061 ( .A1(n11655), .A2(n11528), .ZN(n11529) );
  INV_X1 U14062 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n15206) );
  AND2_X1 U14063 ( .A1(n11531), .A2(n15206), .ZN(n11532) );
  OR2_X1 U14064 ( .A1(n11532), .A2(n11546), .ZN(n14043) );
  INV_X1 U14065 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n11535) );
  NAND2_X1 U14066 ( .A1(n11599), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11534) );
  NAND2_X1 U14067 ( .A1(n11657), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n11533) );
  OAI211_X1 U14068 ( .C1(n11662), .C2(n11535), .A(n11534), .B(n11533), .ZN(
        n11536) );
  INV_X1 U14069 ( .A(n11536), .ZN(n11537) );
  OAI21_X1 U14070 ( .B1(n14043), .B2(n11553), .A(n11537), .ZN(n14194) );
  MUX2_X1 U14071 ( .A(n14187), .B(n14194), .S(n6443), .Z(n11540) );
  MUX2_X1 U14072 ( .A(n14187), .B(n14194), .S(n11422), .Z(n11538) );
  INV_X1 U14073 ( .A(n11540), .ZN(n11541) );
  NOR2_X1 U14074 ( .A1(n11546), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11547) );
  OR2_X1 U14075 ( .A1(n11562), .A2(n11547), .ZN(n14032) );
  INV_X1 U14076 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n11550) );
  NAND2_X1 U14077 ( .A1(n11599), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11549) );
  NAND2_X1 U14078 ( .A1(n11657), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n11548) );
  OAI211_X1 U14079 ( .C1(n11550), .C2(n11662), .A(n11549), .B(n11548), .ZN(
        n11551) );
  INV_X1 U14080 ( .A(n11551), .ZN(n11552) );
  OAI21_X1 U14081 ( .B1(n14032), .B2(n11553), .A(n11552), .ZN(n14047) );
  NAND2_X1 U14082 ( .A1(n11556), .A2(n11557), .ZN(n11555) );
  MUX2_X1 U14083 ( .A(n14180), .B(n14047), .S(n6443), .Z(n11554) );
  NAND2_X1 U14084 ( .A1(n11555), .A2(n11554), .ZN(n11561) );
  INV_X1 U14085 ( .A(n11557), .ZN(n11558) );
  NAND2_X1 U14086 ( .A1(n11559), .A2(n11558), .ZN(n11560) );
  OR2_X1 U14087 ( .A1(n11562), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11563) );
  NAND2_X1 U14088 ( .A1(n11562), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11576) );
  AND2_X1 U14089 ( .A1(n11563), .A2(n11576), .ZN(n13686) );
  NAND2_X1 U14090 ( .A1(n13686), .A2(n11646), .ZN(n11569) );
  INV_X1 U14091 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n11566) );
  NAND2_X1 U14092 ( .A1(n11599), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n11565) );
  NAND2_X1 U14093 ( .A1(n11657), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n11564) );
  OAI211_X1 U14094 ( .C1(n11662), .C2(n11566), .A(n11565), .B(n11564), .ZN(
        n11567) );
  INV_X1 U14095 ( .A(n11567), .ZN(n11568) );
  NAND2_X1 U14096 ( .A1(n11569), .A2(n11568), .ZN(n13888) );
  NAND2_X1 U14097 ( .A1(n14273), .A2(n11641), .ZN(n11571) );
  INV_X1 U14098 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n14277) );
  OR2_X1 U14099 ( .A1(n11655), .A2(n14277), .ZN(n11570) );
  MUX2_X1 U14100 ( .A(n13888), .B(n14175), .S(n11422), .Z(n11573) );
  MUX2_X1 U14101 ( .A(n13888), .B(n14175), .S(n6443), .Z(n11572) );
  INV_X1 U14102 ( .A(n11573), .ZN(n11574) );
  NAND2_X1 U14103 ( .A1(n11614), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n11580) );
  NAND2_X1 U14104 ( .A1(n11599), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11579) );
  INV_X1 U14105 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13751) );
  INV_X1 U14106 ( .A(n11576), .ZN(n11575) );
  NAND2_X1 U14107 ( .A1(n11575), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n11589) );
  AOI21_X1 U14108 ( .B1(n13751), .B2(n11576), .A(n11588), .ZN(n14001) );
  NAND2_X1 U14109 ( .A1(n11646), .A2(n14001), .ZN(n11578) );
  NAND2_X1 U14110 ( .A1(n11657), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n11577) );
  NAND4_X1 U14111 ( .A1(n11580), .A2(n11579), .A3(n11578), .A4(n11577), .ZN(
        n14154) );
  OR2_X1 U14112 ( .A1(n11655), .A2(n11582), .ZN(n11583) );
  MUX2_X1 U14113 ( .A(n14154), .B(n14170), .S(n6443), .Z(n11586) );
  MUX2_X1 U14114 ( .A(n14170), .B(n14154), .S(n6443), .Z(n11585) );
  INV_X1 U14115 ( .A(n11586), .ZN(n11587) );
  NAND2_X1 U14116 ( .A1(n11614), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n11593) );
  NAND2_X1 U14117 ( .A1(n11599), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n11592) );
  INV_X1 U14118 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13720) );
  NAND2_X1 U14119 ( .A1(n11588), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n11600) );
  INV_X1 U14120 ( .A(n11600), .ZN(n11601) );
  AOI21_X1 U14121 ( .B1(n13720), .B2(n11589), .A(n11601), .ZN(n13984) );
  NAND2_X1 U14122 ( .A1(n11646), .A2(n13984), .ZN(n11591) );
  NAND2_X1 U14123 ( .A1(n11657), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n11590) );
  NAND4_X1 U14124 ( .A1(n11593), .A2(n11592), .A3(n11591), .A4(n11590), .ZN(
        n14004) );
  NAND2_X1 U14125 ( .A1(n13664), .A2(n11641), .ZN(n11595) );
  OR2_X1 U14126 ( .A1(n11655), .A2(n14271), .ZN(n11594) );
  MUX2_X1 U14127 ( .A(n14004), .B(n13983), .S(n11422), .Z(n11598) );
  MUX2_X1 U14128 ( .A(n14004), .B(n13983), .S(n6443), .Z(n11596) );
  NAND2_X1 U14129 ( .A1(n11599), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n11606) );
  NAND2_X1 U14130 ( .A1(n11614), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n11605) );
  INV_X1 U14131 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13785) );
  NAND2_X1 U14132 ( .A1(n13785), .A2(n11600), .ZN(n11602) );
  NAND2_X1 U14133 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n11601), .ZN(n11616) );
  AND2_X1 U14134 ( .A1(n11602), .A2(n11616), .ZN(n13786) );
  NAND2_X1 U14135 ( .A1(n11646), .A2(n13786), .ZN(n11604) );
  NAND2_X1 U14136 ( .A1(n11657), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n11603) );
  NAND4_X1 U14137 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n14155) );
  NAND2_X1 U14138 ( .A1(n13661), .A2(n11641), .ZN(n11608) );
  OR2_X1 U14139 ( .A1(n11655), .A2(n14265), .ZN(n11607) );
  MUX2_X1 U14140 ( .A(n14155), .B(n14150), .S(n6443), .Z(n11611) );
  MUX2_X1 U14141 ( .A(n14155), .B(n14150), .S(n11609), .Z(n11610) );
  OR2_X1 U14142 ( .A1(n11655), .A2(n11612), .ZN(n11613) );
  NAND2_X1 U14143 ( .A1(n11614), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n11621) );
  NAND2_X1 U14144 ( .A1(n11599), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n11620) );
  INV_X1 U14145 ( .A(n11616), .ZN(n11615) );
  NAND2_X1 U14146 ( .A1(n11615), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n11627) );
  INV_X1 U14147 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13677) );
  NAND2_X1 U14148 ( .A1(n11616), .A2(n13677), .ZN(n11617) );
  NAND2_X1 U14149 ( .A1(n10112), .A2(n13948), .ZN(n11619) );
  NAND2_X1 U14150 ( .A1(n11657), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n11618) );
  NAND4_X1 U14151 ( .A1(n11621), .A2(n11620), .A3(n11619), .A4(n11618), .ZN(
        n13967) );
  MUX2_X1 U14152 ( .A(n13967), .B(n14142), .S(n6443), .Z(n11622) );
  INV_X1 U14153 ( .A(n11624), .ZN(n11625) );
  INV_X1 U14154 ( .A(n11637), .ZN(n11636) );
  NAND2_X1 U14155 ( .A1(n9899), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n11632) );
  NAND2_X1 U14156 ( .A1(n11599), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n11631) );
  INV_X1 U14157 ( .A(n11627), .ZN(n11626) );
  NAND2_X1 U14158 ( .A1(n11626), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13916) );
  INV_X1 U14159 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n11873) );
  NAND2_X1 U14160 ( .A1(n11627), .A2(n11873), .ZN(n11628) );
  NAND2_X1 U14161 ( .A1(n11646), .A2(n11874), .ZN(n11630) );
  NAND2_X1 U14162 ( .A1(n11657), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n11629) );
  NAND2_X1 U14163 ( .A1(n14261), .A2(n11641), .ZN(n11634) );
  OR2_X1 U14164 ( .A1(n11655), .A2(n14264), .ZN(n11633) );
  MUX2_X1 U14165 ( .A(n14138), .B(n14132), .S(n6443), .Z(n11638) );
  MUX2_X1 U14166 ( .A(n13937), .B(n14120), .S(n6443), .Z(n11635) );
  OAI21_X1 U14167 ( .B1(n11636), .B2(n11638), .A(n11635), .ZN(n11640) );
  NAND2_X1 U14168 ( .A1(n11636), .A2(n11638), .ZN(n11639) );
  NAND2_X1 U14169 ( .A1(n11642), .A2(n11641), .ZN(n11644) );
  OR2_X1 U14170 ( .A1(n11655), .A2(n14260), .ZN(n11643) );
  NAND2_X1 U14171 ( .A1(n11614), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n11650) );
  NAND2_X1 U14172 ( .A1(n11599), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n11649) );
  INV_X1 U14173 ( .A(n13916), .ZN(n11645) );
  NAND2_X1 U14174 ( .A1(n11646), .A2(n11645), .ZN(n11648) );
  NAND2_X1 U14175 ( .A1(n11657), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n11647) );
  NAND4_X1 U14176 ( .A1(n11650), .A2(n11649), .A3(n11648), .A4(n11647), .ZN(
        n13928) );
  MUX2_X1 U14177 ( .A(n13909), .B(n13928), .S(n6443), .Z(n11669) );
  INV_X1 U14178 ( .A(n11651), .ZN(n11652) );
  INV_X1 U14179 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15172) );
  INV_X1 U14180 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n11661) );
  NAND2_X1 U14181 ( .A1(n11657), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n11660) );
  NAND2_X1 U14182 ( .A1(n11599), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n11659) );
  OAI211_X1 U14183 ( .C1(n11662), .C2(n11661), .A(n11660), .B(n11659), .ZN(
        n13912) );
  OAI22_X1 U14184 ( .A1(n13870), .A2(n6443), .B1(n9609), .B2(n11663), .ZN(
        n11664) );
  AOI22_X1 U14185 ( .A1(n13866), .A2(n6443), .B1(n13912), .B2(n11664), .ZN(
        n11670) );
  OAI21_X1 U14186 ( .B1(n13807), .B2(n11665), .A(n13912), .ZN(n11666) );
  MUX2_X1 U14187 ( .A(n14118), .B(n11666), .S(n6443), .Z(n11671) );
  INV_X1 U14188 ( .A(n11671), .ZN(n11667) );
  INV_X1 U14189 ( .A(n13928), .ZN(n11875) );
  INV_X1 U14190 ( .A(n13909), .ZN(n14123) );
  MUX2_X1 U14191 ( .A(n11875), .B(n14123), .S(n6443), .Z(n11668) );
  INV_X1 U14192 ( .A(n11670), .ZN(n11672) );
  XNOR2_X1 U14193 ( .A(n14150), .B(n14139), .ZN(n13971) );
  XNOR2_X1 U14194 ( .A(n13983), .B(n14166), .ZN(n13979) );
  XNOR2_X1 U14195 ( .A(n14170), .B(n14154), .ZN(n13997) );
  INV_X1 U14196 ( .A(n14047), .ZN(n14184) );
  INV_X1 U14197 ( .A(n14194), .ZN(n13770) );
  NAND2_X1 U14198 ( .A1(n14049), .A2(n13770), .ZN(n13885) );
  NAND2_X1 U14199 ( .A1(n14187), .A2(n14194), .ZN(n11673) );
  XNOR2_X1 U14200 ( .A(n14069), .B(n14203), .ZN(n14058) );
  NAND2_X1 U14201 ( .A1(n14214), .A2(n14202), .ZN(n11674) );
  NOR4_X1 U14202 ( .A1(n11677), .A2(n14698), .A3(n11676), .A4(n11675), .ZN(
        n11681) );
  NAND4_X1 U14203 ( .A1(n11679), .A2(n11680), .A3(n11681), .A4(n11678), .ZN(
        n11683) );
  NOR4_X1 U14204 ( .A1(n11684), .A2(n11683), .A3(n14677), .A4(n11682), .ZN(
        n11686) );
  NAND4_X1 U14205 ( .A1(n11687), .A2(n11686), .A3(n14532), .A4(n11685), .ZN(
        n11688) );
  NOR4_X1 U14206 ( .A1(n11690), .A2(n11689), .A3(n14433), .A4(n11688), .ZN(
        n11693) );
  NAND4_X1 U14207 ( .A1(n14099), .A2(n11693), .A3(n11692), .A4(n11691), .ZN(
        n11694) );
  NOR4_X1 U14208 ( .A1(n13884), .A2(n14078), .A3(n14058), .A4(n11694), .ZN(
        n11695) );
  XNOR2_X1 U14209 ( .A(n14175), .B(n13888), .ZN(n14012) );
  NAND4_X1 U14210 ( .A1(n13997), .A2(n6630), .A3(n11695), .A4(n14012), .ZN(
        n11696) );
  NOR4_X1 U14211 ( .A1(n13908), .A2(n13971), .A3(n13979), .A4(n11696), .ZN(
        n11701) );
  NOR2_X1 U14212 ( .A1(n11697), .A2(n7365), .ZN(n11700) );
  XNOR2_X1 U14213 ( .A(n13867), .B(n13870), .ZN(n11714) );
  INV_X1 U14214 ( .A(n11714), .ZN(n11699) );
  NAND2_X1 U14215 ( .A1(n13937), .A2(n14120), .ZN(n13893) );
  NAND4_X1 U14216 ( .A1(n11701), .A2(n11700), .A3(n11699), .A4(n13932), .ZN(
        n11702) );
  NOR3_X1 U14217 ( .A1(n14115), .A2(n13807), .A3(n11704), .ZN(n11707) );
  NOR3_X1 U14218 ( .A1(n11706), .A2(n13807), .A3(n11713), .ZN(n11705) );
  AOI21_X1 U14219 ( .B1(n11707), .B2(n11706), .A(n11705), .ZN(n11711) );
  XOR2_X1 U14220 ( .A(n11713), .B(n11708), .Z(n11709) );
  NAND4_X1 U14221 ( .A1(n11709), .A2(n14115), .A3(n13807), .A4(n11712), .ZN(
        n11710) );
  OAI211_X1 U14222 ( .C1(n7447), .C2(n11712), .A(n11711), .B(n11710), .ZN(
        n11716) );
  AOI211_X1 U14223 ( .C1(n11718), .C2(n11717), .A(n11716), .B(n11715), .ZN(
        n11723) );
  NAND3_X1 U14224 ( .A1(n11720), .A2(n11719), .A3(n14766), .ZN(n11721) );
  OAI211_X1 U14225 ( .C1(n14279), .C2(n14274), .A(n11721), .B(P1_B_REG_SCAN_IN), .ZN(n11722) );
  OAI21_X1 U14226 ( .B1(n11723), .B2(n14274), .A(n11722), .ZN(P1_U3242) );
  OAI22_X1 U14227 ( .A1(n13490), .A2(n11725), .B1(n11724), .B2(n13487), .ZN(
        n11728) );
  NOR2_X1 U14228 ( .A1(n11726), .A2(n13410), .ZN(n11727) );
  AOI211_X1 U14229 ( .C1(n13493), .C2(n12037), .A(n11728), .B(n11727), .ZN(
        n11731) );
  OR2_X1 U14230 ( .A1(n11729), .A2(n15079), .ZN(n11730) );
  OAI211_X1 U14231 ( .C1(n11732), .C2(n13474), .A(n11731), .B(n11730), .ZN(
        P2_U3236) );
  INV_X1 U14232 ( .A(SI_30_), .ZN(n12283) );
  NAND2_X1 U14233 ( .A1(n14260), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11733) );
  NAND2_X1 U14234 ( .A1(n15172), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12273) );
  INV_X1 U14235 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12138) );
  NAND2_X1 U14236 ( .A1(n12138), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n11735) );
  AND2_X1 U14237 ( .A1(n12273), .A2(n11735), .ZN(n11736) );
  NAND2_X1 U14238 ( .A1(n11737), .A2(n11736), .ZN(n12274) );
  OAI21_X1 U14239 ( .B1(n11737), .B2(n11736), .A(n12274), .ZN(n12282) );
  OAI222_X1 U14240 ( .A1(n11738), .A2(P3_U3151), .B1(n12995), .B2(n12283), 
        .C1(n12997), .C2(n12282), .ZN(P3_U3265) );
  INV_X1 U14241 ( .A(n11739), .ZN(n11741) );
  AOI22_X1 U14242 ( .A1(n6612), .A2(n11801), .B1(n11863), .B2(n14404), .ZN(
        n11747) );
  NAND2_X1 U14243 ( .A1(n14538), .A2(n11858), .ZN(n11745) );
  NAND2_X1 U14244 ( .A1(n14404), .A2(n11801), .ZN(n11744) );
  NAND2_X1 U14245 ( .A1(n11745), .A2(n11744), .ZN(n11746) );
  XNOR2_X1 U14246 ( .A(n11746), .B(n11861), .ZN(n11749) );
  XOR2_X1 U14247 ( .A(n11747), .B(n11749), .Z(n14523) );
  INV_X1 U14248 ( .A(n11747), .ZN(n11748) );
  AND2_X1 U14249 ( .A1(n11863), .A2(n14519), .ZN(n11750) );
  AOI21_X1 U14250 ( .B1(n13712), .B2(n11801), .A(n11750), .ZN(n11759) );
  NAND2_X1 U14251 ( .A1(n13712), .A2(n11858), .ZN(n11752) );
  NAND2_X1 U14252 ( .A1(n14519), .A2(n11801), .ZN(n11751) );
  NAND2_X1 U14253 ( .A1(n11752), .A2(n11751), .ZN(n11753) );
  XNOR2_X1 U14254 ( .A(n11753), .B(n11861), .ZN(n11761) );
  XOR2_X1 U14255 ( .A(n11759), .B(n11761), .Z(n13711) );
  INV_X1 U14256 ( .A(n13711), .ZN(n11754) );
  NAND2_X1 U14257 ( .A1(n14570), .A2(n11858), .ZN(n11756) );
  NAND2_X1 U14258 ( .A1(n14558), .A2(n11801), .ZN(n11755) );
  NAND2_X1 U14259 ( .A1(n11756), .A2(n11755), .ZN(n11757) );
  INV_X2 U14260 ( .A(n6452), .ZN(n11861) );
  XNOR2_X1 U14261 ( .A(n11757), .B(n11861), .ZN(n11763) );
  AND2_X1 U14262 ( .A1(n11863), .A2(n14558), .ZN(n11758) );
  AOI21_X1 U14263 ( .B1(n14570), .B2(n11801), .A(n11758), .ZN(n11764) );
  XNOR2_X1 U14264 ( .A(n11763), .B(n11764), .ZN(n14513) );
  INV_X1 U14265 ( .A(n11759), .ZN(n11760) );
  NAND2_X1 U14266 ( .A1(n11761), .A2(n11760), .ZN(n14511) );
  NAND2_X1 U14267 ( .A1(n13708), .A2(n11762), .ZN(n14512) );
  INV_X1 U14268 ( .A(n11763), .ZN(n11765) );
  NAND2_X1 U14269 ( .A1(n11765), .A2(n11764), .ZN(n11766) );
  NAND2_X1 U14270 ( .A1(n14512), .A2(n11766), .ZN(n14498) );
  INV_X1 U14271 ( .A(n11767), .ZN(n14562) );
  OAI22_X1 U14272 ( .A1(n14562), .A2(n11867), .B1(n14421), .B2(n9799), .ZN(
        n11775) );
  NAND2_X1 U14273 ( .A1(n11767), .A2(n11858), .ZN(n11769) );
  OR2_X1 U14274 ( .A1(n14421), .A2(n11867), .ZN(n11768) );
  NAND2_X1 U14275 ( .A1(n11769), .A2(n11768), .ZN(n11770) );
  XNOR2_X1 U14276 ( .A(n11770), .B(n11861), .ZN(n11776) );
  XOR2_X1 U14277 ( .A(n11775), .B(n11776), .Z(n14499) );
  NAND2_X1 U14278 ( .A1(n14498), .A2(n14499), .ZN(n13793) );
  NAND2_X1 U14279 ( .A1(n13804), .A2(n11858), .ZN(n11772) );
  OR2_X1 U14280 ( .A1(n14501), .A2(n11867), .ZN(n11771) );
  NAND2_X1 U14281 ( .A1(n11772), .A2(n11771), .ZN(n11773) );
  XNOR2_X1 U14282 ( .A(n11773), .B(n6452), .ZN(n13795) );
  NOR2_X1 U14283 ( .A1(n14501), .A2(n9799), .ZN(n11774) );
  AOI21_X1 U14284 ( .B1(n13804), .B2(n11801), .A(n11774), .ZN(n13794) );
  NOR2_X1 U14285 ( .A1(n11776), .A2(n11775), .ZN(n13791) );
  AOI21_X1 U14286 ( .B1(n13795), .B2(n13794), .A(n13791), .ZN(n11777) );
  INV_X1 U14287 ( .A(n13795), .ZN(n11779) );
  INV_X1 U14288 ( .A(n13794), .ZN(n11778) );
  NAND2_X1 U14289 ( .A1(n11779), .A2(n11778), .ZN(n11780) );
  AOI22_X1 U14290 ( .A1(n14227), .A2(n11858), .B1(n11801), .B2(n14547), .ZN(
        n11781) );
  XNOR2_X1 U14291 ( .A(n11781), .B(n11861), .ZN(n11784) );
  AOI22_X1 U14292 ( .A1(n14227), .A2(n11801), .B1(n11863), .B2(n14547), .ZN(
        n11783) );
  XNOR2_X1 U14293 ( .A(n11784), .B(n11783), .ZN(n13729) );
  NAND2_X1 U14294 ( .A1(n11784), .A2(n11783), .ZN(n11785) );
  NAND2_X1 U14295 ( .A1(n13727), .A2(n11785), .ZN(n13739) );
  OR2_X1 U14296 ( .A1(n14221), .A2(n11867), .ZN(n11787) );
  NAND2_X1 U14297 ( .A1(n14093), .A2(n11863), .ZN(n11786) );
  NAND2_X1 U14298 ( .A1(n11787), .A2(n11786), .ZN(n11790) );
  OAI22_X1 U14299 ( .A1(n14221), .A2(n10169), .B1(n14210), .B2(n11867), .ZN(
        n11788) );
  XNOR2_X1 U14300 ( .A(n11788), .B(n11861), .ZN(n11789) );
  XOR2_X1 U14301 ( .A(n11790), .B(n11789), .Z(n13740) );
  NAND2_X1 U14302 ( .A1(n13739), .A2(n13740), .ZN(n13738) );
  INV_X1 U14303 ( .A(n11789), .ZN(n11792) );
  INV_X1 U14304 ( .A(n11790), .ZN(n11791) );
  NAND2_X1 U14305 ( .A1(n11792), .A2(n11791), .ZN(n11793) );
  NAND2_X1 U14306 ( .A1(n13738), .A2(n11793), .ZN(n13777) );
  OAI22_X1 U14307 ( .A1(n14097), .A2(n11867), .B1(n14202), .B2(n9799), .ZN(
        n11796) );
  OAI22_X1 U14308 ( .A1(n14097), .A2(n10169), .B1(n14202), .B2(n11867), .ZN(
        n11794) );
  XNOR2_X1 U14309 ( .A(n11794), .B(n11861), .ZN(n11795) );
  XOR2_X1 U14310 ( .A(n11796), .B(n11795), .Z(n13776) );
  INV_X1 U14311 ( .A(n11795), .ZN(n11798) );
  INV_X1 U14312 ( .A(n11796), .ZN(n11797) );
  NAND2_X1 U14313 ( .A1(n11798), .A2(n11797), .ZN(n11799) );
  NOR2_X1 U14314 ( .A1(n14211), .A2(n9799), .ZN(n11800) );
  AOI21_X1 U14315 ( .B1(n14205), .B2(n11801), .A(n11800), .ZN(n11806) );
  NAND2_X1 U14316 ( .A1(n14205), .A2(n11858), .ZN(n11803) );
  OR2_X1 U14317 ( .A1(n14211), .A2(n11867), .ZN(n11802) );
  NAND2_X1 U14318 ( .A1(n11803), .A2(n11802), .ZN(n11804) );
  XNOR2_X1 U14319 ( .A(n11804), .B(n11861), .ZN(n11805) );
  XOR2_X1 U14320 ( .A(n11806), .B(n11805), .Z(n13691) );
  INV_X1 U14321 ( .A(n11805), .ZN(n11807) );
  OR2_X1 U14322 ( .A1(n11807), .A2(n11806), .ZN(n11808) );
  NAND2_X1 U14323 ( .A1(n13693), .A2(n11808), .ZN(n13759) );
  OAI22_X1 U14324 ( .A1(n14197), .A2(n11867), .B1(n14203), .B2(n9799), .ZN(
        n11810) );
  OAI22_X1 U14325 ( .A1(n14197), .A2(n10169), .B1(n14203), .B2(n11867), .ZN(
        n11809) );
  XNOR2_X1 U14326 ( .A(n11809), .B(n11861), .ZN(n11811) );
  XOR2_X1 U14327 ( .A(n11810), .B(n11811), .Z(n13758) );
  NAND2_X1 U14328 ( .A1(n11811), .A2(n11810), .ZN(n11812) );
  OAI22_X1 U14329 ( .A1(n14049), .A2(n10169), .B1(n13770), .B2(n11867), .ZN(
        n11813) );
  XNOR2_X1 U14330 ( .A(n11813), .B(n11861), .ZN(n11815) );
  OAI22_X1 U14331 ( .A1(n14049), .A2(n11867), .B1(n13770), .B2(n9799), .ZN(
        n11816) );
  XNOR2_X1 U14332 ( .A(n11815), .B(n11816), .ZN(n13703) );
  INV_X1 U14333 ( .A(n13703), .ZN(n11814) );
  INV_X1 U14334 ( .A(n11815), .ZN(n11818) );
  INV_X1 U14335 ( .A(n11816), .ZN(n11817) );
  NAND2_X1 U14336 ( .A1(n11818), .A2(n11817), .ZN(n11819) );
  NAND2_X1 U14337 ( .A1(n13700), .A2(n11819), .ZN(n13767) );
  OAI22_X1 U14338 ( .A1(n13775), .A2(n11867), .B1(n14184), .B2(n9799), .ZN(
        n11824) );
  NAND2_X1 U14339 ( .A1(n14180), .A2(n11858), .ZN(n11821) );
  NAND2_X1 U14340 ( .A1(n14047), .A2(n11801), .ZN(n11820) );
  NAND2_X1 U14341 ( .A1(n11821), .A2(n11820), .ZN(n11822) );
  XNOR2_X1 U14342 ( .A(n11822), .B(n11861), .ZN(n11823) );
  XOR2_X1 U14343 ( .A(n11824), .B(n11823), .Z(n13768) );
  INV_X1 U14344 ( .A(n11823), .ZN(n11826) );
  INV_X1 U14345 ( .A(n11824), .ZN(n11825) );
  NAND2_X1 U14346 ( .A1(n11826), .A2(n11825), .ZN(n11827) );
  NAND2_X1 U14347 ( .A1(n14175), .A2(n11858), .ZN(n11829) );
  NAND2_X1 U14348 ( .A1(n13888), .A2(n11801), .ZN(n11828) );
  NAND2_X1 U14349 ( .A1(n11829), .A2(n11828), .ZN(n11830) );
  XNOR2_X1 U14350 ( .A(n11830), .B(n11861), .ZN(n11831) );
  AOI22_X1 U14351 ( .A1(n14175), .A2(n11801), .B1(n11863), .B2(n13888), .ZN(
        n11832) );
  XNOR2_X1 U14352 ( .A(n11831), .B(n11832), .ZN(n13683) );
  INV_X1 U14353 ( .A(n11831), .ZN(n11833) );
  NAND2_X1 U14354 ( .A1(n14170), .A2(n11858), .ZN(n11835) );
  NAND2_X1 U14355 ( .A1(n14154), .A2(n11801), .ZN(n11834) );
  NAND2_X1 U14356 ( .A1(n11835), .A2(n11834), .ZN(n11836) );
  XNOR2_X1 U14357 ( .A(n11836), .B(n11861), .ZN(n11837) );
  AOI22_X1 U14358 ( .A1(n14170), .A2(n11801), .B1(n11863), .B2(n14154), .ZN(
        n11838) );
  NAND2_X1 U14359 ( .A1(n13749), .A2(n13750), .ZN(n11841) );
  INV_X1 U14360 ( .A(n11837), .ZN(n11839) );
  NAND2_X1 U14361 ( .A1(n11839), .A2(n11838), .ZN(n11840) );
  NAND2_X1 U14362 ( .A1(n11841), .A2(n11840), .ZN(n13718) );
  NAND2_X1 U14363 ( .A1(n13983), .A2(n11858), .ZN(n11843) );
  NAND2_X1 U14364 ( .A1(n14004), .A2(n11801), .ZN(n11842) );
  NAND2_X1 U14365 ( .A1(n11843), .A2(n11842), .ZN(n11844) );
  XNOR2_X1 U14366 ( .A(n11844), .B(n11861), .ZN(n11845) );
  AOI22_X1 U14367 ( .A1(n13983), .A2(n11801), .B1(n11863), .B2(n14004), .ZN(
        n11846) );
  XNOR2_X1 U14368 ( .A(n11845), .B(n11846), .ZN(n13719) );
  NAND2_X1 U14369 ( .A1(n13718), .A2(n13719), .ZN(n11849) );
  INV_X1 U14370 ( .A(n11845), .ZN(n11847) );
  NAND2_X1 U14371 ( .A1(n11847), .A2(n11846), .ZN(n11848) );
  NAND2_X1 U14372 ( .A1(n11849), .A2(n11848), .ZN(n13783) );
  NAND2_X1 U14373 ( .A1(n14150), .A2(n11858), .ZN(n11851) );
  NAND2_X1 U14374 ( .A1(n14155), .A2(n11801), .ZN(n11850) );
  NAND2_X1 U14375 ( .A1(n11851), .A2(n11850), .ZN(n11852) );
  XNOR2_X1 U14376 ( .A(n11852), .B(n11861), .ZN(n11853) );
  AOI22_X1 U14377 ( .A1(n14150), .A2(n11801), .B1(n11863), .B2(n14155), .ZN(
        n11854) );
  XNOR2_X1 U14378 ( .A(n11853), .B(n11854), .ZN(n13784) );
  NAND2_X1 U14379 ( .A1(n13783), .A2(n13784), .ZN(n11857) );
  INV_X1 U14380 ( .A(n11853), .ZN(n11855) );
  NAND2_X1 U14381 ( .A1(n11855), .A2(n11854), .ZN(n11856) );
  NAND2_X1 U14382 ( .A1(n14142), .A2(n11858), .ZN(n11860) );
  NAND2_X1 U14383 ( .A1(n13967), .A2(n11801), .ZN(n11859) );
  NAND2_X1 U14384 ( .A1(n11860), .A2(n11859), .ZN(n11862) );
  XNOR2_X1 U14385 ( .A(n11862), .B(n11861), .ZN(n11864) );
  AOI22_X1 U14386 ( .A1(n14142), .A2(n11801), .B1(n11863), .B2(n13967), .ZN(
        n11865) );
  XNOR2_X1 U14387 ( .A(n11864), .B(n11865), .ZN(n13676) );
  INV_X1 U14388 ( .A(n11864), .ZN(n11866) );
  AOI22_X1 U14389 ( .A1(n13675), .A2(n13676), .B1(n11866), .B2(n11865), .ZN(
        n11872) );
  OAI22_X1 U14390 ( .A1(n14132), .A2(n10169), .B1(n14138), .B2(n11867), .ZN(
        n11870) );
  OAI22_X1 U14391 ( .A1(n14132), .A2(n11867), .B1(n14138), .B2(n9799), .ZN(
        n11868) );
  XNOR2_X1 U14392 ( .A(n11868), .B(n11861), .ZN(n11869) );
  XOR2_X1 U14393 ( .A(n11870), .B(n11869), .Z(n11871) );
  XNOR2_X1 U14394 ( .A(n11872), .B(n11871), .ZN(n11879) );
  OAI22_X1 U14395 ( .A1(n14503), .A2(n14147), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11873), .ZN(n11877) );
  INV_X1 U14396 ( .A(n11874), .ZN(n13934) );
  OAI22_X1 U14397 ( .A1(n14502), .A2(n11875), .B1(n14628), .B2(n13934), .ZN(
        n11876) );
  AOI211_X1 U14398 ( .C1(n13937), .C2(n14525), .A(n11877), .B(n11876), .ZN(
        n11878) );
  OAI21_X1 U14399 ( .B1(n11879), .B2(n14620), .A(n11878), .ZN(P1_U3220) );
  NAND2_X1 U14400 ( .A1(n15077), .A2(n11882), .ZN(n11926) );
  NAND2_X1 U14401 ( .A1(n11883), .A2(n6595), .ZN(n11884) );
  MUX2_X1 U14402 ( .A(n8917), .B(n11885), .S(n12030), .Z(n11888) );
  MUX2_X1 U14403 ( .A(n8917), .B(n11885), .S(n12032), .Z(n11886) );
  OAI211_X1 U14404 ( .C1(n11889), .C2(n11888), .A(n11887), .B(n12095), .ZN(
        n11895) );
  OAI21_X1 U14405 ( .B1(n13146), .B2(n12032), .A(n11890), .ZN(n11893) );
  NAND2_X1 U14406 ( .A1(n13146), .A2(n12032), .ZN(n11891) );
  NAND2_X1 U14407 ( .A1(n11891), .A2(n14865), .ZN(n11892) );
  NAND2_X1 U14408 ( .A1(n11893), .A2(n11892), .ZN(n11894) );
  NAND2_X1 U14409 ( .A1(n11895), .A2(n11894), .ZN(n11901) );
  MUX2_X1 U14410 ( .A(n13145), .B(n15068), .S(n12030), .Z(n11900) );
  NAND2_X1 U14411 ( .A1(n11901), .A2(n11900), .ZN(n11897) );
  NAND2_X1 U14412 ( .A1(n11897), .A2(n11896), .ZN(n11899) );
  OAI211_X1 U14413 ( .C1(n11901), .C2(n11900), .A(n11899), .B(n11898), .ZN(
        n11907) );
  OAI21_X1 U14414 ( .B1(n13144), .B2(n12032), .A(n14872), .ZN(n11905) );
  NAND2_X1 U14415 ( .A1(n13144), .A2(n12032), .ZN(n11903) );
  NAND2_X1 U14416 ( .A1(n11903), .A2(n11902), .ZN(n11904) );
  NAND2_X1 U14417 ( .A1(n11905), .A2(n11904), .ZN(n11906) );
  MUX2_X1 U14418 ( .A(n13143), .B(n11908), .S(n12030), .Z(n11912) );
  NAND2_X1 U14419 ( .A1(n11910), .A2(n11909), .ZN(n11911) );
  OAI211_X1 U14420 ( .C1(n11913), .C2(n11912), .A(n11911), .B(n12102), .ZN(
        n11917) );
  AND2_X1 U14421 ( .A1(n13142), .A2(n12032), .ZN(n11915) );
  OAI21_X1 U14422 ( .B1(n13142), .B2(n12032), .A(n13104), .ZN(n11914) );
  OAI21_X1 U14423 ( .B1(n11915), .B2(n13104), .A(n11914), .ZN(n11916) );
  NAND2_X1 U14424 ( .A1(n11917), .A2(n11916), .ZN(n11920) );
  MUX2_X1 U14425 ( .A(n13141), .B(n11918), .S(n12030), .Z(n11921) );
  MUX2_X1 U14426 ( .A(n13141), .B(n11918), .S(n12032), .Z(n11919) );
  AND2_X1 U14427 ( .A1(n13140), .A2(n12032), .ZN(n11924) );
  OAI21_X1 U14428 ( .B1(n13140), .B2(n12032), .A(n11923), .ZN(n11922) );
  OAI21_X1 U14429 ( .B1(n11924), .B2(n11923), .A(n11922), .ZN(n11925) );
  MUX2_X1 U14430 ( .A(n13139), .B(n13492), .S(n12030), .Z(n11930) );
  NAND2_X1 U14431 ( .A1(n11929), .A2(n11930), .ZN(n11928) );
  MUX2_X1 U14432 ( .A(n13139), .B(n13492), .S(n12031), .Z(n11927) );
  NAND2_X1 U14433 ( .A1(n11928), .A2(n11927), .ZN(n11934) );
  INV_X1 U14434 ( .A(n11929), .ZN(n11932) );
  INV_X1 U14435 ( .A(n11930), .ZN(n11931) );
  NAND2_X1 U14436 ( .A1(n11932), .A2(n11931), .ZN(n11933) );
  MUX2_X1 U14437 ( .A(n13138), .B(n13479), .S(n12031), .Z(n11938) );
  NAND2_X1 U14438 ( .A1(n11937), .A2(n11938), .ZN(n11936) );
  MUX2_X1 U14439 ( .A(n13138), .B(n13479), .S(n12030), .Z(n11935) );
  INV_X1 U14440 ( .A(n11937), .ZN(n11940) );
  INV_X1 U14441 ( .A(n11938), .ZN(n11939) );
  MUX2_X1 U14442 ( .A(n13137), .B(n13600), .S(n12030), .Z(n11942) );
  MUX2_X1 U14443 ( .A(n13137), .B(n13600), .S(n12031), .Z(n11941) );
  INV_X1 U14444 ( .A(n11942), .ZN(n11943) );
  MUX2_X1 U14445 ( .A(n13136), .B(n11944), .S(n12031), .Z(n11948) );
  NAND2_X1 U14446 ( .A1(n11947), .A2(n11948), .ZN(n11946) );
  MUX2_X1 U14447 ( .A(n13136), .B(n11944), .S(n12077), .Z(n11945) );
  NAND2_X1 U14448 ( .A1(n11946), .A2(n11945), .ZN(n11952) );
  INV_X1 U14449 ( .A(n11947), .ZN(n11950) );
  INV_X1 U14450 ( .A(n11948), .ZN(n11949) );
  NAND2_X1 U14451 ( .A1(n11950), .A2(n11949), .ZN(n11951) );
  MUX2_X1 U14452 ( .A(n13135), .B(n13645), .S(n12077), .Z(n11956) );
  NAND2_X1 U14453 ( .A1(n11955), .A2(n11956), .ZN(n11954) );
  MUX2_X1 U14454 ( .A(n13135), .B(n13645), .S(n12031), .Z(n11953) );
  NAND2_X1 U14455 ( .A1(n11954), .A2(n11953), .ZN(n11960) );
  INV_X1 U14456 ( .A(n11955), .ZN(n11958) );
  INV_X1 U14457 ( .A(n11956), .ZN(n11957) );
  NAND2_X1 U14458 ( .A1(n11958), .A2(n11957), .ZN(n11959) );
  MUX2_X1 U14459 ( .A(n13134), .B(n13589), .S(n12031), .Z(n11964) );
  NAND2_X1 U14460 ( .A1(n11963), .A2(n11964), .ZN(n11962) );
  MUX2_X1 U14461 ( .A(n13134), .B(n13589), .S(n12077), .Z(n11961) );
  NAND2_X1 U14462 ( .A1(n11962), .A2(n11961), .ZN(n11968) );
  INV_X1 U14463 ( .A(n11963), .ZN(n11966) );
  INV_X1 U14464 ( .A(n11964), .ZN(n11965) );
  NAND2_X1 U14465 ( .A1(n11966), .A2(n11965), .ZN(n11967) );
  MUX2_X1 U14466 ( .A(n13425), .B(n13580), .S(n12030), .Z(n11970) );
  MUX2_X1 U14467 ( .A(n13425), .B(n13580), .S(n12031), .Z(n11969) );
  INV_X1 U14468 ( .A(n11970), .ZN(n11971) );
  MUX2_X1 U14469 ( .A(n13133), .B(n13577), .S(n12031), .Z(n11975) );
  NAND2_X1 U14470 ( .A1(n11974), .A2(n11975), .ZN(n11973) );
  MUX2_X1 U14471 ( .A(n13133), .B(n13577), .S(n12030), .Z(n11972) );
  NAND2_X1 U14472 ( .A1(n11973), .A2(n11972), .ZN(n11979) );
  INV_X1 U14473 ( .A(n11974), .ZN(n11977) );
  INV_X1 U14474 ( .A(n11975), .ZN(n11976) );
  NAND2_X1 U14475 ( .A1(n11977), .A2(n11976), .ZN(n11978) );
  MUX2_X1 U14476 ( .A(n13428), .B(n13634), .S(n12077), .Z(n11981) );
  INV_X1 U14477 ( .A(n11981), .ZN(n11982) );
  MUX2_X1 U14478 ( .A(n13132), .B(n13562), .S(n12031), .Z(n11986) );
  NAND2_X1 U14479 ( .A1(n11985), .A2(n11986), .ZN(n11984) );
  MUX2_X1 U14480 ( .A(n13132), .B(n13562), .S(n12077), .Z(n11983) );
  NAND2_X1 U14481 ( .A1(n11984), .A2(n11983), .ZN(n11990) );
  INV_X1 U14482 ( .A(n11985), .ZN(n11988) );
  INV_X1 U14483 ( .A(n11986), .ZN(n11987) );
  NAND2_X1 U14484 ( .A1(n11988), .A2(n11987), .ZN(n11989) );
  MUX2_X1 U14485 ( .A(n13386), .B(n13559), .S(n12077), .Z(n11992) );
  MUX2_X1 U14486 ( .A(n13386), .B(n13559), .S(n12031), .Z(n11991) );
  INV_X1 U14487 ( .A(n11992), .ZN(n11993) );
  MUX2_X1 U14488 ( .A(n13131), .B(n13553), .S(n12077), .Z(n11994) );
  INV_X1 U14489 ( .A(n11995), .ZN(n11998) );
  INV_X1 U14490 ( .A(n11996), .ZN(n11997) );
  MUX2_X1 U14491 ( .A(n13549), .B(n13353), .S(n12031), .Z(n12000) );
  MUX2_X1 U14492 ( .A(n13353), .B(n13549), .S(n12031), .Z(n11999) );
  MUX2_X1 U14493 ( .A(n13626), .B(n13130), .S(n12077), .Z(n12004) );
  NAND2_X1 U14494 ( .A1(n12003), .A2(n12004), .ZN(n12002) );
  MUX2_X1 U14495 ( .A(n13626), .B(n13130), .S(n12031), .Z(n12001) );
  NAND2_X1 U14496 ( .A1(n12002), .A2(n12001), .ZN(n12008) );
  INV_X1 U14497 ( .A(n12003), .ZN(n12006) );
  INV_X1 U14498 ( .A(n12004), .ZN(n12005) );
  NAND2_X1 U14499 ( .A1(n12006), .A2(n12005), .ZN(n12007) );
  MUX2_X1 U14500 ( .A(n13129), .B(n13313), .S(n12077), .Z(n12010) );
  INV_X1 U14501 ( .A(n12010), .ZN(n12011) );
  NAND2_X1 U14502 ( .A1(n12014), .A2(n12015), .ZN(n12013) );
  MUX2_X1 U14503 ( .A(n13529), .B(n13128), .S(n12031), .Z(n12012) );
  NAND2_X1 U14504 ( .A1(n12013), .A2(n12012), .ZN(n12019) );
  INV_X1 U14505 ( .A(n12014), .ZN(n12017) );
  INV_X1 U14506 ( .A(n12015), .ZN(n12016) );
  NAND2_X1 U14507 ( .A1(n12017), .A2(n12016), .ZN(n12018) );
  MUX2_X1 U14508 ( .A(n13127), .B(n13525), .S(n12077), .Z(n12023) );
  NAND2_X1 U14509 ( .A1(n12022), .A2(n12023), .ZN(n12021) );
  MUX2_X1 U14510 ( .A(n13127), .B(n13525), .S(n12031), .Z(n12020) );
  NAND2_X1 U14511 ( .A1(n12021), .A2(n12020), .ZN(n12027) );
  INV_X1 U14512 ( .A(n12022), .ZN(n12025) );
  INV_X1 U14513 ( .A(n12023), .ZN(n12024) );
  NAND2_X1 U14514 ( .A1(n12025), .A2(n12024), .ZN(n12026) );
  MUX2_X1 U14515 ( .A(n13245), .B(n13520), .S(n12031), .Z(n12035) );
  NAND2_X1 U14516 ( .A1(n12036), .A2(n12035), .ZN(n12029) );
  MUX2_X1 U14517 ( .A(n13245), .B(n13520), .S(n12077), .Z(n12028) );
  MUX2_X1 U14518 ( .A(n13253), .B(n13114), .S(n12030), .Z(n12054) );
  MUX2_X1 U14519 ( .A(n13514), .B(n13126), .S(n12031), .Z(n12053) );
  NAND2_X1 U14520 ( .A1(n12054), .A2(n12053), .ZN(n12034) );
  MUX2_X1 U14521 ( .A(n13244), .B(n13512), .S(n12031), .Z(n12039) );
  INV_X1 U14522 ( .A(n12039), .ZN(n12033) );
  NAND2_X1 U14523 ( .A1(n12033), .A2(n12038), .ZN(n12057) );
  MUX2_X1 U14524 ( .A(n12037), .B(n13125), .S(n12077), .Z(n12071) );
  INV_X1 U14525 ( .A(n12071), .ZN(n12051) );
  MUX2_X1 U14526 ( .A(n13125), .B(n12037), .S(n12077), .Z(n12070) );
  INV_X1 U14527 ( .A(n12038), .ZN(n12040) );
  NAND2_X1 U14528 ( .A1(n12040), .A2(n12039), .ZN(n12050) );
  NAND2_X1 U14529 ( .A1(n14254), .A2(n12059), .ZN(n12042) );
  INV_X1 U14530 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13650) );
  OR2_X1 U14531 ( .A1(n12061), .A2(n13650), .ZN(n12041) );
  INV_X1 U14532 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n12048) );
  NAND2_X1 U14533 ( .A1(n6601), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n12047) );
  INV_X1 U14534 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n12044) );
  OR2_X1 U14535 ( .A1(n6614), .A2(n12044), .ZN(n12046) );
  OAI211_X1 U14536 ( .C1(n12049), .C2(n12048), .A(n12047), .B(n12046), .ZN(
        n13218) );
  XNOR2_X1 U14537 ( .A(n13501), .B(n13218), .ZN(n12128) );
  OAI211_X1 U14538 ( .C1(n12051), .C2(n12070), .A(n12050), .B(n12128), .ZN(
        n12052) );
  INV_X1 U14539 ( .A(n12053), .ZN(n12056) );
  INV_X1 U14540 ( .A(n12054), .ZN(n12055) );
  NAND3_X1 U14541 ( .A1(n12057), .A2(n12056), .A3(n12055), .ZN(n12058) );
  NAND2_X1 U14542 ( .A1(n12060), .A2(n12059), .ZN(n12063) );
  OR2_X1 U14543 ( .A1(n12061), .A2(n12138), .ZN(n12062) );
  MUX2_X1 U14544 ( .A(n13610), .B(n13124), .S(n12077), .Z(n12076) );
  OAI211_X1 U14545 ( .C1(n12065), .C2(n12097), .A(n8101), .B(n12064), .ZN(
        n12066) );
  AOI21_X1 U14546 ( .B1(n13218), .B2(n12031), .A(n12066), .ZN(n12068) );
  INV_X1 U14547 ( .A(n13124), .ZN(n12067) );
  NOR2_X1 U14548 ( .A1(n12068), .A2(n12067), .ZN(n12069) );
  AOI21_X1 U14549 ( .B1(n13610), .B2(n12077), .A(n12069), .ZN(n12075) );
  INV_X1 U14550 ( .A(n12070), .ZN(n12072) );
  OAI22_X1 U14551 ( .A1(n12076), .A2(n12075), .B1(n12072), .B2(n12071), .ZN(
        n12073) );
  NAND2_X1 U14552 ( .A1(n12073), .A2(n12128), .ZN(n12074) );
  NAND2_X1 U14553 ( .A1(n12076), .A2(n12075), .ZN(n12081) );
  AND2_X1 U14554 ( .A1(n13218), .A2(n12077), .ZN(n12079) );
  NOR2_X1 U14555 ( .A1(n13218), .A2(n12077), .ZN(n12078) );
  MUX2_X1 U14556 ( .A(n12079), .B(n12078), .S(n13501), .Z(n12080) );
  MUX2_X1 U14557 ( .A(n8102), .B(n8101), .S(n12097), .Z(n12082) );
  NAND2_X1 U14558 ( .A1(n12082), .A2(n6689), .ZN(n12083) );
  NAND2_X1 U14559 ( .A1(n12084), .A2(n12083), .ZN(n12089) );
  NOR2_X1 U14560 ( .A1(n8102), .A2(n6595), .ZN(n12086) );
  AOI211_X1 U14561 ( .C1(n8101), .C2(n13312), .A(n12086), .B(n12132), .ZN(
        n12087) );
  NAND2_X1 U14562 ( .A1(n12089), .A2(n12088), .ZN(n12137) );
  NOR2_X1 U14563 ( .A1(n12090), .A2(P2_U3088), .ZN(n12131) );
  INV_X1 U14564 ( .A(n12131), .ZN(n13669) );
  XNOR2_X1 U14565 ( .A(n13610), .B(n13124), .ZN(n12126) );
  XNOR2_X1 U14566 ( .A(n13589), .B(n12093), .ZN(n13457) );
  NAND4_X1 U14567 ( .A1(n14855), .A2(n12097), .A3(n12096), .A4(n12095), .ZN(
        n12100) );
  NOR3_X1 U14568 ( .A1(n12100), .A2(n12099), .A3(n12098), .ZN(n12103) );
  NAND4_X1 U14569 ( .A1(n12104), .A2(n12103), .A3(n12102), .A4(n12101), .ZN(
        n12105) );
  NOR2_X1 U14570 ( .A1(n7107), .A2(n12105), .ZN(n12108) );
  NAND4_X1 U14571 ( .A1(n12109), .A2(n12108), .A3(n12107), .A4(n12106), .ZN(
        n12110) );
  OR4_X1 U14572 ( .A1(n13440), .A2(n12112), .A3(n12111), .A4(n12110), .ZN(
        n12113) );
  OR4_X1 U14573 ( .A1(n13411), .A2(n13419), .A3(n13457), .A4(n12113), .ZN(
        n12114) );
  NOR2_X1 U14574 ( .A1(n13384), .A2(n12114), .ZN(n12117) );
  XNOR2_X1 U14575 ( .A(n13553), .B(n13131), .ZN(n13352) );
  NAND2_X1 U14576 ( .A1(n12116), .A2(n12115), .ZN(n13366) );
  NAND4_X1 U14577 ( .A1(n13338), .A2(n12117), .A3(n13352), .A4(n13366), .ZN(
        n12118) );
  NOR2_X1 U14578 ( .A1(n12119), .A2(n12118), .ZN(n12120) );
  NAND4_X1 U14579 ( .A1(n13285), .A2(n12121), .A3(n13315), .A4(n12120), .ZN(
        n12122) );
  NOR2_X1 U14580 ( .A1(n12123), .A2(n12122), .ZN(n12125) );
  AND4_X1 U14581 ( .A1(n12126), .A2(n12125), .A3(n12124), .A4(n13258), .ZN(
        n12127) );
  NAND3_X1 U14582 ( .A1(n12128), .A2(n12127), .A3(n13233), .ZN(n12129) );
  XNOR2_X1 U14583 ( .A(n12129), .B(n6689), .ZN(n12130) );
  NAND4_X1 U14584 ( .A1(n14854), .A2(n12133), .A3(n12132), .A4(n13426), .ZN(
        n12134) );
  OAI211_X1 U14585 ( .C1(n8102), .C2(n13669), .A(n12134), .B(P2_B_REG_SCAN_IN), 
        .ZN(n12135) );
  OAI211_X1 U14586 ( .C1(n12137), .C2(n13669), .A(n12136), .B(n12135), .ZN(
        P2_U3328) );
  XNOR2_X1 U14587 ( .A(n12461), .B(n12139), .ZN(n12147) );
  INV_X1 U14588 ( .A(n12147), .ZN(n12140) );
  NAND2_X1 U14589 ( .A1(n12140), .A2(n12216), .ZN(n12154) );
  INV_X1 U14590 ( .A(n12141), .ZN(n12142) );
  NAND4_X1 U14591 ( .A1(n12153), .A2(n12142), .A3(n12216), .A4(n12147), .ZN(
        n12152) );
  AOI22_X1 U14592 ( .A1(n12489), .A2(n12264), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12144) );
  NAND2_X1 U14593 ( .A1(n12635), .A2(n12243), .ZN(n12143) );
  OAI211_X1 U14594 ( .C1(n12145), .C2(n12261), .A(n12144), .B(n12143), .ZN(
        n12149) );
  NOR4_X1 U14595 ( .A1(n12147), .A2(n14886), .A3(n12146), .A4(n12489), .ZN(
        n12148) );
  AOI211_X1 U14596 ( .C1(n12150), .C2(n12268), .A(n12149), .B(n12148), .ZN(
        n12151) );
  OAI211_X1 U14597 ( .C1(n12154), .C2(n12153), .A(n12152), .B(n12151), .ZN(
        P3_U3160) );
  INV_X1 U14598 ( .A(n12155), .ZN(n12156) );
  OAI222_X1 U14599 ( .A1(P3_U3151), .A2(n12602), .B1(n12997), .B2(n12156), 
        .C1(n7635), .C2(n12995), .ZN(P3_U3268) );
  XOR2_X1 U14600 ( .A(n12158), .B(n12157), .Z(n12166) );
  INV_X1 U14601 ( .A(n12976), .ZN(n12164) );
  NOR2_X1 U14602 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12159), .ZN(n12524) );
  NOR2_X1 U14603 ( .A1(n12160), .A2(n12261), .ZN(n12161) );
  AOI211_X1 U14604 ( .C1(n12264), .C2(n12821), .A(n12524), .B(n12161), .ZN(
        n12162) );
  OAI21_X1 U14605 ( .B1(n12826), .B2(n12266), .A(n12162), .ZN(n12163) );
  AOI21_X1 U14606 ( .B1(n12164), .B2(n12268), .A(n12163), .ZN(n12165) );
  OAI21_X1 U14607 ( .B1(n12166), .B2(n14886), .A(n12165), .ZN(P3_U3155) );
  INV_X1 U14608 ( .A(n12169), .ZN(n12215) );
  AOI21_X1 U14609 ( .B1(n12685), .B2(n12167), .A(n12215), .ZN(n12174) );
  AOI22_X1 U14610 ( .A1(n12702), .A2(n12264), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12171) );
  NAND2_X1 U14611 ( .A1(n12243), .A2(n12711), .ZN(n12170) );
  OAI211_X1 U14612 ( .C1(n12705), .C2(n12261), .A(n12171), .B(n12170), .ZN(
        n12172) );
  AOI21_X1 U14613 ( .B1(n12706), .B2(n12268), .A(n12172), .ZN(n12173) );
  OAI21_X1 U14614 ( .B1(n12174), .B2(n14886), .A(n12173), .ZN(P3_U3156) );
  XOR2_X1 U14615 ( .A(n12176), .B(n12175), .Z(n12177) );
  NAND2_X1 U14616 ( .A1(n12177), .A2(n12216), .ZN(n12181) );
  NAND2_X1 U14617 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12611)
         );
  OAI21_X1 U14618 ( .B1(n12733), .B2(n12261), .A(n12611), .ZN(n12179) );
  NOR2_X1 U14619 ( .A1(n12266), .A2(n12759), .ZN(n12178) );
  AOI211_X1 U14620 ( .C1(n12264), .C2(n12781), .A(n12179), .B(n12178), .ZN(
        n12180) );
  OAI211_X1 U14621 ( .C1(n14891), .C2(n12962), .A(n12181), .B(n12180), .ZN(
        P3_U3159) );
  INV_X1 U14622 ( .A(n12182), .ZN(n12954) );
  INV_X1 U14623 ( .A(n12183), .ZN(n12185) );
  NOR3_X1 U14624 ( .A1(n6480), .A2(n12185), .A3(n12184), .ZN(n12188) );
  OR2_X1 U14625 ( .A1(n12186), .A2(n6485), .ZN(n12187) );
  OAI21_X1 U14626 ( .B1(n12188), .B2(n12187), .A(n12216), .ZN(n12192) );
  AOI22_X1 U14627 ( .A1(n12755), .A2(n12264), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12189) );
  OAI21_X1 U14628 ( .B1(n12734), .B2(n12261), .A(n12189), .ZN(n12190) );
  AOI21_X1 U14629 ( .B1(n12737), .B2(n12243), .A(n12190), .ZN(n12191) );
  OAI211_X1 U14630 ( .C1(n12954), .C2(n14891), .A(n12192), .B(n12191), .ZN(
        P3_U3163) );
  XNOR2_X1 U14631 ( .A(n12194), .B(n12193), .ZN(n12200) );
  NOR2_X1 U14632 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12195), .ZN(n12547) );
  NOR2_X1 U14633 ( .A1(n12769), .A2(n12261), .ZN(n12196) );
  AOI211_X1 U14634 ( .C1(n12264), .C2(n12820), .A(n12547), .B(n12196), .ZN(
        n12197) );
  OAI21_X1 U14635 ( .B1(n12794), .B2(n12266), .A(n12197), .ZN(n12198) );
  AOI21_X1 U14636 ( .B1(n12914), .B2(n12268), .A(n12198), .ZN(n12199) );
  OAI21_X1 U14637 ( .B1(n12200), .B2(n14886), .A(n12199), .ZN(P3_U3166) );
  INV_X1 U14638 ( .A(n12202), .ZN(n12203) );
  AOI21_X1 U14639 ( .B1(n12204), .B2(n12201), .A(n12203), .ZN(n12210) );
  NAND2_X1 U14640 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12566)
         );
  OAI21_X1 U14641 ( .B1(n12205), .B2(n12261), .A(n12566), .ZN(n12206) );
  AOI21_X1 U14642 ( .B1(n12264), .B2(n12805), .A(n12206), .ZN(n12207) );
  OAI21_X1 U14643 ( .B1(n12783), .B2(n12266), .A(n12207), .ZN(n12208) );
  AOI21_X1 U14644 ( .B1(n12910), .B2(n12268), .A(n12208), .ZN(n12209) );
  OAI21_X1 U14645 ( .B1(n12210), .B2(n14886), .A(n12209), .ZN(P3_U3168) );
  INV_X1 U14646 ( .A(n12211), .ZN(n12943) );
  INV_X1 U14647 ( .A(n12212), .ZN(n12214) );
  NOR3_X1 U14648 ( .A1(n12215), .A2(n12214), .A3(n12213), .ZN(n12218) );
  OAI21_X1 U14649 ( .B1(n12218), .B2(n12217), .A(n12216), .ZN(n12222) );
  AOI22_X1 U14650 ( .A1(n12686), .A2(n14888), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12219) );
  OAI21_X1 U14651 ( .B1(n12719), .B2(n12227), .A(n12219), .ZN(n12220) );
  AOI21_X1 U14652 ( .B1(n12694), .B2(n12243), .A(n12220), .ZN(n12221) );
  OAI211_X1 U14653 ( .C1(n12943), .C2(n14891), .A(n12222), .B(n12221), .ZN(
        P3_U3169) );
  AOI21_X1 U14654 ( .B1(n12224), .B2(n12223), .A(n6480), .ZN(n12230) );
  NAND2_X1 U14655 ( .A1(n12243), .A2(n12748), .ZN(n12226) );
  AOI22_X1 U14656 ( .A1(n14888), .A2(n12490), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12225) );
  OAI211_X1 U14657 ( .C1(n12770), .C2(n12227), .A(n12226), .B(n12225), .ZN(
        n12228) );
  AOI21_X1 U14658 ( .B1(n12747), .B2(n12268), .A(n12228), .ZN(n12229) );
  OAI21_X1 U14659 ( .B1(n12230), .B2(n14886), .A(n12229), .ZN(P3_U3173) );
  NOR2_X1 U14660 ( .A1(n12231), .A2(n6579), .ZN(n12232) );
  XNOR2_X1 U14661 ( .A(n12233), .B(n12232), .ZN(n12239) );
  AND2_X1 U14662 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n14993) );
  NOR2_X1 U14663 ( .A1(n12234), .A2(n12261), .ZN(n12235) );
  AOI211_X1 U14664 ( .C1(n12264), .C2(n12843), .A(n14993), .B(n12235), .ZN(
        n12236) );
  OAI21_X1 U14665 ( .B1(n12848), .B2(n12266), .A(n12236), .ZN(n12237) );
  AOI21_X1 U14666 ( .B1(n12847), .B2(n12268), .A(n12237), .ZN(n12238) );
  OAI21_X1 U14667 ( .B1(n12239), .B2(n14886), .A(n12238), .ZN(P3_U3174) );
  INV_X1 U14668 ( .A(n12241), .ZN(n12242) );
  AOI21_X1 U14669 ( .B1(n12702), .B2(n12240), .A(n12242), .ZN(n12248) );
  AOI22_X1 U14670 ( .A1(n12264), .A2(n12490), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12245) );
  NAND2_X1 U14671 ( .A1(n12243), .A2(n12723), .ZN(n12244) );
  OAI211_X1 U14672 ( .C1(n12719), .C2(n12261), .A(n12245), .B(n12244), .ZN(
        n12246) );
  AOI21_X1 U14673 ( .B1(n12722), .B2(n12268), .A(n12246), .ZN(n12247) );
  OAI21_X1 U14674 ( .B1(n12248), .B2(n14886), .A(n12247), .ZN(P3_U3175) );
  INV_X1 U14675 ( .A(n12249), .ZN(n12966) );
  AOI21_X1 U14676 ( .B1(n12251), .B2(n12250), .A(n14886), .ZN(n12253) );
  NAND2_X1 U14677 ( .A1(n12253), .A2(n12252), .ZN(n12257) );
  NAND2_X1 U14678 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12583)
         );
  OAI21_X1 U14679 ( .B1(n12770), .B2(n12261), .A(n12583), .ZN(n12255) );
  NOR2_X1 U14680 ( .A1(n12266), .A2(n12774), .ZN(n12254) );
  AOI211_X1 U14681 ( .C1(n12264), .C2(n12792), .A(n12255), .B(n12254), .ZN(
        n12256) );
  OAI211_X1 U14682 ( .C1(n12966), .C2(n14891), .A(n12257), .B(n12256), .ZN(
        P3_U3178) );
  XNOR2_X1 U14683 ( .A(n12258), .B(n12820), .ZN(n12259) );
  XNOR2_X1 U14684 ( .A(n12260), .B(n12259), .ZN(n12270) );
  AND2_X1 U14685 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n14469) );
  NOR2_X1 U14686 ( .A1(n12262), .A2(n12261), .ZN(n12263) );
  AOI211_X1 U14687 ( .C1(n12264), .C2(n12842), .A(n14469), .B(n12263), .ZN(
        n12265) );
  OAI21_X1 U14688 ( .B1(n12812), .B2(n12266), .A(n12265), .ZN(n12267) );
  AOI21_X1 U14689 ( .B1(n12811), .B2(n12268), .A(n12267), .ZN(n12269) );
  OAI21_X1 U14690 ( .B1(n12270), .B2(n14886), .A(n12269), .ZN(P3_U3181) );
  INV_X1 U14691 ( .A(n12271), .ZN(n12272) );
  NAND2_X1 U14692 ( .A1(n12274), .A2(n12273), .ZN(n12276) );
  XNOR2_X1 U14693 ( .A(n13650), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n12275) );
  XNOR2_X1 U14694 ( .A(n12276), .B(n12275), .ZN(n12983) );
  NAND2_X1 U14695 ( .A1(n12983), .A2(n12277), .ZN(n12279) );
  INV_X1 U14696 ( .A(SI_31_), .ZN(n12989) );
  OR2_X1 U14697 ( .A1(n8258), .A2(n12989), .ZN(n12278) );
  OR2_X1 U14698 ( .A1(n12290), .A2(n12280), .ZN(n12287) );
  OR2_X1 U14699 ( .A1(n12282), .A2(n12281), .ZN(n12285) );
  OR2_X1 U14700 ( .A1(n8258), .A2(n12283), .ZN(n12284) );
  NAND2_X1 U14701 ( .A1(n14474), .A2(n12289), .ZN(n12286) );
  NAND2_X1 U14702 ( .A1(n12287), .A2(n12286), .ZN(n12296) );
  INV_X1 U14703 ( .A(n14474), .ZN(n12628) );
  OAI21_X1 U14704 ( .B1(n12628), .B2(n12624), .A(n12464), .ZN(n12288) );
  NOR2_X1 U14705 ( .A1(n12296), .A2(n12288), .ZN(n12293) );
  NOR2_X1 U14706 ( .A1(n14474), .A2(n12289), .ZN(n12318) );
  XNOR2_X1 U14707 ( .A(n12295), .B(n12612), .ZN(n12480) );
  INV_X1 U14708 ( .A(n12296), .ZN(n12472) );
  INV_X1 U14709 ( .A(n12461), .ZN(n12454) );
  NAND2_X1 U14710 ( .A1(n12450), .A2(n12449), .ZN(n12655) );
  INV_X1 U14711 ( .A(n12655), .ZN(n12315) );
  NAND2_X1 U14712 ( .A1(n12430), .A2(n12431), .ZN(n12720) );
  INV_X1 U14713 ( .A(n12731), .ZN(n12735) );
  NOR2_X1 U14714 ( .A1(n12720), .A2(n12735), .ZN(n12297) );
  AND2_X1 U14715 ( .A1(n12707), .A2(n12297), .ZN(n12429) );
  INV_X1 U14716 ( .A(n12429), .ZN(n12312) );
  INV_X1 U14717 ( .A(n9979), .ZN(n12299) );
  NAND4_X1 U14718 ( .A1(n12300), .A2(n12299), .A3(n12298), .A4(n12346), .ZN(
        n12303) );
  INV_X1 U14719 ( .A(n12301), .ZN(n12374) );
  NAND3_X1 U14720 ( .A1(n14887), .A2(n12374), .A3(n12363), .ZN(n12302) );
  NOR2_X1 U14721 ( .A1(n12303), .A2(n12302), .ZN(n12307) );
  INV_X1 U14722 ( .A(n12304), .ZN(n12385) );
  AND3_X1 U14723 ( .A1(n12385), .A2(n12344), .A3(n12305), .ZN(n12306) );
  AND4_X1 U14724 ( .A1(n12307), .A2(n12855), .A3(n12306), .A4(n12369), .ZN(
        n12308) );
  INV_X1 U14725 ( .A(n12839), .ZN(n12835) );
  NAND4_X1 U14726 ( .A1(n12308), .A2(n8437), .A3(n12382), .A4(n12835), .ZN(
        n12309) );
  NOR2_X1 U14727 ( .A1(n12309), .A2(n12803), .ZN(n12310) );
  NAND4_X1 U14728 ( .A1(n12772), .A2(n12798), .A3(n12788), .A4(n12310), .ZN(
        n12311) );
  OR4_X1 U14729 ( .A1(n12312), .A2(n12743), .A3(n7446), .A4(n12311), .ZN(
        n12313) );
  NOR2_X1 U14730 ( .A1(n12689), .A2(n12313), .ZN(n12314) );
  NAND4_X1 U14731 ( .A1(n12452), .A2(n12672), .A3(n12315), .A4(n12314), .ZN(
        n12316) );
  NOR3_X1 U14732 ( .A1(n12317), .A2(n12454), .A3(n12316), .ZN(n12320) );
  INV_X1 U14733 ( .A(n12318), .ZN(n12467) );
  INV_X1 U14734 ( .A(n12470), .ZN(n12319) );
  MUX2_X1 U14735 ( .A(n12322), .B(n12321), .S(n12457), .Z(n12428) );
  MUX2_X1 U14736 ( .A(n12331), .B(n12326), .S(n12457), .Z(n12335) );
  NAND2_X1 U14737 ( .A1(n12325), .A2(n12323), .ZN(n12324) );
  NAND2_X1 U14738 ( .A1(n12324), .A2(n12457), .ZN(n12328) );
  NAND3_X1 U14739 ( .A1(n12326), .A2(n12325), .A3(n12484), .ZN(n12327) );
  NAND2_X1 U14740 ( .A1(n12328), .A2(n12327), .ZN(n12333) );
  NAND2_X1 U14741 ( .A1(n12330), .A2(n12329), .ZN(n12332) );
  NAND3_X1 U14742 ( .A1(n12333), .A2(n12332), .A3(n12331), .ZN(n12334) );
  NAND3_X1 U14743 ( .A1(n12335), .A2(n12305), .A3(n12334), .ZN(n12339) );
  NAND2_X1 U14744 ( .A1(n12499), .A2(n8789), .ZN(n12336) );
  NAND2_X1 U14745 ( .A1(n12345), .A2(n12336), .ZN(n12337) );
  NAND2_X1 U14746 ( .A1(n12337), .A2(n12460), .ZN(n12338) );
  NAND2_X1 U14747 ( .A1(n12339), .A2(n12338), .ZN(n12343) );
  AOI21_X1 U14748 ( .B1(n12342), .B2(n12340), .A(n12460), .ZN(n12341) );
  AOI21_X1 U14749 ( .B1(n12343), .B2(n12342), .A(n12341), .ZN(n12348) );
  OAI21_X1 U14750 ( .B1(n12460), .B2(n12345), .A(n12344), .ZN(n12347) );
  OAI21_X1 U14751 ( .B1(n12348), .B2(n12347), .A(n12346), .ZN(n12358) );
  NAND2_X1 U14752 ( .A1(n12360), .A2(n12349), .ZN(n12352) );
  NAND2_X1 U14753 ( .A1(n12352), .A2(n12457), .ZN(n12357) );
  NAND2_X1 U14754 ( .A1(n12350), .A2(n12457), .ZN(n12351) );
  NOR2_X1 U14755 ( .A1(n12352), .A2(n12351), .ZN(n12355) );
  AND2_X1 U14756 ( .A1(n12353), .A2(n12460), .ZN(n12354) );
  MUX2_X1 U14757 ( .A(n12355), .B(n12354), .S(n15012), .Z(n12356) );
  AOI21_X1 U14758 ( .B1(n12358), .B2(n12357), .A(n12356), .ZN(n12365) );
  AOI21_X1 U14759 ( .B1(n12361), .B2(n12359), .A(n12457), .ZN(n12364) );
  MUX2_X1 U14760 ( .A(n12361), .B(n12360), .S(n12460), .Z(n12362) );
  OAI211_X1 U14761 ( .C1(n12365), .C2(n12364), .A(n12363), .B(n12362), .ZN(
        n12370) );
  MUX2_X1 U14762 ( .A(n12367), .B(n12366), .S(n12460), .Z(n12368) );
  NAND3_X1 U14763 ( .A1(n12370), .A2(n12369), .A3(n12368), .ZN(n12375) );
  NAND2_X1 U14764 ( .A1(n12494), .A2(n15032), .ZN(n12371) );
  MUX2_X1 U14765 ( .A(n12372), .B(n12371), .S(n12460), .Z(n12373) );
  NAND3_X1 U14766 ( .A1(n12375), .A2(n12374), .A3(n12373), .ZN(n12379) );
  MUX2_X1 U14767 ( .A(n12377), .B(n12376), .S(n12457), .Z(n12378) );
  NAND2_X1 U14768 ( .A1(n12379), .A2(n12378), .ZN(n12386) );
  MUX2_X1 U14769 ( .A(n12381), .B(n12380), .S(n12457), .Z(n12383) );
  NAND2_X1 U14770 ( .A1(n12383), .A2(n12382), .ZN(n12384) );
  AOI21_X1 U14771 ( .B1(n12386), .B2(n12385), .A(n12384), .ZN(n12395) );
  NAND2_X1 U14772 ( .A1(n12392), .A2(n12387), .ZN(n12390) );
  OAI21_X1 U14773 ( .B1(n12859), .B2(n12388), .A(n12391), .ZN(n12389) );
  MUX2_X1 U14774 ( .A(n12390), .B(n12389), .S(n12460), .Z(n12394) );
  MUX2_X1 U14775 ( .A(n12392), .B(n12391), .S(n12457), .Z(n12393) );
  OAI211_X1 U14776 ( .C1(n12395), .C2(n12394), .A(n12835), .B(n12393), .ZN(
        n12399) );
  MUX2_X1 U14777 ( .A(n12397), .B(n12396), .S(n12457), .Z(n12398) );
  NAND4_X1 U14778 ( .A1(n12399), .A2(n12810), .A3(n8437), .A4(n12398), .ZN(
        n12404) );
  OAI211_X1 U14779 ( .C1(n12803), .C2(n12401), .A(n12409), .B(n12400), .ZN(
        n12402) );
  NAND2_X1 U14780 ( .A1(n12402), .A2(n12457), .ZN(n12403) );
  AOI21_X1 U14781 ( .B1(n12404), .B2(n12403), .A(n7043), .ZN(n12411) );
  OAI211_X1 U14782 ( .C1(n12803), .C2(n12407), .A(n12406), .B(n12405), .ZN(
        n12408) );
  AND2_X1 U14783 ( .A1(n12408), .A2(n12460), .ZN(n12410) );
  OAI22_X1 U14784 ( .A1(n12411), .A2(n12410), .B1(n12409), .B2(n12457), .ZN(
        n12417) );
  INV_X1 U14785 ( .A(n12412), .ZN(n12413) );
  NAND2_X1 U14786 ( .A1(n12418), .A2(n12413), .ZN(n12414) );
  NAND4_X1 U14787 ( .A1(n12424), .A2(n12460), .A3(n12415), .A4(n12414), .ZN(
        n12420) );
  AOI22_X1 U14788 ( .A1(n12417), .A2(n12788), .B1(n12416), .B2(n12420), .ZN(
        n12422) );
  NAND3_X1 U14789 ( .A1(n12423), .A2(n12418), .A3(n12457), .ZN(n12419) );
  NAND2_X1 U14790 ( .A1(n12420), .A2(n12419), .ZN(n12421) );
  OAI21_X1 U14791 ( .B1(n12422), .B2(n8690), .A(n12421), .ZN(n12426) );
  MUX2_X1 U14792 ( .A(n12424), .B(n12423), .S(n12460), .Z(n12425) );
  NAND3_X1 U14793 ( .A1(n12426), .A2(n8539), .A3(n12425), .ZN(n12427) );
  NAND3_X1 U14794 ( .A1(n12429), .A2(n12428), .A3(n12427), .ZN(n12439) );
  MUX2_X1 U14795 ( .A(n12431), .B(n12430), .S(n12460), .Z(n12436) );
  INV_X1 U14796 ( .A(n12720), .ZN(n12716) );
  MUX2_X1 U14797 ( .A(n12433), .B(n12432), .S(n12460), .Z(n12434) );
  NAND2_X1 U14798 ( .A1(n12716), .A2(n12434), .ZN(n12435) );
  NAND3_X1 U14799 ( .A1(n12707), .A2(n12436), .A3(n12435), .ZN(n12438) );
  NAND3_X1 U14800 ( .A1(n12706), .A2(n12719), .A3(n12460), .ZN(n12437) );
  AND3_X1 U14801 ( .A1(n12439), .A2(n12438), .A3(n12437), .ZN(n12444) );
  XNOR2_X1 U14802 ( .A(n12440), .B(n12460), .ZN(n12441) );
  OR2_X1 U14803 ( .A1(n12442), .A2(n12441), .ZN(n12443) );
  OAI211_X1 U14804 ( .C1(n12444), .C2(n12689), .A(n12672), .B(n12443), .ZN(
        n12448) );
  MUX2_X1 U14805 ( .A(n12446), .B(n12445), .S(n12457), .Z(n12447) );
  AND2_X1 U14806 ( .A1(n12448), .A2(n12447), .ZN(n12453) );
  MUX2_X1 U14807 ( .A(n12450), .B(n12449), .S(n12457), .Z(n12451) );
  OAI211_X1 U14808 ( .C1(n12453), .C2(n12655), .A(n12452), .B(n12451), .ZN(
        n12459) );
  AOI21_X1 U14809 ( .B1(n12455), .B2(n12459), .A(n12454), .ZN(n12466) );
  OAI21_X1 U14810 ( .B1(n12458), .B2(n12457), .A(n12456), .ZN(n12465) );
  INV_X1 U14811 ( .A(n12459), .ZN(n12462) );
  NAND3_X1 U14812 ( .A1(n12462), .A2(n12461), .A3(n12460), .ZN(n12463) );
  OAI211_X1 U14813 ( .C1(n12466), .C2(n12465), .A(n12464), .B(n12463), .ZN(
        n12469) );
  NAND3_X1 U14814 ( .A1(n12469), .A2(n12468), .A3(n12467), .ZN(n12471) );
  AOI21_X1 U14815 ( .B1(n12472), .B2(n12471), .A(n12470), .ZN(n12473) );
  AOI21_X1 U14816 ( .B1(n12480), .B2(n12479), .A(n12478), .ZN(n12487) );
  NAND3_X1 U14817 ( .A1(n12482), .A2(n12481), .A3(n12602), .ZN(n12483) );
  OAI211_X1 U14818 ( .C1(n12484), .C2(n12486), .A(n12483), .B(P3_B_REG_SCAN_IN), .ZN(n12485) );
  OAI21_X1 U14819 ( .B1(n12487), .B2(n12486), .A(n12485), .ZN(P3_U3296) );
  MUX2_X1 U14820 ( .A(n12488), .B(P3_DATAO_REG_29__SCAN_IN), .S(n12500), .Z(
        P3_U3520) );
  MUX2_X1 U14821 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12489), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14822 ( .A(n12668), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12500), .Z(
        P3_U3517) );
  MUX2_X1 U14823 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12686), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14824 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12667), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14825 ( .A(n12685), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12500), .Z(
        P3_U3514) );
  MUX2_X1 U14826 ( .A(n12702), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12500), .Z(
        P3_U3513) );
  MUX2_X1 U14827 ( .A(n12490), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12500), .Z(
        P3_U3512) );
  MUX2_X1 U14828 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12755), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14829 ( .A(n12491), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12500), .Z(
        P3_U3510) );
  MUX2_X1 U14830 ( .A(n12781), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12500), .Z(
        P3_U3509) );
  MUX2_X1 U14831 ( .A(n12805), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12500), .Z(
        P3_U3507) );
  MUX2_X1 U14832 ( .A(n12820), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12500), .Z(
        P3_U3506) );
  MUX2_X1 U14833 ( .A(n12842), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12500), .Z(
        P3_U3505) );
  MUX2_X1 U14834 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12821), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14835 ( .A(n12843), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12500), .Z(
        P3_U3503) );
  MUX2_X1 U14836 ( .A(n12492), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12500), .Z(
        P3_U3501) );
  MUX2_X1 U14837 ( .A(n12493), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12500), .Z(
        P3_U3500) );
  MUX2_X1 U14838 ( .A(n12494), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12500), .Z(
        P3_U3499) );
  MUX2_X1 U14839 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12495), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14840 ( .A(n12496), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12500), .Z(
        P3_U3497) );
  MUX2_X1 U14841 ( .A(n12497), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12500), .Z(
        P3_U3496) );
  MUX2_X1 U14842 ( .A(n12498), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12500), .Z(
        P3_U3494) );
  MUX2_X1 U14843 ( .A(n12499), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12500), .Z(
        P3_U3493) );
  MUX2_X1 U14844 ( .A(n10042), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12500), .Z(
        P3_U3492) );
  MUX2_X1 U14845 ( .A(n8666), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12500), .Z(
        P3_U3491) );
  NAND2_X1 U14846 ( .A1(n12527), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12551) );
  OAI21_X1 U14847 ( .B1(n12527), .B2(P3_REG1_REG_14__SCAN_IN), .A(n12551), 
        .ZN(n12520) );
  AOI21_X1 U14848 ( .B1(n12505), .B2(n12520), .A(n12549), .ZN(n12531) );
  NAND2_X1 U14849 ( .A1(n12527), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12539) );
  OAI21_X1 U14850 ( .B1(n12527), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12539), 
        .ZN(n12532) );
  XNOR2_X1 U14851 ( .A(n12533), .B(n12532), .ZN(n12529) );
  MUX2_X1 U14852 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12602), .Z(n12512) );
  NOR2_X1 U14853 ( .A1(n12512), .A2(n14980), .ZN(n12522) );
  XNOR2_X1 U14854 ( .A(n12512), .B(n14980), .ZN(n14986) );
  OR2_X1 U14855 ( .A1(n12514), .A2(n12513), .ZN(n12519) );
  INV_X1 U14856 ( .A(n12515), .ZN(n12517) );
  NAND2_X1 U14857 ( .A1(n12519), .A2(n12518), .ZN(n14985) );
  MUX2_X1 U14858 ( .A(n12532), .B(n12520), .S(n12602), .Z(n12521) );
  OAI21_X1 U14859 ( .B1(n12522), .B2(n14984), .A(n12521), .ZN(n12523) );
  NAND3_X1 U14860 ( .A1(n12523), .A2(n14945), .A3(n12541), .ZN(n12526) );
  AOI21_X1 U14861 ( .B1(n14972), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12524), 
        .ZN(n12525) );
  OAI211_X1 U14862 ( .C1(n14979), .C2(n12527), .A(n12526), .B(n12525), .ZN(
        n12528) );
  AOI21_X1 U14863 ( .B1(n12529), .B2(n14897), .A(n12528), .ZN(n12530) );
  OAI21_X1 U14864 ( .B1(n12531), .B2(n14989), .A(n12530), .ZN(P3_U3196) );
  NAND2_X1 U14865 ( .A1(n12539), .A2(n12534), .ZN(n12535) );
  INV_X1 U14866 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14455) );
  INV_X1 U14867 ( .A(n12555), .ZN(n14400) );
  INV_X1 U14868 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12536) );
  AOI22_X1 U14869 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12555), .B1(n14400), 
        .B2(n12536), .ZN(n12537) );
  AOI21_X1 U14870 ( .B1(n12538), .B2(n12537), .A(n12564), .ZN(n12563) );
  MUX2_X1 U14871 ( .A(n12539), .B(n12551), .S(n12602), .Z(n12540) );
  MUX2_X1 U14872 ( .A(n14455), .B(n14460), .S(n12602), .Z(n14461) );
  MUX2_X1 U14873 ( .A(n12536), .B(n12554), .S(n12602), .Z(n12543) );
  NAND2_X1 U14874 ( .A1(n12543), .A2(n12555), .ZN(n12567) );
  MUX2_X1 U14875 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12602), .Z(n12544) );
  AND2_X1 U14876 ( .A1(n12544), .A2(n14400), .ZN(n12568) );
  INV_X1 U14877 ( .A(n12568), .ZN(n12545) );
  NAND2_X1 U14878 ( .A1(n12567), .A2(n12545), .ZN(n12546) );
  XNOR2_X1 U14879 ( .A(n6453), .B(n12546), .ZN(n12561) );
  AOI21_X1 U14880 ( .B1(n14972), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n12547), 
        .ZN(n12548) );
  OAI21_X1 U14881 ( .B1(n14979), .B2(n14400), .A(n12548), .ZN(n12560) );
  AOI22_X1 U14882 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12555), .B1(n14400), 
        .B2(n12554), .ZN(n12556) );
  AOI21_X1 U14883 ( .B1(n12557), .B2(n12556), .A(n12573), .ZN(n12558) );
  NOR2_X1 U14884 ( .A1(n12558), .A2(n14989), .ZN(n12559) );
  AOI211_X1 U14885 ( .C1(n14945), .C2(n12561), .A(n12560), .B(n12559), .ZN(
        n12562) );
  OAI21_X1 U14886 ( .B1(n12563), .B2(n14995), .A(n12562), .ZN(P3_U3198) );
  AOI21_X1 U14887 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n14400), .A(n12564), 
        .ZN(n12580) );
  XNOR2_X1 U14888 ( .A(n12591), .B(n12580), .ZN(n12565) );
  AOI21_X1 U14889 ( .B1(n12565), .B2(n12784), .A(n12581), .ZN(n12579) );
  INV_X1 U14890 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14385) );
  OAI21_X1 U14891 ( .B1(n14978), .B2(n14385), .A(n12566), .ZN(n12572) );
  MUX2_X1 U14892 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12602), .Z(n12586) );
  XNOR2_X1 U14893 ( .A(n12586), .B(n12585), .ZN(n12569) );
  AOI211_X1 U14894 ( .C1(n12570), .C2(n12569), .A(n12584), .B(n14987), .ZN(
        n12571) );
  AOI211_X1 U14895 ( .C1(n14944), .C2(n12591), .A(n12572), .B(n12571), .ZN(
        n12578) );
  XNOR2_X1 U14896 ( .A(n12591), .B(n12590), .ZN(n12574) );
  AOI21_X1 U14897 ( .B1(n12575), .B2(n12574), .A(n12592), .ZN(n12576) );
  OR2_X1 U14898 ( .A1(n12576), .A2(n14989), .ZN(n12577) );
  OAI211_X1 U14899 ( .C1(n12579), .C2(n14995), .A(n12578), .B(n12577), .ZN(
        P3_U3199) );
  NAND2_X1 U14900 ( .A1(n12594), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12599) );
  OAI21_X1 U14901 ( .B1(n12594), .B2(P3_REG2_REG_18__SCAN_IN), .A(n12599), 
        .ZN(n12582) );
  AOI21_X1 U14902 ( .B1(n6550), .B2(n12582), .A(n12600), .ZN(n12598) );
  INV_X1 U14903 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14449) );
  OAI21_X1 U14904 ( .B1(n14978), .B2(n14449), .A(n12583), .ZN(n12589) );
  MUX2_X1 U14905 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12602), .Z(n12588) );
  XNOR2_X1 U14906 ( .A(n12607), .B(n12606), .ZN(n12587) );
  NOR2_X1 U14907 ( .A1(n12587), .A2(n12588), .ZN(n12605) );
  NOR2_X1 U14908 ( .A1(n12591), .A2(n12590), .ZN(n12593) );
  NAND2_X1 U14909 ( .A1(n12594), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12613) );
  OAI21_X1 U14910 ( .B1(n12594), .B2(P3_REG1_REG_18__SCAN_IN), .A(n12613), 
        .ZN(n12595) );
  AOI21_X1 U14911 ( .B1(n6547), .B2(n12595), .A(n12614), .ZN(n12596) );
  OR2_X1 U14912 ( .A1(n12596), .A2(n14989), .ZN(n12597) );
  MUX2_X1 U14913 ( .A(P3_REG2_REG_19__SCAN_IN), .B(n12760), .S(n12612), .Z(
        n12604) );
  XNOR2_X1 U14914 ( .A(n12601), .B(n12604), .ZN(n12619) );
  XNOR2_X1 U14915 ( .A(n12612), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12616) );
  INV_X1 U14916 ( .A(n12616), .ZN(n12603) );
  MUX2_X1 U14917 ( .A(n12604), .B(n12603), .S(n12602), .Z(n12609) );
  AOI21_X1 U14918 ( .B1(n12607), .B2(n12606), .A(n12605), .ZN(n12608) );
  NAND2_X1 U14919 ( .A1(n14972), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12610) );
  OAI211_X1 U14920 ( .C1(n14979), .C2(n12612), .A(n12611), .B(n12610), .ZN(
        n12617) );
  INV_X1 U14921 ( .A(n12620), .ZN(n12621) );
  NAND2_X1 U14922 ( .A1(n12621), .A2(n12828), .ZN(n12630) );
  INV_X1 U14923 ( .A(n12622), .ZN(n12623) );
  NAND2_X1 U14924 ( .A1(n12624), .A2(n12623), .ZN(n14472) );
  AOI21_X1 U14925 ( .B1(n12630), .B2(n14472), .A(n12868), .ZN(n12626) );
  AOI21_X1 U14926 ( .B1(n12833), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12626), 
        .ZN(n12625) );
  OAI21_X1 U14927 ( .B1(n12931), .B2(n12866), .A(n12625), .ZN(P3_U3202) );
  AOI21_X1 U14928 ( .B1(n12833), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12626), 
        .ZN(n12627) );
  OAI21_X1 U14929 ( .B1(n12628), .B2(n12866), .A(n12627), .ZN(P3_U3203) );
  NAND2_X1 U14930 ( .A1(n12833), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n12629) );
  OAI211_X1 U14931 ( .C1(n12631), .C2(n12866), .A(n12630), .B(n12629), .ZN(
        n12632) );
  AOI21_X1 U14932 ( .B1(n12633), .B2(n12831), .A(n12632), .ZN(n12634) );
  OAI21_X1 U14933 ( .B1(n6481), .B2(n12833), .A(n12634), .ZN(P3_U3204) );
  AOI22_X1 U14934 ( .A1(n12635), .A2(n12828), .B1(n12833), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12636) );
  OAI21_X1 U14935 ( .B1(n12637), .B2(n12866), .A(n12636), .ZN(n12638) );
  AOI21_X1 U14936 ( .B1(n12639), .B2(n12831), .A(n12638), .ZN(n12640) );
  OAI21_X1 U14937 ( .B1(n12641), .B2(n12833), .A(n12640), .ZN(P3_U3205) );
  INV_X1 U14938 ( .A(n12642), .ZN(n12650) );
  AOI22_X1 U14939 ( .A1(n12643), .A2(n12828), .B1(n12833), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12644) );
  OAI21_X1 U14940 ( .B1(n12645), .B2(n12866), .A(n12644), .ZN(n12646) );
  AOI21_X1 U14941 ( .B1(n12648), .B2(n12647), .A(n12646), .ZN(n12649) );
  OAI21_X1 U14942 ( .B1(n12650), .B2(n12833), .A(n12649), .ZN(P3_U3206) );
  NAND2_X1 U14943 ( .A1(n12664), .A2(n12651), .ZN(n12652) );
  INV_X1 U14944 ( .A(n12874), .ZN(n12660) );
  XOR2_X1 U14945 ( .A(n12655), .B(n12654), .Z(n12875) );
  AOI22_X1 U14946 ( .A1(n12656), .A2(n12828), .B1(n12868), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12657) );
  OAI21_X1 U14947 ( .B1(n12935), .B2(n12866), .A(n12657), .ZN(n12658) );
  AOI21_X1 U14948 ( .B1(n12875), .B2(n12831), .A(n12658), .ZN(n12659) );
  OAI21_X1 U14949 ( .B1(n12660), .B2(n12833), .A(n12659), .ZN(P3_U3207) );
  OR2_X1 U14950 ( .A1(n12661), .A2(n12662), .ZN(n12680) );
  NAND2_X1 U14951 ( .A1(n12680), .A2(n12663), .ZN(n12666) );
  OAI211_X1 U14952 ( .C1(n12666), .C2(n12665), .A(n12664), .B(n12837), .ZN(
        n12670) );
  AOI22_X1 U14953 ( .A1(n12668), .A2(n12841), .B1(n12667), .B2(n12844), .ZN(
        n12669) );
  NAND2_X1 U14954 ( .A1(n12670), .A2(n12669), .ZN(n12878) );
  INV_X1 U14955 ( .A(n12878), .ZN(n12678) );
  OAI21_X1 U14956 ( .B1(n12673), .B2(n12672), .A(n12671), .ZN(n12879) );
  AOI22_X1 U14957 ( .A1(n12868), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n12674), 
        .B2(n12828), .ZN(n12675) );
  OAI21_X1 U14958 ( .B1(n12939), .B2(n12866), .A(n12675), .ZN(n12676) );
  AOI21_X1 U14959 ( .B1(n12879), .B2(n12831), .A(n12676), .ZN(n12677) );
  OAI21_X1 U14960 ( .B1(n12678), .B2(n12868), .A(n12677), .ZN(P3_U3208) );
  AND2_X1 U14961 ( .A1(n12680), .A2(n12679), .ZN(n12684) );
  OR2_X1 U14962 ( .A1(n12661), .A2(n12707), .ZN(n12699) );
  NAND3_X1 U14963 ( .A1(n12699), .A2(n12682), .A3(n12681), .ZN(n12683) );
  NAND3_X1 U14964 ( .A1(n12684), .A2(n12837), .A3(n12683), .ZN(n12688) );
  AOI22_X1 U14965 ( .A1(n12686), .A2(n12841), .B1(n12844), .B2(n12685), .ZN(
        n12687) );
  NAND2_X1 U14966 ( .A1(n12688), .A2(n12687), .ZN(n12882) );
  INV_X1 U14967 ( .A(n12882), .ZN(n12698) );
  INV_X1 U14968 ( .A(n12709), .ZN(n12691) );
  OAI21_X1 U14969 ( .B1(n12691), .B2(n12690), .A(n12689), .ZN(n12693) );
  NAND2_X1 U14970 ( .A1(n12693), .A2(n12692), .ZN(n12883) );
  AOI22_X1 U14971 ( .A1(n12868), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n12828), 
        .B2(n12694), .ZN(n12695) );
  OAI21_X1 U14972 ( .B1(n12943), .B2(n12866), .A(n12695), .ZN(n12696) );
  AOI21_X1 U14973 ( .B1(n12883), .B2(n12831), .A(n12696), .ZN(n12697) );
  OAI21_X1 U14974 ( .B1(n12698), .B2(n12868), .A(n12697), .ZN(P3_U3209) );
  INV_X1 U14975 ( .A(n12661), .ZN(n12701) );
  INV_X1 U14976 ( .A(n12707), .ZN(n12700) );
  OAI211_X1 U14977 ( .C1(n12701), .C2(n12700), .A(n12699), .B(n12837), .ZN(
        n12704) );
  NAND2_X1 U14978 ( .A1(n12702), .A2(n12844), .ZN(n12703) );
  OAI211_X1 U14979 ( .C1(n12705), .C2(n12862), .A(n12704), .B(n12703), .ZN(
        n12886) );
  INV_X1 U14980 ( .A(n12706), .ZN(n12947) );
  OR2_X1 U14981 ( .A1(n12708), .A2(n12707), .ZN(n12710) );
  AND2_X1 U14982 ( .A1(n12710), .A2(n12709), .ZN(n12887) );
  NAND2_X1 U14983 ( .A1(n12887), .A2(n12831), .ZN(n12713) );
  AOI22_X1 U14984 ( .A1(n12868), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n12828), 
        .B2(n12711), .ZN(n12712) );
  OAI211_X1 U14985 ( .C1(n12947), .C2(n12866), .A(n12713), .B(n12712), .ZN(
        n12714) );
  AOI21_X1 U14986 ( .B1(n12886), .B2(n12863), .A(n12714), .ZN(n12715) );
  INV_X1 U14987 ( .A(n12715), .ZN(P3_U3210) );
  XNOR2_X1 U14988 ( .A(n12717), .B(n12716), .ZN(n12718) );
  OAI222_X1 U14989 ( .A1(n12862), .A2(n12719), .B1(n12860), .B2(n12745), .C1(
        n12858), .C2(n12718), .ZN(n12890) );
  INV_X1 U14990 ( .A(n12890), .ZN(n12727) );
  XNOR2_X1 U14991 ( .A(n12721), .B(n12720), .ZN(n12891) );
  INV_X1 U14992 ( .A(n12722), .ZN(n12951) );
  AOI22_X1 U14993 ( .A1(n12868), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n12828), 
        .B2(n12723), .ZN(n12724) );
  OAI21_X1 U14994 ( .B1(n12951), .B2(n12866), .A(n12724), .ZN(n12725) );
  AOI21_X1 U14995 ( .B1(n12891), .B2(n12831), .A(n12725), .ZN(n12726) );
  OAI21_X1 U14996 ( .B1(n12727), .B2(n12868), .A(n12726), .ZN(P3_U3211) );
  INV_X1 U14997 ( .A(n12728), .ZN(n12729) );
  AOI21_X1 U14998 ( .B1(n12731), .B2(n12730), .A(n12729), .ZN(n12732) );
  OAI222_X1 U14999 ( .A1(n12862), .A2(n12734), .B1(n12860), .B2(n12733), .C1(
        n12858), .C2(n12732), .ZN(n12894) );
  INV_X1 U15000 ( .A(n12894), .ZN(n12741) );
  XNOR2_X1 U15001 ( .A(n12736), .B(n12735), .ZN(n12895) );
  AOI22_X1 U15002 ( .A1(n12868), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n12828), 
        .B2(n12737), .ZN(n12738) );
  OAI21_X1 U15003 ( .B1(n12954), .B2(n12866), .A(n12738), .ZN(n12739) );
  AOI21_X1 U15004 ( .B1(n12895), .B2(n12831), .A(n12739), .ZN(n12740) );
  OAI21_X1 U15005 ( .B1(n12741), .B2(n12868), .A(n12740), .ZN(P3_U3212) );
  XNOR2_X1 U15006 ( .A(n12742), .B(n12743), .ZN(n12744) );
  OAI222_X1 U15007 ( .A1(n12862), .A2(n12745), .B1(n12860), .B2(n12770), .C1(
        n12744), .C2(n12858), .ZN(n12898) );
  INV_X1 U15008 ( .A(n12898), .ZN(n12752) );
  XNOR2_X1 U15009 ( .A(n12746), .B(n8539), .ZN(n12899) );
  INV_X1 U15010 ( .A(n12747), .ZN(n12958) );
  AOI22_X1 U15011 ( .A1(n12868), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n12828), 
        .B2(n12748), .ZN(n12749) );
  OAI21_X1 U15012 ( .B1(n12958), .B2(n12866), .A(n12749), .ZN(n12750) );
  AOI21_X1 U15013 ( .B1(n12899), .B2(n12831), .A(n12750), .ZN(n12751) );
  OAI21_X1 U15014 ( .B1(n12752), .B2(n12868), .A(n12751), .ZN(P3_U3213) );
  OAI211_X1 U15015 ( .C1(n12754), .C2(n7446), .A(n12837), .B(n12753), .ZN(
        n12757) );
  AOI22_X1 U15016 ( .A1(n12755), .A2(n12841), .B1(n12844), .B2(n12781), .ZN(
        n12756) );
  NAND2_X1 U15017 ( .A1(n12757), .A2(n12756), .ZN(n12902) );
  INV_X1 U15018 ( .A(n12902), .ZN(n12764) );
  XNOR2_X1 U15019 ( .A(n12758), .B(n7446), .ZN(n12903) );
  NOR2_X1 U15020 ( .A1(n12962), .A2(n12866), .ZN(n12762) );
  OAI22_X1 U15021 ( .A1(n12863), .A2(n12760), .B1(n12759), .B2(n12864), .ZN(
        n12761) );
  AOI211_X1 U15022 ( .C1(n12903), .C2(n12831), .A(n12762), .B(n12761), .ZN(
        n12763) );
  OAI21_X1 U15023 ( .B1(n12764), .B2(n12868), .A(n12763), .ZN(P3_U3214) );
  INV_X1 U15024 ( .A(n12765), .ZN(n12766) );
  AOI21_X1 U15025 ( .B1(n12772), .B2(n12767), .A(n12766), .ZN(n12768) );
  OAI222_X1 U15026 ( .A1(n12862), .A2(n12770), .B1(n12860), .B2(n12769), .C1(
        n12858), .C2(n12768), .ZN(n12906) );
  INV_X1 U15027 ( .A(n12906), .ZN(n12779) );
  NAND2_X1 U15028 ( .A1(n12786), .A2(n12771), .ZN(n12773) );
  XNOR2_X1 U15029 ( .A(n12773), .B(n12772), .ZN(n12907) );
  NOR2_X1 U15030 ( .A1(n12966), .A2(n12866), .ZN(n12777) );
  INV_X1 U15031 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12775) );
  OAI22_X1 U15032 ( .A1(n12863), .A2(n12775), .B1(n12774), .B2(n12864), .ZN(
        n12776) );
  AOI211_X1 U15033 ( .C1(n12907), .C2(n12831), .A(n12777), .B(n12776), .ZN(
        n12778) );
  OAI21_X1 U15034 ( .B1(n12779), .B2(n12868), .A(n12778), .ZN(P3_U3215) );
  XNOR2_X1 U15035 ( .A(n12780), .B(n12788), .ZN(n12782) );
  AOI222_X1 U15036 ( .A1(n12837), .A2(n12782), .B1(n12781), .B2(n12841), .C1(
        n12805), .C2(n12844), .ZN(n12913) );
  OAI22_X1 U15037 ( .A1(n12863), .A2(n12784), .B1(n12783), .B2(n12864), .ZN(
        n12785) );
  AOI21_X1 U15038 ( .B1(n12910), .B2(n12796), .A(n12785), .ZN(n12790) );
  OAI21_X1 U15039 ( .B1(n12788), .B2(n12787), .A(n12786), .ZN(n12911) );
  NAND2_X1 U15040 ( .A1(n12911), .A2(n12831), .ZN(n12789) );
  OAI211_X1 U15041 ( .C1(n12913), .C2(n12833), .A(n12790), .B(n12789), .ZN(
        P3_U3216) );
  XNOR2_X1 U15042 ( .A(n6639), .B(n12798), .ZN(n12793) );
  AOI222_X1 U15043 ( .A1(n12837), .A2(n12793), .B1(n12820), .B2(n12844), .C1(
        n12792), .C2(n12841), .ZN(n12917) );
  OAI22_X1 U15044 ( .A1(n12863), .A2(n12536), .B1(n12794), .B2(n12864), .ZN(
        n12795) );
  AOI21_X1 U15045 ( .B1(n12914), .B2(n12796), .A(n12795), .ZN(n12801) );
  OAI21_X1 U15046 ( .B1(n12799), .B2(n12798), .A(n12797), .ZN(n12915) );
  NAND2_X1 U15047 ( .A1(n12915), .A2(n12831), .ZN(n12800) );
  OAI211_X1 U15048 ( .C1(n12917), .C2(n12868), .A(n12801), .B(n12800), .ZN(
        P3_U3217) );
  OAI211_X1 U15049 ( .C1(n12804), .C2(n12803), .A(n12802), .B(n12837), .ZN(
        n12807) );
  AOI22_X1 U15050 ( .A1(n12844), .A2(n12842), .B1(n12805), .B2(n12841), .ZN(
        n12806) );
  NAND2_X1 U15051 ( .A1(n12807), .A2(n12806), .ZN(n12918) );
  INV_X1 U15052 ( .A(n12918), .ZN(n12817) );
  OAI21_X1 U15053 ( .B1(n12810), .B2(n12809), .A(n12808), .ZN(n12919) );
  INV_X1 U15054 ( .A(n12811), .ZN(n12972) );
  INV_X1 U15055 ( .A(n12812), .ZN(n12813) );
  AOI22_X1 U15056 ( .A1(n12833), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n12828), 
        .B2(n12813), .ZN(n12814) );
  OAI21_X1 U15057 ( .B1(n12972), .B2(n12866), .A(n12814), .ZN(n12815) );
  AOI21_X1 U15058 ( .B1(n12919), .B2(n12831), .A(n12815), .ZN(n12816) );
  OAI21_X1 U15059 ( .B1(n12817), .B2(n12833), .A(n12816), .ZN(P3_U3218) );
  OAI211_X1 U15060 ( .C1(n12819), .C2(n12824), .A(n12818), .B(n12837), .ZN(
        n12823) );
  AOI22_X1 U15061 ( .A1(n12821), .A2(n12844), .B1(n12841), .B2(n12820), .ZN(
        n12822) );
  NAND2_X1 U15062 ( .A1(n12823), .A2(n12822), .ZN(n12921) );
  INV_X1 U15063 ( .A(n12921), .ZN(n12834) );
  XNOR2_X1 U15064 ( .A(n12825), .B(n12824), .ZN(n12922) );
  INV_X1 U15065 ( .A(n12826), .ZN(n12827) );
  AOI22_X1 U15066 ( .A1(n12833), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n12828), 
        .B2(n12827), .ZN(n12829) );
  OAI21_X1 U15067 ( .B1(n12976), .B2(n12866), .A(n12829), .ZN(n12830) );
  AOI21_X1 U15068 ( .B1(n12922), .B2(n12831), .A(n12830), .ZN(n12832) );
  OAI21_X1 U15069 ( .B1(n12834), .B2(n12833), .A(n12832), .ZN(P3_U3219) );
  XNOR2_X1 U15070 ( .A(n12836), .B(n12835), .ZN(n12926) );
  INV_X1 U15071 ( .A(n12926), .ZN(n12853) );
  OAI211_X1 U15072 ( .C1(n12840), .C2(n12839), .A(n12838), .B(n12837), .ZN(
        n12846) );
  AOI22_X1 U15073 ( .A1(n12844), .A2(n12843), .B1(n12842), .B2(n12841), .ZN(
        n12845) );
  NAND2_X1 U15074 ( .A1(n12846), .A2(n12845), .ZN(n12925) );
  INV_X1 U15075 ( .A(n12847), .ZN(n12980) );
  NOR2_X1 U15076 ( .A1(n12980), .A2(n12866), .ZN(n12851) );
  OAI22_X1 U15077 ( .A1(n12863), .A2(n12849), .B1(n12848), .B2(n12864), .ZN(
        n12850) );
  AOI211_X1 U15078 ( .C1(n12925), .C2(n12863), .A(n12851), .B(n12850), .ZN(
        n12852) );
  OAI21_X1 U15079 ( .B1(n12872), .B2(n12853), .A(n12852), .ZN(P3_U3220) );
  XNOR2_X1 U15080 ( .A(n12854), .B(n12855), .ZN(n14480) );
  INV_X1 U15081 ( .A(n14480), .ZN(n12871) );
  XNOR2_X1 U15082 ( .A(n12856), .B(n12855), .ZN(n12857) );
  OAI222_X1 U15083 ( .A1(n12862), .A2(n12861), .B1(n12860), .B2(n12859), .C1(
        n12858), .C2(n12857), .ZN(n14478) );
  NAND2_X1 U15084 ( .A1(n14478), .A2(n12863), .ZN(n12870) );
  OAI22_X1 U15085 ( .A1(n12866), .A2(n14477), .B1(n12865), .B2(n12864), .ZN(
        n12867) );
  AOI21_X1 U15086 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n12868), .A(n12867), 
        .ZN(n12869) );
  OAI211_X1 U15087 ( .C1(n12872), .C2(n12871), .A(n12870), .B(n12869), .ZN(
        P3_U3221) );
  MUX2_X1 U15088 ( .A(n14472), .B(n10396), .S(n15064), .Z(n12873) );
  OAI21_X1 U15089 ( .B1(n12931), .B2(n12928), .A(n12873), .ZN(P3_U3490) );
  OAI21_X1 U15090 ( .B1(n12935), .B2(n12928), .A(n12877), .ZN(P3_U3485) );
  AOI21_X1 U15091 ( .B1(n15049), .B2(n12879), .A(n12878), .ZN(n12936) );
  MUX2_X1 U15092 ( .A(n12880), .B(n12936), .S(n15066), .Z(n12881) );
  OAI21_X1 U15093 ( .B1(n12939), .B2(n12928), .A(n12881), .ZN(P3_U3484) );
  INV_X1 U15094 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12884) );
  AOI21_X1 U15095 ( .B1(n15049), .B2(n12883), .A(n12882), .ZN(n12940) );
  MUX2_X1 U15096 ( .A(n12884), .B(n12940), .S(n15066), .Z(n12885) );
  OAI21_X1 U15097 ( .B1(n12943), .B2(n12928), .A(n12885), .ZN(P3_U3483) );
  AOI21_X1 U15098 ( .B1(n12887), .B2(n15049), .A(n12886), .ZN(n12944) );
  MUX2_X1 U15099 ( .A(n12888), .B(n12944), .S(n15066), .Z(n12889) );
  OAI21_X1 U15100 ( .B1(n12947), .B2(n12928), .A(n12889), .ZN(P3_U3482) );
  INV_X1 U15101 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12892) );
  AOI21_X1 U15102 ( .B1(n15049), .B2(n12891), .A(n12890), .ZN(n12948) );
  MUX2_X1 U15103 ( .A(n12892), .B(n12948), .S(n15066), .Z(n12893) );
  OAI21_X1 U15104 ( .B1(n12951), .B2(n12928), .A(n12893), .ZN(P3_U3481) );
  AOI21_X1 U15105 ( .B1(n15049), .B2(n12895), .A(n12894), .ZN(n12952) );
  MUX2_X1 U15106 ( .A(n12896), .B(n12952), .S(n15066), .Z(n12897) );
  OAI21_X1 U15107 ( .B1(n12954), .B2(n12928), .A(n12897), .ZN(P3_U3480) );
  AOI21_X1 U15108 ( .B1(n12899), .B2(n15049), .A(n12898), .ZN(n12955) );
  MUX2_X1 U15109 ( .A(n12900), .B(n12955), .S(n15066), .Z(n12901) );
  OAI21_X1 U15110 ( .B1(n12958), .B2(n12928), .A(n12901), .ZN(P3_U3479) );
  INV_X1 U15111 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12904) );
  AOI21_X1 U15112 ( .B1(n15049), .B2(n12903), .A(n12902), .ZN(n12959) );
  MUX2_X1 U15113 ( .A(n12904), .B(n12959), .S(n15066), .Z(n12905) );
  OAI21_X1 U15114 ( .B1(n12928), .B2(n12962), .A(n12905), .ZN(P3_U3478) );
  AOI21_X1 U15115 ( .B1(n12907), .B2(n15049), .A(n12906), .ZN(n12963) );
  MUX2_X1 U15116 ( .A(n12908), .B(n12963), .S(n15066), .Z(n12909) );
  OAI21_X1 U15117 ( .B1(n12966), .B2(n12928), .A(n12909), .ZN(P3_U3477) );
  AOI22_X1 U15118 ( .A1(n12911), .A2(n15049), .B1(n15007), .B2(n12910), .ZN(
        n12912) );
  NAND2_X1 U15119 ( .A1(n12913), .A2(n12912), .ZN(n12967) );
  MUX2_X1 U15120 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12967), .S(n15066), .Z(
        P3_U3476) );
  AOI22_X1 U15121 ( .A1(n12915), .A2(n15049), .B1(n15007), .B2(n12914), .ZN(
        n12916) );
  NAND2_X1 U15122 ( .A1(n12917), .A2(n12916), .ZN(n12968) );
  MUX2_X1 U15123 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n12968), .S(n15066), .Z(
        P3_U3475) );
  AOI21_X1 U15124 ( .B1(n15049), .B2(n12919), .A(n12918), .ZN(n12969) );
  MUX2_X1 U15125 ( .A(n14460), .B(n12969), .S(n15066), .Z(n12920) );
  OAI21_X1 U15126 ( .B1(n12972), .B2(n12928), .A(n12920), .ZN(P3_U3474) );
  AOI21_X1 U15127 ( .B1(n15049), .B2(n12922), .A(n12921), .ZN(n12973) );
  MUX2_X1 U15128 ( .A(n12923), .B(n12973), .S(n15066), .Z(n12924) );
  OAI21_X1 U15129 ( .B1(n12928), .B2(n12976), .A(n12924), .ZN(P3_U3473) );
  AOI21_X1 U15130 ( .B1(n12926), .B2(n15049), .A(n12925), .ZN(n12977) );
  MUX2_X1 U15131 ( .A(n14983), .B(n12977), .S(n15066), .Z(n12927) );
  OAI21_X1 U15132 ( .B1(n12980), .B2(n12928), .A(n12927), .ZN(P3_U3472) );
  MUX2_X1 U15133 ( .A(n14472), .B(n12929), .S(n15050), .Z(n12930) );
  OAI21_X1 U15134 ( .B1(n12931), .B2(n12979), .A(n12930), .ZN(P3_U3458) );
  INV_X1 U15135 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12933) );
  MUX2_X1 U15136 ( .A(n12933), .B(n12932), .S(n15052), .Z(n12934) );
  OAI21_X1 U15137 ( .B1(n12935), .B2(n12979), .A(n12934), .ZN(P3_U3453) );
  INV_X1 U15138 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12937) );
  MUX2_X1 U15139 ( .A(n12937), .B(n12936), .S(n15052), .Z(n12938) );
  OAI21_X1 U15140 ( .B1(n12939), .B2(n12979), .A(n12938), .ZN(P3_U3452) );
  INV_X1 U15141 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12941) );
  MUX2_X1 U15142 ( .A(n12941), .B(n12940), .S(n15052), .Z(n12942) );
  OAI21_X1 U15143 ( .B1(n12943), .B2(n12979), .A(n12942), .ZN(P3_U3451) );
  INV_X1 U15144 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12945) );
  MUX2_X1 U15145 ( .A(n12945), .B(n12944), .S(n15052), .Z(n12946) );
  OAI21_X1 U15146 ( .B1(n12947), .B2(n12979), .A(n12946), .ZN(P3_U3450) );
  INV_X1 U15147 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12949) );
  MUX2_X1 U15148 ( .A(n12949), .B(n12948), .S(n15052), .Z(n12950) );
  OAI21_X1 U15149 ( .B1(n12951), .B2(n12979), .A(n12950), .ZN(P3_U3449) );
  MUX2_X1 U15150 ( .A(n15207), .B(n12952), .S(n15052), .Z(n12953) );
  OAI21_X1 U15151 ( .B1(n12954), .B2(n12979), .A(n12953), .ZN(P3_U3448) );
  MUX2_X1 U15152 ( .A(n12956), .B(n12955), .S(n15052), .Z(n12957) );
  OAI21_X1 U15153 ( .B1(n12958), .B2(n12979), .A(n12957), .ZN(P3_U3447) );
  INV_X1 U15154 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12960) );
  MUX2_X1 U15155 ( .A(n12960), .B(n12959), .S(n15052), .Z(n12961) );
  OAI21_X1 U15156 ( .B1(n12979), .B2(n12962), .A(n12961), .ZN(P3_U3446) );
  INV_X1 U15157 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12964) );
  MUX2_X1 U15158 ( .A(n12964), .B(n12963), .S(n15052), .Z(n12965) );
  OAI21_X1 U15159 ( .B1(n12966), .B2(n12979), .A(n12965), .ZN(P3_U3444) );
  MUX2_X1 U15160 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n12967), .S(n15052), .Z(
        P3_U3441) );
  MUX2_X1 U15161 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n12968), .S(n15052), .Z(
        P3_U3438) );
  INV_X1 U15162 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12970) );
  MUX2_X1 U15163 ( .A(n12970), .B(n12969), .S(n15052), .Z(n12971) );
  OAI21_X1 U15164 ( .B1(n12972), .B2(n12979), .A(n12971), .ZN(P3_U3435) );
  INV_X1 U15165 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12974) );
  MUX2_X1 U15166 ( .A(n12974), .B(n12973), .S(n15052), .Z(n12975) );
  OAI21_X1 U15167 ( .B1(n12979), .B2(n12976), .A(n12975), .ZN(P3_U3432) );
  MUX2_X1 U15168 ( .A(n15159), .B(n12977), .S(n15052), .Z(n12978) );
  OAI21_X1 U15169 ( .B1(n12980), .B2(n12979), .A(n12978), .ZN(P3_U3429) );
  MUX2_X1 U15170 ( .A(P3_D_REG_0__SCAN_IN), .B(n12982), .S(n12981), .Z(
        P3_U3376) );
  NAND2_X1 U15171 ( .A1(n12983), .A2(n14397), .ZN(n12988) );
  INV_X1 U15172 ( .A(n12984), .ZN(n12986) );
  OR4_X1 U15173 ( .A1(n12986), .A2(P3_IR_REG_30__SCAN_IN), .A3(n12985), .A4(
        P3_U3151), .ZN(n12987) );
  OAI211_X1 U15174 ( .C1(n12989), .C2(n12995), .A(n12988), .B(n12987), .ZN(
        P3_U3264) );
  INV_X1 U15175 ( .A(n12990), .ZN(n12991) );
  OAI222_X1 U15176 ( .A1(n12995), .A2(n12992), .B1(P3_U3151), .B2(n8187), .C1(
        n12997), .C2(n12991), .ZN(P3_U3266) );
  INV_X1 U15177 ( .A(n12993), .ZN(n12996) );
  OAI222_X1 U15178 ( .A1(n12997), .A2(n12996), .B1(n12995), .B2(n12994), .C1(
        P3_U3151), .C2(n8664), .ZN(P3_U3267) );
  XNOR2_X1 U15179 ( .A(n12999), .B(n12998), .ZN(n13005) );
  OAI22_X1 U15180 ( .A1(n13093), .A2(n13001), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13000), .ZN(n13003) );
  OAI22_X1 U15181 ( .A1(n13072), .A2(n13031), .B1(n13118), .B2(n13251), .ZN(
        n13002) );
  AOI211_X1 U15182 ( .C1(n13514), .C2(n13120), .A(n13003), .B(n13002), .ZN(
        n13004) );
  OAI21_X1 U15183 ( .B1(n13005), .B2(n13122), .A(n13004), .ZN(P2_U3186) );
  OAI21_X1 U15184 ( .B1(n13008), .B2(n13007), .A(n13006), .ZN(n13009) );
  NAND2_X1 U15185 ( .A1(n13009), .A2(n13098), .ZN(n13015) );
  INV_X1 U15186 ( .A(n13306), .ZN(n13013) );
  INV_X1 U15187 ( .A(n13118), .ZN(n13089) );
  AND2_X1 U15188 ( .A1(n13128), .A2(n13427), .ZN(n13010) );
  AOI21_X1 U15189 ( .B1(n13130), .B2(n13426), .A(n13010), .ZN(n13309) );
  INV_X1 U15190 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13011) );
  OAI22_X1 U15191 ( .A1(n13309), .A2(n13082), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13011), .ZN(n13012) );
  AOI21_X1 U15192 ( .B1(n13013), .B2(n13089), .A(n13012), .ZN(n13014) );
  OAI211_X1 U15193 ( .C1(n6914), .C2(n13077), .A(n13015), .B(n13014), .ZN(
        P2_U3188) );
  AOI21_X1 U15194 ( .B1(n13016), .B2(n13017), .A(n6565), .ZN(n13021) );
  AOI22_X1 U15195 ( .A1(n13131), .A2(n13427), .B1(n13426), .B2(n13132), .ZN(
        n13368) );
  NAND2_X1 U15196 ( .A1(n13089), .A2(n13372), .ZN(n13018) );
  NAND2_X1 U15197 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13210)
         );
  OAI211_X1 U15198 ( .C1(n13368), .C2(n13082), .A(n13018), .B(n13210), .ZN(
        n13019) );
  AOI21_X1 U15199 ( .B1(n13559), .B2(n13120), .A(n13019), .ZN(n13020) );
  OAI21_X1 U15200 ( .B1(n13021), .B2(n13122), .A(n13020), .ZN(P2_U3191) );
  XNOR2_X1 U15201 ( .A(n13023), .B(n13022), .ZN(n13028) );
  AOI22_X1 U15202 ( .A1(n13130), .A2(n13427), .B1(n13426), .B2(n13131), .ZN(
        n13340) );
  OAI22_X1 U15203 ( .A1(n13340), .A2(n13082), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13024), .ZN(n13026) );
  NOR2_X1 U15204 ( .A1(n6918), .A2(n13077), .ZN(n13025) );
  AOI211_X1 U15205 ( .C1(n13089), .C2(n13343), .A(n13026), .B(n13025), .ZN(
        n13027) );
  OAI21_X1 U15206 ( .B1(n13028), .B2(n13122), .A(n13027), .ZN(P2_U3195) );
  XNOR2_X1 U15207 ( .A(n13030), .B(n13029), .ZN(n13036) );
  OAI22_X1 U15208 ( .A1(n13032), .A2(n13464), .B1(n13031), .B2(n13462), .ZN(
        n13279) );
  AOI22_X1 U15209 ( .A1(n13116), .A2(n13279), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13033) );
  OAI21_X1 U15210 ( .B1(n13282), .B2(n13118), .A(n13033), .ZN(n13034) );
  AOI21_X1 U15211 ( .B1(n13525), .B2(n13120), .A(n13034), .ZN(n13035) );
  OAI21_X1 U15212 ( .B1(n13036), .B2(n13122), .A(n13035), .ZN(P2_U3197) );
  INV_X1 U15213 ( .A(n13038), .ZN(n13039) );
  AOI21_X1 U15214 ( .B1(n13040), .B2(n13037), .A(n13039), .ZN(n13045) );
  OAI21_X1 U15215 ( .B1(n13093), .B2(n13388), .A(n13041), .ZN(n13043) );
  OAI22_X1 U15216 ( .A1(n13072), .A2(n13461), .B1(n13118), .B2(n13431), .ZN(
        n13042) );
  AOI211_X1 U15217 ( .C1(n13577), .C2(n13120), .A(n13043), .B(n13042), .ZN(
        n13044) );
  OAI21_X1 U15218 ( .B1(n13045), .B2(n13122), .A(n13044), .ZN(P2_U3198) );
  OAI21_X1 U15219 ( .B1(n13048), .B2(n13047), .A(n13046), .ZN(n13049) );
  NAND2_X1 U15220 ( .A1(n13049), .A2(n13098), .ZN(n13056) );
  NAND2_X1 U15221 ( .A1(n13132), .A2(n13427), .ZN(n13051) );
  NAND2_X1 U15222 ( .A1(n13133), .A2(n13426), .ZN(n13050) );
  NAND2_X1 U15223 ( .A1(n13051), .A2(n13050), .ZN(n13413) );
  INV_X1 U15224 ( .A(n13052), .ZN(n13054) );
  NOR2_X1 U15225 ( .A1(n13118), .A2(n13406), .ZN(n13053) );
  AOI211_X1 U15226 ( .C1(n13116), .C2(n13413), .A(n13054), .B(n13053), .ZN(
        n13055) );
  OAI211_X1 U15227 ( .C1(n13405), .C2(n13077), .A(n13056), .B(n13055), .ZN(
        P2_U3200) );
  NAND2_X1 U15228 ( .A1(n13129), .A2(n13426), .ZN(n13058) );
  NAND2_X1 U15229 ( .A1(n13127), .A2(n13427), .ZN(n13057) );
  NAND2_X1 U15230 ( .A1(n13058), .A2(n13057), .ZN(n13531) );
  AOI22_X1 U15231 ( .A1(n13531), .A2(n13116), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13059) );
  OAI21_X1 U15232 ( .B1(n13291), .B2(n13118), .A(n13059), .ZN(n13065) );
  INV_X1 U15233 ( .A(n13060), .ZN(n13061) );
  AOI211_X1 U15234 ( .C1(n13063), .C2(n13062), .A(n13122), .B(n13061), .ZN(
        n13064) );
  AOI211_X1 U15235 ( .C1(n13529), .C2(n13120), .A(n13065), .B(n13064), .ZN(
        n13066) );
  INV_X1 U15236 ( .A(n13066), .ZN(P2_U3201) );
  OAI21_X1 U15237 ( .B1(n13069), .B2(n13068), .A(n13067), .ZN(n13070) );
  NAND2_X1 U15238 ( .A1(n13070), .A2(n13098), .ZN(n13076) );
  NOR2_X1 U15239 ( .A1(n13071), .A2(n13093), .ZN(n13074) );
  OAI22_X1 U15240 ( .A1(n13072), .A2(n13094), .B1(n13118), .B2(n13355), .ZN(
        n13073) );
  AOI211_X1 U15241 ( .C1(P2_REG3_REG_20__SCAN_IN), .C2(P2_U3088), .A(n13074), 
        .B(n13073), .ZN(n13075) );
  OAI211_X1 U15242 ( .C1(n8103), .C2(n13077), .A(n13076), .B(n13075), .ZN(
        P2_U3205) );
  XNOR2_X1 U15243 ( .A(n13078), .B(n13079), .ZN(n13086) );
  NOR2_X1 U15244 ( .A1(n13118), .A2(n13329), .ZN(n13084) );
  AND2_X1 U15245 ( .A1(n13353), .A2(n13426), .ZN(n13080) );
  AOI21_X1 U15246 ( .B1(n13129), .B2(n13427), .A(n13080), .ZN(n13320) );
  OAI22_X1 U15247 ( .A1(n13320), .A2(n13082), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13081), .ZN(n13083) );
  AOI211_X1 U15248 ( .C1(n13626), .C2(n13120), .A(n13084), .B(n13083), .ZN(
        n13085) );
  OAI21_X1 U15249 ( .B1(n13086), .B2(n13122), .A(n13085), .ZN(P2_U3207) );
  XNOR2_X1 U15250 ( .A(n13088), .B(n13087), .ZN(n13097) );
  AOI22_X1 U15251 ( .A1(n13090), .A2(n13428), .B1(n13089), .B2(n13396), .ZN(
        n13092) );
  OAI211_X1 U15252 ( .C1(n13094), .C2(n13093), .A(n13092), .B(n13091), .ZN(
        n13095) );
  AOI21_X1 U15253 ( .B1(n13562), .B2(n13120), .A(n13095), .ZN(n13096) );
  OAI21_X1 U15254 ( .B1(n13097), .B2(n13122), .A(n13096), .ZN(P2_U3210) );
  OAI211_X1 U15255 ( .C1(n13101), .C2(n13100), .A(n13099), .B(n13098), .ZN(
        n13109) );
  INV_X1 U15256 ( .A(n13102), .ZN(n13103) );
  AOI22_X1 U15257 ( .A1(n13116), .A2(n13103), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13108) );
  NAND2_X1 U15258 ( .A1(n13120), .A2(n13104), .ZN(n13107) );
  OR2_X1 U15259 ( .A1(n13118), .A2(n13105), .ZN(n13106) );
  NAND4_X1 U15260 ( .A1(n13109), .A2(n13108), .A3(n13107), .A4(n13106), .ZN(
        P2_U3211) );
  INV_X1 U15261 ( .A(n13110), .ZN(n13111) );
  AOI21_X1 U15262 ( .B1(n13113), .B2(n13112), .A(n13111), .ZN(n13123) );
  OAI22_X1 U15263 ( .A1(n13115), .A2(n13464), .B1(n13114), .B2(n13462), .ZN(
        n13264) );
  AOI22_X1 U15264 ( .A1(n13116), .A2(n13264), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13117) );
  OAI21_X1 U15265 ( .B1(n13267), .B2(n13118), .A(n13117), .ZN(n13119) );
  AOI21_X1 U15266 ( .B1(n13520), .B2(n13120), .A(n13119), .ZN(n13121) );
  OAI21_X1 U15267 ( .B1(n13123), .B2(n13122), .A(n13121), .ZN(P2_U3212) );
  MUX2_X1 U15268 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13218), .S(n6445), .Z(
        P2_U3562) );
  MUX2_X1 U15269 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13124), .S(n6445), .Z(
        P2_U3561) );
  MUX2_X1 U15270 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13125), .S(n6445), .Z(
        P2_U3560) );
  MUX2_X1 U15271 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13244), .S(n6445), .Z(
        P2_U3559) );
  MUX2_X1 U15272 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13126), .S(n6445), .Z(
        P2_U3558) );
  MUX2_X1 U15273 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13245), .S(n6445), .Z(
        P2_U3557) );
  MUX2_X1 U15274 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13127), .S(n6445), .Z(
        P2_U3556) );
  MUX2_X1 U15275 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13128), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15276 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13129), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15277 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13130), .S(n6445), .Z(
        P2_U3553) );
  MUX2_X1 U15278 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13353), .S(n6445), .Z(
        P2_U3552) );
  MUX2_X1 U15279 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13131), .S(n6445), .Z(
        P2_U3551) );
  MUX2_X1 U15280 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13386), .S(n6445), .Z(
        P2_U3550) );
  MUX2_X1 U15281 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13132), .S(n6445), .Z(
        P2_U3549) );
  MUX2_X1 U15282 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13428), .S(n6445), .Z(
        P2_U3548) );
  MUX2_X1 U15283 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13133), .S(n6445), .Z(
        P2_U3547) );
  MUX2_X1 U15284 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13425), .S(n6445), .Z(
        P2_U3546) );
  MUX2_X1 U15285 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13134), .S(n6445), .Z(
        P2_U3545) );
  MUX2_X1 U15286 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13135), .S(n6445), .Z(
        P2_U3544) );
  MUX2_X1 U15287 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13136), .S(n6445), .Z(
        P2_U3543) );
  MUX2_X1 U15288 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13137), .S(n6445), .Z(
        P2_U3542) );
  MUX2_X1 U15289 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13138), .S(n6445), .Z(
        P2_U3541) );
  MUX2_X1 U15290 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13139), .S(n6445), .Z(
        P2_U3540) );
  MUX2_X1 U15291 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13140), .S(n6445), .Z(
        P2_U3539) );
  MUX2_X1 U15292 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13141), .S(n6445), .Z(
        P2_U3538) );
  MUX2_X1 U15293 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13142), .S(n6445), .Z(
        P2_U3537) );
  MUX2_X1 U15294 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13143), .S(n6445), .Z(
        P2_U3536) );
  MUX2_X1 U15295 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13144), .S(n6445), .Z(
        P2_U3535) );
  MUX2_X1 U15296 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13145), .S(n6445), .Z(
        P2_U3534) );
  MUX2_X1 U15297 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13146), .S(n6445), .Z(
        P2_U3533) );
  MUX2_X1 U15298 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8917), .S(n6445), .Z(
        P2_U3532) );
  MUX2_X1 U15299 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n11881), .S(n6445), .Z(
        P2_U3531) );
  INV_X1 U15300 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n13148) );
  OAI21_X1 U15301 ( .B1(n13211), .B2(n13148), .A(n13147), .ZN(n13149) );
  AOI21_X1 U15302 ( .B1(n13153), .B2(n14822), .A(n13149), .ZN(n13159) );
  MUX2_X1 U15303 ( .A(n9441), .B(P2_REG1_REG_7__SCAN_IN), .S(n13153), .Z(
        n13150) );
  NAND3_X1 U15304 ( .A1(n14798), .A2(n13151), .A3(n13150), .ZN(n13152) );
  NAND3_X1 U15305 ( .A1(n14827), .A2(n13171), .A3(n13152), .ZN(n13158) );
  MUX2_X1 U15306 ( .A(n9469), .B(P2_REG2_REG_7__SCAN_IN), .S(n13153), .Z(
        n13154) );
  NAND3_X1 U15307 ( .A1(n14795), .A2(n13155), .A3(n13154), .ZN(n13156) );
  NAND3_X1 U15308 ( .A1(n14824), .A2(n13165), .A3(n13156), .ZN(n13157) );
  NAND3_X1 U15309 ( .A1(n13159), .A2(n13158), .A3(n13157), .ZN(P2_U3221) );
  INV_X1 U15310 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n13161) );
  OAI21_X1 U15311 ( .B1(n13211), .B2(n13161), .A(n13160), .ZN(n13162) );
  AOI21_X1 U15312 ( .B1(n13168), .B2(n14822), .A(n13162), .ZN(n13176) );
  MUX2_X1 U15313 ( .A(n10576), .B(P2_REG2_REG_8__SCAN_IN), .S(n13168), .Z(
        n13163) );
  NAND3_X1 U15314 ( .A1(n13165), .A2(n13164), .A3(n13163), .ZN(n13166) );
  NAND3_X1 U15315 ( .A1(n14824), .A2(n13167), .A3(n13166), .ZN(n13175) );
  MUX2_X1 U15316 ( .A(n9444), .B(P2_REG1_REG_8__SCAN_IN), .S(n13168), .Z(
        n13169) );
  NAND3_X1 U15317 ( .A1(n13171), .A2(n13170), .A3(n13169), .ZN(n13172) );
  NAND3_X1 U15318 ( .A1(n14827), .A2(n13173), .A3(n13172), .ZN(n13174) );
  NAND3_X1 U15319 ( .A1(n13176), .A2(n13175), .A3(n13174), .ZN(P2_U3222) );
  NOR3_X1 U15320 ( .A1(n14806), .A2(n13489), .A3(n13183), .ZN(n13180) );
  INV_X1 U15321 ( .A(n13177), .ZN(n13187) );
  NOR3_X1 U15322 ( .A1(n14812), .A2(n13178), .A3(n13187), .ZN(n13179) );
  OR3_X1 U15323 ( .A1(n14822), .A2(n13180), .A3(n13179), .ZN(n13185) );
  OAI21_X1 U15324 ( .B1(n13183), .B2(n13182), .A(n13181), .ZN(n13184) );
  AOI22_X1 U15325 ( .A1(n13185), .A2(n13186), .B1(n14824), .B2(n13184), .ZN(
        n13193) );
  NAND2_X1 U15326 ( .A1(n14820), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n13191) );
  NOR3_X1 U15327 ( .A1(n13187), .A2(n13186), .A3(P2_REG1_REG_9__SCAN_IN), .ZN(
        n13188) );
  OAI21_X1 U15328 ( .B1(n13189), .B2(n13188), .A(n14827), .ZN(n13190) );
  NAND4_X1 U15329 ( .A1(n13193), .A2(n13192), .A3(n13191), .A4(n13190), .ZN(
        P2_U3223) );
  NOR2_X1 U15330 ( .A1(n13195), .A2(n13194), .ZN(n13196) );
  XNOR2_X1 U15331 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13196), .ZN(n13204) );
  OR2_X1 U15332 ( .A1(n13198), .A2(n13197), .ZN(n13202) );
  NAND2_X1 U15333 ( .A1(n13200), .A2(n13199), .ZN(n13201) );
  NAND2_X1 U15334 ( .A1(n13202), .A2(n13201), .ZN(n13203) );
  XNOR2_X1 U15335 ( .A(n13203), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13205) );
  OAI22_X1 U15336 ( .A1(n13204), .A2(n14806), .B1(n13205), .B2(n14812), .ZN(
        n13209) );
  NAND2_X1 U15337 ( .A1(n13204), .A2(n14824), .ZN(n13207) );
  AOI21_X1 U15338 ( .B1(n13205), .B2(n14827), .A(n14822), .ZN(n13206) );
  NAND2_X1 U15339 ( .A1(n13207), .A2(n13206), .ZN(n13208) );
  MUX2_X1 U15340 ( .A(n13209), .B(n13208), .S(n6689), .Z(n13213) );
  OAI21_X1 U15341 ( .B1(n13211), .B2(n7516), .A(n13210), .ZN(n13212) );
  XNOR2_X1 U15342 ( .A(n13222), .B(n13607), .ZN(n13216) );
  NAND2_X1 U15343 ( .A1(n13216), .A2(n8927), .ZN(n13500) );
  NAND2_X1 U15344 ( .A1(n13218), .A2(n13217), .ZN(n13502) );
  NOR2_X1 U15345 ( .A1(n15079), .A2(n13502), .ZN(n13225) );
  AOI21_X1 U15346 ( .B1(n15079), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13225), 
        .ZN(n13220) );
  NAND2_X1 U15347 ( .A1(n13501), .A2(n13493), .ZN(n13219) );
  OAI211_X1 U15348 ( .C1(n13500), .C2(n13410), .A(n13220), .B(n13219), .ZN(
        P2_U3234) );
  AOI21_X1 U15349 ( .B1(n13221), .B2(n13610), .A(n13465), .ZN(n13223) );
  NAND2_X1 U15350 ( .A1(n13223), .A2(n13222), .ZN(n13503) );
  NOR2_X1 U15351 ( .A1(n13490), .A2(n13224), .ZN(n13226) );
  AOI211_X1 U15352 ( .C1(n13610), .C2(n13493), .A(n13226), .B(n13225), .ZN(
        n13227) );
  OAI21_X1 U15353 ( .B1(n13503), .B2(n13410), .A(n13227), .ZN(P2_U3235) );
  OAI211_X1 U15354 ( .C1(n13234), .C2(n13233), .A(n13232), .B(n13421), .ZN(
        n13237) );
  INV_X1 U15355 ( .A(n13235), .ZN(n13236) );
  OAI211_X1 U15356 ( .C1(n13613), .C2(n13250), .A(n8927), .B(n13238), .ZN(
        n13506) );
  OAI22_X1 U15357 ( .A1(n13506), .A2(n6689), .B1(n13487), .B2(n13239), .ZN(
        n13240) );
  OAI21_X1 U15358 ( .B1(n6649), .B2(n13240), .A(n13490), .ZN(n13242) );
  AOI22_X1 U15359 ( .A1(n13512), .A2(n13493), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n15079), .ZN(n13241) );
  OAI211_X1 U15360 ( .C1(n13474), .C2(n13508), .A(n13242), .B(n13241), .ZN(
        P2_U3237) );
  XNOR2_X1 U15361 ( .A(n13258), .B(n13243), .ZN(n13246) );
  AOI222_X1 U15362 ( .A1(n13421), .A2(n13246), .B1(n13245), .B2(n13426), .C1(
        n13244), .C2(n13427), .ZN(n13518) );
  NAND2_X1 U15363 ( .A1(n13514), .A2(n13247), .ZN(n13248) );
  NAND2_X1 U15364 ( .A1(n13248), .A2(n8927), .ZN(n13249) );
  NOR2_X1 U15365 ( .A1(n13250), .A2(n13249), .ZN(n13513) );
  OAI22_X1 U15366 ( .A1(n13490), .A2(n13252), .B1(n13251), .B2(n13487), .ZN(
        n13255) );
  NOR2_X1 U15367 ( .A1(n13253), .A2(n14839), .ZN(n13254) );
  AOI211_X1 U15368 ( .C1(n13513), .C2(n14833), .A(n13255), .B(n13254), .ZN(
        n13260) );
  NAND2_X1 U15369 ( .A1(n13258), .A2(n13257), .ZN(n13515) );
  NAND3_X1 U15370 ( .A1(n13256), .A2(n13515), .A3(n14842), .ZN(n13259) );
  OAI211_X1 U15371 ( .C1(n13518), .C2(n15079), .A(n13260), .B(n13259), .ZN(
        P2_U3238) );
  AOI211_X1 U15372 ( .C1(n13520), .C2(n13275), .A(n13262), .B(n13261), .ZN(
        n13519) );
  XNOR2_X1 U15373 ( .A(n13263), .B(n13269), .ZN(n13265) );
  AOI21_X1 U15374 ( .B1(n13265), .B2(n13421), .A(n13264), .ZN(n13521) );
  INV_X1 U15375 ( .A(n13521), .ZN(n13266) );
  AOI21_X1 U15376 ( .B1(n13519), .B2(n6688), .A(n13266), .ZN(n13274) );
  OAI22_X1 U15377 ( .A1(n13490), .A2(n13268), .B1(n13267), .B2(n13487), .ZN(
        n13272) );
  XNOR2_X1 U15378 ( .A(n13270), .B(n13269), .ZN(n13523) );
  NOR2_X1 U15379 ( .A1(n13523), .A2(n13474), .ZN(n13271) );
  AOI211_X1 U15380 ( .C1(n13493), .C2(n13520), .A(n13272), .B(n13271), .ZN(
        n13273) );
  OAI21_X1 U15381 ( .B1(n15079), .B2(n13274), .A(n13273), .ZN(P2_U3239) );
  INV_X1 U15382 ( .A(n13293), .ZN(n13277) );
  INV_X1 U15383 ( .A(n13275), .ZN(n13276) );
  AOI211_X1 U15384 ( .C1(n13525), .C2(n13277), .A(n13465), .B(n13276), .ZN(
        n13524) );
  XNOR2_X1 U15385 ( .A(n13278), .B(n13285), .ZN(n13280) );
  AOI21_X1 U15386 ( .B1(n13280), .B2(n13421), .A(n13279), .ZN(n13527) );
  INV_X1 U15387 ( .A(n13527), .ZN(n13281) );
  AOI21_X1 U15388 ( .B1(n13524), .B2(n13312), .A(n13281), .ZN(n13289) );
  OAI22_X1 U15389 ( .A1(n13490), .A2(n13283), .B1(n13282), .B2(n13487), .ZN(
        n13287) );
  XOR2_X1 U15390 ( .A(n13285), .B(n13284), .Z(n13528) );
  NOR2_X1 U15391 ( .A1(n13528), .A2(n13474), .ZN(n13286) );
  AOI211_X1 U15392 ( .C1(n13493), .C2(n13525), .A(n13287), .B(n13286), .ZN(
        n13288) );
  OAI21_X1 U15393 ( .B1(n15079), .B2(n13289), .A(n13288), .ZN(P2_U3240) );
  XNOR2_X1 U15394 ( .A(n13290), .B(n13295), .ZN(n13530) );
  OAI22_X1 U15395 ( .A1(n13490), .A2(n13292), .B1(n13291), .B2(n13487), .ZN(
        n13302) );
  AOI211_X1 U15396 ( .C1(n13529), .C2(n13304), .A(n13465), .B(n13293), .ZN(
        n13533) );
  INV_X1 U15397 ( .A(n13307), .ZN(n13297) );
  INV_X1 U15398 ( .A(n13294), .ZN(n13296) );
  OAI21_X1 U15399 ( .B1(n13297), .B2(n13296), .A(n13295), .ZN(n13299) );
  AOI21_X1 U15400 ( .B1(n13299), .B2(n13298), .A(n13459), .ZN(n13532) );
  AOI211_X1 U15401 ( .C1(n13533), .C2(n6688), .A(n13531), .B(n13532), .ZN(
        n13300) );
  NOR2_X1 U15402 ( .A1(n13300), .A2(n15079), .ZN(n13301) );
  AOI211_X1 U15403 ( .C1(n13493), .C2(n13529), .A(n13302), .B(n13301), .ZN(
        n13303) );
  OAI21_X1 U15404 ( .B1(n13474), .B2(n13530), .A(n13303), .ZN(P2_U3241) );
  INV_X1 U15405 ( .A(n13304), .ZN(n13305) );
  AOI211_X1 U15406 ( .C1(n13313), .C2(n13328), .A(n13465), .B(n13305), .ZN(
        n13537) );
  NOR2_X1 U15407 ( .A1(n13306), .A2(n13487), .ZN(n13311) );
  OAI211_X1 U15408 ( .C1(n13315), .C2(n13308), .A(n13307), .B(n13421), .ZN(
        n13310) );
  NAND2_X1 U15409 ( .A1(n13310), .A2(n13309), .ZN(n13538) );
  AOI211_X1 U15410 ( .C1(n13537), .C2(n13312), .A(n13311), .B(n13538), .ZN(
        n13318) );
  AOI22_X1 U15411 ( .A1(n13313), .A2(n13493), .B1(n15079), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n13317) );
  XNOR2_X1 U15412 ( .A(n13314), .B(n13315), .ZN(n13539) );
  NAND2_X1 U15413 ( .A1(n13539), .A2(n14842), .ZN(n13316) );
  OAI211_X1 U15414 ( .C1(n13318), .C2(n15079), .A(n13317), .B(n13316), .ZN(
        P2_U3242) );
  XNOR2_X1 U15415 ( .A(n13323), .B(n13319), .ZN(n13322) );
  INV_X1 U15416 ( .A(n13320), .ZN(n13321) );
  AOI21_X1 U15417 ( .B1(n13322), .B2(n13421), .A(n13321), .ZN(n13543) );
  NAND2_X1 U15418 ( .A1(n13324), .A2(n13323), .ZN(n13325) );
  NAND2_X1 U15419 ( .A1(n13326), .A2(n13325), .ZN(n13544) );
  INV_X1 U15420 ( .A(n13544), .ZN(n13334) );
  AOI21_X1 U15421 ( .B1(n13626), .B2(n6919), .A(n13465), .ZN(n13327) );
  NAND2_X1 U15422 ( .A1(n13328), .A2(n13327), .ZN(n13542) );
  INV_X1 U15423 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13330) );
  OAI22_X1 U15424 ( .A1(n13490), .A2(n13330), .B1(n13329), .B2(n13487), .ZN(
        n13331) );
  AOI21_X1 U15425 ( .B1(n13626), .B2(n13493), .A(n13331), .ZN(n13332) );
  OAI21_X1 U15426 ( .B1(n13542), .B2(n13410), .A(n13332), .ZN(n13333) );
  AOI21_X1 U15427 ( .B1(n13334), .B2(n14842), .A(n13333), .ZN(n13335) );
  OAI21_X1 U15428 ( .B1(n15079), .B2(n13543), .A(n13335), .ZN(P2_U3243) );
  XNOR2_X1 U15429 ( .A(n13336), .B(n13338), .ZN(n13551) );
  AND2_X1 U15430 ( .A1(n13351), .A2(n13352), .ZN(n13349) );
  NOR2_X1 U15431 ( .A1(n13349), .A2(n13337), .ZN(n13339) );
  XNOR2_X1 U15432 ( .A(n13339), .B(n13338), .ZN(n13341) );
  OAI21_X1 U15433 ( .B1(n13341), .B2(n13459), .A(n13340), .ZN(n13547) );
  NAND2_X1 U15434 ( .A1(n13547), .A2(n13490), .ZN(n13347) );
  AOI211_X1 U15435 ( .C1(n13549), .C2(n13359), .A(n13465), .B(n13342), .ZN(
        n13548) );
  INV_X1 U15436 ( .A(n13487), .ZN(n15071) );
  AOI22_X1 U15437 ( .A1(n15079), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13343), 
        .B2(n15071), .ZN(n13344) );
  OAI21_X1 U15438 ( .B1(n6918), .B2(n14839), .A(n13344), .ZN(n13345) );
  AOI21_X1 U15439 ( .B1(n13548), .B2(n14833), .A(n13345), .ZN(n13346) );
  OAI211_X1 U15440 ( .C1(n13551), .C2(n13474), .A(n13347), .B(n13346), .ZN(
        P2_U3244) );
  XNOR2_X1 U15441 ( .A(n13348), .B(n13352), .ZN(n13556) );
  INV_X1 U15442 ( .A(n13349), .ZN(n13350) );
  OAI21_X1 U15443 ( .B1(n13352), .B2(n13351), .A(n13350), .ZN(n13354) );
  AOI222_X1 U15444 ( .A1(n13421), .A2(n13354), .B1(n13353), .B2(n13427), .C1(
        n13386), .C2(n13426), .ZN(n13555) );
  INV_X1 U15445 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n13356) );
  OAI22_X1 U15446 ( .A1(n13490), .A2(n13356), .B1(n13355), .B2(n13487), .ZN(
        n13357) );
  AOI21_X1 U15447 ( .B1(n13553), .B2(n13493), .A(n13357), .ZN(n13362) );
  AOI21_X1 U15448 ( .B1(n13553), .B2(n13370), .A(n13465), .ZN(n13360) );
  AND2_X1 U15449 ( .A1(n13360), .A2(n13359), .ZN(n13552) );
  NAND2_X1 U15450 ( .A1(n13552), .A2(n14833), .ZN(n13361) );
  OAI211_X1 U15451 ( .C1(n13555), .C2(n15079), .A(n13362), .B(n13361), .ZN(
        n13363) );
  INV_X1 U15452 ( .A(n13363), .ZN(n13364) );
  OAI21_X1 U15453 ( .B1(n13474), .B2(n13556), .A(n13364), .ZN(P2_U3245) );
  XNOR2_X1 U15454 ( .A(n13365), .B(n13366), .ZN(n13561) );
  XOR2_X1 U15455 ( .A(n13367), .B(n13366), .Z(n13369) );
  OAI21_X1 U15456 ( .B1(n13369), .B2(n13459), .A(n13368), .ZN(n13557) );
  NAND2_X1 U15457 ( .A1(n13557), .A2(n13490), .ZN(n13378) );
  AOI21_X1 U15458 ( .B1(n13559), .B2(n13394), .A(n13465), .ZN(n13371) );
  AND2_X1 U15459 ( .A1(n13371), .A2(n13370), .ZN(n13558) );
  INV_X1 U15460 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13375) );
  NAND2_X1 U15461 ( .A1(n13559), .A2(n13493), .ZN(n13374) );
  NAND2_X1 U15462 ( .A1(n15071), .A2(n13372), .ZN(n13373) );
  OAI211_X1 U15463 ( .C1(n13490), .C2(n13375), .A(n13374), .B(n13373), .ZN(
        n13376) );
  AOI21_X1 U15464 ( .B1(n13558), .B2(n14833), .A(n13376), .ZN(n13377) );
  OAI211_X1 U15465 ( .C1(n13474), .C2(n13561), .A(n13378), .B(n13377), .ZN(
        P2_U3246) );
  NAND2_X1 U15466 ( .A1(n13379), .A2(n13380), .ZN(n13381) );
  NAND2_X1 U15467 ( .A1(n13382), .A2(n13381), .ZN(n13566) );
  NAND2_X1 U15468 ( .A1(n13566), .A2(n13383), .ZN(n13392) );
  XNOR2_X1 U15469 ( .A(n13385), .B(n13384), .ZN(n13390) );
  NAND2_X1 U15470 ( .A1(n13386), .A2(n13427), .ZN(n13387) );
  OAI21_X1 U15471 ( .B1(n13388), .B2(n13464), .A(n13387), .ZN(n13389) );
  AOI21_X1 U15472 ( .B1(n13390), .B2(n13421), .A(n13389), .ZN(n13391) );
  INV_X1 U15473 ( .A(n13393), .ZN(n13400) );
  AOI21_X1 U15474 ( .B1(n13562), .B2(n13404), .A(n13465), .ZN(n13395) );
  NAND2_X1 U15475 ( .A1(n13395), .A2(n13394), .ZN(n13563) );
  AOI22_X1 U15476 ( .A1(n15079), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13396), 
        .B2(n15071), .ZN(n13398) );
  NAND2_X1 U15477 ( .A1(n13562), .A2(n13493), .ZN(n13397) );
  OAI211_X1 U15478 ( .C1(n13563), .C2(n13410), .A(n13398), .B(n13397), .ZN(
        n13399) );
  AOI21_X1 U15479 ( .B1(n13566), .B2(n13400), .A(n13399), .ZN(n13401) );
  OAI21_X1 U15480 ( .B1(n13568), .B2(n15079), .A(n13401), .ZN(P2_U3247) );
  INV_X1 U15481 ( .A(n13411), .ZN(n13402) );
  XNOR2_X1 U15482 ( .A(n13403), .B(n13402), .ZN(n13569) );
  OAI211_X1 U15483 ( .C1(n13435), .C2(n13405), .A(n13404), .B(n8927), .ZN(
        n13570) );
  OAI22_X1 U15484 ( .A1(n13490), .A2(n13407), .B1(n13406), .B2(n13487), .ZN(
        n13408) );
  AOI21_X1 U15485 ( .B1(n13634), .B2(n13493), .A(n13408), .ZN(n13409) );
  OAI21_X1 U15486 ( .B1(n13570), .B2(n13410), .A(n13409), .ZN(n13416) );
  XNOR2_X1 U15487 ( .A(n13412), .B(n13411), .ZN(n13414) );
  AOI21_X1 U15488 ( .B1(n13414), .B2(n13421), .A(n13413), .ZN(n13571) );
  NOR2_X1 U15489 ( .A1(n13571), .A2(n15079), .ZN(n13415) );
  AOI211_X1 U15490 ( .C1(n14842), .C2(n13569), .A(n13416), .B(n13415), .ZN(
        n13417) );
  INV_X1 U15491 ( .A(n13417), .ZN(P2_U3248) );
  OAI21_X1 U15492 ( .B1(n13420), .B2(n13419), .A(n13418), .ZN(n13579) );
  OAI211_X1 U15493 ( .C1(n13424), .C2(n13423), .A(n13422), .B(n13421), .ZN(
        n13430) );
  AOI22_X1 U15494 ( .A1(n13428), .A2(n13427), .B1(n13426), .B2(n13425), .ZN(
        n13429) );
  NAND2_X1 U15495 ( .A1(n13430), .A2(n13429), .ZN(n13575) );
  NOR2_X1 U15496 ( .A1(n13487), .A2(n13431), .ZN(n13432) );
  OAI21_X1 U15497 ( .B1(n13575), .B2(n13432), .A(n13490), .ZN(n13439) );
  NAND2_X1 U15498 ( .A1(n13450), .A2(n13577), .ZN(n13433) );
  NAND2_X1 U15499 ( .A1(n13433), .A2(n8927), .ZN(n13434) );
  NOR2_X1 U15500 ( .A1(n13435), .A2(n13434), .ZN(n13576) );
  INV_X1 U15501 ( .A(n13577), .ZN(n13436) );
  OAI22_X1 U15502 ( .A1(n13436), .A2(n14839), .B1(n13490), .B2(n10410), .ZN(
        n13437) );
  AOI21_X1 U15503 ( .B1(n13576), .B2(n14833), .A(n13437), .ZN(n13438) );
  OAI211_X1 U15504 ( .C1(n13579), .C2(n13474), .A(n13439), .B(n13438), .ZN(
        P2_U3249) );
  XNOR2_X1 U15505 ( .A(n13441), .B(n13440), .ZN(n13443) );
  OAI21_X1 U15506 ( .B1(n13443), .B2(n13459), .A(n13442), .ZN(n13581) );
  NAND2_X1 U15507 ( .A1(n13581), .A2(n13490), .ZN(n13455) );
  OAI22_X1 U15508 ( .A1(n13490), .A2(n13445), .B1(n13444), .B2(n13487), .ZN(
        n13446) );
  AOI21_X1 U15509 ( .B1(n13580), .B2(n13493), .A(n13446), .ZN(n13454) );
  XNOR2_X1 U15510 ( .A(n13448), .B(n13447), .ZN(n13583) );
  NAND2_X1 U15511 ( .A1(n13583), .A2(n14842), .ZN(n13453) );
  AOI21_X1 U15512 ( .B1(n6929), .B2(n13580), .A(n13465), .ZN(n13451) );
  AND2_X1 U15513 ( .A1(n13451), .A2(n13450), .ZN(n13582) );
  NAND2_X1 U15514 ( .A1(n13582), .A2(n14833), .ZN(n13452) );
  NAND4_X1 U15515 ( .A1(n13455), .A2(n13454), .A3(n13453), .A4(n13452), .ZN(
        P2_U3250) );
  XOR2_X1 U15516 ( .A(n13456), .B(n13457), .Z(n13591) );
  XOR2_X1 U15517 ( .A(n13458), .B(n13457), .Z(n13460) );
  OAI222_X1 U15518 ( .A1(n13464), .A2(n13463), .B1(n13462), .B2(n13461), .C1(
        n13460), .C2(n13459), .ZN(n13587) );
  NAND2_X1 U15519 ( .A1(n13587), .A2(n13490), .ZN(n13473) );
  AOI211_X1 U15520 ( .C1(n13589), .C2(n13466), .A(n13465), .B(n13449), .ZN(
        n13588) );
  INV_X1 U15521 ( .A(n13467), .ZN(n13468) );
  AOI22_X1 U15522 ( .A1(n15079), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n13468), 
        .B2(n15071), .ZN(n13469) );
  OAI21_X1 U15523 ( .B1(n13470), .B2(n14839), .A(n13469), .ZN(n13471) );
  AOI21_X1 U15524 ( .B1(n13588), .B2(n14833), .A(n13471), .ZN(n13472) );
  OAI211_X1 U15525 ( .C1(n13591), .C2(n13474), .A(n13473), .B(n13472), .ZN(
        P2_U3251) );
  NAND2_X1 U15526 ( .A1(n13475), .A2(n13490), .ZN(n13485) );
  OAI22_X1 U15527 ( .A1(n13490), .A2(n13477), .B1(n13476), .B2(n13487), .ZN(
        n13478) );
  AOI21_X1 U15528 ( .B1(n13479), .B2(n13493), .A(n13478), .ZN(n13484) );
  NAND2_X1 U15529 ( .A1(n13480), .A2(n14842), .ZN(n13483) );
  NAND2_X1 U15530 ( .A1(n13481), .A2(n14833), .ZN(n13482) );
  NAND4_X1 U15531 ( .A1(n13485), .A2(n13484), .A3(n13483), .A4(n13482), .ZN(
        P2_U3255) );
  NAND2_X1 U15532 ( .A1(n13486), .A2(n13490), .ZN(n13499) );
  OAI22_X1 U15533 ( .A1(n13490), .A2(n13489), .B1(n13488), .B2(n13487), .ZN(
        n13491) );
  AOI21_X1 U15534 ( .B1(n13493), .B2(n13492), .A(n13491), .ZN(n13498) );
  NAND2_X1 U15535 ( .A1(n13494), .A2(n14842), .ZN(n13497) );
  NAND2_X1 U15536 ( .A1(n13495), .A2(n14833), .ZN(n13496) );
  NAND4_X1 U15537 ( .A1(n13499), .A2(n13498), .A3(n13497), .A4(n13496), .ZN(
        P2_U3256) );
  NAND2_X1 U15538 ( .A1(n13503), .A2(n13502), .ZN(n13608) );
  MUX2_X1 U15539 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13608), .S(n14885), .Z(
        n13504) );
  AOI21_X1 U15540 ( .B1(n13596), .B2(n13610), .A(n13504), .ZN(n13505) );
  INV_X1 U15541 ( .A(n13505), .ZN(P2_U3529) );
  OAI21_X1 U15542 ( .B1(n13508), .B2(n13603), .A(n13507), .ZN(n13612) );
  AOI21_X1 U15543 ( .B1(n14873), .B2(n13514), .A(n13513), .ZN(n13517) );
  NAND3_X1 U15544 ( .A1(n13256), .A2(n13584), .A3(n13515), .ZN(n13516) );
  NAND3_X1 U15545 ( .A1(n13518), .A2(n13517), .A3(n13516), .ZN(n13614) );
  MUX2_X1 U15546 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13614), .S(n14885), .Z(
        P2_U3526) );
  AOI21_X1 U15547 ( .B1(n14873), .B2(n13520), .A(n13519), .ZN(n13522) );
  OAI211_X1 U15548 ( .C1(n13603), .C2(n13523), .A(n13522), .B(n13521), .ZN(
        n13615) );
  MUX2_X1 U15549 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13615), .S(n14885), .Z(
        P2_U3525) );
  AOI21_X1 U15550 ( .B1(n14873), .B2(n13525), .A(n13524), .ZN(n13526) );
  OAI211_X1 U15551 ( .C1(n13528), .C2(n13603), .A(n13527), .B(n13526), .ZN(
        n13616) );
  MUX2_X1 U15552 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13616), .S(n14885), .Z(
        P2_U3524) );
  INV_X1 U15553 ( .A(n13529), .ZN(n13620) );
  NOR2_X1 U15554 ( .A1(n13530), .A2(n13603), .ZN(n13534) );
  NOR4_X1 U15555 ( .A1(n13534), .A2(n13533), .A3(n13532), .A4(n13531), .ZN(
        n13617) );
  MUX2_X1 U15556 ( .A(n13535), .B(n13617), .S(n14885), .Z(n13536) );
  OAI21_X1 U15557 ( .B1(n13620), .B2(n8170), .A(n13536), .ZN(P2_U3523) );
  AOI211_X1 U15558 ( .C1(n13539), .C2(n13584), .A(n13538), .B(n13537), .ZN(
        n13621) );
  MUX2_X1 U15559 ( .A(n13540), .B(n13621), .S(n14885), .Z(n13541) );
  OAI21_X1 U15560 ( .B1(n6914), .B2(n8170), .A(n13541), .ZN(P2_U3522) );
  OAI211_X1 U15561 ( .C1(n13544), .C2(n13603), .A(n13543), .B(n13542), .ZN(
        n13624) );
  MUX2_X1 U15562 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13624), .S(n14885), .Z(
        n13545) );
  AOI21_X1 U15563 ( .B1(n13596), .B2(n13626), .A(n13545), .ZN(n13546) );
  INV_X1 U15564 ( .A(n13546), .ZN(P2_U3521) );
  AOI211_X1 U15565 ( .C1(n14873), .C2(n13549), .A(n13548), .B(n13547), .ZN(
        n13550) );
  OAI21_X1 U15566 ( .B1(n13603), .B2(n13551), .A(n13550), .ZN(n13628) );
  MUX2_X1 U15567 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13628), .S(n14885), .Z(
        P2_U3520) );
  AOI21_X1 U15568 ( .B1(n14873), .B2(n13553), .A(n13552), .ZN(n13554) );
  OAI211_X1 U15569 ( .C1(n13603), .C2(n13556), .A(n13555), .B(n13554), .ZN(
        n13629) );
  MUX2_X1 U15570 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13629), .S(n14885), .Z(
        P2_U3519) );
  AOI211_X1 U15571 ( .C1(n14873), .C2(n13559), .A(n13558), .B(n13557), .ZN(
        n13560) );
  OAI21_X1 U15572 ( .B1(n13603), .B2(n13561), .A(n13560), .ZN(n13630) );
  MUX2_X1 U15573 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13630), .S(n14885), .Z(
        P2_U3518) );
  INV_X1 U15574 ( .A(n13562), .ZN(n13564) );
  OAI21_X1 U15575 ( .B1(n13564), .B2(n14864), .A(n13563), .ZN(n13565) );
  AOI21_X1 U15576 ( .B1(n13566), .B2(n14869), .A(n13565), .ZN(n13567) );
  NAND2_X1 U15577 ( .A1(n13568), .A2(n13567), .ZN(n13631) );
  MUX2_X1 U15578 ( .A(n13631), .B(P2_REG1_REG_18__SCAN_IN), .S(n14883), .Z(
        P2_U3517) );
  NAND2_X1 U15579 ( .A1(n13569), .A2(n13584), .ZN(n13572) );
  NAND3_X1 U15580 ( .A1(n13572), .A2(n13571), .A3(n13570), .ZN(n13632) );
  MUX2_X1 U15581 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13632), .S(n14885), .Z(
        n13573) );
  AOI21_X1 U15582 ( .B1(n13596), .B2(n13634), .A(n13573), .ZN(n13574) );
  INV_X1 U15583 ( .A(n13574), .ZN(P2_U3516) );
  AOI211_X1 U15584 ( .C1(n14873), .C2(n13577), .A(n13576), .B(n13575), .ZN(
        n13578) );
  OAI21_X1 U15585 ( .B1(n13603), .B2(n13579), .A(n13578), .ZN(n13636) );
  MUX2_X1 U15586 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13636), .S(n14885), .Z(
        P2_U3515) );
  INV_X1 U15587 ( .A(n13580), .ZN(n13641) );
  AOI211_X1 U15588 ( .C1(n13584), .C2(n13583), .A(n13582), .B(n13581), .ZN(
        n13637) );
  MUX2_X1 U15589 ( .A(n13585), .B(n13637), .S(n14885), .Z(n13586) );
  OAI21_X1 U15590 ( .B1(n13641), .B2(n8170), .A(n13586), .ZN(P2_U3514) );
  AOI211_X1 U15591 ( .C1(n14873), .C2(n13589), .A(n13588), .B(n13587), .ZN(
        n13590) );
  OAI21_X1 U15592 ( .B1(n13603), .B2(n13591), .A(n13590), .ZN(n13642) );
  MUX2_X1 U15593 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13642), .S(n14885), .Z(
        P2_U3513) );
  OAI211_X1 U15594 ( .C1(n13603), .C2(n13594), .A(n13593), .B(n13592), .ZN(
        n13643) );
  MUX2_X1 U15595 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n13643), .S(n14885), .Z(
        n13595) );
  AOI21_X1 U15596 ( .B1(n13596), .B2(n13645), .A(n13595), .ZN(n13597) );
  INV_X1 U15597 ( .A(n13597), .ZN(P2_U3512) );
  AOI211_X1 U15598 ( .C1(n14873), .C2(n13600), .A(n13599), .B(n13598), .ZN(
        n13601) );
  OAI21_X1 U15599 ( .B1(n13603), .B2(n13602), .A(n13601), .ZN(n13648) );
  MUX2_X1 U15600 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n13648), .S(n14885), .Z(
        P2_U3510) );
  MUX2_X1 U15601 ( .A(n13604), .B(P2_REG0_REG_31__SCAN_IN), .S(n14879), .Z(
        n13605) );
  INV_X1 U15602 ( .A(n13605), .ZN(n13606) );
  OAI21_X1 U15603 ( .B1(n13607), .B2(n13640), .A(n13606), .ZN(P2_U3498) );
  MUX2_X1 U15604 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13608), .S(n14880), .Z(
        n13609) );
  AOI21_X1 U15605 ( .B1(n13646), .B2(n13610), .A(n13609), .ZN(n13611) );
  INV_X1 U15606 ( .A(n13611), .ZN(P2_U3497) );
  MUX2_X1 U15607 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13614), .S(n14880), .Z(
        P2_U3494) );
  MUX2_X1 U15608 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13615), .S(n14880), .Z(
        P2_U3493) );
  MUX2_X1 U15609 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13616), .S(n14880), .Z(
        P2_U3492) );
  INV_X1 U15610 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n13618) );
  MUX2_X1 U15611 ( .A(n13618), .B(n13617), .S(n14880), .Z(n13619) );
  OAI21_X1 U15612 ( .B1(n13620), .B2(n13640), .A(n13619), .ZN(P2_U3491) );
  INV_X1 U15613 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n13622) );
  MUX2_X1 U15614 ( .A(n13622), .B(n13621), .S(n14880), .Z(n13623) );
  OAI21_X1 U15615 ( .B1(n6914), .B2(n13640), .A(n13623), .ZN(P2_U3490) );
  MUX2_X1 U15616 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13624), .S(n14880), .Z(
        n13625) );
  AOI21_X1 U15617 ( .B1(n13646), .B2(n13626), .A(n13625), .ZN(n13627) );
  INV_X1 U15618 ( .A(n13627), .ZN(P2_U3489) );
  MUX2_X1 U15619 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13628), .S(n14880), .Z(
        P2_U3488) );
  MUX2_X1 U15620 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13629), .S(n14880), .Z(
        P2_U3487) );
  MUX2_X1 U15621 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13630), .S(n14880), .Z(
        P2_U3486) );
  MUX2_X1 U15622 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13631), .S(n14880), .Z(
        P2_U3484) );
  MUX2_X1 U15623 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13632), .S(n14880), .Z(
        n13633) );
  AOI21_X1 U15624 ( .B1(n13646), .B2(n13634), .A(n13633), .ZN(n13635) );
  INV_X1 U15625 ( .A(n13635), .ZN(P2_U3481) );
  MUX2_X1 U15626 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13636), .S(n14880), .Z(
        P2_U3478) );
  MUX2_X1 U15627 ( .A(n13638), .B(n13637), .S(n14880), .Z(n13639) );
  OAI21_X1 U15628 ( .B1(n13641), .B2(n13640), .A(n13639), .ZN(P2_U3475) );
  MUX2_X1 U15629 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13642), .S(n14880), .Z(
        P2_U3472) );
  MUX2_X1 U15630 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n13643), .S(n14880), .Z(
        n13644) );
  AOI21_X1 U15631 ( .B1(n13646), .B2(n13645), .A(n13644), .ZN(n13647) );
  INV_X1 U15632 ( .A(n13647), .ZN(P2_U3469) );
  MUX2_X1 U15633 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n13648), .S(n14880), .Z(
        P2_U3463) );
  NAND3_X1 U15634 ( .A1(n13649), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13651) );
  OAI22_X1 U15635 ( .A1(n13652), .A2(n13651), .B1(n13650), .B2(n13671), .ZN(
        n13653) );
  AOI21_X1 U15636 ( .B1(n14254), .B2(n13668), .A(n13653), .ZN(n13654) );
  INV_X1 U15637 ( .A(n13654), .ZN(P2_U3296) );
  NAND2_X1 U15638 ( .A1(n14261), .A2(n13668), .ZN(n13656) );
  OAI211_X1 U15639 ( .C1(n13657), .C2(n13671), .A(n13656), .B(n13655), .ZN(
        P2_U3299) );
  OAI222_X1 U15640 ( .A1(n13671), .A2(n13660), .B1(n13666), .B2(n13659), .C1(
        n13658), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U15641 ( .A(n13661), .ZN(n14266) );
  OAI222_X1 U15642 ( .A1(P2_U3088), .A2(n13663), .B1(n13666), .B2(n14266), 
        .C1(n13662), .C2(n13671), .ZN(P2_U3301) );
  INV_X1 U15643 ( .A(n13664), .ZN(n14269) );
  OAI222_X1 U15644 ( .A1(n13671), .A2(n13667), .B1(n13666), .B2(n14269), .C1(
        P2_U3088), .C2(n13665), .ZN(P2_U3302) );
  NAND2_X1 U15645 ( .A1(n14273), .A2(n13668), .ZN(n13670) );
  OAI211_X1 U15646 ( .C1(n13672), .C2(n13671), .A(n13670), .B(n13669), .ZN(
        P2_U3304) );
  MUX2_X1 U15647 ( .A(n13674), .B(n13673), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3327) );
  XOR2_X1 U15648 ( .A(n13676), .B(n13675), .Z(n13682) );
  OAI22_X1 U15649 ( .A1(n14503), .A2(n14139), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13677), .ZN(n13680) );
  INV_X1 U15650 ( .A(n13948), .ZN(n13678) );
  OAI22_X1 U15651 ( .A1(n14502), .A2(n14138), .B1(n14628), .B2(n13678), .ZN(
        n13679) );
  AOI211_X1 U15652 ( .C1(n14142), .C2(n14525), .A(n13680), .B(n13679), .ZN(
        n13681) );
  OAI21_X1 U15653 ( .B1(n13682), .B2(n14620), .A(n13681), .ZN(P1_U3214) );
  XOR2_X1 U15654 ( .A(n13684), .B(n13683), .Z(n13690) );
  INV_X1 U15655 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13685) );
  OAI22_X1 U15656 ( .A1(n14184), .A2(n14503), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13685), .ZN(n13688) );
  INV_X1 U15657 ( .A(n13686), .ZN(n14018) );
  INV_X1 U15658 ( .A(n14154), .ZN(n13987) );
  OAI22_X1 U15659 ( .A1(n14018), .A2(n14628), .B1(n13987), .B2(n14502), .ZN(
        n13687) );
  AOI211_X1 U15660 ( .C1(n14175), .C2(n14525), .A(n13688), .B(n13687), .ZN(
        n13689) );
  OAI21_X1 U15661 ( .B1(n13690), .B2(n14620), .A(n13689), .ZN(P1_U3216) );
  AOI21_X1 U15662 ( .B1(n13692), .B2(n13691), .A(n14620), .ZN(n13694) );
  NAND2_X1 U15663 ( .A1(n13694), .A2(n13693), .ZN(n13699) );
  NOR2_X1 U15664 ( .A1(n13695), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13863) );
  INV_X1 U15665 ( .A(n14074), .ZN(n13696) );
  OAI22_X1 U15666 ( .A1(n14503), .A2(n14202), .B1(n14628), .B2(n13696), .ZN(
        n13697) );
  AOI211_X1 U15667 ( .C1(n13746), .C2(n13899), .A(n13863), .B(n13697), .ZN(
        n13698) );
  OAI211_X1 U15668 ( .C1(n6952), .C2(n14500), .A(n13699), .B(n13698), .ZN(
        P1_U3219) );
  INV_X1 U15669 ( .A(n13700), .ZN(n13701) );
  AOI21_X1 U15670 ( .B1(n13703), .B2(n13702), .A(n13701), .ZN(n13707) );
  OAI22_X1 U15671 ( .A1(n14184), .A2(n14502), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15206), .ZN(n13705) );
  OAI22_X1 U15672 ( .A1(n14503), .A2(n14203), .B1(n14628), .B2(n14043), .ZN(
        n13704) );
  AOI211_X1 U15673 ( .C1(n14187), .C2(n14525), .A(n13705), .B(n13704), .ZN(
        n13706) );
  OAI21_X1 U15674 ( .B1(n13707), .B2(n14620), .A(n13706), .ZN(P1_U3223) );
  INV_X1 U15675 ( .A(n13708), .ZN(n13709) );
  AOI211_X1 U15676 ( .C1(n13711), .C2(n13710), .A(n14620), .B(n13709), .ZN(
        n13717) );
  INV_X1 U15677 ( .A(n13712), .ZN(n14407) );
  AOI22_X1 U15678 ( .A1(n13746), .A2(n14558), .B1(P1_REG3_REG_12__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13715) );
  INV_X1 U15679 ( .A(n14503), .ZN(n13800) );
  AOI22_X1 U15680 ( .A1(n13800), .A2(n14404), .B1(n13713), .B2(n13798), .ZN(
        n13714) );
  OAI211_X1 U15681 ( .C1(n14407), .C2(n14500), .A(n13715), .B(n13714), .ZN(
        n13716) );
  OR2_X1 U15682 ( .A1(n13717), .A2(n13716), .ZN(P1_U3224) );
  XOR2_X1 U15683 ( .A(n13719), .B(n13718), .Z(n13725) );
  OAI22_X1 U15684 ( .A1(n14503), .A2(n13987), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13720), .ZN(n13723) );
  INV_X1 U15685 ( .A(n13984), .ZN(n13721) );
  OAI22_X1 U15686 ( .A1(n14502), .A2(n14139), .B1(n14628), .B2(n13721), .ZN(
        n13722) );
  AOI211_X1 U15687 ( .C1(n13983), .C2(n14525), .A(n13723), .B(n13722), .ZN(
        n13724) );
  OAI21_X1 U15688 ( .B1(n13725), .B2(n14620), .A(n13724), .ZN(P1_U3225) );
  INV_X1 U15689 ( .A(n13727), .ZN(n13728) );
  AOI21_X1 U15690 ( .B1(n13729), .B2(n13726), .A(n13728), .ZN(n13737) );
  NAND2_X1 U15691 ( .A1(n13798), .A2(n13730), .ZN(n13732) );
  OAI211_X1 U15692 ( .C1(n13734), .C2(n13733), .A(n13732), .B(n13731), .ZN(
        n13735) );
  AOI21_X1 U15693 ( .B1(n14227), .B2(n14525), .A(n13735), .ZN(n13736) );
  OAI21_X1 U15694 ( .B1(n13737), .B2(n14620), .A(n13736), .ZN(P1_U3226) );
  OAI21_X1 U15695 ( .B1(n13740), .B2(n13739), .A(n13738), .ZN(n13741) );
  NAND2_X1 U15696 ( .A1(n13741), .A2(n14527), .ZN(n13748) );
  INV_X1 U15697 ( .A(n13742), .ZN(n13745) );
  OAI22_X1 U15698 ( .A1(n14503), .A2(n13802), .B1(n14628), .B2(n13743), .ZN(
        n13744) );
  AOI211_X1 U15699 ( .C1(n13746), .C2(n14218), .A(n13745), .B(n13744), .ZN(
        n13747) );
  OAI211_X1 U15700 ( .C1(n14221), .C2(n14500), .A(n13748), .B(n13747), .ZN(
        P1_U3228) );
  XOR2_X1 U15701 ( .A(n13750), .B(n13749), .Z(n13756) );
  INV_X1 U15702 ( .A(n13888), .ZN(n14167) );
  OAI22_X1 U15703 ( .A1(n14167), .A2(n14503), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13751), .ZN(n13754) );
  INV_X1 U15704 ( .A(n14001), .ZN(n13752) );
  OAI22_X1 U15705 ( .A1(n14502), .A2(n14166), .B1(n14628), .B2(n13752), .ZN(
        n13753) );
  AOI211_X1 U15706 ( .C1(n14170), .C2(n14525), .A(n13754), .B(n13753), .ZN(
        n13755) );
  OAI21_X1 U15707 ( .B1(n13756), .B2(n14620), .A(n13755), .ZN(P1_U3229) );
  OAI211_X1 U15708 ( .C1(n13759), .C2(n13758), .A(n13757), .B(n14527), .ZN(
        n13765) );
  OAI22_X1 U15709 ( .A1(n13770), .A2(n14502), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13760), .ZN(n13763) );
  INV_X1 U15710 ( .A(n14060), .ZN(n13761) );
  OAI22_X1 U15711 ( .A1(n14503), .A2(n14211), .B1(n14628), .B2(n13761), .ZN(
        n13762) );
  NOR2_X1 U15712 ( .A1(n13763), .A2(n13762), .ZN(n13764) );
  OAI211_X1 U15713 ( .C1(n14197), .C2(n14500), .A(n13765), .B(n13764), .ZN(
        P1_U3233) );
  OAI21_X1 U15714 ( .B1(n13768), .B2(n13767), .A(n13766), .ZN(n13769) );
  NAND2_X1 U15715 ( .A1(n13769), .A2(n14527), .ZN(n13774) );
  OAI22_X1 U15716 ( .A1(n14167), .A2(n14420), .B1(n13770), .B2(n14209), .ZN(
        n14034) );
  INV_X1 U15717 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13771) );
  OAI22_X1 U15718 ( .A1(n14032), .A2(n14628), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13771), .ZN(n13772) );
  AOI21_X1 U15719 ( .B1(n14034), .B2(n14625), .A(n13772), .ZN(n13773) );
  OAI211_X1 U15720 ( .C1(n14500), .C2(n13775), .A(n13774), .B(n13773), .ZN(
        P1_U3235) );
  XOR2_X1 U15721 ( .A(n13777), .B(n13776), .Z(n13782) );
  AOI22_X1 U15722 ( .A1(n13800), .A2(n14093), .B1(n14089), .B2(n13798), .ZN(
        n13779) );
  OAI211_X1 U15723 ( .C1(n14211), .C2(n14502), .A(n13779), .B(n13778), .ZN(
        n13780) );
  AOI21_X1 U15724 ( .B1(n14214), .B2(n14525), .A(n13780), .ZN(n13781) );
  OAI21_X1 U15725 ( .B1(n13782), .B2(n14620), .A(n13781), .ZN(P1_U3238) );
  XOR2_X1 U15726 ( .A(n13784), .B(n13783), .Z(n13790) );
  OAI22_X1 U15727 ( .A1(n14503), .A2(n14166), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13785), .ZN(n13788) );
  INV_X1 U15728 ( .A(n13786), .ZN(n13963) );
  OAI22_X1 U15729 ( .A1(n14502), .A2(n14147), .B1(n14628), .B2(n13963), .ZN(
        n13787) );
  AOI211_X1 U15730 ( .C1(n14150), .C2(n14525), .A(n13788), .B(n13787), .ZN(
        n13789) );
  OAI21_X1 U15731 ( .B1(n13790), .B2(n14620), .A(n13789), .ZN(P1_U3240) );
  INV_X1 U15732 ( .A(n13791), .ZN(n13792) );
  NAND2_X1 U15733 ( .A1(n13793), .A2(n13792), .ZN(n13797) );
  XNOR2_X1 U15734 ( .A(n13795), .B(n13794), .ZN(n13796) );
  XNOR2_X1 U15735 ( .A(n13797), .B(n13796), .ZN(n13806) );
  AOI22_X1 U15736 ( .A1(n13800), .A2(n14548), .B1(n13799), .B2(n13798), .ZN(
        n13801) );
  NAND2_X1 U15737 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14672)
         );
  OAI211_X1 U15738 ( .C1(n13802), .C2(n14502), .A(n13801), .B(n14672), .ZN(
        n13803) );
  AOI21_X1 U15739 ( .B1(n13804), .B2(n14525), .A(n13803), .ZN(n13805) );
  OAI21_X1 U15740 ( .B1(n13806), .B2(n14620), .A(n13805), .ZN(P1_U3241) );
  MUX2_X1 U15741 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13807), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15742 ( .A(n13912), .B(P1_DATAO_REG_30__SCAN_IN), .S(n13817), .Z(
        P1_U3590) );
  MUX2_X1 U15743 ( .A(n13928), .B(P1_DATAO_REG_29__SCAN_IN), .S(n13817), .Z(
        P1_U3589) );
  MUX2_X1 U15744 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14120), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15745 ( .A(n13967), .B(P1_DATAO_REG_27__SCAN_IN), .S(n13817), .Z(
        P1_U3587) );
  MUX2_X1 U15746 ( .A(n14155), .B(P1_DATAO_REG_26__SCAN_IN), .S(n13817), .Z(
        P1_U3586) );
  MUX2_X1 U15747 ( .A(n14004), .B(P1_DATAO_REG_25__SCAN_IN), .S(n13817), .Z(
        P1_U3585) );
  MUX2_X1 U15748 ( .A(n14154), .B(P1_DATAO_REG_24__SCAN_IN), .S(n13817), .Z(
        P1_U3584) );
  MUX2_X1 U15749 ( .A(n13888), .B(P1_DATAO_REG_23__SCAN_IN), .S(n13817), .Z(
        P1_U3583) );
  MUX2_X1 U15750 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14047), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15751 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14194), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15752 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13899), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15753 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14193), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15754 ( .A(n14218), .B(P1_DATAO_REG_18__SCAN_IN), .S(n13817), .Z(
        P1_U3578) );
  MUX2_X1 U15755 ( .A(n14093), .B(P1_DATAO_REG_17__SCAN_IN), .S(n13817), .Z(
        P1_U3577) );
  MUX2_X1 U15756 ( .A(n14547), .B(P1_DATAO_REG_16__SCAN_IN), .S(n13817), .Z(
        P1_U3576) );
  MUX2_X1 U15757 ( .A(n14559), .B(P1_DATAO_REG_15__SCAN_IN), .S(n13817), .Z(
        P1_U3575) );
  MUX2_X1 U15758 ( .A(n14548), .B(P1_DATAO_REG_14__SCAN_IN), .S(n13817), .Z(
        P1_U3574) );
  MUX2_X1 U15759 ( .A(n14558), .B(P1_DATAO_REG_13__SCAN_IN), .S(n13817), .Z(
        P1_U3573) );
  MUX2_X1 U15760 ( .A(n14519), .B(P1_DATAO_REG_12__SCAN_IN), .S(n13817), .Z(
        P1_U3572) );
  MUX2_X1 U15761 ( .A(n14404), .B(P1_DATAO_REG_11__SCAN_IN), .S(n13817), .Z(
        P1_U3571) );
  MUX2_X1 U15762 ( .A(n14520), .B(P1_DATAO_REG_10__SCAN_IN), .S(n13817), .Z(
        P1_U3570) );
  MUX2_X1 U15763 ( .A(n14765), .B(P1_DATAO_REG_9__SCAN_IN), .S(n13817), .Z(
        P1_U3569) );
  MUX2_X1 U15764 ( .A(n13808), .B(P1_DATAO_REG_8__SCAN_IN), .S(n13817), .Z(
        P1_U3568) );
  MUX2_X1 U15765 ( .A(n14744), .B(P1_DATAO_REG_7__SCAN_IN), .S(n13817), .Z(
        P1_U3567) );
  MUX2_X1 U15766 ( .A(n13809), .B(P1_DATAO_REG_6__SCAN_IN), .S(n13817), .Z(
        P1_U3566) );
  MUX2_X1 U15767 ( .A(n13810), .B(P1_DATAO_REG_5__SCAN_IN), .S(n13817), .Z(
        P1_U3565) );
  MUX2_X1 U15768 ( .A(n6446), .B(P1_DATAO_REG_4__SCAN_IN), .S(n13817), .Z(
        P1_U3564) );
  MUX2_X1 U15769 ( .A(n13811), .B(P1_DATAO_REG_3__SCAN_IN), .S(n13817), .Z(
        P1_U3563) );
  MUX2_X1 U15770 ( .A(n13812), .B(P1_DATAO_REG_2__SCAN_IN), .S(n13817), .Z(
        P1_U3562) );
  MUX2_X1 U15771 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13813), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15772 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9693), .S(P1_U4016), .Z(
        P1_U3560) );
  MUX2_X1 U15773 ( .A(n13815), .B(n13814), .S(n14631), .Z(n13820) );
  INV_X1 U15774 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n13818) );
  OAI21_X1 U15775 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n14631), .A(n13816), .ZN(
        n14629) );
  AOI21_X1 U15776 ( .B1(n13818), .B2(n14629), .A(n13817), .ZN(n13819) );
  OAI21_X1 U15777 ( .B1(n13820), .B2(n14262), .A(n13819), .ZN(n14659) );
  AOI22_X1 U15778 ( .A1(n14633), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13830) );
  INV_X1 U15779 ( .A(n13840), .ZN(n13821) );
  AOI211_X1 U15780 ( .C1(n13823), .C2(n13822), .A(n13821), .B(n14666), .ZN(
        n13827) );
  AOI211_X1 U15781 ( .C1(n13825), .C2(n13824), .A(n13837), .B(n14668), .ZN(
        n13826) );
  AOI211_X1 U15782 ( .C1(n14657), .C2(n13828), .A(n13827), .B(n13826), .ZN(
        n13829) );
  NAND3_X1 U15783 ( .A1(n14659), .A2(n13830), .A3(n13829), .ZN(P1_U3245) );
  AND2_X1 U15784 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n14616) );
  NOR2_X1 U15785 ( .A1(n14670), .A2(n13833), .ZN(n13831) );
  AOI211_X1 U15786 ( .C1(n14633), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n14616), .B(
        n13831), .ZN(n13845) );
  INV_X1 U15787 ( .A(n13832), .ZN(n13835) );
  MUX2_X1 U15788 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9309), .S(n13833), .Z(
        n13834) );
  NAND2_X1 U15789 ( .A1(n13835), .A2(n13834), .ZN(n13836) );
  OAI211_X1 U15790 ( .C1(n13837), .C2(n13836), .A(n14652), .B(n14649), .ZN(
        n13844) );
  INV_X1 U15791 ( .A(n14645), .ZN(n13842) );
  NAND3_X1 U15792 ( .A1(n13840), .A2(n13839), .A3(n13838), .ZN(n13841) );
  NAND3_X1 U15793 ( .A1(n14643), .A2(n13842), .A3(n13841), .ZN(n13843) );
  NAND3_X1 U15794 ( .A1(n13845), .A2(n13844), .A3(n13843), .ZN(P1_U3246) );
  NAND2_X1 U15795 ( .A1(n13846), .A2(n13851), .ZN(n13847) );
  NAND2_X1 U15796 ( .A1(n13848), .A2(n13847), .ZN(n13850) );
  XNOR2_X1 U15797 ( .A(n13850), .B(n13849), .ZN(n13860) );
  NAND2_X1 U15798 ( .A1(n13852), .A2(n13851), .ZN(n13853) );
  NAND2_X1 U15799 ( .A1(n13854), .A2(n13853), .ZN(n13855) );
  XOR2_X1 U15800 ( .A(n13855), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13859) );
  INV_X1 U15801 ( .A(n13859), .ZN(n13856) );
  NAND2_X1 U15802 ( .A1(n13856), .A2(n14643), .ZN(n13857) );
  OAI211_X1 U15803 ( .C1(n13860), .C2(n14668), .A(n13857), .B(n14670), .ZN(
        n13858) );
  INV_X1 U15804 ( .A(n13858), .ZN(n13862) );
  AOI22_X1 U15805 ( .A1(n13860), .A2(n14652), .B1(n14643), .B2(n13859), .ZN(
        n13861) );
  MUX2_X1 U15806 ( .A(n13862), .B(n13861), .S(n14022), .Z(n13865) );
  INV_X1 U15807 ( .A(n13863), .ZN(n13864) );
  OAI211_X1 U15808 ( .C1(n7515), .C2(n14674), .A(n13865), .B(n13864), .ZN(
        P1_U3262) );
  INV_X1 U15809 ( .A(n14150), .ZN(n13969) );
  INV_X1 U15810 ( .A(n14175), .ZN(n14020) );
  OR2_X1 U15811 ( .A1(n14187), .A2(n14065), .ZN(n14041) );
  XNOR2_X1 U15812 ( .A(n13873), .B(n13867), .ZN(n13868) );
  NAND2_X1 U15813 ( .A1(n13868), .A2(n14686), .ZN(n14114) );
  INV_X1 U15814 ( .A(P1_B_REG_SCAN_IN), .ZN(n13869) );
  OAI21_X1 U15815 ( .B1(n14631), .B2(n13869), .A(n14745), .ZN(n13913) );
  OR2_X1 U15816 ( .A1(n13870), .A2(n13913), .ZN(n14116) );
  NOR2_X1 U15817 ( .A1(n14704), .A2(n14116), .ZN(n13876) );
  NOR2_X1 U15818 ( .A1(n14115), .A2(n14096), .ZN(n13871) );
  AOI211_X1 U15819 ( .C1(n14704), .C2(P1_REG2_REG_31__SCAN_IN), .A(n13876), 
        .B(n13871), .ZN(n13872) );
  OAI21_X1 U15820 ( .B1(n14114), .B2(n14066), .A(n13872), .ZN(P1_U3263) );
  OAI211_X1 U15821 ( .C1(n14118), .C2(n6958), .A(n13874), .B(n14686), .ZN(
        n14117) );
  NOR2_X1 U15822 ( .A1(n14118), .A2(n14096), .ZN(n13875) );
  AOI211_X1 U15823 ( .C1(n14704), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13876), 
        .B(n13875), .ZN(n13877) );
  OAI21_X1 U15824 ( .B1(n14117), .B2(n14066), .A(n13877), .ZN(P1_U3264) );
  OR2_X1 U15825 ( .A1(n14221), .A2(n14210), .ZN(n13879) );
  NAND2_X1 U15826 ( .A1(n13880), .A2(n13879), .ZN(n14085) );
  OR2_X1 U15827 ( .A1(n14197), .A2(n14203), .ZN(n13883) );
  NAND2_X1 U15828 ( .A1(n14175), .A2(n13888), .ZN(n13889) );
  INV_X1 U15829 ( .A(n13979), .ZN(n13992) );
  NAND2_X1 U15830 ( .A1(n14150), .A2(n14155), .ZN(n13890) );
  INV_X1 U15831 ( .A(n14142), .ZN(n13951) );
  NAND2_X1 U15832 ( .A1(n13951), .A2(n14147), .ZN(n13892) );
  NAND2_X1 U15833 ( .A1(n14221), .A2(n14093), .ZN(n13895) );
  NAND2_X1 U15834 ( .A1(n14100), .A2(n14099), .ZN(n14098) );
  AND2_X2 U15835 ( .A1(n14098), .A2(n13897), .ZN(n14080) );
  NAND2_X1 U15836 ( .A1(n14205), .A2(n14211), .ZN(n13898) );
  NAND2_X1 U15837 ( .A1(n14197), .A2(n13899), .ZN(n13900) );
  NAND2_X1 U15838 ( .A1(n14049), .A2(n14194), .ZN(n13901) );
  NAND2_X1 U15839 ( .A1(n14180), .A2(n14184), .ZN(n13903) );
  AND2_X1 U15840 ( .A1(n14175), .A2(n14167), .ZN(n13904) );
  NAND2_X1 U15841 ( .A1(n13983), .A2(n14166), .ZN(n13905) );
  INV_X1 U15842 ( .A(n13971), .ZN(n13958) );
  NAND2_X1 U15843 ( .A1(n13959), .A2(n13958), .ZN(n13907) );
  NAND2_X1 U15844 ( .A1(n14150), .A2(n14139), .ZN(n13906) );
  NAND2_X2 U15845 ( .A1(n13907), .A2(n13906), .ZN(n13955) );
  AOI21_X1 U15846 ( .B1(n13931), .B2(n13909), .A(n14572), .ZN(n13911) );
  NAND2_X1 U15847 ( .A1(n13911), .A2(n13910), .ZN(n14122) );
  NOR2_X1 U15848 ( .A1(n14122), .A2(n14066), .ZN(n13923) );
  INV_X1 U15849 ( .A(n13912), .ZN(n13914) );
  NOR2_X1 U15850 ( .A1(n13914), .A2(n13913), .ZN(n14119) );
  NAND2_X1 U15851 ( .A1(n14119), .A2(n13915), .ZN(n13918) );
  OAI22_X1 U15852 ( .A1(n13918), .A2(n13917), .B1(n13916), .B2(n14706), .ZN(
        n13920) );
  NOR2_X1 U15853 ( .A1(n14064), .A2(n14138), .ZN(n13919) );
  AOI211_X1 U15854 ( .C1(n14704), .C2(P1_REG2_REG_29__SCAN_IN), .A(n13920), 
        .B(n13919), .ZN(n13921) );
  OAI21_X1 U15855 ( .B1(n14123), .B2(n14096), .A(n13921), .ZN(n13922) );
  AOI211_X1 U15856 ( .C1(n14125), .C2(n14434), .A(n13923), .B(n13922), .ZN(
        n13924) );
  OAI21_X1 U15857 ( .B1(n14128), .B2(n14700), .A(n13924), .ZN(P1_U3356) );
  XNOR2_X1 U15858 ( .A(n13926), .B(n13925), .ZN(n13927) );
  NAND2_X1 U15859 ( .A1(n13927), .A2(n14763), .ZN(n13930) );
  AOI22_X1 U15860 ( .A1(n14745), .A2(n13928), .B1(n13967), .B2(n14766), .ZN(
        n13929) );
  NAND2_X1 U15861 ( .A1(n13930), .A2(n13929), .ZN(n14129) );
  OAI211_X1 U15862 ( .C1(n14132), .C2(n13947), .A(n14686), .B(n13931), .ZN(
        n14134) );
  NAND2_X1 U15863 ( .A1(n13933), .A2(n13932), .ZN(n14131) );
  NAND3_X1 U15864 ( .A1(n14131), .A2(n14544), .A3(n14130), .ZN(n13939) );
  INV_X1 U15865 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n13935) );
  OAI22_X1 U15866 ( .A1(n14437), .A2(n13935), .B1(n13934), .B2(n14706), .ZN(
        n13936) );
  AOI21_X1 U15867 ( .B1(n13937), .B2(n14683), .A(n13936), .ZN(n13938) );
  OAI211_X1 U15868 ( .C1(n14066), .C2(n14134), .A(n13939), .B(n13938), .ZN(
        n13940) );
  AOI21_X1 U15869 ( .B1(n14129), .B2(n14437), .A(n13940), .ZN(n13941) );
  INV_X1 U15870 ( .A(n13941), .ZN(P1_U3265) );
  INV_X1 U15871 ( .A(n13942), .ZN(n13943) );
  NAND2_X1 U15872 ( .A1(n14142), .A2(n13961), .ZN(n13945) );
  NAND2_X1 U15873 ( .A1(n13945), .A2(n14686), .ZN(n13946) );
  NOR2_X1 U15874 ( .A1(n13947), .A2(n13946), .ZN(n14140) );
  AOI22_X1 U15875 ( .A1(n14704), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13948), 
        .B2(n14682), .ZN(n13950) );
  NAND2_X1 U15876 ( .A1(n14061), .A2(n14120), .ZN(n13949) );
  OAI211_X1 U15877 ( .C1(n14139), .C2(n14064), .A(n13950), .B(n13949), .ZN(
        n13953) );
  NOR2_X1 U15878 ( .A1(n13951), .A2(n14096), .ZN(n13952) );
  AOI211_X1 U15879 ( .C1(n14140), .C2(n14690), .A(n13953), .B(n13952), .ZN(
        n13957) );
  XNOR2_X1 U15880 ( .A(n13955), .B(n13954), .ZN(n14143) );
  NAND2_X1 U15881 ( .A1(n14143), .A2(n14434), .ZN(n13956) );
  OAI211_X1 U15882 ( .C1(n14146), .C2(n14700), .A(n13957), .B(n13956), .ZN(
        P1_U3266) );
  XNOR2_X1 U15883 ( .A(n13959), .B(n13958), .ZN(n13960) );
  NAND2_X1 U15884 ( .A1(n13960), .A2(n14763), .ZN(n14151) );
  INV_X1 U15885 ( .A(n13961), .ZN(n13962) );
  AOI211_X1 U15886 ( .C1(n14150), .C2(n6942), .A(n14572), .B(n13962), .ZN(
        n14148) );
  INV_X1 U15887 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n13964) );
  OAI22_X1 U15888 ( .A1(n14437), .A2(n13964), .B1(n13963), .B2(n14706), .ZN(
        n13966) );
  NOR2_X1 U15889 ( .A1(n14064), .A2(n14166), .ZN(n13965) );
  AOI211_X1 U15890 ( .C1(n14061), .C2(n13967), .A(n13966), .B(n13965), .ZN(
        n13968) );
  OAI21_X1 U15891 ( .B1(n13969), .B2(n14096), .A(n13968), .ZN(n13974) );
  OAI21_X1 U15892 ( .B1(n13972), .B2(n13971), .A(n13970), .ZN(n14153) );
  NOR2_X1 U15893 ( .A1(n14153), .A2(n14700), .ZN(n13973) );
  AOI211_X1 U15894 ( .C1(n14148), .C2(n14690), .A(n13974), .B(n13973), .ZN(
        n13975) );
  OAI21_X1 U15895 ( .B1(n14704), .B2(n14151), .A(n13975), .ZN(P1_U3267) );
  INV_X1 U15896 ( .A(n13976), .ZN(n13977) );
  AOI21_X1 U15897 ( .B1(n13979), .B2(n13978), .A(n13977), .ZN(n14163) );
  NAND2_X1 U15898 ( .A1(n13999), .A2(n13983), .ZN(n13980) );
  NAND2_X1 U15899 ( .A1(n13980), .A2(n14686), .ZN(n13981) );
  OR2_X1 U15900 ( .A1(n13982), .A2(n13981), .ZN(n14157) );
  INV_X1 U15901 ( .A(n14157), .ZN(n13991) );
  NAND2_X1 U15902 ( .A1(n14704), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n13986) );
  NAND2_X1 U15903 ( .A1(n13984), .A2(n14682), .ZN(n13985) );
  OAI211_X1 U15904 ( .C1(n14064), .C2(n13987), .A(n13986), .B(n13985), .ZN(
        n13988) );
  AOI21_X1 U15905 ( .B1(n14061), .B2(n14155), .A(n13988), .ZN(n13989) );
  OAI21_X1 U15906 ( .B1(n6940), .B2(n14096), .A(n13989), .ZN(n13990) );
  AOI21_X1 U15907 ( .B1(n13991), .B2(n14690), .A(n13990), .ZN(n13995) );
  NAND2_X1 U15908 ( .A1(n13993), .A2(n13992), .ZN(n14159) );
  NAND3_X1 U15909 ( .A1(n14160), .A2(n14159), .A3(n14544), .ZN(n13994) );
  OAI211_X1 U15910 ( .C1(n14163), .C2(n14701), .A(n13995), .B(n13994), .ZN(
        P1_U3268) );
  XOR2_X1 U15911 ( .A(n13997), .B(n13996), .Z(n14173) );
  OR2_X1 U15912 ( .A1(n13998), .A2(n13997), .ZN(n14165) );
  NAND3_X1 U15913 ( .A1(n14165), .A2(n14164), .A3(n14434), .ZN(n14008) );
  AOI21_X1 U15914 ( .B1(n14015), .B2(n14170), .A(n14572), .ZN(n14000) );
  AND2_X1 U15915 ( .A1(n14000), .A2(n13999), .ZN(n14168) );
  AOI22_X1 U15916 ( .A1(n14704), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14001), 
        .B2(n14682), .ZN(n14002) );
  OAI21_X1 U15917 ( .B1(n14167), .B2(n14064), .A(n14002), .ZN(n14003) );
  AOI21_X1 U15918 ( .B1(n14061), .B2(n14004), .A(n14003), .ZN(n14005) );
  OAI21_X1 U15919 ( .B1(n6941), .B2(n14096), .A(n14005), .ZN(n14006) );
  AOI21_X1 U15920 ( .B1(n14168), .B2(n14690), .A(n14006), .ZN(n14007) );
  OAI211_X1 U15921 ( .C1(n14173), .C2(n14700), .A(n14008), .B(n14007), .ZN(
        P1_U3269) );
  INV_X1 U15922 ( .A(n14009), .ZN(n14024) );
  OAI21_X1 U15923 ( .B1(n14011), .B2(n7351), .A(n6628), .ZN(n14178) );
  XNOR2_X1 U15924 ( .A(n6608), .B(n14012), .ZN(n14014) );
  AOI222_X1 U15925 ( .A1(n14763), .A2(n14014), .B1(n14047), .B2(n14766), .C1(
        n14154), .C2(n14745), .ZN(n14177) );
  INV_X1 U15926 ( .A(n14029), .ZN(n14017) );
  INV_X1 U15927 ( .A(n14015), .ZN(n14016) );
  AOI211_X1 U15928 ( .C1(n14175), .C2(n14017), .A(n14572), .B(n14016), .ZN(
        n14174) );
  OAI22_X1 U15929 ( .A1(n14020), .A2(n14019), .B1(n14018), .B2(n14706), .ZN(
        n14021) );
  AOI21_X1 U15930 ( .B1(n14174), .B2(n14022), .A(n14021), .ZN(n14023) );
  OAI211_X1 U15931 ( .C1(n14024), .C2(n14178), .A(n14177), .B(n14023), .ZN(
        n14025) );
  MUX2_X1 U15932 ( .A(P1_REG2_REG_23__SCAN_IN), .B(n14025), .S(n14437), .Z(
        P1_U3270) );
  XNOR2_X1 U15933 ( .A(n14026), .B(n6630), .ZN(n14183) );
  NAND2_X1 U15934 ( .A1(n14180), .A2(n14041), .ZN(n14027) );
  NAND2_X1 U15935 ( .A1(n14027), .A2(n14686), .ZN(n14028) );
  NOR2_X1 U15936 ( .A1(n14029), .A2(n14028), .ZN(n14179) );
  NAND2_X1 U15937 ( .A1(n14180), .A2(n14683), .ZN(n14031) );
  NAND2_X1 U15938 ( .A1(n14704), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n14030) );
  OAI211_X1 U15939 ( .C1(n14706), .C2(n14032), .A(n14031), .B(n14030), .ZN(
        n14037) );
  OAI21_X1 U15940 ( .B1(n6439), .B2(n6630), .A(n14033), .ZN(n14035) );
  AOI21_X1 U15941 ( .B1(n14035), .B2(n14763), .A(n14034), .ZN(n14182) );
  NOR2_X1 U15942 ( .A1(n14182), .A2(n14704), .ZN(n14036) );
  AOI211_X1 U15943 ( .C1(n14179), .C2(n14690), .A(n14037), .B(n14036), .ZN(
        n14038) );
  OAI21_X1 U15944 ( .B1(n14183), .B2(n14700), .A(n14038), .ZN(P1_U3271) );
  OAI211_X1 U15945 ( .C1(n14040), .C2(n14053), .A(n14763), .B(n14039), .ZN(
        n14188) );
  INV_X1 U15946 ( .A(n14041), .ZN(n14042) );
  AOI211_X1 U15947 ( .C1(n14187), .C2(n14065), .A(n14572), .B(n14042), .ZN(
        n14185) );
  INV_X1 U15948 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14044) );
  OAI22_X1 U15949 ( .A1(n14437), .A2(n14044), .B1(n14043), .B2(n14706), .ZN(
        n14046) );
  NOR2_X1 U15950 ( .A1(n14064), .A2(n14203), .ZN(n14045) );
  AOI211_X1 U15951 ( .C1(n14061), .C2(n14047), .A(n14046), .B(n14045), .ZN(
        n14048) );
  OAI21_X1 U15952 ( .B1(n14049), .B2(n14096), .A(n14048), .ZN(n14055) );
  INV_X1 U15953 ( .A(n14051), .ZN(n14052) );
  AOI21_X1 U15954 ( .B1(n14053), .B2(n14050), .A(n14052), .ZN(n14190) );
  NOR2_X1 U15955 ( .A1(n14190), .A2(n14700), .ZN(n14054) );
  AOI211_X1 U15956 ( .C1(n14185), .C2(n14690), .A(n14055), .B(n14054), .ZN(
        n14056) );
  OAI21_X1 U15957 ( .B1(n14704), .B2(n14188), .A(n14056), .ZN(P1_U3272) );
  OAI21_X1 U15958 ( .B1(n7437), .B2(n14058), .A(n14057), .ZN(n14201) );
  NAND2_X1 U15959 ( .A1(n14059), .A2(n14058), .ZN(n14191) );
  NAND3_X1 U15960 ( .A1(n14192), .A2(n14191), .A3(n14434), .ZN(n14071) );
  AOI22_X1 U15961 ( .A1(n14704), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14060), 
        .B2(n14682), .ZN(n14063) );
  NAND2_X1 U15962 ( .A1(n14061), .A2(n14194), .ZN(n14062) );
  OAI211_X1 U15963 ( .C1(n14211), .C2(n14064), .A(n14063), .B(n14062), .ZN(
        n14068) );
  OAI211_X1 U15964 ( .C1(n14197), .C2(n6558), .A(n14686), .B(n14065), .ZN(
        n14196) );
  NOR2_X1 U15965 ( .A1(n14196), .A2(n14066), .ZN(n14067) );
  AOI211_X1 U15966 ( .C1(n14683), .C2(n14069), .A(n14068), .B(n14067), .ZN(
        n14070) );
  OAI211_X1 U15967 ( .C1(n14201), .C2(n14700), .A(n14071), .B(n14070), .ZN(
        P1_U3273) );
  XOR2_X1 U15968 ( .A(n14072), .B(n14078), .Z(n14208) );
  AND2_X1 U15969 ( .A1(n14205), .A2(n14087), .ZN(n14073) );
  AOI22_X1 U15970 ( .A1(n14704), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14074), 
        .B2(n14682), .ZN(n14075) );
  OAI21_X1 U15971 ( .B1(n14091), .B2(n14203), .A(n14075), .ZN(n14076) );
  AOI21_X1 U15972 ( .B1(n14094), .B2(n14218), .A(n14076), .ZN(n14077) );
  OAI21_X1 U15973 ( .B1(n6952), .B2(n14096), .A(n14077), .ZN(n14083) );
  OAI21_X1 U15974 ( .B1(n14080), .B2(n6771), .A(n14079), .ZN(n14081) );
  NAND2_X1 U15975 ( .A1(n14081), .A2(n14763), .ZN(n14207) );
  NOR2_X1 U15976 ( .A1(n14207), .A2(n14704), .ZN(n14082) );
  AOI211_X1 U15977 ( .C1(n6469), .C2(n14690), .A(n14083), .B(n14082), .ZN(
        n14084) );
  OAI21_X1 U15978 ( .B1(n14700), .B2(n14208), .A(n14084), .ZN(P1_U3274) );
  XOR2_X1 U15979 ( .A(n14085), .B(n14099), .Z(n14217) );
  OR2_X1 U15980 ( .A1(n14097), .A2(n14086), .ZN(n14088) );
  AND3_X1 U15981 ( .A1(n14686), .A2(n14088), .A3(n14087), .ZN(n14212) );
  AOI22_X1 U15982 ( .A1(n14704), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14089), 
        .B2(n14682), .ZN(n14090) );
  OAI21_X1 U15983 ( .B1(n14091), .B2(n14211), .A(n14090), .ZN(n14092) );
  AOI21_X1 U15984 ( .B1(n14094), .B2(n14093), .A(n14092), .ZN(n14095) );
  OAI21_X1 U15985 ( .B1(n14097), .B2(n14096), .A(n14095), .ZN(n14102) );
  OAI211_X1 U15986 ( .C1(n14100), .C2(n14099), .A(n14098), .B(n14763), .ZN(
        n14215) );
  NOR2_X1 U15987 ( .A1(n14215), .A2(n14704), .ZN(n14101) );
  AOI211_X1 U15988 ( .C1(n14212), .C2(n14690), .A(n14102), .B(n14101), .ZN(
        n14103) );
  OAI21_X1 U15989 ( .B1(n14700), .B2(n14217), .A(n14103), .ZN(P1_U3275) );
  MUX2_X1 U15990 ( .A(n14104), .B(P1_REG2_REG_1__SCAN_IN), .S(n14704), .Z(
        n14105) );
  INV_X1 U15991 ( .A(n14105), .ZN(n14113) );
  INV_X1 U15992 ( .A(n14106), .ZN(n14107) );
  AND2_X1 U15993 ( .A1(n14437), .A2(n14107), .ZN(n14691) );
  AOI22_X1 U15994 ( .A1(n14691), .A2(n14108), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n14682), .ZN(n14112) );
  AOI22_X1 U15995 ( .A1(n14110), .A2(n14690), .B1(n14683), .B2(n14109), .ZN(
        n14111) );
  NAND3_X1 U15996 ( .A1(n14113), .A2(n14112), .A3(n14111), .ZN(P1_U3292) );
  OAI211_X1 U15997 ( .C1(n14115), .C2(n14748), .A(n14114), .B(n14116), .ZN(
        n14233) );
  MUX2_X1 U15998 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14233), .S(n14790), .Z(
        P1_U3559) );
  OAI211_X1 U15999 ( .C1(n14118), .C2(n14748), .A(n14117), .B(n14116), .ZN(
        n14234) );
  MUX2_X1 U16000 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14234), .S(n14790), .Z(
        P1_U3558) );
  AOI21_X1 U16001 ( .B1(n14766), .B2(n14120), .A(n14119), .ZN(n14121) );
  OAI211_X1 U16002 ( .C1(n14123), .C2(n14748), .A(n14122), .B(n14121), .ZN(
        n14124) );
  NAND2_X1 U16003 ( .A1(n14125), .A2(n14763), .ZN(n14126) );
  OAI211_X1 U16004 ( .C1(n14128), .C2(n14755), .A(n14127), .B(n14126), .ZN(
        n14235) );
  MUX2_X1 U16005 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14235), .S(n14790), .Z(
        P1_U3557) );
  INV_X1 U16006 ( .A(n14129), .ZN(n14137) );
  NAND3_X1 U16007 ( .A1(n14131), .A2(n14774), .A3(n14130), .ZN(n14136) );
  MUX2_X1 U16008 ( .A(n14236), .B(P1_REG1_REG_28__SCAN_IN), .S(n14787), .Z(
        P1_U3556) );
  OAI22_X1 U16009 ( .A1(n14139), .A2(n14209), .B1(n14138), .B2(n14420), .ZN(
        n14141) );
  AOI211_X1 U16010 ( .C1(n14142), .C2(n14767), .A(n14141), .B(n14140), .ZN(
        n14145) );
  NAND2_X1 U16011 ( .A1(n14143), .A2(n14763), .ZN(n14144) );
  MUX2_X1 U16012 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14237), .S(n14790), .Z(
        P1_U3555) );
  OAI22_X1 U16013 ( .A1(n14147), .A2(n14420), .B1(n14166), .B2(n14209), .ZN(
        n14149) );
  AOI211_X1 U16014 ( .C1(n14150), .C2(n14767), .A(n14149), .B(n14148), .ZN(
        n14152) );
  OAI211_X1 U16015 ( .C1(n14755), .C2(n14153), .A(n14152), .B(n14151), .ZN(
        n14238) );
  MUX2_X1 U16016 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14238), .S(n14790), .Z(
        P1_U3554) );
  AOI22_X1 U16017 ( .A1(n14745), .A2(n14155), .B1(n14154), .B2(n14766), .ZN(
        n14156) );
  OAI211_X1 U16018 ( .C1(n6940), .C2(n14748), .A(n14157), .B(n14156), .ZN(
        n14158) );
  INV_X1 U16019 ( .A(n14158), .ZN(n14162) );
  NAND3_X1 U16020 ( .A1(n14160), .A2(n14159), .A3(n14774), .ZN(n14161) );
  OAI211_X1 U16021 ( .C1(n14163), .C2(n14574), .A(n14162), .B(n14161), .ZN(
        n14239) );
  MUX2_X1 U16022 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14239), .S(n14790), .Z(
        P1_U3553) );
  NAND3_X1 U16023 ( .A1(n14165), .A2(n14763), .A3(n14164), .ZN(n14172) );
  OAI22_X1 U16024 ( .A1(n14167), .A2(n14209), .B1(n14166), .B2(n14420), .ZN(
        n14169) );
  AOI211_X1 U16025 ( .C1(n14170), .C2(n14767), .A(n14169), .B(n14168), .ZN(
        n14171) );
  OAI211_X1 U16026 ( .C1(n14755), .C2(n14173), .A(n14172), .B(n14171), .ZN(
        n14240) );
  MUX2_X1 U16027 ( .A(n14240), .B(P1_REG1_REG_24__SCAN_IN), .S(n14787), .Z(
        P1_U3552) );
  AOI21_X1 U16028 ( .B1(n14175), .B2(n14767), .A(n14174), .ZN(n14176) );
  OAI211_X1 U16029 ( .C1(n14755), .C2(n14178), .A(n14177), .B(n14176), .ZN(
        n14241) );
  MUX2_X1 U16030 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14241), .S(n14790), .Z(
        P1_U3551) );
  AOI21_X1 U16031 ( .B1(n14180), .B2(n14767), .A(n14179), .ZN(n14181) );
  OAI211_X1 U16032 ( .C1(n14755), .C2(n14183), .A(n14182), .B(n14181), .ZN(
        n14242) );
  MUX2_X1 U16033 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14242), .S(n14790), .Z(
        P1_U3550) );
  OAI22_X1 U16034 ( .A1(n14184), .A2(n14420), .B1(n14203), .B2(n14209), .ZN(
        n14186) );
  AOI211_X1 U16035 ( .C1(n14187), .C2(n14767), .A(n14186), .B(n14185), .ZN(
        n14189) );
  OAI211_X1 U16036 ( .C1(n14190), .C2(n14755), .A(n14189), .B(n14188), .ZN(
        n14243) );
  MUX2_X1 U16037 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14243), .S(n14790), .Z(
        P1_U3549) );
  NAND3_X1 U16038 ( .A1(n14192), .A2(n14763), .A3(n14191), .ZN(n14200) );
  AOI22_X1 U16039 ( .A1(n14194), .A2(n14745), .B1(n14766), .B2(n14193), .ZN(
        n14195) );
  OAI211_X1 U16040 ( .C1(n14197), .C2(n14748), .A(n14196), .B(n14195), .ZN(
        n14198) );
  INV_X1 U16041 ( .A(n14198), .ZN(n14199) );
  OAI211_X1 U16042 ( .C1(n14755), .C2(n14201), .A(n14200), .B(n14199), .ZN(
        n14244) );
  MUX2_X1 U16043 ( .A(n14244), .B(P1_REG1_REG_20__SCAN_IN), .S(n14787), .Z(
        P1_U3548) );
  OAI22_X1 U16044 ( .A1(n14203), .A2(n14420), .B1(n14202), .B2(n14209), .ZN(
        n14204) );
  AOI211_X1 U16045 ( .C1(n14205), .C2(n14767), .A(n14204), .B(n6469), .ZN(
        n14206) );
  OAI211_X1 U16046 ( .C1(n14755), .C2(n14208), .A(n14207), .B(n14206), .ZN(
        n14245) );
  MUX2_X1 U16047 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14245), .S(n14790), .Z(
        P1_U3547) );
  OAI22_X1 U16048 ( .A1(n14211), .A2(n14420), .B1(n14210), .B2(n14209), .ZN(
        n14213) );
  AOI211_X1 U16049 ( .C1(n14214), .C2(n14767), .A(n14213), .B(n14212), .ZN(
        n14216) );
  OAI211_X1 U16050 ( .C1(n14217), .C2(n14755), .A(n14216), .B(n14215), .ZN(
        n14246) );
  MUX2_X1 U16051 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14246), .S(n14790), .Z(
        P1_U3546) );
  AOI22_X1 U16052 ( .A1(n14218), .A2(n14745), .B1(n14766), .B2(n14547), .ZN(
        n14219) );
  OAI211_X1 U16053 ( .C1(n14221), .C2(n14748), .A(n14220), .B(n14219), .ZN(
        n14222) );
  AOI21_X1 U16054 ( .B1(n14223), .B2(n14763), .A(n14222), .ZN(n14224) );
  OAI21_X1 U16055 ( .B1(n14755), .B2(n14225), .A(n14224), .ZN(n14247) );
  MUX2_X1 U16056 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14247), .S(n14790), .Z(
        P1_U3545) );
  AOI21_X1 U16057 ( .B1(n14227), .B2(n14767), .A(n14226), .ZN(n14228) );
  OAI211_X1 U16058 ( .C1(n14755), .C2(n14230), .A(n14229), .B(n14228), .ZN(
        n14248) );
  MUX2_X1 U16059 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14248), .S(n14790), .Z(
        P1_U3544) );
  MUX2_X1 U16060 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n14231), .S(n14790), .Z(
        P1_U3533) );
  MUX2_X1 U16061 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n14232), .S(n14790), .Z(
        P1_U3528) );
  MUX2_X1 U16062 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14233), .S(n6444), .Z(
        P1_U3527) );
  MUX2_X1 U16063 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14234), .S(n6444), .Z(
        P1_U3526) );
  MUX2_X1 U16064 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14235), .S(n6444), .Z(
        P1_U3525) );
  MUX2_X1 U16065 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14236), .S(n6444), .Z(
        P1_U3524) );
  MUX2_X1 U16066 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14237), .S(n6444), .Z(
        P1_U3523) );
  MUX2_X1 U16067 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14238), .S(n6444), .Z(
        P1_U3522) );
  MUX2_X1 U16068 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14239), .S(n6444), .Z(
        P1_U3521) );
  MUX2_X1 U16069 ( .A(n14240), .B(P1_REG0_REG_24__SCAN_IN), .S(n14775), .Z(
        P1_U3520) );
  MUX2_X1 U16070 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14241), .S(n6444), .Z(
        P1_U3519) );
  MUX2_X1 U16071 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14242), .S(n6444), .Z(
        P1_U3518) );
  MUX2_X1 U16072 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14243), .S(n6444), .Z(
        P1_U3517) );
  MUX2_X1 U16073 ( .A(n14244), .B(P1_REG0_REG_20__SCAN_IN), .S(n14775), .Z(
        P1_U3516) );
  MUX2_X1 U16074 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14245), .S(n6444), .Z(
        P1_U3515) );
  MUX2_X1 U16075 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14246), .S(n6444), .Z(
        P1_U3513) );
  MUX2_X1 U16076 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14247), .S(n6444), .Z(
        P1_U3510) );
  MUX2_X1 U16077 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14248), .S(n6444), .Z(
        P1_U3507) );
  INV_X1 U16078 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14250) );
  NAND3_X1 U16079 ( .A1(n14250), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n14252) );
  OAI22_X1 U16080 ( .A1(n14249), .A2(n14252), .B1(n14251), .B2(n14276), .ZN(
        n14253) );
  AOI21_X1 U16081 ( .B1(n14254), .B2(n14272), .A(n14253), .ZN(n14255) );
  INV_X1 U16082 ( .A(n14255), .ZN(P1_U3324) );
  OAI222_X1 U16083 ( .A1(n14276), .A2(n15172), .B1(n14270), .B2(n14257), .C1(
        n14256), .C2(P1_U3086), .ZN(P1_U3325) );
  OAI222_X1 U16084 ( .A1(n14276), .A2(n14260), .B1(n14270), .B2(n14259), .C1(
        n14258), .C2(P1_U3086), .ZN(P1_U3326) );
  INV_X1 U16085 ( .A(n14261), .ZN(n14263) );
  OAI222_X1 U16086 ( .A1(n14276), .A2(n14264), .B1(n14270), .B2(n14263), .C1(
        P1_U3086), .C2(n14262), .ZN(P1_U3327) );
  OAI222_X1 U16087 ( .A1(n14267), .A2(P1_U3086), .B1(n14270), .B2(n14266), 
        .C1(n14265), .C2(n14276), .ZN(P1_U3329) );
  INV_X1 U16088 ( .A(n9272), .ZN(n14268) );
  OAI222_X1 U16089 ( .A1(n14276), .A2(n14271), .B1(n14270), .B2(n14269), .C1(
        n14268), .C2(P1_U3086), .ZN(P1_U3330) );
  NAND2_X1 U16090 ( .A1(n14273), .A2(n14272), .ZN(n14275) );
  OAI211_X1 U16091 ( .C1(n14277), .C2(n14276), .A(n14275), .B(n14274), .ZN(
        P1_U3332) );
  MUX2_X1 U16092 ( .A(n14279), .B(n14278), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16093 ( .A(n14280), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16094 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14316) );
  INV_X1 U16095 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15108) );
  INV_X1 U16096 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14977) );
  INV_X1 U16097 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14308) );
  INV_X1 U16098 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14306) );
  XOR2_X1 U16099 ( .A(n15218), .B(n14306), .Z(n14325) );
  INV_X1 U16100 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14302) );
  XNOR2_X1 U16101 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n14360) );
  INV_X1 U16102 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14300) );
  NOR2_X1 U16103 ( .A1(n14334), .A2(n14333), .ZN(n14282) );
  NOR2_X1 U16104 ( .A1(n14285), .A2(n14286), .ZN(n14288) );
  NOR2_X1 U16105 ( .A1(n14289), .A2(n14935), .ZN(n14291) );
  NOR2_X2 U16106 ( .A1(n14291), .A2(n14290), .ZN(n14349) );
  INV_X1 U16107 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14292) );
  NOR2_X1 U16108 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14292), .ZN(n14294) );
  INV_X1 U16109 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14293) );
  NOR2_X1 U16110 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14295), .ZN(n14298) );
  XNOR2_X1 U16111 ( .A(n14300), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n14329) );
  NAND2_X1 U16112 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14303), .ZN(n14327) );
  NAND2_X1 U16113 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n14327), .ZN(n14304) );
  NAND2_X1 U16114 ( .A1(n14326), .A2(n14304), .ZN(n14324) );
  XNOR2_X1 U16115 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n14368) );
  NAND2_X1 U16116 ( .A1(n14369), .A2(n14368), .ZN(n14307) );
  OAI21_X1 U16117 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14308), .A(n14307), 
        .ZN(n14309) );
  INV_X1 U16118 ( .A(n14309), .ZN(n14323) );
  AND2_X1 U16119 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14977), .ZN(n14310) );
  INV_X1 U16120 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14311) );
  NOR2_X1 U16121 ( .A1(n14311), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n14312) );
  OAI22_X1 U16122 ( .A1(n15108), .A2(P3_ADDR_REG_14__SCAN_IN), .B1(n14374), 
        .B2(n14312), .ZN(n14379) );
  INV_X1 U16123 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14675) );
  NOR2_X1 U16124 ( .A1(n14675), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n14313) );
  INV_X1 U16125 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14456) );
  OAI22_X1 U16126 ( .A1(n14379), .A2(n14313), .B1(n14456), .B2(
        P1_ADDR_REG_15__SCAN_IN), .ZN(n14381) );
  INV_X1 U16127 ( .A(n14381), .ZN(n14315) );
  OR2_X1 U16128 ( .A1(n14316), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n14314) );
  AOI22_X1 U16129 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14316), .B1(n14315), 
        .B2(n14314), .ZN(n14317) );
  INV_X1 U16130 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14318) );
  NAND2_X1 U16131 ( .A1(n14317), .A2(n14318), .ZN(n14320) );
  XOR2_X1 U16132 ( .A(n14318), .B(n14317), .Z(n14384) );
  NAND2_X1 U16133 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14384), .ZN(n14319) );
  NAND2_X1 U16134 ( .A1(n14320), .A2(n14319), .ZN(n14446) );
  NOR2_X1 U16135 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n14449), .ZN(n14321) );
  AOI21_X1 U16136 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n14449), .A(n14321), 
        .ZN(n14447) );
  XNOR2_X1 U16137 ( .A(n14446), .B(n14447), .ZN(n14445) );
  INV_X1 U16138 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14442) );
  INV_X1 U16139 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14613) );
  INV_X1 U16140 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14608) );
  XOR2_X1 U16141 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n14322) );
  XNOR2_X1 U16142 ( .A(n14323), .B(n14322), .ZN(n14599) );
  XOR2_X1 U16143 ( .A(n14325), .B(n14324), .Z(n14595) );
  NAND2_X1 U16144 ( .A1(n14327), .A2(n14326), .ZN(n14328) );
  XOR2_X1 U16145 ( .A(n14330), .B(n14329), .Z(n14358) );
  XNOR2_X1 U16146 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n14331), .ZN(n14332) );
  NAND2_X1 U16147 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14332), .ZN(n14345) );
  INV_X1 U16148 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14392) );
  XNOR2_X1 U16149 ( .A(n14334), .B(n14333), .ZN(n14390) );
  NAND2_X1 U16150 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14338), .ZN(n14340) );
  AOI21_X1 U16151 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14337), .A(n14336), .ZN(
        n15242) );
  NOR2_X1 U16152 ( .A1(n15242), .A2(n9531), .ZN(n15250) );
  XOR2_X1 U16153 ( .A(n14338), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15249) );
  NAND2_X1 U16154 ( .A1(n15250), .A2(n15249), .ZN(n14339) );
  NAND2_X1 U16155 ( .A1(n14390), .A2(n14391), .ZN(n14341) );
  NOR2_X1 U16156 ( .A1(n14390), .A2(n14391), .ZN(n14389) );
  XNOR2_X1 U16157 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14342), .ZN(n15247) );
  NOR2_X1 U16158 ( .A1(n15246), .A2(n15247), .ZN(n14344) );
  INV_X1 U16159 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n14343) );
  NAND2_X1 U16160 ( .A1(n15246), .A2(n15247), .ZN(n15245) );
  OAI21_X1 U16161 ( .B1(n14344), .B2(n14343), .A(n15245), .ZN(n15239) );
  XNOR2_X1 U16162 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n14350) );
  XOR2_X1 U16163 ( .A(n14350), .B(n14349), .Z(n14394) );
  NAND2_X1 U16164 ( .A1(n14351), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14352) );
  NAND2_X1 U16165 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14353), .ZN(n14356) );
  XNOR2_X1 U16166 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14354), .ZN(n15243) );
  NAND2_X1 U16167 ( .A1(n15244), .A2(n15243), .ZN(n14355) );
  XNOR2_X1 U16168 ( .A(n14360), .B(n14359), .ZN(n14362) );
  NAND2_X1 U16169 ( .A1(n14361), .A2(n14362), .ZN(n14363) );
  NAND2_X1 U16170 ( .A1(n14403), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n14367) );
  NAND2_X1 U16171 ( .A1(n14365), .A2(n14364), .ZN(n14366) );
  INV_X1 U16172 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n15130) );
  NAND2_X1 U16173 ( .A1(n14595), .A2(n14596), .ZN(n14594) );
  XNOR2_X1 U16174 ( .A(n14369), .B(n14368), .ZN(n14370) );
  AND2_X1 U16175 ( .A1(n14600), .A2(n14599), .ZN(n14373) );
  OAI21_X1 U16176 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(n14373), .A(n14372), 
        .ZN(n14377) );
  XNOR2_X1 U16177 ( .A(P1_ADDR_REG_14__SCAN_IN), .B(P3_ADDR_REG_14__SCAN_IN), 
        .ZN(n14375) );
  XOR2_X1 U16178 ( .A(n14375), .B(n14374), .Z(n14376) );
  XOR2_X1 U16179 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .Z(n14378) );
  XNOR2_X1 U16180 ( .A(n14379), .B(n14378), .ZN(n14606) );
  AOI21_X2 U16181 ( .B1(n14608), .B2(n14380), .A(n14605), .ZN(n14611) );
  XNOR2_X1 U16182 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(P3_ADDR_REG_16__SCAN_IN), 
        .ZN(n14382) );
  XNOR2_X1 U16183 ( .A(n14382), .B(n14381), .ZN(n14612) );
  NAND2_X1 U16184 ( .A1(n14611), .A2(n14612), .ZN(n14383) );
  NOR2_X1 U16185 ( .A1(n14611), .A2(n14612), .ZN(n14610) );
  AOI21_X2 U16186 ( .B1(n14613), .B2(n14383), .A(n14610), .ZN(n14441) );
  XOR2_X1 U16187 ( .A(n14385), .B(n14384), .Z(n14440) );
  NAND2_X1 U16188 ( .A1(n14441), .A2(n14440), .ZN(n14386) );
  XNOR2_X1 U16189 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14444), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16190 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14387) );
  OAI21_X1 U16191 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14387), 
        .ZN(U28) );
  AOI21_X1 U16192 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14388) );
  OAI21_X1 U16193 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14388), 
        .ZN(U29) );
  AOI21_X1 U16194 ( .B1(n14391), .B2(n14390), .A(n14389), .ZN(n14393) );
  XNOR2_X1 U16195 ( .A(n14393), .B(n14392), .ZN(SUB_1596_U61) );
  XOR2_X1 U16196 ( .A(n14395), .B(n14394), .Z(SUB_1596_U57) );
  AOI22_X1 U16197 ( .A1(n14398), .A2(n14397), .B1(SI_16_), .B2(n14396), .ZN(
        n14399) );
  OAI21_X1 U16198 ( .B1(P3_U3151), .B2(n14400), .A(n14399), .ZN(P3_U3279) );
  XNOR2_X1 U16199 ( .A(n14401), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16200 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14402), .Z(SUB_1596_U54) );
  XOR2_X1 U16201 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14403), .Z(SUB_1596_U70)
         );
  AOI22_X1 U16202 ( .A1(n14745), .A2(n14558), .B1(n14404), .B2(n14766), .ZN(
        n14405) );
  OAI211_X1 U16203 ( .C1(n14407), .C2(n14748), .A(n14406), .B(n14405), .ZN(
        n14408) );
  INV_X1 U16204 ( .A(n14408), .ZN(n14409) );
  OAI211_X1 U16205 ( .C1(n14411), .C2(n14730), .A(n14410), .B(n14409), .ZN(
        n14412) );
  AOI21_X1 U16206 ( .B1(n14733), .B2(n14413), .A(n14412), .ZN(n14415) );
  INV_X1 U16207 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14414) );
  AOI22_X1 U16208 ( .A1(n6444), .A2(n14415), .B1(n14414), .B2(n14775), .ZN(
        P1_U3495) );
  AOI22_X1 U16209 ( .A1(n14790), .A2(n14415), .B1(n9661), .B2(n14787), .ZN(
        P1_U3540) );
  NAND2_X1 U16210 ( .A1(n14416), .A2(n14570), .ZN(n14417) );
  NAND2_X1 U16211 ( .A1(n14418), .A2(n14417), .ZN(n14573) );
  OR2_X1 U16212 ( .A1(n14421), .A2(n14420), .ZN(n14423) );
  NAND2_X1 U16213 ( .A1(n14519), .A2(n14766), .ZN(n14422) );
  NAND2_X1 U16214 ( .A1(n14423), .A2(n14422), .ZN(n14569) );
  INV_X1 U16215 ( .A(n14569), .ZN(n14424) );
  OAI21_X1 U16216 ( .B1(n14518), .B2(n14706), .A(n14424), .ZN(n14425) );
  AOI21_X1 U16217 ( .B1(n14570), .B2(n14426), .A(n14425), .ZN(n14427) );
  OAI21_X1 U16218 ( .B1(n14573), .B2(n14419), .A(n14427), .ZN(n14428) );
  INV_X1 U16219 ( .A(n14428), .ZN(n14438) );
  OAI21_X1 U16220 ( .B1(n14431), .B2(n14430), .A(n14429), .ZN(n14575) );
  INV_X1 U16221 ( .A(n14575), .ZN(n14435) );
  XNOR2_X1 U16222 ( .A(n14432), .B(n14433), .ZN(n14578) );
  AOI22_X1 U16223 ( .A1(n14435), .A2(n14434), .B1(n14544), .B2(n14578), .ZN(
        n14436) );
  OAI221_X1 U16224 ( .B1(n14704), .B2(n14438), .C1(n14437), .C2(n9971), .A(
        n14436), .ZN(P1_U3280) );
  AOI21_X1 U16225 ( .B1(n14441), .B2(n14440), .A(n14439), .ZN(n14443) );
  XNOR2_X1 U16226 ( .A(n14443), .B(n14442), .ZN(SUB_1596_U63) );
  NAND2_X1 U16227 ( .A1(n14447), .A2(n14446), .ZN(n14448) );
  OAI21_X1 U16228 ( .B1(n14449), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n14448), 
        .ZN(n14452) );
  XNOR2_X1 U16229 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14450) );
  XNOR2_X1 U16230 ( .A(n14450), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n14451) );
  AOI21_X1 U16231 ( .B1(n14455), .B2(n14454), .A(n14453), .ZN(n14471) );
  OAI22_X1 U16232 ( .A1(n14457), .A2(n14979), .B1(n14978), .B2(n14456), .ZN(
        n14468) );
  AOI21_X1 U16233 ( .B1(n14460), .B2(n14459), .A(n14458), .ZN(n14466) );
  NOR2_X1 U16234 ( .A1(n14462), .A2(n14461), .ZN(n14463) );
  OAI21_X1 U16235 ( .B1(n14464), .B2(n14463), .A(n14945), .ZN(n14465) );
  OAI21_X1 U16236 ( .B1(n14466), .B2(n14989), .A(n14465), .ZN(n14467) );
  NOR3_X1 U16237 ( .A1(n14469), .A2(n14468), .A3(n14467), .ZN(n14470) );
  OAI21_X1 U16238 ( .B1(n14471), .B2(n14995), .A(n14470), .ZN(P3_U3197) );
  INV_X1 U16239 ( .A(n14472), .ZN(n14473) );
  AOI21_X1 U16240 ( .B1(n14474), .B2(n15007), .A(n14473), .ZN(n14486) );
  INV_X1 U16241 ( .A(n14486), .ZN(n14475) );
  OAI22_X1 U16242 ( .A1(n15064), .A2(n14475), .B1(P3_REG1_REG_30__SCAN_IN), 
        .B2(n15066), .ZN(n14476) );
  INV_X1 U16243 ( .A(n14476), .ZN(P3_U3489) );
  NOR2_X1 U16244 ( .A1(n14477), .A2(n15044), .ZN(n14479) );
  AOI211_X1 U16245 ( .C1(n14480), .C2(n15049), .A(n14479), .B(n14478), .ZN(
        n14488) );
  AOI22_X1 U16246 ( .A1(n15066), .A2(n14488), .B1(n11066), .B2(n15064), .ZN(
        P3_U3471) );
  NOR2_X1 U16247 ( .A1(n14481), .A2(n15044), .ZN(n14483) );
  AOI211_X1 U16248 ( .C1(n14484), .C2(n15049), .A(n14483), .B(n14482), .ZN(
        n14490) );
  AOI22_X1 U16249 ( .A1(n15066), .A2(n14490), .B1(n11003), .B2(n15064), .ZN(
        P3_U3470) );
  AOI22_X1 U16250 ( .A1(n15052), .A2(n14486), .B1(n14485), .B2(n15050), .ZN(
        P3_U3457) );
  INV_X1 U16251 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14487) );
  AOI22_X1 U16252 ( .A1(n15052), .A2(n14488), .B1(n14487), .B2(n15050), .ZN(
        P3_U3426) );
  INV_X1 U16253 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14489) );
  AOI22_X1 U16254 ( .A1(n15052), .A2(n14490), .B1(n14489), .B2(n15050), .ZN(
        P3_U3423) );
  INV_X1 U16255 ( .A(n14491), .ZN(n14496) );
  OAI21_X1 U16256 ( .B1(n14493), .B2(n14864), .A(n14492), .ZN(n14495) );
  AOI211_X1 U16257 ( .C1(n14869), .C2(n14496), .A(n14495), .B(n14494), .ZN(
        n14497) );
  AOI22_X1 U16258 ( .A1(n14885), .A2(n14497), .B1(n15112), .B2(n14883), .ZN(
        P2_U3511) );
  AOI22_X1 U16259 ( .A1(n14880), .A2(n14497), .B1(n7842), .B2(n14879), .ZN(
        P2_U3466) );
  XNOR2_X1 U16260 ( .A(n14498), .B(n14499), .ZN(n14507) );
  NOR2_X1 U16261 ( .A1(n14562), .A2(n14500), .ZN(n14506) );
  OAI22_X1 U16262 ( .A1(n14504), .A2(n14503), .B1(n14502), .B2(n14501), .ZN(
        n14505) );
  AOI211_X1 U16263 ( .C1(n14507), .C2(n14527), .A(n14506), .B(n14505), .ZN(
        n14509) );
  OAI211_X1 U16264 ( .C1(n14628), .C2(n14510), .A(n14509), .B(n14508), .ZN(
        P1_U3215) );
  AND2_X1 U16265 ( .A1(n13708), .A2(n14511), .ZN(n14514) );
  OAI21_X1 U16266 ( .B1(n14514), .B2(n14513), .A(n14512), .ZN(n14515) );
  AOI222_X1 U16267 ( .A1(n14569), .A2(n14625), .B1(n14515), .B2(n14527), .C1(
        n14570), .C2(n14525), .ZN(n14517) );
  OAI211_X1 U16268 ( .C1(n14628), .C2(n14518), .A(n14517), .B(n14516), .ZN(
        P1_U3234) );
  NAND2_X1 U16269 ( .A1(n14519), .A2(n14745), .ZN(n14522) );
  NAND2_X1 U16270 ( .A1(n14520), .A2(n14766), .ZN(n14521) );
  NAND2_X1 U16271 ( .A1(n14522), .A2(n14521), .ZN(n14534) );
  XNOR2_X1 U16272 ( .A(n14524), .B(n14523), .ZN(n14526) );
  AOI222_X1 U16273 ( .A1(n14534), .A2(n14625), .B1(n14527), .B2(n14526), .C1(
        n6612), .C2(n14525), .ZN(n14529) );
  OAI211_X1 U16274 ( .C1(n14628), .C2(n14530), .A(n14529), .B(n14528), .ZN(
        P1_U3236) );
  NOR2_X1 U16275 ( .A1(n14532), .A2(n7384), .ZN(n14533) );
  AOI21_X1 U16276 ( .B1(n14762), .B2(n14533), .A(n14574), .ZN(n14535) );
  AOI21_X1 U16277 ( .B1(n14536), .B2(n14535), .A(n14534), .ZN(n14581) );
  AOI222_X1 U16278 ( .A1(n6612), .A2(n14683), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n14704), .C1(n14682), .C2(n14537), .ZN(n14546) );
  XNOR2_X1 U16279 ( .A(n14539), .B(n14540), .ZN(n14584) );
  OAI211_X1 U16280 ( .C1(n14542), .C2(n14582), .A(n14686), .B(n14541), .ZN(
        n14580) );
  INV_X1 U16281 ( .A(n14580), .ZN(n14543) );
  AOI22_X1 U16282 ( .A1(n14584), .A2(n14544), .B1(n14690), .B2(n14543), .ZN(
        n14545) );
  OAI211_X1 U16283 ( .C1(n14704), .C2(n14581), .A(n14546), .B(n14545), .ZN(
        P1_U3282) );
  AOI22_X1 U16284 ( .A1(n14548), .A2(n14766), .B1(n14745), .B2(n14547), .ZN(
        n14549) );
  OAI211_X1 U16285 ( .C1(n14551), .C2(n14748), .A(n14550), .B(n14549), .ZN(
        n14554) );
  NOR2_X1 U16286 ( .A1(n14552), .A2(n14574), .ZN(n14553) );
  AOI211_X1 U16287 ( .C1(n14774), .C2(n14555), .A(n14554), .B(n14553), .ZN(
        n14587) );
  INV_X1 U16288 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14556) );
  AOI22_X1 U16289 ( .A1(n14790), .A2(n14587), .B1(n14556), .B2(n14787), .ZN(
        P1_U3543) );
  AND2_X1 U16290 ( .A1(n14557), .A2(n14774), .ZN(n14567) );
  AOI22_X1 U16291 ( .A1(n14559), .A2(n14745), .B1(n14766), .B2(n14558), .ZN(
        n14560) );
  OAI211_X1 U16292 ( .C1(n14562), .C2(n14748), .A(n14561), .B(n14560), .ZN(
        n14565) );
  INV_X1 U16293 ( .A(n14563), .ZN(n14564) );
  AOI211_X1 U16294 ( .C1(n14567), .C2(n14566), .A(n14565), .B(n14564), .ZN(
        n14589) );
  AOI22_X1 U16295 ( .A1(n14790), .A2(n14589), .B1(n14568), .B2(n14787), .ZN(
        P1_U3542) );
  AOI21_X1 U16296 ( .B1(n14570), .B2(n14767), .A(n14569), .ZN(n14571) );
  OAI21_X1 U16297 ( .B1(n14573), .B2(n14572), .A(n14571), .ZN(n14577) );
  NOR2_X1 U16298 ( .A1(n14575), .A2(n14574), .ZN(n14576) );
  AOI211_X1 U16299 ( .C1(n14578), .C2(n14774), .A(n14577), .B(n14576), .ZN(
        n14591) );
  AOI22_X1 U16300 ( .A1(n14790), .A2(n14591), .B1(n14579), .B2(n14787), .ZN(
        P1_U3541) );
  OAI211_X1 U16301 ( .C1(n14582), .C2(n14748), .A(n14581), .B(n14580), .ZN(
        n14583) );
  AOI21_X1 U16302 ( .B1(n14584), .B2(n14774), .A(n14583), .ZN(n14593) );
  AOI22_X1 U16303 ( .A1(n14790), .A2(n14593), .B1(n14585), .B2(n14787), .ZN(
        P1_U3539) );
  INV_X1 U16304 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14586) );
  AOI22_X1 U16305 ( .A1(n6444), .A2(n14587), .B1(n14586), .B2(n14775), .ZN(
        P1_U3504) );
  INV_X1 U16306 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14588) );
  AOI22_X1 U16307 ( .A1(n6444), .A2(n14589), .B1(n14588), .B2(n14775), .ZN(
        P1_U3501) );
  INV_X1 U16308 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14590) );
  AOI22_X1 U16309 ( .A1(n6444), .A2(n14591), .B1(n14590), .B2(n14775), .ZN(
        P1_U3498) );
  INV_X1 U16310 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14592) );
  AOI22_X1 U16311 ( .A1(n6444), .A2(n14593), .B1(n14592), .B2(n14775), .ZN(
        P1_U3492) );
  OAI21_X1 U16312 ( .B1(n14596), .B2(n14595), .A(n14594), .ZN(n14597) );
  XNOR2_X1 U16313 ( .A(n14597), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  XNOR2_X1 U16314 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n14598), .ZN(SUB_1596_U68)
         );
  XOR2_X1 U16315 ( .A(n14601), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  NOR2_X1 U16316 ( .A1(n14603), .A2(n14602), .ZN(n14604) );
  XOR2_X1 U16317 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n14604), .Z(SUB_1596_U66)
         );
  AOI21_X1 U16318 ( .B1(n14607), .B2(n14606), .A(n14605), .ZN(n14609) );
  XNOR2_X1 U16319 ( .A(n14609), .B(n14608), .ZN(SUB_1596_U65) );
  AOI21_X1 U16320 ( .B1(n14612), .B2(n14611), .A(n14610), .ZN(n14614) );
  XNOR2_X1 U16321 ( .A(n14614), .B(n14613), .ZN(SUB_1596_U64) );
  NAND2_X1 U16322 ( .A1(n14767), .A2(n14615), .ZN(n14710) );
  INV_X1 U16323 ( .A(n14710), .ZN(n14617) );
  AOI21_X1 U16324 ( .B1(n14618), .B2(n14617), .A(n14616), .ZN(n14627) );
  AOI211_X1 U16325 ( .C1(n14622), .C2(n14621), .A(n14620), .B(n14619), .ZN(
        n14623) );
  AOI21_X1 U16326 ( .B1(n14625), .B2(n14624), .A(n14623), .ZN(n14626) );
  OAI211_X1 U16327 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n14628), .A(n14627), .B(
        n14626), .ZN(P1_U3218) );
  INV_X1 U16328 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n14630) );
  AOI21_X1 U16329 ( .B1(n14631), .B2(n14630), .A(n14629), .ZN(n14632) );
  XNOR2_X1 U16330 ( .A(n14632), .B(P1_IR_REG_0__SCAN_IN), .ZN(n14636) );
  AOI22_X1 U16331 ( .A1(n14633), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14634) );
  OAI21_X1 U16332 ( .B1(n14636), .B2(n14635), .A(n14634), .ZN(P1_U3243) );
  INV_X1 U16333 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14638) );
  OAI21_X1 U16334 ( .B1(n14674), .B2(n14638), .A(n14637), .ZN(n14656) );
  MUX2_X1 U16335 ( .A(n9887), .B(P1_REG2_REG_4__SCAN_IN), .S(n14658), .Z(
        n14641) );
  INV_X1 U16336 ( .A(n14639), .ZN(n14640) );
  NAND2_X1 U16337 ( .A1(n14641), .A2(n14640), .ZN(n14644) );
  OAI211_X1 U16338 ( .C1(n14645), .C2(n14644), .A(n14643), .B(n14642), .ZN(
        n14654) );
  INV_X1 U16339 ( .A(n14646), .ZN(n14651) );
  NAND3_X1 U16340 ( .A1(n14649), .A2(n14648), .A3(n14647), .ZN(n14650) );
  NAND3_X1 U16341 ( .A1(n14652), .A2(n14651), .A3(n14650), .ZN(n14653) );
  NAND2_X1 U16342 ( .A1(n14654), .A2(n14653), .ZN(n14655) );
  AOI211_X1 U16343 ( .C1(n14658), .C2(n14657), .A(n14656), .B(n14655), .ZN(
        n14660) );
  NAND2_X1 U16344 ( .A1(n14660), .A2(n14659), .ZN(P1_U3247) );
  AOI21_X1 U16345 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n14662), .A(n14661), 
        .ZN(n14667) );
  AOI21_X1 U16346 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14664), .A(n14663), 
        .ZN(n14665) );
  OAI222_X1 U16347 ( .A1(n14670), .A2(n14669), .B1(n14668), .B2(n14667), .C1(
        n14666), .C2(n14665), .ZN(n14671) );
  INV_X1 U16348 ( .A(n14671), .ZN(n14673) );
  OAI211_X1 U16349 ( .C1(n14675), .C2(n14674), .A(n14673), .B(n14672), .ZN(
        P1_U3258) );
  XNOR2_X1 U16350 ( .A(n14676), .B(n14677), .ZN(n14740) );
  INV_X1 U16351 ( .A(n14736), .ZN(n14680) );
  XNOR2_X1 U16352 ( .A(n14678), .B(n14677), .ZN(n14679) );
  AND2_X1 U16353 ( .A1(n14679), .A2(n14763), .ZN(n14738) );
  AOI211_X1 U16354 ( .C1(n14733), .C2(n14740), .A(n14680), .B(n14738), .ZN(
        n14694) );
  AOI222_X1 U16355 ( .A1(n14684), .A2(n14683), .B1(P1_REG2_REG_7__SCAN_IN), 
        .B2(n14704), .C1(n14682), .C2(n14681), .ZN(n14693) );
  OAI211_X1 U16356 ( .C1(n14688), .C2(n14687), .A(n14686), .B(n14685), .ZN(
        n14737) );
  INV_X1 U16357 ( .A(n14737), .ZN(n14689) );
  AOI22_X1 U16358 ( .A1(n14740), .A2(n14691), .B1(n14690), .B2(n14689), .ZN(
        n14692) );
  OAI211_X1 U16359 ( .C1(n14704), .C2(n14694), .A(n14693), .B(n14692), .ZN(
        P1_U3286) );
  INV_X1 U16360 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n15110) );
  OAI21_X1 U16361 ( .B1(n14697), .B2(n14696), .A(n14695), .ZN(n14703) );
  INV_X1 U16362 ( .A(n14698), .ZN(n14699) );
  AOI21_X1 U16363 ( .B1(n14701), .B2(n14700), .A(n14699), .ZN(n14702) );
  AOI221_X1 U16364 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n14704), .C1(n14703), 
        .C2(n14437), .A(n14702), .ZN(n14705) );
  OAI21_X1 U16365 ( .B1(n15110), .B2(n14706), .A(n14705), .ZN(P1_U3293) );
  AND2_X1 U16366 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14708), .ZN(P1_U3294) );
  AND2_X1 U16367 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14708), .ZN(P1_U3295) );
  AND2_X1 U16368 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14708), .ZN(P1_U3296) );
  AND2_X1 U16369 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14708), .ZN(P1_U3297) );
  AND2_X1 U16370 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14708), .ZN(P1_U3298) );
  INV_X1 U16371 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n15204) );
  NOR2_X1 U16372 ( .A1(n14707), .A2(n15204), .ZN(P1_U3299) );
  AND2_X1 U16373 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14708), .ZN(P1_U3300) );
  AND2_X1 U16374 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14708), .ZN(P1_U3301) );
  AND2_X1 U16375 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14708), .ZN(P1_U3302) );
  AND2_X1 U16376 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14708), .ZN(P1_U3303) );
  AND2_X1 U16377 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14708), .ZN(P1_U3304) );
  AND2_X1 U16378 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14708), .ZN(P1_U3305) );
  AND2_X1 U16379 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14708), .ZN(P1_U3306) );
  AND2_X1 U16380 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14708), .ZN(P1_U3307) );
  AND2_X1 U16381 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14708), .ZN(P1_U3308) );
  AND2_X1 U16382 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14708), .ZN(P1_U3309) );
  AND2_X1 U16383 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14708), .ZN(P1_U3310) );
  AND2_X1 U16384 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14708), .ZN(P1_U3311) );
  AND2_X1 U16385 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14708), .ZN(P1_U3312) );
  AND2_X1 U16386 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14708), .ZN(P1_U3313) );
  AND2_X1 U16387 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14708), .ZN(P1_U3314) );
  AND2_X1 U16388 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14708), .ZN(P1_U3315) );
  AND2_X1 U16389 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14708), .ZN(P1_U3316) );
  INV_X1 U16390 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15173) );
  NOR2_X1 U16391 ( .A1(n14707), .A2(n15173), .ZN(P1_U3317) );
  AND2_X1 U16392 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14708), .ZN(P1_U3318) );
  AND2_X1 U16393 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14708), .ZN(P1_U3319) );
  AND2_X1 U16394 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14708), .ZN(P1_U3320) );
  AND2_X1 U16395 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14708), .ZN(P1_U3321) );
  AND2_X1 U16396 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14708), .ZN(P1_U3322) );
  AND2_X1 U16397 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14708), .ZN(P1_U3323) );
  NAND2_X1 U16398 ( .A1(n14709), .A2(n14774), .ZN(n14713) );
  NAND4_X1 U16399 ( .A1(n14713), .A2(n14712), .A3(n14711), .A4(n14710), .ZN(
        n14714) );
  AOI21_X1 U16400 ( .B1(n14715), .B2(n14763), .A(n14714), .ZN(n14777) );
  INV_X1 U16401 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14716) );
  AOI22_X1 U16402 ( .A1(n6444), .A2(n14777), .B1(n14716), .B2(n14775), .ZN(
        P1_U3468) );
  INV_X1 U16403 ( .A(n14717), .ZN(n14723) );
  OR4_X1 U16404 ( .A1(n14721), .A2(n14720), .A3(n14719), .A4(n14718), .ZN(
        n14722) );
  AOI21_X1 U16405 ( .B1(n14723), .B2(n14774), .A(n14722), .ZN(n14779) );
  INV_X1 U16406 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14724) );
  AOI22_X1 U16407 ( .A1(n6444), .A2(n14779), .B1(n14724), .B2(n14775), .ZN(
        P1_U3471) );
  INV_X1 U16408 ( .A(n14729), .ZN(n14732) );
  AOI211_X1 U16409 ( .C1(n14727), .C2(n14767), .A(n14726), .B(n14725), .ZN(
        n14728) );
  OAI21_X1 U16410 ( .B1(n14730), .B2(n14729), .A(n14728), .ZN(n14731) );
  AOI21_X1 U16411 ( .B1(n14733), .B2(n14732), .A(n14731), .ZN(n14781) );
  INV_X1 U16412 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14734) );
  AOI22_X1 U16413 ( .A1(n6444), .A2(n14781), .B1(n14734), .B2(n14775), .ZN(
        P1_U3477) );
  NAND3_X1 U16414 ( .A1(n14737), .A2(n14736), .A3(n14735), .ZN(n14739) );
  AOI211_X1 U16415 ( .C1(n14740), .C2(n14774), .A(n14739), .B(n14738), .ZN(
        n14783) );
  INV_X1 U16416 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14741) );
  AOI22_X1 U16417 ( .A1(n6444), .A2(n14783), .B1(n14741), .B2(n14775), .ZN(
        P1_U3480) );
  INV_X1 U16418 ( .A(n14742), .ZN(n14753) );
  INV_X1 U16419 ( .A(n14743), .ZN(n14747) );
  AOI22_X1 U16420 ( .A1(n14745), .A2(n14765), .B1(n14744), .B2(n14766), .ZN(
        n14746) );
  OAI211_X1 U16421 ( .C1(n14749), .C2(n14748), .A(n14747), .B(n14746), .ZN(
        n14752) );
  INV_X1 U16422 ( .A(n14750), .ZN(n14751) );
  AOI211_X1 U16423 ( .C1(n14753), .C2(n14774), .A(n14752), .B(n14751), .ZN(
        n14784) );
  INV_X1 U16424 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14754) );
  AOI22_X1 U16425 ( .A1(n6444), .A2(n14784), .B1(n14754), .B2(n14775), .ZN(
        P1_U3483) );
  NOR2_X1 U16426 ( .A1(n14756), .A2(n14755), .ZN(n14760) );
  NOR4_X1 U16427 ( .A1(n14760), .A2(n14759), .A3(n14758), .A4(n14757), .ZN(
        n14786) );
  INV_X1 U16428 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14761) );
  AOI22_X1 U16429 ( .A1(n6444), .A2(n14786), .B1(n14761), .B2(n14775), .ZN(
        P1_U3486) );
  NAND3_X1 U16430 ( .A1(n14764), .A2(n14763), .A3(n14762), .ZN(n14771) );
  AOI22_X1 U16431 ( .A1(n14768), .A2(n14767), .B1(n14766), .B2(n14765), .ZN(
        n14769) );
  NAND3_X1 U16432 ( .A1(n14771), .A2(n14770), .A3(n14769), .ZN(n14772) );
  AOI21_X1 U16433 ( .B1(n14774), .B2(n14773), .A(n14772), .ZN(n14789) );
  INV_X1 U16434 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14776) );
  AOI22_X1 U16435 ( .A1(n6444), .A2(n14789), .B1(n14776), .B2(n14775), .ZN(
        P1_U3489) );
  AOI22_X1 U16436 ( .A1(n14790), .A2(n14777), .B1(n9309), .B2(n14787), .ZN(
        P1_U3531) );
  AOI22_X1 U16437 ( .A1(n14790), .A2(n14779), .B1(n14778), .B2(n14787), .ZN(
        P1_U3532) );
  AOI22_X1 U16438 ( .A1(n14790), .A2(n14781), .B1(n14780), .B2(n14787), .ZN(
        P1_U3534) );
  AOI22_X1 U16439 ( .A1(n14790), .A2(n14783), .B1(n14782), .B2(n14787), .ZN(
        P1_U3535) );
  AOI22_X1 U16440 ( .A1(n14790), .A2(n14784), .B1(n9352), .B2(n14787), .ZN(
        P1_U3536) );
  AOI22_X1 U16441 ( .A1(n14790), .A2(n14786), .B1(n14785), .B2(n14787), .ZN(
        P1_U3537) );
  AOI22_X1 U16442 ( .A1(n14790), .A2(n14789), .B1(n14788), .B2(n14787), .ZN(
        P1_U3538) );
  NOR2_X1 U16443 ( .A1(n14820), .A2(P2_U3947), .ZN(P2_U3087) );
  INV_X1 U16444 ( .A(n14791), .ZN(n14793) );
  OAI21_X1 U16445 ( .B1(n14793), .B2(n14792), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14794) );
  OAI21_X1 U16446 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n14794), .ZN(n14804) );
  OAI211_X1 U16447 ( .C1(n14797), .C2(n14796), .A(n14824), .B(n14795), .ZN(
        n14803) );
  OAI211_X1 U16448 ( .C1(n14800), .C2(n14799), .A(n14827), .B(n14798), .ZN(
        n14802) );
  NAND2_X1 U16449 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n14820), .ZN(n14801) );
  NAND4_X1 U16450 ( .A1(n14804), .A2(n14803), .A3(n14802), .A4(n14801), .ZN(
        P2_U3220) );
  AOI22_X1 U16451 ( .A1(n14820), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n14819) );
  NAND2_X1 U16452 ( .A1(n14822), .A2(n14805), .ZN(n14818) );
  AOI21_X1 U16453 ( .B1(n14808), .B2(n14807), .A(n14806), .ZN(n14810) );
  NAND2_X1 U16454 ( .A1(n14810), .A2(n14809), .ZN(n14817) );
  AOI211_X1 U16455 ( .C1(n14814), .C2(n14813), .A(n14812), .B(n14811), .ZN(
        n14815) );
  INV_X1 U16456 ( .A(n14815), .ZN(n14816) );
  NAND4_X1 U16457 ( .A1(n14819), .A2(n14818), .A3(n14817), .A4(n14816), .ZN(
        P2_U3227) );
  AOI22_X1 U16458 ( .A1(n14820), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14832) );
  NAND2_X1 U16459 ( .A1(n14822), .A2(n14821), .ZN(n14831) );
  OAI211_X1 U16460 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n14825), .A(n14824), 
        .B(n14823), .ZN(n14830) );
  OAI211_X1 U16461 ( .C1(n14828), .C2(P2_REG1_REG_15__SCAN_IN), .A(n14827), 
        .B(n14826), .ZN(n14829) );
  NAND4_X1 U16462 ( .A1(n14832), .A2(n14831), .A3(n14830), .A4(n14829), .ZN(
        P2_U3229) );
  NAND2_X1 U16463 ( .A1(n14834), .A2(n14833), .ZN(n14838) );
  INV_X1 U16464 ( .A(n14835), .ZN(n14836) );
  AOI22_X1 U16465 ( .A1(n15079), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n14836), 
        .B2(n15071), .ZN(n14837) );
  OAI211_X1 U16466 ( .C1(n14840), .C2(n14839), .A(n14838), .B(n14837), .ZN(
        n14841) );
  AOI21_X1 U16467 ( .B1(n14843), .B2(n14842), .A(n14841), .ZN(n14844) );
  OAI21_X1 U16468 ( .B1(n15079), .B2(n14845), .A(n14844), .ZN(P2_U3258) );
  AND2_X1 U16469 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14848), .ZN(P2_U3266) );
  INV_X1 U16470 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15149) );
  NOR2_X1 U16471 ( .A1(n14847), .A2(n15149), .ZN(P2_U3267) );
  INV_X1 U16472 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15143) );
  NOR2_X1 U16473 ( .A1(n14847), .A2(n15143), .ZN(P2_U3268) );
  AND2_X1 U16474 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14848), .ZN(P2_U3269) );
  AND2_X1 U16475 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14848), .ZN(P2_U3270) );
  AND2_X1 U16476 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14848), .ZN(P2_U3271) );
  AND2_X1 U16477 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14848), .ZN(P2_U3272) );
  AND2_X1 U16478 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14848), .ZN(P2_U3273) );
  AND2_X1 U16479 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14848), .ZN(P2_U3274) );
  AND2_X1 U16480 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14848), .ZN(P2_U3275) );
  AND2_X1 U16481 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14848), .ZN(P2_U3276) );
  AND2_X1 U16482 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14848), .ZN(P2_U3277) );
  AND2_X1 U16483 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14848), .ZN(P2_U3278) );
  AND2_X1 U16484 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14848), .ZN(P2_U3279) );
  AND2_X1 U16485 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14848), .ZN(P2_U3280) );
  AND2_X1 U16486 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14848), .ZN(P2_U3281) );
  INV_X1 U16487 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15187) );
  NOR2_X1 U16488 ( .A1(n14847), .A2(n15187), .ZN(P2_U3282) );
  AND2_X1 U16489 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14848), .ZN(P2_U3283) );
  AND2_X1 U16490 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14848), .ZN(P2_U3284) );
  AND2_X1 U16491 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14848), .ZN(P2_U3285) );
  AND2_X1 U16492 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14848), .ZN(P2_U3286) );
  AND2_X1 U16493 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14848), .ZN(P2_U3287) );
  AND2_X1 U16494 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14848), .ZN(P2_U3288) );
  AND2_X1 U16495 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14848), .ZN(P2_U3289) );
  AND2_X1 U16496 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14848), .ZN(P2_U3290) );
  AND2_X1 U16497 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14848), .ZN(P2_U3291) );
  AND2_X1 U16498 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14848), .ZN(P2_U3292) );
  AND2_X1 U16499 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14848), .ZN(P2_U3293) );
  AND2_X1 U16500 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14848), .ZN(P2_U3294) );
  AND2_X1 U16501 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14848), .ZN(P2_U3295) );
  AOI22_X1 U16502 ( .A1(n14854), .A2(n14850), .B1(n14849), .B2(n14851), .ZN(
        P2_U3416) );
  AOI22_X1 U16503 ( .A1(n14854), .A2(n14853), .B1(n14852), .B2(n14851), .ZN(
        P2_U3417) );
  NOR2_X1 U16504 ( .A1(n14855), .A2(n14876), .ZN(n14858) );
  INV_X1 U16505 ( .A(n14856), .ZN(n14857) );
  AOI211_X1 U16506 ( .C1(n14860), .C2(n14859), .A(n14858), .B(n14857), .ZN(
        n14881) );
  INV_X1 U16507 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14861) );
  AOI22_X1 U16508 ( .A1(n14880), .A2(n14881), .B1(n14861), .B2(n14879), .ZN(
        P2_U3430) );
  INV_X1 U16509 ( .A(n14862), .ZN(n14868) );
  OAI21_X1 U16510 ( .B1(n14865), .B2(n14864), .A(n14863), .ZN(n14867) );
  AOI211_X1 U16511 ( .C1(n14869), .C2(n14868), .A(n14867), .B(n14866), .ZN(
        n14882) );
  INV_X1 U16512 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14870) );
  AOI22_X1 U16513 ( .A1(n14880), .A2(n14882), .B1(n14870), .B2(n14879), .ZN(
        P2_U3436) );
  AOI21_X1 U16514 ( .B1(n14873), .B2(n14872), .A(n14871), .ZN(n14874) );
  OAI211_X1 U16515 ( .C1(n14877), .C2(n14876), .A(n14875), .B(n14874), .ZN(
        n14878) );
  INV_X1 U16516 ( .A(n14878), .ZN(n14884) );
  AOI22_X1 U16517 ( .A1(n14880), .A2(n14884), .B1(n7704), .B2(n14879), .ZN(
        P2_U3442) );
  AOI22_X1 U16518 ( .A1(n14885), .A2(n14881), .B1(n9526), .B2(n14883), .ZN(
        P2_U3499) );
  AOI22_X1 U16519 ( .A1(n14885), .A2(n14882), .B1(n9427), .B2(n14883), .ZN(
        P2_U3501) );
  AOI22_X1 U16520 ( .A1(n14885), .A2(n14884), .B1(n9433), .B2(n14883), .ZN(
        P2_U3503) );
  NOR2_X1 U16521 ( .A1(P3_U3897), .A2(n14972), .ZN(P3_U3150) );
  OR2_X1 U16522 ( .A1(n14887), .A2(n14886), .ZN(n14890) );
  NAND2_X1 U16523 ( .A1(n14888), .A2(n10042), .ZN(n14889) );
  OAI211_X1 U16524 ( .C1(n14892), .C2(n14891), .A(n14890), .B(n14889), .ZN(
        n14893) );
  INV_X1 U16525 ( .A(n14893), .ZN(n14894) );
  OAI21_X1 U16526 ( .B1(n14895), .B2(n8190), .A(n14894), .ZN(P3_U3172) );
  AOI22_X1 U16527 ( .A1(n14944), .A2(P3_IR_REG_0__SCAN_IN), .B1(n14972), .B2(
        P3_ADDR_REG_0__SCAN_IN), .ZN(n14903) );
  NOR3_X1 U16528 ( .A1(n14897), .A2(n14896), .A3(n14945), .ZN(n14901) );
  AOI21_X1 U16529 ( .B1(n15107), .B2(n14899), .A(n14898), .ZN(n14900) );
  OR2_X1 U16530 ( .A1(n14901), .A2(n14900), .ZN(n14902) );
  OAI211_X1 U16531 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n8190), .A(n14903), .B(
        n14902), .ZN(P3_U3182) );
  XNOR2_X1 U16532 ( .A(n14905), .B(n14904), .ZN(n14915) );
  NOR2_X1 U16533 ( .A1(n14979), .A2(n14906), .ZN(n14914) );
  AOI21_X1 U16534 ( .B1(n14908), .B2(n10563), .A(n14907), .ZN(n14912) );
  AOI21_X1 U16535 ( .B1(n14910), .B2(n15055), .A(n14909), .ZN(n14911) );
  OAI22_X1 U16536 ( .A1(n14912), .A2(n14995), .B1(n14989), .B2(n14911), .ZN(
        n14913) );
  AOI211_X1 U16537 ( .C1(n14915), .C2(n14945), .A(n14914), .B(n14913), .ZN(
        n14917) );
  OAI211_X1 U16538 ( .C1(n14918), .C2(n14978), .A(n14917), .B(n14916), .ZN(
        P3_U3185) );
  OAI21_X1 U16539 ( .B1(n14921), .B2(n14920), .A(n14919), .ZN(n14932) );
  NOR2_X1 U16540 ( .A1(n14979), .A2(n14922), .ZN(n14931) );
  AOI21_X1 U16541 ( .B1(n14925), .B2(n14924), .A(n14923), .ZN(n14929) );
  AOI21_X1 U16542 ( .B1(n14927), .B2(n8268), .A(n14926), .ZN(n14928) );
  OAI22_X1 U16543 ( .A1(n14929), .A2(n14995), .B1(n14989), .B2(n14928), .ZN(
        n14930) );
  AOI211_X1 U16544 ( .C1(n14932), .C2(n14945), .A(n14931), .B(n14930), .ZN(
        n14934) );
  OAI211_X1 U16545 ( .C1(n14935), .C2(n14978), .A(n14934), .B(n14933), .ZN(
        P3_U3187) );
  INV_X1 U16546 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n14953) );
  AOI21_X1 U16547 ( .B1(n8301), .B2(n14937), .A(n14936), .ZN(n14949) );
  AOI21_X1 U16548 ( .B1(n8296), .B2(n14939), .A(n14938), .ZN(n14940) );
  OR2_X1 U16549 ( .A1(n14940), .A2(n14995), .ZN(n14948) );
  OAI21_X1 U16550 ( .B1(n14943), .B2(n14942), .A(n14941), .ZN(n14946) );
  AOI22_X1 U16551 ( .A1(n14946), .A2(n14945), .B1(n14944), .B2(n7145), .ZN(
        n14947) );
  OAI211_X1 U16552 ( .C1(n14949), .C2(n14989), .A(n14948), .B(n14947), .ZN(
        n14950) );
  INV_X1 U16553 ( .A(n14950), .ZN(n14952) );
  OAI211_X1 U16554 ( .C1(n14953), .C2(n14978), .A(n14952), .B(n14951), .ZN(
        P3_U3189) );
  INV_X1 U16555 ( .A(n14954), .ZN(n14955) );
  AOI21_X1 U16556 ( .B1(n14957), .B2(n14956), .A(n14955), .ZN(n14974) );
  INV_X1 U16557 ( .A(n14958), .ZN(n14959) );
  AOI21_X1 U16558 ( .B1(n14961), .B2(n14960), .A(n14959), .ZN(n14963) );
  OAI21_X1 U16559 ( .B1(n14963), .B2(n14989), .A(n14962), .ZN(n14971) );
  AOI21_X1 U16560 ( .B1(n14966), .B2(n14965), .A(n14964), .ZN(n14969) );
  INV_X1 U16561 ( .A(n14967), .ZN(n14968) );
  OAI22_X1 U16562 ( .A1(n14969), .A2(n14987), .B1(n14968), .B2(n14979), .ZN(
        n14970) );
  AOI211_X1 U16563 ( .C1(n14972), .C2(P3_ADDR_REG_10__SCAN_IN), .A(n14971), 
        .B(n14970), .ZN(n14973) );
  OAI21_X1 U16564 ( .B1(n14974), .B2(n14995), .A(n14973), .ZN(P3_U3192) );
  AOI21_X1 U16565 ( .B1(n12849), .B2(n14976), .A(n14975), .ZN(n14996) );
  OAI22_X1 U16566 ( .A1(n14980), .A2(n14979), .B1(n14978), .B2(n14977), .ZN(
        n14992) );
  AOI21_X1 U16567 ( .B1(n14983), .B2(n14982), .A(n14981), .ZN(n14990) );
  AOI21_X1 U16568 ( .B1(n14986), .B2(n14985), .A(n14984), .ZN(n14988) );
  OAI22_X1 U16569 ( .A1(n14990), .A2(n14989), .B1(n14988), .B2(n14987), .ZN(
        n14991) );
  NOR3_X1 U16570 ( .A1(n14993), .A2(n14992), .A3(n14991), .ZN(n14994) );
  OAI21_X1 U16571 ( .B1(n14996), .B2(n14995), .A(n14994), .ZN(P3_U3195) );
  INV_X1 U16572 ( .A(n14997), .ZN(n15000) );
  AOI211_X1 U16573 ( .C1(n15036), .C2(n15000), .A(n14999), .B(n14998), .ZN(
        n15053) );
  AOI22_X1 U16574 ( .A1(n15052), .A2(n15053), .B1(n8206), .B2(n15050), .ZN(
        P3_U3393) );
  INV_X1 U16575 ( .A(n15001), .ZN(n15004) );
  AOI211_X1 U16576 ( .C1(n15004), .C2(n15036), .A(n15003), .B(n15002), .ZN(
        n15054) );
  INV_X1 U16577 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15005) );
  AOI22_X1 U16578 ( .A1(n15052), .A2(n15054), .B1(n15005), .B2(n15050), .ZN(
        P3_U3396) );
  AOI22_X1 U16579 ( .A1(n15008), .A2(n15036), .B1(n15007), .B2(n15006), .ZN(
        n15009) );
  AND2_X1 U16580 ( .A1(n15010), .A2(n15009), .ZN(n15056) );
  INV_X1 U16581 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15011) );
  AOI22_X1 U16582 ( .A1(n15052), .A2(n15056), .B1(n15011), .B2(n15050), .ZN(
        P3_U3399) );
  OAI22_X1 U16583 ( .A1(n15013), .A2(n15039), .B1(n15044), .B2(n15012), .ZN(
        n15014) );
  NOR2_X1 U16584 ( .A1(n15015), .A2(n15014), .ZN(n15057) );
  INV_X1 U16585 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15016) );
  AOI22_X1 U16586 ( .A1(n15052), .A2(n15057), .B1(n15016), .B2(n15050), .ZN(
        P3_U3402) );
  NOR2_X1 U16587 ( .A1(n15017), .A2(n15044), .ZN(n15019) );
  AOI211_X1 U16588 ( .C1(n15020), .C2(n15036), .A(n15019), .B(n15018), .ZN(
        n15058) );
  INV_X1 U16589 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15021) );
  AOI22_X1 U16590 ( .A1(n15052), .A2(n15058), .B1(n15021), .B2(n15050), .ZN(
        P3_U3405) );
  NOR2_X1 U16591 ( .A1(n15022), .A2(n15044), .ZN(n15024) );
  AOI211_X1 U16592 ( .C1(n15025), .C2(n15036), .A(n15024), .B(n15023), .ZN(
        n15059) );
  INV_X1 U16593 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15026) );
  AOI22_X1 U16594 ( .A1(n15052), .A2(n15059), .B1(n15026), .B2(n15050), .ZN(
        P3_U3408) );
  OAI22_X1 U16595 ( .A1(n15028), .A2(n15039), .B1(n15044), .B2(n15027), .ZN(
        n15029) );
  NOR2_X1 U16596 ( .A1(n15030), .A2(n15029), .ZN(n15060) );
  INV_X1 U16597 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15031) );
  AOI22_X1 U16598 ( .A1(n15052), .A2(n15060), .B1(n15031), .B2(n15050), .ZN(
        P3_U3411) );
  NOR2_X1 U16599 ( .A1(n15032), .A2(n15044), .ZN(n15034) );
  AOI211_X1 U16600 ( .C1(n15036), .C2(n15035), .A(n15034), .B(n15033), .ZN(
        n15061) );
  INV_X1 U16601 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15037) );
  AOI22_X1 U16602 ( .A1(n15052), .A2(n15061), .B1(n15037), .B2(n15050), .ZN(
        P3_U3414) );
  OAI22_X1 U16603 ( .A1(n15040), .A2(n15039), .B1(n15044), .B2(n15038), .ZN(
        n15041) );
  NOR2_X1 U16604 ( .A1(n15042), .A2(n15041), .ZN(n15063) );
  INV_X1 U16605 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15043) );
  AOI22_X1 U16606 ( .A1(n15052), .A2(n15063), .B1(n15043), .B2(n15050), .ZN(
        P3_U3417) );
  NOR2_X1 U16607 ( .A1(n15045), .A2(n15044), .ZN(n15047) );
  AOI211_X1 U16608 ( .C1(n15049), .C2(n15048), .A(n15047), .B(n15046), .ZN(
        n15065) );
  INV_X1 U16609 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15051) );
  AOI22_X1 U16610 ( .A1(n15052), .A2(n15065), .B1(n15051), .B2(n15050), .ZN(
        P3_U3420) );
  AOI22_X1 U16611 ( .A1(n15066), .A2(n15053), .B1(n9774), .B2(n15064), .ZN(
        P3_U3460) );
  AOI22_X1 U16612 ( .A1(n15066), .A2(n15054), .B1(n9923), .B2(n15064), .ZN(
        P3_U3461) );
  AOI22_X1 U16613 ( .A1(n15066), .A2(n15056), .B1(n15055), .B2(n15064), .ZN(
        P3_U3462) );
  AOI22_X1 U16614 ( .A1(n15066), .A2(n15057), .B1(n9925), .B2(n15064), .ZN(
        P3_U3463) );
  AOI22_X1 U16615 ( .A1(n15066), .A2(n15058), .B1(n8268), .B2(n15064), .ZN(
        P3_U3464) );
  AOI22_X1 U16616 ( .A1(n15066), .A2(n15059), .B1(n10188), .B2(n15064), .ZN(
        P3_U3465) );
  AOI22_X1 U16617 ( .A1(n15066), .A2(n15060), .B1(n8301), .B2(n15064), .ZN(
        P3_U3466) );
  AOI22_X1 U16618 ( .A1(n15066), .A2(n15061), .B1(n10522), .B2(n15064), .ZN(
        P3_U3467) );
  AOI22_X1 U16619 ( .A1(n15066), .A2(n15063), .B1(n15062), .B2(n15064), .ZN(
        P3_U3468) );
  AOI22_X1 U16620 ( .A1(n15066), .A2(n15065), .B1(n10997), .B2(n15064), .ZN(
        P3_U3469) );
  INV_X1 U16621 ( .A(n15067), .ZN(n15073) );
  AOI22_X1 U16622 ( .A1(n15071), .A2(n15070), .B1(n15069), .B2(n15068), .ZN(
        n15072) );
  OAI21_X1 U16623 ( .B1(n15073), .B2(n6689), .A(n15072), .ZN(n15075) );
  AOI211_X1 U16624 ( .C1(n15077), .C2(n15076), .A(n15075), .B(n15074), .ZN(
        n15078) );
  AOI22_X1 U16625 ( .A1(n15079), .A2(n9461), .B1(n15078), .B2(n13490), .ZN(
        n15238) );
  NOR4_X1 U16626 ( .A1(n15080), .A2(P1_IR_REG_25__SCAN_IN), .A3(
        P2_IR_REG_20__SCAN_IN), .A4(P1_REG0_REG_25__SCAN_IN), .ZN(n15084) );
  INV_X1 U16627 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n15193) );
  NAND4_X1 U16628 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n15189), .A3(n15186), 
        .A4(n15193), .ZN(n15081) );
  NOR3_X1 U16629 ( .A1(n15192), .A2(n15082), .A3(n15081), .ZN(n15083) );
  NAND4_X1 U16630 ( .A1(n15084), .A2(P2_IR_REG_29__SCAN_IN), .A3(
        P2_REG2_REG_31__SCAN_IN), .A4(n15083), .ZN(n15086) );
  NAND4_X1 U16631 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), 
        .A3(P2_D_REG_15__SCAN_IN), .A4(n15149), .ZN(n15085) );
  NOR2_X1 U16632 ( .A1(n15086), .A2(n15085), .ZN(n15105) );
  NOR4_X1 U16633 ( .A1(SI_22_), .A2(P1_REG2_REG_14__SCAN_IN), .A3(n15087), 
        .A4(n15221), .ZN(n15104) );
  NOR4_X1 U16634 ( .A1(n15172), .A2(n14782), .A3(P2_REG3_REG_11__SCAN_IN), 
        .A4(P3_REG2_REG_1__SCAN_IN), .ZN(n15090) );
  NAND4_X1 U16635 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P2_REG1_REG_14__SCAN_IN), 
        .A3(P1_REG2_REG_16__SCAN_IN), .A4(n15218), .ZN(n15088) );
  NOR3_X1 U16636 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_DATAO_REG_4__SCAN_IN), 
        .A3(n15088), .ZN(n15089) );
  AND4_X1 U16637 ( .A1(n15090), .A2(P3_D_REG_1__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(n15089), .ZN(n15103) );
  NAND4_X1 U16638 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(
        P3_DATAO_REG_17__SCAN_IN), .A3(P3_DATAO_REG_31__SCAN_IN), .A4(n15122), 
        .ZN(n15101) );
  NOR4_X1 U16639 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .A3(n13268), .A4(n15207), .ZN(n15093) );
  NOR3_X1 U16640 ( .A1(P3_DATAO_REG_30__SCAN_IN), .A2(n15130), .A3(n15133), 
        .ZN(n15092) );
  NOR4_X1 U16641 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P2_DATAO_REG_13__SCAN_IN), 
        .A3(P1_REG3_REG_0__SCAN_IN), .A4(P1_ADDR_REG_14__SCAN_IN), .ZN(n15091)
         );
  NAND4_X1 U16642 ( .A1(P3_D_REG_11__SCAN_IN), .A2(n15093), .A3(n15092), .A4(
        n15091), .ZN(n15100) );
  NAND4_X1 U16643 ( .A1(P3_D_REG_28__SCAN_IN), .A2(P3_REG2_REG_17__SCAN_IN), 
        .A3(P2_REG0_REG_14__SCAN_IN), .A4(P1_REG2_REG_0__SCAN_IN), .ZN(n15099)
         );
  NOR3_X1 U16644 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_20__SCAN_IN), 
        .A3(P2_REG1_REG_12__SCAN_IN), .ZN(n15097) );
  INV_X1 U16645 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n15158) );
  NOR4_X1 U16646 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(P2_DATAO_REG_20__SCAN_IN), 
        .A3(n15159), .A4(n15158), .ZN(n15096) );
  NOR4_X1 U16647 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P2_REG0_REG_30__SCAN_IN), .A4(n15094), .ZN(n15095) );
  NAND4_X1 U16648 ( .A1(P1_REG2_REG_25__SCAN_IN), .A2(n15097), .A3(n15096), 
        .A4(n15095), .ZN(n15098) );
  NOR4_X1 U16649 ( .A1(n15101), .A2(n15100), .A3(n15099), .A4(n15098), .ZN(
        n15102) );
  NAND4_X1 U16650 ( .A1(n15105), .A2(n15104), .A3(n15103), .A4(n15102), .ZN(
        n15236) );
  AOI22_X1 U16651 ( .A1(n15108), .A2(keyinput12), .B1(n15107), .B2(keyinput21), 
        .ZN(n15106) );
  OAI221_X1 U16652 ( .B1(n15108), .B2(keyinput12), .C1(n15107), .C2(keyinput21), .A(n15106), .ZN(n15120) );
  AOI22_X1 U16653 ( .A1(n15111), .A2(keyinput60), .B1(keyinput9), .B2(n15110), 
        .ZN(n15109) );
  OAI221_X1 U16654 ( .B1(n15111), .B2(keyinput60), .C1(n15110), .C2(keyinput9), 
        .A(n15109), .ZN(n15119) );
  XOR2_X1 U16655 ( .A(n15112), .B(keyinput30), .Z(n15117) );
  INV_X1 U16656 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n15113) );
  XOR2_X1 U16657 ( .A(n15113), .B(keyinput51), .Z(n15116) );
  XNOR2_X1 U16658 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput28), .ZN(n15115) );
  XNOR2_X1 U16659 ( .A(P3_IR_REG_31__SCAN_IN), .B(keyinput11), .ZN(n15114) );
  NAND4_X1 U16660 ( .A1(n15117), .A2(n15116), .A3(n15115), .A4(n15114), .ZN(
        n15118) );
  NOR3_X1 U16661 ( .A1(n15120), .A2(n15119), .A3(n15118), .ZN(n15170) );
  AOI22_X1 U16662 ( .A1(n15082), .A2(keyinput17), .B1(n15122), .B2(keyinput6), 
        .ZN(n15121) );
  OAI221_X1 U16663 ( .B1(n15082), .B2(keyinput17), .C1(n15122), .C2(keyinput6), 
        .A(n15121), .ZN(n15127) );
  XNOR2_X1 U16664 ( .A(n15123), .B(keyinput37), .ZN(n15126) );
  XNOR2_X1 U16665 ( .A(n15124), .B(keyinput22), .ZN(n15125) );
  OR3_X1 U16666 ( .A1(n15127), .A2(n15126), .A3(n15125), .ZN(n15136) );
  INV_X1 U16667 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n15129) );
  AOI22_X1 U16668 ( .A1(n15130), .A2(keyinput1), .B1(keyinput10), .B2(n15129), 
        .ZN(n15128) );
  OAI221_X1 U16669 ( .B1(n15130), .B2(keyinput1), .C1(n15129), .C2(keyinput10), 
        .A(n15128), .ZN(n15135) );
  INV_X1 U16670 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n15132) );
  AOI22_X1 U16671 ( .A1(n15133), .A2(keyinput23), .B1(n15132), .B2(keyinput5), 
        .ZN(n15131) );
  OAI221_X1 U16672 ( .B1(n15133), .B2(keyinput23), .C1(n15132), .C2(keyinput5), 
        .A(n15131), .ZN(n15134) );
  NOR3_X1 U16673 ( .A1(n15136), .A2(n15135), .A3(n15134), .ZN(n15169) );
  INV_X1 U16674 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n15139) );
  INV_X1 U16675 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n15138) );
  AOI22_X1 U16676 ( .A1(n15139), .A2(keyinput3), .B1(keyinput33), .B2(n15138), 
        .ZN(n15137) );
  OAI221_X1 U16677 ( .B1(n15139), .B2(keyinput3), .C1(n15138), .C2(keyinput33), 
        .A(n15137), .ZN(n15140) );
  INV_X1 U16678 ( .A(n15140), .ZN(n15153) );
  AOI22_X1 U16679 ( .A1(n15143), .A2(keyinput38), .B1(n15142), .B2(keyinput2), 
        .ZN(n15141) );
  OAI221_X1 U16680 ( .B1(n15143), .B2(keyinput38), .C1(n15142), .C2(keyinput2), 
        .A(n15141), .ZN(n15144) );
  INV_X1 U16681 ( .A(n15144), .ZN(n15152) );
  XNOR2_X1 U16682 ( .A(P3_IR_REG_16__SCAN_IN), .B(keyinput20), .ZN(n15147) );
  XNOR2_X1 U16683 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput35), .ZN(n15146) );
  XNOR2_X1 U16684 ( .A(keyinput15), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n15145) );
  AND3_X1 U16685 ( .A1(n15147), .A2(n15146), .A3(n15145), .ZN(n15151) );
  INV_X1 U16686 ( .A(keyinput34), .ZN(n15148) );
  XNOR2_X1 U16687 ( .A(n15149), .B(n15148), .ZN(n15150) );
  AND4_X1 U16688 ( .A1(n15153), .A2(n15152), .A3(n15151), .A4(n15150), .ZN(
        n15168) );
  INV_X1 U16689 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n15156) );
  AOI22_X1 U16690 ( .A1(n15156), .A2(keyinput50), .B1(keyinput8), .B2(n15155), 
        .ZN(n15154) );
  OAI221_X1 U16691 ( .B1(n15156), .B2(keyinput50), .C1(n15155), .C2(keyinput8), 
        .A(n15154), .ZN(n15166) );
  AOI22_X1 U16692 ( .A1(n15159), .A2(keyinput58), .B1(keyinput62), .B2(n15158), 
        .ZN(n15157) );
  OAI221_X1 U16693 ( .B1(n15159), .B2(keyinput58), .C1(n15158), .C2(keyinput62), .A(n15157), .ZN(n15165) );
  XOR2_X1 U16694 ( .A(n12784), .B(keyinput31), .Z(n15163) );
  XNOR2_X1 U16695 ( .A(P1_REG2_REG_0__SCAN_IN), .B(keyinput18), .ZN(n15162) );
  XNOR2_X1 U16696 ( .A(P2_REG0_REG_14__SCAN_IN), .B(keyinput42), .ZN(n15161)
         );
  XNOR2_X1 U16697 ( .A(P3_IR_REG_20__SCAN_IN), .B(keyinput61), .ZN(n15160) );
  NAND4_X1 U16698 ( .A1(n15163), .A2(n15162), .A3(n15161), .A4(n15160), .ZN(
        n15164) );
  NOR3_X1 U16699 ( .A1(n15166), .A2(n15165), .A3(n15164), .ZN(n15167) );
  NAND4_X1 U16700 ( .A1(n15170), .A2(n15169), .A3(n15168), .A4(n15167), .ZN(
        n15234) );
  AOI22_X1 U16701 ( .A1(n15173), .A2(keyinput55), .B1(keyinput26), .B2(n15172), 
        .ZN(n15171) );
  OAI221_X1 U16702 ( .B1(n15173), .B2(keyinput55), .C1(n15172), .C2(keyinput26), .A(n15171), .ZN(n15184) );
  INV_X1 U16703 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n15176) );
  AOI22_X1 U16704 ( .A1(n15176), .A2(keyinput46), .B1(n15175), .B2(keyinput29), 
        .ZN(n15174) );
  OAI221_X1 U16705 ( .B1(n15176), .B2(keyinput46), .C1(n15175), .C2(keyinput29), .A(n15174), .ZN(n15183) );
  XOR2_X1 U16706 ( .A(n15177), .B(keyinput0), .Z(n15181) );
  XNOR2_X1 U16707 ( .A(keyinput27), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n15180) );
  XNOR2_X1 U16708 ( .A(P3_REG2_REG_1__SCAN_IN), .B(keyinput53), .ZN(n15179) );
  XNOR2_X1 U16709 ( .A(P3_IR_REG_21__SCAN_IN), .B(keyinput32), .ZN(n15178) );
  NAND4_X1 U16710 ( .A1(n15181), .A2(n15180), .A3(n15179), .A4(n15178), .ZN(
        n15182) );
  NOR3_X1 U16711 ( .A1(n15184), .A2(n15183), .A3(n15182), .ZN(n15232) );
  AOI22_X1 U16712 ( .A1(n15187), .A2(keyinput40), .B1(keyinput16), .B2(n15186), 
        .ZN(n15185) );
  OAI221_X1 U16713 ( .B1(n15187), .B2(keyinput40), .C1(n15186), .C2(keyinput16), .A(n15185), .ZN(n15199) );
  AOI22_X1 U16714 ( .A1(n15190), .A2(keyinput39), .B1(keyinput49), .B2(n15189), 
        .ZN(n15188) );
  OAI221_X1 U16715 ( .B1(n15190), .B2(keyinput39), .C1(n15189), .C2(keyinput49), .A(n15188), .ZN(n15198) );
  AOI22_X1 U16716 ( .A1(n15193), .A2(keyinput43), .B1(n15192), .B2(keyinput7), 
        .ZN(n15191) );
  OAI221_X1 U16717 ( .B1(n15193), .B2(keyinput43), .C1(n15192), .C2(keyinput7), 
        .A(n15191), .ZN(n15197) );
  XOR2_X1 U16718 ( .A(n12044), .B(keyinput44), .Z(n15195) );
  XNOR2_X1 U16719 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput25), .ZN(n15194) );
  NAND2_X1 U16720 ( .A1(n15195), .A2(n15194), .ZN(n15196) );
  NOR4_X1 U16721 ( .A1(n15199), .A2(n15198), .A3(n15197), .A4(n15196), .ZN(
        n15231) );
  AOI22_X1 U16722 ( .A1(n15202), .A2(keyinput45), .B1(keyinput57), .B2(n15201), 
        .ZN(n15200) );
  OAI221_X1 U16723 ( .B1(n15202), .B2(keyinput45), .C1(n15201), .C2(keyinput57), .A(n15200), .ZN(n15213) );
  AOI22_X1 U16724 ( .A1(n15204), .A2(keyinput59), .B1(n13268), .B2(keyinput4), 
        .ZN(n15203) );
  OAI221_X1 U16725 ( .B1(n15204), .B2(keyinput59), .C1(n13268), .C2(keyinput4), 
        .A(n15203), .ZN(n15212) );
  AOI22_X1 U16726 ( .A1(n15207), .A2(keyinput41), .B1(keyinput36), .B2(n15206), 
        .ZN(n15205) );
  OAI221_X1 U16727 ( .B1(n15207), .B2(keyinput41), .C1(n15206), .C2(keyinput36), .A(n15205), .ZN(n15211) );
  XNOR2_X1 U16728 ( .A(P2_REG1_REG_14__SCAN_IN), .B(keyinput48), .ZN(n15209)
         );
  XNOR2_X1 U16729 ( .A(P1_REG3_REG_7__SCAN_IN), .B(keyinput14), .ZN(n15208) );
  NAND2_X1 U16730 ( .A1(n15209), .A2(n15208), .ZN(n15210) );
  NOR4_X1 U16731 ( .A1(n15213), .A2(n15212), .A3(n15211), .A4(n15210), .ZN(
        n15230) );
  AOI22_X1 U16732 ( .A1(n15216), .A2(keyinput19), .B1(n15215), .B2(keyinput47), 
        .ZN(n15214) );
  OAI221_X1 U16733 ( .B1(n15216), .B2(keyinput19), .C1(n15215), .C2(keyinput47), .A(n15214), .ZN(n15228) );
  INV_X1 U16734 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n15219) );
  AOI22_X1 U16735 ( .A1(n15219), .A2(keyinput63), .B1(keyinput56), .B2(n15218), 
        .ZN(n15217) );
  OAI221_X1 U16736 ( .B1(n15219), .B2(keyinput63), .C1(n15218), .C2(keyinput56), .A(n15217), .ZN(n15227) );
  AOI22_X1 U16737 ( .A1(n15222), .A2(keyinput13), .B1(keyinput52), .B2(n15221), 
        .ZN(n15220) );
  OAI221_X1 U16738 ( .B1(n15222), .B2(keyinput13), .C1(n15221), .C2(keyinput52), .A(n15220), .ZN(n15226) );
  XNOR2_X1 U16739 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput54), .ZN(n15224)
         );
  XNOR2_X1 U16740 ( .A(SI_19_), .B(keyinput24), .ZN(n15223) );
  NAND2_X1 U16741 ( .A1(n15224), .A2(n15223), .ZN(n15225) );
  NOR4_X1 U16742 ( .A1(n15228), .A2(n15227), .A3(n15226), .A4(n15225), .ZN(
        n15229) );
  NAND4_X1 U16743 ( .A1(n15232), .A2(n15231), .A3(n15230), .A4(n15229), .ZN(
        n15233) );
  NOR2_X1 U16744 ( .A1(n15234), .A2(n15233), .ZN(n15235) );
  XOR2_X1 U16745 ( .A(n15236), .B(n15235), .Z(n15237) );
  XNOR2_X1 U16746 ( .A(n15238), .B(n15237), .ZN(P2_U3262) );
  XOR2_X1 U16747 ( .A(n15240), .B(n15239), .Z(SUB_1596_U59) );
  XNOR2_X1 U16748 ( .A(n15241), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16749 ( .B1(n15242), .B2(n9531), .A(n15250), .ZN(SUB_1596_U53) );
  XOR2_X1 U16750 ( .A(n15244), .B(n15243), .Z(SUB_1596_U56) );
  OAI21_X1 U16751 ( .B1(n15247), .B2(n15246), .A(n15245), .ZN(n15248) );
  XNOR2_X1 U16752 ( .A(n15248), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U16753 ( .A(n15250), .B(n15249), .Z(SUB_1596_U5) );
  CLKBUF_X1 U7202 ( .A(n11422), .Z(n11609) );
  CLKBUF_X1 U7208 ( .A(n12791), .Z(n6639) );
  CLKBUF_X1 U7224 ( .A(n12043), .Z(n6441) );
  INV_X1 U7249 ( .A(n12049), .ZN(n8093) );
  NAND2_X1 U7251 ( .A1(n10453), .A2(n7764), .ZN(n10501) );
  CLKBUF_X1 U7265 ( .A(n7627), .Z(n7476) );
  CLKBUF_X1 U7266 ( .A(n9734), .Z(n11657) );
  XNOR2_X1 U7789 ( .A(n7642), .B(n7641), .ZN(n11324) );
endmodule

