

module b22_C_gen_AntiSAT_k_128_2 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225;

  OAI21_X1 U7216 ( .B1(n11768), .B2(n11757), .A(n14779), .ZN(n13244) );
  INV_X2 U7217 ( .A(n11850), .ZN(n13412) );
  AND2_X1 U7218 ( .A1(n10194), .A2(n10079), .ZN(n10148) );
  BUF_X1 U7219 ( .A(n10204), .Z(n6487) );
  NAND2_X1 U7221 ( .A1(n10561), .A2(n11228), .ZN(n10760) );
  CLKBUF_X1 U7222 ( .A(n8214), .Z(n10076) );
  INV_X1 U7223 ( .A(n8068), .ZN(n7592) );
  NAND2_X1 U7224 ( .A1(n9132), .A2(n7191), .ZN(n10490) );
  BUF_X1 U7225 ( .A(n9136), .Z(n9569) );
  NAND2_X1 U7226 ( .A1(n9091), .A2(n9099), .ZN(n11165) );
  XNOR2_X1 U7227 ( .A(n14034), .B(n14141), .ZN(n14015) );
  OR2_X2 U7228 ( .A1(n9467), .A2(n9466), .ZN(n7418) );
  INV_X2 U7229 ( .A(n12107), .ZN(n12146) );
  INV_X1 U7230 ( .A(n8663), .ZN(n12182) );
  BUF_X1 U7231 ( .A(n10204), .Z(n6488) );
  INV_X1 U7232 ( .A(n9819), .ZN(n7943) );
  AND2_X1 U7233 ( .A1(n13270), .A2(n12015), .ZN(n13470) );
  MUX2_X1 U7234 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7471), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n7472) );
  INV_X1 U7235 ( .A(n12105), .ZN(n12147) );
  INV_X1 U7236 ( .A(n8420), .ZN(n8887) );
  INV_X1 U7237 ( .A(n8463), .ZN(n12181) );
  INV_X1 U7238 ( .A(n6469), .ZN(n6474) );
  INV_X1 U7239 ( .A(n13753), .ZN(n14543) );
  INV_X2 U7240 ( .A(n10760), .ZN(n11850) );
  CLKBUF_X3 U7241 ( .A(n10065), .Z(n6477) );
  INV_X1 U7242 ( .A(n10875), .ZN(n12520) );
  AOI211_X1 U7243 ( .C1(n12629), .C2(n14964), .A(n12628), .B(n12627), .ZN(
        n12630) );
  AND2_X1 U7244 ( .A1(n6769), .A2(n6532), .ZN(n14355) );
  INV_X1 U7245 ( .A(n12813), .ZN(n12891) );
  INV_X2 U7246 ( .A(n12541), .ZN(n12601) );
  INV_X1 U7247 ( .A(n14586), .ZN(n10220) );
  AND4_X1 U7248 ( .A1(n6844), .A2(n6843), .A3(n8279), .A4(n8270), .ZN(n6468)
         );
  NAND2_X1 U7249 ( .A1(n7454), .A2(n7456), .ZN(n6469) );
  OR2_X1 U7250 ( .A1(n7798), .A2(n7797), .ZN(n6470) );
  NAND2_X2 U7251 ( .A1(n10067), .A2(n10332), .ZN(n7516) );
  NAND4_X2 U7252 ( .A1(n7521), .A2(n7524), .A3(n7522), .A4(n7523), .ZN(n10068)
         );
  NAND2_X2 U7253 ( .A1(n13728), .A2(n13727), .ZN(n13726) );
  NAND2_X2 U7254 ( .A1(n13057), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8384) );
  CLKBUF_X2 U7255 ( .A(n10071), .Z(n6471) );
  XNOR2_X2 U7256 ( .A(n14202), .B(n14201), .ZN(n14239) );
  NAND2_X2 U7257 ( .A1(n14199), .A2(n14200), .ZN(n14202) );
  NAND3_X2 U7258 ( .A1(n8394), .A2(n8393), .A3(n6718), .ZN(n12523) );
  XNOR2_X1 U7259 ( .A(n13202), .B(n10078), .ZN(n10071) );
  NAND4_X2 U7260 ( .A1(n7505), .A2(n7504), .A3(n7503), .A4(n7502), .ZN(n13202)
         );
  NOR2_X2 U7261 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n8416) );
  CLKBUF_X3 U7262 ( .A(n9584), .Z(n6472) );
  NAND2_X1 U7263 ( .A1(n6638), .A2(n9102), .ZN(n9584) );
  AOI21_X2 U7264 ( .B1(n12397), .B2(n12396), .A(n8972), .ZN(n12490) );
  NAND2_X2 U7265 ( .A1(n7261), .A2(n6550), .ZN(n12397) );
  OAI21_X2 U7266 ( .B1(n14029), .B2(n11898), .A(n11897), .ZN(n14016) );
  AOI21_X2 U7267 ( .B1(n12062), .B2(n14152), .A(n11896), .ZN(n14029) );
  AOI21_X2 U7268 ( .B1(n13976), .B2(n11902), .A(n6554), .ZN(n13952) );
  NAND2_X2 U7269 ( .A1(n13979), .A2(n6805), .ZN(n13976) );
  NOR2_X2 U7270 ( .A1(n11835), .A2(n11834), .ZN(n11925) );
  XNOR2_X2 U7271 ( .A(n14197), .B(n6691), .ZN(n14252) );
  NAND2_X2 U7272 ( .A1(n14195), .A2(n6692), .ZN(n14197) );
  BUF_X2 U7273 ( .A(n8187), .Z(n6473) );
  NAND2_X1 U7274 ( .A1(n7456), .A2(n13582), .ZN(n8187) );
  OAI21_X2 U7275 ( .B1(n11539), .B2(n8543), .A(n11538), .ZN(n12528) );
  AOI21_X2 U7276 ( .B1(n7108), .B2(n6828), .A(n6509), .ZN(n6827) );
  OAI21_X4 U7277 ( .B1(n10067), .B2(n10066), .A(n13257), .ZN(n10179) );
  NOR2_X2 U7278 ( .A1(n10178), .A2(n6476), .ZN(n10067) );
  XNOR2_X1 U7280 ( .A(n6871), .B(n8362), .ZN(n12610) );
  OAI21_X2 U7281 ( .B1(n8096), .B2(n8095), .A(n8094), .ZN(n8119) );
  NOR2_X2 U7282 ( .A1(n14283), .A2(n14284), .ZN(n14288) );
  INV_X2 U7283 ( .A(n6469), .ZN(n6475) );
  NAND2_X4 U7284 ( .A1(n12370), .A2(n11867), .ZN(n8890) );
  OAI222_X1 U7285 ( .A1(P3_U3151), .A2(n12370), .B1(n13067), .B2(n12372), .C1(
        n15145), .C2(n13059), .ZN(P3_U3265) );
  AND2_X4 U7286 ( .A1(n8388), .A2(n12370), .ZN(n12172) );
  XNOR2_X2 U7287 ( .A(n8384), .B(n13058), .ZN(n12370) );
  CLKBUF_X1 U7288 ( .A(n10065), .Z(n6476) );
  XNOR2_X1 U7289 ( .A(n7487), .B(P2_IR_REG_22__SCAN_IN), .ZN(n10065) );
  XNOR2_X1 U7290 ( .A(n10347), .B(n10360), .ZN(n10404) );
  XNOR2_X2 U7291 ( .A(n8406), .B(n8405), .ZN(n10360) );
  XNOR2_X2 U7292 ( .A(n9077), .B(n14174), .ZN(n9080) );
  NAND2_X2 U7293 ( .A1(n14173), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9077) );
  OAI22_X2 U7294 ( .A1(n14869), .A2(n15011), .B1(n11393), .B2(n11411), .ZN(
        n14888) );
  NAND2_X4 U7295 ( .A1(n8389), .A2(n11867), .ZN(n8420) );
  XNOR2_X2 U7296 ( .A(n8387), .B(n8386), .ZN(n11867) );
  XOR2_X2 U7297 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n14255), .Z(n14256) );
  XNOR2_X2 U7298 ( .A(n14204), .B(n6961), .ZN(n14255) );
  INV_X1 U7299 ( .A(n7530), .ZN(n6478) );
  NAND2_X2 U7300 ( .A1(n7468), .A2(n7467), .ZN(n7510) );
  NOR2_X1 U7301 ( .A1(n11340), .A2(n7019), .ZN(n7018) );
  AND2_X1 U7302 ( .A1(n11278), .A2(n8789), .ZN(n8791) );
  NAND2_X1 U7303 ( .A1(n7684), .A2(n7683), .ZN(n10790) );
  NAND2_X1 U7304 ( .A1(n14795), .A2(n10115), .ZN(n13385) );
  CLKBUF_X2 U7305 ( .A(P2_U3947), .Z(n6480) );
  OAI211_X1 U7306 ( .C1(SI_9_), .C2(n8663), .A(n8508), .B(n8507), .ZN(n12270)
         );
  INV_X4 U7307 ( .A(n10798), .ZN(n12379) );
  INV_X1 U7308 ( .A(n13459), .ZN(n7048) );
  CLKBUF_X2 U7309 ( .A(n6481), .Z(n8111) );
  INV_X1 U7310 ( .A(n10197), .ZN(n10204) );
  INV_X1 U7311 ( .A(n13752), .ZN(n13711) );
  INV_X4 U7312 ( .A(n12106), .ZN(n10630) );
  BUF_X1 U7313 ( .A(n8776), .Z(n6484) );
  INV_X4 U7314 ( .A(n12172), .ZN(n8779) );
  BUF_X1 U7315 ( .A(n8776), .Z(n6485) );
  INV_X2 U7316 ( .A(n9579), .ZN(n9148) );
  NAND2_X1 U7317 ( .A1(n8389), .A2(n8388), .ZN(n8776) );
  INV_X4 U7318 ( .A(n7556), .ZN(n8210) );
  INV_X4 U7319 ( .A(n9133), .ZN(n9579) );
  INV_X4 U7320 ( .A(n8187), .ZN(n6479) );
  INV_X2 U7321 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X2 U7322 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8357) );
  OR2_X1 U7323 ( .A1(n8265), .A2(n8264), .ZN(n7283) );
  NOR2_X1 U7324 ( .A1(n13484), .A2(n6669), .ZN(n6668) );
  AOI21_X1 U7325 ( .B1(n13281), .B2(n13280), .A(n13279), .ZN(n13477) );
  AOI21_X1 U7326 ( .B1(n8896), .B2(n12878), .A(n8895), .ZN(n12378) );
  AOI22_X1 U7327 ( .A1(n13847), .A2(n14549), .B1(n14033), .B2(n13872), .ZN(
        n14075) );
  NOR2_X1 U7328 ( .A1(n13294), .A2(n7010), .ZN(n13277) );
  OAI21_X1 U7329 ( .B1(n6569), .B2(n7371), .A(n7372), .ZN(n7960) );
  NAND2_X1 U7330 ( .A1(n13319), .A2(n13318), .ZN(n13317) );
  INV_X1 U7331 ( .A(n7105), .ZN(n13163) );
  AOI21_X1 U7332 ( .B1(n9047), .B2(n9046), .A(n12499), .ZN(n9048) );
  NAND2_X1 U7333 ( .A1(n13347), .A2(n6529), .ZN(n13325) );
  NAND2_X1 U7334 ( .A1(n6786), .A2(n6785), .ZN(n13629) );
  OR2_X1 U7335 ( .A1(n13345), .A2(n13344), .ZN(n13347) );
  NAND2_X1 U7336 ( .A1(n13124), .A2(n11951), .ZN(n13106) );
  AND2_X1 U7337 ( .A1(n6953), .A2(n6952), .ZN(n6894) );
  AND2_X1 U7338 ( .A1(n13510), .A2(n12004), .ZN(n13367) );
  AOI21_X1 U7339 ( .B1(n6869), .B2(n12649), .A(n6867), .ZN(n6866) );
  AOI21_X1 U7340 ( .B1(n11906), .B2(n7189), .A(n7188), .ZN(n7187) );
  NAND2_X1 U7341 ( .A1(n12695), .A2(n8726), .ZN(n12697) );
  AND2_X1 U7342 ( .A1(n13845), .A2(n9599), .ZN(n11906) );
  NAND2_X1 U7343 ( .A1(n13669), .A2(n13668), .ZN(n13667) );
  AND2_X1 U7344 ( .A1(n7217), .A2(n6581), .ZN(n7216) );
  OR3_X1 U7345 ( .A1(n13854), .A2(n11908), .A3(n14058), .ZN(n14077) );
  NAND2_X1 U7346 ( .A1(n8162), .A2(n8161), .ZN(n13475) );
  NAND2_X1 U7347 ( .A1(n11982), .A2(n11981), .ZN(n13407) );
  NAND2_X1 U7348 ( .A1(n8750), .A2(n8749), .ZN(n12339) );
  NAND2_X1 U7349 ( .A1(n6960), .A2(n6959), .ZN(n14475) );
  NAND2_X1 U7350 ( .A1(n9536), .A2(n9535), .ZN(n14084) );
  NAND2_X1 U7351 ( .A1(n9522), .A2(n9521), .ZN(n14089) );
  NAND2_X1 U7352 ( .A1(n9504), .A2(n9503), .ZN(n14095) );
  XNOR2_X1 U7353 ( .A(n11923), .B(n11924), .ZN(n11835) );
  NAND2_X1 U7354 ( .A1(n12433), .A2(n8976), .ZN(n12466) );
  OAI21_X1 U7355 ( .B1(n8698), .B2(n8697), .A(n8333), .ZN(n8708) );
  OR2_X1 U7356 ( .A1(n6523), .A2(n12771), .ZN(n12755) );
  NAND2_X1 U7357 ( .A1(n7977), .A2(n7976), .ZN(n13523) );
  NAND2_X1 U7358 ( .A1(n8678), .A2(n8677), .ZN(n12954) );
  NAND2_X1 U7359 ( .A1(n11800), .A2(n11799), .ZN(n14427) );
  INV_X1 U7360 ( .A(n11742), .ZN(n11743) );
  OAI21_X1 U7361 ( .B1(n10915), .B2(n6808), .A(n6806), .ZN(n11362) );
  CLKBUF_X1 U7362 ( .A(n14377), .Z(n6677) );
  NAND2_X1 U7363 ( .A1(n8666), .A2(n8665), .ZN(n13034) );
  NAND2_X1 U7364 ( .A1(n13706), .A2(n11019), .ZN(n11024) );
  OAI21_X1 U7365 ( .B1(n10943), .B2(n10907), .A(n10909), .ZN(n10956) );
  AND2_X1 U7366 ( .A1(n11344), .A2(n7271), .ZN(n11586) );
  OR2_X1 U7367 ( .A1(n7629), .A2(n7399), .ZN(n7401) );
  NAND2_X1 U7368 ( .A1(n7807), .A2(n7806), .ZN(n14670) );
  NAND2_X1 U7369 ( .A1(n9273), .A2(n9272), .ZN(n11605) );
  NAND2_X1 U7370 ( .A1(n7734), .A2(n7733), .ZN(n11072) );
  AND2_X1 U7371 ( .A1(n8797), .A2(n11558), .ZN(n8798) );
  NAND2_X1 U7372 ( .A1(n7716), .A2(n7715), .ZN(n10887) );
  AND2_X1 U7373 ( .A1(n8679), .A2(n8668), .ZN(n12781) );
  NAND2_X1 U7374 ( .A1(n14760), .A2(n14759), .ZN(n14758) );
  XNOR2_X1 U7375 ( .A(n10635), .B(n10632), .ZN(n10672) );
  NOR2_X1 U7376 ( .A1(n10629), .A2(n7411), .ZN(n10635) );
  NAND2_X1 U7377 ( .A1(n7705), .A2(n7704), .ZN(n7760) );
  NAND2_X1 U7378 ( .A1(n9240), .A2(n9239), .ZN(n11200) );
  AND2_X2 U7379 ( .A1(n10139), .A2(n10336), .ZN(n14835) );
  INV_X1 U7380 ( .A(n10685), .ZN(n10692) );
  NAND2_X2 U7381 ( .A1(n7639), .A2(n7638), .ZN(n14815) );
  NAND2_X1 U7382 ( .A1(n6957), .A2(n6956), .ZN(n10602) );
  NAND2_X1 U7383 ( .A1(n7618), .A2(n7617), .ZN(n14808) );
  NAND2_X2 U7384 ( .A1(n9169), .A2(n9168), .ZN(n10674) );
  NAND2_X2 U7385 ( .A1(n7590), .A2(n7589), .ZN(n14802) );
  NAND2_X1 U7386 ( .A1(n6970), .A2(n14263), .ZN(n14264) );
  AND2_X1 U7387 ( .A1(n7659), .A2(n7636), .ZN(n9742) );
  NAND2_X2 U7388 ( .A1(n10476), .A2(n14526), .ZN(n14576) );
  NAND2_X1 U7389 ( .A1(n7635), .A2(n7634), .ZN(n7659) );
  NOR2_X1 U7390 ( .A1(n14258), .A2(n14259), .ZN(n14260) );
  NAND2_X1 U7391 ( .A1(n7561), .A2(n7560), .ZN(n10843) );
  NAND2_X1 U7392 ( .A1(n7537), .A2(n6954), .ZN(n13459) );
  NAND2_X1 U7393 ( .A1(n9160), .A2(n9159), .ZN(n14554) );
  INV_X1 U7394 ( .A(n11101), .ZN(n12515) );
  XNOR2_X1 U7395 ( .A(n11395), .B(n11422), .ZN(n14906) );
  INV_X2 U7396 ( .A(n7591), .ZN(n6481) );
  NAND4_X1 U7397 ( .A1(n7624), .A2(n7623), .A3(n7622), .A4(n7621), .ZN(n13199)
         );
  NAND3_X1 U7398 ( .A1(n9174), .A2(n9172), .A3(n6547), .ZN(n13753) );
  NAND2_X1 U7399 ( .A1(n6689), .A2(n14254), .ZN(n14257) );
  INV_X2 U7400 ( .A(n9584), .ZN(n9143) );
  INV_X2 U7401 ( .A(n7592), .ZN(n8184) );
  AND4_X1 U7402 ( .A1(n9108), .A2(n9107), .A3(n9106), .A4(n9105), .ZN(n10014)
         );
  INV_X2 U7403 ( .A(n13738), .ZN(P1_U4016) );
  OR2_X1 U7404 ( .A1(n8515), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8529) );
  AND3_X1 U7405 ( .A1(n8398), .A2(n8397), .A3(n6717), .ZN(n12219) );
  INV_X2 U7406 ( .A(n9569), .ZN(n9575) );
  CLKBUF_X3 U7407 ( .A(n9137), .Z(n9567) );
  INV_X2 U7408 ( .A(n9111), .ZN(n9153) );
  AND2_X1 U7409 ( .A1(n7482), .A2(n7481), .ZN(n8214) );
  NAND2_X2 U7410 ( .A1(n10254), .A2(n9678), .ZN(n8663) );
  INV_X1 U7411 ( .A(n11867), .ZN(n8388) );
  NAND2_X2 U7412 ( .A1(n7455), .A2(n13582), .ZN(n8185) );
  NAND2_X1 U7413 ( .A1(n9587), .A2(n11168), .ZN(n6638) );
  NAND2_X1 U7414 ( .A1(n7455), .A2(n7454), .ZN(n8068) );
  OR3_X1 U7415 ( .A1(n11857), .A2(n11860), .A3(n14188), .ZN(n10323) );
  CLKBUF_X1 U7416 ( .A(n9130), .Z(n9580) );
  XNOR2_X1 U7417 ( .A(n9656), .B(n9655), .ZN(n11857) );
  NAND2_X1 U7418 ( .A1(n6490), .A2(n9678), .ZN(n9130) );
  NAND2_X1 U7419 ( .A1(n7486), .A2(n7485), .ZN(n11228) );
  INV_X1 U7420 ( .A(n10332), .ZN(n13257) );
  NAND2_X2 U7421 ( .A1(n13068), .A2(n12610), .ZN(n10254) );
  AND3_X1 U7422 ( .A1(n7483), .A2(n7498), .A3(n7497), .ZN(n10332) );
  NAND2_X1 U7423 ( .A1(n8361), .A2(n8385), .ZN(n13068) );
  NAND2_X1 U7424 ( .A1(n8385), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U7425 ( .A1(n7451), .A2(n7450), .ZN(n13582) );
  OAI21_X1 U7426 ( .B1(n9654), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9656) );
  AOI22_X1 U7427 ( .A1(n10443), .A2(P3_REG1_REG_3__SCAN_IN), .B1(n10442), .B2(
        n10441), .ZN(n11391) );
  NAND2_X1 U7428 ( .A1(n8266), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7487) );
  XNOR2_X1 U7429 ( .A(n10441), .B(n10437), .ZN(n10443) );
  XNOR2_X1 U7430 ( .A(n9101), .B(n9100), .ZN(n11168) );
  AOI21_X1 U7431 ( .B1(n14251), .B2(n14250), .A(n14308), .ZN(n15220) );
  XNOR2_X1 U7432 ( .A(n9097), .B(P1_IR_REG_21__SCAN_IN), .ZN(n10238) );
  NAND2_X1 U7433 ( .A1(n13577), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7453) );
  NAND2_X1 U7434 ( .A1(n6986), .A2(n6985), .ZN(n13577) );
  NOR2_X1 U7435 ( .A1(n7483), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n7484) );
  NAND2_X2 U7436 ( .A1(n9678), .A2(P2_U3088), .ZN(n13587) );
  XNOR2_X1 U7437 ( .A(n9079), .B(n9075), .ZN(n11865) );
  MUX2_X1 U7438 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9070), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n9071) );
  OR2_X1 U7439 ( .A1(n7782), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n7826) );
  AND2_X1 U7440 ( .A1(n8360), .A2(n8359), .ZN(n8383) );
  AND2_X1 U7441 ( .A1(n6934), .A2(n7275), .ZN(n8360) );
  OAI21_X1 U7442 ( .B1(n8842), .B2(n6936), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n6871) );
  NAND2_X1 U7443 ( .A1(n9067), .A2(n9066), .ZN(n9663) );
  OAI21_X1 U7444 ( .B1(n6804), .B2(n9094), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9095) );
  NOR2_X1 U7445 ( .A1(n6518), .A2(n6935), .ZN(n6934) );
  OAI21_X1 U7446 ( .B1(n6804), .B2(n7351), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9090) );
  INV_X1 U7447 ( .A(n6804), .ZN(n9092) );
  AND2_X1 U7448 ( .A1(n6696), .A2(n6695), .ZN(n7275) );
  NAND3_X1 U7449 ( .A1(n9351), .A2(n7206), .A3(n9058), .ZN(n6804) );
  INV_X1 U7450 ( .A(n9216), .ZN(n7206) );
  BUF_X4 U7451 ( .A(n10378), .Z(n6483) );
  AND2_X1 U7452 ( .A1(n9350), .A2(n9058), .ZN(n7203) );
  NOR2_X1 U7454 ( .A1(n9657), .A2(n9065), .ZN(n7205) );
  AND2_X1 U7455 ( .A1(n7410), .A2(n6526), .ZN(n7274) );
  AND4_X1 U7456 ( .A1(n9053), .A2(n9052), .A3(n9051), .A4(n9306), .ZN(n9350)
         );
  NAND2_X1 U7457 ( .A1(n7441), .A2(n7440), .ZN(n7442) );
  AND2_X1 U7458 ( .A1(n6975), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14245) );
  INV_X1 U7459 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13262) );
  NOR2_X1 U7460 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n9052) );
  NOR2_X1 U7461 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n7434) );
  NOR2_X1 U7462 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n9051) );
  INV_X1 U7463 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8581) );
  NOR2_X1 U7464 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n8347) );
  NOR2_X1 U7465 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n6838) );
  NOR2_X1 U7466 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n6917) );
  NOR2_X2 U7467 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n6915) );
  NOR2_X1 U7468 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8346) );
  NOR2_X1 U7469 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n7432) );
  NOR2_X1 U7470 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n9060) );
  NOR2_X1 U7471 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n7433) );
  INV_X1 U7472 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7461) );
  NOR2_X1 U7473 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7430) );
  INV_X1 U7474 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9388) );
  XNOR2_X1 U7475 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n14244) );
  INV_X1 U7476 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9306) );
  INV_X1 U7477 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8521) );
  INV_X1 U7478 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8763) );
  INV_X4 U7479 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7480 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8563) );
  INV_X1 U7481 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8270) );
  INV_X1 U7482 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9655) );
  NOR2_X1 U7483 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n9061) );
  NOR2_X1 U7484 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n9062) );
  NOR2_X1 U7485 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n7258) );
  AOI21_X1 U7486 ( .B1(n9436), .B2(n9437), .A(n6634), .ZN(n6686) );
  OR2_X2 U7487 ( .A1(n12551), .A2(n6760), .ZN(n6759) );
  NAND2_X1 U7488 ( .A1(n13885), .A2(n13886), .ZN(n13884) );
  OAI22_X1 U7489 ( .A1(n7729), .A2(n7379), .B1(n7728), .B2(n7727), .ZN(n7748)
         );
  OAI222_X1 U7490 ( .A1(n13587), .A2(n14182), .B1(P2_U3088), .B2(n7456), .C1(
        n12165), .C2(n13593), .ZN(P2_U3297) );
  OAI21_X2 U7491 ( .B1(n12007), .B2(n13487), .A(n13317), .ZN(n13295) );
  OR2_X2 U7492 ( .A1(n10804), .A2(n12521), .ZN(n6851) );
  OR2_X1 U7493 ( .A1(n8416), .A2(n8357), .ZN(n8417) );
  NOR2_X2 U7494 ( .A1(n11925), .A2(n6847), .ZN(n14383) );
  NOR2_X2 U7495 ( .A1(n14555), .A2(n10674), .ZN(n10466) );
  OAI21_X2 U7496 ( .B1(n14292), .B2(n14463), .A(n14460), .ZN(n14467) );
  XNOR2_X1 U7497 ( .A(n9095), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14189) );
  BUF_X4 U7498 ( .A(n10197), .Z(n11963) );
  NOR2_X2 U7499 ( .A1(n11781), .A2(n14388), .ZN(n11849) );
  INV_X1 U7500 ( .A(n7556), .ZN(n6486) );
  INV_X2 U7501 ( .A(n6481), .ZN(n8223) );
  INV_X2 U7502 ( .A(n6481), .ZN(n8222) );
  NAND2_X1 U7503 ( .A1(n9666), .A2(n9665), .ZN(n6489) );
  NAND2_X1 U7504 ( .A1(n9666), .A2(n9665), .ZN(n6490) );
  CLKBUF_X1 U7505 ( .A(n14048), .Z(n6491) );
  OAI21_X1 U7506 ( .B1(n9436), .B2(n9437), .A(n6563), .ZN(n6685) );
  INV_X2 U7507 ( .A(n10078), .ZN(n10194) );
  NAND3_X2 U7508 ( .A1(n7515), .A2(n7052), .A3(n7050), .ZN(n10078) );
  NOR2_X2 U7509 ( .A1(n10701), .A2(n14607), .ZN(n10936) );
  INV_X1 U7510 ( .A(n9111), .ZN(n6492) );
  NAND2_X1 U7511 ( .A1(n6489), .A2(n7530), .ZN(n9111) );
  NOR2_X1 U7512 ( .A1(n8808), .A2(n6858), .ZN(n6857) );
  INV_X1 U7513 ( .A(n8807), .ZN(n6858) );
  NAND2_X1 U7514 ( .A1(n7871), .A2(n15094), .ZN(n7894) );
  NAND2_X1 U7515 ( .A1(n7851), .A2(n15068), .ZN(n7869) );
  NOR2_X1 U7516 ( .A1(n8350), .A2(n8349), .ZN(n6695) );
  NOR2_X1 U7517 ( .A1(n13936), .A2(n7199), .ZN(n7198) );
  INV_X1 U7518 ( .A(n6484), .ZN(n8754) );
  NAND2_X1 U7519 ( .A1(n9819), .A2(n9678), .ZN(n7556) );
  OAI21_X1 U7520 ( .B1(n9147), .B2(n9146), .A(n9145), .ZN(n9162) );
  NAND2_X1 U7521 ( .A1(n6688), .A2(n6687), .ZN(n9274) );
  NAND2_X1 U7522 ( .A1(n9262), .A2(n9264), .ZN(n6687) );
  NAND2_X1 U7523 ( .A1(n7387), .A2(n7386), .ZN(n7385) );
  INV_X1 U7524 ( .A(n7865), .ZN(n7387) );
  INV_X1 U7525 ( .A(n7864), .ZN(n7386) );
  AOI21_X1 U7526 ( .B1(n6714), .B2(n6715), .A(n6546), .ZN(n6713) );
  INV_X1 U7527 ( .A(n6716), .ZN(n6715) );
  OAI21_X1 U7528 ( .B1(n6705), .B2(n12329), .A(n6702), .ZN(n7153) );
  INV_X1 U7529 ( .A(n6703), .ZN(n6702) );
  AOI21_X1 U7530 ( .B1(n12328), .B2(n6706), .A(n6606), .ZN(n6705) );
  OAI21_X1 U7531 ( .B1(n12331), .B2(n12332), .A(n6704), .ZN(n6703) );
  AND2_X1 U7532 ( .A1(n7362), .A2(n7369), .ZN(n7361) );
  INV_X1 U7533 ( .A(n8075), .ZN(n7369) );
  NAND2_X1 U7534 ( .A1(n8076), .A2(n7363), .ZN(n7362) );
  NOR2_X1 U7535 ( .A1(n8076), .A2(n7363), .ZN(n7360) );
  INV_X1 U7536 ( .A(n7921), .ZN(n7318) );
  INV_X1 U7537 ( .A(n7145), .ZN(n6734) );
  INV_X1 U7538 ( .A(n8035), .ZN(n6663) );
  NAND2_X1 U7539 ( .A1(n7896), .A2(n10088), .ZN(n7921) );
  INV_X1 U7540 ( .A(n7780), .ZN(n7298) );
  NOR2_X1 U7541 ( .A1(n13001), .A2(n12188), .ZN(n12352) );
  INV_X1 U7542 ( .A(n12370), .ZN(n8389) );
  NOR2_X1 U7543 ( .A1(n8818), .A2(n6863), .ZN(n6862) );
  INV_X1 U7544 ( .A(n8816), .ZN(n6863) );
  OR2_X1 U7545 ( .A1(n12748), .A2(n12759), .ZN(n12324) );
  NOR2_X1 U7546 ( .A1(n6907), .A2(n12333), .ZN(n6906) );
  INV_X1 U7547 ( .A(n12330), .ZN(n6907) );
  NAND2_X1 U7548 ( .A1(n12677), .A2(n8737), .ZN(n6905) );
  INV_X1 U7549 ( .A(n8879), .ZN(n8881) );
  INV_X1 U7550 ( .A(n8308), .ZN(n7148) );
  INV_X1 U7551 ( .A(n6740), .ZN(n6739) );
  OAI21_X1 U7552 ( .B1(n8450), .B2(n6741), .A(n8298), .ZN(n6740) );
  AND2_X1 U7553 ( .A1(n7137), .A2(n8299), .ZN(n7136) );
  INV_X1 U7554 ( .A(n8474), .ZN(n7137) );
  NOR2_X1 U7555 ( .A1(n13487), .A2(n13335), .ZN(n6949) );
  OAI21_X1 U7556 ( .B1(n11326), .B2(n7015), .A(n7013), .ZN(n11654) );
  INV_X1 U7557 ( .A(n12138), .ZN(n7336) );
  NAND2_X1 U7558 ( .A1(n10672), .A2(n10673), .ZN(n6778) );
  NAND2_X1 U7559 ( .A1(n7187), .A2(n7190), .ZN(n7185) );
  NOR2_X1 U7560 ( .A1(n14102), .A2(n14108), .ZN(n6945) );
  NAND2_X1 U7561 ( .A1(n9082), .A2(n11865), .ZN(n9137) );
  INV_X1 U7562 ( .A(n9080), .ZN(n9082) );
  NAND2_X1 U7563 ( .A1(n6647), .A2(n6621), .ZN(n8158) );
  INV_X1 U7564 ( .A(n8178), .ZN(n6647) );
  INV_X1 U7565 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9064) );
  NAND2_X1 U7566 ( .A1(n9066), .A2(n7357), .ZN(n7356) );
  INV_X1 U7567 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7357) );
  NAND2_X1 U7568 ( .A1(n7870), .A2(n7869), .ZN(n7893) );
  AND2_X1 U7569 ( .A1(n7894), .A2(n7873), .ZN(n7892) );
  NAND2_X1 U7570 ( .A1(n7290), .A2(n7289), .ZN(n7824) );
  AOI21_X1 U7571 ( .B1(n7292), .B2(n7294), .A(n6566), .ZN(n7289) );
  INV_X1 U7572 ( .A(n7532), .ZN(n7531) );
  NAND2_X1 U7573 ( .A1(n7529), .A2(SI_2_), .ZN(n7553) );
  NAND2_X1 U7574 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n6693), .ZN(n6692) );
  INV_X1 U7575 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6693) );
  OR2_X1 U7576 ( .A1(n8679), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8701) );
  OR2_X1 U7577 ( .A1(n13015), .A2(n12651), .ZN(n7414) );
  OR2_X1 U7578 ( .A1(n9001), .A2(n12679), .ZN(n8827) );
  NOR2_X1 U7579 ( .A1(n12852), .A2(n6853), .ZN(n6852) );
  INV_X1 U7580 ( .A(n6855), .ZN(n6853) );
  NAND2_X1 U7581 ( .A1(n11684), .A2(n8802), .ZN(n12902) );
  NAND2_X1 U7582 ( .A1(n8847), .A2(n8846), .ZN(n9759) );
  INV_X1 U7583 ( .A(n7274), .ZN(n6935) );
  NAND2_X1 U7584 ( .A1(n8838), .A2(n8355), .ZN(n8836) );
  AND2_X1 U7585 ( .A1(n8304), .A2(n8303), .ZN(n8488) );
  AND2_X1 U7586 ( .A1(n14373), .A2(n11830), .ZN(n7112) );
  NAND2_X1 U7587 ( .A1(n7097), .A2(n7098), .ZN(n6836) );
  AND2_X1 U7588 ( .A1(n10850), .A2(n7099), .ZN(n7098) );
  NAND2_X1 U7589 ( .A1(n7102), .A2(n7100), .ZN(n7099) );
  AND2_X1 U7590 ( .A1(n10076), .A2(n6477), .ZN(n10119) );
  XOR2_X1 U7591 ( .A(n13177), .B(n13304), .Z(n13299) );
  NOR2_X1 U7592 ( .A1(n12006), .A2(n7070), .ZN(n7069) );
  INV_X1 U7593 ( .A(n7073), .ZN(n7070) );
  OR2_X1 U7594 ( .A1(n13523), .A2(n11983), .ZN(n6992) );
  OR2_X1 U7595 ( .A1(n13406), .A2(n12000), .ZN(n12002) );
  NOR2_X1 U7596 ( .A1(n11179), .A2(n7061), .ZN(n7060) );
  INV_X1 U7597 ( .A(n11073), .ZN(n7061) );
  INV_X1 U7598 ( .A(n10185), .ZN(n7046) );
  NAND2_X1 U7599 ( .A1(n6471), .A2(n10070), .ZN(n10145) );
  NOR2_X1 U7600 ( .A1(n9712), .A2(n7530), .ZN(n7051) );
  NAND2_X1 U7601 ( .A1(n8146), .A2(n8145), .ZN(n13471) );
  NAND2_X1 U7602 ( .A1(n7994), .A2(n7993), .ZN(n13518) );
  INV_X1 U7603 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7447) );
  NAND2_X1 U7604 ( .A1(n13698), .A2(n13699), .ZN(n7344) );
  AND2_X1 U7605 ( .A1(n13596), .A2(n7335), .ZN(n7334) );
  OR2_X1 U7606 ( .A1(n13719), .A2(n7336), .ZN(n7335) );
  NAND2_X1 U7607 ( .A1(n13667), .A2(n7338), .ZN(n13619) );
  NOR2_X1 U7608 ( .A1(n13621), .A2(n7339), .ZN(n7338) );
  INV_X1 U7609 ( .A(n12100), .ZN(n7339) );
  INV_X1 U7610 ( .A(n7340), .ZN(n6790) );
  INV_X1 U7611 ( .A(n6626), .ZN(n6777) );
  OR2_X1 U7612 ( .A1(n7322), .A2(n10016), .ZN(n12105) );
  NAND2_X1 U7613 ( .A1(n10229), .A2(n10323), .ZN(n7322) );
  NAND2_X2 U7614 ( .A1(n10323), .A2(n10016), .ZN(n12106) );
  NAND2_X1 U7615 ( .A1(n9562), .A2(n9560), .ZN(n7122) );
  INV_X2 U7616 ( .A(n9441), .ZN(n9547) );
  INV_X1 U7617 ( .A(n14071), .ZN(n13855) );
  OR2_X1 U7618 ( .A1(n7224), .A2(n7222), .ZN(n7221) );
  INV_X1 U7619 ( .A(n7227), .ZN(n7222) );
  INV_X1 U7620 ( .A(n7225), .ZN(n7224) );
  OAI21_X1 U7621 ( .B1(n13910), .B2(n7226), .A(n13883), .ZN(n7225) );
  OAI21_X1 U7622 ( .B1(n13911), .B2(n13910), .A(n6531), .ZN(n13885) );
  NAND2_X1 U7623 ( .A1(n14108), .A2(n13954), .ZN(n7233) );
  NOR2_X1 U7624 ( .A1(n13935), .A2(n7232), .ZN(n7231) );
  INV_X1 U7625 ( .A(n7235), .ZN(n7232) );
  NAND2_X2 U7626 ( .A1(n9666), .A2(n9665), .ZN(n9733) );
  AND2_X1 U7627 ( .A1(n14411), .A2(n13743), .ZN(n11715) );
  XNOR2_X1 U7628 ( .A(n14411), .B(n13743), .ZN(n11711) );
  NAND2_X1 U7629 ( .A1(n11370), .A2(n14443), .ZN(n11678) );
  NAND2_X1 U7630 ( .A1(n11816), .A2(n14421), .ZN(n11366) );
  INV_X2 U7631 ( .A(n9130), .ZN(n9415) );
  OAI21_X1 U7632 ( .B1(n9461), .B2(n8041), .A(n8040), .ZN(n8060) );
  XNOR2_X1 U7633 ( .A(n9650), .B(n9649), .ZN(n10322) );
  INV_X1 U7634 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9649) );
  AOI21_X1 U7635 ( .B1(n7760), .B2(n7759), .A(n6508), .ZN(n7781) );
  OAI21_X1 U7636 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14225), .A(n14224), .ZN(
        n14290) );
  NAND2_X1 U7637 ( .A1(n8878), .A2(n7413), .ZN(n8886) );
  INV_X1 U7638 ( .A(n14664), .ZN(n14384) );
  XNOR2_X1 U7639 ( .A(n12011), .B(n11990), .ZN(n13473) );
  AOI21_X1 U7640 ( .B1(n11995), .B2(n13437), .A(n11994), .ZN(n13472) );
  NAND2_X1 U7641 ( .A1(n11993), .A2(n11992), .ZN(n11994) );
  OAI211_X1 U7642 ( .C1(n13295), .C2(n7005), .A(n7003), .B(n7002), .ZN(n11995)
         );
  OR2_X1 U7643 ( .A1(n10337), .A2(n10333), .ZN(n7500) );
  MUX2_X1 U7644 ( .A(n9164), .B(n9163), .S(n14554), .Z(n9165) );
  OR2_X1 U7645 ( .A1(n9195), .A2(n7128), .ZN(n7127) );
  INV_X1 U7646 ( .A(n9194), .ZN(n7128) );
  OR2_X1 U7647 ( .A1(n7654), .A2(n7655), .ZN(n7656) );
  OAI21_X1 U7648 ( .B1(n7675), .B2(n7392), .A(n6655), .ZN(n7697) );
  AND2_X1 U7649 ( .A1(n7391), .A2(n6584), .ZN(n6655) );
  NOR2_X1 U7650 ( .A1(n9291), .A2(n9290), .ZN(n9312) );
  NOR2_X1 U7651 ( .A1(n6530), .A2(n7116), .ZN(n7115) );
  INV_X1 U7652 ( .A(n9413), .ZN(n7116) );
  NOR2_X1 U7653 ( .A1(n9400), .A2(n11898), .ZN(n7117) );
  INV_X1 U7654 ( .A(n11897), .ZN(n7118) );
  AOI21_X1 U7655 ( .B1(n6726), .B2(n12286), .A(n12285), .ZN(n6725) );
  OAI22_X1 U7656 ( .A1(n12283), .A2(n12901), .B1(n12346), .B2(n12282), .ZN(
        n6726) );
  INV_X1 U7657 ( .A(n9435), .ZN(n6634) );
  OAI21_X1 U7658 ( .B1(n7866), .B2(n7388), .A(n6656), .ZN(n7890) );
  AND2_X1 U7659 ( .A1(n6657), .A2(n7385), .ZN(n6656) );
  AOI21_X1 U7660 ( .B1(n12294), .B2(n12293), .A(n6722), .ZN(n12292) );
  AND2_X1 U7661 ( .A1(n12509), .A2(n13046), .ZN(n6722) );
  INV_X1 U7662 ( .A(n7936), .ZN(n7374) );
  INV_X1 U7663 ( .A(n7935), .ZN(n7373) );
  AOI21_X1 U7664 ( .B1(n6713), .B2(n6711), .A(n6578), .ZN(n6710) );
  INV_X1 U7665 ( .A(n6714), .ZN(n6711) );
  INV_X1 U7666 ( .A(n6713), .ZN(n6712) );
  NAND2_X1 U7667 ( .A1(n9494), .A2(n7125), .ZN(n7124) );
  NAND2_X1 U7668 ( .A1(n12338), .A2(n7153), .ZN(n7150) );
  NOR2_X1 U7669 ( .A1(n6507), .A2(n12312), .ZN(n7149) );
  NAND2_X1 U7670 ( .A1(n12335), .A2(n7153), .ZN(n7152) );
  INV_X1 U7671 ( .A(n7820), .ZN(n7821) );
  INV_X1 U7672 ( .A(n8266), .ZN(n7480) );
  NOR2_X1 U7673 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n7479) );
  INV_X1 U7674 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7441) );
  INV_X1 U7675 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7440) );
  NAND2_X1 U7676 ( .A1(n8063), .A2(n8062), .ZN(n8079) );
  NAND2_X1 U7677 ( .A1(n8060), .A2(n8059), .ZN(n8063) );
  AND2_X1 U7678 ( .A1(n7313), .A2(n6618), .ZN(n6885) );
  INV_X1 U7679 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9054) );
  INV_X1 U7680 ( .A(n7849), .ZN(n7299) );
  AOI21_X1 U7681 ( .B1(n7297), .B2(n7295), .A(n7293), .ZN(n7292) );
  INV_X1 U7682 ( .A(n7800), .ZN(n7293) );
  INV_X1 U7683 ( .A(n7295), .ZN(n7294) );
  OAI21_X1 U7684 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14217), .A(n14216), .ZN(
        n14218) );
  INV_X1 U7685 ( .A(n6851), .ZN(n8922) );
  INV_X1 U7686 ( .A(n12218), .ZN(n12367) );
  OR2_X1 U7687 ( .A1(n14958), .A2(n14957), .ZN(n7028) );
  OR3_X1 U7688 ( .A1(n8751), .A2(P3_REG3_REG_27__SCAN_IN), .A3(
        P3_REG3_REG_26__SCAN_IN), .ZN(n8752) );
  INV_X1 U7689 ( .A(n12698), .ZN(n12329) );
  NOR2_X1 U7690 ( .A1(n8673), .A2(n6933), .ZN(n6932) );
  INV_X1 U7691 ( .A(n12306), .ZN(n6933) );
  AOI21_X1 U7692 ( .B1(n6857), .B2(n12886), .A(n6611), .ZN(n6855) );
  NAND2_X1 U7693 ( .A1(n6922), .A2(n6923), .ZN(n6921) );
  INV_X1 U7694 ( .A(n6924), .ZN(n6922) );
  NOR2_X1 U7695 ( .A1(n12263), .A2(n8794), .ZN(n8795) );
  INV_X1 U7696 ( .A(n6913), .ZN(n6912) );
  OAI21_X1 U7697 ( .B1(n12240), .B2(n6914), .A(n12245), .ZN(n6913) );
  INV_X1 U7698 ( .A(n12242), .ZN(n6914) );
  NAND2_X1 U7699 ( .A1(n12970), .A2(n6932), .ZN(n6931) );
  NAND2_X1 U7700 ( .A1(n12809), .A2(n12808), .ZN(n12795) );
  NOR2_X1 U7701 ( .A1(n8341), .A2(n6752), .ZN(n6751) );
  INV_X1 U7702 ( .A(n8340), .ZN(n6752) );
  INV_X1 U7703 ( .A(n8339), .ZN(n6749) );
  NOR2_X1 U7704 ( .A1(n8761), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n8765) );
  OR2_X1 U7705 ( .A1(n8633), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n8761) );
  AND2_X1 U7706 ( .A1(n10432), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8314) );
  INV_X1 U7707 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8310) );
  INV_X1 U7708 ( .A(n13113), .ZN(n7096) );
  AOI21_X1 U7709 ( .B1(n7359), .B2(n6505), .A(n6575), .ZN(n7358) );
  INV_X1 U7710 ( .A(n13582), .ZN(n7454) );
  INV_X1 U7711 ( .A(n7456), .ZN(n7455) );
  OAI21_X1 U7712 ( .B1(n7010), .B2(n7008), .A(n6561), .ZN(n7007) );
  INV_X1 U7713 ( .A(n13299), .ZN(n7008) );
  OAI21_X1 U7714 ( .B1(n13475), .B2(n13176), .A(n12010), .ZN(n7012) );
  NOR2_X1 U7715 ( .A1(n6539), .A2(n6990), .ZN(n6989) );
  INV_X1 U7716 ( .A(n6992), .ZN(n6990) );
  INV_X1 U7717 ( .A(n7020), .ZN(n7019) );
  AND2_X1 U7718 ( .A1(n10576), .A2(n10657), .ZN(n6996) );
  AND2_X1 U7719 ( .A1(n13299), .A2(n6533), .ZN(n7067) );
  NOR2_X1 U7720 ( .A1(n7435), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n6839) );
  OR2_X1 U7721 ( .A1(n7681), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n7707) );
  INV_X1 U7722 ( .A(n12111), .ZN(n7343) );
  INV_X1 U7723 ( .A(n11889), .ZN(n7189) );
  INV_X1 U7724 ( .A(n13845), .ZN(n7188) );
  NAND2_X1 U7725 ( .A1(n13870), .A2(n11889), .ZN(n11890) );
  NAND2_X1 U7726 ( .A1(n14089), .A2(n13871), .ZN(n7227) );
  INV_X1 U7727 ( .A(n11715), .ZN(n7242) );
  AND2_X1 U7728 ( .A1(n11738), .A2(n9604), .ZN(n11736) );
  NOR2_X1 U7729 ( .A1(n11711), .A2(n7245), .ZN(n7244) );
  INV_X1 U7730 ( .A(n11672), .ZN(n7245) );
  OAI21_X1 U7731 ( .B1(n7406), .B2(n10490), .A(n10234), .ZN(n10223) );
  NAND2_X1 U7732 ( .A1(n9080), .A2(n11865), .ZN(n9136) );
  NOR2_X1 U7733 ( .A1(n14089), .A2(n6942), .ZN(n6941) );
  INV_X1 U7734 ( .A(n6943), .ZN(n6942) );
  NAND2_X1 U7735 ( .A1(n10906), .A2(n10905), .ZN(n10943) );
  INV_X1 U7736 ( .A(n7310), .ZN(n7309) );
  INV_X1 U7737 ( .A(n8143), .ZN(n7312) );
  NAND2_X1 U7738 ( .A1(n8158), .A2(n8123), .ZN(n8127) );
  NAND2_X1 U7739 ( .A1(n8121), .A2(n8120), .ZN(n8178) );
  OAI21_X1 U7740 ( .B1(n8119), .B2(n15171), .A(n8118), .ZN(n8121) );
  XNOR2_X1 U7741 ( .A(n8079), .B(SI_24_), .ZN(n8077) );
  NOR2_X1 U7742 ( .A1(n7353), .A2(n7351), .ZN(n7350) );
  INV_X1 U7743 ( .A(n9096), .ZN(n7353) );
  AND2_X1 U7744 ( .A1(n7921), .A2(n7898), .ZN(n7919) );
  NAND2_X1 U7745 ( .A1(n7895), .A2(n7894), .ZN(n7920) );
  INV_X1 U7746 ( .A(n6890), .ZN(n6889) );
  OAI21_X1 U7747 ( .B1(n7824), .B2(n7823), .A(n7822), .ZN(n6890) );
  AOI21_X1 U7748 ( .B1(n7677), .B2(n7288), .A(n7287), .ZN(n7286) );
  INV_X1 U7749 ( .A(n7658), .ZN(n7288) );
  INV_X1 U7750 ( .A(n7679), .ZN(n7287) );
  OAI21_X1 U7751 ( .B1(n9678), .B2(n9688), .A(n6676), .ZN(n7583) );
  NAND2_X1 U7752 ( .A1(n6478), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6676) );
  INV_X1 U7753 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14240) );
  INV_X1 U7754 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14209) );
  INV_X1 U7755 ( .A(n8992), .ZN(n7253) );
  NAND2_X1 U7756 ( .A1(n6681), .A2(n6680), .ZN(n8509) );
  INV_X1 U7757 ( .A(n8482), .ZN(n6681) );
  NOR2_X2 U7758 ( .A1(n8408), .A2(n8407), .ZN(n10804) );
  NAND2_X1 U7759 ( .A1(n12449), .A2(n12450), .ZN(n7270) );
  NAND2_X1 U7760 ( .A1(n12523), .A2(n12219), .ZN(n12227) );
  OAI21_X1 U7761 ( .B1(n8979), .B2(n8978), .A(n8977), .ZN(n12412) );
  AOI21_X1 U7762 ( .B1(n7268), .B2(n7266), .A(n7265), .ZN(n7264) );
  INV_X1 U7763 ( .A(n7268), .ZN(n7267) );
  INV_X1 U7764 ( .A(n8986), .ZN(n7265) );
  AND4_X1 U7765 ( .A1(n8449), .A2(n8448), .A3(n8447), .A4(n8446), .ZN(n8936)
         );
  XNOR2_X1 U7766 ( .A(n11406), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n10447) );
  NOR2_X1 U7767 ( .A1(n14874), .A2(n11382), .ZN(n11383) );
  NAND2_X1 U7768 ( .A1(n14925), .A2(n14924), .ZN(n14923) );
  OR2_X1 U7769 ( .A1(n14911), .A2(n6762), .ZN(n6761) );
  NOR2_X1 U7770 ( .A1(n11428), .A2(n11639), .ZN(n6762) );
  OR2_X1 U7771 ( .A1(n12572), .A2(n12573), .ZN(n7024) );
  INV_X1 U7772 ( .A(n6759), .ZN(n12571) );
  NAND2_X1 U7773 ( .A1(n7275), .A2(n6526), .ZN(n8633) );
  AND2_X1 U7774 ( .A1(n6767), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6763) );
  AOI21_X1 U7775 ( .B1(n6901), .B2(n6900), .A(n6507), .ZN(n6899) );
  INV_X1 U7776 ( .A(n6906), .ZN(n6900) );
  OR2_X1 U7777 ( .A1(n12334), .A2(n6507), .ZN(n12663) );
  NAND2_X1 U7778 ( .A1(n8380), .A2(n8379), .ZN(n8751) );
  INV_X1 U7779 ( .A(n8731), .ZN(n8380) );
  XNOR2_X1 U7780 ( .A(n12702), .B(n12408), .ZN(n12698) );
  NOR2_X1 U7781 ( .A1(n8822), .A2(n6861), .ZN(n6860) );
  AND2_X1 U7782 ( .A1(n12714), .A2(n12713), .ZN(n12729) );
  NAND2_X1 U7783 ( .A1(n8696), .A2(n12324), .ZN(n12712) );
  AND2_X1 U7784 ( .A1(n12763), .A2(n12755), .ZN(n8819) );
  NAND2_X1 U7785 ( .A1(n8817), .A2(n6862), .ZN(n12741) );
  AND4_X1 U7786 ( .A1(n8684), .A2(n8683), .A3(n8682), .A4(n8681), .ZN(n12774)
         );
  OR2_X1 U7787 ( .A1(n12967), .A2(n12775), .ZN(n12306) );
  OR2_X1 U7788 ( .A1(n12736), .A2(n12789), .ZN(n12787) );
  AND4_X1 U7789 ( .A1(n8593), .A2(n8592), .A3(n8591), .A4(n8590), .ZN(n12862)
         );
  OR2_X1 U7790 ( .A1(n12288), .A2(n12206), .ZN(n12866) );
  AND4_X1 U7791 ( .A1(n8549), .A2(n8548), .A3(n8547), .A4(n8546), .ZN(n12907)
         );
  AND4_X1 U7792 ( .A1(n8520), .A2(n8519), .A3(n8518), .A4(n8517), .ZN(n12905)
         );
  NAND2_X1 U7793 ( .A1(n8496), .A2(n12265), .ZN(n11565) );
  AND4_X1 U7794 ( .A1(n8460), .A2(n8459), .A3(n8458), .A4(n8457), .ZN(n11516)
         );
  NAND2_X1 U7795 ( .A1(n6679), .A2(n6678), .ZN(n8468) );
  INV_X1 U7796 ( .A(n8455), .ZN(n6679) );
  AND2_X1 U7797 ( .A1(n12249), .A2(n12248), .ZN(n12245) );
  NOR2_X1 U7798 ( .A1(n8454), .A2(n8453), .ZN(n11282) );
  NAND2_X1 U7799 ( .A1(n10820), .A2(n12241), .ZN(n11216) );
  AND4_X1 U7800 ( .A1(n8436), .A2(n8435), .A3(n8434), .A4(n8433), .ZN(n10825)
         );
  NAND2_X1 U7801 ( .A1(n10821), .A2(n12198), .ZN(n10820) );
  NAND2_X1 U7802 ( .A1(n8830), .A2(n12346), .ZN(n12906) );
  OR2_X1 U7803 ( .A1(n8890), .A2(n8409), .ZN(n8411) );
  INV_X1 U7804 ( .A(n12846), .ZN(n12908) );
  NAND2_X1 U7805 ( .A1(n8741), .A2(n8740), .ZN(n9001) );
  AND2_X1 U7806 ( .A1(n13055), .A2(n9672), .ZN(n10714) );
  AND2_X1 U7807 ( .A1(n8829), .A2(n12346), .ZN(n12846) );
  INV_X1 U7808 ( .A(n12878), .ZN(n12903) );
  OAI21_X1 U7809 ( .B1(n12162), .B2(n12161), .A(n12164), .ZN(n12180) );
  INV_X1 U7810 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8386) );
  OAI21_X1 U7811 ( .B1(n8748), .B2(n8342), .A(n8343), .ZN(n8879) );
  NAND2_X1 U7812 ( .A1(n8338), .A2(n7162), .ZN(n8728) );
  NOR2_X1 U7813 ( .A1(n8842), .A2(P3_IR_REG_24__SCAN_IN), .ZN(n8838) );
  NAND2_X1 U7814 ( .A1(n8337), .A2(n7163), .ZN(n7162) );
  OR2_X1 U7815 ( .A1(n8336), .A2(n11777), .ZN(n8338) );
  NAND2_X1 U7816 ( .A1(n8688), .A2(n8332), .ZN(n8698) );
  NAND2_X1 U7817 ( .A1(n8768), .A2(n8770), .ZN(n8833) );
  AND2_X1 U7818 ( .A1(n8765), .A2(n8762), .ZN(n8768) );
  INV_X1 U7819 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8762) );
  INV_X1 U7820 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8770) );
  NAND2_X1 U7821 ( .A1(n8686), .A2(n8685), .ZN(n8688) );
  OR2_X1 U7822 ( .A1(n8674), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8676) );
  NAND2_X1 U7823 ( .A1(n8646), .A2(n8645), .ZN(n8648) );
  NAND2_X1 U7824 ( .A1(n8616), .A2(n8319), .ZN(n8629) );
  INV_X1 U7825 ( .A(n8597), .ZN(n7160) );
  OR2_X1 U7826 ( .A1(n8579), .A2(n8314), .ZN(n7159) );
  AOI21_X1 U7827 ( .B1(n7146), .B2(n7148), .A(n6570), .ZN(n7145) );
  AND2_X1 U7828 ( .A1(n8308), .A2(n8307), .ZN(n8523) );
  NAND2_X1 U7829 ( .A1(n8524), .A2(n8523), .ZN(n8526) );
  NAND2_X1 U7830 ( .A1(n6736), .A2(n6735), .ZN(n8491) );
  AOI21_X1 U7831 ( .B1(n6497), .B2(n6741), .A(n7134), .ZN(n6735) );
  NAND2_X1 U7832 ( .A1(n6737), .A2(n6739), .ZN(n8300) );
  OR2_X1 U7833 ( .A1(n8451), .A2(n6741), .ZN(n6737) );
  NAND2_X1 U7834 ( .A1(n8300), .A2(n7136), .ZN(n8477) );
  NAND2_X1 U7835 ( .A1(n6728), .A2(n8292), .ZN(n8438) );
  INV_X1 U7836 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7277) );
  NAND2_X1 U7837 ( .A1(n8285), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U7838 ( .A1(n7829), .A2(n7828), .ZN(n14377) );
  NAND2_X1 U7839 ( .A1(n7096), .A2(n7095), .ZN(n7094) );
  INV_X1 U7840 ( .A(n13112), .ZN(n7095) );
  XNOR2_X1 U7841 ( .A(n14815), .B(n6487), .ZN(n10509) );
  OAI21_X2 U7842 ( .B1(n11829), .B2(n7111), .A(n7109), .ZN(n11923) );
  INV_X1 U7843 ( .A(n7112), .ZN(n7111) );
  AOI21_X1 U7844 ( .B1(n7112), .B2(n7110), .A(n6567), .ZN(n7109) );
  NOR2_X1 U7845 ( .A1(n8259), .A2(n10076), .ZN(n7281) );
  NAND2_X1 U7846 ( .A1(n7484), .A2(n7477), .ZN(n8266) );
  NAND2_X1 U7847 ( .A1(n6479), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7457) );
  NOR2_X1 U7848 ( .A1(n13475), .A2(n6947), .ZN(n6946) );
  INV_X1 U7849 ( .A(n6948), .ZN(n6947) );
  NAND2_X1 U7850 ( .A1(n13475), .A2(n13176), .ZN(n12010) );
  INV_X1 U7851 ( .A(n7004), .ZN(n7002) );
  AOI22_X1 U7852 ( .A1(n6891), .A2(n7006), .B1(n7007), .B2(n12012), .ZN(n7004)
         );
  NAND2_X1 U7853 ( .A1(n7010), .A2(n12012), .ZN(n6891) );
  NAND2_X1 U7854 ( .A1(n13356), .A2(n6949), .ZN(n13310) );
  NAND2_X1 U7855 ( .A1(n13356), .A2(n13491), .ZN(n13331) );
  NAND2_X1 U7856 ( .A1(n13496), .A2(n13180), .ZN(n7073) );
  NOR2_X1 U7857 ( .A1(n13340), .A2(n7072), .ZN(n7071) );
  INV_X1 U7858 ( .A(n12005), .ZN(n7072) );
  NAND2_X1 U7859 ( .A1(n11987), .A2(n11986), .ZN(n13363) );
  OR2_X1 U7860 ( .A1(n13447), .A2(n13448), .ZN(n13445) );
  NAND2_X1 U7861 ( .A1(n11975), .A2(n7001), .ZN(n7000) );
  INV_X1 U7862 ( .A(n11841), .ZN(n7001) );
  NAND2_X1 U7863 ( .A1(n11658), .A2(n11657), .ZN(n11842) );
  AND2_X1 U7864 ( .A1(n11656), .A2(n11647), .ZN(n7081) );
  NAND2_X1 U7865 ( .A1(n11646), .A2(n11645), .ZN(n11786) );
  NOR2_X1 U7866 ( .A1(n7831), .A2(n7830), .ZN(n7858) );
  NAND2_X1 U7867 ( .A1(n7055), .A2(n7053), .ZN(n11339) );
  AOI21_X1 U7868 ( .B1(n7057), .B2(n7059), .A(n7054), .ZN(n7053) );
  INV_X1 U7869 ( .A(n11297), .ZN(n7054) );
  NAND2_X1 U7870 ( .A1(n11071), .A2(n11070), .ZN(n11074) );
  AOI21_X1 U7871 ( .B1(n6980), .B2(n10723), .A(n6560), .ZN(n6978) );
  INV_X1 U7872 ( .A(n6980), .ZN(n6979) );
  AND2_X1 U7873 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7619) );
  NAND2_X1 U7874 ( .A1(n10166), .A2(n10165), .ZN(n10169) );
  INV_X1 U7875 ( .A(n13430), .ZN(n13437) );
  NOR2_X1 U7876 ( .A1(n13203), .A2(n10079), .ZN(n10070) );
  AND2_X1 U7877 ( .A1(n10332), .A2(n11228), .ZN(n10338) );
  AND2_X1 U7878 ( .A1(n7068), .A2(n6533), .ZN(n13300) );
  NAND2_X1 U7879 ( .A1(n7068), .A2(n7067), .ZN(n13479) );
  NAND2_X1 U7880 ( .A1(n7925), .A2(n7924), .ZN(n13532) );
  AND2_X1 U7881 ( .A1(n9823), .A2(n9818), .ZN(n10129) );
  INV_X1 U7882 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8279) );
  XNOR2_X1 U7883 ( .A(n8275), .B(P2_IR_REG_25__SCAN_IN), .ZN(n10044) );
  OR2_X1 U7884 ( .A1(n8273), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n8277) );
  NAND2_X1 U7885 ( .A1(n6662), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n6661) );
  NAND2_X1 U7886 ( .A1(n7483), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6662) );
  AOI21_X1 U7887 ( .B1(n7334), .B2(n7336), .A(n6577), .ZN(n7333) );
  NOR2_X1 U7888 ( .A1(n10016), .A2(n10015), .ZN(n12042) );
  NAND2_X1 U7889 ( .A1(n13726), .A2(n7325), .ZN(n13638) );
  INV_X1 U7890 ( .A(n7342), .ZN(n7341) );
  OAI21_X1 U7891 ( .B1(n13690), .B2(n7343), .A(n13603), .ZN(n7342) );
  NOR2_X1 U7892 ( .A1(n9959), .A2(n7321), .ZN(n9962) );
  NOR2_X1 U7893 ( .A1(n14047), .A2(n12105), .ZN(n7321) );
  NAND2_X1 U7894 ( .A1(n9958), .A2(n9957), .ZN(n9959) );
  NAND2_X1 U7895 ( .A1(n9960), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n9957) );
  NAND2_X1 U7896 ( .A1(n9961), .A2(n6802), .ZN(n10021) );
  INV_X1 U7897 ( .A(n6801), .ZN(n6802) );
  OAI21_X1 U7898 ( .B1(n12107), .B2(n10218), .A(n6803), .ZN(n6801) );
  INV_X1 U7899 ( .A(n12036), .ZN(n6784) );
  INV_X1 U7900 ( .A(n6783), .ZN(n6782) );
  OAI21_X1 U7901 ( .B1(n6519), .B2(n6784), .A(n13680), .ZN(n6783) );
  AND2_X1 U7902 ( .A1(n12061), .A2(n7326), .ZN(n7325) );
  INV_X1 U7903 ( .A(n13640), .ZN(n7326) );
  NAND2_X1 U7904 ( .A1(n13651), .A2(n6797), .ZN(n6796) );
  INV_X1 U7905 ( .A(n12070), .ZN(n6797) );
  NAND2_X1 U7906 ( .A1(n6776), .A2(n6774), .ZN(n13706) );
  AND2_X1 U7907 ( .A1(n13707), .A2(n6775), .ZN(n6774) );
  NAND2_X1 U7908 ( .A1(n6777), .A2(n11012), .ZN(n6775) );
  NAND2_X1 U7909 ( .A1(n9640), .A2(n9639), .ZN(n9641) );
  INV_X1 U7910 ( .A(n9631), .ZN(n9640) );
  INV_X1 U7911 ( .A(n9638), .ZN(n9639) );
  NAND2_X1 U7912 ( .A1(n11890), .A2(n11906), .ZN(n13846) );
  NAND2_X1 U7913 ( .A1(n7415), .A2(n7227), .ZN(n7223) );
  NAND2_X1 U7914 ( .A1(n11888), .A2(n9602), .ZN(n13883) );
  OR2_X1 U7915 ( .A1(n14102), .A2(n13741), .ZN(n11903) );
  NAND2_X1 U7916 ( .A1(n13900), .A2(n13910), .ZN(n13899) );
  NAND2_X1 U7917 ( .A1(n7195), .A2(n6534), .ZN(n13917) );
  NAND2_X1 U7918 ( .A1(n13963), .A2(n13622), .ZN(n7235) );
  OR2_X1 U7919 ( .A1(n14130), .A2(n13623), .ZN(n6805) );
  NAND2_X1 U7920 ( .A1(n7178), .A2(n11884), .ZN(n7174) );
  OR2_X1 U7921 ( .A1(n7175), .A2(n7173), .ZN(n7172) );
  INV_X1 U7922 ( .A(n7178), .ZN(n7173) );
  AND2_X1 U7923 ( .A1(n7176), .A2(n14015), .ZN(n7175) );
  OR2_X1 U7924 ( .A1(n14031), .A2(n7177), .ZN(n7176) );
  NAND2_X1 U7925 ( .A1(n6517), .A2(n14031), .ZN(n14030) );
  OR2_X1 U7926 ( .A1(n12053), .A2(n12057), .ZN(n11738) );
  NOR2_X1 U7927 ( .A1(n6815), .A2(n6814), .ZN(n6817) );
  INV_X1 U7928 ( .A(n11739), .ZN(n6815) );
  INV_X1 U7929 ( .A(n11736), .ZN(n11733) );
  AND2_X1 U7930 ( .A1(n11673), .A2(n7244), .ZN(n11716) );
  NAND2_X1 U7931 ( .A1(n11369), .A2(n11368), .ZN(n11673) );
  AND4_X1 U7932 ( .A1(n9334), .A2(n9333), .A3(n9332), .A4(n9331), .ZN(n12038)
         );
  INV_X1 U7933 ( .A(n6807), .ZN(n6806) );
  OAI21_X1 U7934 ( .B1(n6808), .B2(n11109), .A(n11313), .ZN(n6807) );
  OR2_X1 U7935 ( .A1(n14431), .A2(n13746), .ZN(n11306) );
  AND2_X1 U7936 ( .A1(n7213), .A2(n10996), .ZN(n7212) );
  OR2_X1 U7937 ( .A1(n10955), .A2(n7214), .ZN(n7213) );
  INV_X1 U7938 ( .A(n10921), .ZN(n7214) );
  CLKBUF_X1 U7939 ( .A(n10951), .Z(n6644) );
  NAND2_X1 U7940 ( .A1(n6644), .A2(n10955), .ZN(n10950) );
  AND3_X1 U7941 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n9200) );
  NAND2_X1 U7942 ( .A1(n14541), .A2(n10226), .ZN(n14540) );
  INV_X1 U7943 ( .A(n14556), .ZN(n14058) );
  INV_X1 U7944 ( .A(n14562), .ZN(n14055) );
  OR2_X1 U7945 ( .A1(n10216), .A2(n9665), .ZN(n14542) );
  AND2_X2 U7946 ( .A1(n9193), .A2(n9192), .ZN(n10685) );
  XNOR2_X1 U7947 ( .A(n8208), .B(n7307), .ZN(n12159) );
  OAI21_X1 U7948 ( .B1(n8127), .B2(n7312), .A(n7310), .ZN(n8208) );
  INV_X1 U7949 ( .A(n7356), .ZN(n7354) );
  INV_X1 U7950 ( .A(n9067), .ZN(n9659) );
  XNOR2_X1 U7951 ( .A(n8039), .B(SI_22_), .ZN(n9461) );
  XNOR2_X1 U7952 ( .A(n7992), .B(n7991), .ZN(n11256) );
  NAND2_X1 U7953 ( .A1(n7291), .A2(n7295), .ZN(n7801) );
  NAND2_X1 U7954 ( .A1(n7760), .A2(n7296), .ZN(n7291) );
  NAND2_X1 U7955 ( .A1(n7284), .A2(n7553), .ZN(n7533) );
  INV_X1 U7956 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n6691) );
  OAI21_X1 U7957 ( .B1(n14317), .B2(n14316), .A(P2_ADDR_REG_9__SCAN_IN), .ZN(
        n6671) );
  OAI21_X1 U7958 ( .B1(n14459), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n6522), .ZN(
        n6964) );
  AOI22_X1 U7959 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14289), .B1(n14290), 
        .B2(n14227), .ZN(n14237) );
  AOI21_X1 U7960 ( .B1(n11170), .B2(n8956), .A(n7407), .ZN(n11231) );
  NAND2_X1 U7961 ( .A1(n11231), .A2(n7273), .ZN(n11344) );
  AND2_X1 U7962 ( .A1(n8959), .A2(n11345), .ZN(n7273) );
  NOR2_X1 U7963 ( .A1(n12523), .A2(n12219), .ZN(n12222) );
  NAND2_X1 U7964 ( .A1(n12365), .A2(n9027), .ZN(n12479) );
  AND3_X1 U7965 ( .A1(n8695), .A2(n8694), .A3(n8693), .ZN(n12759) );
  AND4_X1 U7966 ( .A1(n8535), .A2(n8534), .A3(n8533), .A4(n8532), .ZN(n12876)
         );
  INV_X1 U7967 ( .A(n12503), .ZN(n12665) );
  AND2_X1 U7968 ( .A1(n12509), .A2(n8971), .ZN(n8972) );
  XNOR2_X1 U7969 ( .A(n12194), .B(n12193), .ZN(n6701) );
  NAND2_X1 U7970 ( .A1(n12190), .A2(n12189), .ZN(n12191) );
  INV_X1 U7971 ( .A(n7144), .ZN(n6699) );
  AND3_X1 U7972 ( .A1(n12190), .A2(n6755), .A3(n6754), .ZN(n12217) );
  XNOR2_X1 U7973 ( .A(n11383), .B(n11422), .ZN(n14894) );
  NAND2_X1 U7974 ( .A1(n14344), .A2(n6694), .ZN(n12622) );
  OR2_X1 U7975 ( .A1(n14342), .A2(n12972), .ZN(n6694) );
  NOR2_X1 U7976 ( .A1(n12608), .A2(n7045), .ZN(n7038) );
  INV_X1 U7977 ( .A(n7039), .ZN(n7036) );
  INV_X1 U7978 ( .A(n13001), .ZN(n12638) );
  NAND2_X1 U7979 ( .A1(n8710), .A2(n8709), .ZN(n12721) );
  OAI211_X1 U7980 ( .C1(n9716), .C2(n8463), .A(n8467), .B(n8466), .ZN(n11358)
         );
  INV_X1 U7981 ( .A(n12219), .ZN(n10811) );
  AND2_X1 U7982 ( .A1(n8851), .A2(n8850), .ZN(n13054) );
  OR2_X1 U7983 ( .A1(n9759), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8851) );
  AND2_X1 U7984 ( .A1(n8849), .A2(n8848), .ZN(n13056) );
  OR2_X1 U7985 ( .A1(n9759), .A2(P3_D_REG_0__SCAN_IN), .ZN(n8849) );
  INV_X1 U7986 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13058) );
  MUX2_X1 U7987 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8358), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n8361) );
  INV_X1 U7988 ( .A(SI_11_), .ZN(n15202) );
  NAND2_X1 U7989 ( .A1(n11829), .A2(n11828), .ZN(n14662) );
  NAND2_X1 U7990 ( .A1(n14662), .A2(n7112), .ZN(n14372) );
  INV_X1 U7991 ( .A(n10862), .ZN(n10863) );
  NAND2_X1 U7992 ( .A1(n7945), .A2(n7944), .ZN(n13528) );
  AOI21_X1 U7993 ( .B1(n7106), .B2(n13165), .A(n11962), .ZN(n7104) );
  NAND2_X1 U7994 ( .A1(n13106), .A2(n13105), .ZN(n13104) );
  NAND2_X1 U7995 ( .A1(n7878), .A2(n7877), .ZN(n14388) );
  NAND3_X1 U7996 ( .A1(n11917), .A2(n6830), .A3(n10203), .ZN(n6832) );
  INV_X1 U7997 ( .A(n10289), .ZN(n6830) );
  NAND2_X1 U7998 ( .A1(n6835), .A2(n6834), .ZN(n6833) );
  INV_X1 U7999 ( .A(n10287), .ZN(n6834) );
  INV_X1 U8000 ( .A(n10288), .ZN(n6835) );
  XNOR2_X1 U8001 ( .A(n11944), .B(n11943), .ZN(n13149) );
  NAND2_X1 U8002 ( .A1(n10330), .A2(n10121), .ZN(n14664) );
  NAND2_X1 U8003 ( .A1(n7857), .A2(n7856), .ZN(n13546) );
  NAND2_X1 U8004 ( .A1(n7764), .A2(n7763), .ZN(n11183) );
  NAND2_X1 U8005 ( .A1(n6544), .A2(n8281), .ZN(n7052) );
  NAND2_X1 U8006 ( .A1(n9819), .A2(n7051), .ZN(n7050) );
  AND2_X1 U8007 ( .A1(n13432), .A2(n13257), .ZN(n13455) );
  OAI211_X1 U8008 ( .C1(n13473), .C2(n14812), .A(n13472), .B(n6894), .ZN(
        n13559) );
  NAND2_X1 U8009 ( .A1(n13471), .A2(n14816), .ZN(n6952) );
  INV_X1 U8010 ( .A(n13470), .ZN(n6953) );
  AND2_X1 U8011 ( .A1(n6542), .A2(n7443), .ZN(n6985) );
  INV_X1 U8012 ( .A(n7474), .ZN(n6986) );
  NAND2_X1 U8013 ( .A1(n6793), .A2(n12138), .ZN(n6792) );
  NAND2_X1 U8014 ( .A1(n13718), .A2(n13719), .ZN(n6793) );
  INV_X1 U8015 ( .A(n13596), .ZN(n6791) );
  NAND2_X1 U8016 ( .A1(n9478), .A2(n9477), .ZN(n14108) );
  AND2_X1 U8017 ( .A1(n11606), .A2(n6501), .ZN(n6798) );
  OR2_X1 U8018 ( .A1(n10317), .A2(n10316), .ZN(n10318) );
  NAND2_X1 U8019 ( .A1(n7344), .A2(n6551), .ZN(n13612) );
  AOI21_X1 U8020 ( .B1(n6788), .B2(n6790), .A(n6557), .ZN(n6785) );
  AND2_X1 U8021 ( .A1(n9339), .A2(n9338), .ZN(n14443) );
  NAND2_X1 U8022 ( .A1(n9971), .A2(n9970), .ZN(n14426) );
  NAND2_X1 U8023 ( .A1(n10325), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14436) );
  AND2_X1 U8024 ( .A1(n11472), .A2(n14606), .ZN(n14432) );
  INV_X1 U8025 ( .A(n9561), .ZN(n13739) );
  INV_X1 U8026 ( .A(n11165), .ZN(n13826) );
  NAND2_X1 U8027 ( .A1(n9073), .A2(n9072), .ZN(n14071) );
  NAND2_X1 U8028 ( .A1(n7179), .A2(n6639), .ZN(n13847) );
  NOR2_X1 U8029 ( .A1(n6640), .A2(n6562), .ZN(n6639) );
  NAND2_X1 U8030 ( .A1(n9319), .A2(n9318), .ZN(n14411) );
  NAND2_X1 U8031 ( .A1(n11165), .A2(n14576), .ZN(n13947) );
  INV_X1 U8032 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14174) );
  INV_X1 U8033 ( .A(n14271), .ZN(n6966) );
  XNOR2_X1 U8034 ( .A(n14288), .B(n14287), .ZN(n14459) );
  NAND2_X1 U8035 ( .A1(n14462), .A2(n14461), .ZN(n14460) );
  INV_X1 U8036 ( .A(n14297), .ZN(n6959) );
  INV_X1 U8037 ( .A(n14298), .ZN(n6960) );
  NAND2_X1 U8038 ( .A1(n15018), .A2(n15017), .ZN(n15019) );
  OAI21_X1 U8039 ( .B1(n15018), .B2(n15017), .A(n14305), .ZN(n6969) );
  NAND2_X1 U8040 ( .A1(n10337), .A2(n10333), .ZN(n6977) );
  NAND2_X1 U8041 ( .A1(n7627), .A2(n7628), .ZN(n7402) );
  NAND2_X1 U8042 ( .A1(n7400), .A2(n7405), .ZN(n7404) );
  INV_X1 U8043 ( .A(n7628), .ZN(n7405) );
  INV_X1 U8044 ( .A(n7627), .ZN(n7400) );
  INV_X1 U8045 ( .A(n7674), .ZN(n7393) );
  AOI21_X1 U8046 ( .B1(n7392), .B2(n7391), .A(n6584), .ZN(n7390) );
  NOR2_X1 U8047 ( .A1(n7381), .A2(n7380), .ZN(n7379) );
  INV_X1 U8048 ( .A(n7728), .ZN(n7381) );
  INV_X1 U8049 ( .A(n9275), .ZN(n6636) );
  INV_X1 U8050 ( .A(n7775), .ZN(n7395) );
  AND2_X1 U8051 ( .A1(n11711), .A2(n9343), .ZN(n9344) );
  INV_X1 U8052 ( .A(n7889), .ZN(n6657) );
  NAND2_X1 U8053 ( .A1(n7384), .A2(n7889), .ZN(n7383) );
  NAND2_X1 U8054 ( .A1(n7388), .A2(n7385), .ZN(n7384) );
  AND2_X1 U8055 ( .A1(n7864), .A2(n7865), .ZN(n7388) );
  AOI21_X1 U8056 ( .B1(n7115), .B2(n6506), .A(n7168), .ZN(n7114) );
  NAND2_X1 U8057 ( .A1(n6724), .A2(n6723), .ZN(n12294) );
  NOR2_X1 U8058 ( .A1(n12866), .A2(n12287), .ZN(n6723) );
  INV_X1 U8059 ( .A(n6725), .ZN(n6724) );
  AOI21_X1 U8060 ( .B1(n6716), .B2(n12211), .A(n12796), .ZN(n6714) );
  NAND2_X1 U8061 ( .A1(n7374), .A2(n7373), .ZN(n7372) );
  NAND2_X1 U8062 ( .A1(n7918), .A2(n6556), .ZN(n7371) );
  INV_X1 U8063 ( .A(n9479), .ZN(n6645) );
  INV_X1 U8064 ( .A(n9480), .ZN(n6646) );
  AOI21_X1 U8065 ( .B1(n6710), .B2(n6712), .A(n6576), .ZN(n6709) );
  NOR2_X1 U8066 ( .A1(n6707), .A2(n12706), .ZN(n6706) );
  INV_X1 U8067 ( .A(n12327), .ZN(n6707) );
  NAND2_X1 U8068 ( .A1(n7398), .A2(n6608), .ZN(n7397) );
  NAND2_X1 U8069 ( .A1(n9523), .A2(n9525), .ZN(n7120) );
  NAND2_X1 U8070 ( .A1(n7152), .A2(n7151), .ZN(n6721) );
  NAND2_X1 U8071 ( .A1(n7150), .A2(n7149), .ZN(n6720) );
  NOR2_X1 U8072 ( .A1(n12334), .A2(n12346), .ZN(n7151) );
  INV_X1 U8073 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8348) );
  INV_X1 U8074 ( .A(n8325), .ZN(n7142) );
  INV_X1 U8075 ( .A(n8327), .ZN(n7141) );
  INV_X1 U8076 ( .A(n8660), .ZN(n7143) );
  INV_X1 U8077 ( .A(n8645), .ZN(n7139) );
  NAND2_X1 U8078 ( .A1(n7365), .A2(n8076), .ZN(n7364) );
  INV_X1 U8079 ( .A(n7366), .ZN(n7365) );
  NOR2_X1 U8080 ( .A1(n8055), .A2(n7370), .ZN(n7366) );
  INV_X1 U8081 ( .A(n8115), .ZN(n7367) );
  INV_X1 U8082 ( .A(n8114), .ZN(n7368) );
  INV_X1 U8083 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6843) );
  AOI21_X1 U8084 ( .B1(n7316), .B2(n7318), .A(n7314), .ZN(n7313) );
  INV_X1 U8085 ( .A(n7975), .ZN(n7314) );
  NAND2_X1 U8086 ( .A1(n7730), .A2(SI_10_), .ZN(n7755) );
  INV_X1 U8087 ( .A(P2_RD_REG_SCAN_IN), .ZN(n14307) );
  INV_X1 U8088 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7465) );
  INV_X1 U8089 ( .A(n12450), .ZN(n7266) );
  NAND2_X1 U8090 ( .A1(n14886), .A2(n11394), .ZN(n11395) );
  INV_X1 U8091 ( .A(n7022), .ZN(n6768) );
  INV_X1 U8092 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8351) );
  INV_X1 U8093 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7276) );
  INV_X1 U8094 ( .A(n7045), .ZN(n7043) );
  NAND2_X1 U8095 ( .A1(n8885), .A2(n7131), .ZN(n12354) );
  AND2_X1 U8096 ( .A1(n7132), .A2(n8884), .ZN(n7131) );
  NAND2_X1 U8097 ( .A1(n7133), .A2(n12384), .ZN(n12350) );
  OR2_X1 U8098 ( .A1(n12391), .A2(n12652), .ZN(n8899) );
  AND2_X1 U8099 ( .A1(n12698), .A2(n12696), .ZN(n12332) );
  INV_X1 U8100 ( .A(n8824), .ZN(n6861) );
  INV_X1 U8101 ( .A(n12320), .ZN(n6926) );
  INV_X1 U8102 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n15136) );
  NOR2_X1 U8103 ( .A1(n8622), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n6682) );
  NOR2_X1 U8104 ( .A1(n8587), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8374) );
  INV_X1 U8105 ( .A(n6857), .ZN(n6856) );
  NOR2_X1 U8106 ( .A1(n8529), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n6683) );
  OR2_X1 U8107 ( .A1(n11174), .A2(n8792), .ZN(n6924) );
  OR2_X1 U8108 ( .A1(n9759), .A2(n8863), .ZN(n8902) );
  NOR2_X1 U8109 ( .A1(n12763), .A2(n6930), .ZN(n6929) );
  INV_X1 U8110 ( .A(n12316), .ZN(n6930) );
  NAND2_X1 U8111 ( .A1(n8708), .A2(n8707), .ZN(n6729) );
  AOI21_X1 U8112 ( .B1(n7138), .B2(n6747), .A(n6746), .ZN(n6745) );
  INV_X1 U8113 ( .A(n8322), .ZN(n6747) );
  INV_X1 U8114 ( .A(n7140), .ZN(n6746) );
  AOI21_X1 U8115 ( .B1(n8660), .B2(n7142), .A(n7141), .ZN(n7140) );
  INV_X1 U8116 ( .A(n7275), .ZN(n8617) );
  INV_X1 U8117 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8561) );
  INV_X1 U8118 ( .A(n6733), .ZN(n6732) );
  AOI21_X1 U8119 ( .B1(n6733), .B2(n6734), .A(n6614), .ZN(n6731) );
  AOI21_X1 U8120 ( .B1(n7145), .B2(n7147), .A(n8553), .ZN(n6733) );
  NOR2_X1 U8121 ( .A1(n8550), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n8562) );
  OR2_X1 U8122 ( .A1(n8492), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8501) );
  INV_X1 U8123 ( .A(n8297), .ZN(n6741) );
  AOI21_X1 U8124 ( .B1(n13089), .B2(n6515), .A(n7089), .ZN(n7088) );
  INV_X1 U8125 ( .A(n13134), .ZN(n7089) );
  NAND2_X1 U8126 ( .A1(n7085), .A2(n7087), .ZN(n7082) );
  INV_X1 U8127 ( .A(n11828), .ZN(n7110) );
  NAND2_X1 U8128 ( .A1(n6572), .A2(n7319), .ZN(n8232) );
  NAND2_X1 U8129 ( .A1(n6588), .A2(n7320), .ZN(n7319) );
  NOR2_X1 U8130 ( .A1(n8200), .A2(n8201), .ZN(n7320) );
  NAND2_X1 U8131 ( .A1(n8141), .A2(n8140), .ZN(n8236) );
  INV_X1 U8132 ( .A(n7007), .ZN(n7006) );
  AND2_X1 U8133 ( .A1(n6949), .A2(n13483), .ZN(n6948) );
  AND2_X1 U8134 ( .A1(n7926), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7946) );
  INV_X1 U8135 ( .A(n11178), .ZN(n7059) );
  INV_X1 U8136 ( .A(n7058), .ZN(n7057) );
  OAI21_X1 U8137 ( .B1(n7060), .B2(n7059), .A(n11295), .ZN(n7058) );
  NOR2_X1 U8138 ( .A1(n10888), .A2(n6981), .ZN(n6980) );
  INV_X1 U8139 ( .A(n10730), .ZN(n6981) );
  NAND2_X1 U8140 ( .A1(n6994), .A2(n10657), .ZN(n6993) );
  INV_X1 U8141 ( .A(n7442), .ZN(n6841) );
  NOR2_X1 U8142 ( .A1(n7480), .A2(n7479), .ZN(n7481) );
  INV_X1 U8143 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7661) );
  NAND2_X1 U8144 ( .A1(n9960), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6803) );
  NOR2_X1 U8145 ( .A1(n10636), .A2(n6771), .ZN(n6770) );
  INV_X1 U8146 ( .A(n11012), .ZN(n6771) );
  OR2_X1 U8147 ( .A1(n7221), .A2(n7218), .ZN(n7217) );
  INV_X1 U8148 ( .A(n7223), .ZN(n7220) );
  NOR2_X1 U8149 ( .A1(n14095), .A2(n6944), .ZN(n6943) );
  INV_X1 U8150 ( .A(n6945), .ZN(n6944) );
  NOR2_X1 U8151 ( .A1(n7197), .A2(n7201), .ZN(n7194) );
  AND2_X1 U8152 ( .A1(n14108), .A2(n11886), .ZN(n7201) );
  INV_X1 U8153 ( .A(n9439), .ZN(n9455) );
  NOR2_X1 U8154 ( .A1(n7170), .A2(n6813), .ZN(n6812) );
  AND2_X1 U8155 ( .A1(n6814), .A2(n11882), .ZN(n6813) );
  NAND2_X1 U8156 ( .A1(n7171), .A2(n13996), .ZN(n7170) );
  INV_X1 U8157 ( .A(n7174), .ZN(n7171) );
  INV_X1 U8158 ( .A(n7172), .ZN(n6642) );
  NAND2_X1 U8159 ( .A1(n11741), .A2(n11738), .ZN(n6814) );
  NAND2_X1 U8160 ( .A1(n11310), .A2(n6809), .ZN(n6808) );
  INV_X1 U8161 ( .A(n10228), .ZN(n7208) );
  XNOR2_X1 U8162 ( .A(n10685), .B(n13711), .ZN(n10690) );
  NAND2_X1 U8163 ( .A1(n6940), .A2(n11899), .ZN(n14003) );
  AOI21_X1 U8164 ( .B1(n8143), .B2(n7311), .A(n6624), .ZN(n7310) );
  INV_X1 U8165 ( .A(n8126), .ZN(n7311) );
  OAI21_X1 U8166 ( .B1(n8077), .B2(n7302), .A(n8080), .ZN(n8096) );
  INV_X1 U8167 ( .A(n8078), .ZN(n7302) );
  OAI21_X1 U8168 ( .B1(n7920), .B2(n6884), .A(n6882), .ZN(n8039) );
  AOI21_X1 U8169 ( .B1(n6885), .B2(n7317), .A(n6883), .ZN(n6882) );
  INV_X1 U8170 ( .A(n6885), .ZN(n6884) );
  INV_X1 U8171 ( .A(n8020), .ZN(n6883) );
  INV_X1 U8172 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9056) );
  INV_X1 U8173 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9055) );
  NAND2_X1 U8174 ( .A1(n6886), .A2(n7313), .ZN(n8021) );
  NAND2_X1 U8175 ( .A1(n7920), .A2(n7316), .ZN(n6886) );
  NAND2_X1 U8176 ( .A1(n7315), .A2(n7921), .ZN(n7969) );
  XNOR2_X1 U8177 ( .A(n7969), .B(SI_18_), .ZN(n7938) );
  NAND2_X1 U8178 ( .A1(n6887), .A2(n6888), .ZN(n7868) );
  AOI21_X1 U8179 ( .B1(n7823), .B2(n6494), .A(n6573), .ZN(n6888) );
  AND2_X1 U8180 ( .A1(n7869), .A2(n7853), .ZN(n7867) );
  AOI21_X1 U8181 ( .B1(n6508), .B2(n7298), .A(n6568), .ZN(n7295) );
  NOR2_X1 U8182 ( .A1(n9237), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9352) );
  INV_X1 U8183 ( .A(SI_2_), .ZN(n7527) );
  NAND2_X1 U8184 ( .A1(n6962), .A2(n14203), .ZN(n14204) );
  INV_X1 U8185 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n6961) );
  OAI21_X1 U8186 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n14209), .A(n14208), .ZN(
        n14210) );
  OAI21_X1 U8187 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14223), .A(n14222), .ZN(
        n14286) );
  NOR2_X1 U8188 ( .A1(n7263), .A2(n8966), .ZN(n7262) );
  INV_X1 U8189 ( .A(n8966), .ZN(n7260) );
  NOR2_X1 U8190 ( .A1(n12420), .A2(n7269), .ZN(n7268) );
  INV_X1 U8191 ( .A(n8984), .ZN(n7269) );
  OR2_X1 U8192 ( .A1(n8983), .A2(n12774), .ZN(n8984) );
  INV_X1 U8193 ( .A(n8701), .ZN(n8378) );
  NOR2_X1 U8194 ( .A1(n7272), .A2(n8963), .ZN(n7271) );
  INV_X1 U8195 ( .A(n8962), .ZN(n7272) );
  NOR2_X1 U8196 ( .A1(n8419), .A2(n8418), .ZN(n11062) );
  NAND2_X1 U8197 ( .A1(n6850), .A2(n6849), .ZN(n10746) );
  NAND2_X1 U8198 ( .A1(n10743), .A2(n10798), .ZN(n6849) );
  NAND2_X1 U8199 ( .A1(n7252), .A2(n6612), .ZN(n12474) );
  NAND2_X1 U8200 ( .A1(n7256), .A2(n12728), .ZN(n7251) );
  NOR2_X1 U8201 ( .A1(n12216), .A2(n12352), .ZN(n6754) );
  AND2_X1 U8202 ( .A1(n12178), .A2(n12177), .ZN(n12632) );
  AND4_X1 U8203 ( .A1(n8473), .A2(n8472), .A3(n8471), .A4(n8470), .ZN(n11101)
         );
  OAI21_X1 U8204 ( .B1(n8779), .B2(n10352), .A(n8395), .ZN(n6719) );
  NAND2_X1 U8205 ( .A1(n7026), .A2(n10448), .ZN(n10386) );
  NAND2_X1 U8206 ( .A1(n6758), .A2(n10447), .ZN(n6757) );
  AND3_X1 U8207 ( .A1(n7026), .A2(n10448), .A3(P3_REG2_REG_3__SCAN_IN), .ZN(
        n6758) );
  NAND2_X1 U8208 ( .A1(n14923), .A2(n11397), .ZN(n11398) );
  NOR2_X1 U8209 ( .A1(n14930), .A2(n11387), .ZN(n14958) );
  INV_X1 U8210 ( .A(n6761), .ZN(n11386) );
  INV_X1 U8211 ( .A(n7028), .ZN(n14956) );
  INV_X1 U8212 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14223) );
  AND2_X1 U8213 ( .A1(n7028), .A2(n7027), .ZN(n11478) );
  NAND2_X1 U8214 ( .A1(n14969), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7027) );
  AOI21_X1 U8215 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n11545), .A(n11536), .ZN(
        n12524) );
  XNOR2_X1 U8216 ( .A(n12528), .B(n12538), .ZN(n11540) );
  NAND2_X1 U8217 ( .A1(n11540), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n12530) );
  AND2_X1 U8218 ( .A1(n12558), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n6760) );
  OR2_X1 U8219 ( .A1(n14330), .A2(n6768), .ZN(n6767) );
  NAND2_X1 U8220 ( .A1(n6764), .A2(n6628), .ZN(n6766) );
  INV_X1 U8221 ( .A(n12597), .ZN(n6764) );
  NAND2_X1 U8222 ( .A1(n12597), .A2(n12618), .ZN(n6765) );
  NAND2_X1 U8223 ( .A1(n14345), .A2(n14346), .ZN(n14344) );
  NOR2_X1 U8224 ( .A1(n12617), .A2(n12825), .ZN(n7022) );
  NOR2_X1 U8225 ( .A1(n14342), .A2(n12600), .ZN(n7045) );
  NAND2_X1 U8226 ( .A1(n7041), .A2(n7040), .ZN(n7039) );
  NAND2_X1 U8227 ( .A1(n12608), .A2(n7043), .ZN(n7040) );
  NAND2_X1 U8228 ( .A1(n7042), .A2(n12611), .ZN(n7041) );
  NAND2_X1 U8229 ( .A1(n14354), .A2(n7043), .ZN(n7042) );
  NAND2_X1 U8230 ( .A1(n6870), .A2(n6869), .ZN(n8878) );
  OR2_X1 U8231 ( .A1(n13007), .A2(n12652), .ZN(n7413) );
  AND2_X1 U8232 ( .A1(n12380), .A2(n6582), .ZN(n6869) );
  OAI21_X1 U8233 ( .B1(n12380), .B2(n6582), .A(n12878), .ZN(n6867) );
  NAND2_X1 U8234 ( .A1(n12347), .A2(n6897), .ZN(n6868) );
  INV_X1 U8235 ( .A(n12334), .ZN(n6903) );
  NAND2_X1 U8236 ( .A1(n6898), .A2(n6896), .ZN(n12648) );
  AOI21_X1 U8237 ( .B1(n6899), .B2(n6902), .A(n6897), .ZN(n6896) );
  NAND2_X1 U8238 ( .A1(n12697), .A2(n6899), .ZN(n6898) );
  OR2_X1 U8239 ( .A1(n12721), .A2(n12728), .ZN(n12696) );
  AND2_X1 U8240 ( .A1(n12324), .A2(n12323), .ZN(n12743) );
  OAI21_X1 U8241 ( .B1(n12970), .B2(n6928), .A(n6925), .ZN(n12747) );
  INV_X1 U8242 ( .A(n6929), .ZN(n6928) );
  AOI21_X1 U8243 ( .B1(n6929), .B2(n6927), .A(n6926), .ZN(n6925) );
  INV_X1 U8244 ( .A(n6932), .ZN(n6927) );
  NAND2_X1 U8245 ( .A1(n8376), .A2(n8375), .ZN(n8679) );
  INV_X1 U8246 ( .A(n8667), .ZN(n8376) );
  OR2_X1 U8247 ( .A1(n8653), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U8248 ( .A1(n8817), .A2(n8816), .ZN(n12736) );
  AND4_X1 U8249 ( .A1(n8644), .A2(n8643), .A3(n8642), .A4(n8641), .ZN(n12791)
         );
  NAND2_X1 U8250 ( .A1(n6682), .A2(n15136), .ZN(n8653) );
  NAND2_X1 U8251 ( .A1(n8374), .A2(n8373), .ZN(n8622) );
  INV_X1 U8252 ( .A(n6682), .ZN(n8638) );
  INV_X1 U8253 ( .A(n8813), .ZN(n12821) );
  AND2_X1 U8254 ( .A1(n12291), .A2(n12299), .ZN(n12833) );
  INV_X1 U8255 ( .A(n8374), .ZN(n8606) );
  NAND2_X1 U8256 ( .A1(n6854), .A2(n6855), .ZN(n12842) );
  OAI22_X1 U8257 ( .A1(n11565), .A2(n6918), .B1(n6920), .B2(n8558), .ZN(n12864) );
  AND2_X1 U8258 ( .A1(n8559), .A2(n6921), .ZN(n6920) );
  NAND2_X1 U8259 ( .A1(n8557), .A2(n6923), .ZN(n6918) );
  NAND2_X1 U8260 ( .A1(n6683), .A2(n15111), .ZN(n8569) );
  INV_X1 U8261 ( .A(n6683), .ZN(n8544) );
  INV_X1 U8262 ( .A(n12899), .ZN(n12901) );
  AND2_X1 U8263 ( .A1(n12279), .A2(n12284), .ZN(n12899) );
  NAND2_X1 U8264 ( .A1(n8371), .A2(n8370), .ZN(n8515) );
  INV_X1 U8265 ( .A(n8509), .ZN(n8371) );
  NOR2_X1 U8266 ( .A1(n8528), .A2(n8527), .ZN(n12275) );
  NAND2_X1 U8267 ( .A1(n6919), .A2(n6923), .ZN(n12893) );
  NAND2_X1 U8268 ( .A1(n11565), .A2(n6924), .ZN(n6919) );
  INV_X1 U8269 ( .A(n12200), .ZN(n12268) );
  AND4_X2 U8270 ( .A1(n8487), .A2(n8486), .A3(n8485), .A4(n8484), .ZN(n11562)
         );
  INV_X1 U8271 ( .A(n8468), .ZN(n8369) );
  AOI21_X1 U8272 ( .B1(n6912), .B2(n6914), .A(n6909), .ZN(n6908) );
  INV_X1 U8273 ( .A(n12249), .ZN(n6909) );
  AND2_X1 U8274 ( .A1(n12255), .A2(n12256), .ZN(n12197) );
  INV_X1 U8275 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8367) );
  INV_X1 U8276 ( .A(n12906), .ZN(n12847) );
  INV_X1 U8277 ( .A(n10538), .ZN(n12221) );
  NAND2_X1 U8278 ( .A1(n6904), .A2(n6905), .ZN(n12664) );
  NAND2_X1 U8279 ( .A1(n8730), .A2(n8729), .ZN(n12933) );
  NAND2_X1 U8280 ( .A1(n6931), .A2(n6929), .ZN(n12957) );
  NAND2_X1 U8281 ( .A1(n6931), .A2(n12316), .ZN(n12764) );
  NAND2_X1 U8282 ( .A1(n8621), .A2(n8620), .ZN(n12978) );
  OR2_X1 U8283 ( .A1(n10010), .A2(n8463), .ZN(n8621) );
  OR2_X1 U8284 ( .A1(n8903), .A2(n8906), .ZN(n9020) );
  NAND2_X1 U8285 ( .A1(n6756), .A2(n8883), .ZN(n12162) );
  NAND2_X1 U8286 ( .A1(n8881), .A2(n8880), .ZN(n6756) );
  AOI21_X1 U8287 ( .B1(n6751), .B2(n6749), .A(n6630), .ZN(n6748) );
  INV_X1 U8288 ( .A(n6751), .ZN(n6750) );
  NAND2_X1 U8289 ( .A1(n7258), .A2(n8843), .ZN(n6936) );
  INV_X1 U8290 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8834) );
  OAI21_X1 U8291 ( .B1(n8833), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8835) );
  XNOR2_X1 U8292 ( .A(n8767), .B(P3_IR_REG_20__SCAN_IN), .ZN(n8904) );
  XNOR2_X1 U8293 ( .A(n8662), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12609) );
  NAND2_X1 U8294 ( .A1(n6727), .A2(n7157), .ZN(n8614) );
  AOI21_X1 U8295 ( .B1(n6604), .B2(n8314), .A(n7158), .ZN(n7157) );
  INV_X1 U8296 ( .A(n8317), .ZN(n7158) );
  AND2_X1 U8297 ( .A1(n8319), .A2(n8318), .ZN(n8613) );
  NAND2_X1 U8298 ( .A1(n8614), .A2(n8613), .ZN(n8616) );
  INV_X1 U8299 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8539) );
  OR2_X1 U8300 ( .A1(n8538), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n8550) );
  AND2_X1 U8301 ( .A1(n8306), .A2(n8305), .ZN(n8497) );
  NAND2_X1 U8302 ( .A1(n8498), .A2(n8497), .ZN(n8500) );
  NOR2_X1 U8303 ( .A1(n8501), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8505) );
  OR2_X1 U8304 ( .A1(n8464), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8492) );
  INV_X1 U8305 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n6916) );
  AND2_X1 U8306 ( .A1(n8294), .A2(n8293), .ZN(n8437) );
  NAND2_X1 U8307 ( .A1(n7129), .A2(n8289), .ZN(n8426) );
  INV_X1 U8308 ( .A(n7108), .ZN(n6829) );
  INV_X1 U8309 ( .A(n11959), .ZN(n7107) );
  NAND2_X1 U8310 ( .A1(n6827), .A2(n6829), .ZN(n6825) );
  NAND2_X1 U8311 ( .A1(n6515), .A2(n13087), .ZN(n7090) );
  INV_X1 U8312 ( .A(n7088), .ZN(n7087) );
  AND2_X1 U8313 ( .A1(n7086), .A2(n13097), .ZN(n7085) );
  NAND2_X1 U8314 ( .A1(n7088), .A2(n7090), .ZN(n7086) );
  NOR2_X1 U8315 ( .A1(n7903), .A2(n13117), .ZN(n7926) );
  OR2_X1 U8316 ( .A1(n7880), .A2(n7879), .ZN(n7903) );
  NOR2_X1 U8317 ( .A1(n10759), .A2(n10756), .ZN(n7102) );
  OR2_X1 U8318 ( .A1(n10758), .A2(n7101), .ZN(n7100) );
  INV_X1 U8319 ( .A(n10756), .ZN(n7101) );
  NAND2_X1 U8320 ( .A1(n7946), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n7996) );
  OR2_X1 U8321 ( .A1(n7787), .A2(n7786), .ZN(n7808) );
  AND2_X1 U8322 ( .A1(n7735), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7765) );
  AND2_X1 U8323 ( .A1(n7094), .A2(n6590), .ZN(n7092) );
  NAND2_X1 U8324 ( .A1(n13104), .A2(n6837), .ZN(n7105) );
  NOR2_X1 U8325 ( .A1(n13165), .A2(n11954), .ZN(n6837) );
  NOR2_X1 U8326 ( .A1(n10136), .A2(n10137), .ZN(n10125) );
  INV_X1 U8327 ( .A(n10338), .ZN(n7282) );
  OR2_X1 U8328 ( .A1(n8184), .A2(n10563), .ZN(n7624) );
  NAND2_X1 U8329 ( .A1(n6479), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7503) );
  AOI21_X1 U8330 ( .B1(n13210), .B2(P2_REG2_REG_4__SCAN_IN), .A(n13207), .ZN(
        n14716) );
  AOI21_X1 U8331 ( .B1(n10980), .B2(P2_REG2_REG_10__SCAN_IN), .A(n10973), .ZN(
        n13220) );
  XNOR2_X1 U8332 ( .A(n11761), .B(n11750), .ZN(n10977) );
  OR2_X1 U8333 ( .A1(n7826), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n7854) );
  NAND2_X1 U8334 ( .A1(n8213), .A2(n8212), .ZN(n13269) );
  NAND2_X1 U8335 ( .A1(n7006), .A2(n12012), .ZN(n7005) );
  AOI21_X1 U8336 ( .B1(n7067), .B2(n13318), .A(n6574), .ZN(n7065) );
  INV_X1 U8337 ( .A(n7012), .ZN(n13283) );
  INV_X1 U8338 ( .A(n13278), .ZN(n7011) );
  AND2_X1 U8339 ( .A1(n13335), .A2(n11989), .ZN(n6675) );
  INV_X1 U8340 ( .A(n8066), .ZN(n8067) );
  NAND2_X1 U8341 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n8067), .ZN(n8101) );
  NAND2_X1 U8342 ( .A1(n6988), .A2(n6987), .ZN(n13378) );
  AOI21_X1 U8343 ( .B1(n6989), .B2(n11984), .A(n6541), .ZN(n6987) );
  AOI21_X1 U8344 ( .B1(n13448), .B2(n6496), .A(n7077), .ZN(n7076) );
  NOR2_X1 U8345 ( .A1(n13425), .A2(n11999), .ZN(n7077) );
  AOI21_X1 U8346 ( .B1(n7081), .B2(n7079), .A(n6500), .ZN(n7078) );
  INV_X1 U8347 ( .A(n7081), .ZN(n7080) );
  NAND2_X1 U8348 ( .A1(n11649), .A2(n11648), .ZN(n11781) );
  AOI21_X1 U8349 ( .B1(n7018), .B2(n11325), .A(n6565), .ZN(n7017) );
  OR2_X1 U8350 ( .A1(n7808), .A2(n14658), .ZN(n7831) );
  OR2_X1 U8351 ( .A1(n14670), .A2(n11328), .ZN(n7020) );
  OR2_X1 U8352 ( .A1(n11326), .A2(n11325), .ZN(n7021) );
  NAND2_X1 U8353 ( .A1(n7018), .A2(n7021), .ZN(n11652) );
  NOR2_X1 U8354 ( .A1(n11083), .A2(n11183), .ZN(n11192) );
  OR2_X1 U8355 ( .A1(n10894), .A2(n11072), .ZN(n11083) );
  INV_X1 U8356 ( .A(n11070), .ZN(n6983) );
  OR2_X1 U8357 ( .A1(n7685), .A2(n9980), .ZN(n7718) );
  NOR2_X1 U8358 ( .A1(n7718), .A2(n7717), .ZN(n7735) );
  NAND2_X1 U8359 ( .A1(n10728), .A2(n10727), .ZN(n6982) );
  NAND2_X1 U8360 ( .A1(n10734), .A2(n10737), .ZN(n10894) );
  NAND2_X1 U8361 ( .A1(n10575), .A2(n10576), .ZN(n6997) );
  INV_X1 U8362 ( .A(n10573), .ZN(n10574) );
  NAND2_X1 U8363 ( .A1(n10574), .A2(n6994), .ZN(n10652) );
  AND2_X1 U8364 ( .A1(n10542), .A2(n8241), .ZN(n10608) );
  XNOR2_X1 U8365 ( .A(n10843), .B(n10545), .ZN(n10167) );
  INV_X1 U8366 ( .A(n10160), .ZN(n6957) );
  NAND2_X1 U8367 ( .A1(n10145), .A2(n10144), .ZN(n10163) );
  NAND2_X1 U8368 ( .A1(n7049), .A2(n12003), .ZN(n13384) );
  NAND2_X1 U8369 ( .A1(n9742), .A2(n8210), .ZN(n7639) );
  NAND2_X1 U8370 ( .A1(n10561), .A2(n10077), .ZN(n14837) );
  INV_X1 U8371 ( .A(n14837), .ZN(n14816) );
  NAND2_X1 U8372 ( .A1(n10047), .A2(n10046), .ZN(n14790) );
  XNOR2_X1 U8373 ( .A(n8268), .B(n8270), .ZN(n9818) );
  OR2_X1 U8374 ( .A1(n7707), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n7709) );
  INV_X1 U8375 ( .A(n9454), .ZN(n9471) );
  INV_X1 U8376 ( .A(n13740), .ZN(n13721) );
  NOR2_X1 U8377 ( .A1(n11208), .A2(n7349), .ZN(n7348) );
  INV_X1 U8378 ( .A(n11205), .ZN(n7349) );
  OAI22_X1 U8379 ( .A1(n10220), .A2(n12107), .B1(n14563), .B2(n12106), .ZN(
        n10017) );
  INV_X1 U8380 ( .A(n9485), .ZN(n9497) );
  INV_X1 U8381 ( .A(n6789), .ZN(n6788) );
  OAI21_X1 U8382 ( .B1(n6790), .B2(n7341), .A(n13661), .ZN(n6789) );
  AOI21_X1 U8383 ( .B1(n7341), .B2(n7343), .A(n6555), .ZN(n7340) );
  NAND2_X1 U8384 ( .A1(n9956), .A2(n10323), .ZN(n12107) );
  NAND2_X1 U8385 ( .A1(n7346), .A2(n6520), .ZN(n7345) );
  INV_X1 U8386 ( .A(n7348), .ZN(n7346) );
  OR2_X1 U8387 ( .A1(n9419), .A2(n9418), .ZN(n9426) );
  NAND2_X1 U8388 ( .A1(n13689), .A2(n13690), .ZN(n13688) );
  INV_X1 U8389 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9278) );
  NAND2_X1 U8390 ( .A1(n9393), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9407) );
  OR2_X1 U8391 ( .A1(n9329), .A2(n9320), .ZN(n9357) );
  INV_X1 U8392 ( .A(n9567), .ZN(n9574) );
  OR2_X1 U8393 ( .A1(n9569), .A2(n6649), .ZN(n9150) );
  NOR2_X1 U8394 ( .A1(n13870), .A2(n7186), .ZN(n6640) );
  NAND2_X1 U8395 ( .A1(n11906), .A2(n13851), .ZN(n7186) );
  NAND2_X1 U8396 ( .A1(n7184), .A2(n7185), .ZN(n7183) );
  NAND2_X1 U8397 ( .A1(n7187), .A2(n13851), .ZN(n7182) );
  INV_X1 U8398 ( .A(n7187), .ZN(n7181) );
  NAND2_X1 U8399 ( .A1(n6822), .A2(n7218), .ZN(n13870) );
  NAND2_X1 U8400 ( .A1(n13884), .A2(n11888), .ZN(n6822) );
  NAND2_X1 U8401 ( .A1(n13872), .A2(n14055), .ZN(n6820) );
  INV_X1 U8402 ( .A(n9470), .ZN(n9486) );
  NAND2_X1 U8403 ( .A1(n13958), .A2(n6945), .ZN(n13924) );
  AND2_X1 U8404 ( .A1(n7193), .A2(n7194), .ZN(n13919) );
  NAND2_X1 U8405 ( .A1(n13958), .A2(n13942), .ZN(n13941) );
  AND2_X1 U8406 ( .A1(n7169), .A2(n7167), .ZN(n13981) );
  AOI21_X1 U8407 ( .B1(n6642), .B2(n13996), .A(n6641), .ZN(n7167) );
  OAI21_X1 U8408 ( .B1(n11739), .B2(n6816), .A(n6812), .ZN(n7169) );
  INV_X1 U8409 ( .A(n11885), .ZN(n6641) );
  NAND2_X1 U8410 ( .A1(n13981), .A2(n13980), .ZN(n13979) );
  NAND2_X1 U8411 ( .A1(n11899), .A2(n13654), .ZN(n7229) );
  AND2_X1 U8412 ( .A1(n11897), .A2(n9603), .ZN(n14028) );
  NAND2_X1 U8413 ( .A1(n7241), .A2(n6498), .ZN(n7240) );
  NAND2_X1 U8414 ( .A1(n11733), .A2(n7242), .ZN(n7241) );
  INV_X1 U8415 ( .A(n14443), .ZN(n11671) );
  OR3_X1 U8416 ( .A1(n9279), .A2(n9277), .A3(n9278), .ZN(n9299) );
  INV_X1 U8417 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11811) );
  NOR2_X1 U8418 ( .A1(n9299), .A2(n11811), .ZN(n9327) );
  NAND2_X1 U8419 ( .A1(n6811), .A2(n6810), .ZN(n11110) );
  INV_X1 U8420 ( .A(n10924), .ZN(n6810) );
  INV_X1 U8421 ( .A(n10915), .ZN(n6811) );
  NAND2_X1 U8422 ( .A1(n11005), .A2(n11004), .ZN(n11003) );
  AOI21_X1 U8423 ( .B1(n10956), .B2(n10911), .A(n10910), .ZN(n10997) );
  NAND2_X1 U8424 ( .A1(n10323), .A2(n9731), .ZN(n10475) );
  NAND2_X1 U8425 ( .A1(n10466), .A2(n10685), .ZN(n10701) );
  INV_X1 U8426 ( .A(n10690), .ZN(n10689) );
  NAND2_X1 U8427 ( .A1(n10479), .A2(n10234), .ZN(n14541) );
  NAND2_X1 U8428 ( .A1(n6938), .A2(n6937), .ZN(n14555) );
  NAND2_X1 U8429 ( .A1(n10222), .A2(n10221), .ZN(n10478) );
  NAND2_X1 U8430 ( .A1(n10219), .A2(n14060), .ZN(n10222) );
  NOR2_X1 U8431 ( .A1(n14586), .A2(n14565), .ZN(n14048) );
  NOR2_X1 U8432 ( .A1(n7530), .A2(n7508), .ZN(n7238) );
  OR2_X1 U8433 ( .A1(n9137), .A2(n9115), .ZN(n9116) );
  CLKBUF_X1 U8434 ( .A(n10014), .Z(n14563) );
  AND2_X1 U8435 ( .A1(n9565), .A2(n9564), .ZN(n14065) );
  AND2_X1 U8436 ( .A1(n9582), .A2(n9581), .ZN(n14068) );
  AND2_X1 U8437 ( .A1(n13877), .A2(n13876), .ZN(n14083) );
  NAND2_X1 U8438 ( .A1(n9434), .A2(n9433), .ZN(n14130) );
  AND2_X1 U8439 ( .A1(n9382), .A2(n9381), .ZN(n14152) );
  AND2_X1 U8440 ( .A1(n14568), .A2(n9953), .ZN(n14636) );
  INV_X1 U8441 ( .A(n14606), .ZN(n14640) );
  NOR2_X1 U8442 ( .A1(n7309), .A2(n8209), .ZN(n7308) );
  INV_X1 U8443 ( .A(n7305), .ZN(n7304) );
  OAI22_X1 U8444 ( .A1(n7309), .A2(n7306), .B1(n15145), .B2(n8131), .ZN(n7305)
         );
  NAND2_X1 U8445 ( .A1(n7312), .A2(n7307), .ZN(n7306) );
  NOR2_X1 U8446 ( .A1(n7356), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n7355) );
  XNOR2_X1 U8447 ( .A(n8144), .B(n8143), .ZN(n11864) );
  XNOR2_X1 U8448 ( .A(n8160), .B(n8159), .ZN(n12032) );
  XNOR2_X1 U8449 ( .A(n8178), .B(n8177), .ZN(n13589) );
  NAND2_X1 U8450 ( .A1(n9092), .A2(n9388), .ZN(n9402) );
  NOR2_X1 U8451 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n9647) );
  NOR2_X1 U8452 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n9096) );
  XNOR2_X1 U8453 ( .A(n7938), .B(n7966), .ZN(n11105) );
  NAND2_X1 U8454 ( .A1(n6890), .A2(SI_14_), .ZN(n7825) );
  NAND2_X1 U8455 ( .A1(n6889), .A2(n7301), .ZN(n7300) );
  OAI21_X1 U8456 ( .B1(n7659), .B2(n7676), .A(n7286), .ZN(n7700) );
  AND2_X1 U8457 ( .A1(n6823), .A2(n7631), .ZN(n9717) );
  NOR2_X1 U8458 ( .A1(n7615), .A2(n6879), .ZN(n6824) );
  NAND2_X1 U8459 ( .A1(n6876), .A2(n7579), .ZN(n6881) );
  NAND2_X1 U8460 ( .A1(n6880), .A2(n6881), .ZN(n7612) );
  INV_X1 U8461 ( .A(n7584), .ZN(n6880) );
  NAND2_X1 U8462 ( .A1(n6974), .A2(n6972), .ZN(n14243) );
  NAND2_X1 U8463 ( .A1(n6973), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6972) );
  INV_X1 U8464 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6973) );
  XOR2_X1 U8465 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n14196), .Z(n14242) );
  OAI21_X1 U8466 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n14215), .A(n14214), .ZN(
        n14274) );
  OAI21_X1 U8467 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14229), .A(n14228), .ZN(
        n14235) );
  NAND2_X1 U8468 ( .A1(n11033), .A2(n8942), .ZN(n11127) );
  NAND2_X1 U8469 ( .A1(n7256), .A2(n12440), .ZN(n12405) );
  NAND2_X1 U8470 ( .A1(n7270), .A2(n8984), .ZN(n12419) );
  NAND2_X1 U8471 ( .A1(n8690), .A2(n8689), .ZN(n12748) );
  OR2_X1 U8472 ( .A1(n10539), .A2(n8463), .ZN(n8690) );
  NOR2_X1 U8473 ( .A1(n11620), .A2(n11621), .ZN(n11619) );
  AND4_X1 U8474 ( .A1(n8627), .A2(n8626), .A3(n8625), .A4(n8624), .ZN(n12832)
         );
  AND2_X1 U8475 ( .A1(n11033), .A2(n11032), .ZN(n11093) );
  NAND2_X1 U8476 ( .A1(n8980), .A2(n12508), .ZN(n8981) );
  NAND2_X1 U8477 ( .A1(n8700), .A2(n8699), .ZN(n12730) );
  AND2_X1 U8478 ( .A1(n8949), .A2(n11094), .ZN(n11097) );
  NAND2_X1 U8479 ( .A1(n9025), .A2(n9024), .ZN(n12482) );
  INV_X1 U8480 ( .A(n12477), .ZN(n12499) );
  NAND2_X1 U8481 ( .A1(n8759), .A2(n8758), .ZN(n12503) );
  NAND2_X1 U8482 ( .A1(n8746), .A2(n8745), .ZN(n12679) );
  INV_X1 U8483 ( .A(n12791), .ZN(n12818) );
  INV_X1 U8484 ( .A(n12832), .ZN(n12805) );
  INV_X1 U8485 ( .A(n12862), .ZN(n12509) );
  INV_X1 U8486 ( .A(n12876), .ZN(n12511) );
  INV_X1 U8487 ( .A(n11516), .ZN(n12516) );
  INV_X1 U8488 ( .A(n8936), .ZN(n12517) );
  INV_X1 U8489 ( .A(n10825), .ZN(n12518) );
  INV_X1 U8490 ( .A(P3_U3897), .ZN(n12522) );
  INV_X1 U8491 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14246) );
  AND2_X1 U8492 ( .A1(n7025), .A2(n6757), .ZN(n11379) );
  AND2_X1 U8493 ( .A1(n14856), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n14857) );
  NOR2_X1 U8494 ( .A1(n14894), .A2(n11421), .ZN(n14893) );
  NAND2_X1 U8495 ( .A1(n7031), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7030) );
  NAND2_X1 U8496 ( .A1(n11384), .A2(n7031), .ZN(n7029) );
  INV_X1 U8497 ( .A(n14912), .ZN(n7031) );
  XNOR2_X1 U8498 ( .A(n6761), .B(n14938), .ZN(n14931) );
  NOR2_X1 U8499 ( .A1(n14931), .A2(n11434), .ZN(n14930) );
  XNOR2_X1 U8500 ( .A(n11478), .B(n11479), .ZN(n11389) );
  XNOR2_X1 U8501 ( .A(n12524), .B(n12538), .ZN(n11537) );
  NOR2_X1 U8502 ( .A1(n11537), .A2(n8568), .ZN(n12525) );
  OAI21_X1 U8503 ( .B1(n11537), .B2(n7033), .A(n7032), .ZN(n12551) );
  NAND2_X1 U8504 ( .A1(n12542), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7033) );
  NAND2_X1 U8505 ( .A1(n12526), .A2(n12542), .ZN(n7032) );
  XNOR2_X1 U8506 ( .A(n6759), .B(n12577), .ZN(n12552) );
  NOR2_X1 U8507 ( .A1(n12552), .A2(n12553), .ZN(n12572) );
  AND2_X1 U8508 ( .A1(n7024), .A2(n7023), .ZN(n12597) );
  INV_X1 U8509 ( .A(n12574), .ZN(n7023) );
  INV_X1 U8510 ( .A(n7024), .ZN(n12575) );
  NAND2_X1 U8511 ( .A1(n7039), .A2(n7044), .ZN(n7037) );
  OR2_X1 U8512 ( .A1(n12611), .A2(n14354), .ZN(n7044) );
  NAND2_X1 U8513 ( .A1(n12697), .A2(n12330), .ZN(n12682) );
  NAND2_X1 U8514 ( .A1(n7156), .A2(n6619), .ZN(n12702) );
  NAND2_X1 U8515 ( .A1(n6623), .A2(n7530), .ZN(n7156) );
  NAND2_X1 U8516 ( .A1(n9678), .A2(n7155), .ZN(n7154) );
  NAND2_X1 U8517 ( .A1(n12741), .A2(n8822), .ZN(n12726) );
  OR2_X1 U8518 ( .A1(n10456), .A2(n8463), .ZN(n8678) );
  AND2_X1 U8519 ( .A1(n12778), .A2(n12777), .ZN(n12963) );
  NAND2_X1 U8520 ( .A1(n12970), .A2(n12306), .ZN(n12780) );
  NAND2_X1 U8521 ( .A1(n8652), .A2(n8651), .ZN(n12967) );
  NAND2_X1 U8522 ( .A1(n12874), .A2(n12207), .ZN(n6859) );
  NAND2_X1 U8523 ( .A1(n6911), .A2(n12242), .ZN(n11276) );
  NAND2_X1 U8524 ( .A1(n11216), .A2(n12240), .ZN(n6911) );
  NAND2_X1 U8525 ( .A1(n12656), .A2(n10819), .ZN(n12888) );
  INV_X1 U8526 ( .A(n12870), .ZN(n12801) );
  NAND2_X1 U8527 ( .A1(n10714), .A2(n10713), .ZN(n12910) );
  NAND2_X1 U8528 ( .A1(n12914), .A2(n12979), .ZN(n12870) );
  NAND2_X1 U8529 ( .A1(n12171), .A2(n12170), .ZN(n12997) );
  NAND2_X1 U8530 ( .A1(n12184), .A2(n12183), .ZN(n13001) );
  INV_X1 U8531 ( .A(n12339), .ZN(n13011) );
  INV_X1 U8532 ( .A(n9001), .ZN(n13015) );
  OR2_X1 U8533 ( .A1(n12945), .A2(n12944), .ZN(n13018) );
  NAND2_X1 U8534 ( .A1(n8586), .A2(n8585), .ZN(n13046) );
  NAND2_X1 U8535 ( .A1(n8567), .A2(n8566), .ZN(n13052) );
  OR2_X1 U8536 ( .A1(n8663), .A2(n9714), .ZN(n6717) );
  AND2_X1 U8537 ( .A1(n10252), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13055) );
  INV_X1 U8538 ( .A(SI_26_), .ZN(n15171) );
  NAND2_X1 U8539 ( .A1(n6753), .A2(n8340), .ZN(n8739) );
  XNOR2_X1 U8540 ( .A(n8837), .B(n8356), .ZN(n11535) );
  XNOR2_X1 U8541 ( .A(n8844), .B(n8843), .ZN(n11255) );
  XNOR2_X1 U8542 ( .A(n8764), .B(n8763), .ZN(n12218) );
  INV_X1 U8543 ( .A(SI_20_), .ZN(n15090) );
  INV_X1 U8544 ( .A(n8904), .ZN(n10455) );
  NAND2_X1 U8545 ( .A1(n8648), .A2(n8325), .ZN(n8661) );
  INV_X1 U8546 ( .A(SI_17_), .ZN(n10088) );
  INV_X1 U8547 ( .A(SI_16_), .ZN(n15094) );
  INV_X1 U8548 ( .A(SI_15_), .ZN(n15068) );
  NAND2_X1 U8549 ( .A1(n7159), .A2(n6604), .ZN(n8600) );
  NAND2_X1 U8550 ( .A1(n7159), .A2(n8315), .ZN(n8598) );
  INV_X1 U8551 ( .A(n12588), .ZN(n12577) );
  INV_X1 U8552 ( .A(SI_12_), .ZN(n9724) );
  OAI21_X1 U8553 ( .B1(n6730), .B2(n7147), .A(n7145), .ZN(n8554) );
  NAND2_X1 U8554 ( .A1(n8526), .A2(n8308), .ZN(n8537) );
  NAND2_X1 U8555 ( .A1(n8477), .A2(n8302), .ZN(n8489) );
  NAND2_X1 U8556 ( .A1(n8300), .A2(n8299), .ZN(n8475) );
  NAND2_X1 U8557 ( .A1(n6738), .A2(n8297), .ZN(n8462) );
  NAND2_X1 U8558 ( .A1(n8451), .A2(n8450), .ZN(n6738) );
  INV_X1 U8559 ( .A(n11415), .ZN(n14882) );
  NAND2_X1 U8560 ( .A1(n6915), .A2(n6917), .ZN(n8439) );
  INV_X1 U8561 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8345) );
  OR2_X1 U8562 ( .A1(n8280), .A2(n13595), .ZN(n9823) );
  INV_X1 U8563 ( .A(n9818), .ZN(n9822) );
  OAI21_X1 U8564 ( .B1(n6829), .B2(n10298), .A(n6827), .ZN(n10522) );
  NOR2_X1 U8565 ( .A1(n13163), .A2(n11959), .ZN(n13073) );
  NAND2_X1 U8566 ( .A1(n7105), .A2(n7106), .ZN(n13071) );
  NAND2_X1 U8567 ( .A1(n6836), .A2(n10855), .ZN(n10861) );
  NAND2_X1 U8568 ( .A1(n13153), .A2(n6845), .ZN(n13091) );
  NAND2_X1 U8569 ( .A1(n11933), .A2(n6846), .ZN(n6845) );
  INV_X1 U8570 ( .A(n11934), .ZN(n6846) );
  INV_X1 U8571 ( .A(n7083), .ZN(n13098) );
  AOI21_X1 U8572 ( .B1(n13091), .B2(n7084), .A(n7087), .ZN(n7083) );
  INV_X1 U8573 ( .A(n7090), .ZN(n7084) );
  OAI21_X1 U8574 ( .B1(n13091), .B2(n7087), .A(n7085), .ZN(n13096) );
  INV_X1 U8575 ( .A(n11242), .ZN(n11243) );
  AND2_X1 U8576 ( .A1(n11927), .A2(n11926), .ZN(n6847) );
  NAND2_X1 U8577 ( .A1(n14383), .A2(n14382), .ZN(n14381) );
  NAND2_X1 U8578 ( .A1(n10298), .A2(n10299), .ZN(n10420) );
  NAND2_X1 U8579 ( .A1(n7093), .A2(n7094), .ZN(n13115) );
  OAI21_X1 U8580 ( .B1(n10757), .B2(n7102), .A(n7100), .ZN(n10851) );
  AOI21_X1 U8581 ( .B1(n13091), .B2(n13087), .A(n13089), .ZN(n13136) );
  NOR2_X1 U8582 ( .A1(n13149), .A2(n13148), .ZN(n13147) );
  NAND2_X1 U8583 ( .A1(n7093), .A2(n7091), .ZN(n13153) );
  AND2_X1 U8584 ( .A1(n13154), .A2(n7092), .ZN(n7091) );
  AND2_X1 U8585 ( .A1(n7093), .A2(n7092), .ZN(n13155) );
  NAND2_X1 U8586 ( .A1(n10420), .A2(n10419), .ZN(n10506) );
  NAND2_X1 U8587 ( .A1(n13104), .A2(n11955), .ZN(n13164) );
  NAND2_X1 U8588 ( .A1(n8099), .A2(n8098), .ZN(n13487) );
  AND2_X1 U8589 ( .A1(n10119), .A2(n8282), .ZN(n13166) );
  OR2_X1 U8590 ( .A1(n6473), .A2(n7520), .ZN(n7521) );
  OR2_X1 U8591 ( .A1(n8068), .A2(n7519), .ZN(n7524) );
  NAND2_X1 U8592 ( .A1(n7592), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7458) );
  XNOR2_X1 U8593 ( .A(n7506), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9903) );
  OAI21_X1 U8594 ( .B1(n10030), .B2(n9856), .A(n9855), .ZN(n9978) );
  XNOR2_X1 U8595 ( .A(n13247), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n13254) );
  INV_X1 U8596 ( .A(n13254), .ZN(n13256) );
  INV_X1 U8597 ( .A(n13269), .ZN(n13469) );
  AND2_X1 U8598 ( .A1(n7074), .A2(n7073), .ZN(n13330) );
  OR2_X1 U8599 ( .A1(n13343), .A2(n13342), .ZN(n13499) );
  NAND2_X1 U8600 ( .A1(n13366), .A2(n12005), .ZN(n13341) );
  NAND2_X1 U8601 ( .A1(n8065), .A2(n8064), .ZN(n13496) );
  NAND2_X1 U8602 ( .A1(n8043), .A2(n8042), .ZN(n13505) );
  NAND2_X1 U8603 ( .A1(n8023), .A2(n8022), .ZN(n13511) );
  NAND2_X1 U8604 ( .A1(n6991), .A2(n6992), .ZN(n13396) );
  OR2_X1 U8605 ( .A1(n13407), .A2(n11984), .ZN(n6991) );
  NAND2_X1 U8606 ( .A1(n13445), .A2(n11998), .ZN(n13421) );
  NAND2_X1 U8607 ( .A1(n7902), .A2(n7901), .ZN(n13537) );
  NAND2_X1 U8608 ( .A1(n11842), .A2(n11841), .ZN(n11976) );
  NAND2_X1 U8609 ( .A1(n11786), .A2(n7081), .ZN(n11845) );
  NAND2_X1 U8610 ( .A1(n11074), .A2(n7060), .ZN(n7056) );
  NAND2_X1 U8611 ( .A1(n7785), .A2(n7784), .ZN(n11290) );
  NAND2_X1 U8612 ( .A1(n11074), .A2(n11073), .ZN(n11180) );
  INV_X1 U8613 ( .A(n14808), .ZN(n10570) );
  INV_X1 U8614 ( .A(n13455), .ZN(n13391) );
  AOI21_X1 U8615 ( .B1(n7557), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n6955), .ZN(
        n6954) );
  NOR2_X1 U8616 ( .A1(n9819), .A2(n14681), .ZN(n6955) );
  INV_X1 U8617 ( .A(n13443), .ZN(n13460) );
  NAND2_X1 U8618 ( .A1(n13482), .A2(n6668), .ZN(n13561) );
  NAND2_X1 U8619 ( .A1(n13481), .A2(n6607), .ZN(n6669) );
  AND2_X1 U8620 ( .A1(n10129), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14795) );
  INV_X1 U8621 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n7452) );
  NAND2_X1 U8622 ( .A1(n7473), .A2(n7446), .ZN(n7451) );
  NOR2_X1 U8623 ( .A1(n7448), .A2(n7445), .ZN(n7446) );
  XNOR2_X1 U8624 ( .A(n8279), .B(n8278), .ZN(n13595) );
  OAI21_X1 U8625 ( .B1(n8277), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8278) );
  INV_X1 U8626 ( .A(n10076), .ZN(n11257) );
  NAND2_X1 U8627 ( .A1(n6661), .A2(n6659), .ZN(n7486) );
  NAND2_X1 U8628 ( .A1(n6660), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6659) );
  INV_X1 U8629 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10814) );
  INV_X1 U8630 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10682) );
  INV_X1 U8631 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10535) );
  INV_X1 U8632 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10431) );
  INV_X1 U8633 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10111) );
  INV_X1 U8634 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10086) );
  INV_X1 U8635 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9762) );
  INV_X1 U8636 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9756) );
  INV_X1 U8637 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9752) );
  INV_X1 U8638 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9749) );
  INV_X1 U8639 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9743) );
  INV_X1 U8640 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9719) );
  INV_X1 U8641 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9690) );
  INV_X1 U8642 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9687) );
  INV_X1 U8643 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9676) );
  NAND2_X1 U8644 ( .A1(n11024), .A2(n11023), .ZN(n11206) );
  NAND2_X1 U8645 ( .A1(n6781), .A2(n6540), .ZN(n14409) );
  NAND2_X1 U8646 ( .A1(n6782), .A2(n6784), .ZN(n6780) );
  NAND2_X1 U8647 ( .A1(n13688), .A2(n12111), .ZN(n13602) );
  AND2_X1 U8648 ( .A1(n6799), .A2(n6501), .ZN(n11607) );
  NAND2_X1 U8649 ( .A1(n7344), .A2(n12084), .ZN(n13610) );
  NAND2_X1 U8650 ( .A1(n12151), .A2(n7331), .ZN(n7330) );
  INV_X1 U8651 ( .A(n7334), .ZN(n7331) );
  NAND2_X1 U8652 ( .A1(n7333), .A2(n12151), .ZN(n7332) );
  NAND2_X1 U8653 ( .A1(n11206), .A2(n11205), .ZN(n11207) );
  OR2_X1 U8654 ( .A1(n10021), .A2(n12042), .ZN(n10022) );
  NAND2_X1 U8655 ( .A1(n9449), .A2(n9448), .ZN(n14121) );
  AND2_X1 U8656 ( .A1(n9310), .A2(n9309), .ZN(n11816) );
  NAND2_X1 U8657 ( .A1(n14427), .A2(n6519), .ZN(n12037) );
  NAND2_X1 U8658 ( .A1(n14427), .A2(n11804), .ZN(n11806) );
  NAND2_X1 U8659 ( .A1(n13726), .A2(n12061), .ZN(n13637) );
  INV_X1 U8660 ( .A(n14152), .ZN(n13646) );
  NAND2_X1 U8661 ( .A1(n13649), .A2(n13651), .ZN(n13650) );
  NAND2_X1 U8662 ( .A1(n6787), .A2(n7340), .ZN(n13660) );
  NAND2_X1 U8663 ( .A1(n13689), .A2(n7341), .ZN(n6787) );
  NAND2_X1 U8664 ( .A1(n9493), .A2(n9492), .ZN(n14102) );
  INV_X1 U8665 ( .A(n6799), .ZN(n11600) );
  NAND2_X1 U8666 ( .A1(n13612), .A2(n12093), .ZN(n13669) );
  NAND2_X1 U8667 ( .A1(n12037), .A2(n12036), .ZN(n13679) );
  INV_X1 U8668 ( .A(n13747), .ZN(n14420) );
  INV_X1 U8669 ( .A(n10316), .ZN(n10315) );
  INV_X1 U8670 ( .A(n13672), .ZN(n14414) );
  AND2_X1 U8671 ( .A1(n6796), .A2(n12077), .ZN(n6795) );
  OAI21_X1 U8672 ( .B1(n6778), .B2(n6777), .A(n6772), .ZN(n13708) );
  INV_X1 U8673 ( .A(n6773), .ZN(n6772) );
  OAI21_X1 U8674 ( .B1(n6779), .B2(n6777), .A(n11012), .ZN(n6773) );
  NOR2_X1 U8675 ( .A1(n9642), .A2(n9641), .ZN(n9643) );
  NAND2_X1 U8676 ( .A1(n6635), .A2(n6552), .ZN(n9645) );
  AND4_X1 U8677 ( .A1(n9365), .A2(n9364), .A3(n9363), .A4(n9362), .ZN(n12057)
         );
  OR2_X1 U8678 ( .A1(n9671), .A2(n10323), .ZN(n13738) );
  NAND4_X1 U8679 ( .A1(n9189), .A2(n9188), .A3(n9187), .A4(n9186), .ZN(n13752)
         );
  INV_X1 U8680 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7462) );
  INV_X1 U8681 ( .A(n14065), .ZN(n13838) );
  INV_X1 U8682 ( .A(n14068), .ZN(n13842) );
  NAND2_X1 U8683 ( .A1(n11893), .A2(n11892), .ZN(n11894) );
  AOI21_X1 U8684 ( .B1(n6821), .B2(n14549), .A(n6818), .ZN(n14086) );
  NAND2_X1 U8685 ( .A1(n6820), .A2(n6819), .ZN(n6818) );
  OAI21_X1 U8686 ( .B1(n7218), .B2(n6822), .A(n13870), .ZN(n6821) );
  NAND2_X1 U8687 ( .A1(n13871), .A2(n14033), .ZN(n6819) );
  OAI21_X1 U8688 ( .B1(n13900), .B2(n7223), .A(n7221), .ZN(n13869) );
  NAND2_X1 U8689 ( .A1(n13899), .A2(n7415), .ZN(n13882) );
  AND2_X1 U8690 ( .A1(n7234), .A2(n7233), .ZN(n13916) );
  NAND2_X1 U8691 ( .A1(n7193), .A2(n7196), .ZN(n13939) );
  AOI21_X1 U8692 ( .B1(n13952), .B2(n13951), .A(n7200), .ZN(n13937) );
  NAND2_X1 U8693 ( .A1(n13956), .A2(n7235), .ZN(n13934) );
  INV_X1 U8694 ( .A(n14121), .ZN(n13973) );
  NAND2_X1 U8695 ( .A1(n7166), .A2(n7172), .ZN(n13997) );
  OR2_X1 U8696 ( .A1(n6517), .A2(n7174), .ZN(n7166) );
  NAND2_X1 U8697 ( .A1(n14030), .A2(n11884), .ZN(n14012) );
  NOR2_X1 U8698 ( .A1(n11716), .A2(n11715), .ZN(n11734) );
  NAND2_X1 U8699 ( .A1(n11673), .A2(n11672), .ZN(n11674) );
  NAND2_X1 U8700 ( .A1(n9288), .A2(n9287), .ZN(n14431) );
  OAI21_X1 U8701 ( .B1(n6644), .B2(n7214), .A(n7212), .ZN(n10994) );
  NAND2_X1 U8702 ( .A1(n10950), .A2(n10921), .ZN(n10995) );
  NAND2_X1 U8703 ( .A1(n14540), .A2(n10236), .ZN(n10458) );
  NAND2_X1 U8704 ( .A1(n7209), .A2(n10228), .ZN(n10464) );
  NAND2_X1 U8705 ( .A1(n14544), .A2(n10227), .ZN(n7209) );
  NOR2_X1 U8706 ( .A1(n9130), .A2(n9674), .ZN(n7192) );
  AND2_X1 U8707 ( .A1(n14576), .A2(n10495), .ZN(n14571) );
  INV_X1 U8708 ( .A(n13947), .ZN(n14558) );
  AND2_X1 U8709 ( .A1(n14576), .A2(n10487), .ZN(n14550) );
  AND2_X2 U8710 ( .A1(n10247), .A2(n13858), .ZN(n14657) );
  AND2_X1 U8711 ( .A1(n14073), .A2(n14072), .ZN(n14074) );
  AND2_X2 U8712 ( .A1(n10247), .A2(n10473), .ZN(n14646) );
  NAND2_X1 U8713 ( .A1(n7204), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9069) );
  NAND2_X1 U8714 ( .A1(n9663), .A2(n9662), .ZN(n14188) );
  NAND2_X1 U8715 ( .A1(n9088), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n9091) );
  INV_X1 U8716 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11107) );
  INV_X1 U8717 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10815) );
  INV_X1 U8718 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10683) );
  INV_X1 U8719 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10432) );
  INV_X1 U8720 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10109) );
  INV_X1 U8721 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9892) );
  INV_X1 U8722 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9764) );
  INV_X1 U8723 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9757) );
  INV_X1 U8724 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9753) );
  INV_X1 U8725 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9747) );
  INV_X1 U8726 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9744) );
  NAND2_X1 U8727 ( .A1(n7525), .A2(n6527), .ZN(n7513) );
  NAND2_X1 U8728 ( .A1(n14248), .A2(n14249), .ZN(n14310) );
  XNOR2_X1 U8729 ( .A(n14241), .B(n6643), .ZN(n15213) );
  INV_X1 U8730 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6643) );
  OAI21_X1 U8731 ( .B1(n14253), .B2(n15222), .A(n15219), .ZN(n15212) );
  INV_X1 U8732 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6971) );
  XNOR2_X1 U8733 ( .A(n14264), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15218) );
  NAND2_X1 U8734 ( .A1(n6965), .A2(n14272), .ZN(n14317) );
  AND2_X1 U8735 ( .A1(n14277), .A2(n14276), .ZN(n14319) );
  AND2_X1 U8736 ( .A1(n6964), .A2(n6963), .ZN(n14292) );
  AND2_X1 U8737 ( .A1(n11231), .A2(n8959), .ZN(n11346) );
  NAND2_X1 U8738 ( .A1(n6516), .A2(n6495), .ZN(n6700) );
  NAND2_X1 U8739 ( .A1(n14353), .A2(n7037), .ZN(n7035) );
  AND2_X1 U8740 ( .A1(n9036), .A2(n9035), .ZN(n9037) );
  NAND2_X1 U8741 ( .A1(n9034), .A2(n15016), .ZN(n9038) );
  AOI21_X1 U8742 ( .B1(n12391), .B2(n8875), .A(n8874), .ZN(n8876) );
  AND2_X1 U8743 ( .A1(n14662), .A2(n11830), .ZN(n14374) );
  NAND2_X1 U8744 ( .A1(n11917), .A2(n10203), .ZN(n10290) );
  NAND2_X1 U8745 ( .A1(n6832), .A2(n6833), .ZN(n10398) );
  INV_X1 U8746 ( .A(n12022), .ZN(n12023) );
  OAI21_X1 U8747 ( .B1(n13473), .B2(n13449), .A(n12021), .ZN(n12022) );
  AOI21_X1 U8748 ( .B1(n13470), .B2(n13455), .A(n12020), .ZN(n12021) );
  NAND2_X1 U8749 ( .A1(n14853), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6950) );
  NAND2_X1 U8750 ( .A1(n13559), .A2(n14855), .ZN(n6951) );
  NAND2_X1 U8751 ( .A1(n6893), .A2(n6892), .ZN(P2_U3496) );
  OR2_X1 U8752 ( .A1(n14835), .A2(n8149), .ZN(n6892) );
  NAND2_X1 U8753 ( .A1(n13559), .A2(n14835), .ZN(n6893) );
  XNOR2_X1 U8754 ( .A(n6792), .B(n6791), .ZN(n13601) );
  OAI21_X1 U8755 ( .B1(n14182), .B2(n14183), .A(n7323), .ZN(P1_U3325) );
  INV_X1 U8756 ( .A(n7324), .ZN(n7323) );
  INV_X1 U8757 ( .A(n14475), .ZN(n14474) );
  XNOR2_X1 U8758 ( .A(n15211), .B(n15206), .ZN(n6967) );
  NAND2_X1 U8759 ( .A1(n15019), .A2(n6969), .ZN(n6968) );
  NAND2_X1 U8760 ( .A1(n12363), .A2(n12362), .ZN(n6493) );
  AND2_X1 U8761 ( .A1(n7822), .A2(n6503), .ZN(n6494) );
  AND2_X1 U8762 ( .A1(n12368), .A2(n12369), .ZN(n6495) );
  INV_X1 U8763 ( .A(n7147), .ZN(n7146) );
  OAI21_X1 U8764 ( .B1(n8523), .B2(n7148), .A(n8309), .ZN(n7147) );
  INV_X1 U8765 ( .A(n13951), .ZN(n7199) );
  XNOR2_X1 U8766 ( .A(n12339), .B(n12503), .ZN(n12649) );
  INV_X1 U8767 ( .A(n12649), .ZN(n6897) );
  INV_X1 U8768 ( .A(n9134), .ZN(n9441) );
  INV_X1 U8769 ( .A(n10337), .ZN(n10079) );
  AND2_X1 U8770 ( .A1(n6537), .A2(n11998), .ZN(n6496) );
  AND2_X1 U8771 ( .A1(n6739), .A2(n8302), .ZN(n6497) );
  OR2_X1 U8772 ( .A1(n12053), .A2(n11732), .ZN(n6498) );
  XOR2_X1 U8773 ( .A(n7469), .B(n8285), .Z(n6499) );
  AND2_X1 U8774 ( .A1(n14388), .A2(n13188), .ZN(n6500) );
  NAND2_X1 U8775 ( .A1(n11599), .A2(n11598), .ZN(n6501) );
  NOR2_X1 U8776 ( .A1(n7255), .A2(n7254), .ZN(n6502) );
  OR2_X1 U8777 ( .A1(n7299), .A2(n7301), .ZN(n6503) );
  AND3_X1 U8778 ( .A1(n6468), .A2(n7438), .A3(n6842), .ZN(n6504) );
  INV_X1 U8779 ( .A(n13996), .ZN(n7168) );
  AND2_X1 U8780 ( .A1(n9423), .A2(n11885), .ZN(n13996) );
  NOR2_X1 U8781 ( .A1(n7360), .A2(n7361), .ZN(n6505) );
  NAND2_X1 U8782 ( .A1(n14015), .A2(n6553), .ZN(n6506) );
  AND2_X1 U8783 ( .A1(n9001), .A2(n12651), .ZN(n6507) );
  NOR2_X1 U8784 ( .A1(n8057), .A2(n8056), .ZN(n7363) );
  NOR2_X1 U8785 ( .A1(n7758), .A2(n7757), .ZN(n6508) );
  AND2_X1 U8786 ( .A1(n10512), .A2(n10511), .ZN(n6509) );
  OAI21_X1 U8787 ( .B1(n12997), .B2(n12632), .A(n12185), .ZN(n12356) );
  INV_X1 U8788 ( .A(n12356), .ZN(n6755) );
  AND2_X1 U8789 ( .A1(n6564), .A2(n7000), .ZN(n6510) );
  AND2_X1 U8790 ( .A1(n10863), .A2(n10855), .ZN(n6511) );
  AND2_X1 U8791 ( .A1(n7345), .A2(n6800), .ZN(n6512) );
  INV_X1 U8792 ( .A(n12677), .ZN(n6704) );
  NAND2_X1 U8793 ( .A1(n14190), .A2(n9733), .ZN(n13963) );
  AND3_X1 U8794 ( .A1(n8715), .A2(n8714), .A3(n8713), .ZN(n12728) );
  AND2_X1 U8795 ( .A1(n14353), .A2(n6629), .ZN(n6513) );
  AND2_X1 U8796 ( .A1(n12368), .A2(n12195), .ZN(n6514) );
  INV_X1 U8797 ( .A(n14554), .ZN(n6937) );
  OR2_X1 U8798 ( .A1(n11938), .A2(n11937), .ZN(n6515) );
  OR2_X1 U8799 ( .A1(n6701), .A2(n12369), .ZN(n6516) );
  INV_X1 U8800 ( .A(n10223), .ZN(n10233) );
  INV_X1 U8801 ( .A(n14047), .ZN(n14049) );
  INV_X1 U8802 ( .A(n13362), .ZN(n6976) );
  NAND2_X1 U8803 ( .A1(n7439), .A2(n7438), .ZN(n7587) );
  NOR2_X1 U8804 ( .A1(n6817), .A2(n6816), .ZN(n6517) );
  OR2_X1 U8805 ( .A1(n6936), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n6518) );
  AND2_X1 U8806 ( .A1(n11808), .A2(n11804), .ZN(n6519) );
  INV_X1 U8807 ( .A(n12151), .ZN(n7337) );
  NAND2_X1 U8808 ( .A1(n11460), .A2(n11459), .ZN(n6520) );
  AND2_X1 U8809 ( .A1(n7673), .A2(n7672), .ZN(n6521) );
  NAND2_X1 U8810 ( .A1(n7253), .A2(n7257), .ZN(n7256) );
  OR2_X1 U8811 ( .A1(n14288), .A2(n14287), .ZN(n6522) );
  NOR2_X1 U8812 ( .A1(n13034), .A2(n12792), .ZN(n6523) );
  AND2_X1 U8813 ( .A1(n13958), .A2(n6943), .ZN(n6524) );
  AND2_X1 U8814 ( .A1(n7460), .A2(n7457), .ZN(n6525) );
  NAND2_X1 U8815 ( .A1(n12131), .A2(n12130), .ZN(n13718) );
  AND2_X1 U8816 ( .A1(n8351), .A2(n7276), .ZN(n6526) );
  NAND2_X1 U8817 ( .A1(n13957), .A2(n7199), .ZN(n13956) );
  OR2_X1 U8818 ( .A1(n7509), .A2(SI_1_), .ZN(n6527) );
  INV_X1 U8819 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n14196) );
  INV_X1 U8820 ( .A(n6902), .ZN(n6901) );
  NAND2_X1 U8821 ( .A1(n6905), .A2(n6903), .ZN(n6902) );
  NAND2_X1 U8822 ( .A1(n8085), .A2(n8084), .ZN(n13335) );
  INV_X1 U8823 ( .A(n13851), .ZN(n7184) );
  OR2_X1 U8824 ( .A1(n15018), .A2(n15017), .ZN(n6528) );
  OR2_X1 U8825 ( .A1(n13133), .A2(n13180), .ZN(n6529) );
  AND2_X1 U8826 ( .A1(n14015), .A2(n7117), .ZN(n6530) );
  INV_X1 U8827 ( .A(n11905), .ZN(n7218) );
  NAND2_X1 U8828 ( .A1(n13667), .A2(n12100), .ZN(n13618) );
  INV_X1 U8829 ( .A(n9495), .ZN(n7125) );
  OR2_X1 U8830 ( .A1(n11904), .A2(n13920), .ZN(n6531) );
  OR2_X1 U8831 ( .A1(n14330), .A2(n12599), .ZN(n6532) );
  NAND2_X1 U8832 ( .A1(n13312), .A2(n12007), .ZN(n6533) );
  AND2_X1 U8833 ( .A1(n7194), .A2(n13918), .ZN(n6534) );
  AND2_X1 U8834 ( .A1(n7096), .A2(n14382), .ZN(n6535) );
  AND2_X1 U8835 ( .A1(n6862), .A2(n8824), .ZN(n6536) );
  OR2_X1 U8836 ( .A1(n13528), .A2(n13185), .ZN(n6537) );
  NAND2_X1 U8837 ( .A1(n13356), .A2(n6948), .ZN(n6538) );
  NAND2_X1 U8838 ( .A1(n8416), .A2(n7277), .ZN(n8427) );
  NOR2_X1 U8839 ( .A1(n13518), .A2(n13143), .ZN(n6539) );
  INV_X1 U8840 ( .A(n7317), .ZN(n7316) );
  OAI21_X1 U8841 ( .B1(n7919), .B2(n7318), .A(n7968), .ZN(n7317) );
  AND2_X1 U8842 ( .A1(n12049), .A2(n6780), .ZN(n6540) );
  NOR2_X1 U8843 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n7491) );
  INV_X1 U8844 ( .A(n8302), .ZN(n7135) );
  AND2_X1 U8845 ( .A1(n13518), .A2(n13143), .ZN(n6541) );
  NAND2_X1 U8846 ( .A1(n7583), .A2(SI_4_), .ZN(n7611) );
  AND2_X1 U8847 ( .A1(n7447), .A2(n7448), .ZN(n6542) );
  NAND2_X1 U8848 ( .A1(n8180), .A2(n8179), .ZN(n13304) );
  INV_X1 U8849 ( .A(n13304), .ZN(n13483) );
  AND2_X1 U8850 ( .A1(n8235), .A2(n8234), .ZN(n6543) );
  INV_X1 U8851 ( .A(n12053), .ZN(n14439) );
  NAND2_X1 U8852 ( .A1(n9355), .A2(n9354), .ZN(n12053) );
  INV_X1 U8853 ( .A(n7489), .ZN(n6840) );
  AND2_X1 U8854 ( .A1(n13590), .A2(n9903), .ZN(n6544) );
  INV_X1 U8855 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7448) );
  AND2_X1 U8856 ( .A1(n6664), .A2(n6663), .ZN(n6545) );
  NAND2_X1 U8857 ( .A1(n8899), .A2(n8898), .ZN(n12380) );
  AND2_X1 U8858 ( .A1(n12315), .A2(n12314), .ZN(n6546) );
  AND2_X1 U8859 ( .A1(n9173), .A2(n9171), .ZN(n6547) );
  AND2_X1 U8860 ( .A1(n7439), .A2(n6841), .ZN(n6548) );
  AND2_X1 U8861 ( .A1(n7270), .A2(n7268), .ZN(n6549) );
  AND2_X1 U8862 ( .A1(n7259), .A2(n8970), .ZN(n6550) );
  AND2_X1 U8863 ( .A1(n12089), .A2(n12084), .ZN(n6551) );
  INV_X1 U8864 ( .A(n11884), .ZN(n7177) );
  NOR2_X1 U8865 ( .A1(n9628), .A2(n9625), .ZN(n6552) );
  OR2_X1 U8866 ( .A1(n9399), .A2(n7118), .ZN(n6553) );
  AND2_X1 U8867 ( .A1(n13973), .A2(n13953), .ZN(n6554) );
  AND2_X1 U8868 ( .A1(n12117), .A2(n12116), .ZN(n6555) );
  INV_X1 U8869 ( .A(n7197), .ZN(n7196) );
  NOR2_X1 U8870 ( .A1(n13936), .A2(n7202), .ZN(n7197) );
  NAND2_X1 U8871 ( .A1(n7935), .A2(n7936), .ZN(n6556) );
  NAND2_X1 U8872 ( .A1(n11174), .A2(n8792), .ZN(n6923) );
  AND2_X1 U8873 ( .A1(n12123), .A2(n12122), .ZN(n6557) );
  INV_X1 U8874 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8843) );
  NAND2_X1 U8875 ( .A1(n12740), .A2(n12741), .ZN(n6558) );
  AND2_X1 U8876 ( .A1(n6516), .A2(n12368), .ZN(n6559) );
  NOR2_X1 U8877 ( .A1(n10887), .A2(n10886), .ZN(n6560) );
  NAND2_X1 U8878 ( .A1(n8500), .A2(n8306), .ZN(n8524) );
  NAND2_X1 U8879 ( .A1(n12014), .A2(n13176), .ZN(n6561) );
  INV_X1 U8880 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8355) );
  AND2_X1 U8881 ( .A1(n7183), .A2(n7182), .ZN(n6562) );
  INV_X1 U8882 ( .A(n7202), .ZN(n7200) );
  NAND2_X1 U8883 ( .A1(n8136), .A2(n8135), .ZN(n13263) );
  INV_X1 U8884 ( .A(n13263), .ZN(n8141) );
  OR2_X1 U8885 ( .A1(n9452), .A2(n9450), .ZN(n6563) );
  INV_X1 U8886 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7352) );
  OR2_X1 U8887 ( .A1(n13537), .A2(n11974), .ZN(n6564) );
  AND2_X1 U8888 ( .A1(n14377), .A2(n11779), .ZN(n6565) );
  AND2_X1 U8889 ( .A1(n7802), .A2(n9724), .ZN(n6566) );
  AND2_X1 U8890 ( .A1(n11833), .A2(n11832), .ZN(n6567) );
  AND2_X1 U8891 ( .A1(n7779), .A2(n15202), .ZN(n6568) );
  AND2_X1 U8892 ( .A1(n7917), .A2(n7916), .ZN(n6569) );
  INV_X1 U8893 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9074) );
  AND2_X1 U8894 ( .A1(n9892), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U8895 ( .A1(n9388), .A2(n7352), .ZN(n7351) );
  INV_X1 U8896 ( .A(n11906), .ZN(n7190) );
  INV_X1 U8897 ( .A(n11882), .ZN(n6816) );
  OAI21_X1 U8898 ( .B1(n7136), .B2(n7135), .A(n8488), .ZN(n7134) );
  AND2_X1 U8899 ( .A1(n7239), .A2(n7236), .ZN(n6571) );
  AND2_X1 U8900 ( .A1(n8231), .A2(n8230), .ZN(n6572) );
  AND2_X1 U8901 ( .A1(n7299), .A2(n7301), .ZN(n6573) );
  INV_X1 U8902 ( .A(n10229), .ZN(n14564) );
  INV_X1 U8903 ( .A(n7297), .ZN(n7296) );
  NAND2_X1 U8904 ( .A1(n7298), .A2(n7759), .ZN(n7297) );
  INV_X1 U8905 ( .A(n7415), .ZN(n7226) );
  NOR2_X1 U8906 ( .A1(n13483), .A2(n12009), .ZN(n6574) );
  AND2_X1 U8907 ( .A1(n7368), .A2(n7367), .ZN(n6575) );
  INV_X1 U8908 ( .A(n7010), .ZN(n7009) );
  NAND2_X1 U8909 ( .A1(n7012), .A2(n7011), .ZN(n7010) );
  AND2_X1 U8910 ( .A1(n12306), .A2(n12313), .ZN(n12789) );
  NAND2_X1 U8911 ( .A1(n12322), .A2(n12743), .ZN(n6576) );
  AND2_X1 U8912 ( .A1(n12145), .A2(n12144), .ZN(n6577) );
  NAND2_X1 U8913 ( .A1(n12319), .A2(n12318), .ZN(n6578) );
  AND2_X1 U8914 ( .A1(n11985), .A2(n12003), .ZN(n6579) );
  NAND2_X1 U8915 ( .A1(n8992), .A2(n8991), .ZN(n12440) );
  INV_X1 U8916 ( .A(n12440), .ZN(n7254) );
  AND4_X1 U8917 ( .A1(n6915), .A2(n10351), .A3(n8406), .A4(n6916), .ZN(n6580)
         );
  OR2_X1 U8918 ( .A1(n14084), .A2(n13740), .ZN(n6581) );
  NAND2_X1 U8919 ( .A1(n13011), .A2(n12665), .ZN(n6582) );
  AND2_X1 U8920 ( .A1(n6520), .A2(n11023), .ZN(n6583) );
  AND2_X1 U8921 ( .A1(n7693), .A2(n7692), .ZN(n6584) );
  OR2_X1 U8922 ( .A1(n7775), .A2(n7777), .ZN(n6585) );
  NOR2_X1 U8923 ( .A1(n13546), .A2(n11659), .ZN(n6586) );
  INV_X1 U8924 ( .A(n7727), .ZN(n7380) );
  AND2_X1 U8925 ( .A1(n11168), .A2(n10238), .ZN(n10016) );
  AOI22_X1 U8926 ( .A1(n7360), .A2(n7366), .B1(n7361), .B2(n7364), .ZN(n7359)
         );
  AND2_X1 U8927 ( .A1(n7244), .A2(n6498), .ZN(n6587) );
  AND2_X1 U8928 ( .A1(n8257), .A2(n8174), .ZN(n6588) );
  INV_X1 U8929 ( .A(n10236), .ZN(n7165) );
  AND2_X1 U8930 ( .A1(n11657), .A2(n11975), .ZN(n6589) );
  NAND2_X1 U8931 ( .A1(n11932), .A2(n11931), .ZN(n6590) );
  AND2_X1 U8932 ( .A1(n13915), .A2(n7233), .ZN(n6591) );
  AND2_X1 U8933 ( .A1(n12997), .A2(n12632), .ZN(n12357) );
  INV_X1 U8934 ( .A(n12357), .ZN(n12190) );
  OR2_X1 U8935 ( .A1(n9525), .A2(n9523), .ZN(n6592) );
  OR2_X1 U8936 ( .A1(n9264), .A2(n9262), .ZN(n6593) );
  OR2_X1 U8937 ( .A1(n9560), .A2(n9562), .ZN(n6594) );
  AND2_X1 U8938 ( .A1(n7337), .A2(n7334), .ZN(n6595) );
  AND2_X1 U8939 ( .A1(n9140), .A2(n9141), .ZN(n6596) );
  OR2_X1 U8940 ( .A1(n7818), .A2(n7819), .ZN(n6597) );
  OR2_X1 U8941 ( .A1(n7395), .A2(n7776), .ZN(n6598) );
  OR2_X1 U8942 ( .A1(n9494), .A2(n7125), .ZN(n6599) );
  OR2_X1 U8943 ( .A1(n7378), .A2(n7377), .ZN(n6600) );
  AND2_X1 U8944 ( .A1(n7009), .A2(n11990), .ZN(n6601) );
  OR2_X1 U8945 ( .A1(n7398), .A2(n6608), .ZN(n6602) );
  AND2_X1 U8946 ( .A1(n13072), .A2(n7107), .ZN(n7106) );
  AND2_X1 U8947 ( .A1(n7082), .A2(n11942), .ZN(n6603) );
  INV_X1 U8948 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6660) );
  INV_X1 U8949 ( .A(n8968), .ZN(n7263) );
  INV_X1 U8950 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7438) );
  INV_X1 U8951 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8285) );
  INV_X1 U8952 ( .A(n12508), .ZN(n12792) );
  NAND2_X1 U8953 ( .A1(n14383), .A2(n6535), .ZN(n7093) );
  AND2_X1 U8954 ( .A1(n7160), .A2(n8315), .ZN(n6604) );
  OAI21_X1 U8955 ( .B1(n14427), .B2(n6784), .A(n6782), .ZN(n13678) );
  OR2_X1 U8956 ( .A1(n11247), .A2(n11248), .ZN(n11829) );
  AND4_X1 U8957 ( .A1(n9305), .A2(n9304), .A3(n9303), .A4(n9302), .ZN(n14421)
         );
  AND2_X1 U8958 ( .A1(n12178), .A2(n8782), .ZN(n12384) );
  INV_X1 U8959 ( .A(n12384), .ZN(n7132) );
  NAND2_X1 U8960 ( .A1(n6859), .A2(n8807), .ZN(n12860) );
  INV_X1 U8961 ( .A(n6940), .ZN(n14038) );
  INV_X1 U8962 ( .A(n11428), .ZN(n14919) );
  NOR2_X1 U8963 ( .A1(n8617), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U8964 ( .A1(n13638), .A2(n12070), .ZN(n13649) );
  AND2_X1 U8965 ( .A1(n11739), .A2(n11738), .ZN(n6605) );
  AND3_X1 U8966 ( .A1(n12721), .A2(n12728), .A3(n12346), .ZN(n6606) );
  OR2_X1 U8967 ( .A1(n13483), .A2(n14837), .ZN(n6607) );
  AND2_X1 U8968 ( .A1(n7985), .A2(n7984), .ZN(n6608) );
  NOR2_X1 U8969 ( .A1(n12525), .A2(n12526), .ZN(n6609) );
  NOR2_X1 U8970 ( .A1(n11633), .A2(n12263), .ZN(n6610) );
  NOR2_X1 U8971 ( .A1(n13440), .A2(n13532), .ZN(n6958) );
  INV_X1 U8972 ( .A(n7133), .ZN(n12375) );
  INV_X1 U8973 ( .A(n6939), .ZN(n14002) );
  NOR2_X1 U8974 ( .A1(n14003), .A2(n14136), .ZN(n6939) );
  INV_X1 U8975 ( .A(n12875), .ZN(n8969) );
  AND4_X1 U8976 ( .A1(n8574), .A2(n8573), .A3(n8572), .A4(n8571), .ZN(n12875)
         );
  AND2_X1 U8977 ( .A1(n13052), .A2(n12875), .ZN(n6611) );
  INV_X1 U8978 ( .A(SI_14_), .ZN(n7301) );
  AND2_X1 U8979 ( .A1(n12441), .A2(n8999), .ZN(n6612) );
  INV_X1 U8980 ( .A(n12391), .ZN(n13007) );
  NAND2_X1 U8981 ( .A1(n8364), .A2(n8363), .ZN(n12391) );
  AND2_X1 U8982 ( .A1(n7021), .A2(n7020), .ZN(n6613) );
  AND2_X1 U8983 ( .A1(n8310), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n6614) );
  AND2_X1 U8984 ( .A1(n6999), .A2(n6510), .ZN(n6615) );
  AND2_X1 U8985 ( .A1(n6745), .A2(n6743), .ZN(n6616) );
  NOR2_X1 U8986 ( .A1(n7139), .A2(n7143), .ZN(n7138) );
  AND2_X1 U8987 ( .A1(n11786), .A2(n11647), .ZN(n6617) );
  AND2_X1 U8988 ( .A1(n7423), .A2(n7424), .ZN(n6618) );
  INV_X1 U8989 ( .A(n11645), .ZN(n7079) );
  XNOR2_X1 U8990 ( .A(n14815), .B(n13198), .ZN(n7063) );
  NAND2_X1 U8991 ( .A1(n7056), .A2(n11178), .ZN(n11296) );
  NAND2_X1 U8992 ( .A1(n10652), .A2(n10651), .ZN(n10767) );
  NAND2_X1 U8993 ( .A1(n11110), .A2(n11109), .ZN(n11311) );
  NAND2_X1 U8994 ( .A1(n6982), .A2(n10730), .ZN(n10889) );
  AND2_X1 U8995 ( .A1(n6653), .A2(n7154), .ZN(n6619) );
  NOR2_X1 U8996 ( .A1(n11619), .A2(n8966), .ZN(n6620) );
  INV_X1 U8997 ( .A(n10636), .ZN(n6779) );
  INV_X1 U8998 ( .A(n12312), .ZN(n12346) );
  NAND2_X1 U8999 ( .A1(n12367), .A2(n12221), .ZN(n12312) );
  OR2_X1 U9000 ( .A1(n8175), .A2(SI_27_), .ZN(n6621) );
  AND2_X1 U9001 ( .A1(n11206), .A2(n7348), .ZN(n6622) );
  NAND2_X1 U9002 ( .A1(n8720), .A2(n8719), .ZN(n6623) );
  AND2_X1 U9003 ( .A1(n8129), .A2(n11869), .ZN(n6624) );
  AND2_X1 U9004 ( .A1(n6778), .A2(n6779), .ZN(n6625) );
  NAND2_X1 U9005 ( .A1(n7472), .A2(n7473), .ZN(n8281) );
  INV_X1 U9006 ( .A(n8209), .ZN(n7307) );
  AND2_X2 U9007 ( .A1(n10139), .A2(n10128), .ZN(n14855) );
  INV_X1 U9008 ( .A(n6471), .ZN(n10064) );
  INV_X1 U9009 ( .A(n12617), .ZN(n12598) );
  INV_X1 U9010 ( .A(n10843), .ZN(n6956) );
  OR2_X1 U9011 ( .A1(n10643), .A2(n10642), .ZN(n6626) );
  INV_X1 U9012 ( .A(n14553), .ZN(n6938) );
  NOR2_X1 U9013 ( .A1(n14893), .A2(n11384), .ZN(n6627) );
  INV_X1 U9014 ( .A(n14330), .ZN(n12618) );
  AND2_X1 U9015 ( .A1(n14330), .A2(n6768), .ZN(n6628) );
  OR2_X1 U9016 ( .A1(n7036), .A2(n7038), .ZN(n6629) );
  AND2_X1 U9017 ( .A1(n13594), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6630) );
  INV_X1 U9018 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n6678) );
  INV_X1 U9019 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n6680) );
  INV_X1 U9020 ( .A(SI_24_), .ZN(n7155) );
  INV_X1 U9021 ( .A(n14342), .ZN(n12614) );
  OR2_X1 U9022 ( .A1(n10386), .A2(n10829), .ZN(n6631) );
  INV_X1 U9023 ( .A(n13761), .ZN(n7237) );
  AND2_X1 U9024 ( .A1(n8403), .A2(n8396), .ZN(n6632) );
  INV_X1 U9025 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6743) );
  INV_X1 U9026 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6975) );
  INV_X1 U9027 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6649) );
  AND2_X1 U9028 ( .A1(n14141), .A2(n14034), .ZN(n7228) );
  AOI21_X2 U9029 ( .B1(n14294), .B2(n14293), .A(n14469), .ZN(n14298) );
  NOR2_X1 U9030 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n14319), .ZN(n14278) );
  OAI21_X1 U9031 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n14299), .A(n14322), .ZN(
        n15018) );
  XNOR2_X1 U9032 ( .A(n14260), .B(n6971), .ZN(n14313) );
  NAND2_X1 U9033 ( .A1(n14476), .A2(n14477), .ZN(n14473) );
  NAND2_X1 U9034 ( .A1(n6671), .A2(n14315), .ZN(n14277) );
  XNOR2_X1 U9035 ( .A(n14270), .B(n6966), .ZN(n14314) );
  NAND2_X1 U9036 ( .A1(n15019), .A2(n6528), .ZN(n6670) );
  NAND2_X1 U9037 ( .A1(n14298), .A2(n14297), .ZN(n14476) );
  NAND2_X1 U9038 ( .A1(n14313), .A2(n14312), .ZN(n6970) );
  NAND2_X1 U9039 ( .A1(n14473), .A2(n14475), .ZN(n14324) );
  NAND2_X1 U9040 ( .A1(n14314), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n6965) );
  NAND2_X1 U9041 ( .A1(n14239), .A2(n14240), .ZN(n6962) );
  NOR2_X1 U9042 ( .A1(n14471), .A2(n14470), .ZN(n14469) );
  OAI21_X1 U9043 ( .B1(n14467), .B2(n14466), .A(P2_ADDR_REG_14__SCAN_IN), .ZN(
        n6690) );
  XNOR2_X1 U9044 ( .A(n14282), .B(n14281), .ZN(n14458) );
  NAND2_X1 U9045 ( .A1(n7207), .A2(n6633), .ZN(n10465) );
  NAND3_X1 U9046 ( .A1(n14544), .A2(n10462), .A3(n10227), .ZN(n6633) );
  NAND2_X1 U9047 ( .A1(n11367), .A2(n11366), .ZN(n11369) );
  NAND2_X1 U9048 ( .A1(n10933), .A2(n10920), .ZN(n10951) );
  NAND2_X1 U9049 ( .A1(n14000), .A2(n11901), .ZN(n13983) );
  OAI21_X1 U9050 ( .B1(n13900), .B2(n7219), .A(n7216), .ZN(n7215) );
  AND3_X2 U9051 ( .A1(n9139), .A2(n9138), .A3(n6596), .ZN(n7406) );
  NAND2_X1 U9052 ( .A1(n9468), .A2(n7418), .ZN(n9480) );
  INV_X1 U9053 ( .A(n9598), .ZN(n6635) );
  INV_X1 U9054 ( .A(n9274), .ZN(n6637) );
  NAND2_X1 U9055 ( .A1(n6674), .A2(n6672), .ZN(n9147) );
  OAI21_X1 U9056 ( .B1(n6686), .B2(n6685), .A(n7119), .ZN(n9467) );
  NAND2_X1 U9057 ( .A1(n9372), .A2(n7408), .ZN(n9385) );
  NAND2_X1 U9058 ( .A1(n6637), .A2(n6636), .ZN(n9294) );
  OAI21_X1 U9059 ( .B1(n9385), .B2(n9384), .A(n9383), .ZN(n9387) );
  NAND2_X1 U9060 ( .A1(n9229), .A2(n9228), .ZN(n9243) );
  INV_X1 U9061 ( .A(n10014), .ZN(n13755) );
  NAND2_X1 U9062 ( .A1(n6646), .A2(n6645), .ZN(n9484) );
  NAND2_X1 U9063 ( .A1(n7123), .A2(n7124), .ZN(n9507) );
  NAND2_X1 U9064 ( .A1(n6652), .A2(n7120), .ZN(n9539) );
  NAND2_X1 U9065 ( .A1(n9206), .A2(n9205), .ZN(n9223) );
  AOI21_X1 U9066 ( .B1(n9298), .B2(n9297), .A(n9296), .ZN(n9311) );
  NAND2_X1 U9067 ( .A1(n9507), .A2(n9508), .ZN(n9506) );
  NAND2_X1 U9068 ( .A1(n9539), .A2(n9540), .ZN(n9538) );
  OR2_X2 U9069 ( .A1(n9080), .A2(n11865), .ZN(n9134) );
  AOI21_X1 U9070 ( .B1(n7286), .B2(n7676), .A(n7699), .ZN(n7285) );
  NAND2_X4 U9071 ( .A1(n9405), .A2(n9404), .ZN(n14141) );
  NAND2_X1 U9072 ( .A1(n13952), .A2(n7198), .ZN(n7195) );
  INV_X1 U9073 ( .A(n7067), .ZN(n7066) );
  NAND2_X1 U9074 ( .A1(n6951), .A2(n6950), .ZN(P2_U3528) );
  NAND2_X1 U9075 ( .A1(n13284), .A2(n13283), .ZN(n13282) );
  XNOR2_X1 U9076 ( .A(n14239), .B(n14240), .ZN(n14241) );
  NAND2_X1 U9077 ( .A1(n14243), .A2(n14242), .ZN(n14195) );
  NAND2_X1 U9078 ( .A1(n14465), .A2(n6690), .ZN(n14471) );
  XNOR2_X1 U9079 ( .A(n6968), .B(n6967), .ZN(SUB_1596_U4) );
  NOR2_X2 U9080 ( .A1(n11735), .A2(n11741), .ZN(n11896) );
  OAI21_X1 U9081 ( .B1(n10463), .B2(n7208), .A(n10462), .ZN(n7207) );
  NAND2_X1 U9082 ( .A1(n13126), .A2(n13125), .ZN(n13124) );
  NOR2_X1 U9083 ( .A1(n13851), .A2(n7181), .ZN(n7180) );
  NAND2_X1 U9084 ( .A1(n6603), .A2(n6648), .ZN(n11944) );
  NAND2_X1 U9085 ( .A1(n13091), .A2(n7085), .ZN(n6648) );
  NAND3_X1 U9086 ( .A1(n9483), .A2(n9484), .A3(n6599), .ZN(n7123) );
  NAND2_X1 U9087 ( .A1(n6872), .A2(n7701), .ZN(n7705) );
  NAND3_X1 U9088 ( .A1(n9127), .A2(n9605), .A3(n9143), .ZN(n9128) );
  OR2_X1 U9089 ( .A1(n9111), .A2(n9712), .ZN(n9112) );
  NAND2_X1 U9090 ( .A1(n7528), .A2(n7527), .ZN(n7284) );
  NAND2_X1 U9091 ( .A1(n7612), .A2(n6824), .ZN(n6823) );
  INV_X1 U9092 ( .A(n6673), .ZN(n6672) );
  NAND3_X1 U9093 ( .A1(n6651), .A2(n6650), .A3(n6594), .ZN(n7121) );
  NAND2_X1 U9094 ( .A1(n9559), .A2(n9558), .ZN(n6650) );
  NAND2_X1 U9095 ( .A1(n9555), .A2(n9554), .ZN(n6651) );
  INV_X1 U9096 ( .A(n9370), .ZN(n6666) );
  NAND2_X1 U9097 ( .A1(n8791), .A2(n8790), .ZN(n11514) );
  NAND3_X1 U9098 ( .A1(n9182), .A2(n9181), .A3(n7126), .ZN(n6665) );
  NAND3_X1 U9099 ( .A1(n9512), .A2(n9511), .A3(n6592), .ZN(n6652) );
  NAND2_X1 U9100 ( .A1(n7274), .A2(n7275), .ZN(n8842) );
  NAND2_X2 U9101 ( .A1(n8828), .A2(n7414), .ZN(n12647) );
  NAND2_X1 U9102 ( .A1(n9126), .A2(n9125), .ZN(n6674) );
  AOI21_X2 U9103 ( .B1(n11056), .B2(n8785), .A(n8784), .ZN(n10823) );
  NAND2_X1 U9104 ( .A1(n14049), .A2(n10218), .ZN(n9606) );
  AOI211_X2 U9105 ( .C1(n8817), .C2(n6536), .A(n6860), .B(n8823), .ZN(n12707)
         );
  OAI21_X1 U9107 ( .B1(n12655), .B2(n12903), .A(n12654), .ZN(n12925) );
  OAI21_X1 U9108 ( .B1(n6545), .B2(n6654), .A(n7358), .ZN(n8117) );
  OAI21_X1 U9109 ( .B1(n8037), .B2(n8036), .A(n7359), .ZN(n6654) );
  NAND2_X1 U9110 ( .A1(n7401), .A2(n7404), .ZN(n7654) );
  NAND2_X1 U9111 ( .A1(n6658), .A2(n8269), .ZN(n7278) );
  NAND3_X1 U9112 ( .A1(n7280), .A2(n7283), .A3(n7279), .ZN(n6658) );
  INV_X2 U9113 ( .A(n7516), .ZN(n7591) );
  NAND2_X1 U9114 ( .A1(n8037), .A2(n8036), .ZN(n6664) );
  NAND2_X1 U9115 ( .A1(n6665), .A2(n7127), .ZN(n9207) );
  NAND2_X1 U9116 ( .A1(n6667), .A2(n6666), .ZN(n9372) );
  NAND2_X1 U9117 ( .A1(n9371), .A2(n11738), .ZN(n6667) );
  NAND2_X1 U9118 ( .A1(n7212), .A2(n7214), .ZN(n7210) );
  AOI21_X2 U9119 ( .B1(n7230), .B2(n7229), .A(n7228), .ZN(n14001) );
  INV_X1 U9120 ( .A(n7215), .ZN(n11907) );
  OR2_X1 U9121 ( .A1(n7635), .A2(n7634), .ZN(n7636) );
  NAND2_X1 U9122 ( .A1(n13394), .A2(n13395), .ZN(n7049) );
  INV_X1 U9123 ( .A(n6881), .ZN(n7585) );
  AOI21_X1 U9124 ( .B1(n11339), .B2(n11338), .A(n11337), .ZN(n11341) );
  NAND2_X1 U9125 ( .A1(n7074), .A2(n7069), .ZN(n13328) );
  OAI21_X1 U9126 ( .B1(n11646), .B2(n7080), .A(n7078), .ZN(n11847) );
  NAND3_X1 U9127 ( .A1(n7064), .A2(n7062), .A3(n10653), .ZN(n10655) );
  NOR2_X2 U9128 ( .A1(n14278), .A2(n14320), .ZN(n14282) );
  NAND2_X1 U9129 ( .A1(n14467), .A2(n14466), .ZN(n14465) );
  XNOR2_X1 U9130 ( .A(n6670), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  AND3_X2 U9131 ( .A1(n7203), .A2(n7205), .A3(n7206), .ZN(n9067) );
  NAND2_X2 U9132 ( .A1(n13590), .A2(n8281), .ZN(n9819) );
  XNOR2_X2 U9133 ( .A(n7475), .B(n7443), .ZN(n13590) );
  OR2_X2 U9134 ( .A1(n11330), .A2(n14670), .ZN(n11331) );
  NOR2_X4 U9135 ( .A1(n13496), .A2(n13372), .ZN(n13356) );
  NAND2_X1 U9136 ( .A1(n14001), .A2(n7168), .ZN(n14000) );
  NAND2_X1 U9137 ( .A1(n11849), .A2(n13123), .ZN(n13440) );
  INV_X1 U9138 ( .A(n6958), .ZN(n13439) );
  NAND2_X1 U9139 ( .A1(n7243), .A2(n7240), .ZN(n11735) );
  INV_X1 U9140 ( .A(n14016), .ZN(n7230) );
  NOR2_X2 U9141 ( .A1(n13413), .A2(n13518), .ZN(n13399) );
  NAND2_X1 U9142 ( .A1(n10570), .A2(n10601), .ZN(n10582) );
  NAND2_X1 U9143 ( .A1(n7234), .A2(n6591), .ZN(n13914) );
  NAND3_X1 U9144 ( .A1(n7476), .A2(n6504), .A3(n6548), .ZN(n7474) );
  NAND2_X1 U9145 ( .A1(n12820), .A2(n12300), .ZN(n12809) );
  INV_X4 U9146 ( .A(n8890), .ZN(n12173) );
  NAND2_X2 U9147 ( .A1(n12795), .A2(n8659), .ZN(n12970) );
  NAND2_X1 U9148 ( .A1(n12864), .A2(n8577), .ZN(n12851) );
  INV_X1 U9149 ( .A(n8785), .ZN(n12224) );
  NAND2_X1 U9150 ( .A1(n8596), .A2(n8595), .ZN(n12834) );
  NAND2_X1 U9151 ( .A1(n6910), .A2(n6908), .ZN(n11352) );
  NAND2_X1 U9152 ( .A1(n9544), .A2(n9543), .ZN(n9556) );
  NAND2_X1 U9153 ( .A1(n9274), .A2(n9275), .ZN(n9293) );
  OAI21_X1 U9154 ( .B1(n9143), .B2(n9605), .A(n9128), .ZN(n6673) );
  OAI21_X1 U9155 ( .B1(n8924), .B2(n8925), .A(n10748), .ZN(n8934) );
  OAI21_X2 U9156 ( .B1(n12490), .B2(n12486), .A(n12487), .ZN(n12428) );
  INV_X1 U9157 ( .A(n8464), .ZN(n6696) );
  NAND3_X1 U9158 ( .A1(n6917), .A2(n6848), .A3(n6915), .ZN(n8464) );
  NAND2_X1 U9159 ( .A1(n8989), .A2(n12745), .ZN(n12456) );
  OAI21_X1 U9160 ( .B1(n12449), .B2(n7267), .A(n7264), .ZN(n8988) );
  NOR2_X2 U9161 ( .A1(n13295), .A2(n13299), .ZN(n13294) );
  NAND2_X1 U9162 ( .A1(n7300), .A2(n7825), .ZN(n7850) );
  AOI21_X2 U9163 ( .B1(n13325), .B2(n12006), .A(n6675), .ZN(n13319) );
  OAI21_X1 U9164 ( .B1(n12690), .B2(n8826), .A(n12676), .ZN(n12662) );
  OAI21_X1 U9165 ( .B1(n12942), .B2(n12728), .A(n12705), .ZN(n12688) );
  OR2_X2 U9166 ( .A1(n12647), .A2(n12649), .ZN(n6870) );
  NAND4_X1 U9167 ( .A1(n6877), .A2(n6878), .A3(n7615), .A4(n6684), .ZN(n7631)
         );
  NAND3_X1 U9168 ( .A1(n7611), .A2(n7578), .A3(n7579), .ZN(n6684) );
  NAND2_X1 U9169 ( .A1(n13846), .A2(n11891), .ZN(n11895) );
  NAND2_X1 U9170 ( .A1(n7121), .A2(n7122), .ZN(n9598) );
  NAND3_X1 U9171 ( .A1(n9248), .A2(n9247), .A3(n6593), .ZN(n6688) );
  NAND2_X1 U9172 ( .A1(n15213), .A2(n15212), .ZN(n6689) );
  NOR2_X1 U9173 ( .A1(n14324), .A2(n14323), .ZN(n14299) );
  NAND2_X1 U9174 ( .A1(n14244), .A2(n14245), .ZN(n6974) );
  OAI21_X2 U9175 ( .B1(n12617), .B2(n12616), .A(n12615), .ZN(n12619) );
  AND3_X1 U9176 ( .A1(n6698), .A2(n6697), .A3(n6700), .ZN(P3_U3296) );
  NAND3_X1 U9177 ( .A1(n6699), .A2(n6559), .A3(n6493), .ZN(n6697) );
  NAND3_X1 U9178 ( .A1(n6699), .A2(n6514), .A3(n6493), .ZN(n6698) );
  NAND2_X1 U9179 ( .A1(n6708), .A2(n6709), .ZN(n12326) );
  NAND2_X1 U9180 ( .A1(n12311), .A2(n6710), .ZN(n6708) );
  NAND2_X1 U9181 ( .A1(n12315), .A2(n12310), .ZN(n6716) );
  INV_X1 U9182 ( .A(n12227), .ZN(n12226) );
  INV_X1 U9183 ( .A(n6719), .ZN(n6718) );
  NAND3_X1 U9184 ( .A1(n6721), .A2(n6720), .A3(n12649), .ZN(n12345) );
  NAND2_X1 U9185 ( .A1(n8579), .A2(n6604), .ZN(n6727) );
  NAND2_X1 U9186 ( .A1(n8438), .A2(n8437), .ZN(n8295) );
  NAND2_X1 U9187 ( .A1(n8426), .A2(n8291), .ZN(n6728) );
  NAND2_X1 U9188 ( .A1(n6729), .A2(n8335), .ZN(n8336) );
  INV_X1 U9189 ( .A(n8524), .ZN(n6730) );
  OAI21_X1 U9190 ( .B1(n6730), .B2(n6732), .A(n6731), .ZN(n8311) );
  NAND2_X1 U9191 ( .A1(n8451), .A2(n6497), .ZN(n6736) );
  INV_X1 U9192 ( .A(n8323), .ZN(n6742) );
  NAND2_X1 U9193 ( .A1(n6742), .A2(n7138), .ZN(n6744) );
  NAND2_X1 U9194 ( .A1(n6744), .A2(n6745), .ZN(n8328) );
  NAND2_X1 U9195 ( .A1(n8323), .A2(n8322), .ZN(n8646) );
  NAND2_X1 U9196 ( .A1(n6744), .A2(n6616), .ZN(n8329) );
  NAND2_X1 U9197 ( .A1(n8728), .A2(n8339), .ZN(n6753) );
  OAI21_X1 U9198 ( .B1(n8728), .B2(n6750), .A(n6748), .ZN(n8748) );
  NAND3_X1 U9199 ( .A1(n6757), .A2(n7025), .A3(n11378), .ZN(n11380) );
  NOR2_X1 U9200 ( .A1(n12597), .A2(n7022), .ZN(n12599) );
  NAND3_X1 U9201 ( .A1(n6766), .A2(n6763), .A3(n6765), .ZN(n6769) );
  NAND3_X1 U9202 ( .A1(n6766), .A2(n6767), .A3(n6765), .ZN(n14327) );
  INV_X1 U9203 ( .A(n6769), .ZN(n14326) );
  NAND2_X1 U9204 ( .A1(n6778), .A2(n6770), .ZN(n6776) );
  NAND2_X1 U9205 ( .A1(n14427), .A2(n6782), .ZN(n6781) );
  NAND2_X1 U9206 ( .A1(n13689), .A2(n6788), .ZN(n6786) );
  NAND2_X1 U9207 ( .A1(n6794), .A2(n6795), .ZN(n13698) );
  NAND3_X1 U9208 ( .A1(n13726), .A2(n7325), .A3(n13651), .ZN(n6794) );
  NAND2_X1 U9209 ( .A1(n7347), .A2(n6512), .ZN(n6799) );
  NAND2_X1 U9210 ( .A1(n6799), .A2(n6798), .ZN(n11800) );
  NAND2_X1 U9211 ( .A1(n7347), .A2(n7345), .ZN(n11465) );
  INV_X1 U9212 ( .A(n11464), .ZN(n6800) );
  NAND3_X1 U9213 ( .A1(n9155), .A2(n9059), .A3(n9060), .ZN(n9216) );
  NAND2_X1 U9214 ( .A1(n10924), .A2(n11109), .ZN(n6809) );
  INV_X1 U9215 ( .A(n6817), .ZN(n11883) );
  NAND2_X1 U9216 ( .A1(n6827), .A2(n10298), .ZN(n6826) );
  NAND3_X1 U9217 ( .A1(n6826), .A2(n10521), .A3(n6825), .ZN(n10527) );
  INV_X1 U9218 ( .A(n10299), .ZN(n6828) );
  NAND2_X1 U9219 ( .A1(n6832), .A2(n6831), .ZN(n10395) );
  AND2_X1 U9220 ( .A1(n10296), .A2(n6833), .ZN(n6831) );
  NAND2_X1 U9221 ( .A1(n6836), .A2(n6511), .ZN(n11245) );
  NOR2_X1 U9222 ( .A1(n7489), .A2(n7435), .ZN(n7476) );
  NAND3_X1 U9223 ( .A1(n7431), .A2(n7430), .A3(n6838), .ZN(n7489) );
  NAND4_X1 U9224 ( .A1(n6504), .A2(n6840), .A3(n6839), .A4(n6548), .ZN(n7470)
         );
  INV_X1 U9225 ( .A(n7558), .ZN(n7439) );
  AND2_X1 U9226 ( .A1(n6660), .A2(n7436), .ZN(n6842) );
  NOR2_X1 U9227 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n6844) );
  MUX2_X1 U9228 ( .A(P2_IR_REG_0__SCAN_IN), .B(n6499), .S(n9819), .Z(n10337)
         );
  NOR2_X1 U9229 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .ZN(
        n6848) );
  NAND2_X2 U9230 ( .A1(n12229), .A2(n6851), .ZN(n12202) );
  OR2_X1 U9231 ( .A1(n8922), .A2(n10798), .ZN(n8930) );
  OR2_X1 U9232 ( .A1(n8922), .A2(n10798), .ZN(n6850) );
  NAND2_X1 U9233 ( .A1(n12228), .A2(n6851), .ZN(n12231) );
  NAND2_X1 U9234 ( .A1(n10745), .A2(n6851), .ZN(n11055) );
  NAND2_X1 U9235 ( .A1(n12223), .A2(n6851), .ZN(n12225) );
  NAND2_X1 U9236 ( .A1(n6854), .A2(n6852), .ZN(n12844) );
  OR2_X2 U9237 ( .A1(n12874), .A2(n6856), .ZN(n6854) );
  AOI21_X2 U9238 ( .B1(n11514), .B2(n8801), .A(n7421), .ZN(n11685) );
  OR2_X1 U9239 ( .A1(n12647), .A2(n6868), .ZN(n6865) );
  NAND3_X1 U9240 ( .A1(n6865), .A2(n6864), .A3(n6866), .ZN(n8832) );
  NAND2_X1 U9241 ( .A1(n12647), .A2(n6869), .ZN(n6864) );
  INV_X1 U9242 ( .A(n6870), .ZN(n12646) );
  NAND2_X1 U9243 ( .A1(n6873), .A2(n7285), .ZN(n6872) );
  NAND2_X1 U9244 ( .A1(n7659), .A2(n7286), .ZN(n6873) );
  NAND3_X1 U9245 ( .A1(n6527), .A2(n7525), .A3(n7511), .ZN(n7526) );
  AND2_X1 U9246 ( .A1(n6874), .A2(SI_0_), .ZN(n7511) );
  MUX2_X1 U9247 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(P1_DATAO_REG_0__SCAN_IN), 
        .S(n7510), .Z(n6874) );
  NAND2_X1 U9248 ( .A1(n7509), .A2(SI_1_), .ZN(n7525) );
  NAND2_X1 U9249 ( .A1(n6875), .A2(n7611), .ZN(n6877) );
  NOR2_X1 U9250 ( .A1(n7582), .A2(n7580), .ZN(n6875) );
  NAND2_X1 U9251 ( .A1(n7582), .A2(n7581), .ZN(n6876) );
  NAND2_X1 U9252 ( .A1(n7584), .A2(n7611), .ZN(n6878) );
  INV_X1 U9253 ( .A(n7611), .ZN(n6879) );
  NAND2_X1 U9254 ( .A1(n7824), .A2(n6494), .ZN(n6887) );
  OR2_X1 U9255 ( .A1(n12697), .A2(n6902), .ZN(n6895) );
  NAND2_X1 U9256 ( .A1(n12697), .A2(n6906), .ZN(n6904) );
  NAND2_X1 U9257 ( .A1(n6895), .A2(n6899), .ZN(n12650) );
  NAND2_X1 U9258 ( .A1(n11216), .A2(n6912), .ZN(n6910) );
  MUX2_X1 U9259 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14191), .S(n9733), .Z(n14565)
         );
  NAND2_X2 U9260 ( .A1(n9071), .A2(n7204), .ZN(n9666) );
  OR2_X2 U9261 ( .A1(n11717), .A2(n12053), .ZN(n11742) );
  OR2_X2 U9262 ( .A1(n11678), .A2(n14411), .ZN(n11717) );
  NOR2_X2 U9263 ( .A1(n11118), .A2(n14431), .ZN(n11318) );
  OR2_X2 U9264 ( .A1(n11003), .A2(n11605), .ZN(n11118) );
  NOR2_X2 U9265 ( .A1(n10952), .A2(n11200), .ZN(n11005) );
  NOR2_X2 U9266 ( .A1(n14002), .A2(n14130), .ZN(n13986) );
  NOR2_X2 U9267 ( .A1(n14037), .A2(n14147), .ZN(n6940) );
  NAND2_X1 U9268 ( .A1(n13958), .A2(n6941), .ZN(n13894) );
  NAND2_X1 U9269 ( .A1(n13356), .A2(n6946), .ZN(n13288) );
  NOR2_X2 U9270 ( .A1(n10582), .A2(n14815), .ZN(n10769) );
  NOR2_X2 U9271 ( .A1(n10602), .A2(n14802), .ZN(n10601) );
  NOR2_X2 U9272 ( .A1(n13439), .A2(n13528), .ZN(n13411) );
  NOR2_X2 U9273 ( .A1(n10768), .A2(n10790), .ZN(n10734) );
  INV_X1 U9274 ( .A(n6964), .ZN(n14462) );
  INV_X1 U9275 ( .A(n14461), .ZN(n6963) );
  NOR2_X2 U9276 ( .A1(n14266), .A2(n14267), .ZN(n14270) );
  OAI21_X2 U9277 ( .B1(n13363), .B2(n6976), .A(n11988), .ZN(n13345) );
  NAND2_X1 U9278 ( .A1(n13203), .A2(n10337), .ZN(n10185) );
  NAND2_X1 U9279 ( .A1(n13203), .A2(n10079), .ZN(n8242) );
  NAND3_X1 U9280 ( .A1(n7516), .A2(n13203), .A3(n6977), .ZN(n7499) );
  NAND3_X2 U9281 ( .A1(n6525), .A2(n7458), .A3(n7459), .ZN(n13203) );
  OAI21_X2 U9282 ( .B1(n10728), .B2(n6979), .A(n6978), .ZN(n10891) );
  NAND2_X1 U9283 ( .A1(n6984), .A2(n6983), .ZN(n11076) );
  INV_X1 U9284 ( .A(n10891), .ZN(n6984) );
  NAND2_X1 U9285 ( .A1(n13407), .A2(n6989), .ZN(n6988) );
  NAND3_X1 U9286 ( .A1(n6995), .A2(n10659), .A3(n6993), .ZN(n10662) );
  INV_X1 U9287 ( .A(n7063), .ZN(n6994) );
  NAND2_X1 U9288 ( .A1(n10575), .A2(n6996), .ZN(n6995) );
  NAND2_X1 U9289 ( .A1(n10658), .A2(n10657), .ZN(n10774) );
  NAND2_X1 U9290 ( .A1(n6997), .A2(n7063), .ZN(n10658) );
  NAND2_X1 U9291 ( .A1(n6999), .A2(n6998), .ZN(n11980) );
  NAND2_X1 U9292 ( .A1(n11658), .A2(n6589), .ZN(n6999) );
  AND2_X1 U9293 ( .A1(n11977), .A2(n6510), .ZN(n6998) );
  NAND2_X1 U9294 ( .A1(n13295), .A2(n6601), .ZN(n7003) );
  AOI21_X1 U9295 ( .B1(n7017), .B2(n7014), .A(n6586), .ZN(n7013) );
  INV_X1 U9296 ( .A(n7018), .ZN(n7014) );
  INV_X1 U9297 ( .A(n7017), .ZN(n7015) );
  NAND2_X1 U9298 ( .A1(n7016), .A2(n7017), .ZN(n11778) );
  NAND2_X1 U9299 ( .A1(n11326), .A2(n7018), .ZN(n7016) );
  NAND2_X1 U9300 ( .A1(n10446), .A2(n10447), .ZN(n7025) );
  OR2_X1 U9301 ( .A1(n10385), .A2(n10442), .ZN(n7026) );
  NAND2_X1 U9302 ( .A1(n10385), .A2(n10442), .ZN(n10448) );
  OAI21_X1 U9303 ( .B1(n14894), .B2(n7030), .A(n7029), .ZN(n14911) );
  NAND2_X1 U9304 ( .A1(n14355), .A2(n6513), .ZN(n7034) );
  OAI211_X1 U9305 ( .C1(n14355), .C2(n7035), .A(n7034), .B(n12630), .ZN(
        P3_U3201) );
  NOR2_X1 U9306 ( .A1(n14355), .A2(n14354), .ZN(n14356) );
  NOR2_X1 U9307 ( .A1(n11481), .A2(n11480), .ZN(n11483) );
  NOR2_X1 U9308 ( .A1(n12912), .A2(n11389), .ZN(n11480) );
  NAND2_X1 U9309 ( .A1(n10550), .A2(n10549), .ZN(n10575) );
  NAND2_X1 U9310 ( .A1(n11078), .A2(n11077), .ZN(n11185) );
  OR2_X1 U9311 ( .A1(n8185), .A2(n9847), .ZN(n7505) );
  NAND2_X1 U9312 ( .A1(n10169), .A2(n10168), .ZN(n10609) );
  NOR2_X1 U9313 ( .A1(n11483), .A2(n11482), .ZN(n11536) );
  NAND2_X1 U9314 ( .A1(n11076), .A2(n11075), .ZN(n11078) );
  XNOR2_X1 U9315 ( .A(n11380), .B(n11411), .ZN(n14856) );
  NOR2_X2 U9316 ( .A1(n7587), .A2(n7442), .ZN(n7488) );
  OAI21_X1 U9317 ( .B1(n6471), .B2(n7046), .A(n10140), .ZN(n7047) );
  NAND2_X1 U9318 ( .A1(n7047), .A2(n10142), .ZN(n10157) );
  XNOR2_X1 U9319 ( .A(n7048), .B(n10068), .ZN(n10142) );
  NAND2_X1 U9320 ( .A1(n10141), .A2(n10140), .ZN(n10143) );
  NAND2_X1 U9321 ( .A1(n10064), .A2(n10185), .ZN(n10141) );
  INV_X1 U9322 ( .A(n10142), .ZN(n10162) );
  NAND2_X1 U9323 ( .A1(n7049), .A2(n6579), .ZN(n13510) );
  NAND2_X1 U9324 ( .A1(n11074), .A2(n7057), .ZN(n7055) );
  NAND2_X1 U9325 ( .A1(n7063), .A2(n10651), .ZN(n7062) );
  NAND2_X1 U9326 ( .A1(n10573), .A2(n10651), .ZN(n7064) );
  OAI21_X1 U9327 ( .B1(n13309), .B2(n7066), .A(n7065), .ZN(n13284) );
  NAND2_X1 U9328 ( .A1(n13309), .A2(n12008), .ZN(n7068) );
  NAND2_X1 U9329 ( .A1(n13366), .A2(n7071), .ZN(n7074) );
  INV_X1 U9330 ( .A(n7074), .ZN(n13342) );
  NAND2_X1 U9331 ( .A1(n13447), .A2(n6496), .ZN(n7075) );
  NAND2_X1 U9332 ( .A1(n7075), .A2(n7076), .ZN(n13406) );
  NAND2_X1 U9333 ( .A1(n10757), .A2(n7100), .ZN(n7097) );
  NAND2_X1 U9334 ( .A1(n7103), .A2(n7104), .ZN(n11967) );
  NAND2_X1 U9335 ( .A1(n13164), .A2(n7106), .ZN(n7103) );
  AND2_X1 U9336 ( .A1(n10508), .A2(n10419), .ZN(n7108) );
  NAND2_X1 U9337 ( .A1(n9401), .A2(n7115), .ZN(n7113) );
  NAND2_X1 U9338 ( .A1(n7113), .A2(n7114), .ZN(n9425) );
  NAND2_X1 U9339 ( .A1(n9450), .A2(n9452), .ZN(n7119) );
  OR2_X1 U9340 ( .A1(n9194), .A2(n9196), .ZN(n7126) );
  NAND2_X1 U9341 ( .A1(n8415), .A2(n8414), .ZN(n7129) );
  NAND2_X1 U9342 ( .A1(n7130), .A2(n8287), .ZN(n8415) );
  NAND2_X1 U9343 ( .A1(n8286), .A2(n8404), .ZN(n7130) );
  NAND2_X1 U9344 ( .A1(n8885), .A2(n8884), .ZN(n7133) );
  OAI22_X1 U9345 ( .A1(n12361), .A2(n12360), .B1(n12363), .B2(n12359), .ZN(
        n7144) );
  INV_X1 U9346 ( .A(n7162), .ZN(n7161) );
  NAND2_X1 U9347 ( .A1(n7161), .A2(n8338), .ZN(n8720) );
  NAND2_X1 U9348 ( .A1(n8338), .A2(n8337), .ZN(n8718) );
  INV_X1 U9349 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7163) );
  OAI211_X1 U9350 ( .C1(n10226), .C2(n7165), .A(n7164), .B(n10457), .ZN(n10460) );
  NAND3_X1 U9351 ( .A1(n10479), .A2(n10234), .A3(n10236), .ZN(n7164) );
  NAND2_X1 U9352 ( .A1(n11899), .A2(n14034), .ZN(n7178) );
  NAND2_X1 U9353 ( .A1(n13870), .A2(n7180), .ZN(n7179) );
  AOI21_X1 U9354 ( .B1(n9414), .B2(n13775), .A(n7192), .ZN(n7191) );
  CLKBUF_X1 U9355 ( .A(n7195), .Z(n7193) );
  NAND2_X1 U9356 ( .A1(n14115), .A2(n13622), .ZN(n7202) );
  NAND4_X1 U9357 ( .A1(n7203), .A2(n7206), .A3(n7354), .A4(n7205), .ZN(n7204)
         );
  NAND2_X1 U9358 ( .A1(n9605), .A2(n10230), .ZN(n10219) );
  NAND2_X1 U9359 ( .A1(n13755), .A2(n10220), .ZN(n9605) );
  NAND2_X1 U9360 ( .A1(n10951), .A2(n7212), .ZN(n7211) );
  NAND3_X1 U9361 ( .A1(n7211), .A2(n10923), .A3(n7210), .ZN(n10925) );
  NAND2_X1 U9362 ( .A1(n7220), .A2(n11905), .ZN(n7219) );
  NAND2_X1 U9363 ( .A1(n13956), .A2(n7231), .ZN(n7234) );
  INV_X1 U9364 ( .A(n7234), .ZN(n13933) );
  NAND2_X1 U9365 ( .A1(n9733), .A2(n7238), .ZN(n7236) );
  XNOR2_X2 U9366 ( .A(n9069), .B(n9074), .ZN(n9665) );
  NAND3_X1 U9367 ( .A1(n9666), .A2(n9665), .A3(n7237), .ZN(n7239) );
  NAND2_X1 U9368 ( .A1(n11673), .A2(n6587), .ZN(n7243) );
  NAND2_X1 U9369 ( .A1(n7246), .A2(n9033), .ZN(P3_U3154) );
  NAND2_X1 U9370 ( .A1(n7247), .A2(n12477), .ZN(n7246) );
  NAND2_X1 U9371 ( .A1(n7248), .A2(n12394), .ZN(n7247) );
  NAND2_X1 U9372 ( .A1(n9008), .A2(n9007), .ZN(n12394) );
  NAND2_X1 U9373 ( .A1(n7250), .A2(n7249), .ZN(n7248) );
  INV_X1 U9374 ( .A(n9009), .ZN(n7249) );
  NAND2_X1 U9375 ( .A1(n9008), .A2(n9006), .ZN(n7250) );
  NAND2_X1 U9376 ( .A1(n7251), .A2(n12440), .ZN(n7252) );
  NAND2_X1 U9377 ( .A1(n7255), .A2(n12440), .ZN(n9043) );
  NAND2_X1 U9378 ( .A1(n7256), .A2(n12728), .ZN(n7255) );
  INV_X1 U9379 ( .A(n8991), .ZN(n7257) );
  NAND2_X1 U9380 ( .A1(n11620), .A2(n7262), .ZN(n7261) );
  NAND3_X1 U9381 ( .A1(n8968), .A2(n11621), .A3(n7260), .ZN(n7259) );
  NAND2_X1 U9382 ( .A1(n11344), .A2(n8962), .ZN(n8964) );
  NAND2_X1 U9383 ( .A1(n7278), .A2(n8284), .ZN(P2_U3328) );
  NAND2_X1 U9384 ( .A1(n8265), .A2(n8263), .ZN(n7279) );
  OAI21_X1 U9385 ( .B1(n8265), .B2(n7282), .A(n7281), .ZN(n7280) );
  NAND3_X1 U9386 ( .A1(n7284), .A2(n7553), .A3(n7531), .ZN(n7554) );
  NAND2_X1 U9387 ( .A1(n7659), .A2(n7658), .ZN(n7678) );
  NAND2_X1 U9388 ( .A1(n7760), .A2(n7292), .ZN(n7290) );
  NAND2_X1 U9389 ( .A1(n7868), .A2(n7867), .ZN(n7870) );
  NAND2_X1 U9390 ( .A1(n8127), .A2(n7308), .ZN(n7303) );
  NAND2_X1 U9391 ( .A1(n7303), .A2(n7304), .ZN(n8134) );
  NAND2_X1 U9392 ( .A1(n8127), .A2(n8126), .ZN(n8144) );
  NAND2_X1 U9393 ( .A1(n7920), .A2(n7919), .ZN(n7315) );
  AND2_X2 U9394 ( .A1(n9081), .A2(n9080), .ZN(n9133) );
  OAI22_X1 U9395 ( .A1(n9080), .A2(P1_U3086), .B1(n14181), .B2(n14180), .ZN(
        n7324) );
  OAI211_X1 U9396 ( .C1(n13718), .C2(n7332), .A(n7328), .B(n7327), .ZN(n12158)
         );
  NAND2_X1 U9397 ( .A1(n13718), .A2(n6595), .ZN(n7327) );
  OAI21_X1 U9398 ( .B1(n7333), .B2(n7337), .A(n7329), .ZN(n7328) );
  NAND2_X1 U9399 ( .A1(n7333), .A2(n7330), .ZN(n7329) );
  NAND2_X1 U9400 ( .A1(n11024), .A2(n6583), .ZN(n7347) );
  NAND2_X1 U9401 ( .A1(n9092), .A2(n7350), .ZN(n9646) );
  INV_X1 U9402 ( .A(n9646), .ZN(n9648) );
  NAND2_X1 U9403 ( .A1(n9067), .A2(n7355), .ZN(n9078) );
  INV_X1 U9404 ( .A(n9078), .ZN(n9076) );
  INV_X1 U9405 ( .A(n8056), .ZN(n7370) );
  NAND2_X1 U9406 ( .A1(n7375), .A2(n6597), .ZN(n7843) );
  NAND3_X1 U9407 ( .A1(n7376), .A2(n6470), .A3(n6600), .ZN(n7375) );
  INV_X1 U9408 ( .A(n7799), .ZN(n7376) );
  INV_X1 U9409 ( .A(n7819), .ZN(n7377) );
  INV_X1 U9410 ( .A(n7818), .ZN(n7378) );
  NAND2_X1 U9411 ( .A1(n7748), .A2(n7749), .ZN(n7747) );
  AOI21_X1 U9412 ( .B1(n7866), .B2(n7385), .A(n7383), .ZN(n7382) );
  INV_X1 U9413 ( .A(n7382), .ZN(n7888) );
  NAND2_X1 U9414 ( .A1(n7389), .A2(n7390), .ZN(n7696) );
  NAND2_X1 U9415 ( .A1(n7675), .A2(n7391), .ZN(n7389) );
  NAND2_X1 U9416 ( .A1(n6521), .A2(n7393), .ZN(n7391) );
  NOR2_X1 U9417 ( .A1(n6521), .A2(n7393), .ZN(n7392) );
  NAND2_X1 U9418 ( .A1(n7394), .A2(n6598), .ZN(n7798) );
  NAND3_X1 U9419 ( .A1(n7753), .A2(n6585), .A3(n7752), .ZN(n7394) );
  NAND2_X1 U9420 ( .A1(n7396), .A2(n7397), .ZN(n8010) );
  NAND3_X1 U9421 ( .A1(n7965), .A2(n7964), .A3(n6602), .ZN(n7396) );
  INV_X1 U9422 ( .A(n7986), .ZN(n7398) );
  INV_X1 U9423 ( .A(n7402), .ZN(n7399) );
  NAND2_X1 U9424 ( .A1(n7629), .A2(n7404), .ZN(n7403) );
  NAND3_X1 U9425 ( .A1(n7403), .A2(n7655), .A3(n7402), .ZN(n7653) );
  NAND4_X2 U9426 ( .A1(n8402), .A2(n8401), .A3(n8400), .A4(n8399), .ZN(n12521)
         );
  NAND2_X1 U9427 ( .A1(n8313), .A2(n8312), .ZN(n8579) );
  AOI21_X1 U9428 ( .B1(n13079), .B2(n13080), .A(n7417), .ZN(n13126) );
  AND4_X2 U9429 ( .A1(n8413), .A2(n8412), .A3(n8411), .A4(n8410), .ZN(n10875)
         );
  INV_X1 U9430 ( .A(n10188), .ZN(n10186) );
  AND4_X2 U9431 ( .A1(n9116), .A2(n9119), .A3(n9117), .A4(n9118), .ZN(n14047)
         );
  OR2_X1 U9432 ( .A1(n8360), .A2(n8357), .ZN(n8358) );
  NAND2_X1 U9433 ( .A1(n9598), .A2(n9597), .ZN(n9644) );
  NAND2_X1 U9434 ( .A1(n9098), .A2(n10238), .ZN(n9102) );
  XNOR2_X1 U9435 ( .A(n8311), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8560) );
  OAI22_X1 U9436 ( .A1(n14595), .A2(n12106), .B1(n7406), .B2(n12105), .ZN(
        n10316) );
  INV_X1 U9437 ( .A(n8929), .ZN(n10872) );
  NAND2_X1 U9438 ( .A1(n9133), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9118) );
  NAND2_X1 U9439 ( .A1(n12456), .A2(n8990), .ZN(n8992) );
  NOR2_X1 U9440 ( .A1(n10309), .A2(n10020), .ZN(n10025) );
  AND2_X1 U9441 ( .A1(n10019), .A2(n10018), .ZN(n10020) );
  INV_X1 U9442 ( .A(n8185), .ZN(n8215) );
  OR2_X1 U9443 ( .A1(n8185), .A2(n9894), .ZN(n7459) );
  OR2_X1 U9444 ( .A1(n8950), .A2(n11097), .ZN(n11126) );
  XNOR2_X1 U9445 ( .A(n8935), .B(n8936), .ZN(n11154) );
  OR2_X1 U9446 ( .A1(n12192), .A2(n12191), .ZN(n12194) );
  OAI21_X2 U9447 ( .B1(n11586), .B2(n12876), .A(n11587), .ZN(n11620) );
  NAND2_X1 U9448 ( .A1(n12435), .A2(n12434), .ZN(n12433) );
  OAI222_X1 U9449 ( .A1(P3_U3151), .A2(n12601), .B1(n13067), .B2(n11617), .C1(
        n15059), .C2(n13059), .ZN(P3_U3268) );
  OAI21_X1 U9450 ( .B1(n8239), .B2(n6543), .A(n8238), .ZN(n8265) );
  INV_X1 U9451 ( .A(n7406), .ZN(n14054) );
  NOR2_X1 U9452 ( .A1(n8955), .A2(n11171), .ZN(n7407) );
  OR2_X1 U9453 ( .A1(n9604), .A2(n9585), .ZN(n7408) );
  AND2_X1 U9454 ( .A1(n9367), .A2(n9585), .ZN(n7409) );
  AND4_X1 U9455 ( .A1(n8354), .A2(n8353), .A3(n8763), .A4(n8352), .ZN(n7410)
         );
  AND2_X1 U9456 ( .A1(n10628), .A2(n10627), .ZN(n7411) );
  AND2_X1 U9457 ( .A1(n6588), .A2(n8199), .ZN(n7412) );
  OR2_X1 U9458 ( .A1(n11904), .A2(n13720), .ZN(n7415) );
  INV_X1 U9459 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7445) );
  AND2_X2 U9460 ( .A1(n8872), .A2(n8871), .ZN(n15016) );
  NAND2_X1 U9461 ( .A1(n11152), .A2(n8947), .ZN(n7416) );
  AND2_X1 U9462 ( .A1(n11947), .A2(n11946), .ZN(n7417) );
  INV_X1 U9463 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9075) );
  INV_X1 U9464 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7477) );
  AND2_X1 U9465 ( .A1(n7831), .A2(n7830), .ZN(n7419) );
  OAI211_X1 U9466 ( .C1(n8890), .C2(n13020), .A(n8706), .B(n8705), .ZN(n12708)
         );
  XOR2_X1 U9467 ( .A(n12187), .B(n12196), .Z(n7420) );
  NOR2_X1 U9468 ( .A1(n8800), .A2(n11556), .ZN(n7421) );
  INV_X1 U9469 ( .A(n12996), .ZN(n8875) );
  INV_X1 U9470 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8370) );
  AND2_X1 U9471 ( .A1(n9150), .A2(n9149), .ZN(n7422) );
  NAND2_X1 U9472 ( .A1(n15004), .A2(n12979), .ZN(n13053) );
  INV_X1 U9473 ( .A(n13053), .ZN(n8912) );
  INV_X1 U9474 ( .A(n7557), .ZN(n7713) );
  OR2_X1 U9475 ( .A1(n8016), .A2(SI_20_), .ZN(n7423) );
  INV_X1 U9476 ( .A(n12038), .ZN(n13744) );
  INV_X1 U9477 ( .A(n11816), .ZN(n11503) );
  INV_X1 U9478 ( .A(n12789), .ZN(n12796) );
  INV_X4 U9479 ( .A(n7530), .ZN(n9678) );
  INV_X1 U9480 ( .A(n12706), .ZN(n12716) );
  OR2_X1 U9481 ( .A1(n8018), .A2(SI_21_), .ZN(n7424) );
  AND2_X1 U9482 ( .A1(n11944), .A2(n11943), .ZN(n7425) );
  INV_X1 U9483 ( .A(n11985), .ZN(n13383) );
  AND4_X1 U9484 ( .A1(n11711), .A2(n9349), .A3(n9348), .A4(n9347), .ZN(n7426)
         );
  INV_X1 U9485 ( .A(n11649), .ZN(n11783) );
  INV_X1 U9486 ( .A(n12609), .ZN(n12193) );
  AND2_X1 U9487 ( .A1(n10818), .A2(n12924), .ZN(n14977) );
  INV_X1 U9488 ( .A(n13411), .ZN(n13422) );
  OR2_X1 U9489 ( .A1(n13048), .A2(n13047), .ZN(P3_U3432) );
  OR2_X1 U9490 ( .A1(n12991), .A2(n12990), .ZN(P3_U3473) );
  AND2_X1 U9491 ( .A1(n14075), .A2(n14074), .ZN(n7429) );
  NAND2_X1 U9492 ( .A1(n7406), .A2(n9143), .ZN(n9144) );
  NAND2_X1 U9493 ( .A1(n7610), .A2(n7609), .ZN(n7629) );
  NAND2_X1 U9494 ( .A1(n7698), .A2(n7697), .ZN(n7729) );
  NOR2_X1 U9495 ( .A1(n7426), .A2(n7409), .ZN(n9368) );
  INV_X1 U9496 ( .A(n9399), .ZN(n9400) );
  NAND2_X1 U9497 ( .A1(n7848), .A2(n7847), .ZN(n7866) );
  INV_X1 U9498 ( .A(n7915), .ZN(n7916) );
  XNOR2_X1 U9499 ( .A(n11165), .B(n14189), .ZN(n9098) );
  INV_X1 U9500 ( .A(n9098), .ZN(n9587) );
  INV_X1 U9501 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8352) );
  INV_X1 U9502 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n7436) );
  INV_X1 U9503 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9057) );
  INV_X1 U9504 ( .A(n13265), .ZN(n8140) );
  AND4_X1 U9505 ( .A1(n9057), .A2(n9056), .A3(n9055), .A4(n9054), .ZN(n9058)
         );
  NAND2_X1 U9506 ( .A1(n12352), .A2(n12997), .ZN(n12189) );
  NAND2_X1 U9507 ( .A1(n14054), .A2(n10630), .ZN(n10312) );
  NAND2_X1 U9508 ( .A1(n14443), .A2(n12038), .ZN(n11672) );
  INV_X1 U9509 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7508) );
  AND2_X1 U9510 ( .A1(n11032), .A2(n8943), .ZN(n8941) );
  NAND2_X1 U9511 ( .A1(n8938), .A2(n8947), .ZN(n8948) );
  INV_X1 U9512 ( .A(n11406), .ZN(n11377) );
  NAND2_X1 U9513 ( .A1(n12844), .A2(n8809), .ZN(n12829) );
  INV_X1 U9514 ( .A(n12197), .ZN(n8790) );
  INV_X1 U9515 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7717) );
  INV_X1 U9516 ( .A(n13475), .ZN(n12014) );
  INV_X1 U9517 ( .A(n14021), .ZN(n11900) );
  NOR2_X1 U9518 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n9059) );
  AND2_X1 U9519 ( .A1(n11092), .A2(n8941), .ZN(n8942) );
  OAI21_X1 U9520 ( .B1(n12466), .B2(n12464), .A(n12806), .ZN(n8977) );
  OR2_X1 U9521 ( .A1(n8711), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8721) );
  INV_X1 U9522 ( .A(n9018), .ZN(n9027) );
  NAND2_X1 U9523 ( .A1(n11377), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n11378) );
  INV_X1 U9524 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n15111) );
  OR2_X1 U9525 ( .A1(n12702), .A2(n12408), .ZN(n8825) );
  INV_X1 U9526 ( .A(n14977), .ZN(n8900) );
  INV_X1 U9527 ( .A(n10818), .ZN(n12667) );
  OR2_X1 U9528 ( .A1(n8907), .A2(n8906), .ZN(n9018) );
  INV_X1 U9529 ( .A(n10397), .ZN(n10296) );
  OR2_X1 U9530 ( .A1(n7996), .A2(n7995), .ZN(n8025) );
  NAND2_X1 U9531 ( .A1(n7765), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7787) );
  INV_X1 U9532 ( .A(n12012), .ZN(n11990) );
  INV_X1 U9533 ( .A(n13523), .ZN(n12013) );
  INV_X1 U9534 ( .A(n13546), .ZN(n11648) );
  INV_X1 U9535 ( .A(n11656), .ZN(n11657) );
  NOR2_X1 U9536 ( .A1(n8266), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8271) );
  OR2_X1 U9537 ( .A1(n7899), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n7922) );
  INV_X1 U9538 ( .A(n11201), .ZN(n11204) );
  NAND2_X1 U9539 ( .A1(n9455), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9454) );
  INV_X1 U9540 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9356) );
  INV_X1 U9541 ( .A(n11865), .ZN(n9081) );
  OR2_X1 U9542 ( .A1(n9407), .A2(n9406), .ZN(n9419) );
  AND2_X1 U9543 ( .A1(n9374), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9393) );
  INV_X1 U9544 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9066) );
  INV_X1 U9545 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14217) );
  INV_X1 U9546 ( .A(n12679), .ZN(n12651) );
  OR2_X1 U9547 ( .A1(n8721), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8731) );
  AND2_X1 U9548 ( .A1(n8965), .A2(n12907), .ZN(n8966) );
  NAND2_X1 U9549 ( .A1(n8378), .A2(n8377), .ZN(n8711) );
  OR2_X1 U9550 ( .A1(n8975), .A2(n12791), .ZN(n8976) );
  INV_X1 U9551 ( .A(n11064), .ZN(n12359) );
  OR2_X1 U9552 ( .A1(n8779), .A2(n15011), .ZN(n8448) );
  INV_X1 U9553 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14201) );
  INV_X1 U9554 ( .A(n12529), .ZN(n12538) );
  AND2_X1 U9555 ( .A1(n10262), .A2(n10255), .ZN(n10259) );
  NAND2_X1 U9556 ( .A1(n12692), .A2(n8825), .ZN(n12678) );
  AND2_X1 U9557 ( .A1(n12797), .A2(n12796), .ZN(n12968) );
  INV_X1 U9558 ( .A(n12211), .ZN(n12808) );
  INV_X1 U9559 ( .A(n12207), .ZN(n12886) );
  AND2_X1 U9560 ( .A1(n10455), .A2(n12609), .ZN(n11064) );
  OR2_X1 U9561 ( .A1(n8463), .A2(n6632), .ZN(n8398) );
  NAND2_X1 U9562 ( .A1(n7420), .A2(n8900), .ZN(n8901) );
  NAND2_X1 U9563 ( .A1(n12218), .A2(n10538), .ZN(n12941) );
  AND2_X1 U9564 ( .A1(n8325), .A2(n8324), .ZN(n8645) );
  OR2_X1 U9565 ( .A1(n8580), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8601) );
  AND2_X1 U9566 ( .A1(n8297), .A2(n8296), .ZN(n8450) );
  OAI22_X1 U9567 ( .A1(n10185), .A2(n11850), .B1(n10337), .B2(n11963), .ZN(
        n10188) );
  INV_X1 U9568 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n13117) );
  AND2_X1 U9569 ( .A1(n10119), .A2(n8281), .ZN(n13167) );
  INV_X1 U9570 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n14658) );
  AND2_X1 U9571 ( .A1(n10203), .A2(n10202), .ZN(n11919) );
  OR2_X1 U9572 ( .A1(n8183), .A2(n8163), .ZN(n12016) );
  NOR2_X1 U9573 ( .A1(n8025), .A2(n8024), .ZN(n8044) );
  INV_X1 U9574 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9980) );
  OR2_X1 U9575 ( .A1(n10101), .A2(n10100), .ZN(n13225) );
  INV_X1 U9576 ( .A(n12006), .ZN(n13329) );
  NAND2_X1 U9577 ( .A1(n13411), .A2(n12013), .ZN(n13413) );
  NAND2_X1 U9578 ( .A1(n11334), .A2(n10562), .ZN(n13443) );
  INV_X1 U9579 ( .A(n10114), .ZN(n10115) );
  INV_X1 U9580 ( .A(n11839), .ZN(n11846) );
  AND2_X1 U9581 ( .A1(n10073), .A2(n10072), .ZN(n13430) );
  INV_X1 U9582 ( .A(n14840), .ZN(n14819) );
  INV_X2 U9583 ( .A(n7510), .ZN(n7530) );
  NAND2_X1 U9584 ( .A1(n11018), .A2(n11017), .ZN(n11019) );
  INV_X1 U9585 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9320) );
  INV_X1 U9586 ( .A(n13611), .ZN(n12089) );
  INV_X2 U9587 ( .A(n9733), .ZN(n9414) );
  NOR2_X1 U9588 ( .A1(n10635), .A2(n10634), .ZN(n10636) );
  INV_X1 U9589 ( .A(n9972), .ZN(n10321) );
  NOR2_X1 U9590 ( .A1(n9357), .A2(n9356), .ZN(n9374) );
  NOR2_X1 U9591 ( .A1(n9426), .A2(n13671), .ZN(n9438) );
  OR2_X1 U9592 ( .A1(n9136), .A2(n9103), .ZN(n9108) );
  INV_X1 U9593 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14198) );
  INV_X1 U9594 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14219) );
  INV_X1 U9595 ( .A(n11168), .ZN(n10239) );
  INV_X1 U9596 ( .A(n14032), .ZN(n12062) );
  INV_X1 U9597 ( .A(n14550), .ZN(n14530) );
  INV_X1 U9598 ( .A(n10233), .ZN(n10477) );
  AND3_X1 U9599 ( .A1(n10214), .A2(n10213), .A3(n10321), .ZN(n13862) );
  OR2_X1 U9600 ( .A1(n10216), .A2(n9973), .ZN(n14562) );
  INV_X1 U9601 ( .A(n10922), .ZN(n10996) );
  AND2_X1 U9602 ( .A1(n11168), .A2(n13826), .ZN(n14568) );
  OR2_X1 U9603 ( .A1(n11857), .A2(P1_B_REG_SCAN_IN), .ZN(n9727) );
  INV_X1 U9604 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9089) );
  OR2_X1 U9605 ( .A1(n9258), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n9285) );
  OR3_X1 U9606 ( .A1(n11535), .A2(n11477), .A3(n11255), .ZN(n9672) );
  OAI21_X1 U9607 ( .B1(n13011), .B2(n12485), .A(n9031), .ZN(n9032) );
  NAND2_X1 U9608 ( .A1(n8637), .A2(n8636), .ZN(n12974) );
  INV_X1 U9609 ( .A(n12479), .ZN(n12493) );
  AND2_X1 U9610 ( .A1(n9010), .A2(n10714), .ZN(n12477) );
  AOI21_X1 U9611 ( .B1(n12683), .B2(n8754), .A(n8736), .ZN(n12690) );
  AND4_X1 U9612 ( .A1(n8658), .A2(n8657), .A3(n8656), .A4(n8655), .ZN(n12775)
         );
  INV_X1 U9613 ( .A(n12623), .ZN(n14954) );
  AND2_X1 U9614 ( .A1(P3_U3897), .A2(n13068), .ZN(n14964) );
  NAND2_X1 U9615 ( .A1(n12688), .A2(n12329), .ZN(n12692) );
  OR2_X1 U9616 ( .A1(n10712), .A2(n10711), .ZN(n10715) );
  NAND2_X1 U9617 ( .A1(n8905), .A2(n12195), .ZN(n12878) );
  NOR2_X1 U9618 ( .A1(n10715), .A2(n11064), .ZN(n12914) );
  NAND2_X1 U9619 ( .A1(n15014), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9035) );
  AND2_X1 U9620 ( .A1(n8870), .A2(n8869), .ZN(n8871) );
  NAND2_X1 U9621 ( .A1(n12378), .A2(n8901), .ZN(n9034) );
  INV_X1 U9622 ( .A(n12941), .ZN(n12979) );
  OR2_X1 U9623 ( .A1(n9020), .A2(n9013), .ZN(n8911) );
  INV_X1 U9624 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8362) );
  XNOR2_X1 U9625 ( .A(n8835), .B(n8834), .ZN(n10252) );
  AND2_X1 U9626 ( .A1(n8327), .A2(n8326), .ZN(n8660) );
  INV_X1 U9627 ( .A(n13070), .ZN(n9693) );
  INV_X1 U9628 ( .A(n6474), .ZN(n8219) );
  INV_X1 U9629 ( .A(n14746), .ZN(n14783) );
  OAI21_X1 U9630 ( .B1(n9823), .B2(n9822), .A(n9821), .ZN(n9854) );
  INV_X1 U9631 ( .A(n12008), .ZN(n13318) );
  INV_X1 U9632 ( .A(n13453), .ZN(n13432) );
  INV_X1 U9633 ( .A(n13453), .ZN(n11334) );
  AND2_X1 U9634 ( .A1(n10338), .A2(n11456), .ZN(n14840) );
  AND2_X1 U9635 ( .A1(n10179), .A2(n14819), .ZN(n14812) );
  INV_X1 U9636 ( .A(n14812), .ZN(n14833) );
  AND2_X1 U9637 ( .A1(n10138), .A2(n10137), .ZN(n10336) );
  NAND2_X1 U9638 ( .A1(n9955), .A2(n10486), .ZN(n14606) );
  AND2_X1 U9639 ( .A1(n10324), .A2(n9965), .ZN(n11472) );
  INV_X1 U9640 ( .A(n14426), .ZN(n14412) );
  AND4_X1 U9641 ( .A1(n9460), .A2(n9459), .A3(n9458), .A4(n9457), .ZN(n13622)
         );
  NAND2_X1 U9642 ( .A1(n9148), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9152) );
  INV_X1 U9643 ( .A(n14517), .ZN(n14490) );
  AND2_X1 U9644 ( .A1(n9791), .A2(n9777), .ZN(n14483) );
  AND2_X1 U9645 ( .A1(n9791), .A2(n9665), .ZN(n14492) );
  OAI22_X1 U9646 ( .A1(n13983), .A2(n13980), .B1(n13623), .B2(n13677), .ZN(
        n13966) );
  INV_X1 U9647 ( .A(n14542), .ZN(n14033) );
  OR2_X1 U9648 ( .A1(n10475), .A2(n10474), .ZN(n14526) );
  AND2_X1 U9649 ( .A1(n9939), .A2(n9938), .ZN(n13858) );
  INV_X1 U9650 ( .A(n14549), .ZN(n14580) );
  INV_X1 U9651 ( .A(n14644), .ZN(n14581) );
  NAND2_X1 U9652 ( .A1(n14609), .A2(n14545), .ZN(n14644) );
  INV_X1 U9653 ( .A(n13858), .ZN(n10473) );
  NAND3_X1 U9654 ( .A1(n9727), .A2(n9726), .A3(n9725), .ZN(n9952) );
  INV_X1 U9655 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9100) );
  XNOR2_X1 U9656 ( .A(n15205), .B(n15204), .ZN(n15206) );
  AND2_X1 U9657 ( .A1(n10262), .A2(n10261), .ZN(n14943) );
  INV_X1 U9658 ( .A(n12482), .ZN(n12495) );
  NAND2_X1 U9659 ( .A1(n9012), .A2(n9011), .ZN(n12485) );
  AOI21_X1 U9660 ( .B1(n12640), .B2(n8754), .A(n8392), .ZN(n12652) );
  INV_X1 U9661 ( .A(n12775), .ZN(n12806) );
  INV_X1 U9662 ( .A(n14964), .ZN(n14939) );
  INV_X1 U9663 ( .A(n14943), .ZN(n14975) );
  INV_X1 U9664 ( .A(n14353), .ZN(n14959) );
  AND2_X1 U9665 ( .A1(n10715), .A2(n12910), .ZN(n12786) );
  AND2_X1 U9666 ( .A1(n11687), .A2(n11686), .ZN(n15003) );
  INV_X1 U9667 ( .A(n12888), .ZN(n12918) );
  NAND2_X1 U9668 ( .A1(n15016), .A2(n12979), .ZN(n12996) );
  INV_X1 U9669 ( .A(n15016), .ZN(n15014) );
  AND2_X1 U9670 ( .A1(n8915), .A2(n8914), .ZN(n8916) );
  INV_X2 U9671 ( .A(n15006), .ZN(n15004) );
  AND2_X1 U9672 ( .A1(n8911), .A2(n8910), .ZN(n15006) );
  NAND2_X1 U9673 ( .A1(n13055), .A2(n9759), .ZN(n9760) );
  INV_X1 U9674 ( .A(SI_29_), .ZN(n11869) );
  INV_X1 U9675 ( .A(SI_18_), .ZN(n15126) );
  INV_X1 U9676 ( .A(n11539), .ZN(n11545) );
  INV_X1 U9677 ( .A(n14752), .ZN(n14775) );
  INV_X1 U9678 ( .A(n13335), .ZN(n13491) );
  OR2_X1 U9679 ( .A1(n10205), .A2(P2_U3088), .ZN(n14672) );
  INV_X1 U9680 ( .A(n14669), .ZN(n13162) );
  INV_X1 U9681 ( .A(n14776), .ZN(n14707) );
  INV_X1 U9682 ( .A(n14778), .ZN(n14713) );
  AND2_X1 U9683 ( .A1(n11191), .A2(n11190), .ZN(n14403) );
  NAND2_X1 U9684 ( .A1(n11334), .A2(n10544), .ZN(n13449) );
  AND2_X2 U9685 ( .A1(n10331), .A2(n13385), .ZN(n13453) );
  INV_X1 U9686 ( .A(n14855), .ZN(n14853) );
  AND2_X1 U9687 ( .A1(n14403), .A2(n14402), .ZN(n14405) );
  AND2_X1 U9688 ( .A1(n14843), .A2(n14842), .ZN(n14854) );
  NAND2_X1 U9689 ( .A1(n10113), .A2(n14795), .ZN(n14793) );
  INV_X1 U9690 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11777) );
  INV_X1 U9691 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11106) );
  INV_X1 U9692 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9891) );
  OR2_X1 U9693 ( .A1(n9668), .A2(n9667), .ZN(n9669) );
  OR2_X1 U9694 ( .A1(n9378), .A2(n9377), .ZN(n14032) );
  OR2_X1 U9695 ( .A1(n9774), .A2(n9773), .ZN(n14517) );
  INV_X1 U9696 ( .A(n14492), .ZN(n14521) );
  INV_X1 U9697 ( .A(n14571), .ZN(n14536) );
  INV_X1 U9698 ( .A(n14657), .ZN(n14655) );
  INV_X1 U9699 ( .A(n14646), .ZN(n14645) );
  AND2_X1 U9700 ( .A1(n10322), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9731) );
  INV_X1 U9701 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14186) );
  INV_X1 U9702 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10536) );
  AND2_X2 U9703 ( .A1(n13055), .A2(n9673), .ZN(P3_U3897) );
  OAI211_X1 U9704 ( .C1(n12485), .C2(n8826), .A(n9050), .B(n9049), .ZN(
        P3_U3165) );
  NAND2_X1 U9705 ( .A1(n9038), .A2(n9037), .ZN(P3_U3488) );
  NAND2_X1 U9706 ( .A1(n8917), .A2(n8916), .ZN(P3_U3456) );
  NOR3_X1 U9707 ( .A1(n9823), .A2(n9822), .A3(P2_U3088), .ZN(P2_U3947) );
  NOR2_X1 U9708 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7431) );
  NAND4_X1 U9709 ( .A1(n7491), .A2(n7434), .A3(n7433), .A4(n7432), .ZN(n7435)
         );
  NOR2_X2 U9710 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7535) );
  INV_X1 U9711 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7437) );
  NAND2_X1 U9712 ( .A1(n7535), .A2(n7437), .ZN(n7558) );
  INV_X1 U9713 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7443) );
  INV_X1 U9714 ( .A(n7470), .ZN(n7444) );
  NAND2_X1 U9715 ( .A1(n7444), .A2(n7447), .ZN(n7473) );
  NAND2_X1 U9716 ( .A1(n7448), .A2(n7445), .ZN(n7449) );
  AND2_X1 U9717 ( .A1(n13577), .A2(n7449), .ZN(n7450) );
  XNOR2_X2 U9718 ( .A(n7453), .B(n7452), .ZN(n7456) );
  NAND2_X1 U9719 ( .A1(n6474), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7460) );
  INV_X1 U9720 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9894) );
  INV_X1 U9721 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9898) );
  NAND3_X1 U9722 ( .A1(n13262), .A2(n7461), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7463) );
  NAND2_X1 U9723 ( .A1(n7463), .A2(n7462), .ZN(n7468) );
  INV_X1 U9724 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7464) );
  NAND3_X1 U9725 ( .A1(n7465), .A2(n14307), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7466) );
  NAND2_X1 U9726 ( .A1(n7466), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7467) );
  NAND2_X1 U9727 ( .A1(n9678), .A2(SI_0_), .ZN(n7469) );
  NAND2_X1 U9728 ( .A1(n7470), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7471) );
  NAND2_X1 U9729 ( .A1(n7474), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7475) );
  NAND2_X1 U9730 ( .A1(n7476), .A2(n7488), .ZN(n7483) );
  OR2_X1 U9731 ( .A1(n7484), .A2(n7445), .ZN(n7478) );
  OR2_X1 U9732 ( .A1(n7478), .A2(n7477), .ZN(n7482) );
  INV_X1 U9733 ( .A(n7484), .ZN(n7485) );
  NAND2_X1 U9734 ( .A1(n7488), .A2(n6840), .ZN(n7782) );
  AND2_X1 U9735 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n7490) );
  NAND2_X1 U9736 ( .A1(n7826), .A2(n7490), .ZN(n7498) );
  NOR2_X1 U9737 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n7493) );
  INV_X1 U9738 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7492) );
  NAND3_X1 U9739 ( .A1(n7491), .A2(n7493), .A3(n7492), .ZN(n7496) );
  INV_X1 U9740 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7804) );
  NAND2_X1 U9741 ( .A1(n7804), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n7495) );
  XNOR2_X1 U9742 ( .A(P2_IR_REG_31__SCAN_IN), .B(P2_IR_REG_19__SCAN_IN), .ZN(
        n7494) );
  OAI21_X1 U9743 ( .B1(n7496), .B2(n7495), .A(n7494), .ZN(n7497) );
  NAND2_X1 U9744 ( .A1(n8242), .A2(n7591), .ZN(n7501) );
  INV_X1 U9745 ( .A(n10178), .ZN(n10333) );
  NAND3_X1 U9746 ( .A1(n7501), .A2(n7500), .A3(n7499), .ZN(n7545) );
  INV_X1 U9747 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9847) );
  INV_X1 U9748 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10590) );
  OR2_X1 U9749 ( .A1(n8068), .A2(n10590), .ZN(n7504) );
  NAND2_X1 U9750 ( .A1(n6475), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7502) );
  NAND2_X1 U9751 ( .A1(n13202), .A2(n7516), .ZN(n7518) );
  AND2_X2 U9752 ( .A1(n9819), .A2(n7530), .ZN(n7557) );
  NAND2_X1 U9753 ( .A1(n7557), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7515) );
  NAND2_X1 U9754 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7506) );
  NAND2_X1 U9755 ( .A1(n7510), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7507) );
  OAI21_X1 U9756 ( .B1(n7510), .B2(n7508), .A(n7507), .ZN(n7509) );
  INV_X1 U9757 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9120) );
  INV_X1 U9758 ( .A(SI_0_), .ZN(n9714) );
  INV_X1 U9759 ( .A(n7511), .ZN(n7512) );
  NAND2_X1 U9760 ( .A1(n7513), .A2(n7512), .ZN(n7514) );
  NAND2_X1 U9761 ( .A1(n7526), .A2(n7514), .ZN(n9712) );
  NAND2_X1 U9762 ( .A1(n10078), .A2(n7591), .ZN(n7517) );
  NAND2_X1 U9763 ( .A1(n7518), .A2(n7517), .ZN(n7544) );
  INV_X1 U9764 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7519) );
  NAND2_X1 U9765 ( .A1(n6474), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7523) );
  INV_X1 U9766 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n13462) );
  OR2_X1 U9767 ( .A1(n8185), .A2(n13462), .ZN(n7522) );
  INV_X1 U9768 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7520) );
  NAND2_X1 U9769 ( .A1(n10068), .A2(n7516), .ZN(n7539) );
  NAND2_X1 U9770 ( .A1(n7526), .A2(n7525), .ZN(n7529) );
  INV_X1 U9771 ( .A(n7529), .ZN(n7528) );
  INV_X1 U9772 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9674) );
  MUX2_X1 U9773 ( .A(n9674), .B(n9676), .S(n6478), .Z(n7532) );
  NAND2_X1 U9774 ( .A1(n7533), .A2(n7532), .ZN(n7534) );
  AND2_X1 U9775 ( .A1(n7554), .A2(n7534), .ZN(n9129) );
  NAND2_X1 U9776 ( .A1(n9129), .A2(n6486), .ZN(n7537) );
  OR2_X1 U9777 ( .A1(n7535), .A2(n7445), .ZN(n7536) );
  XNOR2_X1 U9778 ( .A(n7536), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9849) );
  NAND2_X1 U9779 ( .A1(n13459), .A2(n8034), .ZN(n7538) );
  AND2_X1 U9780 ( .A1(n7539), .A2(n7538), .ZN(n7547) );
  NAND2_X1 U9781 ( .A1(n10068), .A2(n8034), .ZN(n7541) );
  NAND2_X1 U9782 ( .A1(n13459), .A2(n7516), .ZN(n7540) );
  NAND2_X1 U9783 ( .A1(n7541), .A2(n7540), .ZN(n7546) );
  NAND2_X1 U9784 ( .A1(n7547), .A2(n7546), .ZN(n7542) );
  OAI21_X1 U9785 ( .B1(n7545), .B2(n7544), .A(n7542), .ZN(n7552) );
  AOI22_X1 U9786 ( .A1(n13202), .A2(n7591), .B1(n7516), .B2(n10078), .ZN(n7543) );
  AOI21_X1 U9787 ( .B1(n7545), .B2(n7544), .A(n7543), .ZN(n7551) );
  INV_X1 U9788 ( .A(n7546), .ZN(n7549) );
  INV_X1 U9789 ( .A(n7547), .ZN(n7548) );
  NAND2_X1 U9790 ( .A1(n7549), .A2(n7548), .ZN(n7550) );
  OAI21_X1 U9791 ( .B1(n7552), .B2(n7551), .A(n7550), .ZN(n7572) );
  NAND2_X1 U9792 ( .A1(n7554), .A2(n7553), .ZN(n7582) );
  MUX2_X1 U9793 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n6478), .Z(n7555) );
  NAND2_X1 U9794 ( .A1(n7555), .A2(SI_3_), .ZN(n7579) );
  OAI21_X1 U9795 ( .B1(n7555), .B2(SI_3_), .A(n7579), .ZN(n7578) );
  XNOR2_X1 U9796 ( .A(n7582), .B(n7578), .ZN(n9683) );
  NAND2_X1 U9797 ( .A1(n9683), .A2(n8210), .ZN(n7561) );
  NAND2_X1 U9798 ( .A1(n7558), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7559) );
  XNOR2_X1 U9799 ( .A(n7559), .B(P2_IR_REG_3__SCAN_IN), .ZN(n9851) );
  AOI22_X1 U9800 ( .A1(n7557), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n7943), .B2(
        n9851), .ZN(n7560) );
  INV_X1 U9801 ( .A(n7516), .ZN(n8034) );
  NAND2_X1 U9802 ( .A1(n10843), .A2(n7591), .ZN(n7568) );
  OR2_X1 U9803 ( .A1(n8068), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7566) );
  NAND2_X1 U9804 ( .A1(n6475), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7565) );
  INV_X1 U9805 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9850) );
  OR2_X1 U9806 ( .A1(n8185), .A2(n9850), .ZN(n7564) );
  INV_X1 U9807 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7562) );
  OR2_X1 U9808 ( .A1(n6473), .A2(n7562), .ZN(n7563) );
  NAND4_X1 U9809 ( .A1(n7566), .A2(n7565), .A3(n7564), .A4(n7563), .ZN(n13201)
         );
  NAND2_X1 U9810 ( .A1(n13201), .A2(n6481), .ZN(n7567) );
  NAND2_X1 U9811 ( .A1(n7568), .A2(n7567), .ZN(n7573) );
  NAND2_X1 U9812 ( .A1(n7572), .A2(n7573), .ZN(n7571) );
  INV_X1 U9813 ( .A(n13201), .ZN(n10545) );
  NAND2_X1 U9814 ( .A1(n10843), .A2(n6481), .ZN(n7569) );
  OAI21_X1 U9815 ( .B1(n10545), .B2(n6481), .A(n7569), .ZN(n7570) );
  NAND2_X1 U9816 ( .A1(n7571), .A2(n7570), .ZN(n7577) );
  INV_X1 U9817 ( .A(n7572), .ZN(n7575) );
  INV_X1 U9818 ( .A(n7573), .ZN(n7574) );
  NAND2_X1 U9819 ( .A1(n7575), .A2(n7574), .ZN(n7576) );
  NAND2_X1 U9820 ( .A1(n7577), .A2(n7576), .ZN(n7605) );
  INV_X1 U9821 ( .A(n7578), .ZN(n7581) );
  INV_X1 U9822 ( .A(n7579), .ZN(n7580) );
  OAI21_X1 U9823 ( .B1(n7583), .B2(SI_4_), .A(n7611), .ZN(n7584) );
  NAND2_X1 U9824 ( .A1(n7585), .A2(n7584), .ZN(n7586) );
  NAND2_X1 U9825 ( .A1(n7586), .A2(n7612), .ZN(n9691) );
  OR2_X1 U9826 ( .A1(n9691), .A2(n7556), .ZN(n7590) );
  NAND2_X1 U9827 ( .A1(n7587), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7588) );
  XNOR2_X1 U9828 ( .A(n7588), .B(P2_IR_REG_4__SCAN_IN), .ZN(n13210) );
  AOI22_X1 U9829 ( .A1(n7557), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7943), .B2(
        n13210), .ZN(n7589) );
  NAND2_X1 U9830 ( .A1(n14802), .A2(n6481), .ZN(n7600) );
  NAND2_X1 U9831 ( .A1(n6475), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7598) );
  NOR2_X1 U9832 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7593) );
  NOR2_X1 U9833 ( .A1(n7619), .A2(n7593), .ZN(n10603) );
  NAND2_X1 U9834 ( .A1(n7592), .A2(n10603), .ZN(n7597) );
  INV_X1 U9835 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10613) );
  OR2_X1 U9836 ( .A1(n8185), .A2(n10613), .ZN(n7596) );
  INV_X1 U9837 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7594) );
  OR2_X1 U9838 ( .A1(n6473), .A2(n7594), .ZN(n7595) );
  NAND4_X1 U9839 ( .A1(n7598), .A2(n7597), .A3(n7596), .A4(n7595), .ZN(n13200)
         );
  NAND2_X1 U9840 ( .A1(n13200), .A2(n8222), .ZN(n7599) );
  NAND2_X1 U9841 ( .A1(n7600), .A2(n7599), .ZN(n7606) );
  NAND2_X1 U9842 ( .A1(n7605), .A2(n7606), .ZN(n7604) );
  NAND2_X1 U9843 ( .A1(n14802), .A2(n8222), .ZN(n7602) );
  NAND2_X1 U9844 ( .A1(n13200), .A2(n6481), .ZN(n7601) );
  NAND2_X1 U9845 ( .A1(n7602), .A2(n7601), .ZN(n7603) );
  NAND2_X1 U9846 ( .A1(n7604), .A2(n7603), .ZN(n7610) );
  INV_X1 U9847 ( .A(n7605), .ZN(n7608) );
  INV_X1 U9848 ( .A(n7606), .ZN(n7607) );
  NAND2_X1 U9849 ( .A1(n7608), .A2(n7607), .ZN(n7609) );
  MUX2_X1 U9850 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9678), .Z(n7613) );
  NAND2_X1 U9851 ( .A1(n7613), .A2(SI_5_), .ZN(n7630) );
  OAI21_X1 U9852 ( .B1(n7613), .B2(SI_5_), .A(n7630), .ZN(n7614) );
  INV_X1 U9853 ( .A(n7614), .ZN(n7615) );
  NAND2_X1 U9854 ( .A1(n9717), .A2(n8210), .ZN(n7618) );
  OAI21_X1 U9855 ( .B1(n7587), .B2(P2_IR_REG_4__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7616) );
  XNOR2_X1 U9856 ( .A(n7616), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9852) );
  AOI22_X1 U9857 ( .A1(n7557), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7943), .B2(
        n9852), .ZN(n7617) );
  NAND2_X1 U9858 ( .A1(n14808), .A2(n8222), .ZN(n7626) );
  NAND2_X1 U9859 ( .A1(n7619), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7641) );
  OAI21_X1 U9860 ( .B1(n7619), .B2(P2_REG3_REG_5__SCAN_IN), .A(n7641), .ZN(
        n10563) );
  NAND2_X1 U9861 ( .A1(n6475), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7623) );
  INV_X1 U9862 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10557) );
  OR2_X1 U9863 ( .A1(n8185), .A2(n10557), .ZN(n7622) );
  INV_X1 U9864 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7620) );
  OR2_X1 U9865 ( .A1(n6473), .A2(n7620), .ZN(n7621) );
  NAND2_X1 U9866 ( .A1(n13199), .A2(n6481), .ZN(n7625) );
  NAND2_X1 U9867 ( .A1(n7626), .A2(n7625), .ZN(n7628) );
  AOI22_X1 U9868 ( .A1(n14808), .A2(n6481), .B1(n8222), .B2(n13199), .ZN(n7627) );
  NAND2_X1 U9869 ( .A1(n7631), .A2(n7630), .ZN(n7635) );
  MUX2_X1 U9870 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9678), .Z(n7632) );
  NAND2_X1 U9871 ( .A1(n7632), .A2(SI_6_), .ZN(n7658) );
  OAI21_X1 U9872 ( .B1(SI_6_), .B2(n7632), .A(n7658), .ZN(n7633) );
  INV_X1 U9873 ( .A(n7633), .ZN(n7634) );
  OR2_X1 U9874 ( .A1(n7488), .A2(n7445), .ZN(n7637) );
  XNOR2_X1 U9875 ( .A(n7637), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10035) );
  AOI22_X1 U9876 ( .A1(n7557), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7943), .B2(
        n10035), .ZN(n7638) );
  NAND2_X1 U9877 ( .A1(n14815), .A2(n6481), .ZN(n7649) );
  INV_X1 U9878 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7640) );
  AND2_X1 U9879 ( .A1(n7641), .A2(n7640), .ZN(n7642) );
  NOR2_X1 U9880 ( .A1(n7641), .A2(n7640), .ZN(n7665) );
  OR2_X1 U9881 ( .A1(n7642), .A2(n7665), .ZN(n10583) );
  OR2_X1 U9882 ( .A1(n8184), .A2(n10583), .ZN(n7647) );
  NAND2_X1 U9883 ( .A1(n6474), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7646) );
  INV_X1 U9884 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10580) );
  OR2_X1 U9885 ( .A1(n8185), .A2(n10580), .ZN(n7645) );
  INV_X1 U9886 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7643) );
  OR2_X1 U9887 ( .A1(n6473), .A2(n7643), .ZN(n7644) );
  NAND4_X1 U9888 ( .A1(n7647), .A2(n7646), .A3(n7645), .A4(n7644), .ZN(n13198)
         );
  NAND2_X1 U9889 ( .A1(n13198), .A2(n8222), .ZN(n7648) );
  NAND2_X1 U9890 ( .A1(n7649), .A2(n7648), .ZN(n7655) );
  NAND2_X1 U9891 ( .A1(n14815), .A2(n8222), .ZN(n7651) );
  NAND2_X1 U9892 ( .A1(n13198), .A2(n6481), .ZN(n7650) );
  NAND2_X1 U9893 ( .A1(n7651), .A2(n7650), .ZN(n7652) );
  NAND2_X1 U9894 ( .A1(n7653), .A2(n7652), .ZN(n7657) );
  NAND2_X1 U9895 ( .A1(n7657), .A2(n7656), .ZN(n7675) );
  MUX2_X1 U9896 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6478), .Z(n7660) );
  NAND2_X1 U9897 ( .A1(n7660), .A2(SI_7_), .ZN(n7679) );
  OAI21_X1 U9898 ( .B1(n7660), .B2(SI_7_), .A(n7679), .ZN(n7676) );
  XNOR2_X1 U9899 ( .A(n7678), .B(n7676), .ZN(n9746) );
  NAND2_X1 U9900 ( .A1(n9746), .A2(n8210), .ZN(n7664) );
  NAND2_X1 U9901 ( .A1(n7488), .A2(n7661), .ZN(n7681) );
  NAND2_X1 U9902 ( .A1(n7681), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7662) );
  XNOR2_X1 U9903 ( .A(n7662), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9983) );
  AOI22_X1 U9904 ( .A1(n7557), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7943), .B2(
        n9983), .ZN(n7663) );
  NAND2_X1 U9905 ( .A1(n7664), .A2(n7663), .ZN(n10665) );
  NAND2_X1 U9906 ( .A1(n10665), .A2(n8222), .ZN(n7673) );
  NAND2_X1 U9907 ( .A1(n7665), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7685) );
  OR2_X1 U9908 ( .A1(n7665), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7666) );
  NAND2_X1 U9909 ( .A1(n7685), .A2(n7666), .ZN(n10770) );
  OR2_X1 U9910 ( .A1(n8068), .A2(n10770), .ZN(n7671) );
  NAND2_X1 U9911 ( .A1(n6474), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7670) );
  INV_X1 U9912 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10777) );
  OR2_X1 U9913 ( .A1(n8185), .A2(n10777), .ZN(n7669) );
  INV_X1 U9914 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7667) );
  OR2_X1 U9915 ( .A1(n6473), .A2(n7667), .ZN(n7668) );
  NAND4_X1 U9916 ( .A1(n7671), .A2(n7670), .A3(n7669), .A4(n7668), .ZN(n13197)
         );
  NAND2_X1 U9917 ( .A1(n13197), .A2(n6481), .ZN(n7672) );
  AOI22_X1 U9918 ( .A1(n10665), .A2(n6481), .B1(n8222), .B2(n13197), .ZN(n7674) );
  INV_X1 U9919 ( .A(n7676), .ZN(n7677) );
  MUX2_X1 U9920 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9678), .Z(n7680) );
  NAND2_X1 U9921 ( .A1(n7680), .A2(SI_8_), .ZN(n7701) );
  OAI21_X1 U9922 ( .B1(SI_8_), .B2(n7680), .A(n7701), .ZN(n7699) );
  XNOR2_X1 U9923 ( .A(n7700), .B(n7699), .ZN(n9751) );
  NAND2_X1 U9924 ( .A1(n9751), .A2(n8210), .ZN(n7684) );
  NAND2_X1 U9925 ( .A1(n7707), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7682) );
  XNOR2_X1 U9926 ( .A(n7682), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10094) );
  AOI22_X1 U9927 ( .A1(n7557), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7943), .B2(
        n10094), .ZN(n7683) );
  NAND2_X1 U9928 ( .A1(n10790), .A2(n6481), .ZN(n7693) );
  NAND2_X1 U9929 ( .A1(n7685), .A2(n9980), .ZN(n7686) );
  NAND2_X1 U9930 ( .A1(n7718), .A2(n7686), .ZN(n10787) );
  OR2_X1 U9931 ( .A1(n8184), .A2(n10787), .ZN(n7691) );
  NAND2_X1 U9932 ( .A1(n6475), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7690) );
  INV_X1 U9933 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10788) );
  OR2_X1 U9934 ( .A1(n8185), .A2(n10788), .ZN(n7689) );
  INV_X1 U9935 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7687) );
  OR2_X1 U9936 ( .A1(n6473), .A2(n7687), .ZN(n7688) );
  NAND4_X1 U9937 ( .A1(n7691), .A2(n7690), .A3(n7689), .A4(n7688), .ZN(n13196)
         );
  NAND2_X1 U9938 ( .A1(n13196), .A2(n8222), .ZN(n7692) );
  INV_X1 U9939 ( .A(n13196), .ZN(n10729) );
  NAND2_X1 U9940 ( .A1(n10790), .A2(n8222), .ZN(n7694) );
  OAI21_X1 U9941 ( .B1(n10729), .B2(n8222), .A(n7694), .ZN(n7695) );
  NAND2_X1 U9942 ( .A1(n7696), .A2(n7695), .ZN(n7698) );
  MUX2_X1 U9943 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9678), .Z(n7702) );
  NAND2_X1 U9944 ( .A1(n7702), .A2(SI_9_), .ZN(n7754) );
  OAI21_X1 U9945 ( .B1(n7702), .B2(SI_9_), .A(n7754), .ZN(n7703) );
  INV_X1 U9946 ( .A(n7703), .ZN(n7704) );
  OR2_X1 U9947 ( .A1(n7705), .A2(n7704), .ZN(n7706) );
  NAND2_X1 U9948 ( .A1(n7760), .A2(n7706), .ZN(n9758) );
  OR2_X1 U9949 ( .A1(n9758), .A2(n7556), .ZN(n7716) );
  NAND2_X1 U9950 ( .A1(n7709), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7708) );
  MUX2_X1 U9951 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7708), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n7712) );
  INV_X1 U9952 ( .A(n7709), .ZN(n7711) );
  INV_X1 U9953 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7710) );
  NAND2_X1 U9954 ( .A1(n7711), .A2(n7710), .ZN(n7761) );
  NAND2_X1 U9955 ( .A1(n7712), .A2(n7761), .ZN(n14722) );
  OAI22_X1 U9956 ( .A1(n7713), .A2(n9756), .B1(n9819), .B2(n14722), .ZN(n7714)
         );
  INV_X1 U9957 ( .A(n7714), .ZN(n7715) );
  NAND2_X1 U9958 ( .A1(n10887), .A2(n8222), .ZN(n7726) );
  AND2_X1 U9959 ( .A1(n7718), .A2(n7717), .ZN(n7719) );
  OR2_X1 U9960 ( .A1(n7719), .A2(n7735), .ZN(n10761) );
  OR2_X1 U9961 ( .A1(n8184), .A2(n10761), .ZN(n7724) );
  NAND2_X1 U9962 ( .A1(n6475), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7723) );
  INV_X1 U9963 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10738) );
  OR2_X1 U9964 ( .A1(n8185), .A2(n10738), .ZN(n7722) );
  INV_X1 U9965 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7720) );
  OR2_X1 U9966 ( .A1(n8187), .A2(n7720), .ZN(n7721) );
  NAND4_X1 U9967 ( .A1(n7724), .A2(n7723), .A3(n7722), .A4(n7721), .ZN(n13195)
         );
  NAND2_X1 U9968 ( .A1(n13195), .A2(n6481), .ZN(n7725) );
  NAND2_X1 U9969 ( .A1(n7726), .A2(n7725), .ZN(n7728) );
  AOI22_X1 U9970 ( .A1(n10887), .A2(n6481), .B1(n8222), .B2(n13195), .ZN(n7727) );
  NAND2_X1 U9971 ( .A1(n7760), .A2(n7754), .ZN(n7731) );
  MUX2_X1 U9972 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9678), .Z(n7730) );
  OAI21_X1 U9973 ( .B1(n7730), .B2(SI_10_), .A(n7755), .ZN(n7756) );
  XNOR2_X1 U9974 ( .A(n7731), .B(n7756), .ZN(n9761) );
  NAND2_X1 U9975 ( .A1(n9761), .A2(n8210), .ZN(n7734) );
  NAND2_X1 U9976 ( .A1(n7761), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7732) );
  XNOR2_X1 U9977 ( .A(n7732), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10980) );
  AOI22_X1 U9978 ( .A1(n8211), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n10980), 
        .B2(n7943), .ZN(n7733) );
  NAND2_X1 U9979 ( .A1(n11072), .A2(n6481), .ZN(n7744) );
  NOR2_X1 U9980 ( .A1(n7735), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7736) );
  OR2_X1 U9981 ( .A1(n7765), .A2(n7736), .ZN(n10896) );
  OR2_X1 U9982 ( .A1(n8068), .A2(n10896), .ZN(n7742) );
  NAND2_X1 U9983 ( .A1(n6475), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7741) );
  INV_X1 U9984 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7737) );
  OR2_X1 U9985 ( .A1(n8185), .A2(n7737), .ZN(n7740) );
  INV_X1 U9986 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7738) );
  OR2_X1 U9987 ( .A1(n8187), .A2(n7738), .ZN(n7739) );
  NAND4_X1 U9988 ( .A1(n7742), .A2(n7741), .A3(n7740), .A4(n7739), .ZN(n13194)
         );
  NAND2_X1 U9989 ( .A1(n13194), .A2(n8222), .ZN(n7743) );
  NAND2_X1 U9990 ( .A1(n7744), .A2(n7743), .ZN(n7749) );
  INV_X1 U9991 ( .A(n13194), .ZN(n8246) );
  NAND2_X1 U9992 ( .A1(n11072), .A2(n8222), .ZN(n7745) );
  OAI21_X1 U9993 ( .B1(n8246), .B2(n8222), .A(n7745), .ZN(n7746) );
  NAND2_X1 U9994 ( .A1(n7747), .A2(n7746), .ZN(n7753) );
  INV_X1 U9995 ( .A(n7748), .ZN(n7751) );
  INV_X1 U9996 ( .A(n7749), .ZN(n7750) );
  NAND2_X1 U9997 ( .A1(n7751), .A2(n7750), .ZN(n7752) );
  AND2_X1 U9998 ( .A1(n7754), .A2(n7755), .ZN(n7759) );
  INV_X1 U9999 ( .A(n7755), .ZN(n7758) );
  INV_X1 U10000 ( .A(n7756), .ZN(n7757) );
  MUX2_X1 U10001 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n9678), .Z(n7778) );
  XNOR2_X1 U10002 ( .A(n7778), .B(SI_11_), .ZN(n7780) );
  XNOR2_X1 U10003 ( .A(n7781), .B(n7780), .ZN(n9890) );
  NAND2_X1 U10004 ( .A1(n9890), .A2(n8210), .ZN(n7764) );
  OAI21_X1 U10005 ( .B1(n7761), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7762) );
  XNOR2_X1 U10006 ( .A(n7762), .B(P2_IR_REG_11__SCAN_IN), .ZN(n13228) );
  AOI22_X1 U10007 ( .A1(n13228), .A2(n7943), .B1(n8211), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n7763) );
  NAND2_X1 U10008 ( .A1(n11183), .A2(n8222), .ZN(n7773) );
  OR2_X1 U10009 ( .A1(n7765), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7766) );
  NAND2_X1 U10010 ( .A1(n7787), .A2(n7766), .ZN(n11086) );
  OR2_X1 U10011 ( .A1(n8068), .A2(n11086), .ZN(n7771) );
  NAND2_X1 U10012 ( .A1(n6475), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7770) );
  INV_X1 U10013 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11087) );
  OR2_X1 U10014 ( .A1(n8185), .A2(n11087), .ZN(n7769) );
  INV_X1 U10015 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7767) );
  OR2_X1 U10016 ( .A1(n8187), .A2(n7767), .ZN(n7768) );
  NAND4_X1 U10017 ( .A1(n7771), .A2(n7770), .A3(n7769), .A4(n7768), .ZN(n13193) );
  NAND2_X1 U10018 ( .A1(n13193), .A2(n6481), .ZN(n7772) );
  NAND2_X1 U10019 ( .A1(n7773), .A2(n7772), .ZN(n7776) );
  INV_X1 U10020 ( .A(n13193), .ZN(n11182) );
  NAND2_X1 U10021 ( .A1(n11183), .A2(n6481), .ZN(n7774) );
  OAI21_X1 U10022 ( .B1(n11182), .B2(n6481), .A(n7774), .ZN(n7775) );
  INV_X1 U10023 ( .A(n7776), .ZN(n7777) );
  INV_X1 U10024 ( .A(n7778), .ZN(n7779) );
  MUX2_X1 U10025 ( .A(n8310), .B(n10086), .S(n9678), .Z(n7802) );
  XNOR2_X1 U10026 ( .A(n7802), .B(SI_12_), .ZN(n7800) );
  XNOR2_X1 U10027 ( .A(n7801), .B(n7800), .ZN(n10011) );
  NAND2_X1 U10028 ( .A1(n10011), .A2(n8210), .ZN(n7785) );
  NAND2_X1 U10029 ( .A1(n7782), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7783) );
  XNOR2_X1 U10030 ( .A(n7783), .B(P2_IR_REG_12__SCAN_IN), .ZN(n14749) );
  AOI22_X1 U10031 ( .A1(n8211), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7943), 
        .B2(n14749), .ZN(n7784) );
  NAND2_X1 U10032 ( .A1(n11290), .A2(n8111), .ZN(n7795) );
  INV_X1 U10033 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7786) );
  NAND2_X1 U10034 ( .A1(n7787), .A2(n7786), .ZN(n7788) );
  NAND2_X1 U10035 ( .A1(n7808), .A2(n7788), .ZN(n11251) );
  OR2_X1 U10036 ( .A1(n8184), .A2(n11251), .ZN(n7793) );
  NAND2_X1 U10037 ( .A1(n6474), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7792) );
  INV_X1 U10038 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11193) );
  OR2_X1 U10039 ( .A1(n8185), .A2(n11193), .ZN(n7791) );
  INV_X1 U10040 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7789) );
  OR2_X1 U10041 ( .A1(n6473), .A2(n7789), .ZN(n7790) );
  NAND4_X1 U10042 ( .A1(n7793), .A2(n7792), .A3(n7791), .A4(n7790), .ZN(n13192) );
  NAND2_X1 U10043 ( .A1(n13192), .A2(n8223), .ZN(n7794) );
  NAND2_X1 U10044 ( .A1(n7795), .A2(n7794), .ZN(n7797) );
  AOI22_X1 U10045 ( .A1(n11290), .A2(n8223), .B1(n13192), .B2(n8111), .ZN(
        n7796) );
  AOI21_X1 U10046 ( .B1(n7798), .B2(n7797), .A(n7796), .ZN(n7799) );
  MUX2_X1 U10047 ( .A(n10109), .B(n10111), .S(n9678), .Z(n7820) );
  XNOR2_X1 U10048 ( .A(n7820), .B(SI_13_), .ZN(n7803) );
  XNOR2_X1 U10049 ( .A(n7824), .B(n7803), .ZN(n10108) );
  NAND2_X1 U10050 ( .A1(n10108), .A2(n8210), .ZN(n7807) );
  NAND2_X1 U10051 ( .A1(n7826), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7805) );
  XNOR2_X1 U10052 ( .A(n7805), .B(n7804), .ZN(n10987) );
  INV_X1 U10053 ( .A(n10987), .ZN(n14754) );
  AOI22_X1 U10054 ( .A1(n8211), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7943), 
        .B2(n14754), .ZN(n7806) );
  NAND2_X1 U10055 ( .A1(n14670), .A2(n8223), .ZN(n7817) );
  NAND2_X1 U10056 ( .A1(n7808), .A2(n14658), .ZN(n7809) );
  NAND2_X1 U10057 ( .A1(n7831), .A2(n7809), .ZN(n14673) );
  INV_X1 U10058 ( .A(n14673), .ZN(n7810) );
  NAND2_X1 U10059 ( .A1(n7592), .A2(n7810), .ZN(n7815) );
  NAND2_X1 U10060 ( .A1(n6474), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7814) );
  INV_X1 U10061 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11300) );
  OR2_X1 U10062 ( .A1(n8185), .A2(n11300), .ZN(n7813) );
  INV_X1 U10063 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7811) );
  OR2_X1 U10064 ( .A1(n6473), .A2(n7811), .ZN(n7812) );
  NAND4_X1 U10065 ( .A1(n7815), .A2(n7814), .A3(n7813), .A4(n7812), .ZN(n13191) );
  NAND2_X1 U10066 ( .A1(n13191), .A2(n6481), .ZN(n7816) );
  NAND2_X1 U10067 ( .A1(n7817), .A2(n7816), .ZN(n7819) );
  AOI22_X1 U10068 ( .A1(n14670), .A2(n6481), .B1(n8222), .B2(n13191), .ZN(
        n7818) );
  NOR2_X1 U10069 ( .A1(n7821), .A2(SI_13_), .ZN(n7823) );
  NAND2_X1 U10070 ( .A1(n7821), .A2(SI_13_), .ZN(n7822) );
  MUX2_X1 U10071 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9678), .Z(n7849) );
  XNOR2_X1 U10072 ( .A(n7850), .B(n7849), .ZN(n10430) );
  NAND2_X1 U10073 ( .A1(n10430), .A2(n8210), .ZN(n7829) );
  NAND2_X1 U10074 ( .A1(n7854), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7827) );
  XNOR2_X1 U10075 ( .A(n7827), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U10076 ( .A1(n8211), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7943), 
        .B2(n11751), .ZN(n7828) );
  NAND2_X1 U10077 ( .A1(n6677), .A2(n8111), .ZN(n7838) );
  INV_X1 U10078 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7830) );
  OR2_X1 U10079 ( .A1(n7419), .A2(n7858), .ZN(n14380) );
  INV_X1 U10080 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11760) );
  OR2_X1 U10081 ( .A1(n8219), .A2(n11760), .ZN(n7834) );
  INV_X1 U10082 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7832) );
  OR2_X1 U10083 ( .A1(n6473), .A2(n7832), .ZN(n7833) );
  AND2_X1 U10084 ( .A1(n7834), .A2(n7833), .ZN(n7836) );
  NAND2_X1 U10085 ( .A1(n8215), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7835) );
  OAI211_X1 U10086 ( .C1(n14380), .C2(n8184), .A(n7836), .B(n7835), .ZN(n13190) );
  NAND2_X1 U10087 ( .A1(n13190), .A2(n8223), .ZN(n7837) );
  NAND2_X1 U10088 ( .A1(n7838), .A2(n7837), .ZN(n7844) );
  NAND2_X1 U10089 ( .A1(n7843), .A2(n7844), .ZN(n7842) );
  NAND2_X1 U10090 ( .A1(n6677), .A2(n8223), .ZN(n7840) );
  NAND2_X1 U10091 ( .A1(n13190), .A2(n8111), .ZN(n7839) );
  NAND2_X1 U10092 ( .A1(n7840), .A2(n7839), .ZN(n7841) );
  NAND2_X1 U10093 ( .A1(n7842), .A2(n7841), .ZN(n7848) );
  INV_X1 U10094 ( .A(n7843), .ZN(n7846) );
  INV_X1 U10095 ( .A(n7844), .ZN(n7845) );
  NAND2_X1 U10096 ( .A1(n7846), .A2(n7845), .ZN(n7847) );
  MUX2_X1 U10097 ( .A(n10536), .B(n10535), .S(n9678), .Z(n7851) );
  INV_X1 U10098 ( .A(n7851), .ZN(n7852) );
  NAND2_X1 U10099 ( .A1(n7852), .A2(SI_15_), .ZN(n7853) );
  XNOR2_X1 U10100 ( .A(n7868), .B(n7867), .ZN(n10534) );
  NAND2_X1 U10101 ( .A1(n10534), .A2(n8210), .ZN(n7857) );
  NOR2_X1 U10102 ( .A1(n7854), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n7875) );
  OR2_X1 U10103 ( .A1(n7875), .A2(n7445), .ZN(n7855) );
  XNOR2_X1 U10104 ( .A(n7855), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14765) );
  AOI22_X1 U10105 ( .A1(n14765), .A2(n7943), .B1(n8211), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n7856) );
  NAND2_X1 U10106 ( .A1(n13546), .A2(n8223), .ZN(n7863) );
  NAND2_X1 U10107 ( .A1(n7858), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7880) );
  OR2_X1 U10108 ( .A1(n7858), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7859) );
  NAND2_X1 U10109 ( .A1(n7880), .A2(n7859), .ZN(n11819) );
  AOI22_X1 U10110 ( .A1(n6475), .A2(P2_REG1_REG_15__SCAN_IN), .B1(n8215), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n7861) );
  NAND2_X1 U10111 ( .A1(n6479), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7860) );
  OAI211_X1 U10112 ( .C1(n11819), .C2(n8184), .A(n7861), .B(n7860), .ZN(n13189) );
  NAND2_X1 U10113 ( .A1(n13189), .A2(n8111), .ZN(n7862) );
  NAND2_X1 U10114 ( .A1(n7863), .A2(n7862), .ZN(n7865) );
  AOI22_X1 U10115 ( .A1(n13546), .A2(n8111), .B1(n8223), .B2(n13189), .ZN(
        n7864) );
  MUX2_X1 U10116 ( .A(n10683), .B(n10682), .S(n9678), .Z(n7871) );
  INV_X1 U10117 ( .A(n7871), .ZN(n7872) );
  NAND2_X1 U10118 ( .A1(n7872), .A2(SI_16_), .ZN(n7873) );
  XNOR2_X1 U10119 ( .A(n7893), .B(n7892), .ZN(n10681) );
  NAND2_X1 U10120 ( .A1(n10681), .A2(n8210), .ZN(n7878) );
  INV_X1 U10121 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7874) );
  NAND2_X1 U10122 ( .A1(n7875), .A2(n7874), .ZN(n7899) );
  NAND2_X1 U10123 ( .A1(n7899), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7876) );
  XNOR2_X1 U10124 ( .A(n7876), .B(P2_IR_REG_16__SCAN_IN), .ZN(n13236) );
  AOI22_X1 U10125 ( .A1(n13236), .A2(n7943), .B1(n8211), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n7877) );
  NAND2_X1 U10126 ( .A1(n14388), .A2(n8111), .ZN(n7885) );
  INV_X1 U10127 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7879) );
  NAND2_X1 U10128 ( .A1(n7880), .A2(n7879), .ZN(n7881) );
  NAND2_X1 U10129 ( .A1(n7903), .A2(n7881), .ZN(n14391) );
  AOI22_X1 U10130 ( .A1(n8215), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n6479), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n7883) );
  NAND2_X1 U10131 ( .A1(n6474), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7882) );
  OAI211_X1 U10132 ( .C1(n14391), .C2(n8068), .A(n7883), .B(n7882), .ZN(n13188) );
  NAND2_X1 U10133 ( .A1(n13188), .A2(n8223), .ZN(n7884) );
  NAND2_X1 U10134 ( .A1(n7885), .A2(n7884), .ZN(n7889) );
  INV_X1 U10135 ( .A(n13188), .ZN(n11840) );
  NAND2_X1 U10136 ( .A1(n14388), .A2(n8223), .ZN(n7886) );
  OAI21_X1 U10137 ( .B1(n11840), .B2(n8223), .A(n7886), .ZN(n7887) );
  NAND2_X1 U10138 ( .A1(n7888), .A2(n7887), .ZN(n7891) );
  NAND2_X1 U10139 ( .A1(n7891), .A2(n7890), .ZN(n7914) );
  INV_X1 U10140 ( .A(n7914), .ZN(n7912) );
  NAND2_X1 U10141 ( .A1(n7893), .A2(n7892), .ZN(n7895) );
  MUX2_X1 U10142 ( .A(n10815), .B(n10814), .S(n9678), .Z(n7896) );
  INV_X1 U10143 ( .A(n7896), .ZN(n7897) );
  NAND2_X1 U10144 ( .A1(n7897), .A2(SI_17_), .ZN(n7898) );
  XNOR2_X1 U10145 ( .A(n7920), .B(n7919), .ZN(n10813) );
  NAND2_X1 U10146 ( .A1(n10813), .A2(n8210), .ZN(n7902) );
  NAND2_X1 U10147 ( .A1(n7922), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7900) );
  XNOR2_X1 U10148 ( .A(n7900), .B(P2_IR_REG_17__SCAN_IN), .ZN(n14777) );
  AOI22_X1 U10149 ( .A1(n14777), .A2(n7943), .B1(n8211), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n7901) );
  NAND2_X1 U10150 ( .A1(n13537), .A2(n8223), .ZN(n7910) );
  AND2_X1 U10151 ( .A1(n7903), .A2(n13117), .ZN(n7904) );
  OR2_X1 U10152 ( .A1(n7904), .A2(n7926), .ZN(n13116) );
  INV_X1 U10153 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11767) );
  NAND2_X1 U10154 ( .A1(n6479), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7906) );
  NAND2_X1 U10155 ( .A1(n8215), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7905) );
  OAI211_X1 U10156 ( .C1(n8219), .C2(n11767), .A(n7906), .B(n7905), .ZN(n7907)
         );
  INV_X1 U10157 ( .A(n7907), .ZN(n7908) );
  OAI21_X1 U10158 ( .B1(n13116), .B2(n8184), .A(n7908), .ZN(n13187) );
  NAND2_X1 U10159 ( .A1(n13187), .A2(n8111), .ZN(n7909) );
  NAND2_X1 U10160 ( .A1(n7910), .A2(n7909), .ZN(n7913) );
  INV_X1 U10161 ( .A(n7913), .ZN(n7911) );
  NAND2_X1 U10162 ( .A1(n7912), .A2(n7911), .ZN(n7918) );
  NAND2_X1 U10163 ( .A1(n7914), .A2(n7913), .ZN(n7917) );
  AOI22_X1 U10164 ( .A1(n13537), .A2(n8111), .B1(n8223), .B2(n13187), .ZN(
        n7915) );
  MUX2_X1 U10165 ( .A(n11107), .B(n11106), .S(n9678), .Z(n7966) );
  NAND2_X1 U10166 ( .A1(n11105), .A2(n8210), .ZN(n7925) );
  OAI21_X1 U10167 ( .B1(n7922), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7923) );
  XNOR2_X1 U10168 ( .A(n7923), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13249) );
  AOI22_X1 U10169 ( .A1(n13249), .A2(n7943), .B1(n8211), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n7924) );
  NAND2_X1 U10170 ( .A1(n13532), .A2(n8111), .ZN(n7934) );
  NOR2_X1 U10171 ( .A1(n7926), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7927) );
  OR2_X1 U10172 ( .A1(n7946), .A2(n7927), .ZN(n13156) );
  INV_X1 U10173 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U10174 ( .A1(n8215), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7929) );
  NAND2_X1 U10175 ( .A1(n6479), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7928) );
  OAI211_X1 U10176 ( .C1(n7930), .C2(n8219), .A(n7929), .B(n7928), .ZN(n7931)
         );
  INV_X1 U10177 ( .A(n7931), .ZN(n7932) );
  OAI21_X1 U10178 ( .B1(n13156), .B2(n8184), .A(n7932), .ZN(n13186) );
  NAND2_X1 U10179 ( .A1(n13186), .A2(n8223), .ZN(n7933) );
  NAND2_X1 U10180 ( .A1(n7934), .A2(n7933), .ZN(n7936) );
  AOI22_X1 U10181 ( .A1(n13532), .A2(n8223), .B1(n13186), .B2(n8111), .ZN(
        n7935) );
  INV_X1 U10182 ( .A(n7966), .ZN(n7970) );
  NOR2_X1 U10183 ( .A1(n7969), .A2(n15126), .ZN(n7937) );
  AOI21_X1 U10184 ( .B1(n7938), .B2(n7970), .A(n7937), .ZN(n7942) );
  MUX2_X1 U10185 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9678), .Z(n7939) );
  NAND2_X1 U10186 ( .A1(n7939), .A2(SI_19_), .ZN(n7973) );
  INV_X1 U10187 ( .A(n7939), .ZN(n7940) );
  INV_X1 U10188 ( .A(SI_19_), .ZN(n10154) );
  NAND2_X1 U10189 ( .A1(n7940), .A2(n10154), .ZN(n7971) );
  AND2_X1 U10190 ( .A1(n7973), .A2(n7971), .ZN(n7941) );
  XNOR2_X1 U10191 ( .A(n7942), .B(n7941), .ZN(n11161) );
  NAND2_X1 U10192 ( .A1(n11161), .A2(n8210), .ZN(n7945) );
  AOI22_X1 U10193 ( .A1(n8211), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7943), 
        .B2(n10332), .ZN(n7944) );
  NAND2_X1 U10194 ( .A1(n13528), .A2(n8223), .ZN(n7955) );
  OR2_X1 U10195 ( .A1(n7946), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n7947) );
  AND2_X1 U10196 ( .A1(n7996), .A2(n7947), .ZN(n13423) );
  NAND2_X1 U10197 ( .A1(n13423), .A2(n7592), .ZN(n7953) );
  INV_X1 U10198 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n7950) );
  NAND2_X1 U10199 ( .A1(n6479), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n7949) );
  NAND2_X1 U10200 ( .A1(n8215), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n7948) );
  OAI211_X1 U10201 ( .C1(n8219), .C2(n7950), .A(n7949), .B(n7948), .ZN(n7951)
         );
  INV_X1 U10202 ( .A(n7951), .ZN(n7952) );
  NAND2_X1 U10203 ( .A1(n7953), .A2(n7952), .ZN(n13185) );
  NAND2_X1 U10204 ( .A1(n13185), .A2(n8111), .ZN(n7954) );
  NAND2_X1 U10205 ( .A1(n7955), .A2(n7954), .ZN(n7961) );
  NAND2_X1 U10206 ( .A1(n7960), .A2(n7961), .ZN(n7959) );
  NAND2_X1 U10207 ( .A1(n13528), .A2(n8111), .ZN(n7957) );
  NAND2_X1 U10208 ( .A1(n13185), .A2(n8223), .ZN(n7956) );
  NAND2_X1 U10209 ( .A1(n7957), .A2(n7956), .ZN(n7958) );
  NAND2_X1 U10210 ( .A1(n7959), .A2(n7958), .ZN(n7965) );
  INV_X1 U10211 ( .A(n7960), .ZN(n7963) );
  INV_X1 U10212 ( .A(n7961), .ZN(n7962) );
  NAND2_X1 U10213 ( .A1(n7963), .A2(n7962), .ZN(n7964) );
  OAI21_X1 U10214 ( .B1(n15126), .B2(n7966), .A(n7973), .ZN(n7967) );
  INV_X1 U10215 ( .A(n7967), .ZN(n7968) );
  NOR2_X1 U10216 ( .A1(n7970), .A2(SI_18_), .ZN(n7974) );
  INV_X1 U10217 ( .A(n7971), .ZN(n7972) );
  AOI21_X1 U10218 ( .B1(n7974), .B2(n7973), .A(n7972), .ZN(n7975) );
  XNOR2_X1 U10219 ( .A(n8021), .B(n15090), .ZN(n7987) );
  MUX2_X1 U10220 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n9678), .Z(n8016) );
  XNOR2_X1 U10221 ( .A(n7987), .B(n8016), .ZN(n11166) );
  NAND2_X1 U10222 ( .A1(n11166), .A2(n8210), .ZN(n7977) );
  NAND2_X1 U10223 ( .A1(n8211), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7976) );
  NAND2_X1 U10224 ( .A1(n13523), .A2(n8111), .ZN(n7985) );
  XNOR2_X1 U10225 ( .A(n7996), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n13415) );
  NAND2_X1 U10226 ( .A1(n13415), .A2(n7592), .ZN(n7983) );
  INV_X1 U10227 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n7980) );
  NAND2_X1 U10228 ( .A1(n6479), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n7979) );
  NAND2_X1 U10229 ( .A1(n8215), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n7978) );
  OAI211_X1 U10230 ( .C1(n8219), .C2(n7980), .A(n7979), .B(n7978), .ZN(n7981)
         );
  INV_X1 U10231 ( .A(n7981), .ZN(n7982) );
  NAND2_X1 U10232 ( .A1(n7983), .A2(n7982), .ZN(n13184) );
  NAND2_X1 U10233 ( .A1(n13184), .A2(n8223), .ZN(n7984) );
  AOI22_X1 U10234 ( .A1(n13523), .A2(n8223), .B1(n13184), .B2(n8111), .ZN(
        n7986) );
  INV_X1 U10235 ( .A(n7987), .ZN(n7988) );
  NAND2_X1 U10236 ( .A1(n7988), .A2(n8016), .ZN(n7990) );
  OR2_X1 U10237 ( .A1(n8021), .A2(n15090), .ZN(n7989) );
  NAND2_X1 U10238 ( .A1(n7990), .A2(n7989), .ZN(n7992) );
  MUX2_X1 U10239 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9678), .Z(n8018) );
  XNOR2_X1 U10240 ( .A(n8018), .B(SI_21_), .ZN(n7991) );
  NAND2_X1 U10241 ( .A1(n11256), .A2(n8210), .ZN(n7994) );
  NAND2_X1 U10242 ( .A1(n8211), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7993) );
  NAND2_X1 U10243 ( .A1(n13518), .A2(n8223), .ZN(n8005) );
  INV_X1 U10244 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13137) );
  INV_X1 U10245 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13100) );
  OAI21_X1 U10246 ( .B1(n7996), .B2(n13137), .A(n13100), .ZN(n7997) );
  NAND2_X1 U10247 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n7995) );
  NAND2_X1 U10248 ( .A1(n7997), .A2(n8025), .ZN(n13099) );
  OR2_X1 U10249 ( .A1(n13099), .A2(n8068), .ZN(n8003) );
  INV_X1 U10250 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8000) );
  NAND2_X1 U10251 ( .A1(n6479), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U10252 ( .A1(n8215), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7998) );
  OAI211_X1 U10253 ( .C1(n8219), .C2(n8000), .A(n7999), .B(n7998), .ZN(n8001)
         );
  INV_X1 U10254 ( .A(n8001), .ZN(n8002) );
  NAND2_X1 U10255 ( .A1(n8003), .A2(n8002), .ZN(n13183) );
  NAND2_X1 U10256 ( .A1(n13183), .A2(n8111), .ZN(n8004) );
  NAND2_X1 U10257 ( .A1(n8005), .A2(n8004), .ZN(n8011) );
  NAND2_X1 U10258 ( .A1(n8010), .A2(n8011), .ZN(n8009) );
  NAND2_X1 U10259 ( .A1(n13518), .A2(n8111), .ZN(n8007) );
  NAND2_X1 U10260 ( .A1(n13183), .A2(n8223), .ZN(n8006) );
  NAND2_X1 U10261 ( .A1(n8007), .A2(n8006), .ZN(n8008) );
  NAND2_X1 U10262 ( .A1(n8009), .A2(n8008), .ZN(n8015) );
  INV_X1 U10263 ( .A(n8010), .ZN(n8013) );
  INV_X1 U10264 ( .A(n8011), .ZN(n8012) );
  NAND2_X1 U10265 ( .A1(n8013), .A2(n8012), .ZN(n8014) );
  NAND2_X1 U10266 ( .A1(n8015), .A2(n8014), .ZN(n8037) );
  INV_X1 U10267 ( .A(n8016), .ZN(n8017) );
  NOR2_X1 U10268 ( .A1(n8017), .A2(n15090), .ZN(n8019) );
  AOI22_X1 U10269 ( .A1(n8019), .A2(n7424), .B1(n8018), .B2(SI_21_), .ZN(n8020) );
  MUX2_X1 U10270 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9678), .Z(n8038) );
  XNOR2_X1 U10271 ( .A(n9461), .B(n8038), .ZN(n11455) );
  NAND2_X1 U10272 ( .A1(n11455), .A2(n8210), .ZN(n8023) );
  NAND2_X1 U10273 ( .A1(n8211), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8022) );
  NAND2_X1 U10274 ( .A1(n13511), .A2(n8111), .ZN(n8033) );
  INV_X1 U10275 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8024) );
  AND2_X1 U10276 ( .A1(n8025), .A2(n8024), .ZN(n8026) );
  OR2_X1 U10277 ( .A1(n8026), .A2(n8044), .ZN(n13386) );
  INV_X1 U10278 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8029) );
  NAND2_X1 U10279 ( .A1(n6479), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8028) );
  NAND2_X1 U10280 ( .A1(n8215), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8027) );
  OAI211_X1 U10281 ( .C1(n8219), .C2(n8029), .A(n8028), .B(n8027), .ZN(n8030)
         );
  INV_X1 U10282 ( .A(n8030), .ZN(n8031) );
  OAI21_X1 U10283 ( .B1(n13386), .B2(n8184), .A(n8031), .ZN(n13182) );
  NAND2_X1 U10284 ( .A1(n13182), .A2(n8223), .ZN(n8032) );
  NAND2_X1 U10285 ( .A1(n8033), .A2(n8032), .ZN(n8036) );
  AOI22_X1 U10286 ( .A1(n13511), .A2(n8223), .B1(n13182), .B2(n8111), .ZN(
        n8035) );
  INV_X1 U10287 ( .A(n8038), .ZN(n8041) );
  NAND2_X1 U10288 ( .A1(n8039), .A2(SI_22_), .ZN(n8040) );
  MUX2_X1 U10289 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9678), .Z(n8061) );
  XNOR2_X1 U10290 ( .A(n8061), .B(SI_23_), .ZN(n8058) );
  XNOR2_X1 U10291 ( .A(n8060), .B(n8058), .ZN(n11529) );
  NAND2_X1 U10292 ( .A1(n11529), .A2(n8210), .ZN(n8043) );
  NAND2_X1 U10293 ( .A1(n8211), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8042) );
  NAND2_X1 U10294 ( .A1(n13505), .A2(n8223), .ZN(n8053) );
  OR2_X1 U10295 ( .A1(n8044), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8045) );
  NAND2_X1 U10296 ( .A1(n8044), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8066) );
  NAND2_X1 U10297 ( .A1(n8045), .A2(n8066), .ZN(n13370) );
  OR2_X1 U10298 ( .A1(n13370), .A2(n8068), .ZN(n8051) );
  INV_X1 U10299 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8048) );
  NAND2_X1 U10300 ( .A1(n6479), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8047) );
  NAND2_X1 U10301 ( .A1(n8215), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8046) );
  OAI211_X1 U10302 ( .C1(n8219), .C2(n8048), .A(n8047), .B(n8046), .ZN(n8049)
         );
  INV_X1 U10303 ( .A(n8049), .ZN(n8050) );
  NAND2_X1 U10304 ( .A1(n8051), .A2(n8050), .ZN(n13181) );
  NAND2_X1 U10305 ( .A1(n13181), .A2(n8111), .ZN(n8052) );
  NAND2_X1 U10306 ( .A1(n8053), .A2(n8052), .ZN(n8056) );
  INV_X1 U10307 ( .A(n13181), .ZN(n13145) );
  NAND2_X1 U10308 ( .A1(n13505), .A2(n8111), .ZN(n8054) );
  OAI21_X1 U10309 ( .B1(n13145), .B2(n8111), .A(n8054), .ZN(n8055) );
  INV_X1 U10310 ( .A(n8055), .ZN(n8057) );
  INV_X1 U10311 ( .A(n8058), .ZN(n8059) );
  NAND2_X1 U10312 ( .A1(n8061), .A2(SI_23_), .ZN(n8062) );
  MUX2_X1 U10313 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9678), .Z(n8078) );
  XNOR2_X1 U10314 ( .A(n8077), .B(n8078), .ZN(n11775) );
  NAND2_X1 U10315 ( .A1(n11775), .A2(n8210), .ZN(n8065) );
  NAND2_X1 U10316 ( .A1(n8211), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8064) );
  NAND2_X1 U10317 ( .A1(n13496), .A2(n8111), .ZN(n8074) );
  OAI21_X1 U10318 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n8067), .A(n8101), .ZN(
        n13352) );
  OR2_X1 U10319 ( .A1(n8068), .A2(n13352), .ZN(n8072) );
  NAND2_X1 U10320 ( .A1(n6475), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8071) );
  INV_X1 U10321 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13353) );
  OR2_X1 U10322 ( .A1(n8185), .A2(n13353), .ZN(n8070) );
  INV_X1 U10323 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n13565) );
  OR2_X1 U10324 ( .A1(n8187), .A2(n13565), .ZN(n8069) );
  NAND4_X1 U10325 ( .A1(n8072), .A2(n8071), .A3(n8070), .A4(n8069), .ZN(n13180) );
  NAND2_X1 U10326 ( .A1(n13180), .A2(n8223), .ZN(n8073) );
  NAND2_X1 U10327 ( .A1(n8074), .A2(n8073), .ZN(n8076) );
  AOI22_X1 U10328 ( .A1(n13496), .A2(n8223), .B1(n13180), .B2(n8111), .ZN(
        n8075) );
  NAND2_X1 U10329 ( .A1(n8079), .A2(SI_24_), .ZN(n8080) );
  INV_X1 U10330 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11859) );
  INV_X1 U10331 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11863) );
  MUX2_X1 U10332 ( .A(n11859), .B(n11863), .S(n9678), .Z(n8081) );
  INV_X1 U10333 ( .A(SI_25_), .ZN(n15169) );
  NAND2_X1 U10334 ( .A1(n8081), .A2(n15169), .ZN(n8094) );
  INV_X1 U10335 ( .A(n8081), .ZN(n8082) );
  NAND2_X1 U10336 ( .A1(n8082), .A2(SI_25_), .ZN(n8083) );
  NAND2_X1 U10337 ( .A1(n8094), .A2(n8083), .ZN(n8095) );
  XNOR2_X1 U10338 ( .A(n8096), .B(n8095), .ZN(n11858) );
  NAND2_X1 U10339 ( .A1(n11858), .A2(n8210), .ZN(n8085) );
  NAND2_X1 U10340 ( .A1(n8211), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8084) );
  INV_X1 U10341 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13107) );
  XNOR2_X1 U10342 ( .A(n8101), .B(n13107), .ZN(n13332) );
  OR2_X1 U10343 ( .A1(n8184), .A2(n13332), .ZN(n8090) );
  NAND2_X1 U10344 ( .A1(n6474), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8089) );
  INV_X1 U10345 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13333) );
  OR2_X1 U10346 ( .A1(n8185), .A2(n13333), .ZN(n8088) );
  INV_X1 U10347 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8086) );
  OR2_X1 U10348 ( .A1(n8187), .A2(n8086), .ZN(n8087) );
  NAND4_X1 U10349 ( .A1(n8090), .A2(n8089), .A3(n8088), .A4(n8087), .ZN(n13179) );
  AND2_X1 U10350 ( .A1(n13179), .A2(n8223), .ZN(n8091) );
  AOI21_X1 U10351 ( .B1(n13335), .B2(n8111), .A(n8091), .ZN(n8115) );
  NAND2_X1 U10352 ( .A1(n13335), .A2(n8223), .ZN(n8093) );
  NAND2_X1 U10353 ( .A1(n13179), .A2(n8111), .ZN(n8092) );
  NAND2_X1 U10354 ( .A1(n8093), .A2(n8092), .ZN(n8114) );
  INV_X1 U10355 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13594) );
  MUX2_X1 U10356 ( .A(n14186), .B(n13594), .S(n9678), .Z(n8118) );
  XNOR2_X1 U10357 ( .A(n8118), .B(SI_26_), .ZN(n8097) );
  XNOR2_X1 U10358 ( .A(n8119), .B(n8097), .ZN(n13592) );
  NAND2_X1 U10359 ( .A1(n13592), .A2(n8210), .ZN(n8099) );
  NAND2_X1 U10360 ( .A1(n8211), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8098) );
  INV_X1 U10361 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8100) );
  OAI21_X1 U10362 ( .B1(n8101), .B2(n13107), .A(n8100), .ZN(n8104) );
  INV_X1 U10363 ( .A(n8101), .ZN(n8103) );
  AND2_X1 U10364 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n8102) );
  NAND2_X1 U10365 ( .A1(n8103), .A2(n8102), .ZN(n8181) );
  NAND2_X1 U10366 ( .A1(n8104), .A2(n8181), .ZN(n13313) );
  OR2_X1 U10367 ( .A1(n8184), .A2(n13313), .ZN(n8109) );
  NAND2_X1 U10368 ( .A1(n6474), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8108) );
  INV_X1 U10369 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13314) );
  OR2_X1 U10370 ( .A1(n8185), .A2(n13314), .ZN(n8107) );
  INV_X1 U10371 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8105) );
  OR2_X1 U10372 ( .A1(n6473), .A2(n8105), .ZN(n8106) );
  NAND4_X1 U10373 ( .A1(n8109), .A2(n8108), .A3(n8107), .A4(n8106), .ZN(n13178) );
  AND2_X1 U10374 ( .A1(n13178), .A2(n8223), .ZN(n8110) );
  AOI21_X1 U10375 ( .B1(n13487), .B2(n8111), .A(n8110), .ZN(n8196) );
  NAND2_X1 U10376 ( .A1(n13487), .A2(n8223), .ZN(n8113) );
  NAND2_X1 U10377 ( .A1(n13178), .A2(n8111), .ZN(n8112) );
  NAND2_X1 U10378 ( .A1(n8113), .A2(n8112), .ZN(n8195) );
  AOI22_X1 U10379 ( .A1(n8196), .A2(n8195), .B1(n8115), .B2(n8114), .ZN(n8116)
         );
  NAND2_X1 U10380 ( .A1(n8117), .A2(n8116), .ZN(n8233) );
  NAND2_X1 U10381 ( .A1(n8119), .A2(n15171), .ZN(n8120) );
  MUX2_X1 U10382 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9678), .Z(n8175) );
  MUX2_X1 U10383 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n6478), .Z(n8124) );
  XNOR2_X1 U10384 ( .A(n8124), .B(SI_28_), .ZN(n8159) );
  INV_X1 U10385 ( .A(n8159), .ZN(n8122) );
  NAND2_X1 U10386 ( .A1(n8175), .A2(SI_27_), .ZN(n8157) );
  AND2_X1 U10387 ( .A1(n8122), .A2(n8157), .ZN(n8123) );
  INV_X1 U10388 ( .A(n8124), .ZN(n8125) );
  INV_X1 U10389 ( .A(SI_28_), .ZN(n13069) );
  NAND2_X1 U10390 ( .A1(n8125), .A2(n13069), .ZN(n8126) );
  MUX2_X1 U10391 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n9678), .Z(n8128) );
  XNOR2_X1 U10392 ( .A(n8128), .B(n11869), .ZN(n8143) );
  INV_X1 U10393 ( .A(n8128), .ZN(n8129) );
  MUX2_X1 U10394 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6478), .Z(n8130) );
  XNOR2_X1 U10395 ( .A(n8130), .B(SI_30_), .ZN(n8209) );
  INV_X1 U10396 ( .A(n8130), .ZN(n8131) );
  INV_X1 U10397 ( .A(SI_30_), .ZN(n15145) );
  MUX2_X1 U10398 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9678), .Z(n8132) );
  XNOR2_X1 U10399 ( .A(n8132), .B(SI_31_), .ZN(n8133) );
  XNOR2_X1 U10400 ( .A(n8134), .B(n8133), .ZN(n9563) );
  NAND2_X1 U10401 ( .A1(n9563), .A2(n8210), .ZN(n8136) );
  NAND2_X1 U10402 ( .A1(n8211), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8135) );
  INV_X1 U10403 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8139) );
  NAND2_X1 U10404 ( .A1(n8215), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8138) );
  NAND2_X1 U10405 ( .A1(n6479), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8137) );
  OAI211_X1 U10406 ( .C1(n8219), .C2(n8139), .A(n8138), .B(n8137), .ZN(n13265)
         );
  NAND2_X1 U10407 ( .A1(n13263), .A2(n13265), .ZN(n8142) );
  NAND2_X1 U10408 ( .A1(n8236), .A2(n8142), .ZN(n8257) );
  NAND2_X1 U10409 ( .A1(n11864), .A2(n8210), .ZN(n8146) );
  NAND2_X1 U10410 ( .A1(n8211), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8145) );
  INV_X1 U10411 ( .A(n8181), .ZN(n8147) );
  NAND2_X1 U10412 ( .A1(n8147), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8183) );
  INV_X1 U10413 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8163) );
  OR2_X1 U10414 ( .A1(n8184), .A2(n12016), .ZN(n8153) );
  NAND2_X1 U10415 ( .A1(n6474), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8152) );
  INV_X1 U10416 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8148) );
  OR2_X1 U10417 ( .A1(n8185), .A2(n8148), .ZN(n8151) );
  INV_X1 U10418 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8149) );
  OR2_X1 U10419 ( .A1(n6473), .A2(n8149), .ZN(n8150) );
  NAND4_X1 U10420 ( .A1(n8153), .A2(n8152), .A3(n8151), .A4(n8150), .ZN(n13175) );
  AND2_X1 U10421 ( .A1(n13175), .A2(n8111), .ZN(n8154) );
  AOI21_X1 U10422 ( .B1(n13471), .B2(n8223), .A(n8154), .ZN(n8227) );
  NAND2_X1 U10423 ( .A1(n13471), .A2(n8111), .ZN(n8156) );
  NAND2_X1 U10424 ( .A1(n13175), .A2(n8223), .ZN(n8155) );
  NAND2_X1 U10425 ( .A1(n8156), .A2(n8155), .ZN(n8226) );
  NAND2_X1 U10426 ( .A1(n8227), .A2(n8226), .ZN(n8205) );
  NAND2_X1 U10427 ( .A1(n8158), .A2(n8157), .ZN(n8160) );
  NAND2_X1 U10428 ( .A1(n12032), .A2(n8210), .ZN(n8162) );
  NAND2_X1 U10429 ( .A1(n8211), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8161) );
  NAND2_X1 U10430 ( .A1(n8183), .A2(n8163), .ZN(n8164) );
  NAND2_X1 U10431 ( .A1(n12016), .A2(n8164), .ZN(n13285) );
  OR2_X1 U10432 ( .A1(n8184), .A2(n13285), .ZN(n8169) );
  NAND2_X1 U10433 ( .A1(n6475), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8168) );
  INV_X1 U10434 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13286) );
  OR2_X1 U10435 ( .A1(n8185), .A2(n13286), .ZN(n8167) );
  INV_X1 U10436 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8165) );
  OR2_X1 U10437 ( .A1(n8187), .A2(n8165), .ZN(n8166) );
  NAND4_X1 U10438 ( .A1(n8169), .A2(n8168), .A3(n8167), .A4(n8166), .ZN(n13176) );
  AND2_X1 U10439 ( .A1(n13176), .A2(n8111), .ZN(n8170) );
  AOI21_X1 U10440 ( .B1(n13475), .B2(n8223), .A(n8170), .ZN(n8203) );
  NAND2_X1 U10441 ( .A1(n13475), .A2(n8111), .ZN(n8172) );
  NAND2_X1 U10442 ( .A1(n13176), .A2(n8223), .ZN(n8171) );
  NAND2_X1 U10443 ( .A1(n8172), .A2(n8171), .ZN(n8202) );
  NAND2_X1 U10444 ( .A1(n8203), .A2(n8202), .ZN(n8173) );
  AND2_X1 U10445 ( .A1(n8205), .A2(n8173), .ZN(n8174) );
  INV_X1 U10446 ( .A(n8175), .ZN(n8176) );
  XNOR2_X1 U10447 ( .A(n8176), .B(SI_27_), .ZN(n8177) );
  NAND2_X1 U10448 ( .A1(n13589), .A2(n8210), .ZN(n8180) );
  NAND2_X1 U10449 ( .A1(n8211), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8179) );
  INV_X1 U10450 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13074) );
  NAND2_X1 U10451 ( .A1(n8181), .A2(n13074), .ZN(n8182) );
  NAND2_X1 U10452 ( .A1(n8183), .A2(n8182), .ZN(n13301) );
  OR2_X1 U10453 ( .A1(n8184), .A2(n13301), .ZN(n8191) );
  NAND2_X1 U10454 ( .A1(n6475), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8190) );
  INV_X1 U10455 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13302) );
  OR2_X1 U10456 ( .A1(n8185), .A2(n13302), .ZN(n8189) );
  INV_X1 U10457 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8186) );
  OR2_X1 U10458 ( .A1(n6473), .A2(n8186), .ZN(n8188) );
  NAND4_X1 U10459 ( .A1(n8191), .A2(n8190), .A3(n8189), .A4(n8188), .ZN(n13177) );
  AND2_X1 U10460 ( .A1(n13177), .A2(n8111), .ZN(n8192) );
  AOI21_X1 U10461 ( .B1(n13304), .B2(n8223), .A(n8192), .ZN(n8201) );
  NAND2_X1 U10462 ( .A1(n13304), .A2(n8111), .ZN(n8194) );
  NAND2_X1 U10463 ( .A1(n13177), .A2(n8223), .ZN(n8193) );
  NAND2_X1 U10464 ( .A1(n8194), .A2(n8193), .ZN(n8200) );
  INV_X1 U10465 ( .A(n8195), .ZN(n8198) );
  INV_X1 U10466 ( .A(n8196), .ZN(n8197) );
  AOI22_X1 U10467 ( .A1(n8201), .A2(n8200), .B1(n8198), .B2(n8197), .ZN(n8199)
         );
  INV_X1 U10468 ( .A(n8202), .ZN(n8206) );
  INV_X1 U10469 ( .A(n8203), .ZN(n8204) );
  NAND4_X1 U10470 ( .A1(n8257), .A2(n8206), .A3(n8205), .A4(n8204), .ZN(n8231)
         );
  NAND2_X1 U10471 ( .A1(n13265), .A2(n8223), .ZN(n8207) );
  OAI211_X1 U10472 ( .C1(n8141), .C2(n8223), .A(n8207), .B(n8236), .ZN(n8229)
         );
  NAND2_X1 U10473 ( .A1(n12159), .A2(n8210), .ZN(n8213) );
  NAND2_X1 U10474 ( .A1(n8211), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8212) );
  NAND2_X1 U10475 ( .A1(n13265), .A2(n8111), .ZN(n8237) );
  NAND2_X1 U10476 ( .A1(n10338), .A2(n6477), .ZN(n8262) );
  NAND2_X1 U10477 ( .A1(n13257), .A2(n11228), .ZN(n10077) );
  NAND4_X1 U10478 ( .A1(n8237), .A2(n10076), .A3(n8262), .A4(n10077), .ZN(
        n8220) );
  INV_X1 U10479 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8218) );
  NAND2_X1 U10480 ( .A1(n8215), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8217) );
  NAND2_X1 U10481 ( .A1(n6479), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8216) );
  OAI211_X1 U10482 ( .C1(n8219), .C2(n8218), .A(n8217), .B(n8216), .ZN(n13174)
         );
  AND2_X1 U10483 ( .A1(n8220), .A2(n13174), .ZN(n8221) );
  AOI21_X1 U10484 ( .B1(n13269), .B2(n8223), .A(n8221), .ZN(n8235) );
  NAND2_X1 U10485 ( .A1(n13269), .A2(n8111), .ZN(n8225) );
  NAND2_X1 U10486 ( .A1(n13174), .A2(n8223), .ZN(n8224) );
  NAND2_X1 U10487 ( .A1(n8225), .A2(n8224), .ZN(n8234) );
  OAI22_X1 U10488 ( .A1(n8235), .A2(n8234), .B1(n8227), .B2(n8226), .ZN(n8228)
         );
  NAND2_X1 U10489 ( .A1(n8229), .A2(n8228), .ZN(n8230) );
  AOI21_X1 U10490 ( .B1(n8233), .B2(n7412), .A(n8232), .ZN(n8239) );
  OAI211_X1 U10491 ( .C1(n8141), .C2(n8111), .A(n8237), .B(n8236), .ZN(n8238)
         );
  INV_X1 U10492 ( .A(n13178), .ZN(n12007) );
  XNOR2_X1 U10493 ( .A(n13487), .B(n12007), .ZN(n12008) );
  XNOR2_X1 U10494 ( .A(n13335), .B(n13179), .ZN(n12006) );
  INV_X1 U10495 ( .A(n13182), .ZN(n13082) );
  XNOR2_X1 U10496 ( .A(n13511), .B(n13082), .ZN(n11985) );
  INV_X1 U10497 ( .A(n13183), .ZN(n13143) );
  XNOR2_X1 U10498 ( .A(n13518), .B(n13143), .ZN(n13395) );
  XNOR2_X1 U10499 ( .A(n13528), .B(n13185), .ZN(n13427) );
  XNOR2_X1 U10500 ( .A(n14388), .B(n11840), .ZN(n11656) );
  INV_X1 U10501 ( .A(n13189), .ZN(n11659) );
  XNOR2_X1 U10502 ( .A(n13546), .B(n11659), .ZN(n11645) );
  INV_X1 U10503 ( .A(n13190), .ZN(n11779) );
  XNOR2_X1 U10504 ( .A(n14377), .B(n11779), .ZN(n11340) );
  OR2_X1 U10505 ( .A1(n11290), .A2(n13192), .ZN(n11297) );
  NAND2_X1 U10506 ( .A1(n11290), .A2(n13192), .ZN(n11295) );
  NAND2_X1 U10507 ( .A1(n11297), .A2(n11295), .ZN(n11186) );
  XNOR2_X1 U10508 ( .A(n14670), .B(n13191), .ZN(n11298) );
  XNOR2_X1 U10509 ( .A(n10887), .B(n13195), .ZN(n10731) );
  NAND2_X1 U10510 ( .A1(n10570), .A2(n13199), .ZN(n8240) );
  INV_X1 U10511 ( .A(n13199), .ZN(n10569) );
  NAND2_X1 U10512 ( .A1(n14808), .A2(n10569), .ZN(n10576) );
  NAND2_X1 U10513 ( .A1(n8240), .A2(n10576), .ZN(n10553) );
  INV_X1 U10514 ( .A(n14802), .ZN(n10605) );
  INV_X1 U10515 ( .A(n13200), .ZN(n10548) );
  NAND2_X1 U10516 ( .A1(n10605), .A2(n10548), .ZN(n10542) );
  NAND2_X1 U10517 ( .A1(n14802), .A2(n13200), .ZN(n8241) );
  INV_X1 U10518 ( .A(n11228), .ZN(n10560) );
  INV_X1 U10519 ( .A(n8242), .ZN(n8243) );
  NOR2_X1 U10520 ( .A1(n8243), .A2(n10070), .ZN(n14798) );
  NAND4_X1 U10521 ( .A1(n10162), .A2(n6471), .A3(n10560), .A4(n14798), .ZN(
        n8244) );
  NOR4_X1 U10522 ( .A1(n10553), .A2(n10167), .A3(n10608), .A4(n8244), .ZN(
        n8245) );
  XNOR2_X1 U10523 ( .A(n10665), .B(n13197), .ZN(n10773) );
  NAND4_X1 U10524 ( .A1(n10731), .A2(n8245), .A3(n10773), .A4(n7063), .ZN(
        n8248) );
  XNOR2_X1 U10525 ( .A(n10790), .B(n10729), .ZN(n10723) );
  NAND2_X1 U10526 ( .A1(n11072), .A2(n8246), .ZN(n11075) );
  OR2_X1 U10527 ( .A1(n11072), .A2(n8246), .ZN(n8247) );
  NAND2_X1 U10528 ( .A1(n11075), .A2(n8247), .ZN(n11070) );
  NOR3_X1 U10529 ( .A1(n8248), .A2(n10723), .A3(n11070), .ZN(n8249) );
  XNOR2_X1 U10530 ( .A(n11183), .B(n13193), .ZN(n11077) );
  NAND4_X1 U10531 ( .A1(n11186), .A2(n11298), .A3(n8249), .A4(n11077), .ZN(
        n8250) );
  NOR4_X1 U10532 ( .A1(n11656), .A2(n11645), .A3(n11340), .A4(n8250), .ZN(
        n8251) );
  XNOR2_X1 U10533 ( .A(n13532), .B(n13186), .ZN(n13448) );
  XNOR2_X1 U10534 ( .A(n13537), .B(n13187), .ZN(n11839) );
  NAND4_X1 U10535 ( .A1(n13427), .A2(n8251), .A3(n13448), .A4(n11839), .ZN(
        n8252) );
  INV_X1 U10536 ( .A(n13184), .ZN(n11983) );
  XNOR2_X1 U10537 ( .A(n13523), .B(n11983), .ZN(n13408) );
  NOR4_X1 U10538 ( .A1(n11985), .A2(n13395), .A3(n8252), .A4(n13408), .ZN(
        n8253) );
  XNOR2_X1 U10539 ( .A(n13496), .B(n13180), .ZN(n13340) );
  XNOR2_X1 U10540 ( .A(n13505), .B(n13181), .ZN(n13362) );
  NAND4_X1 U10541 ( .A1(n12006), .A2(n8253), .A3(n13340), .A4(n13362), .ZN(
        n8254) );
  NOR4_X1 U10542 ( .A1(n13299), .A2(n13283), .A3(n12008), .A4(n8254), .ZN(
        n8256) );
  XNOR2_X1 U10543 ( .A(n13269), .B(n13174), .ZN(n8255) );
  XNOR2_X1 U10544 ( .A(n13471), .B(n13175), .ZN(n12012) );
  NAND4_X1 U10545 ( .A1(n8257), .A2(n8256), .A3(n8255), .A4(n12012), .ZN(n8258) );
  XNOR2_X1 U10546 ( .A(n8258), .B(n13257), .ZN(n8259) );
  INV_X1 U10547 ( .A(n10067), .ZN(n8260) );
  OAI211_X1 U10548 ( .C1(n10332), .C2(n11257), .A(n8260), .B(n10077), .ZN(
        n8261) );
  INV_X1 U10549 ( .A(n8261), .ZN(n8264) );
  NAND2_X1 U10550 ( .A1(n10076), .A2(n10560), .ZN(n10072) );
  OAI21_X1 U10551 ( .B1(n10072), .B2(n13257), .A(n8262), .ZN(n8263) );
  INV_X1 U10552 ( .A(n8271), .ZN(n8267) );
  NAND2_X1 U10553 ( .A1(n8267), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8268) );
  INV_X4 U10554 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  OR2_X1 U10555 ( .A1(n9818), .A2(P2_U3088), .ZN(n11526) );
  INV_X1 U10556 ( .A(n11526), .ZN(n8269) );
  NAND2_X1 U10557 ( .A1(n8271), .A2(n8270), .ZN(n8273) );
  NAND2_X1 U10558 ( .A1(n8273), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8272) );
  MUX2_X1 U10559 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8272), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8274) );
  NAND2_X1 U10560 ( .A1(n8274), .A2(n8277), .ZN(n11776) );
  INV_X1 U10561 ( .A(n11776), .ZN(n8276) );
  NAND2_X1 U10562 ( .A1(n8277), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8275) );
  NAND2_X1 U10563 ( .A1(n8276), .A2(n10044), .ZN(n8280) );
  INV_X1 U10564 ( .A(n13590), .ZN(n11991) );
  INV_X1 U10565 ( .A(n10077), .ZN(n10126) );
  INV_X1 U10566 ( .A(n8281), .ZN(n8282) );
  NAND4_X1 U10567 ( .A1(n14795), .A2(n11991), .A3(n10126), .A4(n13166), .ZN(
        n8283) );
  OAI211_X1 U10568 ( .C1(n6477), .C2(n11526), .A(n8283), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8284) );
  XNOR2_X1 U10569 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8404) );
  INV_X1 U10570 ( .A(n8403), .ZN(n8286) );
  INV_X1 U10571 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9711) );
  NAND2_X1 U10572 ( .A1(n9711), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8287) );
  NAND2_X1 U10573 ( .A1(n9676), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8289) );
  NAND2_X1 U10574 ( .A1(n9674), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8288) );
  AND2_X1 U10575 ( .A1(n8289), .A2(n8288), .ZN(n8414) );
  NAND2_X1 U10576 ( .A1(n9687), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8292) );
  INV_X1 U10577 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9684) );
  NAND2_X1 U10578 ( .A1(n9684), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8290) );
  NAND2_X1 U10579 ( .A1(n8292), .A2(n8290), .ZN(n8425) );
  INV_X1 U10580 ( .A(n8425), .ZN(n8291) );
  NAND2_X1 U10581 ( .A1(n9690), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8294) );
  INV_X1 U10582 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9688) );
  NAND2_X1 U10583 ( .A1(n9688), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8293) );
  NAND2_X1 U10584 ( .A1(n8295), .A2(n8294), .ZN(n8451) );
  NAND2_X1 U10585 ( .A1(n9719), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8297) );
  INV_X1 U10586 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9718) );
  NAND2_X1 U10587 ( .A1(n9718), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8296) );
  NAND2_X1 U10588 ( .A1(n9744), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8298) );
  NAND2_X1 U10589 ( .A1(n9743), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8299) );
  NAND2_X1 U10590 ( .A1(n9747), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8302) );
  NAND2_X1 U10591 ( .A1(n9749), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8301) );
  NAND2_X1 U10592 ( .A1(n8302), .A2(n8301), .ZN(n8474) );
  NAND2_X1 U10593 ( .A1(n9753), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8304) );
  NAND2_X1 U10594 ( .A1(n9752), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8303) );
  NAND2_X1 U10595 ( .A1(n8491), .A2(n8304), .ZN(n8498) );
  NAND2_X1 U10596 ( .A1(n9757), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8306) );
  NAND2_X1 U10597 ( .A1(n9756), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8305) );
  NAND2_X1 U10598 ( .A1(n9764), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8308) );
  NAND2_X1 U10599 ( .A1(n9762), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8307) );
  NAND2_X1 U10600 ( .A1(n9891), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8309) );
  XNOR2_X1 U10601 ( .A(n8310), .B(P1_DATAO_REG_12__SCAN_IN), .ZN(n8553) );
  NAND2_X1 U10602 ( .A1(n8560), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8313) );
  NAND2_X1 U10603 ( .A1(n8311), .A2(n10109), .ZN(n8312) );
  NAND2_X1 U10604 ( .A1(n10431), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8315) );
  NAND2_X1 U10605 ( .A1(n10536), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8317) );
  NAND2_X1 U10606 ( .A1(n10535), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8316) );
  NAND2_X1 U10607 ( .A1(n8317), .A2(n8316), .ZN(n8597) );
  NAND2_X1 U10608 ( .A1(n10683), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8319) );
  NAND2_X1 U10609 ( .A1(n10682), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U10610 ( .A1(n10815), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U10611 ( .A1(n10814), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8320) );
  NAND2_X1 U10612 ( .A1(n8322), .A2(n8320), .ZN(n8628) );
  INV_X1 U10613 ( .A(n8628), .ZN(n8321) );
  NAND2_X1 U10614 ( .A1(n8629), .A2(n8321), .ZN(n8323) );
  NAND2_X1 U10615 ( .A1(n11107), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8325) );
  NAND2_X1 U10616 ( .A1(n11106), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8324) );
  INV_X1 U10617 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11163) );
  NAND2_X1 U10618 ( .A1(n11163), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8327) );
  INV_X1 U10619 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11162) );
  NAND2_X1 U10620 ( .A1(n11162), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8326) );
  NAND2_X1 U10621 ( .A1(n8328), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8330) );
  NAND2_X1 U10622 ( .A1(n8330), .A2(n8329), .ZN(n8674) );
  NAND2_X1 U10623 ( .A1(n8676), .A2(n8330), .ZN(n8686) );
  INV_X1 U10624 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11259) );
  NAND2_X1 U10625 ( .A1(n11259), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8332) );
  INV_X1 U10626 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11258) );
  NAND2_X1 U10627 ( .A1(n11258), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8331) );
  AND2_X1 U10628 ( .A1(n8332), .A2(n8331), .ZN(n8685) );
  INV_X1 U10629 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11458) );
  XNOR2_X1 U10630 ( .A(n11458), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8697) );
  NAND2_X1 U10631 ( .A1(n11458), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8333) );
  XNOR2_X1 U10632 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8707) );
  INV_X1 U10633 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8334) );
  NAND2_X1 U10634 ( .A1(n8334), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8335) );
  NAND2_X1 U10635 ( .A1(n8336), .A2(n11777), .ZN(n8337) );
  NAND2_X1 U10636 ( .A1(n11863), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8339) );
  NAND2_X1 U10637 ( .A1(n11859), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8340) );
  AND2_X1 U10638 ( .A1(n14186), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8341) );
  INV_X1 U10639 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13591) );
  AND2_X1 U10640 ( .A1(n13591), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8342) );
  INV_X1 U10641 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14184) );
  NAND2_X1 U10642 ( .A1(n14184), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8343) );
  INV_X1 U10643 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8882) );
  XNOR2_X1 U10644 ( .A(n8882), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n8344) );
  XNOR2_X1 U10645 ( .A(n8879), .B(n8344), .ZN(n13065) );
  NAND4_X1 U10646 ( .A1(n8347), .A2(n8346), .A3(n8561), .A4(n8539), .ZN(n8350)
         );
  NAND4_X1 U10647 ( .A1(n8521), .A2(n8581), .A3(n8563), .A4(n8348), .ZN(n8349)
         );
  NOR2_X1 U10648 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n8354) );
  NOR2_X1 U10649 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), 
        .ZN(n8353) );
  INV_X1 U10650 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8356) );
  INV_X1 U10651 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8359) );
  INV_X1 U10652 ( .A(n8383), .ZN(n8385) );
  NAND2_X2 U10653 ( .A1(n10254), .A2(n7530), .ZN(n8463) );
  NAND2_X1 U10654 ( .A1(n13065), .A2(n12181), .ZN(n8364) );
  NAND2_X1 U10655 ( .A1(n12182), .A2(SI_28_), .ZN(n8363) );
  INV_X1 U10656 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n8366) );
  INV_X1 U10657 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n8365) );
  NAND2_X1 U10658 ( .A1(n8366), .A2(n8365), .ZN(n8443) );
  INV_X1 U10659 ( .A(n8443), .ZN(n8368) );
  NAND2_X1 U10660 ( .A1(n8368), .A2(n8367), .ZN(n8455) );
  NAND2_X1 U10661 ( .A1(n8369), .A2(n15149), .ZN(n8482) );
  INV_X1 U10662 ( .A(n8569), .ZN(n8372) );
  NAND2_X1 U10663 ( .A1(n8372), .A2(n15107), .ZN(n8587) );
  INV_X1 U10664 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8373) );
  INV_X1 U10665 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8375) );
  NOR2_X1 U10666 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(P3_REG3_REG_22__SCAN_IN), 
        .ZN(n8377) );
  INV_X1 U10667 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8379) );
  INV_X1 U10668 ( .A(n8752), .ZN(n8381) );
  NAND2_X1 U10669 ( .A1(n8381), .A2(n15109), .ZN(n12373) );
  NAND2_X1 U10670 ( .A1(n8752), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U10671 ( .A1(n12373), .A2(n8382), .ZN(n12640) );
  NAND2_X1 U10672 ( .A1(n8383), .A2(n8386), .ZN(n13057) );
  INV_X1 U10673 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13005) );
  NAND2_X1 U10674 ( .A1(n12172), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8391) );
  NAND2_X1 U10675 ( .A1(n8887), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8390) );
  OAI211_X1 U10676 ( .C1(n13005), .C2(n8890), .A(n8391), .B(n8390), .ZN(n8392)
         );
  NAND2_X1 U10677 ( .A1(n12391), .A2(n12652), .ZN(n8898) );
  NAND2_X1 U10678 ( .A1(n12173), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8395) );
  INV_X1 U10679 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10716) );
  OR2_X1 U10680 ( .A1(n6484), .A2(n10716), .ZN(n8394) );
  INV_X1 U10681 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10358) );
  OR2_X1 U10682 ( .A1(n8420), .A2(n10358), .ZN(n8393) );
  INV_X1 U10683 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10352) );
  NAND2_X1 U10684 ( .A1(n9120), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8396) );
  INV_X1 U10685 ( .A(n10254), .ZN(n8603) );
  NAND2_X1 U10686 ( .A1(n8603), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n8397) );
  NAND2_X1 U10687 ( .A1(n12173), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U10688 ( .A1(n12172), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8401) );
  INV_X1 U10689 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10877) );
  OR2_X1 U10690 ( .A1(n8776), .A2(n10877), .ZN(n8400) );
  INV_X1 U10691 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10880) );
  OR2_X1 U10692 ( .A1(n8420), .A2(n10880), .ZN(n8399) );
  XNOR2_X1 U10693 ( .A(n8404), .B(n8403), .ZN(n9695) );
  INV_X1 U10694 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8406) );
  NAND2_X1 U10695 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8405) );
  OAI22_X1 U10696 ( .A1(n8463), .A2(n9695), .B1(n10254), .B2(n10360), .ZN(
        n8408) );
  INV_X1 U10697 ( .A(SI_1_), .ZN(n9694) );
  NOR2_X1 U10698 ( .A1(n8663), .A2(n9694), .ZN(n8407) );
  NAND2_X1 U10699 ( .A1(n12521), .A2(n10804), .ZN(n12229) );
  NAND2_X1 U10700 ( .A1(n12222), .A2(n12229), .ZN(n10745) );
  NAND2_X1 U10701 ( .A1(n8887), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8413) );
  INV_X1 U10702 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n11063) );
  OR2_X1 U10703 ( .A1(n6485), .A2(n11063), .ZN(n8412) );
  INV_X1 U10704 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8409) );
  INV_X1 U10705 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10350) );
  OR2_X1 U10706 ( .A1(n8779), .A2(n10350), .ZN(n8410) );
  XNOR2_X1 U10707 ( .A(n8415), .B(n8414), .ZN(n9679) );
  XNOR2_X2 U10708 ( .A(n8417), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10378) );
  OAI22_X1 U10709 ( .A1(n8463), .A2(n9679), .B1(n6483), .B2(n10254), .ZN(n8419) );
  NOR2_X1 U10710 ( .A1(n8663), .A2(SI_2_), .ZN(n8418) );
  NAND2_X1 U10711 ( .A1(n10875), .A2(n11062), .ZN(n12232) );
  INV_X1 U10712 ( .A(n11062), .ZN(n10752) );
  NAND2_X1 U10713 ( .A1(n12520), .A2(n10752), .ZN(n12236) );
  NAND2_X1 U10714 ( .A1(n12232), .A2(n12236), .ZN(n8785) );
  NAND2_X1 U10715 ( .A1(n11055), .A2(n12224), .ZN(n11054) );
  NAND2_X1 U10716 ( .A1(n11054), .A2(n12232), .ZN(n10821) );
  NAND2_X1 U10717 ( .A1(n12173), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8424) );
  OR2_X1 U10718 ( .A1(n6484), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8423) );
  INV_X1 U10719 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10829) );
  OR2_X1 U10720 ( .A1(n8420), .A2(n10829), .ZN(n8422) );
  INV_X1 U10721 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10381) );
  OR2_X1 U10722 ( .A1(n8779), .A2(n10381), .ZN(n8421) );
  NAND4_X1 U10723 ( .A1(n8424), .A2(n8423), .A3(n8422), .A4(n8421), .ZN(n12519) );
  XNOR2_X1 U10724 ( .A(n8426), .B(n8425), .ZN(n9709) );
  NAND2_X1 U10725 ( .A1(n12181), .A2(n9709), .ZN(n8430) );
  NAND2_X1 U10726 ( .A1(n8427), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8428) );
  XNOR2_X1 U10727 ( .A(n8428), .B(n8345), .ZN(n10442) );
  NAND2_X1 U10728 ( .A1(n8603), .A2(n10442), .ZN(n8429) );
  OAI211_X1 U10729 ( .C1(SI_3_), .C2(n8663), .A(n8430), .B(n8429), .ZN(n10969)
         );
  OR2_X1 U10730 ( .A1(n12519), .A2(n10969), .ZN(n12241) );
  NAND2_X1 U10731 ( .A1(n12519), .A2(n10969), .ZN(n12238) );
  NAND2_X1 U10732 ( .A1(n12241), .A2(n12238), .ZN(n8786) );
  INV_X1 U10733 ( .A(n8786), .ZN(n12198) );
  NAND2_X1 U10734 ( .A1(n12172), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8436) );
  INV_X1 U10735 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11376) );
  OR2_X1 U10736 ( .A1(n8420), .A2(n11376), .ZN(n8435) );
  NAND2_X1 U10737 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8431) );
  AND2_X1 U10738 ( .A1(n8443), .A2(n8431), .ZN(n11218) );
  OR2_X1 U10739 ( .A1(n6484), .A2(n11218), .ZN(n8434) );
  INV_X1 U10740 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8432) );
  OR2_X1 U10741 ( .A1(n8890), .A2(n8432), .ZN(n8433) );
  XNOR2_X1 U10742 ( .A(n8438), .B(n8437), .ZN(n9681) );
  NAND2_X1 U10743 ( .A1(n8439), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8440) );
  XNOR2_X1 U10744 ( .A(n8440), .B(P3_IR_REG_4__SCAN_IN), .ZN(n11406) );
  OAI22_X1 U10745 ( .A1(n8463), .A2(n9681), .B1(n11406), .B2(n6653), .ZN(n8442) );
  NOR2_X1 U10746 ( .A1(n8663), .A2(SI_4_), .ZN(n8441) );
  NOR2_X1 U10747 ( .A1(n8442), .A2(n8441), .ZN(n11217) );
  NAND2_X1 U10748 ( .A1(n10825), .A2(n11217), .ZN(n12242) );
  INV_X1 U10749 ( .A(n11217), .ZN(n11037) );
  NAND2_X1 U10750 ( .A1(n12518), .A2(n11037), .ZN(n12243) );
  NAND2_X1 U10751 ( .A1(n12242), .A2(n12243), .ZN(n11220) );
  INV_X1 U10752 ( .A(n11220), .ZN(n12240) );
  NAND2_X1 U10753 ( .A1(n8887), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8449) );
  INV_X1 U10754 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15011) );
  NAND2_X1 U10755 ( .A1(n8443), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8444) );
  AND2_X1 U10756 ( .A1(n8455), .A2(n8444), .ZN(n11283) );
  OR2_X1 U10757 ( .A1(n6485), .A2(n11283), .ZN(n8447) );
  INV_X1 U10758 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n8445) );
  OR2_X1 U10759 ( .A1(n8890), .A2(n8445), .ZN(n8446) );
  XNOR2_X1 U10760 ( .A(n8451), .B(n8450), .ZN(n9701) );
  OR2_X1 U10761 ( .A1(n6580), .A2(n8357), .ZN(n8452) );
  XNOR2_X1 U10762 ( .A(n8452), .B(P3_IR_REG_5__SCAN_IN), .ZN(n11411) );
  OAI22_X1 U10763 ( .A1(n8463), .A2(n9701), .B1(n11411), .B2(n6653), .ZN(n8454) );
  NOR2_X1 U10764 ( .A1(n8663), .A2(SI_5_), .ZN(n8453) );
  NAND2_X1 U10765 ( .A1(n8936), .A2(n11282), .ZN(n12249) );
  INV_X1 U10766 ( .A(n11282), .ZN(n11157) );
  NAND2_X1 U10767 ( .A1(n12517), .A2(n11157), .ZN(n12248) );
  NAND2_X1 U10768 ( .A1(n12173), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8460) );
  INV_X1 U10769 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11413) );
  OR2_X1 U10770 ( .A1(n8779), .A2(n11413), .ZN(n8459) );
  INV_X1 U10771 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11414) );
  OR2_X1 U10772 ( .A1(n8420), .A2(n11414), .ZN(n8458) );
  NAND2_X1 U10773 ( .A1(n8455), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8456) );
  AND2_X1 U10774 ( .A1(n8468), .A2(n8456), .ZN(n11571) );
  OR2_X1 U10775 ( .A1(n6485), .A2(n11571), .ZN(n8457) );
  XNOR2_X1 U10776 ( .A(n9743), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8461) );
  XNOR2_X1 U10777 ( .A(n8462), .B(n8461), .ZN(n9716) );
  NAND2_X1 U10778 ( .A1(n12182), .A2(SI_6_), .ZN(n8467) );
  NAND2_X1 U10779 ( .A1(n8464), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8465) );
  XNOR2_X1 U10780 ( .A(n8465), .B(P3_IR_REG_6__SCAN_IN), .ZN(n11415) );
  NAND2_X1 U10781 ( .A1(n8603), .A2(n11415), .ZN(n8466) );
  NAND2_X1 U10782 ( .A1(n11516), .A2(n11358), .ZN(n12255) );
  INV_X1 U10783 ( .A(n11358), .ZN(n11572) );
  NAND2_X1 U10784 ( .A1(n12516), .A2(n11572), .ZN(n12256) );
  NAND2_X1 U10785 ( .A1(n11352), .A2(n12197), .ZN(n11351) );
  NAND2_X1 U10786 ( .A1(n11351), .A2(n12255), .ZN(n11512) );
  NAND2_X1 U10787 ( .A1(n12173), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8473) );
  INV_X1 U10788 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11420) );
  OR2_X1 U10789 ( .A1(n8779), .A2(n11420), .ZN(n8472) );
  INV_X1 U10790 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11421) );
  OR2_X1 U10791 ( .A1(n8420), .A2(n11421), .ZN(n8471) );
  NAND2_X1 U10792 ( .A1(n8468), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8469) );
  AND2_X1 U10793 ( .A1(n8482), .A2(n8469), .ZN(n11695) );
  OR2_X1 U10794 ( .A1(n6484), .A2(n11695), .ZN(n8470) );
  NAND2_X1 U10795 ( .A1(n8475), .A2(n8474), .ZN(n8476) );
  AND2_X1 U10796 ( .A1(n8477), .A2(n8476), .ZN(n9706) );
  NAND2_X1 U10797 ( .A1(n8492), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8479) );
  INV_X1 U10798 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8478) );
  XNOR2_X1 U10799 ( .A(n8479), .B(n8478), .ZN(n14901) );
  INV_X1 U10800 ( .A(n14901), .ZN(n11422) );
  OAI22_X1 U10801 ( .A1(n8463), .A2(n9706), .B1(n11422), .B2(n6653), .ZN(n8481) );
  NOR2_X1 U10802 ( .A1(n8663), .A2(SI_7_), .ZN(n8480) );
  NOR2_X1 U10803 ( .A1(n8481), .A2(n8480), .ZN(n8793) );
  NAND2_X1 U10804 ( .A1(n11101), .A2(n8793), .ZN(n12260) );
  INV_X1 U10805 ( .A(n8793), .ZN(n11696) );
  NAND2_X1 U10806 ( .A1(n12515), .A2(n11696), .ZN(n12261) );
  NAND2_X1 U10807 ( .A1(n12260), .A2(n12261), .ZN(n11515) );
  INV_X1 U10808 ( .A(n11515), .ZN(n12258) );
  NAND2_X1 U10809 ( .A1(n11512), .A2(n12258), .ZN(n11511) );
  NAND2_X1 U10810 ( .A1(n11511), .A2(n12260), .ZN(n11630) );
  NAND2_X1 U10811 ( .A1(n12173), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8487) );
  INV_X1 U10812 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11427) );
  OR2_X1 U10813 ( .A1(n8779), .A2(n11427), .ZN(n8486) );
  INV_X1 U10814 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11639) );
  OR2_X1 U10815 ( .A1(n8420), .A2(n11639), .ZN(n8485) );
  NAND2_X1 U10816 ( .A1(n8482), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8483) );
  AND2_X1 U10817 ( .A1(n8509), .A2(n8483), .ZN(n11638) );
  OR2_X1 U10818 ( .A1(n6485), .A2(n11638), .ZN(n8484) );
  OR2_X1 U10819 ( .A1(n8489), .A2(n8488), .ZN(n8490) );
  NAND2_X1 U10820 ( .A1(n8491), .A2(n8490), .ZN(n9700) );
  NAND2_X1 U10821 ( .A1(n12182), .A2(SI_8_), .ZN(n8495) );
  NAND2_X1 U10822 ( .A1(n8501), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8493) );
  XNOR2_X1 U10823 ( .A(n8493), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11428) );
  NAND2_X1 U10824 ( .A1(n8603), .A2(n11428), .ZN(n8494) );
  OAI211_X1 U10825 ( .C1(n8463), .C2(n9700), .A(n8495), .B(n8494), .ZN(n11637)
         );
  NAND2_X1 U10826 ( .A1(n11562), .A2(n11637), .ZN(n12265) );
  INV_X1 U10827 ( .A(n11562), .ZN(n12514) );
  INV_X1 U10828 ( .A(n11637), .ZN(n11173) );
  NAND2_X1 U10829 ( .A1(n12514), .A2(n11173), .ZN(n12266) );
  AND2_X2 U10830 ( .A1(n12265), .A2(n12266), .ZN(n12263) );
  NAND2_X1 U10831 ( .A1(n11630), .A2(n12263), .ZN(n8496) );
  OR2_X1 U10832 ( .A1(n8498), .A2(n8497), .ZN(n8499) );
  NAND2_X1 U10833 ( .A1(n8500), .A2(n8499), .ZN(n9704) );
  NAND2_X1 U10834 ( .A1(n12181), .A2(n9704), .ZN(n8508) );
  NOR2_X1 U10835 ( .A1(n8505), .A2(n8357), .ZN(n8502) );
  MUX2_X1 U10836 ( .A(n8357), .B(n8502), .S(P3_IR_REG_9__SCAN_IN), .Z(n8503)
         );
  INV_X1 U10837 ( .A(n8503), .ZN(n8506) );
  INV_X1 U10838 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8504) );
  NAND2_X1 U10839 ( .A1(n8505), .A2(n8504), .ZN(n8538) );
  NAND2_X1 U10840 ( .A1(n8506), .A2(n8538), .ZN(n14938) );
  NAND2_X1 U10841 ( .A1(n8603), .A2(n14938), .ZN(n8507) );
  INV_X1 U10842 ( .A(n12270), .ZN(n8792) );
  NAND2_X1 U10843 ( .A1(n12173), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8514) );
  INV_X1 U10844 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11434) );
  OR2_X1 U10845 ( .A1(n8420), .A2(n11434), .ZN(n8513) );
  NAND2_X1 U10846 ( .A1(n8509), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8510) );
  AND2_X1 U10847 ( .A1(n8515), .A2(n8510), .ZN(n11566) );
  OR2_X1 U10848 ( .A1(n6484), .A2(n11566), .ZN(n8512) );
  INV_X1 U10849 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11433) );
  OR2_X1 U10850 ( .A1(n8779), .A2(n11433), .ZN(n8511) );
  NAND4_X1 U10851 ( .A1(n8514), .A2(n8513), .A3(n8512), .A4(n8511), .ZN(n12513) );
  INV_X1 U10852 ( .A(n12513), .ZN(n11174) );
  NAND2_X1 U10853 ( .A1(n12173), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8520) );
  INV_X1 U10854 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11440) );
  OR2_X1 U10855 ( .A1(n8779), .A2(n11440), .ZN(n8519) );
  INV_X1 U10856 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11691) );
  OR2_X1 U10857 ( .A1(n8420), .A2(n11691), .ZN(n8518) );
  NAND2_X1 U10858 ( .A1(n8515), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8516) );
  AND2_X1 U10859 ( .A1(n8529), .A2(n8516), .ZN(n11690) );
  OR2_X1 U10860 ( .A1(n6485), .A2(n11690), .ZN(n8517) );
  INV_X1 U10861 ( .A(n12905), .ZN(n12512) );
  NAND2_X1 U10862 ( .A1(n8538), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8522) );
  XNOR2_X1 U10863 ( .A(n8522), .B(n8521), .ZN(n14969) );
  INV_X1 U10864 ( .A(n14969), .ZN(n11441) );
  OAI22_X1 U10865 ( .A1(n8663), .A2(SI_10_), .B1(n11441), .B2(n6653), .ZN(
        n8528) );
  OR2_X1 U10866 ( .A1(n8524), .A2(n8523), .ZN(n8525) );
  AND2_X1 U10867 ( .A1(n8526), .A2(n8525), .ZN(n9696) );
  NOR2_X1 U10868 ( .A1(n8463), .A2(n9696), .ZN(n8527) );
  INV_X1 U10869 ( .A(n12275), .ZN(n11347) );
  NAND2_X1 U10870 ( .A1(n12512), .A2(n11347), .ZN(n12892) );
  NAND2_X1 U10871 ( .A1(n12173), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8535) );
  NAND2_X1 U10872 ( .A1(n8529), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8530) );
  AND2_X1 U10873 ( .A1(n8544), .A2(n8530), .ZN(n12911) );
  OR2_X1 U10874 ( .A1(n6484), .A2(n12911), .ZN(n8534) );
  INV_X1 U10875 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12912) );
  OR2_X1 U10876 ( .A1(n8420), .A2(n12912), .ZN(n8533) );
  INV_X1 U10877 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n8531) );
  OR2_X1 U10878 ( .A1(n8779), .A2(n8531), .ZN(n8532) );
  XNOR2_X1 U10879 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8536) );
  XNOR2_X1 U10880 ( .A(n8537), .B(n8536), .ZN(n9713) );
  NAND2_X1 U10881 ( .A1(n12181), .A2(n9713), .ZN(n8542) );
  NAND2_X1 U10882 ( .A1(n8550), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8540) );
  XNOR2_X1 U10883 ( .A(n8540), .B(n8539), .ZN(n11490) );
  NAND2_X1 U10884 ( .A1(n8603), .A2(n11490), .ZN(n8541) );
  OAI211_X1 U10885 ( .C1(SI_11_), .C2(n8663), .A(n8542), .B(n8541), .ZN(n12909) );
  INV_X1 U10886 ( .A(n12909), .ZN(n8804) );
  NAND2_X1 U10887 ( .A1(n12876), .A2(n8804), .ZN(n12279) );
  NAND2_X1 U10888 ( .A1(n12511), .A2(n12909), .ZN(n12284) );
  AND2_X1 U10889 ( .A1(n12892), .A2(n12899), .ZN(n12884) );
  NAND2_X1 U10890 ( .A1(n12173), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8549) );
  INV_X1 U10891 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12882) );
  OR2_X1 U10892 ( .A1(n8420), .A2(n12882), .ZN(n8548) );
  INV_X1 U10893 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n8543) );
  OR2_X1 U10894 ( .A1(n8779), .A2(n8543), .ZN(n8547) );
  NAND2_X1 U10895 ( .A1(n8544), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8545) );
  AND2_X1 U10896 ( .A1(n8569), .A2(n8545), .ZN(n12881) );
  OR2_X1 U10897 ( .A1(n6484), .A2(n12881), .ZN(n8546) );
  OR2_X1 U10898 ( .A1(n8562), .A2(n8357), .ZN(n8551) );
  XNOR2_X1 U10899 ( .A(n8551), .B(P3_IR_REG_12__SCAN_IN), .ZN(n11539) );
  OAI22_X1 U10900 ( .A1(n8663), .A2(n9724), .B1(n6653), .B2(n11545), .ZN(n8552) );
  INV_X1 U10901 ( .A(n8552), .ZN(n8556) );
  XNOR2_X1 U10902 ( .A(n8554), .B(n8553), .ZN(n9722) );
  NAND2_X1 U10903 ( .A1(n12181), .A2(n9722), .ZN(n8555) );
  NAND2_X1 U10904 ( .A1(n8556), .A2(n8555), .ZN(n12880) );
  NAND2_X1 U10905 ( .A1(n12907), .A2(n12880), .ZN(n12863) );
  INV_X1 U10906 ( .A(n12907), .ZN(n12510) );
  INV_X1 U10907 ( .A(n12880), .ZN(n11622) );
  NAND2_X1 U10908 ( .A1(n12510), .A2(n11622), .ZN(n12286) );
  NAND2_X1 U10909 ( .A1(n12863), .A2(n12286), .ZN(n12207) );
  AND2_X1 U10910 ( .A1(n12884), .A2(n12886), .ZN(n8559) );
  NAND2_X1 U10911 ( .A1(n12905), .A2(n12275), .ZN(n12894) );
  OR2_X1 U10912 ( .A1(n12901), .A2(n12894), .ZN(n12896) );
  AND2_X1 U10913 ( .A1(n12896), .A2(n12279), .ZN(n12885) );
  OR2_X1 U10914 ( .A1(n12207), .A2(n12885), .ZN(n8557) );
  INV_X1 U10915 ( .A(n8557), .ZN(n8558) );
  XNOR2_X1 U10916 ( .A(n8560), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9750) );
  NAND2_X1 U10917 ( .A1(n9750), .A2(n12181), .ZN(n8567) );
  NAND2_X1 U10918 ( .A1(n8562), .A2(n8561), .ZN(n8580) );
  NAND2_X1 U10919 ( .A1(n8580), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8564) );
  XNOR2_X1 U10920 ( .A(n8564), .B(n8563), .ZN(n12529) );
  OAI22_X1 U10921 ( .A1(n8663), .A2(SI_13_), .B1(n12538), .B2(n6653), .ZN(
        n8565) );
  INV_X1 U10922 ( .A(n8565), .ZN(n8566) );
  INV_X1 U10923 ( .A(n13052), .ZN(n8575) );
  NAND2_X1 U10924 ( .A1(n12173), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8574) );
  INV_X1 U10925 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12994) );
  OR2_X1 U10926 ( .A1(n8779), .A2(n12994), .ZN(n8573) );
  INV_X1 U10927 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n8568) );
  OR2_X1 U10928 ( .A1(n8420), .A2(n8568), .ZN(n8572) );
  NAND2_X1 U10929 ( .A1(n8569), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8570) );
  AND2_X1 U10930 ( .A1(n8587), .A2(n8570), .ZN(n11725) );
  OR2_X1 U10931 ( .A1(n6485), .A2(n11725), .ZN(n8571) );
  AND2_X1 U10932 ( .A1(n8575), .A2(n12875), .ZN(n12288) );
  INV_X1 U10933 ( .A(n12288), .ZN(n8576) );
  AND2_X1 U10934 ( .A1(n8576), .A2(n12863), .ZN(n8577) );
  XNOR2_X1 U10935 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8578) );
  XNOR2_X1 U10936 ( .A(n8579), .B(n8578), .ZN(n9755) );
  NAND2_X1 U10937 ( .A1(n9755), .A2(n12181), .ZN(n8586) );
  NAND2_X1 U10938 ( .A1(n8601), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8582) );
  XNOR2_X1 U10939 ( .A(n8582), .B(n8581), .ZN(n12558) );
  INV_X1 U10940 ( .A(n12558), .ZN(n8583) );
  OAI22_X1 U10941 ( .A1(n8663), .A2(SI_14_), .B1(n8583), .B2(n6653), .ZN(n8584) );
  INV_X1 U10942 ( .A(n8584), .ZN(n8585) );
  NAND2_X1 U10943 ( .A1(n12172), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8593) );
  INV_X1 U10944 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12856) );
  OR2_X1 U10945 ( .A1(n8420), .A2(n12856), .ZN(n8592) );
  NAND2_X1 U10946 ( .A1(n8587), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8588) );
  AND2_X1 U10947 ( .A1(n8606), .A2(n8588), .ZN(n12855) );
  OR2_X1 U10948 ( .A1(n6485), .A2(n12855), .ZN(n8591) );
  INV_X1 U10949 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n8589) );
  OR2_X1 U10950 ( .A1(n8890), .A2(n8589), .ZN(n8590) );
  XNOR2_X1 U10951 ( .A(n13046), .B(n12862), .ZN(n12852) );
  NAND2_X1 U10952 ( .A1(n13052), .A2(n8969), .ZN(n12850) );
  AND2_X1 U10953 ( .A1(n12852), .A2(n12850), .ZN(n8594) );
  NAND2_X1 U10954 ( .A1(n12851), .A2(n8594), .ZN(n8596) );
  OR2_X1 U10955 ( .A1(n13046), .A2(n12509), .ZN(n8595) );
  NAND2_X1 U10956 ( .A1(n8598), .A2(n8597), .ZN(n8599) );
  NAND2_X1 U10957 ( .A1(n8600), .A2(n8599), .ZN(n9796) );
  OR2_X1 U10958 ( .A1(n9796), .A2(n8463), .ZN(n8605) );
  OAI21_X1 U10959 ( .B1(n8601), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8602) );
  XNOR2_X1 U10960 ( .A(n8602), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12588) );
  AOI22_X1 U10961 ( .A1(n12182), .A2(SI_15_), .B1(n8603), .B2(n12588), .ZN(
        n8604) );
  NAND2_X1 U10962 ( .A1(n8605), .A2(n8604), .ZN(n12835) );
  NAND2_X1 U10963 ( .A1(n12173), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8611) );
  INV_X1 U10964 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12553) );
  OR2_X1 U10965 ( .A1(n8420), .A2(n12553), .ZN(n8610) );
  INV_X1 U10966 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12985) );
  OR2_X1 U10967 ( .A1(n8779), .A2(n12985), .ZN(n8609) );
  NAND2_X1 U10968 ( .A1(n8606), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8607) );
  AND2_X1 U10969 ( .A1(n8622), .A2(n8607), .ZN(n12836) );
  OR2_X1 U10970 ( .A1(n6485), .A2(n12836), .ZN(n8608) );
  NAND4_X1 U10971 ( .A1(n8611), .A2(n8610), .A3(n8609), .A4(n8608), .ZN(n12845) );
  INV_X1 U10972 ( .A(n12845), .ZN(n12398) );
  OR2_X1 U10973 ( .A1(n12835), .A2(n12398), .ZN(n12291) );
  NAND2_X1 U10974 ( .A1(n12835), .A2(n12398), .ZN(n12299) );
  NAND2_X1 U10975 ( .A1(n12834), .A2(n12833), .ZN(n8612) );
  NAND2_X1 U10976 ( .A1(n8612), .A2(n12299), .ZN(n12822) );
  OR2_X1 U10977 ( .A1(n8614), .A2(n8613), .ZN(n8615) );
  NAND2_X1 U10978 ( .A1(n8616), .A2(n8615), .ZN(n10010) );
  NAND2_X1 U10979 ( .A1(n8617), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8618) );
  XNOR2_X1 U10980 ( .A(n8618), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12617) );
  OAI22_X1 U10981 ( .A1(n8663), .A2(n15094), .B1(n6653), .B2(n12598), .ZN(
        n8619) );
  INV_X1 U10982 ( .A(n8619), .ZN(n8620) );
  NAND2_X1 U10983 ( .A1(n12173), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8627) );
  INV_X1 U10984 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12616) );
  OR2_X1 U10985 ( .A1(n8779), .A2(n12616), .ZN(n8626) );
  INV_X1 U10986 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12825) );
  OR2_X1 U10987 ( .A1(n8420), .A2(n12825), .ZN(n8625) );
  NAND2_X1 U10988 ( .A1(n8622), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8623) );
  AND2_X1 U10989 ( .A1(n8638), .A2(n8623), .ZN(n12824) );
  OR2_X1 U10990 ( .A1(n6485), .A2(n12824), .ZN(n8624) );
  OR2_X1 U10991 ( .A1(n12978), .A2(n12832), .ZN(n12290) );
  NAND2_X1 U10992 ( .A1(n12978), .A2(n12832), .ZN(n12300) );
  NAND2_X1 U10993 ( .A1(n12290), .A2(n12300), .ZN(n8813) );
  NAND2_X1 U10994 ( .A1(n12822), .A2(n12821), .ZN(n12820) );
  XNOR2_X1 U10995 ( .A(n8629), .B(n8628), .ZN(n10087) );
  NAND2_X1 U10996 ( .A1(n10087), .A2(n12181), .ZN(n8637) );
  NOR2_X1 U10997 ( .A1(n8630), .A2(n8357), .ZN(n8631) );
  MUX2_X1 U10998 ( .A(n8357), .B(n8631), .S(P3_IR_REG_17__SCAN_IN), .Z(n8632)
         );
  INV_X1 U10999 ( .A(n8632), .ZN(n8634) );
  AND2_X1 U11000 ( .A1(n8634), .A2(n8633), .ZN(n14330) );
  OAI22_X1 U11001 ( .A1(n8663), .A2(n10088), .B1(n6653), .B2(n12618), .ZN(
        n8635) );
  INV_X1 U11002 ( .A(n8635), .ZN(n8636) );
  NAND2_X1 U11003 ( .A1(n12173), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8644) );
  INV_X1 U11004 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12812) );
  OR2_X1 U11005 ( .A1(n8420), .A2(n12812), .ZN(n8643) );
  NAND2_X1 U11006 ( .A1(n8638), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8639) );
  AND2_X1 U11007 ( .A1(n8653), .A2(n8639), .ZN(n12811) );
  OR2_X1 U11008 ( .A1(n6484), .A2(n12811), .ZN(n8642) );
  INV_X1 U11009 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n8640) );
  OR2_X1 U11010 ( .A1(n8779), .A2(n8640), .ZN(n8641) );
  OR2_X1 U11011 ( .A1(n12974), .A2(n12791), .ZN(n12308) );
  NAND2_X1 U11012 ( .A1(n12974), .A2(n12791), .ZN(n12794) );
  NAND2_X1 U11013 ( .A1(n12308), .A2(n12794), .ZN(n12211) );
  OR2_X1 U11014 ( .A1(n8646), .A2(n8645), .ZN(n8647) );
  NAND2_X1 U11015 ( .A1(n8648), .A2(n8647), .ZN(n10112) );
  OR2_X1 U11016 ( .A1(n10112), .A2(n8463), .ZN(n8652) );
  NAND2_X1 U11017 ( .A1(n8633), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8649) );
  XNOR2_X1 U11018 ( .A(n8649), .B(P3_IR_REG_18__SCAN_IN), .ZN(n14342) );
  OAI22_X1 U11019 ( .A1(n8663), .A2(n15126), .B1(n6653), .B2(n12614), .ZN(
        n8650) );
  INV_X1 U11020 ( .A(n8650), .ZN(n8651) );
  NAND2_X1 U11021 ( .A1(n8887), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8658) );
  INV_X1 U11022 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12972) );
  OR2_X1 U11023 ( .A1(n8779), .A2(n12972), .ZN(n8657) );
  NAND2_X1 U11024 ( .A1(n8653), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8654) );
  AND2_X1 U11025 ( .A1(n8667), .A2(n8654), .ZN(n12793) );
  OR2_X1 U11026 ( .A1(n6484), .A2(n12793), .ZN(n8656) );
  INV_X1 U11027 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13036) );
  OR2_X1 U11028 ( .A1(n8890), .A2(n13036), .ZN(n8655) );
  NAND2_X1 U11029 ( .A1(n12967), .A2(n12775), .ZN(n12313) );
  AND2_X1 U11030 ( .A1(n12789), .A2(n12794), .ZN(n8659) );
  XNOR2_X1 U11031 ( .A(n8661), .B(n8660), .ZN(n10155) );
  NAND2_X1 U11032 ( .A1(n10155), .A2(n12181), .ZN(n8666) );
  NAND2_X1 U11033 ( .A1(n8761), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8662) );
  OAI22_X1 U11034 ( .A1(n8663), .A2(SI_19_), .B1(n12609), .B2(n6653), .ZN(
        n8664) );
  INV_X1 U11035 ( .A(n8664), .ZN(n8665) );
  NAND2_X1 U11036 ( .A1(n12173), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8672) );
  INV_X1 U11037 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12782) );
  OR2_X1 U11038 ( .A1(n8420), .A2(n12782), .ZN(n8671) );
  NAND2_X1 U11039 ( .A1(n8667), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8668) );
  OR2_X1 U11040 ( .A1(n6485), .A2(n12781), .ZN(n8670) );
  INV_X1 U11041 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12964) );
  OR2_X1 U11042 ( .A1(n8779), .A2(n12964), .ZN(n8669) );
  NAND4_X1 U11043 ( .A1(n8672), .A2(n8671), .A3(n8670), .A4(n8669), .ZN(n12508) );
  NAND2_X1 U11044 ( .A1(n13034), .A2(n12508), .ZN(n12317) );
  INV_X1 U11045 ( .A(n12317), .ZN(n8673) );
  OR2_X1 U11046 ( .A1(n13034), .A2(n12508), .ZN(n12316) );
  NAND2_X1 U11047 ( .A1(n8674), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U11048 ( .A1(n8676), .A2(n8675), .ZN(n10456) );
  NAND2_X1 U11049 ( .A1(n12182), .A2(SI_20_), .ZN(n8677) );
  NAND2_X1 U11050 ( .A1(n8679), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8680) );
  NAND2_X1 U11051 ( .A1(n8701), .A2(n8680), .ZN(n12760) );
  NAND2_X1 U11052 ( .A1(n8754), .A2(n12760), .ZN(n8684) );
  INV_X1 U11053 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12762) );
  OR2_X1 U11054 ( .A1(n8420), .A2(n12762), .ZN(n8683) );
  INV_X1 U11055 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13028) );
  OR2_X1 U11056 ( .A1(n8890), .A2(n13028), .ZN(n8682) );
  INV_X1 U11057 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12959) );
  OR2_X1 U11058 ( .A1(n8779), .A2(n12959), .ZN(n8681) );
  XNOR2_X1 U11059 ( .A(n12954), .B(n12774), .ZN(n12763) );
  OR2_X1 U11060 ( .A1(n12954), .A2(n12774), .ZN(n12320) );
  OR2_X1 U11061 ( .A1(n8686), .A2(n8685), .ZN(n8687) );
  NAND2_X1 U11062 ( .A1(n8688), .A2(n8687), .ZN(n10539) );
  NAND2_X1 U11063 ( .A1(n12182), .A2(SI_21_), .ZN(n8689) );
  NAND2_X1 U11064 ( .A1(n12172), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8692) );
  NAND2_X1 U11065 ( .A1(n8887), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8691) );
  AND2_X1 U11066 ( .A1(n8692), .A2(n8691), .ZN(n8695) );
  XNOR2_X1 U11067 ( .A(n8701), .B(P3_REG3_REG_21__SCAN_IN), .ZN(n12749) );
  NAND2_X1 U11068 ( .A1(n12749), .A2(n8754), .ZN(n8694) );
  NAND2_X1 U11069 ( .A1(n12173), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8693) );
  NAND2_X1 U11070 ( .A1(n12748), .A2(n12759), .ZN(n12323) );
  NAND2_X1 U11071 ( .A1(n12747), .A2(n12323), .ZN(n8696) );
  XNOR2_X1 U11072 ( .A(n8698), .B(n8697), .ZN(n10721) );
  NAND2_X1 U11073 ( .A1(n10721), .A2(n12181), .ZN(n8700) );
  NAND2_X1 U11074 ( .A1(n12182), .A2(SI_22_), .ZN(n8699) );
  INV_X1 U11075 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13020) );
  OAI21_X1 U11076 ( .B1(n8701), .B2(P3_REG3_REG_21__SCAN_IN), .A(
        P3_REG3_REG_22__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U11077 ( .A1(n8702), .A2(n8711), .ZN(n12731) );
  NAND2_X1 U11078 ( .A1(n12731), .A2(n8754), .ZN(n8706) );
  NAND2_X1 U11079 ( .A1(n12172), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U11080 ( .A1(n8887), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8703) );
  AND2_X1 U11081 ( .A1(n8704), .A2(n8703), .ZN(n8705) );
  INV_X1 U11082 ( .A(n12708), .ZN(n12745) );
  NAND2_X1 U11083 ( .A1(n12730), .A2(n12745), .ZN(n12713) );
  XNOR2_X1 U11084 ( .A(n8708), .B(n8707), .ZN(n10833) );
  NAND2_X1 U11085 ( .A1(n10833), .A2(n12181), .ZN(n8710) );
  NAND2_X1 U11086 ( .A1(n12182), .A2(SI_23_), .ZN(n8709) );
  NAND2_X1 U11087 ( .A1(n8711), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8712) );
  NAND2_X1 U11088 ( .A1(n8721), .A2(n8712), .ZN(n12720) );
  NAND2_X1 U11089 ( .A1(n12720), .A2(n8754), .ZN(n8715) );
  AOI22_X1 U11090 ( .A1(n8887), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n12172), 
        .B2(P3_REG1_REG_23__SCAN_IN), .ZN(n8714) );
  NAND2_X1 U11091 ( .A1(n12173), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U11092 ( .A1(n12721), .A2(n12728), .ZN(n8716) );
  NAND2_X1 U11093 ( .A1(n12696), .A2(n8716), .ZN(n12706) );
  AND2_X1 U11094 ( .A1(n12713), .A2(n12716), .ZN(n8717) );
  NAND2_X1 U11095 ( .A1(n12712), .A2(n8717), .ZN(n12695) );
  NAND2_X1 U11096 ( .A1(n8718), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8719) );
  INV_X1 U11097 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n8725) );
  NAND2_X1 U11098 ( .A1(n8721), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U11099 ( .A1(n8731), .A2(n8722), .ZN(n12700) );
  NAND2_X1 U11100 ( .A1(n12700), .A2(n8754), .ZN(n8724) );
  AOI22_X1 U11101 ( .A1(n8887), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n12172), 
        .B2(P3_REG1_REG_24__SCAN_IN), .ZN(n8723) );
  OAI211_X1 U11102 ( .C1(n8890), .C2(n8725), .A(n8724), .B(n8723), .ZN(n12709)
         );
  OR2_X1 U11103 ( .A1(n12730), .A2(n12745), .ZN(n12714) );
  OR2_X1 U11104 ( .A1(n12706), .A2(n12714), .ZN(n12694) );
  AND2_X1 U11105 ( .A1(n12332), .A2(n12694), .ZN(n8726) );
  INV_X1 U11106 ( .A(n12702), .ZN(n12937) );
  INV_X1 U11107 ( .A(n12709), .ZN(n12408) );
  NAND2_X1 U11108 ( .A1(n12937), .A2(n12408), .ZN(n12330) );
  XNOR2_X1 U11109 ( .A(n11863), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8727) );
  XNOR2_X1 U11110 ( .A(n8728), .B(n8727), .ZN(n11475) );
  NAND2_X1 U11111 ( .A1(n11475), .A2(n12181), .ZN(n8730) );
  NAND2_X1 U11112 ( .A1(n12182), .A2(SI_25_), .ZN(n8729) );
  NAND2_X1 U11113 ( .A1(n8731), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U11114 ( .A1(n8751), .A2(n8732), .ZN(n12683) );
  INV_X1 U11115 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n8735) );
  NAND2_X1 U11116 ( .A1(n12172), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8734) );
  NAND2_X1 U11117 ( .A1(n8887), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8733) );
  OAI211_X1 U11118 ( .C1(n8735), .C2(n8890), .A(n8734), .B(n8733), .ZN(n8736)
         );
  OR2_X1 U11119 ( .A1(n12933), .A2(n12690), .ZN(n12336) );
  NAND2_X1 U11120 ( .A1(n12933), .A2(n12690), .ZN(n8737) );
  NAND2_X1 U11121 ( .A1(n12336), .A2(n8737), .ZN(n12677) );
  INV_X1 U11122 ( .A(n8737), .ZN(n12333) );
  XNOR2_X1 U11123 ( .A(n13594), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n8738) );
  XNOR2_X1 U11124 ( .A(n8739), .B(n8738), .ZN(n11533) );
  NAND2_X1 U11125 ( .A1(n11533), .A2(n12181), .ZN(n8741) );
  NAND2_X1 U11126 ( .A1(n12182), .A2(SI_26_), .ZN(n8740) );
  XNOR2_X1 U11127 ( .A(n8751), .B(P3_REG3_REG_26__SCAN_IN), .ZN(n12671) );
  NAND2_X1 U11128 ( .A1(n12671), .A2(n8754), .ZN(n8746) );
  INV_X1 U11129 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13013) );
  NAND2_X1 U11130 ( .A1(n8887), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U11131 ( .A1(n12172), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8742) );
  OAI211_X1 U11132 ( .C1(n13013), .C2(n8890), .A(n8743), .B(n8742), .ZN(n8744)
         );
  INV_X1 U11133 ( .A(n8744), .ZN(n8745) );
  NOR2_X1 U11134 ( .A1(n9001), .A2(n12651), .ZN(n12334) );
  XNOR2_X1 U11135 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8747) );
  XNOR2_X1 U11136 ( .A(n8748), .B(n8747), .ZN(n11616) );
  NAND2_X1 U11137 ( .A1(n11616), .A2(n12181), .ZN(n8750) );
  NAND2_X1 U11138 ( .A1(n12182), .A2(SI_27_), .ZN(n8749) );
  OAI21_X1 U11139 ( .B1(n8751), .B2(P3_REG3_REG_26__SCAN_IN), .A(
        P3_REG3_REG_27__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U11140 ( .A1(n8753), .A2(n8752), .ZN(n12657) );
  NAND2_X1 U11141 ( .A1(n12657), .A2(n8754), .ZN(n8759) );
  INV_X1 U11142 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13009) );
  NAND2_X1 U11143 ( .A1(n8887), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U11144 ( .A1(n12172), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8755) );
  OAI211_X1 U11145 ( .C1(n8890), .C2(n13009), .A(n8756), .B(n8755), .ZN(n8757)
         );
  INV_X1 U11146 ( .A(n8757), .ZN(n8758) );
  NAND2_X1 U11147 ( .A1(n12339), .A2(n12665), .ZN(n8897) );
  NAND2_X1 U11148 ( .A1(n12648), .A2(n8897), .ZN(n8760) );
  XOR2_X1 U11149 ( .A(n12380), .B(n8760), .Z(n12643) );
  NAND2_X1 U11150 ( .A1(n8833), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8764) );
  INV_X1 U11151 ( .A(n8765), .ZN(n8766) );
  NAND2_X1 U11152 ( .A1(n8766), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8767) );
  OAI21_X1 U11153 ( .B1(n12218), .B2(n8904), .A(n12609), .ZN(n8772) );
  INV_X1 U11154 ( .A(n8768), .ZN(n8769) );
  NAND2_X1 U11155 ( .A1(n8769), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8771) );
  XNOR2_X2 U11156 ( .A(n8771), .B(n8770), .ZN(n10538) );
  NAND2_X1 U11157 ( .A1(n8772), .A2(n10538), .ZN(n8774) );
  OAI21_X1 U11158 ( .B1(n8904), .B2(n12221), .A(n12218), .ZN(n8773) );
  NAND2_X1 U11159 ( .A1(n8774), .A2(n8773), .ZN(n9019) );
  NAND2_X1 U11160 ( .A1(n9019), .A2(n12941), .ZN(n10618) );
  NAND2_X1 U11161 ( .A1(n10455), .A2(n12193), .ZN(n8867) );
  OR2_X1 U11162 ( .A1(n10618), .A2(n8867), .ZN(n8775) );
  OR3_X1 U11163 ( .A1(n12218), .A2(n12609), .A3(n10455), .ZN(n8868) );
  AND2_X1 U11164 ( .A1(n8775), .A2(n8868), .ZN(n10818) );
  NAND2_X1 U11165 ( .A1(n12218), .A2(n11064), .ZN(n12924) );
  OR2_X1 U11166 ( .A1(n12373), .A2(n6484), .ZN(n12178) );
  INV_X1 U11167 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8780) );
  NAND2_X1 U11168 ( .A1(n8887), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8778) );
  NAND2_X1 U11169 ( .A1(n12173), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8777) );
  OAI211_X1 U11170 ( .C1(n8780), .C2(n8779), .A(n8778), .B(n8777), .ZN(n8781)
         );
  INV_X1 U11171 ( .A(n8781), .ZN(n8782) );
  INV_X1 U11172 ( .A(n13068), .ZN(n12364) );
  INV_X1 U11173 ( .A(n12610), .ZN(n12541) );
  NAND2_X1 U11174 ( .A1(n12364), .A2(n12541), .ZN(n10257) );
  NAND2_X1 U11175 ( .A1(n10257), .A2(n6653), .ZN(n8829) );
  INV_X1 U11176 ( .A(n12933), .ZN(n8826) );
  INV_X1 U11177 ( .A(n12721), .ZN(n12942) );
  NAND2_X1 U11178 ( .A1(n12523), .A2(n10811), .ZN(n8929) );
  NAND2_X1 U11179 ( .A1(n12202), .A2(n8929), .ZN(n8783) );
  INV_X1 U11180 ( .A(n12521), .ZN(n11058) );
  NAND2_X1 U11181 ( .A1(n11058), .A2(n10804), .ZN(n10743) );
  NAND2_X1 U11182 ( .A1(n8783), .A2(n10743), .ZN(n11056) );
  NOR2_X1 U11183 ( .A1(n12520), .A2(n11062), .ZN(n8784) );
  NAND2_X1 U11184 ( .A1(n10823), .A2(n8786), .ZN(n10827) );
  INV_X1 U11185 ( .A(n10969), .ZN(n10830) );
  NAND2_X1 U11186 ( .A1(n12519), .A2(n10830), .ZN(n8787) );
  NAND2_X1 U11187 ( .A1(n10827), .A2(n8787), .ZN(n11221) );
  NAND2_X1 U11188 ( .A1(n11221), .A2(n11220), .ZN(n11219) );
  NAND2_X1 U11189 ( .A1(n12518), .A2(n11217), .ZN(n8788) );
  NAND2_X1 U11190 ( .A1(n11219), .A2(n8788), .ZN(n11277) );
  OR2_X2 U11191 ( .A1(n11277), .A2(n12245), .ZN(n11278) );
  NAND2_X1 U11192 ( .A1(n8936), .A2(n11157), .ZN(n8789) );
  NAND2_X1 U11193 ( .A1(n12516), .A2(n11358), .ZN(n11513) );
  NAND2_X1 U11194 ( .A1(n12513), .A2(n8792), .ZN(n8797) );
  XNOR2_X1 U11195 ( .A(n12513), .B(n12270), .ZN(n12200) );
  NAND2_X1 U11196 ( .A1(n11562), .A2(n11173), .ZN(n8799) );
  INV_X1 U11197 ( .A(n8799), .ZN(n8796) );
  NAND2_X1 U11198 ( .A1(n12515), .A2(n8793), .ZN(n11631) );
  INV_X1 U11199 ( .A(n11631), .ZN(n8794) );
  OR2_X1 U11200 ( .A1(n8796), .A2(n8795), .ZN(n11554) );
  OR2_X1 U11201 ( .A1(n12268), .A2(n11554), .ZN(n11558) );
  AND2_X1 U11202 ( .A1(n11513), .A2(n8798), .ZN(n8801) );
  INV_X1 U11203 ( .A(n8798), .ZN(n8800) );
  AND2_X1 U11204 ( .A1(n11515), .A2(n8799), .ZN(n11553) );
  AND2_X1 U11205 ( .A1(n11553), .A2(n12200), .ZN(n11556) );
  NAND2_X1 U11206 ( .A1(n12894), .A2(n12892), .ZN(n12274) );
  NAND2_X1 U11207 ( .A1(n11685), .A2(n12274), .ZN(n11684) );
  NAND2_X1 U11208 ( .A1(n12512), .A2(n12275), .ZN(n8802) );
  NAND2_X1 U11209 ( .A1(n12876), .A2(n12909), .ZN(n8803) );
  NAND2_X1 U11210 ( .A1(n12902), .A2(n8803), .ZN(n8806) );
  NAND2_X1 U11211 ( .A1(n12511), .A2(n8804), .ZN(n8805) );
  NAND2_X1 U11212 ( .A1(n8806), .A2(n8805), .ZN(n12874) );
  NAND2_X1 U11213 ( .A1(n12510), .A2(n12880), .ZN(n8807) );
  NOR2_X1 U11214 ( .A1(n13052), .A2(n12875), .ZN(n8808) );
  OR2_X1 U11215 ( .A1(n13046), .A2(n12862), .ZN(n8809) );
  OR2_X1 U11216 ( .A1(n12835), .A2(n12845), .ZN(n8810) );
  NAND2_X1 U11217 ( .A1(n12829), .A2(n8810), .ZN(n8812) );
  NAND2_X1 U11218 ( .A1(n12835), .A2(n12845), .ZN(n8811) );
  NAND2_X1 U11219 ( .A1(n8812), .A2(n8811), .ZN(n12817) );
  NAND2_X1 U11220 ( .A1(n12817), .A2(n8813), .ZN(n8815) );
  NAND2_X1 U11221 ( .A1(n12978), .A2(n12805), .ZN(n8814) );
  NAND2_X1 U11222 ( .A1(n8815), .A2(n8814), .ZN(n12804) );
  NAND2_X1 U11223 ( .A1(n12804), .A2(n12211), .ZN(n8817) );
  NAND2_X1 U11224 ( .A1(n12974), .A2(n12818), .ZN(n8816) );
  OR2_X1 U11225 ( .A1(n12789), .A2(n6523), .ZN(n12754) );
  INV_X1 U11226 ( .A(n12774), .ZN(n12507) );
  AND2_X1 U11227 ( .A1(n12954), .A2(n12507), .ZN(n8820) );
  OR2_X1 U11228 ( .A1(n12754), .A2(n8820), .ZN(n12737) );
  OR2_X1 U11229 ( .A1(n12737), .A2(n12743), .ZN(n8818) );
  INV_X1 U11230 ( .A(n12759), .ZN(n12506) );
  OR2_X1 U11231 ( .A1(n12748), .A2(n12506), .ZN(n8821) );
  NAND2_X1 U11232 ( .A1(n12316), .A2(n12317), .ZN(n12779) );
  OR2_X1 U11233 ( .A1(n12967), .A2(n12806), .ZN(n12770) );
  AND2_X1 U11234 ( .A1(n12779), .A2(n12770), .ZN(n12771) );
  OR2_X1 U11235 ( .A1(n8820), .A2(n8819), .ZN(n12738) );
  OR2_X1 U11236 ( .A1(n12743), .A2(n12738), .ZN(n12740) );
  AND2_X1 U11237 ( .A1(n8821), .A2(n12740), .ZN(n8822) );
  NAND2_X1 U11238 ( .A1(n12730), .A2(n12708), .ZN(n8824) );
  NOR2_X1 U11239 ( .A1(n12730), .A2(n12708), .ZN(n8823) );
  NAND2_X1 U11240 ( .A1(n12707), .A2(n12706), .ZN(n12705) );
  NAND2_X1 U11241 ( .A1(n12678), .A2(n12677), .ZN(n12676) );
  NAND2_X1 U11242 ( .A1(n12662), .A2(n8827), .ZN(n8828) );
  NAND2_X1 U11243 ( .A1(n12367), .A2(n12609), .ZN(n8905) );
  NAND2_X1 U11244 ( .A1(n12221), .A2(n8904), .ZN(n12195) );
  INV_X1 U11245 ( .A(n8829), .ZN(n8830) );
  NAND2_X1 U11246 ( .A1(n12503), .A2(n12847), .ZN(n8831) );
  OAI211_X1 U11247 ( .C1(n12384), .C2(n12908), .A(n8832), .B(n8831), .ZN(
        n12639) );
  AOI21_X1 U11248 ( .B1(n12643), .B2(n8900), .A(n12639), .ZN(n13004) );
  NAND2_X1 U11249 ( .A1(n8836), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8837) );
  INV_X1 U11250 ( .A(n8838), .ZN(n8839) );
  NAND2_X1 U11251 ( .A1(n8839), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8840) );
  MUX2_X1 U11252 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8840), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8841) );
  NAND2_X1 U11253 ( .A1(n8841), .A2(n8836), .ZN(n11477) );
  NAND2_X1 U11254 ( .A1(n8842), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8844) );
  INV_X1 U11255 ( .A(n11535), .ZN(n8847) );
  XNOR2_X1 U11256 ( .A(n11255), .B(P3_B_REG_SCAN_IN), .ZN(n8845) );
  NAND2_X1 U11257 ( .A1(n11477), .A2(n8845), .ZN(n8846) );
  NAND2_X1 U11258 ( .A1(n11535), .A2(n11255), .ZN(n8848) );
  NAND2_X1 U11259 ( .A1(n11535), .A2(n11477), .ZN(n8850) );
  NAND2_X1 U11260 ( .A1(n13056), .A2(n13054), .ZN(n8903) );
  INV_X1 U11261 ( .A(n13056), .ZN(n8852) );
  INV_X1 U11262 ( .A(n13054), .ZN(n10706) );
  NAND2_X1 U11263 ( .A1(n8852), .A2(n10706), .ZN(n8907) );
  NOR2_X1 U11264 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n8856) );
  NOR4_X1 U11265 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8855) );
  NOR4_X1 U11266 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8854) );
  NOR4_X1 U11267 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8853) );
  NAND4_X1 U11268 ( .A1(n8856), .A2(n8855), .A3(n8854), .A4(n8853), .ZN(n8862)
         );
  NOR4_X1 U11269 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8860) );
  NOR4_X1 U11270 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8859) );
  NOR4_X1 U11271 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8858) );
  NOR4_X1 U11272 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8857) );
  NAND4_X1 U11273 ( .A1(n8860), .A2(n8859), .A3(n8858), .A4(n8857), .ZN(n8861)
         );
  NOR2_X1 U11274 ( .A1(n8862), .A2(n8861), .ZN(n8863) );
  NAND4_X1 U11275 ( .A1(n10714), .A2(n8903), .A3(n8907), .A4(n8902), .ZN(
        n10712) );
  INV_X1 U11276 ( .A(n10712), .ZN(n8872) );
  OAI22_X1 U11277 ( .A1(n12941), .A2(n8904), .B1(n12609), .B2(n12218), .ZN(
        n8864) );
  NAND2_X1 U11278 ( .A1(n8864), .A2(n8867), .ZN(n8865) );
  NAND2_X1 U11279 ( .A1(n8865), .A2(n12312), .ZN(n8866) );
  NAND2_X1 U11280 ( .A1(n8866), .A2(n10706), .ZN(n8870) );
  INV_X1 U11281 ( .A(n8867), .ZN(n12362) );
  OR2_X1 U11282 ( .A1(n12312), .A2(n12362), .ZN(n9015) );
  NAND2_X1 U11283 ( .A1(n12312), .A2(n8868), .ZN(n10708) );
  NAND2_X1 U11284 ( .A1(n9015), .A2(n10708), .ZN(n10707) );
  NAND2_X1 U11285 ( .A1(n10707), .A2(n13054), .ZN(n8869) );
  OR2_X1 U11286 ( .A1(n13004), .A2(n15014), .ZN(n8877) );
  INV_X1 U11287 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n8873) );
  NOR2_X1 U11288 ( .A1(n15016), .A2(n8873), .ZN(n8874) );
  NAND2_X1 U11289 ( .A1(n8877), .A2(n8876), .ZN(P3_U3487) );
  INV_X1 U11290 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12033) );
  NAND2_X1 U11291 ( .A1(n12033), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8880) );
  NAND2_X1 U11292 ( .A1(n8882), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8883) );
  XNOR2_X1 U11293 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12160) );
  XNOR2_X1 U11294 ( .A(n12162), .B(n12160), .ZN(n11866) );
  NAND2_X1 U11295 ( .A1(n11866), .A2(n12181), .ZN(n8885) );
  NAND2_X1 U11296 ( .A1(n12182), .A2(SI_29_), .ZN(n8884) );
  NAND2_X1 U11297 ( .A1(n12354), .A2(n12350), .ZN(n12196) );
  XNOR2_X1 U11298 ( .A(n8886), .B(n12215), .ZN(n8896) );
  INV_X1 U11299 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n8891) );
  NAND2_X1 U11300 ( .A1(n12172), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8889) );
  NAND2_X1 U11301 ( .A1(n8887), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8888) );
  OAI211_X1 U11302 ( .C1(n8891), .C2(n8890), .A(n8889), .B(n8888), .ZN(n8892)
         );
  INV_X1 U11303 ( .A(n8892), .ZN(n8893) );
  AND2_X1 U11304 ( .A1(n12178), .A2(n8893), .ZN(n12188) );
  INV_X1 U11305 ( .A(P3_B_REG_SCAN_IN), .ZN(n8894) );
  OAI21_X1 U11306 ( .B1(n13068), .B2(n8894), .A(n12846), .ZN(n12631) );
  OAI22_X1 U11307 ( .A1(n12652), .A2(n12906), .B1(n12188), .B2(n12631), .ZN(
        n8895) );
  AND2_X1 U11308 ( .A1(n8898), .A2(n8897), .ZN(n12342) );
  INV_X1 U11309 ( .A(n8899), .ZN(n12341) );
  AOI21_X1 U11310 ( .B1(n12648), .B2(n12342), .A(n12341), .ZN(n12187) );
  INV_X1 U11311 ( .A(n8902), .ZN(n8906) );
  NAND2_X1 U11312 ( .A1(n10714), .A2(n12362), .ZN(n9026) );
  OR2_X1 U11313 ( .A1(n9026), .A2(n12312), .ZN(n9013) );
  NAND2_X1 U11314 ( .A1(n10538), .A2(n8904), .ZN(n12360) );
  OR2_X1 U11315 ( .A1(n8905), .A2(n12360), .ZN(n9014) );
  INV_X1 U11316 ( .A(n9019), .ZN(n8908) );
  OAI22_X1 U11317 ( .A1(n9014), .A2(n9020), .B1(n8908), .B2(n9018), .ZN(n8909)
         );
  NAND2_X1 U11318 ( .A1(n8909), .A2(n10714), .ZN(n8910) );
  NAND2_X1 U11319 ( .A1(n9034), .A2(n15004), .ZN(n8917) );
  NAND2_X1 U11320 ( .A1(n7133), .A2(n8912), .ZN(n8915) );
  INV_X1 U11321 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8913) );
  OR2_X1 U11322 ( .A1(n15004), .A2(n8913), .ZN(n8914) );
  INV_X1 U11323 ( .A(n12360), .ZN(n8918) );
  NAND2_X1 U11324 ( .A1(n13056), .A2(n8918), .ZN(n8921) );
  NAND2_X1 U11325 ( .A1(n10538), .A2(n12609), .ZN(n8919) );
  NAND2_X1 U11326 ( .A1(n8919), .A2(n10455), .ZN(n8920) );
  AND2_X4 U11327 ( .A1(n8921), .A2(n8920), .ZN(n10798) );
  XNOR2_X1 U11328 ( .A(n12339), .B(n10798), .ZN(n12387) );
  NOR2_X1 U11329 ( .A1(n12387), .A2(n12503), .ZN(n12382) );
  AOI21_X1 U11330 ( .B1(n12387), .B2(n12503), .A(n12382), .ZN(n9009) );
  XNOR2_X1 U11331 ( .A(n12978), .B(n12379), .ZN(n8974) );
  INV_X1 U11332 ( .A(n10804), .ZN(n10876) );
  NAND3_X1 U11333 ( .A1(n10876), .A2(n10798), .A3(n12521), .ZN(n10744) );
  NAND2_X1 U11334 ( .A1(n10744), .A2(n8929), .ZN(n8926) );
  NOR2_X1 U11335 ( .A1(n8926), .A2(n12379), .ZN(n8925) );
  NAND2_X1 U11336 ( .A1(n8922), .A2(n12379), .ZN(n8923) );
  OAI211_X1 U11337 ( .C1(n10743), .C2(n12379), .A(n8923), .B(n12520), .ZN(
        n8924) );
  XNOR2_X1 U11338 ( .A(n11062), .B(n12379), .ZN(n10748) );
  INV_X1 U11339 ( .A(n10745), .ZN(n8928) );
  INV_X1 U11340 ( .A(n8926), .ZN(n8927) );
  OAI211_X1 U11341 ( .C1(n10875), .C2(n10748), .A(n8928), .B(n8927), .ZN(n8933) );
  NAND3_X1 U11342 ( .A1(n10872), .A2(n10743), .A3(n10798), .ZN(n8931) );
  NAND4_X1 U11343 ( .A1(n8931), .A2(n8930), .A3(n10875), .A4(n10744), .ZN(
        n8932) );
  NAND3_X1 U11344 ( .A1(n8934), .A2(n8933), .A3(n8932), .ZN(n10781) );
  XNOR2_X1 U11345 ( .A(n10969), .B(n12379), .ZN(n8939) );
  XNOR2_X1 U11346 ( .A(n8939), .B(n12519), .ZN(n10780) );
  OR2_X1 U11347 ( .A1(n10781), .A2(n10780), .ZN(n11033) );
  XNOR2_X1 U11348 ( .A(n11217), .B(n10798), .ZN(n8945) );
  XNOR2_X1 U11349 ( .A(n8945), .B(n10825), .ZN(n11034) );
  XNOR2_X1 U11350 ( .A(n11282), .B(n10798), .ZN(n8935) );
  INV_X1 U11351 ( .A(n11154), .ZN(n8938) );
  INV_X1 U11352 ( .A(n8935), .ZN(n8937) );
  NAND2_X1 U11353 ( .A1(n8937), .A2(n8936), .ZN(n8947) );
  AND2_X1 U11354 ( .A1(n11034), .A2(n8948), .ZN(n11092) );
  NAND2_X1 U11355 ( .A1(n8939), .A2(n12519), .ZN(n11032) );
  XNOR2_X1 U11356 ( .A(n11358), .B(n12379), .ZN(n8944) );
  INV_X1 U11357 ( .A(n8944), .ZN(n8940) );
  NAND2_X1 U11358 ( .A1(n12516), .A2(n8940), .ZN(n8943) );
  INV_X1 U11359 ( .A(n8943), .ZN(n8950) );
  XNOR2_X1 U11360 ( .A(n8944), .B(n11516), .ZN(n11095) );
  INV_X1 U11361 ( .A(n11095), .ZN(n8949) );
  INV_X1 U11362 ( .A(n8945), .ZN(n8946) );
  NAND2_X1 U11363 ( .A1(n8946), .A2(n10825), .ZN(n11152) );
  NAND2_X1 U11364 ( .A1(n7416), .A2(n8948), .ZN(n11094) );
  XNOR2_X1 U11365 ( .A(n11515), .B(n10798), .ZN(n11128) );
  NAND3_X1 U11366 ( .A1(n11127), .A2(n11126), .A3(n11128), .ZN(n11170) );
  INV_X1 U11367 ( .A(n11128), .ZN(n8951) );
  NAND2_X1 U11368 ( .A1(n8951), .A2(n12515), .ZN(n11169) );
  XNOR2_X1 U11369 ( .A(n12270), .B(n12379), .ZN(n8957) );
  XNOR2_X1 U11370 ( .A(n8957), .B(n12513), .ZN(n11234) );
  INV_X1 U11371 ( .A(n11234), .ZN(n8952) );
  XNOR2_X1 U11372 ( .A(n11637), .B(n10798), .ZN(n8954) );
  NAND2_X1 U11373 ( .A1(n12514), .A2(n8954), .ZN(n11229) );
  AND2_X1 U11374 ( .A1(n8952), .A2(n11229), .ZN(n8953) );
  AND2_X1 U11375 ( .A1(n11169), .A2(n8953), .ZN(n8956) );
  INV_X1 U11376 ( .A(n8953), .ZN(n8955) );
  XNOR2_X1 U11377 ( .A(n8954), .B(n11562), .ZN(n11171) );
  INV_X1 U11378 ( .A(n8957), .ZN(n8958) );
  NAND2_X1 U11379 ( .A1(n11174), .A2(n8958), .ZN(n8959) );
  XNOR2_X1 U11380 ( .A(n12275), .B(n10798), .ZN(n8960) );
  XNOR2_X1 U11381 ( .A(n8960), .B(n12905), .ZN(n11345) );
  INV_X1 U11382 ( .A(n8960), .ZN(n8961) );
  OR2_X1 U11383 ( .A1(n8961), .A2(n12905), .ZN(n8962) );
  XNOR2_X1 U11384 ( .A(n12909), .B(n12379), .ZN(n8963) );
  NAND2_X1 U11385 ( .A1(n8964), .A2(n8963), .ZN(n11587) );
  XNOR2_X1 U11386 ( .A(n12880), .B(n12379), .ZN(n8965) );
  XNOR2_X1 U11387 ( .A(n8965), .B(n12907), .ZN(n11621) );
  XNOR2_X1 U11388 ( .A(n13052), .B(n12379), .ZN(n11723) );
  INV_X1 U11389 ( .A(n11723), .ZN(n8967) );
  NAND2_X1 U11390 ( .A1(n12875), .A2(n8967), .ZN(n8968) );
  NAND2_X1 U11391 ( .A1(n11723), .A2(n8969), .ZN(n8970) );
  XNOR2_X1 U11392 ( .A(n13046), .B(n12379), .ZN(n8971) );
  XNOR2_X1 U11393 ( .A(n8971), .B(n12862), .ZN(n12396) );
  XNOR2_X1 U11394 ( .A(n12835), .B(n10798), .ZN(n8973) );
  NOR2_X1 U11395 ( .A1(n8973), .A2(n12845), .ZN(n12486) );
  NAND2_X1 U11396 ( .A1(n8973), .A2(n12845), .ZN(n12487) );
  XNOR2_X1 U11397 ( .A(n8974), .B(n12805), .ZN(n12427) );
  NAND2_X1 U11398 ( .A1(n12428), .A2(n12427), .ZN(n12426) );
  OAI21_X1 U11399 ( .B1(n12832), .B2(n8974), .A(n12426), .ZN(n12435) );
  XNOR2_X1 U11400 ( .A(n12974), .B(n12379), .ZN(n8975) );
  XNOR2_X1 U11401 ( .A(n8975), .B(n12818), .ZN(n12434) );
  INV_X1 U11402 ( .A(n12466), .ZN(n8979) );
  XOR2_X1 U11403 ( .A(n12379), .B(n12967), .Z(n12464) );
  INV_X1 U11404 ( .A(n12464), .ZN(n8978) );
  XNOR2_X1 U11405 ( .A(n13034), .B(n12379), .ZN(n8980) );
  XNOR2_X1 U11406 ( .A(n8980), .B(n12792), .ZN(n12413) );
  NAND2_X1 U11407 ( .A1(n12412), .A2(n12413), .ZN(n8982) );
  NAND2_X1 U11408 ( .A1(n8982), .A2(n8981), .ZN(n12449) );
  XNOR2_X1 U11409 ( .A(n12954), .B(n12379), .ZN(n8983) );
  XNOR2_X1 U11410 ( .A(n8983), .B(n12507), .ZN(n12450) );
  XNOR2_X1 U11411 ( .A(n12748), .B(n12379), .ZN(n8985) );
  NAND2_X1 U11412 ( .A1(n8985), .A2(n12759), .ZN(n8986) );
  OAI21_X1 U11413 ( .B1(n8985), .B2(n12759), .A(n8986), .ZN(n12420) );
  XNOR2_X1 U11414 ( .A(n12730), .B(n12379), .ZN(n8987) );
  NAND2_X1 U11415 ( .A1(n8988), .A2(n8987), .ZN(n8990) );
  OAI21_X1 U11416 ( .B1(n8988), .B2(n8987), .A(n8990), .ZN(n12458) );
  INV_X1 U11417 ( .A(n12458), .ZN(n8989) );
  XNOR2_X1 U11418 ( .A(n12721), .B(n12379), .ZN(n8991) );
  INV_X1 U11419 ( .A(n12728), .ZN(n12505) );
  XNOR2_X1 U11420 ( .A(n12702), .B(n10798), .ZN(n8993) );
  NAND2_X1 U11421 ( .A1(n8993), .A2(n12408), .ZN(n9045) );
  INV_X1 U11422 ( .A(n8993), .ZN(n8994) );
  NAND2_X1 U11423 ( .A1(n8994), .A2(n12709), .ZN(n8995) );
  AND2_X1 U11424 ( .A1(n9045), .A2(n8995), .ZN(n12441) );
  XNOR2_X1 U11425 ( .A(n12933), .B(n12379), .ZN(n8996) );
  NAND2_X1 U11426 ( .A1(n8996), .A2(n12690), .ZN(n9000) );
  INV_X1 U11427 ( .A(n8996), .ZN(n8997) );
  INV_X1 U11428 ( .A(n12690), .ZN(n12504) );
  NAND2_X1 U11429 ( .A1(n8997), .A2(n12504), .ZN(n8998) );
  AND2_X1 U11430 ( .A1(n9000), .A2(n8998), .ZN(n8999) );
  INV_X1 U11431 ( .A(n8999), .ZN(n9044) );
  OR2_X1 U11432 ( .A1(n9044), .A2(n9045), .ZN(n9042) );
  AND2_X1 U11433 ( .A1(n9042), .A2(n9000), .ZN(n12473) );
  XNOR2_X1 U11434 ( .A(n9001), .B(n10798), .ZN(n9005) );
  NOR2_X1 U11435 ( .A1(n9005), .A2(n12679), .ZN(n9004) );
  INV_X1 U11436 ( .A(n9004), .ZN(n9003) );
  AND2_X1 U11437 ( .A1(n12473), .A2(n9003), .ZN(n9002) );
  NAND2_X1 U11438 ( .A1(n12474), .A2(n9002), .ZN(n9008) );
  AOI21_X1 U11439 ( .B1(n9005), .B2(n12679), .A(n9004), .ZN(n12475) );
  OR2_X1 U11440 ( .A1(n9004), .A2(n12475), .ZN(n9006) );
  AND2_X1 U11441 ( .A1(n9006), .A2(n9009), .ZN(n9007) );
  OAI22_X1 U11442 ( .A1(n9020), .A2(n10618), .B1(n9018), .B2(n9014), .ZN(n9010) );
  AND2_X1 U11443 ( .A1(n10714), .A2(n12979), .ZN(n9012) );
  NAND2_X1 U11444 ( .A1(n9020), .A2(n12359), .ZN(n9011) );
  OR2_X1 U11445 ( .A1(n9013), .A2(n9027), .ZN(n9025) );
  INV_X1 U11446 ( .A(n9014), .ZN(n9017) );
  NAND3_X1 U11447 ( .A1(n9015), .A2(n9672), .A3(n10252), .ZN(n9016) );
  AOI21_X1 U11448 ( .B1(n9018), .B2(n9017), .A(n9016), .ZN(n9022) );
  NAND2_X1 U11449 ( .A1(n9020), .A2(n9019), .ZN(n9021) );
  NAND2_X1 U11450 ( .A1(n9022), .A2(n9021), .ZN(n9023) );
  NAND2_X1 U11451 ( .A1(n9023), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9024) );
  NOR2_X1 U11452 ( .A1(n12906), .A2(n9026), .ZN(n12365) );
  NOR2_X1 U11453 ( .A1(n12651), .A2(n12479), .ZN(n9030) );
  INV_X1 U11454 ( .A(n9026), .ZN(n9028) );
  NAND3_X1 U11455 ( .A1(n12846), .A2(n9028), .A3(n9027), .ZN(n12491) );
  INV_X1 U11456 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n15078) );
  OAI22_X1 U11457 ( .A1(n12652), .A2(n12491), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15078), .ZN(n9029) );
  AOI211_X1 U11458 ( .C1(n12657), .C2(n12482), .A(n9030), .B(n9029), .ZN(n9031) );
  INV_X1 U11459 ( .A(n9032), .ZN(n9033) );
  NAND2_X1 U11460 ( .A1(n7133), .A2(n8875), .ZN(n9036) );
  AOI22_X1 U11461 ( .A1(n12709), .A2(n12493), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9040) );
  NAND2_X1 U11462 ( .A1(n12683), .A2(n12482), .ZN(n9039) );
  OAI211_X1 U11463 ( .C1(n12651), .C2(n12491), .A(n9040), .B(n9039), .ZN(n9041) );
  INV_X1 U11464 ( .A(n9041), .ZN(n9050) );
  AND2_X1 U11465 ( .A1(n12474), .A2(n9042), .ZN(n9047) );
  NAND2_X1 U11466 ( .A1(n9043), .A2(n12441), .ZN(n12442) );
  NAND3_X1 U11467 ( .A1(n12442), .A2(n9045), .A3(n9044), .ZN(n9046) );
  INV_X1 U11468 ( .A(n9048), .ZN(n9049) );
  NOR2_X1 U11469 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n9053) );
  NOR2_X2 U11470 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9155) );
  NOR2_X1 U11471 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n9063) );
  NAND4_X1 U11472 ( .A1(n9063), .A2(n9062), .A3(n9061), .A4(n9655), .ZN(n9657)
         );
  NAND2_X1 U11473 ( .A1(n9388), .A2(n9064), .ZN(n9065) );
  INV_X1 U11474 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9068) );
  NAND2_X1 U11475 ( .A1(n9663), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9070) );
  NAND2_X1 U11476 ( .A1(n11864), .A2(n9153), .ZN(n9073) );
  INV_X1 U11477 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n12163) );
  OR2_X1 U11478 ( .A1(n9580), .A2(n12163), .ZN(n9072) );
  NAND2_X1 U11479 ( .A1(n9076), .A2(n9075), .ZN(n14173) );
  NAND2_X1 U11480 ( .A1(n9078), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9079) );
  AOI22_X1 U11481 ( .A1(n9148), .A2(P1_REG1_REG_29__SCAN_IN), .B1(n9574), .B2(
        P1_REG2_REG_29__SCAN_IN), .ZN(n9087) );
  NAND2_X1 U11482 ( .A1(n9200), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9230) );
  NAND2_X1 U11483 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n9083) );
  NOR2_X1 U11484 ( .A1(n9230), .A2(n9083), .ZN(n9250) );
  NAND2_X1 U11485 ( .A1(n9250), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9279) );
  INV_X1 U11486 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9277) );
  NAND2_X1 U11487 ( .A1(n9327), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9329) );
  INV_X1 U11488 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9406) );
  INV_X1 U11489 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9418) );
  INV_X1 U11490 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13671) );
  NAND2_X1 U11491 ( .A1(n9438), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9439) );
  NAND2_X1 U11492 ( .A1(n9471), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U11493 ( .A1(n9486), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9485) );
  NAND2_X1 U11494 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n9497), .ZN(n9515) );
  INV_X1 U11495 ( .A(n9515), .ZN(n9084) );
  NAND2_X1 U11496 ( .A1(n9084), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9528) );
  INV_X1 U11497 ( .A(n9528), .ZN(n9085) );
  NAND2_X1 U11498 ( .A1(n9085), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9546) );
  INV_X1 U11499 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n12152) );
  NOR2_X1 U11500 ( .A1(n9546), .A2(n12152), .ZN(n13860) );
  AOI22_X1 U11501 ( .A1(n9575), .A2(P1_REG0_REG_29__SCAN_IN), .B1(n9441), .B2(
        n13860), .ZN(n9086) );
  AND2_X1 U11502 ( .A1(n9087), .A2(n9086), .ZN(n9561) );
  INV_X1 U11503 ( .A(n9090), .ZN(n9088) );
  NAND2_X1 U11504 ( .A1(n9090), .A2(n9089), .ZN(n9099) );
  INV_X1 U11505 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9093) );
  NAND4_X1 U11506 ( .A1(n9096), .A2(n7352), .A3(n9388), .A4(n9093), .ZN(n9094)
         );
  NAND2_X1 U11507 ( .A1(n9646), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9097) );
  NAND2_X1 U11508 ( .A1(n9099), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9101) );
  MUX2_X1 U11509 ( .A(n13855), .B(n9561), .S(n9143), .Z(n9560) );
  INV_X1 U11510 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9103) );
  NAND2_X1 U11511 ( .A1(n9133), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9107) );
  INV_X1 U11512 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n14056) );
  OR2_X1 U11513 ( .A1(n9137), .A2(n14056), .ZN(n9106) );
  INV_X1 U11514 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9104) );
  OR2_X1 U11515 ( .A1(n9134), .A2(n9104), .ZN(n9105) );
  INV_X1 U11516 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9110) );
  NAND2_X1 U11517 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9109) );
  XNOR2_X1 U11518 ( .A(n9110), .B(n9109), .ZN(n13761) );
  NAND2_X2 U11519 ( .A1(n6571), .A2(n9112), .ZN(n14586) );
  INV_X1 U11520 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9113) );
  OR2_X1 U11521 ( .A1(n9136), .A2(n9113), .ZN(n9119) );
  INV_X1 U11522 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9114) );
  OR2_X1 U11523 ( .A1(n9134), .A2(n9114), .ZN(n9117) );
  INV_X1 U11524 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9115) );
  NOR2_X1 U11525 ( .A1(n9678), .A2(n9714), .ZN(n9121) );
  XNOR2_X1 U11526 ( .A(n9121), .B(n9120), .ZN(n14191) );
  INV_X1 U11527 ( .A(n14565), .ZN(n10218) );
  NAND2_X1 U11528 ( .A1(n9606), .A2(n10016), .ZN(n9122) );
  NAND2_X1 U11529 ( .A1(n14047), .A2(n14565), .ZN(n10231) );
  NAND3_X1 U11530 ( .A1(n9122), .A2(n10231), .A3(n6472), .ZN(n9123) );
  NAND2_X1 U11531 ( .A1(n10014), .A2(n14586), .ZN(n10230) );
  NAND2_X1 U11532 ( .A1(n9123), .A2(n10230), .ZN(n9126) );
  INV_X1 U11533 ( .A(n10230), .ZN(n9124) );
  NAND2_X1 U11534 ( .A1(n9124), .A2(n6472), .ZN(n9125) );
  INV_X1 U11535 ( .A(n10231), .ZN(n9127) );
  NAND2_X1 U11536 ( .A1(n9129), .A2(n6492), .ZN(n9132) );
  OR2_X1 U11537 ( .A1(n9155), .A2(n9068), .ZN(n9131) );
  XNOR2_X1 U11538 ( .A(n9131), .B(P1_IR_REG_2__SCAN_IN), .ZN(n13775) );
  NAND2_X1 U11539 ( .A1(n10490), .A2(n9143), .ZN(n9142) );
  NAND2_X1 U11540 ( .A1(n9133), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9141) );
  INV_X1 U11541 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10488) );
  OR2_X1 U11542 ( .A1(n9134), .A2(n10488), .ZN(n9140) );
  INV_X1 U11543 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9135) );
  OR2_X1 U11544 ( .A1(n9569), .A2(n9135), .ZN(n9139) );
  INV_X1 U11545 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9778) );
  OR2_X1 U11546 ( .A1(n9567), .A2(n9778), .ZN(n9138) );
  NAND2_X1 U11547 ( .A1(n9142), .A2(n7406), .ZN(n9146) );
  BUF_X8 U11548 ( .A(n9143), .Z(n9585) );
  OAI21_X1 U11549 ( .B1(n10490), .B2(n9585), .A(n9144), .ZN(n9145) );
  NAND3_X1 U11550 ( .A1(n9147), .A2(n10490), .A3(n9146), .ZN(n9161) );
  INV_X1 U11551 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9780) );
  OR2_X1 U11552 ( .A1(n9567), .A2(n9780), .ZN(n9151) );
  OR2_X1 U11553 ( .A1(n9134), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9149) );
  NAND3_X2 U11554 ( .A1(n9152), .A2(n9151), .A3(n7422), .ZN(n13754) );
  NAND2_X1 U11555 ( .A1(n9683), .A2(n6492), .ZN(n9160) );
  INV_X1 U11556 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9154) );
  NAND2_X1 U11557 ( .A1(n9155), .A2(n9154), .ZN(n9157) );
  NAND2_X1 U11558 ( .A1(n9157), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9156) );
  MUX2_X1 U11559 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9156), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9158) );
  OR2_X1 U11560 ( .A1(n9157), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n9190) );
  AND2_X1 U11561 ( .A1(n9158), .A2(n9190), .ZN(n13788) );
  AOI22_X1 U11562 ( .A1(n9415), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n9414), .B2(
        n13788), .ZN(n9159) );
  XNOR2_X2 U11563 ( .A(n13754), .B(n14554), .ZN(n10226) );
  NAND3_X1 U11564 ( .A1(n9162), .A2(n9161), .A3(n10226), .ZN(n9166) );
  NAND2_X1 U11565 ( .A1(n13754), .A2(n9143), .ZN(n9164) );
  INV_X1 U11566 ( .A(n13754), .ZN(n10235) );
  NAND2_X1 U11567 ( .A1(n10235), .A2(n6472), .ZN(n9163) );
  NAND2_X1 U11568 ( .A1(n9166), .A2(n9165), .ZN(n9177) );
  OR2_X1 U11569 ( .A1(n9691), .A2(n9111), .ZN(n9169) );
  NAND2_X1 U11570 ( .A1(n9190), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9167) );
  XNOR2_X1 U11571 ( .A(n9167), .B(P1_IR_REG_4__SCAN_IN), .ZN(n14491) );
  AOI22_X1 U11572 ( .A1(n9415), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9414), .B2(
        n14491), .ZN(n9168) );
  NAND2_X1 U11573 ( .A1(n9575), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9174) );
  INV_X1 U11574 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9170) );
  OR2_X1 U11575 ( .A1(n9579), .A2(n9170), .ZN(n9173) );
  XNOR2_X1 U11576 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n14527) );
  OR2_X1 U11577 ( .A1(n9547), .A2(n14527), .ZN(n9172) );
  INV_X1 U11578 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n14528) );
  OR2_X1 U11579 ( .A1(n9567), .A2(n14528), .ZN(n9171) );
  MUX2_X1 U11580 ( .A(n10674), .B(n13753), .S(n9585), .Z(n9178) );
  NAND2_X1 U11581 ( .A1(n9177), .A2(n9178), .ZN(n9176) );
  MUX2_X1 U11582 ( .A(n13753), .B(n10674), .S(n9585), .Z(n9175) );
  NAND2_X1 U11583 ( .A1(n9176), .A2(n9175), .ZN(n9182) );
  INV_X1 U11584 ( .A(n9177), .ZN(n9180) );
  INV_X1 U11585 ( .A(n9178), .ZN(n9179) );
  NAND2_X1 U11586 ( .A1(n9180), .A2(n9179), .ZN(n9181) );
  AOI21_X1 U11587 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9183) );
  NOR2_X1 U11588 ( .A1(n9183), .A2(n9200), .ZN(n10648) );
  NAND2_X1 U11589 ( .A1(n9441), .A2(n10648), .ZN(n9189) );
  INV_X1 U11590 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9184) );
  OR2_X1 U11591 ( .A1(n9567), .A2(n9184), .ZN(n9188) );
  OR2_X1 U11592 ( .A1(n9579), .A2(n10470), .ZN(n9187) );
  INV_X1 U11593 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9185) );
  OR2_X1 U11594 ( .A1(n9569), .A2(n9185), .ZN(n9186) );
  NAND2_X1 U11595 ( .A1(n9717), .A2(n9153), .ZN(n9193) );
  OAI21_X1 U11596 ( .B1(n9190), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9191) );
  XNOR2_X1 U11597 ( .A(n9191), .B(P1_IR_REG_5__SCAN_IN), .ZN(n13798) );
  AOI22_X1 U11598 ( .A1(n9415), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9414), .B2(
        n13798), .ZN(n9192) );
  MUX2_X1 U11599 ( .A(n13752), .B(n10692), .S(n9585), .Z(n9195) );
  MUX2_X1 U11600 ( .A(n10692), .B(n13752), .S(n9585), .Z(n9194) );
  INV_X1 U11601 ( .A(n9195), .ZN(n9196) );
  NAND2_X1 U11602 ( .A1(n9742), .A2(n9153), .ZN(n9199) );
  NAND2_X1 U11603 ( .A1(n9216), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9197) );
  XNOR2_X1 U11604 ( .A(n9197), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9797) );
  AOI22_X1 U11605 ( .A1(n9415), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9414), .B2(
        n9797), .ZN(n9198) );
  NAND2_X1 U11606 ( .A1(n9199), .A2(n9198), .ZN(n14607) );
  NAND2_X1 U11607 ( .A1(n9575), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9204) );
  INV_X1 U11608 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9803) );
  OR2_X1 U11609 ( .A1(n9579), .A2(n9803), .ZN(n9203) );
  OAI21_X1 U11610 ( .B1(n9200), .B2(P1_REG3_REG_6__SCAN_IN), .A(n9230), .ZN(
        n13713) );
  OR2_X1 U11611 ( .A1(n9547), .A2(n13713), .ZN(n9202) );
  INV_X1 U11612 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9786) );
  OR2_X1 U11613 ( .A1(n9567), .A2(n9786), .ZN(n9201) );
  NAND4_X1 U11614 ( .A1(n9204), .A2(n9203), .A3(n9202), .A4(n9201), .ZN(n13751) );
  MUX2_X1 U11615 ( .A(n14607), .B(n13751), .S(n9585), .Z(n9208) );
  NAND2_X1 U11616 ( .A1(n9207), .A2(n9208), .ZN(n9206) );
  MUX2_X1 U11617 ( .A(n14607), .B(n13751), .S(n6472), .Z(n9205) );
  INV_X1 U11618 ( .A(n9207), .ZN(n9210) );
  INV_X1 U11619 ( .A(n9208), .ZN(n9209) );
  NAND2_X1 U11620 ( .A1(n9210), .A2(n9209), .ZN(n9226) );
  NAND2_X1 U11621 ( .A1(n9223), .A2(n9226), .ZN(n9220) );
  NAND2_X1 U11622 ( .A1(n9574), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9215) );
  INV_X1 U11623 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9806) );
  OR2_X1 U11624 ( .A1(n9579), .A2(n9806), .ZN(n9214) );
  INV_X1 U11625 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9878) );
  XNOR2_X1 U11626 ( .A(n9230), .B(n9878), .ZN(n11025) );
  OR2_X1 U11627 ( .A1(n9547), .A2(n11025), .ZN(n9213) );
  INV_X1 U11628 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9211) );
  OR2_X1 U11629 ( .A1(n9569), .A2(n9211), .ZN(n9212) );
  NAND4_X1 U11630 ( .A1(n9215), .A2(n9214), .A3(n9213), .A4(n9212), .ZN(n13750) );
  NAND2_X1 U11631 ( .A1(n9746), .A2(n9153), .ZN(n9219) );
  OR2_X1 U11632 ( .A1(n9216), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9237) );
  NAND2_X1 U11633 ( .A1(n9237), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9217) );
  XNOR2_X1 U11634 ( .A(n9217), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9805) );
  AOI22_X1 U11635 ( .A1(n9415), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9414), .B2(
        n9805), .ZN(n9218) );
  NAND2_X1 U11636 ( .A1(n9219), .A2(n9218), .ZN(n11021) );
  MUX2_X1 U11637 ( .A(n13750), .B(n11021), .S(n9585), .Z(n9224) );
  NAND2_X1 U11638 ( .A1(n9220), .A2(n9224), .ZN(n9222) );
  MUX2_X1 U11639 ( .A(n13750), .B(n11021), .S(n6472), .Z(n9221) );
  NAND2_X1 U11640 ( .A1(n9222), .A2(n9221), .ZN(n9229) );
  INV_X1 U11641 ( .A(n9224), .ZN(n9225) );
  AND2_X1 U11642 ( .A1(n9226), .A2(n9225), .ZN(n9227) );
  NAND2_X1 U11643 ( .A1(n9223), .A2(n9227), .ZN(n9228) );
  NAND2_X1 U11644 ( .A1(n9575), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9236) );
  INV_X1 U11645 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9807) );
  OR2_X1 U11646 ( .A1(n9579), .A2(n9807), .ZN(n9235) );
  INV_X1 U11647 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9799) );
  OR2_X1 U11648 ( .A1(n9567), .A2(n9799), .ZN(n9234) );
  INV_X1 U11649 ( .A(n9230), .ZN(n9231) );
  AOI21_X1 U11650 ( .B1(n9231), .B2(P1_REG3_REG_7__SCAN_IN), .A(
        P1_REG3_REG_8__SCAN_IN), .ZN(n9232) );
  OR2_X1 U11651 ( .A1(n9232), .A2(n9250), .ZN(n11212) );
  OR2_X1 U11652 ( .A1(n9547), .A2(n11212), .ZN(n9233) );
  NAND4_X1 U11653 ( .A1(n9236), .A2(n9235), .A3(n9234), .A4(n9233), .ZN(n13749) );
  NAND2_X1 U11654 ( .A1(n9751), .A2(n9153), .ZN(n9240) );
  OR2_X1 U11655 ( .A1(n9352), .A2(n9068), .ZN(n9238) );
  XNOR2_X1 U11656 ( .A(n9238), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9808) );
  AOI22_X1 U11657 ( .A1(n9415), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9414), .B2(
        n9808), .ZN(n9239) );
  MUX2_X1 U11658 ( .A(n13749), .B(n11200), .S(n6472), .Z(n9244) );
  NAND2_X1 U11659 ( .A1(n9243), .A2(n9244), .ZN(n9242) );
  MUX2_X1 U11660 ( .A(n13749), .B(n11200), .S(n9143), .Z(n9241) );
  NAND2_X1 U11661 ( .A1(n9242), .A2(n9241), .ZN(n9248) );
  INV_X1 U11662 ( .A(n9243), .ZN(n9246) );
  INV_X1 U11663 ( .A(n9244), .ZN(n9245) );
  NAND2_X1 U11664 ( .A1(n9246), .A2(n9245), .ZN(n9247) );
  NAND2_X1 U11665 ( .A1(n9575), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9255) );
  INV_X1 U11666 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9249) );
  OR2_X1 U11667 ( .A1(n9579), .A2(n9249), .ZN(n9254) );
  INV_X1 U11668 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11002) );
  OR2_X1 U11669 ( .A1(n9567), .A2(n11002), .ZN(n9253) );
  OR2_X1 U11670 ( .A1(n9250), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9251) );
  NAND2_X1 U11671 ( .A1(n9279), .A2(n9251), .ZN(n11470) );
  OR2_X1 U11672 ( .A1(n9547), .A2(n11470), .ZN(n9252) );
  NAND4_X1 U11673 ( .A1(n9255), .A2(n9254), .A3(n9253), .A4(n9252), .ZN(n13748) );
  OR2_X1 U11674 ( .A1(n9758), .A2(n9111), .ZN(n9261) );
  INV_X1 U11675 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9256) );
  NAND2_X1 U11676 ( .A1(n9352), .A2(n9256), .ZN(n9258) );
  NAND2_X1 U11677 ( .A1(n9258), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9257) );
  MUX2_X1 U11678 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9257), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n9259) );
  AND2_X1 U11679 ( .A1(n9259), .A2(n9285), .ZN(n9909) );
  AOI22_X1 U11680 ( .A1(n9415), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9414), .B2(
        n9909), .ZN(n9260) );
  NAND2_X2 U11681 ( .A1(n9261), .A2(n9260), .ZN(n11466) );
  MUX2_X1 U11682 ( .A(n13748), .B(n11466), .S(n9143), .Z(n9263) );
  MUX2_X1 U11683 ( .A(n11466), .B(n13748), .S(n9585), .Z(n9262) );
  INV_X1 U11684 ( .A(n9263), .ZN(n9264) );
  NAND2_X1 U11685 ( .A1(n9574), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9270) );
  INV_X1 U11686 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9265) );
  OR2_X1 U11687 ( .A1(n9579), .A2(n9265), .ZN(n9269) );
  XNOR2_X1 U11688 ( .A(n9279), .B(n9278), .ZN(n11608) );
  OR2_X1 U11689 ( .A1(n9547), .A2(n11608), .ZN(n9268) );
  INV_X1 U11690 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9266) );
  OR2_X1 U11691 ( .A1(n9569), .A2(n9266), .ZN(n9267) );
  NAND4_X1 U11692 ( .A1(n9270), .A2(n9269), .A3(n9268), .A4(n9267), .ZN(n13747) );
  NAND2_X1 U11693 ( .A1(n9761), .A2(n9153), .ZN(n9273) );
  NAND2_X1 U11694 ( .A1(n9285), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9271) );
  XNOR2_X1 U11695 ( .A(n9271), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9930) );
  AOI22_X1 U11696 ( .A1(n9415), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9414), 
        .B2(n9930), .ZN(n9272) );
  MUX2_X1 U11697 ( .A(n13747), .B(n11605), .S(n6472), .Z(n9275) );
  MUX2_X1 U11698 ( .A(n13747), .B(n11605), .S(n9585), .Z(n9292) );
  AND2_X1 U11699 ( .A1(n9293), .A2(n9292), .ZN(n9291) );
  NAND2_X1 U11700 ( .A1(n9575), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9284) );
  INV_X1 U11701 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9276) );
  OR2_X1 U11702 ( .A1(n9579), .A2(n9276), .ZN(n9283) );
  OAI21_X1 U11703 ( .B1(n9279), .B2(n9278), .A(n9277), .ZN(n9280) );
  NAND2_X1 U11704 ( .A1(n9280), .A2(n9299), .ZN(n14435) );
  OR2_X1 U11705 ( .A1(n9547), .A2(n14435), .ZN(n9282) );
  INV_X1 U11706 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11121) );
  OR2_X1 U11707 ( .A1(n9567), .A2(n11121), .ZN(n9281) );
  NAND4_X1 U11708 ( .A1(n9284), .A2(n9283), .A3(n9282), .A4(n9281), .ZN(n13746) );
  NAND2_X1 U11709 ( .A1(n9890), .A2(n9153), .ZN(n9288) );
  NOR2_X1 U11710 ( .A1(n9285), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n9307) );
  OR2_X1 U11711 ( .A1(n9307), .A2(n9068), .ZN(n9286) );
  XNOR2_X1 U11712 ( .A(n9286), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10001) );
  AOI22_X1 U11713 ( .A1(n9415), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9414), 
        .B2(n10001), .ZN(n9287) );
  MUX2_X1 U11714 ( .A(n13746), .B(n14431), .S(n9585), .Z(n9297) );
  INV_X1 U11715 ( .A(n9297), .ZN(n9289) );
  NAND2_X1 U11716 ( .A1(n9294), .A2(n9289), .ZN(n9290) );
  NAND2_X1 U11717 ( .A1(n9293), .A2(n9292), .ZN(n9295) );
  NAND2_X1 U11718 ( .A1(n9295), .A2(n9294), .ZN(n9298) );
  INV_X1 U11719 ( .A(n13746), .ZN(n11312) );
  INV_X1 U11720 ( .A(n14431), .ZN(n14448) );
  MUX2_X1 U11721 ( .A(n11312), .B(n14448), .S(n6472), .Z(n9296) );
  NAND2_X1 U11722 ( .A1(n9575), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9305) );
  INV_X1 U11723 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11320) );
  OR2_X1 U11724 ( .A1(n9567), .A2(n11320), .ZN(n9304) );
  INV_X1 U11725 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9995) );
  OR2_X1 U11726 ( .A1(n9579), .A2(n9995), .ZN(n9303) );
  INV_X1 U11727 ( .A(n9327), .ZN(n9301) );
  NAND2_X1 U11728 ( .A1(n9299), .A2(n11811), .ZN(n9300) );
  NAND2_X1 U11729 ( .A1(n9301), .A2(n9300), .ZN(n11810) );
  OR2_X1 U11730 ( .A1(n9547), .A2(n11810), .ZN(n9302) );
  NAND2_X1 U11731 ( .A1(n10011), .A2(n9153), .ZN(n9310) );
  NAND2_X1 U11732 ( .A1(n9307), .A2(n9306), .ZN(n9308) );
  NAND2_X1 U11733 ( .A1(n9308), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9314) );
  XNOR2_X1 U11734 ( .A(n9314), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10275) );
  AOI22_X1 U11735 ( .A1(n9415), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n10275), 
        .B2(n9414), .ZN(n9309) );
  MUX2_X1 U11736 ( .A(n14421), .B(n11816), .S(n9585), .Z(n9341) );
  INV_X1 U11737 ( .A(n14421), .ZN(n13745) );
  MUX2_X1 U11738 ( .A(n13745), .B(n11503), .S(n6472), .Z(n9340) );
  OAI22_X1 U11739 ( .A1(n9312), .A2(n9311), .B1(n9341), .B2(n9340), .ZN(n9345)
         );
  NAND2_X1 U11740 ( .A1(n10430), .A2(n9153), .ZN(n9319) );
  INV_X1 U11741 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9313) );
  NAND2_X1 U11742 ( .A1(n9314), .A2(n9313), .ZN(n9315) );
  NAND2_X1 U11743 ( .A1(n9315), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9336) );
  INV_X1 U11744 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9335) );
  NAND2_X1 U11745 ( .A1(n9336), .A2(n9335), .ZN(n9316) );
  NAND2_X1 U11746 ( .A1(n9316), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9317) );
  XNOR2_X1 U11747 ( .A(n9317), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11133) );
  AOI22_X1 U11748 ( .A1(n11133), .A2(n9414), .B1(n9415), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9318) );
  NAND2_X1 U11749 ( .A1(n9575), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9326) );
  NAND2_X1 U11750 ( .A1(n9329), .A2(n9320), .ZN(n9321) );
  NAND2_X1 U11751 ( .A1(n9357), .A2(n9321), .ZN(n14418) );
  OR2_X1 U11752 ( .A1(n9547), .A2(n14418), .ZN(n9325) );
  INV_X1 U11753 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11676) );
  OR2_X1 U11754 ( .A1(n9567), .A2(n11676), .ZN(n9324) );
  INV_X1 U11755 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9322) );
  OR2_X1 U11756 ( .A1(n9579), .A2(n9322), .ZN(n9323) );
  NAND4_X1 U11757 ( .A1(n9326), .A2(n9325), .A3(n9324), .A4(n9323), .ZN(n13743) );
  NAND2_X1 U11758 ( .A1(n9575), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9334) );
  INV_X1 U11759 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10269) );
  OR2_X1 U11760 ( .A1(n9579), .A2(n10269), .ZN(n9333) );
  OR2_X1 U11761 ( .A1(n9327), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9328) );
  NAND2_X1 U11762 ( .A1(n9329), .A2(n9328), .ZN(n13681) );
  OR2_X1 U11763 ( .A1(n9547), .A2(n13681), .ZN(n9332) );
  INV_X1 U11764 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9330) );
  OR2_X1 U11765 ( .A1(n9567), .A2(n9330), .ZN(n9331) );
  NAND2_X1 U11766 ( .A1(n10108), .A2(n9153), .ZN(n9339) );
  XNOR2_X1 U11767 ( .A(n9336), .B(n9335), .ZN(n11881) );
  OAI22_X1 U11768 ( .A1(n11881), .A2(n9733), .B1(n9580), .B2(n10109), .ZN(
        n9337) );
  INV_X1 U11769 ( .A(n9337), .ZN(n9338) );
  MUX2_X1 U11770 ( .A(n12038), .B(n14443), .S(n9585), .Z(n9346) );
  MUX2_X1 U11771 ( .A(n13744), .B(n11671), .S(n6472), .Z(n9342) );
  AOI22_X1 U11772 ( .A1(n9346), .A2(n9342), .B1(n9341), .B2(n9340), .ZN(n9343)
         );
  NAND2_X1 U11773 ( .A1(n9345), .A2(n9344), .ZN(n9369) );
  INV_X1 U11774 ( .A(n9346), .ZN(n9349) );
  NAND2_X1 U11775 ( .A1(n13744), .A2(n9585), .ZN(n9348) );
  NAND2_X1 U11776 ( .A1(n11671), .A2(n6472), .ZN(n9347) );
  INV_X1 U11777 ( .A(n14411), .ZN(n9366) );
  NAND2_X1 U11778 ( .A1(n10534), .A2(n9153), .ZN(n9355) );
  NAND2_X1 U11779 ( .A1(n9352), .A2(n9351), .ZN(n9379) );
  NAND2_X1 U11780 ( .A1(n9379), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9353) );
  XNOR2_X1 U11781 ( .A(n9353), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11142) );
  AOI22_X1 U11782 ( .A1(n9415), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9414), 
        .B2(n11142), .ZN(n9354) );
  AND2_X1 U11783 ( .A1(n9357), .A2(n9356), .ZN(n9358) );
  NOR2_X1 U11784 ( .A1(n9374), .A2(n9358), .ZN(n13734) );
  NAND2_X1 U11785 ( .A1(n9441), .A2(n13734), .ZN(n9365) );
  INV_X1 U11786 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9359) );
  OR2_X1 U11787 ( .A1(n9567), .A2(n9359), .ZN(n9364) );
  INV_X1 U11788 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9360) );
  OR2_X1 U11789 ( .A1(n9579), .A2(n9360), .ZN(n9363) );
  INV_X1 U11790 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9361) );
  OR2_X1 U11791 ( .A1(n9569), .A2(n9361), .ZN(n9362) );
  NAND2_X1 U11792 ( .A1(n12053), .A2(n12057), .ZN(n9604) );
  OAI21_X1 U11793 ( .B1(n9366), .B2(n13743), .A(n9604), .ZN(n9367) );
  NAND2_X1 U11794 ( .A1(n9369), .A2(n9368), .ZN(n9371) );
  INV_X1 U11795 ( .A(n13743), .ZN(n13731) );
  OR2_X1 U11796 ( .A1(n14411), .A2(n13731), .ZN(n11712) );
  AOI21_X1 U11797 ( .B1(n11738), .B2(n11712), .A(n9585), .ZN(n9370) );
  INV_X1 U11798 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11263) );
  NAND2_X1 U11799 ( .A1(n9574), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9373) );
  OAI21_X1 U11800 ( .B1(n9579), .B2(n11263), .A(n9373), .ZN(n9378) );
  NOR2_X1 U11801 ( .A1(n9374), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9375) );
  OR2_X1 U11802 ( .A1(n9393), .A2(n9375), .ZN(n13644) );
  NAND2_X1 U11803 ( .A1(n9575), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9376) );
  OAI21_X1 U11804 ( .B1(n13644), .B2(n9547), .A(n9376), .ZN(n9377) );
  NAND2_X1 U11805 ( .A1(n10681), .A2(n9153), .ZN(n9382) );
  OAI21_X1 U11806 ( .B1(n9379), .B2(P1_IR_REG_15__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9380) );
  XNOR2_X1 U11807 ( .A(n9380), .B(P1_IR_REG_16__SCAN_IN), .ZN(n11145) );
  AOI22_X1 U11808 ( .A1(n9415), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9414), 
        .B2(n11145), .ZN(n9381) );
  MUX2_X1 U11809 ( .A(n12062), .B(n14152), .S(n9585), .Z(n9384) );
  MUX2_X1 U11810 ( .A(n14032), .B(n13646), .S(n6472), .Z(n9383) );
  NAND2_X1 U11811 ( .A1(n9385), .A2(n9384), .ZN(n9386) );
  NAND2_X1 U11812 ( .A1(n9387), .A2(n9386), .ZN(n9401) );
  NAND2_X1 U11813 ( .A1(n10813), .A2(n9153), .ZN(n9392) );
  OR2_X1 U11814 ( .A1(n9092), .A2(n9068), .ZN(n9389) );
  XNOR2_X1 U11815 ( .A(n9389), .B(n9388), .ZN(n13817) );
  INV_X1 U11816 ( .A(n13817), .ZN(n9390) );
  AOI22_X1 U11817 ( .A1(n9415), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9414), 
        .B2(n9390), .ZN(n9391) );
  NAND2_X2 U11818 ( .A1(n9392), .A2(n9391), .ZN(n14147) );
  OR2_X1 U11819 ( .A1(n9393), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9394) );
  NAND2_X1 U11820 ( .A1(n9407), .A2(n9394), .ZN(n14040) );
  INV_X1 U11821 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14041) );
  OR2_X1 U11822 ( .A1(n9567), .A2(n14041), .ZN(n9396) );
  INV_X1 U11823 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n13812) );
  OR2_X1 U11824 ( .A1(n9579), .A2(n13812), .ZN(n9395) );
  AND2_X1 U11825 ( .A1(n9396), .A2(n9395), .ZN(n9398) );
  NAND2_X1 U11826 ( .A1(n9575), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9397) );
  OAI211_X1 U11827 ( .C1(n14040), .C2(n9547), .A(n9398), .B(n9397), .ZN(n14013) );
  AND2_X1 U11828 ( .A1(n14147), .A2(n14013), .ZN(n11898) );
  MUX2_X1 U11829 ( .A(n14013), .B(n14147), .S(n9585), .Z(n9399) );
  OR2_X1 U11830 ( .A1(n14147), .A2(n14013), .ZN(n11897) );
  NAND2_X1 U11831 ( .A1(n11105), .A2(n9153), .ZN(n9405) );
  NAND2_X1 U11832 ( .A1(n9402), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9403) );
  XNOR2_X1 U11833 ( .A(n9403), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13819) );
  AOI22_X1 U11834 ( .A1(n9415), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9414), 
        .B2(n13819), .ZN(n9404) );
  INV_X1 U11835 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14018) );
  NAND2_X1 U11836 ( .A1(n9407), .A2(n9406), .ZN(n9408) );
  NAND2_X1 U11837 ( .A1(n9419), .A2(n9408), .ZN(n14017) );
  OR2_X1 U11838 ( .A1(n14017), .A2(n9547), .ZN(n9410) );
  AOI22_X1 U11839 ( .A1(n9148), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9575), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n9409) );
  OAI211_X1 U11840 ( .C1(n9567), .C2(n14018), .A(n9410), .B(n9409), .ZN(n14034) );
  NAND2_X1 U11841 ( .A1(n14141), .A2(n9585), .ZN(n9412) );
  OR2_X1 U11842 ( .A1(n14141), .A2(n9143), .ZN(n9411) );
  MUX2_X1 U11843 ( .A(n9412), .B(n9411), .S(n14034), .Z(n9413) );
  NAND2_X1 U11844 ( .A1(n11161), .A2(n9153), .ZN(n9417) );
  AOI22_X1 U11845 ( .A1(n9415), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n13826), 
        .B2(n9414), .ZN(n9416) );
  NAND2_X2 U11846 ( .A1(n9417), .A2(n9416), .ZN(n14136) );
  NAND2_X1 U11847 ( .A1(n9419), .A2(n9418), .ZN(n9420) );
  NAND2_X1 U11848 ( .A1(n9426), .A2(n9420), .ZN(n14004) );
  AOI22_X1 U11849 ( .A1(n9148), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n9574), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n9422) );
  NAND2_X1 U11850 ( .A1(n9575), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9421) );
  OAI211_X1 U11851 ( .C1(n14004), .C2(n9547), .A(n9422), .B(n9421), .ZN(n14021) );
  OR2_X1 U11852 ( .A1(n14136), .A2(n11900), .ZN(n9423) );
  NAND2_X1 U11853 ( .A1(n14136), .A2(n11900), .ZN(n11885) );
  MUX2_X1 U11854 ( .A(n11885), .B(n9423), .S(n6472), .Z(n9424) );
  NAND2_X1 U11855 ( .A1(n9425), .A2(n9424), .ZN(n9436) );
  AND2_X1 U11856 ( .A1(n9426), .A2(n13671), .ZN(n9427) );
  OR2_X1 U11857 ( .A1(n9427), .A2(n9438), .ZN(n13987) );
  INV_X1 U11858 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9430) );
  NAND2_X1 U11859 ( .A1(n9574), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9429) );
  NAND2_X1 U11860 ( .A1(n9575), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9428) );
  OAI211_X1 U11861 ( .C1(n9579), .C2(n9430), .A(n9429), .B(n9428), .ZN(n9431)
         );
  INV_X1 U11862 ( .A(n9431), .ZN(n9432) );
  OAI21_X1 U11863 ( .B1(n13987), .B2(n9547), .A(n9432), .ZN(n13998) );
  NAND2_X1 U11864 ( .A1(n11166), .A2(n9153), .ZN(n9434) );
  INV_X1 U11865 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11167) );
  OR2_X1 U11866 ( .A1(n9580), .A2(n11167), .ZN(n9433) );
  MUX2_X1 U11867 ( .A(n13998), .B(n14130), .S(n9585), .Z(n9437) );
  MUX2_X1 U11868 ( .A(n13998), .B(n14130), .S(n6472), .Z(n9435) );
  OR2_X1 U11869 ( .A1(n9438), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9440) );
  AND2_X1 U11870 ( .A1(n9440), .A2(n9439), .ZN(n13969) );
  NAND2_X1 U11871 ( .A1(n13969), .A2(n9441), .ZN(n9447) );
  INV_X1 U11872 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9444) );
  NAND2_X1 U11873 ( .A1(n9574), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9443) );
  NAND2_X1 U11874 ( .A1(n9575), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9442) );
  OAI211_X1 U11875 ( .C1(n9579), .C2(n9444), .A(n9443), .B(n9442), .ZN(n9445)
         );
  INV_X1 U11876 ( .A(n9445), .ZN(n9446) );
  NAND2_X1 U11877 ( .A1(n9447), .A2(n9446), .ZN(n13953) );
  NAND2_X1 U11878 ( .A1(n11256), .A2(n9153), .ZN(n9449) );
  OR2_X1 U11879 ( .A1(n9580), .A2(n11259), .ZN(n9448) );
  MUX2_X1 U11880 ( .A(n13953), .B(n14121), .S(n6472), .Z(n9451) );
  MUX2_X1 U11881 ( .A(n13953), .B(n14121), .S(n9585), .Z(n9450) );
  INV_X1 U11882 ( .A(n9451), .ZN(n9452) );
  NAND2_X1 U11883 ( .A1(n9574), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9460) );
  INV_X1 U11884 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9453) );
  OR2_X1 U11885 ( .A1(n9579), .A2(n9453), .ZN(n9459) );
  OAI21_X1 U11886 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n9455), .A(n9454), .ZN(
        n13692) );
  OR2_X1 U11887 ( .A1(n9547), .A2(n13692), .ZN(n9458) );
  INV_X1 U11888 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9456) );
  OR2_X1 U11889 ( .A1(n9569), .A2(n9456), .ZN(n9457) );
  OR2_X1 U11890 ( .A1(n9461), .A2(n9678), .ZN(n9462) );
  XNOR2_X1 U11891 ( .A(n9462), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14190) );
  MUX2_X1 U11892 ( .A(n13622), .B(n13963), .S(n9585), .Z(n9463) );
  INV_X1 U11893 ( .A(n9463), .ZN(n9466) );
  MUX2_X1 U11894 ( .A(n13963), .B(n13622), .S(n9585), .Z(n9464) );
  AOI21_X1 U11895 ( .B1(n9467), .B2(n9466), .A(n9464), .ZN(n9465) );
  INV_X1 U11896 ( .A(n9465), .ZN(n9468) );
  NAND2_X1 U11897 ( .A1(n9574), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9476) );
  INV_X1 U11898 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9469) );
  OR2_X1 U11899 ( .A1(n9579), .A2(n9469), .ZN(n9475) );
  OAI21_X1 U11900 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n9471), .A(n9470), .ZN(
        n13943) );
  OR2_X1 U11901 ( .A1(n9547), .A2(n13943), .ZN(n9474) );
  INV_X1 U11902 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9472) );
  OR2_X1 U11903 ( .A1(n9569), .A2(n9472), .ZN(n9473) );
  NAND4_X1 U11904 ( .A1(n9476), .A2(n9475), .A3(n9474), .A4(n9473), .ZN(n13954) );
  NAND2_X1 U11905 ( .A1(n11529), .A2(n9153), .ZN(n9478) );
  INV_X1 U11906 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11532) );
  OR2_X1 U11907 ( .A1(n9580), .A2(n11532), .ZN(n9477) );
  MUX2_X1 U11908 ( .A(n13954), .B(n14108), .S(n6472), .Z(n9479) );
  NAND2_X1 U11909 ( .A1(n9480), .A2(n9479), .ZN(n9482) );
  MUX2_X1 U11910 ( .A(n13954), .B(n14108), .S(n9585), .Z(n9481) );
  NAND2_X1 U11911 ( .A1(n9482), .A2(n9481), .ZN(n9483) );
  NAND2_X1 U11912 ( .A1(n9148), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9491) );
  INV_X1 U11913 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n13928) );
  OR2_X1 U11914 ( .A1(n9567), .A2(n13928), .ZN(n9490) );
  OAI21_X1 U11915 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n9486), .A(n9485), .ZN(
        n13927) );
  OR2_X1 U11916 ( .A1(n9547), .A2(n13927), .ZN(n9489) );
  INV_X1 U11917 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9487) );
  OR2_X1 U11918 ( .A1(n9569), .A2(n9487), .ZN(n9488) );
  NAND4_X1 U11919 ( .A1(n9491), .A2(n9490), .A3(n9489), .A4(n9488), .ZN(n13741) );
  NAND2_X1 U11920 ( .A1(n11775), .A2(n9153), .ZN(n9493) );
  OR2_X1 U11921 ( .A1(n9580), .A2(n7163), .ZN(n9492) );
  MUX2_X1 U11922 ( .A(n13741), .B(n14102), .S(n9585), .Z(n9495) );
  MUX2_X1 U11923 ( .A(n13741), .B(n14102), .S(n6472), .Z(n9494) );
  NAND2_X1 U11924 ( .A1(n9574), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9502) );
  INV_X1 U11925 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9496) );
  OR2_X1 U11926 ( .A1(n9579), .A2(n9496), .ZN(n9501) );
  OAI21_X1 U11927 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n9497), .A(n9515), .ZN(
        n13904) );
  OR2_X1 U11928 ( .A1(n9547), .A2(n13904), .ZN(n9500) );
  INV_X1 U11929 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9498) );
  OR2_X1 U11930 ( .A1(n9569), .A2(n9498), .ZN(n9499) );
  NAND4_X1 U11931 ( .A1(n9502), .A2(n9501), .A3(n9500), .A4(n9499), .ZN(n13920) );
  NAND2_X1 U11932 ( .A1(n11858), .A2(n9153), .ZN(n9504) );
  OR2_X1 U11933 ( .A1(n9580), .A2(n11859), .ZN(n9503) );
  MUX2_X1 U11934 ( .A(n13920), .B(n14095), .S(n6472), .Z(n9508) );
  MUX2_X1 U11935 ( .A(n13920), .B(n14095), .S(n9585), .Z(n9505) );
  NAND2_X1 U11936 ( .A1(n9506), .A2(n9505), .ZN(n9512) );
  INV_X1 U11937 ( .A(n9507), .ZN(n9510) );
  INV_X1 U11938 ( .A(n9508), .ZN(n9509) );
  NAND2_X1 U11939 ( .A1(n9510), .A2(n9509), .ZN(n9511) );
  NAND2_X1 U11940 ( .A1(n9148), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9520) );
  INV_X1 U11941 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9513) );
  OR2_X1 U11942 ( .A1(n9569), .A2(n9513), .ZN(n9519) );
  INV_X1 U11943 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9514) );
  NAND2_X1 U11944 ( .A1(n9515), .A2(n9514), .ZN(n9516) );
  NAND2_X1 U11945 ( .A1(n9528), .A2(n9516), .ZN(n13889) );
  OR2_X1 U11946 ( .A1(n9547), .A2(n13889), .ZN(n9518) );
  INV_X1 U11947 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n13890) );
  OR2_X1 U11948 ( .A1(n9567), .A2(n13890), .ZN(n9517) );
  NAND4_X1 U11949 ( .A1(n9520), .A2(n9519), .A3(n9518), .A4(n9517), .ZN(n13871) );
  NAND2_X1 U11950 ( .A1(n13592), .A2(n9153), .ZN(n9522) );
  OR2_X1 U11951 ( .A1(n9580), .A2(n14186), .ZN(n9521) );
  MUX2_X1 U11952 ( .A(n13871), .B(n14089), .S(n9585), .Z(n9524) );
  MUX2_X1 U11953 ( .A(n13871), .B(n14089), .S(n6472), .Z(n9523) );
  INV_X1 U11954 ( .A(n9524), .ZN(n9525) );
  NAND2_X1 U11955 ( .A1(n9574), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9534) );
  INV_X1 U11956 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9526) );
  OR2_X1 U11957 ( .A1(n9579), .A2(n9526), .ZN(n9533) );
  INV_X1 U11958 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9527) );
  NAND2_X1 U11959 ( .A1(n9528), .A2(n9527), .ZN(n9529) );
  NAND2_X1 U11960 ( .A1(n9546), .A2(n9529), .ZN(n13873) );
  OR2_X1 U11961 ( .A1(n9547), .A2(n13873), .ZN(n9532) );
  INV_X1 U11962 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9530) );
  OR2_X1 U11963 ( .A1(n9569), .A2(n9530), .ZN(n9531) );
  NAND4_X1 U11964 ( .A1(n9534), .A2(n9533), .A3(n9532), .A4(n9531), .ZN(n13740) );
  NAND2_X1 U11965 ( .A1(n13589), .A2(n9153), .ZN(n9536) );
  OR2_X1 U11966 ( .A1(n9580), .A2(n14184), .ZN(n9535) );
  MUX2_X1 U11967 ( .A(n13740), .B(n14084), .S(n6472), .Z(n9540) );
  MUX2_X1 U11968 ( .A(n13740), .B(n14084), .S(n9585), .Z(n9537) );
  NAND2_X1 U11969 ( .A1(n9538), .A2(n9537), .ZN(n9544) );
  INV_X1 U11970 ( .A(n9539), .ZN(n9542) );
  INV_X1 U11971 ( .A(n9540), .ZN(n9541) );
  NAND2_X1 U11972 ( .A1(n9542), .A2(n9541), .ZN(n9543) );
  NAND2_X1 U11973 ( .A1(n9148), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9551) );
  INV_X1 U11974 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9545) );
  OR2_X1 U11975 ( .A1(n9569), .A2(n9545), .ZN(n9550) );
  XNOR2_X1 U11976 ( .A(n9546), .B(n12152), .ZN(n12155) );
  OR2_X1 U11977 ( .A1(n9547), .A2(n12155), .ZN(n9549) );
  INV_X1 U11978 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n11909) );
  OR2_X1 U11979 ( .A1(n9567), .A2(n11909), .ZN(n9548) );
  NAND4_X1 U11980 ( .A1(n9551), .A2(n9550), .A3(n9549), .A4(n9548), .ZN(n13872) );
  NAND2_X1 U11981 ( .A1(n12032), .A2(n9153), .ZN(n9553) );
  OR2_X1 U11982 ( .A1(n9580), .A2(n12033), .ZN(n9552) );
  NAND2_X2 U11983 ( .A1(n9553), .A2(n9552), .ZN(n14079) );
  MUX2_X1 U11984 ( .A(n13872), .B(n14079), .S(n9585), .Z(n9557) );
  NAND2_X1 U11985 ( .A1(n9556), .A2(n9557), .ZN(n9555) );
  MUX2_X1 U11986 ( .A(n14079), .B(n13872), .S(n9585), .Z(n9554) );
  INV_X1 U11987 ( .A(n9556), .ZN(n9559) );
  INV_X1 U11988 ( .A(n9557), .ZN(n9558) );
  MUX2_X1 U11989 ( .A(n13739), .B(n14071), .S(n9585), .Z(n9562) );
  NAND2_X1 U11990 ( .A1(n9563), .A2(n9153), .ZN(n9565) );
  INV_X1 U11991 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14175) );
  OR2_X1 U11992 ( .A1(n9580), .A2(n14175), .ZN(n9564) );
  INV_X1 U11993 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9566) );
  OR2_X1 U11994 ( .A1(n9579), .A2(n9566), .ZN(n9572) );
  INV_X1 U11995 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n13833) );
  OR2_X1 U11996 ( .A1(n9567), .A2(n13833), .ZN(n9571) );
  INV_X1 U11997 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9568) );
  OR2_X1 U11998 ( .A1(n9569), .A2(n9568), .ZN(n9570) );
  AND3_X1 U11999 ( .A1(n9572), .A2(n9571), .A3(n9570), .ZN(n9593) );
  INV_X1 U12000 ( .A(n9593), .ZN(n13836) );
  XNOR2_X1 U12001 ( .A(n13838), .B(n13836), .ZN(n9634) );
  INV_X1 U12002 ( .A(n10016), .ZN(n9956) );
  OR2_X1 U12003 ( .A1(n9956), .A2(n11165), .ZN(n10494) );
  NAND2_X1 U12004 ( .A1(n10238), .A2(n14189), .ZN(n10216) );
  OAI21_X1 U12005 ( .B1(n10239), .B2(n14189), .A(n10216), .ZN(n9573) );
  AND2_X1 U12006 ( .A1(n10494), .A2(n9573), .ZN(n9637) );
  NAND2_X1 U12007 ( .A1(n9634), .A2(n9637), .ZN(n9628) );
  INV_X1 U12008 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9578) );
  NAND2_X1 U12009 ( .A1(n9574), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9577) );
  NAND2_X1 U12010 ( .A1(n9575), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9576) );
  OAI211_X1 U12011 ( .C1(n9579), .C2(n9578), .A(n9577), .B(n9576), .ZN(n13857)
         );
  OAI21_X1 U12012 ( .B1(n13836), .B2(n11168), .A(n13857), .ZN(n9583) );
  NAND2_X1 U12013 ( .A1(n12159), .A2(n9153), .ZN(n9582) );
  INV_X1 U12014 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14181) );
  OR2_X1 U12015 ( .A1(n9580), .A2(n14181), .ZN(n9581) );
  MUX2_X1 U12016 ( .A(n9583), .B(n14068), .S(n9585), .Z(n9596) );
  INV_X1 U12017 ( .A(n9596), .ZN(n9592) );
  NAND2_X1 U12018 ( .A1(n13842), .A2(n6472), .ZN(n9590) );
  NAND2_X1 U12019 ( .A1(n13836), .A2(n9585), .ZN(n9586) );
  OAI21_X1 U12020 ( .B1(n10238), .B2(n9587), .A(n9586), .ZN(n9588) );
  NAND2_X1 U12021 ( .A1(n9588), .A2(n13857), .ZN(n9589) );
  NAND2_X1 U12022 ( .A1(n9590), .A2(n9589), .ZN(n9595) );
  INV_X1 U12023 ( .A(n9595), .ZN(n9591) );
  AND2_X1 U12024 ( .A1(n9592), .A2(n9591), .ZN(n9625) );
  MUX2_X1 U12025 ( .A(n14065), .B(n9593), .S(n9143), .Z(n9594) );
  OAI21_X1 U12026 ( .B1(n13838), .B2(n13836), .A(n9594), .ZN(n9635) );
  INV_X1 U12027 ( .A(n10238), .ZN(n11261) );
  AND2_X1 U12028 ( .A1(n10239), .A2(n11261), .ZN(n9954) );
  NOR2_X1 U12029 ( .A1(n9637), .A2(n9954), .ZN(n9632) );
  NAND2_X1 U12030 ( .A1(n9635), .A2(n9632), .ZN(n9630) );
  AND2_X1 U12031 ( .A1(n9596), .A2(n9595), .ZN(n9626) );
  NOR2_X1 U12032 ( .A1(n9630), .A2(n9626), .ZN(n9597) );
  INV_X1 U12033 ( .A(n9634), .ZN(n9621) );
  XNOR2_X1 U12034 ( .A(n13842), .B(n13857), .ZN(n9619) );
  INV_X1 U12035 ( .A(n13872), .ZN(n13848) );
  NAND2_X1 U12036 ( .A1(n14079), .A2(n13848), .ZN(n13845) );
  OR2_X1 U12037 ( .A1(n14079), .A2(n13848), .ZN(n9599) );
  NAND2_X1 U12038 ( .A1(n14084), .A2(n13721), .ZN(n11889) );
  OR2_X1 U12039 ( .A1(n14084), .A2(n13721), .ZN(n9600) );
  NAND2_X1 U12040 ( .A1(n11889), .A2(n9600), .ZN(n11905) );
  XOR2_X1 U12041 ( .A(n13920), .B(n14095), .Z(n13910) );
  INV_X1 U12042 ( .A(n13871), .ZN(n9601) );
  NAND2_X1 U12043 ( .A1(n14089), .A2(n9601), .ZN(n11888) );
  OR2_X1 U12044 ( .A1(n14089), .A2(n9601), .ZN(n9602) );
  XNOR2_X1 U12045 ( .A(n14102), .B(n13741), .ZN(n13918) );
  INV_X1 U12046 ( .A(n13622), .ZN(n13742) );
  XOR2_X1 U12047 ( .A(n13742), .B(n13963), .Z(n13951) );
  INV_X1 U12048 ( .A(n13953), .ZN(n13694) );
  XNOR2_X1 U12049 ( .A(n14121), .B(n13694), .ZN(n13975) );
  INV_X1 U12050 ( .A(n13998), .ZN(n13623) );
  XNOR2_X1 U12051 ( .A(n14130), .B(n13623), .ZN(n13982) );
  INV_X1 U12052 ( .A(n11898), .ZN(n9603) );
  XNOR2_X1 U12053 ( .A(n13646), .B(n12062), .ZN(n11740) );
  XNOR2_X1 U12054 ( .A(n11503), .B(n14421), .ZN(n11314) );
  XNOR2_X1 U12055 ( .A(n11466), .B(n13748), .ZN(n10922) );
  INV_X1 U12056 ( .A(n10674), .ZN(n14529) );
  NAND2_X1 U12057 ( .A1(n14529), .A2(n14543), .ZN(n10461) );
  NAND2_X1 U12058 ( .A1(n10674), .A2(n13753), .ZN(n10462) );
  NAND2_X1 U12059 ( .A1(n10461), .A2(n10462), .ZN(n10237) );
  NAND2_X1 U12060 ( .A1(n7406), .A2(n10490), .ZN(n10234) );
  NAND2_X1 U12061 ( .A1(n10231), .A2(n9606), .ZN(n14584) );
  NOR2_X1 U12062 ( .A1(n10219), .A2(n14584), .ZN(n9607) );
  NAND4_X1 U12063 ( .A1(n10237), .A2(n10233), .A3(n9607), .A4(n10226), .ZN(
        n9608) );
  NOR2_X1 U12064 ( .A1(n10689), .A2(n9608), .ZN(n9609) );
  XNOR2_X1 U12065 ( .A(n11021), .B(n13750), .ZN(n10942) );
  XNOR2_X1 U12066 ( .A(n14607), .B(n13751), .ZN(n10902) );
  NAND4_X1 U12067 ( .A1(n10922), .A2(n9609), .A3(n10942), .A4(n10902), .ZN(
        n9611) );
  XNOR2_X1 U12068 ( .A(n14431), .B(n11312), .ZN(n11309) );
  INV_X1 U12069 ( .A(n13749), .ZN(n10998) );
  XNOR2_X1 U12070 ( .A(n11200), .B(n10998), .ZN(n10955) );
  OR2_X1 U12071 ( .A1(n11605), .A2(n14420), .ZN(n11109) );
  NAND2_X1 U12072 ( .A1(n11605), .A2(n14420), .ZN(n9610) );
  NAND2_X1 U12073 ( .A1(n11109), .A2(n9610), .ZN(n10924) );
  OR4_X1 U12074 ( .A1(n9611), .A2(n11309), .A3(n10955), .A4(n10924), .ZN(n9612) );
  NOR2_X1 U12075 ( .A1(n11314), .A2(n9612), .ZN(n9613) );
  XNOR2_X1 U12076 ( .A(n11671), .B(n13744), .ZN(n11664) );
  NAND4_X1 U12077 ( .A1(n11736), .A2(n9613), .A3(n11711), .A4(n11664), .ZN(
        n9614) );
  OR4_X1 U12078 ( .A1(n7168), .A2(n14028), .A3(n11740), .A4(n9614), .ZN(n9615)
         );
  INV_X1 U12079 ( .A(n14015), .ZN(n14011) );
  NOR4_X1 U12080 ( .A1(n13975), .A2(n13982), .A3(n9615), .A4(n14011), .ZN(
        n9616) );
  XNOR2_X1 U12081 ( .A(n14108), .B(n13954), .ZN(n13935) );
  NAND4_X1 U12082 ( .A1(n13918), .A2(n13951), .A3(n9616), .A4(n13935), .ZN(
        n9617) );
  NOR4_X1 U12083 ( .A1(n11905), .A2(n13910), .A3(n13883), .A4(n9617), .ZN(
        n9618) );
  XNOR2_X1 U12084 ( .A(n14071), .B(n13739), .ZN(n13851) );
  NAND4_X1 U12085 ( .A1(n9619), .A2(n11906), .A3(n9618), .A4(n13851), .ZN(
        n9620) );
  NOR2_X1 U12086 ( .A1(n9621), .A2(n9620), .ZN(n9622) );
  XOR2_X1 U12087 ( .A(n11165), .B(n9622), .Z(n9624) );
  INV_X1 U12088 ( .A(n9954), .ZN(n9623) );
  NOR2_X1 U12089 ( .A1(n9624), .A2(n9623), .ZN(n9642) );
  INV_X1 U12090 ( .A(n9625), .ZN(n9629) );
  INV_X1 U12091 ( .A(n9626), .ZN(n9627) );
  OAI22_X1 U12092 ( .A1(n9630), .A2(n9629), .B1(n9628), .B2(n9627), .ZN(n9631)
         );
  INV_X1 U12093 ( .A(n9632), .ZN(n9633) );
  NOR2_X1 U12094 ( .A1(n9634), .A2(n9633), .ZN(n9636) );
  MUX2_X1 U12095 ( .A(n9637), .B(n9636), .S(n9635), .Z(n9638) );
  NAND3_X1 U12096 ( .A1(n9645), .A2(n9644), .A3(n9643), .ZN(n9653) );
  NAND2_X1 U12097 ( .A1(n9648), .A2(n9647), .ZN(n9654) );
  NAND2_X1 U12098 ( .A1(n9654), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9650) );
  INV_X1 U12099 ( .A(n10322), .ZN(n9651) );
  NAND2_X1 U12100 ( .A1(n9651), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11530) );
  INV_X1 U12101 ( .A(n11530), .ZN(n9652) );
  NAND2_X1 U12102 ( .A1(n9653), .A2(n9652), .ZN(n9670) );
  OAI21_X1 U12103 ( .B1(n9402), .B2(n9657), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9658) );
  MUX2_X1 U12104 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9658), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9660) );
  NAND2_X1 U12105 ( .A1(n9660), .A2(n9659), .ZN(n11860) );
  NAND2_X1 U12106 ( .A1(n9659), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9661) );
  MUX2_X1 U12107 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9661), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n9662) );
  INV_X1 U12108 ( .A(n10216), .ZN(n9967) );
  NAND2_X1 U12109 ( .A1(n11168), .A2(n11165), .ZN(n9664) );
  AND2_X1 U12110 ( .A1(n9967), .A2(n9664), .ZN(n9972) );
  NOR4_X1 U12111 ( .A1(n10475), .A2(n9972), .A3(n14542), .A4(n9666), .ZN(n9668) );
  OAI21_X1 U12112 ( .B1(n11530), .B2(n14189), .A(P1_B_REG_SCAN_IN), .ZN(n9667)
         );
  NAND2_X1 U12113 ( .A1(n9670), .A2(n9669), .ZN(P1_U3242) );
  INV_X1 U12114 ( .A(n9731), .ZN(n9671) );
  INV_X1 U12115 ( .A(n9672), .ZN(n9673) );
  AND2_X1 U12116 ( .A1(n6478), .A2(P1_U3086), .ZN(n10012) );
  INV_X2 U12117 ( .A(n10012), .ZN(n14180) );
  NOR2_X1 U12118 ( .A1(n9678), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14178) );
  INV_X2 U12119 ( .A(n14178), .ZN(n14183) );
  OAI222_X1 U12120 ( .A1(n14180), .A2(n7508), .B1(n14183), .B2(n9712), .C1(
        P1_U3086), .C2(n13761), .ZN(P1_U3354) );
  INV_X1 U12121 ( .A(n13775), .ZN(n9675) );
  INV_X1 U12122 ( .A(n9129), .ZN(n9677) );
  OAI222_X1 U12123 ( .A1(P1_U3086), .A2(n9675), .B1(n14183), .B2(n9677), .C1(
        n9674), .C2(n14180), .ZN(P1_U3353) );
  INV_X1 U12124 ( .A(n9849), .ZN(n14681) );
  NOR2_X1 U12125 ( .A1(n6478), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13585) );
  INV_X2 U12126 ( .A(n13585), .ZN(n13593) );
  OAI222_X1 U12127 ( .A1(P2_U3088), .A2(n14681), .B1(n13587), .B2(n9677), .C1(
        n9676), .C2(n13593), .ZN(P2_U3325) );
  NOR2_X1 U12128 ( .A1(n9678), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13062) );
  NAND2_X1 U12129 ( .A1(n9678), .A2(P3_U3151), .ZN(n13070) );
  AOI222_X1 U12130 ( .A1(n9679), .A2(n13062), .B1(n9693), .B2(SI_2_), .C1(
        n6483), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9680) );
  INV_X1 U12131 ( .A(n9680), .ZN(P3_U3293) );
  AOI222_X1 U12132 ( .A1(n9681), .A2(n13062), .B1(SI_4_), .B2(n9693), .C1(
        n11406), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9682) );
  INV_X1 U12133 ( .A(n9682), .ZN(P3_U3291) );
  INV_X1 U12134 ( .A(n13788), .ZN(n9685) );
  INV_X1 U12135 ( .A(n9683), .ZN(n9686) );
  OAI222_X1 U12136 ( .A1(n9685), .A2(P1_U3086), .B1(n14183), .B2(n9686), .C1(
        n9684), .C2(n14180), .ZN(P1_U3352) );
  INV_X1 U12137 ( .A(n9851), .ZN(n14695) );
  OAI222_X1 U12138 ( .A1(n13593), .A2(n9687), .B1(n13587), .B2(n9686), .C1(
        P2_U3088), .C2(n14695), .ZN(P2_U3324) );
  INV_X1 U12139 ( .A(n14491), .ZN(n9689) );
  OAI222_X1 U12140 ( .A1(P1_U3086), .A2(n9689), .B1(n14183), .B2(n9691), .C1(
        n9688), .C2(n14180), .ZN(P1_U3351) );
  INV_X1 U12141 ( .A(n13210), .ZN(n9692) );
  OAI222_X1 U12142 ( .A1(P2_U3088), .A2(n9692), .B1(n13587), .B2(n9691), .C1(
        n9690), .C2(n13593), .ZN(P2_U3323) );
  INV_X2 U12143 ( .A(n13062), .ZN(n13067) );
  INV_X2 U12144 ( .A(n9693), .ZN(n13059) );
  OAI222_X1 U12145 ( .A1(n13067), .A2(n9695), .B1(n13059), .B2(n9694), .C1(
        P3_U3151), .C2(n10360), .ZN(P3_U3294) );
  INV_X1 U12146 ( .A(SI_10_), .ZN(n9698) );
  INV_X1 U12147 ( .A(n9696), .ZN(n9697) );
  OAI222_X1 U12148 ( .A1(P3_U3151), .A2(n14969), .B1(n13059), .B2(n9698), .C1(
        n13067), .C2(n9697), .ZN(P3_U3285) );
  INV_X1 U12149 ( .A(SI_8_), .ZN(n9699) );
  OAI222_X1 U12150 ( .A1(n13067), .A2(n9700), .B1(n13059), .B2(n9699), .C1(
        P3_U3151), .C2(n14919), .ZN(P3_U3287) );
  INV_X1 U12151 ( .A(n11411), .ZN(n14866) );
  INV_X1 U12152 ( .A(SI_5_), .ZN(n9703) );
  INV_X1 U12153 ( .A(n9701), .ZN(n9702) );
  OAI222_X1 U12154 ( .A1(P3_U3151), .A2(n14866), .B1(n13059), .B2(n9703), .C1(
        n13067), .C2(n9702), .ZN(P3_U3290) );
  INV_X1 U12155 ( .A(SI_9_), .ZN(n9705) );
  OAI222_X1 U12156 ( .A1(P3_U3151), .A2(n14938), .B1(n13059), .B2(n9705), .C1(
        n13067), .C2(n9704), .ZN(P3_U3286) );
  INV_X1 U12157 ( .A(SI_7_), .ZN(n9708) );
  INV_X1 U12158 ( .A(n9706), .ZN(n9707) );
  OAI222_X1 U12159 ( .A1(P3_U3151), .A2(n14901), .B1(n13059), .B2(n9708), .C1(
        n13067), .C2(n9707), .ZN(P3_U3288) );
  INV_X1 U12160 ( .A(SI_3_), .ZN(n9710) );
  OAI222_X1 U12161 ( .A1(P3_U3151), .A2(n10442), .B1(n13059), .B2(n9710), .C1(
        n13067), .C2(n9709), .ZN(P3_U3292) );
  INV_X1 U12162 ( .A(n9903), .ZN(n9848) );
  OAI222_X1 U12163 ( .A1(P2_U3088), .A2(n9848), .B1(n13587), .B2(n9712), .C1(
        n9711), .C2(n13593), .ZN(P2_U3326) );
  OAI222_X1 U12164 ( .A1(n11490), .A2(P3_U3151), .B1(n13067), .B2(n9713), .C1(
        n13059), .C2(n15202), .ZN(P3_U3284) );
  INV_X1 U12165 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10351) );
  OAI222_X1 U12166 ( .A1(P3_U3151), .A2(n10351), .B1(n13067), .B2(n6632), .C1(
        n9714), .C2(n13059), .ZN(P3_U3295) );
  INV_X1 U12167 ( .A(SI_6_), .ZN(n9715) );
  OAI222_X1 U12168 ( .A1(P3_U3151), .A2(n14882), .B1(n13067), .B2(n9716), .C1(
        n9715), .C2(n13059), .ZN(P3_U3289) );
  INV_X1 U12169 ( .A(n13798), .ZN(n9785) );
  INV_X1 U12170 ( .A(n9717), .ZN(n9720) );
  OAI222_X1 U12171 ( .A1(P1_U3086), .A2(n9785), .B1(n14183), .B2(n9720), .C1(
        n9718), .C2(n14180), .ZN(P1_U3350) );
  INV_X1 U12172 ( .A(n9852), .ZN(n14706) );
  OAI222_X1 U12173 ( .A1(P2_U3088), .A2(n14706), .B1(n13587), .B2(n9720), .C1(
        n9719), .C2(n13593), .ZN(P2_U3322) );
  NAND2_X1 U12174 ( .A1(n13738), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9721) );
  OAI21_X1 U12175 ( .B1(n13738), .B2(n12057), .A(n9721), .ZN(P1_U3575) );
  INV_X1 U12176 ( .A(n9722), .ZN(n9723) );
  OAI222_X1 U12177 ( .A1(n13059), .A2(n9724), .B1(n13067), .B2(n9723), .C1(
        n11545), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U12178 ( .A(n10475), .ZN(n9965) );
  NAND3_X1 U12179 ( .A1(n11857), .A2(P1_B_REG_SCAN_IN), .A3(n11860), .ZN(n9726) );
  INV_X1 U12180 ( .A(n14188), .ZN(n9725) );
  NAND2_X1 U12181 ( .A1(n9965), .A2(n9952), .ZN(n14579) );
  INV_X1 U12182 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9729) );
  NAND2_X1 U12183 ( .A1(n11857), .A2(n14188), .ZN(n9938) );
  INV_X1 U12184 ( .A(n9938), .ZN(n9728) );
  AOI22_X1 U12185 ( .A1(n14579), .A2(n9729), .B1(n9731), .B2(n9728), .ZN(
        P1_U3445) );
  INV_X1 U12186 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9732) );
  NAND2_X1 U12187 ( .A1(n11860), .A2(n14188), .ZN(n9940) );
  INV_X1 U12188 ( .A(n9940), .ZN(n9730) );
  AOI22_X1 U12189 ( .A1(n14579), .A2(n9732), .B1(n9731), .B2(n9730), .ZN(
        P1_U3446) );
  NAND2_X1 U12190 ( .A1(n10475), .A2(n11530), .ZN(n9737) );
  NAND2_X1 U12191 ( .A1(n9967), .A2(n10322), .ZN(n9734) );
  NAND2_X1 U12192 ( .A1(n9734), .A2(n9733), .ZN(n9735) );
  AND2_X1 U12193 ( .A1(n9737), .A2(n9735), .ZN(n14494) );
  INV_X1 U12194 ( .A(n14494), .ZN(n14525) );
  INV_X1 U12195 ( .A(n9735), .ZN(n9736) );
  NAND2_X1 U12196 ( .A1(n9737), .A2(n9736), .ZN(n9774) );
  INV_X1 U12197 ( .A(n9774), .ZN(n9791) );
  INV_X1 U12198 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9738) );
  INV_X1 U12199 ( .A(n9665), .ZN(n9973) );
  OAI21_X1 U12200 ( .B1(n9666), .B2(P1_REG2_REG_0__SCAN_IN), .A(n9973), .ZN(
        n13770) );
  AOI21_X1 U12201 ( .B1(n9666), .B2(n9738), .A(n13770), .ZN(n9739) );
  INV_X1 U12202 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n13769) );
  XNOR2_X1 U12203 ( .A(n9739), .B(n13769), .ZN(n9740) );
  AOI22_X1 U12204 ( .A1(n9791), .A2(n9740), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9741) );
  OAI21_X1 U12205 ( .B1(n14525), .B2(n6975), .A(n9741), .ZN(P1_U3243) );
  INV_X1 U12206 ( .A(n10035), .ZN(n10043) );
  INV_X1 U12207 ( .A(n9742), .ZN(n9745) );
  OAI222_X1 U12208 ( .A1(P2_U3088), .A2(n10043), .B1(n13587), .B2(n9745), .C1(
        n9743), .C2(n13593), .ZN(P2_U3321) );
  INV_X1 U12209 ( .A(n9797), .ZN(n9804) );
  OAI222_X1 U12210 ( .A1(P1_U3086), .A2(n9804), .B1(n14183), .B2(n9745), .C1(
        n9744), .C2(n14180), .ZN(P1_U3349) );
  NOR2_X1 U12211 ( .A1(n14494), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12212 ( .A(n9746), .ZN(n9748) );
  INV_X1 U12213 ( .A(n9805), .ZN(n9879) );
  OAI222_X1 U12214 ( .A1(n14180), .A2(n9747), .B1(n14183), .B2(n9748), .C1(
        n9879), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U12215 ( .A(n9983), .ZN(n9860) );
  OAI222_X1 U12216 ( .A1(n13593), .A2(n9749), .B1(n13587), .B2(n9748), .C1(
        P2_U3088), .C2(n9860), .ZN(P2_U3320) );
  INV_X1 U12217 ( .A(SI_13_), .ZN(n15144) );
  OAI222_X1 U12218 ( .A1(P3_U3151), .A2(n12529), .B1(n13059), .B2(n15144), 
        .C1(n13067), .C2(n9750), .ZN(P3_U3282) );
  INV_X1 U12219 ( .A(n9751), .ZN(n9754) );
  INV_X1 U12220 ( .A(n10094), .ZN(n9981) );
  OAI222_X1 U12221 ( .A1(n13593), .A2(n9752), .B1(n13587), .B2(n9754), .C1(
        P2_U3088), .C2(n9981), .ZN(P2_U3319) );
  INV_X1 U12222 ( .A(n9808), .ZN(n9864) );
  OAI222_X1 U12223 ( .A1(n9864), .A2(P1_U3086), .B1(n14183), .B2(n9754), .C1(
        n9753), .C2(n14180), .ZN(P1_U3347) );
  OAI222_X1 U12224 ( .A1(P3_U3151), .A2(n12558), .B1(n13059), .B2(n7301), .C1(
        n13067), .C2(n9755), .ZN(P3_U3281) );
  OAI222_X1 U12225 ( .A1(P2_U3088), .A2(n14722), .B1(n13587), .B2(n9758), .C1(
        n9756), .C2(n13593), .ZN(P2_U3318) );
  INV_X1 U12226 ( .A(n9909), .ZN(n9915) );
  OAI222_X1 U12227 ( .A1(P1_U3086), .A2(n9915), .B1(n14183), .B2(n9758), .C1(
        n9757), .C2(n14180), .ZN(P1_U3346) );
  AND2_X1 U12228 ( .A1(n9760), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12229 ( .A1(n9760), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12230 ( .A1(n9760), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12231 ( .A1(n9760), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12232 ( .A1(n9760), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12233 ( .A1(n9760), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12234 ( .A1(n9760), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12235 ( .A1(n9760), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12236 ( .A1(n9760), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12237 ( .A1(n9760), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12238 ( .A1(n9760), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12239 ( .A1(n9760), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12240 ( .A1(n9760), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12241 ( .A1(n9760), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12242 ( .A1(n9760), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12243 ( .A1(n9760), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12244 ( .A1(n9760), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12245 ( .A1(n9760), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12246 ( .A1(n9760), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12247 ( .A1(n9760), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12248 ( .A1(n9760), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12249 ( .A1(n9760), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12250 ( .A1(n9760), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12251 ( .A1(n9760), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12252 ( .A1(n9760), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12253 ( .A1(n9760), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12254 ( .A1(n9760), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12255 ( .A1(n9760), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12256 ( .A1(n9760), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12257 ( .A1(n9760), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  INV_X1 U12258 ( .A(n9761), .ZN(n9763) );
  INV_X1 U12259 ( .A(n10980), .ZN(n10107) );
  OAI222_X1 U12260 ( .A1(n13593), .A2(n9762), .B1(n13587), .B2(n9763), .C1(
        P2_U3088), .C2(n10107), .ZN(P2_U3317) );
  INV_X1 U12261 ( .A(n9930), .ZN(n9924) );
  OAI222_X1 U12262 ( .A1(n14180), .A2(n9764), .B1(n14183), .B2(n9763), .C1(
        n9924), .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U12263 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9765) );
  MUX2_X1 U12264 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9765), .S(n13775), .Z(
        n13779) );
  INV_X1 U12265 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9766) );
  MUX2_X1 U12266 ( .A(n9766), .B(P1_REG1_REG_1__SCAN_IN), .S(n13761), .Z(n9768) );
  AND2_X1 U12267 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9767) );
  NAND2_X1 U12268 ( .A1(n9768), .A2(n9767), .ZN(n13760) );
  OR2_X1 U12269 ( .A1(n13761), .A2(n9766), .ZN(n9769) );
  NAND2_X1 U12270 ( .A1(n13760), .A2(n9769), .ZN(n13778) );
  NAND2_X1 U12271 ( .A1(n13779), .A2(n13778), .ZN(n13785) );
  NAND2_X1 U12272 ( .A1(n13775), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n13784) );
  NAND2_X1 U12273 ( .A1(n13785), .A2(n13784), .ZN(n9772) );
  INV_X1 U12274 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9770) );
  MUX2_X1 U12275 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9770), .S(n13788), .Z(n9771) );
  NAND2_X1 U12276 ( .A1(n9772), .A2(n9771), .ZN(n14487) );
  NAND2_X1 U12277 ( .A1(n13788), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n14486) );
  MUX2_X1 U12278 ( .A(n9170), .B(P1_REG1_REG_4__SCAN_IN), .S(n14491), .Z(
        n14485) );
  AOI21_X1 U12279 ( .B1(n14487), .B2(n14486), .A(n14485), .ZN(n14484) );
  AOI21_X1 U12280 ( .B1(n14491), .B2(P1_REG1_REG_4__SCAN_IN), .A(n14484), .ZN(
        n13800) );
  INV_X1 U12281 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10470) );
  MUX2_X1 U12282 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10470), .S(n13798), .Z(
        n13801) );
  NAND2_X1 U12283 ( .A1(n13800), .A2(n13801), .ZN(n13799) );
  OAI21_X1 U12284 ( .B1(n13798), .B2(P1_REG1_REG_5__SCAN_IN), .A(n13799), .ZN(
        n9776) );
  MUX2_X1 U12285 ( .A(n9803), .B(P1_REG1_REG_6__SCAN_IN), .S(n9797), .Z(n9775)
         );
  NOR2_X1 U12286 ( .A1(n9776), .A2(n9775), .ZN(n9883) );
  INV_X1 U12287 ( .A(n9666), .ZN(n9773) );
  AOI211_X1 U12288 ( .C1(n9776), .C2(n9775), .A(n9883), .B(n14517), .ZN(n9795)
         );
  NOR2_X1 U12289 ( .A1(n9665), .A2(n9666), .ZN(n9777) );
  INV_X1 U12290 ( .A(n14483), .ZN(n14519) );
  MUX2_X1 U12291 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9778), .S(n13775), .Z(
        n13774) );
  MUX2_X1 U12292 ( .A(n14056), .B(P1_REG2_REG_1__SCAN_IN), .S(n13761), .Z(
        n13757) );
  AND2_X1 U12293 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n13766) );
  NAND2_X1 U12294 ( .A1(n13757), .A2(n13766), .ZN(n13756) );
  OR2_X1 U12295 ( .A1(n13761), .A2(n14056), .ZN(n9779) );
  NAND2_X1 U12296 ( .A1(n13756), .A2(n9779), .ZN(n13773) );
  NAND2_X1 U12297 ( .A1(n13774), .A2(n13773), .ZN(n13790) );
  NAND2_X1 U12298 ( .A1(n13775), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13789) );
  NAND2_X1 U12299 ( .A1(n13790), .A2(n13789), .ZN(n9782) );
  MUX2_X1 U12300 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9780), .S(n13788), .Z(n9781) );
  NAND2_X1 U12301 ( .A1(n9782), .A2(n9781), .ZN(n14480) );
  NAND2_X1 U12302 ( .A1(n13788), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14479) );
  NAND2_X1 U12303 ( .A1(n14480), .A2(n14479), .ZN(n9784) );
  MUX2_X1 U12304 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n14528), .S(n14491), .Z(
        n9783) );
  NAND2_X1 U12305 ( .A1(n9784), .A2(n9783), .ZN(n14482) );
  NAND2_X1 U12306 ( .A1(n14491), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n13805) );
  MUX2_X1 U12307 ( .A(n9184), .B(P1_REG2_REG_5__SCAN_IN), .S(n13798), .Z(
        n13804) );
  AOI21_X1 U12308 ( .B1(n14482), .B2(n13805), .A(n13804), .ZN(n13803) );
  NOR2_X1 U12309 ( .A1(n9785), .A2(n9184), .ZN(n9788) );
  MUX2_X1 U12310 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9786), .S(n9797), .Z(n9787)
         );
  OAI21_X1 U12311 ( .B1(n13803), .B2(n9788), .A(n9787), .ZN(n9876) );
  INV_X1 U12312 ( .A(n9876), .ZN(n9790) );
  NOR3_X1 U12313 ( .A1(n13803), .A2(n9788), .A3(n9787), .ZN(n9789) );
  NOR3_X1 U12314 ( .A1(n14519), .A2(n9790), .A3(n9789), .ZN(n9794) );
  NAND2_X1 U12315 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n13709) );
  NAND2_X1 U12316 ( .A1(n14494), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9792) );
  OAI211_X1 U12317 ( .C1(n14521), .C2(n9804), .A(n13709), .B(n9792), .ZN(n9793) );
  OR3_X1 U12318 ( .A1(n9795), .A2(n9794), .A3(n9793), .ZN(P1_U3249) );
  OAI222_X1 U12319 ( .A1(P3_U3151), .A2(n12577), .B1(n13070), .B2(n15068), 
        .C1(n13067), .C2(n9796), .ZN(P3_U3280) );
  NAND2_X1 U12320 ( .A1(n9797), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9875) );
  INV_X1 U12321 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9798) );
  MUX2_X1 U12322 ( .A(n9798), .B(P1_REG2_REG_7__SCAN_IN), .S(n9805), .Z(n9874)
         );
  AOI21_X1 U12323 ( .B1(n9876), .B2(n9875), .A(n9874), .ZN(n9889) );
  NOR2_X1 U12324 ( .A1(n9879), .A2(n9798), .ZN(n9868) );
  MUX2_X1 U12325 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n9799), .S(n9808), .Z(n9867)
         );
  OAI21_X1 U12326 ( .B1(n9889), .B2(n9868), .A(n9867), .ZN(n9870) );
  NAND2_X1 U12327 ( .A1(n9808), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9801) );
  MUX2_X1 U12328 ( .A(n11002), .B(P1_REG2_REG_9__SCAN_IN), .S(n9909), .Z(n9800) );
  AOI21_X1 U12329 ( .B1(n9870), .B2(n9801), .A(n9800), .ZN(n9921) );
  NAND3_X1 U12330 ( .A1(n9870), .A2(n9801), .A3(n9800), .ZN(n9802) );
  NAND2_X1 U12331 ( .A1(n9802), .A2(n14483), .ZN(n9817) );
  NOR2_X1 U12332 ( .A1(n9804), .A2(n9803), .ZN(n9882) );
  MUX2_X1 U12333 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9806), .S(n9805), .Z(n9881)
         );
  OAI21_X1 U12334 ( .B1(n9883), .B2(n9882), .A(n9881), .ZN(n9885) );
  OAI21_X1 U12335 ( .B1(n9806), .B2(n9879), .A(n9885), .ZN(n9862) );
  MUX2_X1 U12336 ( .A(n9807), .B(P1_REG1_REG_8__SCAN_IN), .S(n9808), .Z(n9863)
         );
  NOR2_X1 U12337 ( .A1(n9862), .A2(n9863), .ZN(n9861) );
  NOR2_X1 U12338 ( .A1(n9808), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9809) );
  MUX2_X1 U12339 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9249), .S(n9909), .Z(n9810)
         );
  OAI21_X1 U12340 ( .B1(n9861), .B2(n9809), .A(n9810), .ZN(n9908) );
  INV_X1 U12341 ( .A(n9908), .ZN(n9812) );
  NOR3_X1 U12342 ( .A1(n9861), .A2(n9810), .A3(n9809), .ZN(n9811) );
  OAI21_X1 U12343 ( .B1(n9812), .B2(n9811), .A(n14490), .ZN(n9816) );
  INV_X1 U12344 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11467) );
  NOR2_X1 U12345 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11467), .ZN(n9814) );
  NOR2_X1 U12346 ( .A1(n14521), .A2(n9915), .ZN(n9813) );
  AOI211_X1 U12347 ( .C1(n14494), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n9814), .B(
        n9813), .ZN(n9815) );
  OAI211_X1 U12348 ( .C1(n9921), .C2(n9817), .A(n9816), .B(n9815), .ZN(
        P1_U3252) );
  NAND2_X1 U12349 ( .A1(n9818), .A2(n10119), .ZN(n9820) );
  NAND2_X1 U12350 ( .A1(n9820), .A2(n9819), .ZN(n9821) );
  AND2_X1 U12351 ( .A1(n9854), .A2(n8281), .ZN(n14680) );
  AND2_X1 U12352 ( .A1(n14680), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14776) );
  OR2_X1 U12353 ( .A1(n9854), .A2(P2_U3088), .ZN(n14752) );
  AND2_X1 U12354 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10515) );
  NOR2_X1 U12355 ( .A1(n8281), .A2(P2_U3088), .ZN(n13584) );
  AND2_X1 U12356 ( .A1(n13584), .A2(n13590), .ZN(n9824) );
  NAND2_X1 U12357 ( .A1(n9854), .A2(n9824), .ZN(n14746) );
  INV_X1 U12358 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9825) );
  MUX2_X1 U12359 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9825), .S(n9849), .Z(n14688) );
  INV_X1 U12360 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9826) );
  MUX2_X1 U12361 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9826), .S(n9903), .Z(n9828)
         );
  AND2_X1 U12362 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9827) );
  NAND2_X1 U12363 ( .A1(n9828), .A2(n9827), .ZN(n9899) );
  NAND2_X1 U12364 ( .A1(n9903), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9829) );
  NAND2_X1 U12365 ( .A1(n9899), .A2(n9829), .ZN(n14689) );
  NAND2_X1 U12366 ( .A1(n14688), .A2(n14689), .ZN(n14687) );
  NAND2_X1 U12367 ( .A1(n9849), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9830) );
  NAND2_X1 U12368 ( .A1(n14687), .A2(n9830), .ZN(n14702) );
  INV_X1 U12369 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9831) );
  MUX2_X1 U12370 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9831), .S(n9851), .Z(n14701) );
  NAND2_X1 U12371 ( .A1(n14702), .A2(n14701), .ZN(n14700) );
  NAND2_X1 U12372 ( .A1(n9851), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n13212) );
  NAND2_X1 U12373 ( .A1(n14700), .A2(n13212), .ZN(n9834) );
  INV_X1 U12374 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9832) );
  MUX2_X1 U12375 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9832), .S(n13210), .Z(n9833) );
  NAND2_X1 U12376 ( .A1(n9834), .A2(n9833), .ZN(n13214) );
  NAND2_X1 U12377 ( .A1(n13210), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9835) );
  NAND2_X1 U12378 ( .A1(n13214), .A2(n9835), .ZN(n14712) );
  INV_X1 U12379 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9836) );
  MUX2_X1 U12380 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9836), .S(n9852), .Z(n14711) );
  NAND2_X1 U12381 ( .A1(n14712), .A2(n14711), .ZN(n14710) );
  NAND2_X1 U12382 ( .A1(n9852), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10037) );
  NAND2_X1 U12383 ( .A1(n14710), .A2(n10037), .ZN(n9839) );
  INV_X1 U12384 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9837) );
  MUX2_X1 U12385 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9837), .S(n10035), .Z(n9838) );
  NAND2_X1 U12386 ( .A1(n9839), .A2(n9838), .ZN(n10039) );
  NAND2_X1 U12387 ( .A1(n10035), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9844) );
  NAND2_X1 U12388 ( .A1(n10039), .A2(n9844), .ZN(n9842) );
  INV_X1 U12389 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9840) );
  MUX2_X1 U12390 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9840), .S(n9983), .Z(n9841)
         );
  NAND2_X1 U12391 ( .A1(n9842), .A2(n9841), .ZN(n9989) );
  MUX2_X1 U12392 ( .A(n9840), .B(P2_REG1_REG_7__SCAN_IN), .S(n9983), .Z(n9843)
         );
  NAND3_X1 U12393 ( .A1(n10039), .A2(n9844), .A3(n9843), .ZN(n9845) );
  AND3_X1 U12394 ( .A1(n14783), .A2(n9989), .A3(n9845), .ZN(n9846) );
  AOI211_X1 U12395 ( .C1(n14775), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n10515), .B(
        n9846), .ZN(n9859) );
  MUX2_X1 U12396 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n9847), .S(n9903), .Z(n9895)
         );
  NAND3_X1 U12397 ( .A1(n9895), .A2(P2_REG2_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n9896) );
  OAI21_X1 U12398 ( .B1(n9847), .B2(n9848), .A(n9896), .ZN(n14686) );
  MUX2_X1 U12399 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n13462), .S(n9849), .Z(
        n14685) );
  NAND2_X1 U12400 ( .A1(n14686), .A2(n14685), .ZN(n14684) );
  OAI21_X1 U12401 ( .B1(n13462), .B2(n14681), .A(n14684), .ZN(n14699) );
  MUX2_X1 U12402 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n9850), .S(n9851), .Z(n14698) );
  NAND2_X1 U12403 ( .A1(n14699), .A2(n14698), .ZN(n14697) );
  NAND2_X1 U12404 ( .A1(n9851), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n13205) );
  MUX2_X1 U12405 ( .A(n10613), .B(P2_REG2_REG_4__SCAN_IN), .S(n13210), .Z(
        n13204) );
  AOI21_X1 U12406 ( .B1(n14697), .B2(n13205), .A(n13204), .ZN(n13207) );
  MUX2_X1 U12407 ( .A(n10557), .B(P2_REG2_REG_5__SCAN_IN), .S(n9852), .Z(
        n14715) );
  NOR2_X1 U12408 ( .A1(n14716), .A2(n14715), .ZN(n14714) );
  AOI21_X1 U12409 ( .B1(n9852), .B2(P2_REG2_REG_5__SCAN_IN), .A(n14714), .ZN(
        n10032) );
  MUX2_X1 U12410 ( .A(n10580), .B(P2_REG2_REG_6__SCAN_IN), .S(n10035), .Z(
        n10031) );
  NOR2_X1 U12411 ( .A1(n10032), .A2(n10031), .ZN(n10030) );
  NOR2_X1 U12412 ( .A1(n10043), .A2(n10580), .ZN(n9856) );
  MUX2_X1 U12413 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10777), .S(n9983), .Z(n9855) );
  AND2_X1 U12414 ( .A1(n13584), .A2(n11991), .ZN(n9853) );
  AND2_X1 U12415 ( .A1(n9854), .A2(n9853), .ZN(n14778) );
  OR3_X1 U12416 ( .A1(n10030), .A2(n9856), .A3(n9855), .ZN(n9857) );
  NAND3_X1 U12417 ( .A1(n9978), .A2(n14778), .A3(n9857), .ZN(n9858) );
  OAI211_X1 U12418 ( .C1(n14707), .C2(n9860), .A(n9859), .B(n9858), .ZN(
        P2_U3221) );
  AOI21_X1 U12419 ( .B1(n9863), .B2(n9862), .A(n9861), .ZN(n9873) );
  AND2_X1 U12420 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9866) );
  NOR2_X1 U12421 ( .A1(n14521), .A2(n9864), .ZN(n9865) );
  AOI211_X1 U12422 ( .C1(n14494), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9866), .B(
        n9865), .ZN(n9872) );
  OR3_X1 U12423 ( .A1(n9889), .A2(n9868), .A3(n9867), .ZN(n9869) );
  NAND3_X1 U12424 ( .A1(n14483), .A2(n9870), .A3(n9869), .ZN(n9871) );
  OAI211_X1 U12425 ( .C1(n9873), .C2(n14517), .A(n9872), .B(n9871), .ZN(
        P1_U3251) );
  NAND3_X1 U12426 ( .A1(n9876), .A2(n9875), .A3(n9874), .ZN(n9877) );
  NAND2_X1 U12427 ( .A1(n14483), .A2(n9877), .ZN(n9888) );
  NOR2_X1 U12428 ( .A1(n9878), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11027) );
  NOR2_X1 U12429 ( .A1(n14521), .A2(n9879), .ZN(n9880) );
  AOI211_X1 U12430 ( .C1(n14494), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n11027), .B(
        n9880), .ZN(n9887) );
  OR3_X1 U12431 ( .A1(n9883), .A2(n9882), .A3(n9881), .ZN(n9884) );
  NAND3_X1 U12432 ( .A1(n9885), .A2(n14490), .A3(n9884), .ZN(n9886) );
  OAI211_X1 U12433 ( .C1(n9889), .C2(n9888), .A(n9887), .B(n9886), .ZN(
        P1_U3250) );
  INV_X1 U12434 ( .A(n9890), .ZN(n9893) );
  INV_X1 U12435 ( .A(n13228), .ZN(n10974) );
  OAI222_X1 U12436 ( .A1(n13593), .A2(n9891), .B1(n13587), .B2(n9893), .C1(
        P2_U3088), .C2(n10974), .ZN(P2_U3316) );
  INV_X1 U12437 ( .A(n10001), .ZN(n9994) );
  OAI222_X1 U12438 ( .A1(n9994), .A2(P1_U3086), .B1(n14183), .B2(n9893), .C1(
        n9892), .C2(n14180), .ZN(P1_U3344) );
  NOR2_X1 U12439 ( .A1(n14713), .A2(n9894), .ZN(n14674) );
  AOI22_X1 U12440 ( .A1(n14674), .A2(P2_IR_REG_0__SCAN_IN), .B1(n14778), .B2(
        n9895), .ZN(n9907) );
  INV_X1 U12441 ( .A(n9896), .ZN(n9906) );
  INV_X1 U12442 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n14845) );
  MUX2_X1 U12443 ( .A(n9826), .B(P2_REG1_REG_1__SCAN_IN), .S(n9903), .Z(n9897)
         );
  OAI21_X1 U12444 ( .B1(n14845), .B2(n9898), .A(n9897), .ZN(n9900) );
  NAND2_X1 U12445 ( .A1(n9900), .A2(n9899), .ZN(n9901) );
  OAI22_X1 U12446 ( .A1(n14746), .A2(n9901), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10590), .ZN(n9902) );
  AOI21_X1 U12447 ( .B1(n14775), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n9902), .ZN(
        n9905) );
  NAND2_X1 U12448 ( .A1(n14776), .A2(n9903), .ZN(n9904) );
  OAI211_X1 U12449 ( .C1(n9907), .C2(n9906), .A(n9905), .B(n9904), .ZN(
        P2_U3215) );
  AND2_X1 U12450 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11612) );
  MUX2_X1 U12451 ( .A(n9265), .B(P1_REG1_REG_10__SCAN_IN), .S(n9930), .Z(n9911) );
  OAI21_X1 U12452 ( .B1(n9909), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9908), .ZN(
        n9910) );
  NOR2_X1 U12453 ( .A1(n9910), .A2(n9911), .ZN(n9929) );
  AOI211_X1 U12454 ( .C1(n9911), .C2(n9910), .A(n14517), .B(n9929), .ZN(n9912)
         );
  INV_X1 U12455 ( .A(n9912), .ZN(n9913) );
  OAI21_X1 U12456 ( .B1(n14219), .B2(n14525), .A(n9913), .ZN(n9914) );
  NOR2_X1 U12457 ( .A1(n11612), .A2(n9914), .ZN(n9923) );
  NOR2_X1 U12458 ( .A1(n9915), .A2(n11002), .ZN(n9919) );
  INV_X1 U12459 ( .A(n9919), .ZN(n9917) );
  INV_X1 U12460 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10928) );
  MUX2_X1 U12461 ( .A(n10928), .B(P1_REG2_REG_10__SCAN_IN), .S(n9930), .Z(
        n9916) );
  NAND2_X1 U12462 ( .A1(n9917), .A2(n9916), .ZN(n9920) );
  MUX2_X1 U12463 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10928), .S(n9930), .Z(
        n9918) );
  OAI21_X1 U12464 ( .B1(n9921), .B2(n9919), .A(n9918), .ZN(n9927) );
  OAI211_X1 U12465 ( .C1(n9921), .C2(n9920), .A(n9927), .B(n14483), .ZN(n9922)
         );
  OAI211_X1 U12466 ( .C1(n14521), .C2(n9924), .A(n9923), .B(n9922), .ZN(
        P1_U3253) );
  NAND2_X1 U12467 ( .A1(n9930), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9926) );
  MUX2_X1 U12468 ( .A(n11121), .B(P1_REG2_REG_11__SCAN_IN), .S(n10001), .Z(
        n9925) );
  AOI21_X1 U12469 ( .B1(n9927), .B2(n9926), .A(n9925), .ZN(n10000) );
  NAND3_X1 U12470 ( .A1(n9927), .A2(n9926), .A3(n9925), .ZN(n9928) );
  NAND2_X1 U12471 ( .A1(n9928), .A2(n14483), .ZN(n9937) );
  MUX2_X1 U12472 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9276), .S(n10001), .Z(
        n9932) );
  AOI21_X1 U12473 ( .B1(n9930), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9929), .ZN(
        n9931) );
  NAND2_X1 U12474 ( .A1(n9931), .A2(n9932), .ZN(n9998) );
  OAI21_X1 U12475 ( .B1(n9932), .B2(n9931), .A(n9998), .ZN(n9933) );
  NAND2_X1 U12476 ( .A1(n9933), .A2(n14490), .ZN(n9936) );
  INV_X1 U12477 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14194) );
  NAND2_X1 U12478 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14433)
         );
  OAI21_X1 U12479 ( .B1(n14525), .B2(n14194), .A(n14433), .ZN(n9934) );
  AOI21_X1 U12480 ( .B1(n10001), .B2(n14492), .A(n9934), .ZN(n9935) );
  OAI211_X1 U12481 ( .C1(n10000), .C2(n9937), .A(n9936), .B(n9935), .ZN(
        P1_U3254) );
  OR2_X1 U12482 ( .A1(n9952), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9939) );
  OR2_X1 U12483 ( .A1(n9952), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9941) );
  AND2_X1 U12484 ( .A1(n9941), .A2(n9940), .ZN(n10213) );
  NAND2_X1 U12485 ( .A1(n13858), .A2(n10213), .ZN(n9963) );
  NOR4_X1 U12486 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9950) );
  NOR4_X1 U12487 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9949) );
  OR4_X1 U12488 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9947) );
  NOR4_X1 U12489 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9945) );
  NOR4_X1 U12490 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9944) );
  NOR4_X1 U12491 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9943) );
  NOR4_X1 U12492 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9942) );
  NAND4_X1 U12493 ( .A1(n9945), .A2(n9944), .A3(n9943), .A4(n9942), .ZN(n9946)
         );
  NOR4_X1 U12494 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9947), .A4(n9946), .ZN(n9948) );
  AND3_X1 U12495 ( .A1(n9950), .A2(n9949), .A3(n9948), .ZN(n9951) );
  NOR2_X1 U12496 ( .A1(n9952), .A2(n9951), .ZN(n9964) );
  INV_X1 U12497 ( .A(n14189), .ZN(n9953) );
  NAND2_X1 U12498 ( .A1(n14636), .A2(n11261), .ZN(n10474) );
  OAI21_X1 U12499 ( .B1(n9963), .B2(n9964), .A(n10474), .ZN(n10324) );
  OR2_X1 U12500 ( .A1(n10238), .A2(n14189), .ZN(n10229) );
  NAND2_X1 U12501 ( .A1(n14564), .A2(n13826), .ZN(n9955) );
  NAND2_X1 U12502 ( .A1(n9954), .A2(n9953), .ZN(n10486) );
  INV_X1 U12503 ( .A(n14432), .ZN(n13737) );
  NAND2_X1 U12504 ( .A1(n10630), .A2(n14565), .ZN(n9958) );
  INV_X1 U12505 ( .A(n10323), .ZN(n9960) );
  OR2_X1 U12506 ( .A1(n14047), .A2(n12106), .ZN(n9961) );
  NAND2_X1 U12507 ( .A1(n9962), .A2(n10021), .ZN(n10023) );
  OAI21_X1 U12508 ( .B1(n9962), .B2(n10021), .A(n10023), .ZN(n13767) );
  INV_X1 U12509 ( .A(n9963), .ZN(n9971) );
  INV_X1 U12510 ( .A(n9964), .ZN(n9966) );
  AND2_X1 U12511 ( .A1(n9966), .A2(n9965), .ZN(n10214) );
  INV_X1 U12512 ( .A(n10214), .ZN(n9969) );
  OR2_X1 U12513 ( .A1(n14606), .A2(n9967), .ZN(n9968) );
  NOR2_X1 U12514 ( .A1(n9969), .A2(n9968), .ZN(n9970) );
  NAND2_X1 U12515 ( .A1(n13862), .A2(n13858), .ZN(n13672) );
  AND2_X1 U12516 ( .A1(n14414), .A2(n14055), .ZN(n13729) );
  AOI22_X1 U12517 ( .A1(n13767), .A2(n14412), .B1(n13729), .B2(n13755), .ZN(
        n9975) );
  NAND2_X1 U12518 ( .A1(n11472), .A2(n10321), .ZN(n12029) );
  NAND2_X1 U12519 ( .A1(n12029), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9974) );
  OAI211_X1 U12520 ( .C1(n13737), .C2(n10218), .A(n9975), .B(n9974), .ZN(
        P1_U3232) );
  NAND2_X1 U12521 ( .A1(n9983), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9977) );
  MUX2_X1 U12522 ( .A(n10788), .B(P2_REG2_REG_8__SCAN_IN), .S(n10094), .Z(
        n9976) );
  AOI21_X1 U12523 ( .B1(n9978), .B2(n9977), .A(n9976), .ZN(n10090) );
  NAND3_X1 U12524 ( .A1(n9978), .A2(n9977), .A3(n9976), .ZN(n9979) );
  NAND2_X1 U12525 ( .A1(n9979), .A2(n14778), .ZN(n9993) );
  NOR2_X1 U12526 ( .A1(n9980), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10529) );
  NOR2_X1 U12527 ( .A1(n14707), .A2(n9981), .ZN(n9982) );
  AOI211_X1 U12528 ( .C1(n14775), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n10529), .B(
        n9982), .ZN(n9992) );
  NAND2_X1 U12529 ( .A1(n9983), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9988) );
  NAND2_X1 U12530 ( .A1(n9989), .A2(n9988), .ZN(n9986) );
  INV_X1 U12531 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9984) );
  MUX2_X1 U12532 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9984), .S(n10094), .Z(n9985) );
  NAND2_X1 U12533 ( .A1(n9986), .A2(n9985), .ZN(n10096) );
  MUX2_X1 U12534 ( .A(n9984), .B(P2_REG1_REG_8__SCAN_IN), .S(n10094), .Z(n9987) );
  NAND3_X1 U12535 ( .A1(n9989), .A2(n9988), .A3(n9987), .ZN(n9990) );
  NAND3_X1 U12536 ( .A1(n14783), .A2(n10096), .A3(n9990), .ZN(n9991) );
  OAI211_X1 U12537 ( .C1(n10090), .C2(n9993), .A(n9992), .B(n9991), .ZN(
        P2_U3222) );
  NAND2_X1 U12538 ( .A1(n9994), .A2(n9276), .ZN(n9996) );
  MUX2_X1 U12539 ( .A(n9995), .B(P1_REG1_REG_12__SCAN_IN), .S(n10275), .Z(
        n9997) );
  AOI21_X1 U12540 ( .B1(n9998), .B2(n9996), .A(n9997), .ZN(n10267) );
  AND3_X1 U12541 ( .A1(n9998), .A2(n9997), .A3(n9996), .ZN(n9999) );
  OAI21_X1 U12542 ( .B1(n10267), .B2(n9999), .A(n14490), .ZN(n10009) );
  MUX2_X1 U12543 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n11320), .S(n10275), .Z(
        n10003) );
  AOI21_X1 U12544 ( .B1(n10001), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10000), 
        .ZN(n10002) );
  NAND2_X1 U12545 ( .A1(n10002), .A2(n10003), .ZN(n10274) );
  OAI21_X1 U12546 ( .B1(n10003), .B2(n10002), .A(n10274), .ZN(n10007) );
  INV_X1 U12547 ( .A(n10275), .ZN(n10268) );
  NOR2_X1 U12548 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11811), .ZN(n10004) );
  AOI21_X1 U12549 ( .B1(n14494), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n10004), 
        .ZN(n10005) );
  OAI21_X1 U12550 ( .B1(n14521), .B2(n10268), .A(n10005), .ZN(n10006) );
  AOI21_X1 U12551 ( .B1(n10007), .B2(n14483), .A(n10006), .ZN(n10008) );
  NAND2_X1 U12552 ( .A1(n10009), .A2(n10008), .ZN(P1_U3255) );
  OAI222_X1 U12553 ( .A1(P3_U3151), .A2(n12598), .B1(n13059), .B2(n15094), 
        .C1(n13067), .C2(n10010), .ZN(P3_U3279) );
  INV_X1 U12554 ( .A(n10011), .ZN(n10085) );
  AOI22_X1 U12555 ( .A1(n10275), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10012), .ZN(n10013) );
  OAI21_X1 U12556 ( .B1(n10085), .B2(n14183), .A(n10013), .ZN(P1_U3343) );
  AND2_X1 U12557 ( .A1(n11165), .A2(n14189), .ZN(n10015) );
  XNOR2_X1 U12558 ( .A(n10017), .B(n12141), .ZN(n10019) );
  OAI22_X1 U12559 ( .A1(n14563), .A2(n12105), .B1(n10220), .B2(n12106), .ZN(
        n10018) );
  NOR2_X1 U12560 ( .A1(n10019), .A2(n10018), .ZN(n10309) );
  NAND2_X1 U12561 ( .A1(n10023), .A2(n10022), .ZN(n10024) );
  NAND2_X1 U12562 ( .A1(n10024), .A2(n10025), .ZN(n10311) );
  OAI21_X1 U12563 ( .B1(n10025), .B2(n10024), .A(n10311), .ZN(n10026) );
  NAND2_X1 U12564 ( .A1(n10026), .A2(n14412), .ZN(n10029) );
  INV_X1 U12565 ( .A(n13729), .ZN(n14422) );
  OR2_X1 U12566 ( .A1(n13672), .A2(n14542), .ZN(n14419) );
  OAI22_X1 U12567 ( .A1(n14422), .A2(n7406), .B1(n14047), .B2(n14419), .ZN(
        n10027) );
  AOI21_X1 U12568 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n12029), .A(n10027), .ZN(
        n10028) );
  OAI211_X1 U12569 ( .C1(n10220), .C2(n13737), .A(n10029), .B(n10028), .ZN(
        P1_U3222) );
  NAND2_X1 U12570 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n10423) );
  AOI211_X1 U12571 ( .C1(n10032), .C2(n10031), .A(n10030), .B(n14713), .ZN(
        n10033) );
  INV_X1 U12572 ( .A(n10033), .ZN(n10034) );
  NAND2_X1 U12573 ( .A1(n10423), .A2(n10034), .ZN(n10041) );
  MUX2_X1 U12574 ( .A(n9837), .B(P2_REG1_REG_6__SCAN_IN), .S(n10035), .Z(
        n10036) );
  NAND3_X1 U12575 ( .A1(n14710), .A2(n10037), .A3(n10036), .ZN(n10038) );
  AND3_X1 U12576 ( .A1(n14783), .A2(n10039), .A3(n10038), .ZN(n10040) );
  AOI211_X1 U12577 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n14775), .A(n10041), .B(
        n10040), .ZN(n10042) );
  OAI21_X1 U12578 ( .B1(n10043), .B2(n14707), .A(n10042), .ZN(P2_U3220) );
  INV_X1 U12579 ( .A(n13595), .ZN(n10047) );
  XNOR2_X1 U12580 ( .A(n11776), .B(P2_B_REG_SCAN_IN), .ZN(n10045) );
  INV_X1 U12581 ( .A(n10044), .ZN(n11861) );
  NAND2_X1 U12582 ( .A1(n10045), .A2(n11861), .ZN(n10046) );
  OR2_X1 U12583 ( .A1(n14790), .A2(P2_D_REG_1__SCAN_IN), .ZN(n10049) );
  NAND2_X1 U12584 ( .A1(n13595), .A2(n11861), .ZN(n10048) );
  AND2_X1 U12585 ( .A1(n10049), .A2(n10048), .ZN(n10113) );
  INV_X1 U12586 ( .A(n10113), .ZN(n10050) );
  INV_X1 U12587 ( .A(n6477), .ZN(n11456) );
  NAND2_X1 U12588 ( .A1(n14840), .A2(n11257), .ZN(n10114) );
  NAND2_X1 U12589 ( .A1(n10050), .A2(n10114), .ZN(n10131) );
  INV_X1 U12590 ( .A(n14795), .ZN(n10051) );
  NOR2_X1 U12591 ( .A1(n10131), .A2(n10051), .ZN(n10139) );
  NOR4_X1 U12592 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n10060) );
  OR4_X1 U12593 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n10057) );
  NOR4_X1 U12594 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n10055) );
  NOR4_X1 U12595 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n10054) );
  NOR4_X1 U12596 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n10053) );
  NOR4_X1 U12597 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n10052) );
  NAND4_X1 U12598 ( .A1(n10055), .A2(n10054), .A3(n10053), .A4(n10052), .ZN(
        n10056) );
  NOR4_X1 U12599 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n10057), .A4(n10056), .ZN(n10059) );
  NOR4_X1 U12600 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n10058) );
  AND3_X1 U12601 ( .A1(n10060), .A2(n10059), .A3(n10058), .ZN(n10061) );
  NOR2_X1 U12602 ( .A1(n14790), .A2(n10061), .ZN(n10136) );
  OR2_X1 U12603 ( .A1(n14790), .A2(P2_D_REG_0__SCAN_IN), .ZN(n10062) );
  NAND2_X1 U12604 ( .A1(n13595), .A2(n11776), .ZN(n14792) );
  NAND2_X1 U12605 ( .A1(n10062), .A2(n14792), .ZN(n10137) );
  INV_X1 U12606 ( .A(n10125), .ZN(n10118) );
  NAND2_X1 U12607 ( .A1(n10114), .A2(n10118), .ZN(n10063) );
  NAND2_X1 U12608 ( .A1(n10119), .A2(n10077), .ZN(n10134) );
  AND2_X1 U12609 ( .A1(n10063), .A2(n10134), .ZN(n10128) );
  OAI21_X1 U12610 ( .B1(n10064), .B2(n10185), .A(n10141), .ZN(n10589) );
  INV_X1 U12611 ( .A(n10589), .ZN(n10083) );
  AND2_X1 U12612 ( .A1(n6477), .A2(n10178), .ZN(n10066) );
  INV_X1 U12613 ( .A(n10179), .ZN(n14823) );
  INV_X1 U12614 ( .A(n13203), .ZN(n10069) );
  INV_X1 U12615 ( .A(n13166), .ZN(n13142) );
  INV_X1 U12616 ( .A(n10068), .ZN(n10164) );
  INV_X1 U12617 ( .A(n13167), .ZN(n13144) );
  OAI22_X1 U12618 ( .A1(n10069), .A2(n13142), .B1(n10164), .B2(n13144), .ZN(
        n10177) );
  INV_X1 U12619 ( .A(n10070), .ZN(n10123) );
  NAND2_X1 U12620 ( .A1(n10064), .A2(n10123), .ZN(n10074) );
  NAND2_X1 U12621 ( .A1(n6477), .A2(n10332), .ZN(n10073) );
  AOI21_X1 U12622 ( .B1(n10074), .B2(n10145), .A(n13430), .ZN(n10075) );
  AOI211_X1 U12623 ( .C1(n14823), .C2(n10589), .A(n10177), .B(n10075), .ZN(
        n10594) );
  NOR2_X2 U12624 ( .A1(n6477), .A2(n10076), .ZN(n10561) );
  NAND2_X1 U12625 ( .A1(n10337), .A2(n10078), .ZN(n10080) );
  NAND2_X1 U12626 ( .A1(n10080), .A2(n11850), .ZN(n10081) );
  NOR2_X1 U12627 ( .A1(n10148), .A2(n10081), .ZN(n10588) );
  AOI21_X1 U12628 ( .B1(n14816), .B2(n10078), .A(n10588), .ZN(n10082) );
  OAI211_X1 U12629 ( .C1(n10083), .C2(n14819), .A(n10594), .B(n10082), .ZN(
        n10595) );
  NAND2_X1 U12630 ( .A1(n10595), .A2(n14855), .ZN(n10084) );
  OAI21_X1 U12631 ( .B1(n14855), .B2(n9826), .A(n10084), .ZN(P2_U3500) );
  INV_X1 U12632 ( .A(n14749), .ZN(n10986) );
  OAI222_X1 U12633 ( .A1(n13593), .A2(n10086), .B1(n13587), .B2(n10085), .C1(
        n10986), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U12634 ( .A(n10087), .ZN(n10089) );
  OAI222_X1 U12635 ( .A1(n12618), .A2(P3_U3151), .B1(n13067), .B2(n10089), 
        .C1(n10088), .C2(n13059), .ZN(P3_U3278) );
  INV_X1 U12636 ( .A(n14722), .ZN(n14730) );
  AOI21_X1 U12637 ( .B1(n10094), .B2(P2_REG2_REG_8__SCAN_IN), .A(n10090), .ZN(
        n14728) );
  MUX2_X1 U12638 ( .A(n10738), .B(P2_REG2_REG_9__SCAN_IN), .S(n14722), .Z(
        n14727) );
  NAND2_X1 U12639 ( .A1(n14728), .A2(n14727), .ZN(n14726) );
  OAI21_X1 U12640 ( .B1(n14730), .B2(P2_REG2_REG_9__SCAN_IN), .A(n14726), .ZN(
        n10092) );
  MUX2_X1 U12641 ( .A(n7737), .B(P2_REG2_REG_10__SCAN_IN), .S(n10980), .Z(
        n10091) );
  NOR2_X1 U12642 ( .A1(n10092), .A2(n10091), .ZN(n10973) );
  AOI211_X1 U12643 ( .C1(n10092), .C2(n10091), .A(n14713), .B(n10973), .ZN(
        n10093) );
  INV_X1 U12644 ( .A(n10093), .ZN(n10106) );
  NAND2_X1 U12645 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n10865)
         );
  INV_X1 U12646 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n14851) );
  MUX2_X1 U12647 ( .A(n14851), .B(P2_REG1_REG_10__SCAN_IN), .S(n10980), .Z(
        n10100) );
  NAND2_X1 U12648 ( .A1(n10094), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10095) );
  NAND2_X1 U12649 ( .A1(n10096), .A2(n10095), .ZN(n14721) );
  INV_X1 U12650 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10097) );
  MUX2_X1 U12651 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10097), .S(n14722), .Z(
        n10098) );
  OR2_X1 U12652 ( .A1(n14721), .A2(n10098), .ZN(n14723) );
  NAND2_X1 U12653 ( .A1(n14722), .A2(n10097), .ZN(n10099) );
  NAND2_X1 U12654 ( .A1(n14723), .A2(n10099), .ZN(n10101) );
  AOI21_X1 U12655 ( .B1(n10100), .B2(n10101), .A(n14746), .ZN(n10102) );
  NAND2_X1 U12656 ( .A1(n10102), .A2(n13225), .ZN(n10103) );
  NAND2_X1 U12657 ( .A1(n10865), .A2(n10103), .ZN(n10104) );
  AOI21_X1 U12658 ( .B1(n14775), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10104), 
        .ZN(n10105) );
  OAI211_X1 U12659 ( .C1(n14707), .C2(n10107), .A(n10106), .B(n10105), .ZN(
        P2_U3224) );
  INV_X1 U12660 ( .A(n10108), .ZN(n10110) );
  OAI222_X1 U12661 ( .A1(P1_U3086), .A2(n11881), .B1(n14183), .B2(n10110), 
        .C1(n10109), .C2(n14180), .ZN(P1_U3342) );
  OAI222_X1 U12662 ( .A1(n13593), .A2(n10111), .B1(n13587), .B2(n10110), .C1(
        n10987), .C2(P2_U3088), .ZN(P2_U3314) );
  OAI222_X1 U12663 ( .A1(P3_U3151), .A2(n12614), .B1(n13070), .B2(n15126), 
        .C1(n13067), .C2(n10112), .ZN(P3_U3277) );
  NAND3_X1 U12664 ( .A1(n10561), .A2(n10560), .A3(n10125), .ZN(n10116) );
  OAI21_X2 U12665 ( .B1(n14793), .B2(n10116), .A(n13385), .ZN(n14669) );
  NAND2_X1 U12666 ( .A1(n13203), .A2(n13412), .ZN(n10117) );
  MUX2_X1 U12667 ( .A(n10117), .B(n13412), .S(n10337), .Z(n10122) );
  INV_X1 U12668 ( .A(n14793), .ZN(n10330) );
  NOR2_X1 U12669 ( .A1(n10119), .A2(n10118), .ZN(n10120) );
  AND2_X1 U12670 ( .A1(n14837), .A2(n10120), .ZN(n10121) );
  AOI21_X1 U12671 ( .B1(n10123), .B2(n10122), .A(n14664), .ZN(n10124) );
  AOI21_X1 U12672 ( .B1(n10337), .B2(n14669), .A(n10124), .ZN(n10133) );
  NAND2_X1 U12673 ( .A1(n10126), .A2(n10125), .ZN(n10127) );
  NOR2_X2 U12674 ( .A1(n14793), .A2(n10127), .ZN(n14386) );
  AND2_X1 U12675 ( .A1(n13202), .A2(n13167), .ZN(n10334) );
  AND2_X1 U12676 ( .A1(n10129), .A2(n10128), .ZN(n10130) );
  AND2_X1 U12677 ( .A1(n10131), .A2(n10130), .ZN(n10205) );
  NAND2_X1 U12678 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10205), .ZN(n11915) );
  AOI22_X1 U12679 ( .A1(n14386), .A2(n10334), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n11915), .ZN(n10132) );
  NAND2_X1 U12680 ( .A1(n10133), .A2(n10132), .ZN(P2_U3204) );
  INV_X1 U12681 ( .A(n10134), .ZN(n10135) );
  NOR2_X1 U12682 ( .A1(n10136), .A2(n10135), .ZN(n10138) );
  INV_X1 U12683 ( .A(n13202), .ZN(n10146) );
  NAND2_X1 U12684 ( .A1(n10146), .A2(n10194), .ZN(n10140) );
  OAI21_X1 U12685 ( .B1(n10143), .B2(n10142), .A(n10157), .ZN(n13456) );
  INV_X1 U12686 ( .A(n13456), .ZN(n10152) );
  NAND2_X1 U12687 ( .A1(n10146), .A2(n10078), .ZN(n10144) );
  XNOR2_X1 U12688 ( .A(n10163), .B(n10162), .ZN(n10147) );
  OAI22_X1 U12689 ( .A1(n10146), .A2(n13142), .B1(n10545), .B2(n13144), .ZN(
        n11916) );
  AOI21_X1 U12690 ( .B1(n10147), .B2(n13437), .A(n11916), .ZN(n13461) );
  NAND2_X1 U12691 ( .A1(n7048), .A2(n10148), .ZN(n10160) );
  INV_X1 U12692 ( .A(n10148), .ZN(n10149) );
  NAND2_X1 U12693 ( .A1(n10149), .A2(n13459), .ZN(n10150) );
  AND3_X1 U12694 ( .A1(n10160), .A2(n10150), .A3(n11850), .ZN(n13454) );
  AOI21_X1 U12695 ( .B1(n14816), .B2(n13459), .A(n13454), .ZN(n10151) );
  OAI211_X1 U12696 ( .C1(n10152), .C2(n14812), .A(n13461), .B(n10151), .ZN(
        n13556) );
  NAND2_X1 U12697 ( .A1(n13556), .A2(n14835), .ZN(n10153) );
  OAI21_X1 U12698 ( .B1(n14835), .B2(n7520), .A(n10153), .ZN(P2_U3436) );
  OAI222_X1 U12699 ( .A1(P3_U3151), .A2(n12193), .B1(n13067), .B2(n10155), 
        .C1(n10154), .C2(n13059), .ZN(P3_U3276) );
  NAND2_X1 U12700 ( .A1(n7048), .A2(n10164), .ZN(n10156) );
  NAND2_X1 U12701 ( .A1(n10157), .A2(n10156), .ZN(n10158) );
  NAND2_X1 U12702 ( .A1(n10158), .A2(n10167), .ZN(n10541) );
  OR2_X1 U12703 ( .A1(n10158), .A2(n10167), .ZN(n10159) );
  NAND2_X1 U12704 ( .A1(n10541), .A2(n10159), .ZN(n10848) );
  AOI21_X1 U12705 ( .B1(n10160), .B2(n10843), .A(n13412), .ZN(n10161) );
  NAND2_X1 U12706 ( .A1(n10161), .A2(n10602), .ZN(n10845) );
  OAI21_X1 U12707 ( .B1(n6956), .B2(n14837), .A(n10845), .ZN(n10175) );
  NAND2_X1 U12708 ( .A1(n10848), .A2(n14823), .ZN(n10174) );
  NAND2_X1 U12709 ( .A1(n10163), .A2(n10162), .ZN(n10166) );
  NAND2_X1 U12710 ( .A1(n10164), .A2(n13459), .ZN(n10165) );
  INV_X1 U12711 ( .A(n10167), .ZN(n10168) );
  OAI21_X1 U12712 ( .B1(n10169), .B2(n10168), .A(n10609), .ZN(n10172) );
  NAND2_X1 U12713 ( .A1(n13200), .A2(n13167), .ZN(n10171) );
  NAND2_X1 U12714 ( .A1(n10068), .A2(n13166), .ZN(n10170) );
  NAND2_X1 U12715 ( .A1(n10171), .A2(n10170), .ZN(n10206) );
  AOI21_X1 U12716 ( .B1(n10172), .B2(n13437), .A(n10206), .ZN(n10173) );
  NAND2_X1 U12717 ( .A1(n10174), .A2(n10173), .ZN(n10842) );
  AOI211_X1 U12718 ( .C1(n14840), .C2(n10848), .A(n10175), .B(n10842), .ZN(
        n10344) );
  NAND2_X1 U12719 ( .A1(n14853), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10176) );
  OAI21_X1 U12720 ( .B1(n10344), .B2(n14853), .A(n10176), .ZN(P2_U3502) );
  AOI22_X1 U12721 ( .A1(n14386), .A2(n10177), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n11915), .ZN(n10193) );
  NAND2_X1 U12722 ( .A1(n10179), .A2(n10178), .ZN(n10197) );
  XNOR2_X1 U12723 ( .A(n10194), .B(n10197), .ZN(n10181) );
  NAND2_X1 U12724 ( .A1(n13202), .A2(n10760), .ZN(n10180) );
  NAND2_X1 U12725 ( .A1(n10181), .A2(n10180), .ZN(n10195) );
  INV_X1 U12726 ( .A(n10180), .ZN(n10183) );
  INV_X1 U12727 ( .A(n10181), .ZN(n10182) );
  NAND2_X1 U12728 ( .A1(n10183), .A2(n10182), .ZN(n10184) );
  NAND2_X1 U12729 ( .A1(n10195), .A2(n10184), .ZN(n10189) );
  INV_X1 U12730 ( .A(n10189), .ZN(n10187) );
  NAND2_X1 U12731 ( .A1(n10187), .A2(n10186), .ZN(n10196) );
  INV_X1 U12732 ( .A(n10196), .ZN(n10191) );
  AND2_X1 U12733 ( .A1(n10189), .A2(n10188), .ZN(n10190) );
  OAI21_X1 U12734 ( .B1(n10191), .B2(n10190), .A(n14384), .ZN(n10192) );
  OAI211_X1 U12735 ( .C1(n13162), .C2(n10194), .A(n10193), .B(n10192), .ZN(
        P2_U3194) );
  NAND2_X1 U12736 ( .A1(n10196), .A2(n10195), .ZN(n11918) );
  XNOR2_X1 U12737 ( .A(n13459), .B(n10204), .ZN(n10198) );
  NAND2_X1 U12738 ( .A1(n10068), .A2(n10760), .ZN(n10199) );
  NAND2_X1 U12739 ( .A1(n10198), .A2(n10199), .ZN(n10203) );
  INV_X1 U12740 ( .A(n10198), .ZN(n10201) );
  INV_X1 U12741 ( .A(n10199), .ZN(n10200) );
  NAND2_X1 U12742 ( .A1(n10201), .A2(n10200), .ZN(n10202) );
  NAND2_X1 U12743 ( .A1(n11918), .A2(n11919), .ZN(n11917) );
  XNOR2_X1 U12744 ( .A(n10843), .B(n6488), .ZN(n10288) );
  NAND2_X1 U12745 ( .A1(n13201), .A2(n10760), .ZN(n10287) );
  XNOR2_X1 U12746 ( .A(n10288), .B(n10287), .ZN(n10289) );
  XNOR2_X1 U12747 ( .A(n10290), .B(n10289), .ZN(n10211) );
  INV_X1 U12748 ( .A(n14672), .ZN(n13159) );
  INV_X1 U12749 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n14694) );
  NAND2_X1 U12750 ( .A1(n14669), .A2(n10843), .ZN(n10208) );
  NAND2_X1 U12751 ( .A1(n14386), .A2(n10206), .ZN(n10207) );
  OAI211_X1 U12752 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n14694), .A(n10208), .B(
        n10207), .ZN(n10209) );
  AOI21_X1 U12753 ( .B1(n13159), .B2(n14694), .A(n10209), .ZN(n10210) );
  OAI21_X1 U12754 ( .B1(n10211), .B2(n14664), .A(n10210), .ZN(P2_U3190) );
  NAND2_X1 U12755 ( .A1(n10474), .A2(n10321), .ZN(n10212) );
  NOR2_X1 U12756 ( .A1(n10213), .A2(n10212), .ZN(n10215) );
  AND2_X1 U12757 ( .A1(n10215), .A2(n10214), .ZN(n10247) );
  INV_X1 U12758 ( .A(n14636), .ZN(n14609) );
  AND2_X1 U12759 ( .A1(n10216), .A2(n11165), .ZN(n10217) );
  NAND2_X1 U12760 ( .A1(n12141), .A2(n10217), .ZN(n14545) );
  OR2_X1 U12761 ( .A1(n14047), .A2(n10218), .ZN(n14060) );
  NAND2_X1 U12762 ( .A1(n14563), .A2(n10220), .ZN(n10221) );
  NAND2_X1 U12763 ( .A1(n10478), .A2(n10223), .ZN(n10225) );
  INV_X2 U12764 ( .A(n10490), .ZN(n14595) );
  NAND2_X1 U12765 ( .A1(n14595), .A2(n7406), .ZN(n10224) );
  NAND2_X1 U12766 ( .A1(n10225), .A2(n10224), .ZN(n14544) );
  INV_X1 U12767 ( .A(n10226), .ZN(n10227) );
  OR2_X1 U12768 ( .A1(n14554), .A2(n13754), .ZN(n10228) );
  XNOR2_X1 U12769 ( .A(n10464), .B(n10237), .ZN(n14535) );
  NAND2_X1 U12770 ( .A1(n14595), .A2(n6491), .ZN(n14553) );
  NOR2_X2 U12771 ( .A1(n10239), .A2(n10229), .ZN(n14556) );
  AOI211_X1 U12772 ( .C1(n10674), .C2(n14555), .A(n14058), .B(n10466), .ZN(
        n14533) );
  AOI21_X1 U12773 ( .B1(n10674), .B2(n14606), .A(n14533), .ZN(n10245) );
  NAND2_X1 U12774 ( .A1(n10231), .A2(n10230), .ZN(n10232) );
  AND2_X1 U12775 ( .A1(n9605), .A2(n10232), .ZN(n10480) );
  NAND2_X1 U12776 ( .A1(n10480), .A2(n10233), .ZN(n10479) );
  NAND2_X1 U12777 ( .A1(n14554), .A2(n10235), .ZN(n10236) );
  XNOR2_X1 U12778 ( .A(n10458), .B(n10237), .ZN(n10244) );
  NAND2_X1 U12779 ( .A1(n10239), .A2(n10238), .ZN(n10241) );
  NAND2_X1 U12780 ( .A1(n13826), .A2(n14189), .ZN(n10240) );
  NAND2_X2 U12781 ( .A1(n10241), .A2(n10240), .ZN(n14549) );
  NAND2_X1 U12782 ( .A1(n13752), .A2(n14055), .ZN(n10243) );
  NAND2_X1 U12783 ( .A1(n13754), .A2(n14033), .ZN(n10242) );
  NAND2_X1 U12784 ( .A1(n10243), .A2(n10242), .ZN(n10675) );
  AOI21_X1 U12785 ( .B1(n10244), .B2(n14549), .A(n10675), .ZN(n14539) );
  OAI211_X1 U12786 ( .C1(n14581), .C2(n14535), .A(n10245), .B(n14539), .ZN(
        n10248) );
  NAND2_X1 U12787 ( .A1(n10248), .A2(n14657), .ZN(n10246) );
  OAI21_X1 U12788 ( .B1(n14657), .B2(n9170), .A(n10246), .ZN(P1_U3532) );
  INV_X1 U12789 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U12790 ( .A1(n10248), .A2(n14646), .ZN(n10249) );
  OAI21_X1 U12791 ( .B1(n14646), .B2(n10250), .A(n10249), .ZN(P1_U3471) );
  OR2_X1 U12792 ( .A1(n10252), .A2(P3_U3151), .ZN(n12369) );
  INV_X1 U12793 ( .A(n12369), .ZN(n10251) );
  OR2_X1 U12794 ( .A1(n10714), .A2(n10251), .ZN(n10262) );
  NAND2_X1 U12795 ( .A1(n12346), .A2(n10252), .ZN(n10253) );
  NAND2_X1 U12796 ( .A1(n6653), .A2(n10253), .ZN(n10261) );
  INV_X1 U12797 ( .A(n10261), .ZN(n10255) );
  INV_X1 U12798 ( .A(n10259), .ZN(n10256) );
  MUX2_X1 U12799 ( .A(n10256), .B(n12522), .S(n12364), .Z(n14970) );
  INV_X1 U12800 ( .A(n10257), .ZN(n10258) );
  AND2_X1 U12801 ( .A1(n10259), .A2(n10258), .ZN(n14353) );
  NAND2_X1 U12802 ( .A1(n10259), .A2(n12601), .ZN(n12623) );
  NAND3_X1 U12803 ( .A1(n14959), .A2(n14939), .A3(n12623), .ZN(n10265) );
  MUX2_X1 U12804 ( .A(n10358), .B(n10352), .S(n12601), .Z(n10260) );
  AND2_X1 U12805 ( .A1(n10260), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10346) );
  INV_X1 U12806 ( .A(n10346), .ZN(n10403) );
  OAI21_X1 U12807 ( .B1(P3_IR_REG_0__SCAN_IN), .B2(n10260), .A(n10403), .ZN(
        n10264) );
  OAI22_X1 U12808 ( .A1(n14975), .A2(n14246), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10716), .ZN(n10263) );
  AOI21_X1 U12809 ( .B1(n10265), .B2(n10264), .A(n10263), .ZN(n10266) );
  OAI21_X1 U12810 ( .B1(n10351), .B2(n14970), .A(n10266), .ZN(P3_U3182) );
  INV_X1 U12811 ( .A(n11133), .ZN(n11141) );
  AOI22_X1 U12812 ( .A1(n11133), .A2(n9322), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n11141), .ZN(n10271) );
  AOI21_X1 U12813 ( .B1(n9995), .B2(n10268), .A(n10267), .ZN(n11876) );
  MUX2_X1 U12814 ( .A(n10269), .B(P1_REG1_REG_13__SCAN_IN), .S(n11881), .Z(
        n11875) );
  NAND2_X1 U12815 ( .A1(n11876), .A2(n11875), .ZN(n11874) );
  OAI21_X1 U12816 ( .B1(n11881), .B2(n10269), .A(n11874), .ZN(n10270) );
  NOR2_X1 U12817 ( .A1(n10271), .A2(n10270), .ZN(n11140) );
  AOI21_X1 U12818 ( .B1(n10271), .B2(n10270), .A(n11140), .ZN(n10281) );
  INV_X1 U12819 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14229) );
  NAND2_X1 U12820 ( .A1(n14492), .A2(n11133), .ZN(n10272) );
  NAND2_X1 U12821 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14416)
         );
  OAI211_X1 U12822 ( .C1(n14229), .C2(n14525), .A(n10272), .B(n14416), .ZN(
        n10273) );
  INV_X1 U12823 ( .A(n10273), .ZN(n10280) );
  OAI21_X1 U12824 ( .B1(n10275), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10274), 
        .ZN(n11871) );
  MUX2_X1 U12825 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n9330), .S(n11881), .Z(
        n11870) );
  OR2_X1 U12826 ( .A1(n11871), .A2(n11870), .ZN(n11872) );
  OAI21_X1 U12827 ( .B1(n9330), .B2(n11881), .A(n11872), .ZN(n10278) );
  MUX2_X1 U12828 ( .A(n11676), .B(P1_REG2_REG_14__SCAN_IN), .S(n11133), .Z(
        n10276) );
  INV_X1 U12829 ( .A(n10276), .ZN(n10277) );
  NAND2_X1 U12830 ( .A1(n10277), .A2(n10278), .ZN(n11134) );
  OAI211_X1 U12831 ( .C1(n10278), .C2(n10277), .A(n14483), .B(n11134), .ZN(
        n10279) );
  OAI211_X1 U12832 ( .C1(n10281), .C2(n14517), .A(n10280), .B(n10279), .ZN(
        P1_U3257) );
  XNOR2_X1 U12833 ( .A(n14808), .B(n6487), .ZN(n10282) );
  NAND2_X1 U12834 ( .A1(n13199), .A2(n10760), .ZN(n10283) );
  NAND2_X1 U12835 ( .A1(n10282), .A2(n10283), .ZN(n10419) );
  INV_X1 U12836 ( .A(n10282), .ZN(n10285) );
  INV_X1 U12837 ( .A(n10283), .ZN(n10284) );
  NAND2_X1 U12838 ( .A1(n10285), .A2(n10284), .ZN(n10286) );
  AND2_X1 U12839 ( .A1(n10419), .A2(n10286), .ZN(n10299) );
  XNOR2_X1 U12840 ( .A(n14802), .B(n6488), .ZN(n10291) );
  NAND2_X1 U12841 ( .A1(n13200), .A2(n10760), .ZN(n10292) );
  NAND2_X1 U12842 ( .A1(n10291), .A2(n10292), .ZN(n10297) );
  INV_X1 U12843 ( .A(n10291), .ZN(n10294) );
  INV_X1 U12844 ( .A(n10292), .ZN(n10293) );
  NAND2_X1 U12845 ( .A1(n10294), .A2(n10293), .ZN(n10295) );
  NAND2_X1 U12846 ( .A1(n10297), .A2(n10295), .ZN(n10397) );
  NAND2_X1 U12847 ( .A1(n10395), .A2(n10297), .ZN(n10298) );
  OAI21_X1 U12848 ( .B1(n10299), .B2(n10298), .A(n10420), .ZN(n10300) );
  NAND2_X1 U12849 ( .A1(n10300), .A2(n14384), .ZN(n10305) );
  NAND2_X1 U12850 ( .A1(n13198), .A2(n13167), .ZN(n10302) );
  NAND2_X1 U12851 ( .A1(n13200), .A2(n13166), .ZN(n10301) );
  NAND2_X1 U12852 ( .A1(n10302), .A2(n10301), .ZN(n10555) );
  AND2_X1 U12853 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n14709) );
  NOR2_X1 U12854 ( .A1(n14672), .A2(n10563), .ZN(n10303) );
  AOI211_X1 U12855 ( .C1(n14386), .C2(n10555), .A(n14709), .B(n10303), .ZN(
        n10304) );
  OAI211_X1 U12856 ( .C1(n10570), .C2(n13162), .A(n10305), .B(n10304), .ZN(
        P2_U3199) );
  AOI22_X1 U12857 ( .A1(n14554), .A2(n10630), .B1(n12147), .B2(n13754), .ZN(
        n10626) );
  NAND2_X1 U12858 ( .A1(n14554), .A2(n12146), .ZN(n10307) );
  NAND2_X1 U12859 ( .A1(n13754), .A2(n10630), .ZN(n10306) );
  NAND2_X1 U12860 ( .A1(n10307), .A2(n10306), .ZN(n10308) );
  XNOR2_X1 U12861 ( .A(n10308), .B(n12141), .ZN(n10627) );
  XOR2_X1 U12862 ( .A(n10626), .B(n10627), .Z(n10320) );
  INV_X1 U12863 ( .A(n10309), .ZN(n10310) );
  NAND2_X1 U12864 ( .A1(n10311), .A2(n10310), .ZN(n12025) );
  NAND2_X1 U12865 ( .A1(n10490), .A2(n12146), .ZN(n10313) );
  NAND2_X1 U12866 ( .A1(n10313), .A2(n10312), .ZN(n10314) );
  XNOR2_X1 U12867 ( .A(n10314), .B(n12141), .ZN(n10317) );
  XNOR2_X1 U12868 ( .A(n10317), .B(n10315), .ZN(n12026) );
  NAND2_X1 U12869 ( .A1(n12025), .A2(n12026), .ZN(n12024) );
  NAND2_X1 U12870 ( .A1(n12024), .A2(n10318), .ZN(n10319) );
  NOR2_X1 U12871 ( .A1(n10319), .A2(n10320), .ZN(n10629) );
  AOI211_X1 U12872 ( .C1(n10320), .C2(n10319), .A(n14426), .B(n10629), .ZN(
        n10329) );
  INV_X1 U12873 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14551) );
  NAND4_X1 U12874 ( .A1(n10324), .A2(n10323), .A3(n10322), .A4(n10321), .ZN(
        n10325) );
  INV_X1 U12875 ( .A(n14436), .ZN(n13733) );
  AOI22_X1 U12876 ( .A1(n14551), .A2(n13733), .B1(n14432), .B2(n14554), .ZN(
        n10327) );
  AOI22_X1 U12877 ( .A1(n13729), .A2(n13753), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10326) );
  OAI211_X1 U12878 ( .C1(n7406), .C2(n14419), .A(n10327), .B(n10326), .ZN(
        n10328) );
  OR2_X1 U12879 ( .A1(n10329), .A2(n10328), .ZN(P1_U3218) );
  NAND2_X1 U12880 ( .A1(n10336), .A2(n10330), .ZN(n10331) );
  NAND2_X1 U12881 ( .A1(n10333), .A2(n10332), .ZN(n10543) );
  OR2_X1 U12882 ( .A1(n13453), .A2(n10543), .ZN(n13361) );
  AOI21_X1 U12883 ( .B1(n13430), .B2(n10179), .A(n14798), .ZN(n10335) );
  NOR2_X1 U12884 ( .A1(n10335), .A2(n10334), .ZN(n14797) );
  INV_X1 U12885 ( .A(n13385), .ZN(n13458) );
  INV_X1 U12886 ( .A(n10336), .ZN(n10339) );
  NAND2_X1 U12887 ( .A1(n10337), .A2(n10561), .ZN(n14796) );
  NOR4_X1 U12888 ( .A1(n10339), .A2(n10338), .A3(n14793), .A4(n14796), .ZN(
        n10340) );
  AOI21_X1 U12889 ( .B1(n13458), .B2(P2_REG3_REG_0__SCAN_IN), .A(n10340), .ZN(
        n10341) );
  OAI21_X1 U12890 ( .B1(n13453), .B2(n14797), .A(n10341), .ZN(n10342) );
  AOI21_X1 U12891 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n13453), .A(n10342), .ZN(
        n10343) );
  OAI21_X1 U12892 ( .B1(n14798), .B2(n13361), .A(n10343), .ZN(P2_U3265) );
  INV_X1 U12893 ( .A(n14835), .ZN(n14844) );
  OR2_X1 U12894 ( .A1(n10344), .A2(n14844), .ZN(n10345) );
  OAI21_X1 U12895 ( .B1(n14835), .B2(n7562), .A(n10345), .ZN(P2_U3439) );
  MUX2_X1 U12896 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12601), .Z(n10374) );
  XNOR2_X1 U12897 ( .A(n10374), .B(n6483), .ZN(n10372) );
  INV_X1 U12898 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10408) );
  MUX2_X1 U12899 ( .A(n10880), .B(n10408), .S(n12601), .Z(n10347) );
  NAND2_X1 U12900 ( .A1(n10404), .A2(n10346), .ZN(n10349) );
  INV_X1 U12901 ( .A(n10360), .ZN(n10416) );
  NAND2_X1 U12902 ( .A1(n10347), .A2(n10416), .ZN(n10348) );
  NAND2_X1 U12903 ( .A1(n10349), .A2(n10348), .ZN(n10373) );
  XOR2_X1 U12904 ( .A(n10372), .B(n10373), .Z(n10371) );
  INV_X1 U12905 ( .A(n14970), .ZN(n14343) );
  MUX2_X1 U12906 ( .A(n10350), .B(P3_REG1_REG_2__SCAN_IN), .S(n6483), .Z(
        n10356) );
  AND2_X1 U12907 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10351), .ZN(n10353) );
  OR3_X1 U12908 ( .A1(n10352), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n10354) );
  OAI21_X1 U12909 ( .B1(n10360), .B2(n10353), .A(n10354), .ZN(n10407) );
  OR2_X1 U12910 ( .A1(n10407), .A2(n10408), .ZN(n10405) );
  NAND2_X1 U12911 ( .A1(n10405), .A2(n10354), .ZN(n10355) );
  NAND2_X1 U12912 ( .A1(n10356), .A2(n10355), .ZN(n10380) );
  OAI21_X1 U12913 ( .B1(n10356), .B2(n10355), .A(n10380), .ZN(n10357) );
  INV_X1 U12914 ( .A(n10357), .ZN(n10368) );
  XNOR2_X1 U12915 ( .A(n6483), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n10363) );
  NOR2_X1 U12916 ( .A1(n10358), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10359) );
  NAND2_X1 U12917 ( .A1(n8416), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10361) );
  OAI21_X1 U12918 ( .B1(n10360), .B2(n10359), .A(n10361), .ZN(n10411) );
  OR2_X1 U12919 ( .A1(n10411), .A2(n10880), .ZN(n10413) );
  NAND2_X1 U12920 ( .A1(n10413), .A2(n10361), .ZN(n10362) );
  NAND2_X1 U12921 ( .A1(n10363), .A2(n10362), .ZN(n10384) );
  OAI21_X1 U12922 ( .B1(n10363), .B2(n10362), .A(n10384), .ZN(n10364) );
  NAND2_X1 U12923 ( .A1(n14353), .A2(n10364), .ZN(n10367) );
  NOR2_X1 U12924 ( .A1(n11063), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10365) );
  AOI21_X1 U12925 ( .B1(n14943), .B2(P3_ADDR_REG_2__SCAN_IN), .A(n10365), .ZN(
        n10366) );
  OAI211_X1 U12926 ( .C1(n10368), .C2(n12623), .A(n10367), .B(n10366), .ZN(
        n10369) );
  AOI21_X1 U12927 ( .B1(n14343), .B2(n6483), .A(n10369), .ZN(n10370) );
  OAI21_X1 U12928 ( .B1(n10371), .B2(n14939), .A(n10370), .ZN(P3_U3184) );
  MUX2_X1 U12929 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12601), .Z(n10436) );
  INV_X1 U12930 ( .A(n10442), .ZN(n10437) );
  XNOR2_X1 U12931 ( .A(n10436), .B(n10437), .ZN(n10434) );
  NAND2_X1 U12932 ( .A1(n10373), .A2(n10372), .ZN(n10377) );
  INV_X1 U12933 ( .A(n10374), .ZN(n10375) );
  NAND2_X1 U12934 ( .A1(n10375), .A2(n6483), .ZN(n10376) );
  NAND2_X1 U12935 ( .A1(n10377), .A2(n10376), .ZN(n10435) );
  XOR2_X1 U12936 ( .A(n10434), .B(n10435), .Z(n10394) );
  INV_X1 U12937 ( .A(n6483), .ZN(n10382) );
  NAND2_X1 U12938 ( .A1(n10382), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10379) );
  NAND2_X1 U12939 ( .A1(n10380), .A2(n10379), .ZN(n10441) );
  XNOR2_X1 U12940 ( .A(n10443), .B(n10381), .ZN(n10391) );
  NAND2_X1 U12941 ( .A1(n10382), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10383) );
  NAND2_X1 U12942 ( .A1(n10384), .A2(n10383), .ZN(n10385) );
  NAND2_X1 U12943 ( .A1(n10386), .A2(n10829), .ZN(n10387) );
  NAND2_X1 U12944 ( .A1(n6631), .A2(n10387), .ZN(n10388) );
  NAND2_X1 U12945 ( .A1(n14353), .A2(n10388), .ZN(n10390) );
  NOR2_X1 U12946 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8365), .ZN(n10784) );
  AOI21_X1 U12947 ( .B1(n14943), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10784), .ZN(
        n10389) );
  OAI211_X1 U12948 ( .C1(n10391), .C2(n12623), .A(n10390), .B(n10389), .ZN(
        n10392) );
  AOI21_X1 U12949 ( .B1(n14343), .B2(n10437), .A(n10392), .ZN(n10393) );
  OAI21_X1 U12950 ( .B1(n10394), .B2(n14939), .A(n10393), .ZN(P3_U3185) );
  INV_X1 U12951 ( .A(n10395), .ZN(n10396) );
  AOI21_X1 U12952 ( .B1(n10398), .B2(n10397), .A(n10396), .ZN(n10402) );
  OAI22_X1 U12953 ( .A1(n10545), .A2(n13142), .B1(n10569), .B2(n13144), .ZN(
        n10611) );
  AND2_X1 U12954 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n13209) );
  AOI21_X1 U12955 ( .B1(n14386), .B2(n10611), .A(n13209), .ZN(n10399) );
  OAI21_X1 U12956 ( .B1(n13162), .B2(n10605), .A(n10399), .ZN(n10400) );
  AOI21_X1 U12957 ( .B1(n10603), .B2(n13159), .A(n10400), .ZN(n10401) );
  OAI21_X1 U12958 ( .B1(n10402), .B2(n14664), .A(n10401), .ZN(P2_U3202) );
  XNOR2_X1 U12959 ( .A(n10404), .B(n10403), .ZN(n10418) );
  INV_X1 U12960 ( .A(n10405), .ZN(n10406) );
  AOI21_X1 U12961 ( .B1(n10408), .B2(n10407), .A(n10406), .ZN(n10410) );
  AOI22_X1 U12962 ( .A1(n14943), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10409) );
  OAI21_X1 U12963 ( .B1(n10410), .B2(n12623), .A(n10409), .ZN(n10415) );
  NAND2_X1 U12964 ( .A1(n10411), .A2(n10880), .ZN(n10412) );
  AOI21_X1 U12965 ( .B1(n10413), .B2(n10412), .A(n14959), .ZN(n10414) );
  AOI211_X1 U12966 ( .C1(n14343), .C2(n10416), .A(n10415), .B(n10414), .ZN(
        n10417) );
  OAI21_X1 U12967 ( .B1(n14939), .B2(n10418), .A(n10417), .ZN(P3_U3183) );
  NAND2_X1 U12968 ( .A1(n13198), .A2(n10760), .ZN(n10510) );
  XNOR2_X1 U12969 ( .A(n10509), .B(n10510), .ZN(n10507) );
  XOR2_X1 U12970 ( .A(n10506), .B(n10507), .Z(n10428) );
  NAND2_X1 U12971 ( .A1(n13197), .A2(n13167), .ZN(n10422) );
  NAND2_X1 U12972 ( .A1(n13199), .A2(n13166), .ZN(n10421) );
  NAND2_X1 U12973 ( .A1(n10422), .A2(n10421), .ZN(n10578) );
  INV_X1 U12974 ( .A(n10423), .ZN(n10424) );
  AOI21_X1 U12975 ( .B1(n14386), .B2(n10578), .A(n10424), .ZN(n10426) );
  NAND2_X1 U12976 ( .A1(n14815), .A2(n14669), .ZN(n10425) );
  OAI211_X1 U12977 ( .C1(n14672), .C2(n10583), .A(n10426), .B(n10425), .ZN(
        n10427) );
  AOI21_X1 U12978 ( .B1(n10428), .B2(n14384), .A(n10427), .ZN(n10429) );
  INV_X1 U12979 ( .A(n10429), .ZN(P2_U3211) );
  INV_X1 U12980 ( .A(n10430), .ZN(n10433) );
  INV_X1 U12981 ( .A(n11751), .ZN(n11761) );
  OAI222_X1 U12982 ( .A1(n13593), .A2(n10431), .B1(n13587), .B2(n10433), .C1(
        n11761), .C2(P2_U3088), .ZN(P2_U3313) );
  OAI222_X1 U12983 ( .A1(P1_U3086), .A2(n11141), .B1(n14183), .B2(n10433), 
        .C1(n10432), .C2(n14180), .ZN(P1_U3341) );
  MUX2_X1 U12984 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12601), .Z(n11405) );
  XNOR2_X1 U12985 ( .A(n11405), .B(n11406), .ZN(n11403) );
  NAND2_X1 U12986 ( .A1(n10435), .A2(n10434), .ZN(n10440) );
  INV_X1 U12987 ( .A(n10436), .ZN(n10438) );
  NAND2_X1 U12988 ( .A1(n10438), .A2(n10437), .ZN(n10439) );
  NAND2_X1 U12989 ( .A1(n10440), .A2(n10439), .ZN(n11404) );
  XOR2_X1 U12990 ( .A(n11403), .B(n11404), .Z(n10454) );
  INV_X1 U12991 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15009) );
  MUX2_X1 U12992 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n15009), .S(n11406), .Z(
        n11390) );
  XNOR2_X1 U12993 ( .A(n11391), .B(n11390), .ZN(n10444) );
  NAND2_X1 U12994 ( .A1(n14954), .A2(n10444), .ZN(n10445) );
  NAND2_X1 U12995 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n11036) );
  OAI211_X1 U12996 ( .C1(n14201), .C2(n14975), .A(n10445), .B(n11036), .ZN(
        n10452) );
  INV_X1 U12997 ( .A(n10448), .ZN(n10446) );
  INV_X1 U12998 ( .A(n10447), .ZN(n10449) );
  NAND3_X1 U12999 ( .A1(n6631), .A2(n10449), .A3(n10448), .ZN(n10450) );
  AOI21_X1 U13000 ( .B1(n11379), .B2(n10450), .A(n14959), .ZN(n10451) );
  AOI211_X1 U13001 ( .C1(n14343), .C2(n11406), .A(n10452), .B(n10451), .ZN(
        n10453) );
  OAI21_X1 U13002 ( .B1(n10454), .B2(n14939), .A(n10453), .ZN(P3_U3186) );
  OAI222_X1 U13003 ( .A1(n13067), .A2(n10456), .B1(n13059), .B2(n15090), .C1(
        P3_U3151), .C2(n10455), .ZN(P3_U3275) );
  NAND2_X1 U13004 ( .A1(n14529), .A2(n13753), .ZN(n10457) );
  NAND2_X1 U13005 ( .A1(n10674), .A2(n14543), .ZN(n10459) );
  NAND2_X1 U13006 ( .A1(n10460), .A2(n10459), .ZN(n10691) );
  XNOR2_X1 U13007 ( .A(n10691), .B(n10689), .ZN(n10505) );
  INV_X1 U13008 ( .A(n10461), .ZN(n10463) );
  NAND2_X1 U13009 ( .A1(n10465), .A2(n10689), .ZN(n10687) );
  OAI21_X1 U13010 ( .B1(n10465), .B2(n10689), .A(n10687), .ZN(n10503) );
  OAI211_X1 U13011 ( .C1(n10685), .C2(n10466), .A(n14556), .B(n10701), .ZN(
        n10501) );
  AOI22_X1 U13012 ( .A1(n14033), .A2(n13753), .B1(n13751), .B2(n14055), .ZN(
        n10497) );
  OAI211_X1 U13013 ( .C1(n10685), .C2(n14640), .A(n10501), .B(n10497), .ZN(
        n10467) );
  AOI21_X1 U13014 ( .B1(n10503), .B2(n14644), .A(n10467), .ZN(n10468) );
  OAI21_X1 U13015 ( .B1(n14580), .B2(n10505), .A(n10468), .ZN(n10471) );
  NAND2_X1 U13016 ( .A1(n10471), .A2(n14657), .ZN(n10469) );
  OAI21_X1 U13017 ( .B1(n14657), .B2(n10470), .A(n10469), .ZN(P1_U3533) );
  NAND2_X1 U13018 ( .A1(n10471), .A2(n14646), .ZN(n10472) );
  OAI21_X1 U13019 ( .B1(n14646), .B2(n9185), .A(n10472), .ZN(P1_U3474) );
  NAND2_X1 U13020 ( .A1(n13862), .A2(n10473), .ZN(n10476) );
  INV_X2 U13021 ( .A(n14576), .ZN(n14578) );
  XNOR2_X1 U13022 ( .A(n10478), .B(n10477), .ZN(n14597) );
  INV_X1 U13023 ( .A(n14545), .ZN(n14593) );
  NAND2_X1 U13024 ( .A1(n14597), .A2(n14593), .ZN(n10485) );
  OAI21_X1 U13025 ( .B1(n10233), .B2(n10480), .A(n10479), .ZN(n10483) );
  OR2_X1 U13026 ( .A1(n14563), .A2(n14542), .ZN(n10482) );
  NAND2_X1 U13027 ( .A1(n13754), .A2(n14055), .ZN(n10481) );
  NAND2_X1 U13028 ( .A1(n10482), .A2(n10481), .ZN(n12028) );
  AOI21_X1 U13029 ( .B1(n10483), .B2(n14549), .A(n12028), .ZN(n10484) );
  AND2_X1 U13030 ( .A1(n10485), .A2(n10484), .ZN(n14599) );
  NOR2_X1 U13031 ( .A1(n14578), .A2(n10494), .ZN(n14559) );
  OAI211_X1 U13032 ( .C1(n14595), .C2(n6491), .A(n14556), .B(n14553), .ZN(
        n14594) );
  INV_X1 U13033 ( .A(n10486), .ZN(n10487) );
  OAI22_X1 U13034 ( .A1(n14576), .A2(n9778), .B1(n10488), .B2(n14526), .ZN(
        n10489) );
  AOI21_X1 U13035 ( .B1(n14550), .B2(n10490), .A(n10489), .ZN(n10491) );
  OAI21_X1 U13036 ( .B1(n13947), .B2(n14594), .A(n10491), .ZN(n10492) );
  AOI21_X1 U13037 ( .B1(n14559), .B2(n14597), .A(n10492), .ZN(n10493) );
  OAI21_X1 U13038 ( .B1(n14578), .B2(n14599), .A(n10493), .ZN(P1_U3291) );
  AND2_X1 U13039 ( .A1(n14576), .A2(n14549), .ZN(n14570) );
  INV_X1 U13040 ( .A(n14570), .ZN(n13995) );
  NAND2_X1 U13041 ( .A1(n14545), .A2(n10494), .ZN(n10495) );
  NOR2_X1 U13042 ( .A1(n14576), .A2(n9184), .ZN(n10499) );
  INV_X1 U13043 ( .A(n10648), .ZN(n10496) );
  OAI22_X1 U13044 ( .A1(n14578), .A2(n10497), .B1(n10496), .B2(n14526), .ZN(
        n10498) );
  AOI211_X1 U13045 ( .C1(n14550), .C2(n10692), .A(n10499), .B(n10498), .ZN(
        n10500) );
  OAI21_X1 U13046 ( .B1(n13947), .B2(n10501), .A(n10500), .ZN(n10502) );
  AOI21_X1 U13047 ( .B1(n14571), .B2(n10503), .A(n10502), .ZN(n10504) );
  OAI21_X1 U13048 ( .B1(n10505), .B2(n13995), .A(n10504), .ZN(P1_U3288) );
  XNOR2_X1 U13049 ( .A(n10665), .B(n11963), .ZN(n10525) );
  NAND2_X1 U13050 ( .A1(n13197), .A2(n13412), .ZN(n10523) );
  XNOR2_X1 U13051 ( .A(n10525), .B(n10523), .ZN(n10521) );
  INV_X1 U13052 ( .A(n10507), .ZN(n10508) );
  INV_X1 U13053 ( .A(n10509), .ZN(n10512) );
  INV_X1 U13054 ( .A(n10510), .ZN(n10511) );
  XOR2_X1 U13055 ( .A(n10521), .B(n10522), .Z(n10519) );
  NAND2_X1 U13056 ( .A1(n10665), .A2(n14669), .ZN(n10517) );
  NAND2_X1 U13057 ( .A1(n13196), .A2(n13167), .ZN(n10514) );
  NAND2_X1 U13058 ( .A1(n13198), .A2(n13166), .ZN(n10513) );
  NAND2_X1 U13059 ( .A1(n10514), .A2(n10513), .ZN(n10775) );
  AOI21_X1 U13060 ( .B1(n14386), .B2(n10775), .A(n10515), .ZN(n10516) );
  OAI211_X1 U13061 ( .C1(n14672), .C2(n10770), .A(n10517), .B(n10516), .ZN(
        n10518) );
  AOI21_X1 U13062 ( .B1(n10519), .B2(n14384), .A(n10518), .ZN(n10520) );
  INV_X1 U13063 ( .A(n10520), .ZN(P2_U3185) );
  INV_X1 U13064 ( .A(n10523), .ZN(n10524) );
  NAND2_X1 U13065 ( .A1(n10525), .A2(n10524), .ZN(n10526) );
  NAND2_X1 U13066 ( .A1(n10527), .A2(n10526), .ZN(n10757) );
  XNOR2_X1 U13067 ( .A(n10790), .B(n11963), .ZN(n10758) );
  NAND2_X1 U13068 ( .A1(n13196), .A2(n13412), .ZN(n10756) );
  XNOR2_X1 U13069 ( .A(n10758), .B(n10756), .ZN(n10528) );
  XNOR2_X1 U13070 ( .A(n10757), .B(n10528), .ZN(n10533) );
  INV_X1 U13071 ( .A(n13197), .ZN(n10660) );
  INV_X1 U13072 ( .A(n13195), .ZN(n10886) );
  OAI22_X1 U13073 ( .A1(n10660), .A2(n13142), .B1(n10886), .B2(n13144), .ZN(
        n10663) );
  AOI21_X1 U13074 ( .B1(n14386), .B2(n10663), .A(n10529), .ZN(n10530) );
  OAI21_X1 U13075 ( .B1(n14672), .B2(n10787), .A(n10530), .ZN(n10531) );
  AOI21_X1 U13076 ( .B1(n10790), .B2(n14669), .A(n10531), .ZN(n10532) );
  OAI21_X1 U13077 ( .B1(n10533), .B2(n14664), .A(n10532), .ZN(P2_U3193) );
  INV_X1 U13078 ( .A(n10534), .ZN(n10537) );
  INV_X1 U13079 ( .A(n14765), .ZN(n11763) );
  OAI222_X1 U13080 ( .A1(n13593), .A2(n10535), .B1(n13587), .B2(n10537), .C1(
        n11763), .C2(P2_U3088), .ZN(P2_U3312) );
  INV_X1 U13081 ( .A(n11142), .ZN(n14507) );
  OAI222_X1 U13082 ( .A1(P1_U3086), .A2(n14507), .B1(n14183), .B2(n10537), 
        .C1(n10536), .C2(n14180), .ZN(P1_U3340) );
  INV_X1 U13083 ( .A(SI_21_), .ZN(n15124) );
  OAI222_X1 U13084 ( .A1(n13067), .A2(n10539), .B1(n13059), .B2(n15124), .C1(
        P3_U3151), .C2(n10538), .ZN(P3_U3274) );
  OR2_X1 U13085 ( .A1(n10843), .A2(n13201), .ZN(n10540) );
  NAND2_X1 U13086 ( .A1(n10541), .A2(n10540), .ZN(n10599) );
  NAND2_X1 U13087 ( .A1(n10599), .A2(n10608), .ZN(n10598) );
  NAND2_X1 U13088 ( .A1(n10598), .A2(n10542), .ZN(n10568) );
  INV_X1 U13089 ( .A(n10553), .ZN(n10549) );
  XNOR2_X1 U13090 ( .A(n10568), .B(n10549), .ZN(n14811) );
  NAND2_X1 U13091 ( .A1(n10179), .A2(n10543), .ZN(n10544) );
  INV_X1 U13092 ( .A(n10608), .ZN(n10547) );
  NAND2_X1 U13093 ( .A1(n10843), .A2(n10545), .ZN(n10607) );
  NAND2_X1 U13094 ( .A1(n10609), .A2(n10607), .ZN(n10546) );
  NAND2_X1 U13095 ( .A1(n10547), .A2(n10546), .ZN(n10551) );
  NAND2_X1 U13096 ( .A1(n14802), .A2(n10548), .ZN(n10552) );
  NAND2_X1 U13097 ( .A1(n10551), .A2(n10552), .ZN(n10550) );
  NAND3_X1 U13098 ( .A1(n10551), .A2(n10553), .A3(n10552), .ZN(n10554) );
  AOI21_X1 U13099 ( .B1(n10575), .B2(n10554), .A(n13430), .ZN(n10556) );
  NOR2_X1 U13100 ( .A1(n10556), .A2(n10555), .ZN(n14809) );
  MUX2_X1 U13101 ( .A(n10557), .B(n14809), .S(n13432), .Z(n10566) );
  INV_X1 U13102 ( .A(n10601), .ZN(n10559) );
  INV_X1 U13103 ( .A(n10582), .ZN(n10558) );
  AOI211_X1 U13104 ( .C1(n14808), .C2(n10559), .A(n13412), .B(n10558), .ZN(
        n14807) );
  AND2_X1 U13105 ( .A1(n10561), .A2(n10560), .ZN(n10562) );
  OAI22_X1 U13106 ( .A1(n13443), .A2(n10570), .B1(n13385), .B2(n10563), .ZN(
        n10564) );
  AOI21_X1 U13107 ( .B1(n14807), .B2(n13455), .A(n10564), .ZN(n10565) );
  OAI211_X1 U13108 ( .C1(n14811), .C2(n13449), .A(n10566), .B(n10565), .ZN(
        P2_U3260) );
  NAND2_X1 U13109 ( .A1(n14808), .A2(n13199), .ZN(n10567) );
  NAND2_X1 U13110 ( .A1(n10568), .A2(n10567), .ZN(n10572) );
  NAND2_X1 U13111 ( .A1(n10570), .A2(n10569), .ZN(n10571) );
  NAND2_X1 U13112 ( .A1(n10572), .A2(n10571), .ZN(n10573) );
  OAI21_X1 U13113 ( .B1(n10574), .B2(n6994), .A(n10652), .ZN(n14818) );
  NAND3_X1 U13114 ( .A1(n6994), .A2(n10576), .A3(n10575), .ZN(n10577) );
  AOI21_X1 U13115 ( .B1(n10658), .B2(n10577), .A(n13430), .ZN(n10579) );
  OR2_X1 U13116 ( .A1(n10579), .A2(n10578), .ZN(n14821) );
  INV_X1 U13117 ( .A(n14821), .ZN(n10581) );
  MUX2_X1 U13118 ( .A(n10581), .B(n10580), .S(n13453), .Z(n10587) );
  AOI211_X1 U13119 ( .C1(n14815), .C2(n10582), .A(n13412), .B(n10769), .ZN(
        n14814) );
  INV_X1 U13120 ( .A(n14815), .ZN(n10584) );
  OAI22_X1 U13121 ( .A1(n13443), .A2(n10584), .B1(n13385), .B2(n10583), .ZN(
        n10585) );
  AOI21_X1 U13122 ( .B1(n14814), .B2(n13455), .A(n10585), .ZN(n10586) );
  OAI211_X1 U13123 ( .C1(n13449), .C2(n14818), .A(n10587), .B(n10586), .ZN(
        P2_U3259) );
  INV_X1 U13124 ( .A(n13361), .ZN(n11197) );
  AOI22_X1 U13125 ( .A1(n11197), .A2(n10589), .B1(n13455), .B2(n10588), .ZN(
        n10593) );
  OAI22_X1 U13126 ( .A1(n11334), .A2(n9847), .B1(n10590), .B2(n13385), .ZN(
        n10591) );
  AOI21_X1 U13127 ( .B1(n13460), .B2(n10078), .A(n10591), .ZN(n10592) );
  OAI211_X1 U13128 ( .C1(n13453), .C2(n10594), .A(n10593), .B(n10592), .ZN(
        P2_U3264) );
  INV_X1 U13129 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10597) );
  NAND2_X1 U13130 ( .A1(n10595), .A2(n14835), .ZN(n10596) );
  OAI21_X1 U13131 ( .B1(n14835), .B2(n10597), .A(n10596), .ZN(P2_U3433) );
  OAI21_X1 U13132 ( .B1(n10599), .B2(n10608), .A(n10598), .ZN(n10600) );
  INV_X1 U13133 ( .A(n10600), .ZN(n14805) );
  AOI211_X1 U13134 ( .C1(n14802), .C2(n10602), .A(n13412), .B(n10601), .ZN(
        n14801) );
  INV_X1 U13135 ( .A(n10603), .ZN(n10604) );
  OAI22_X1 U13136 ( .A1(n13443), .A2(n10605), .B1(n13385), .B2(n10604), .ZN(
        n10606) );
  AOI21_X1 U13137 ( .B1(n13455), .B2(n14801), .A(n10606), .ZN(n10615) );
  NAND3_X1 U13138 ( .A1(n10609), .A2(n10608), .A3(n10607), .ZN(n10610) );
  AOI21_X1 U13139 ( .B1(n10551), .B2(n10610), .A(n13430), .ZN(n10612) );
  NOR2_X1 U13140 ( .A1(n10612), .A2(n10611), .ZN(n14804) );
  MUX2_X1 U13141 ( .A(n10613), .B(n14804), .S(n13432), .Z(n10614) );
  OAI211_X1 U13142 ( .C1(n13449), .C2(n14805), .A(n10615), .B(n10614), .ZN(
        P2_U3261) );
  NOR2_X1 U13143 ( .A1(n12222), .A2(n12226), .ZN(n12199) );
  INV_X1 U13144 ( .A(n12491), .ZN(n12468) );
  INV_X1 U13145 ( .A(n12485), .ZN(n12497) );
  AOI22_X1 U13146 ( .A1(n12468), .A2(n12521), .B1(n12497), .B2(n10811), .ZN(
        n10617) );
  NAND2_X1 U13147 ( .A1(n12495), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10806) );
  NAND2_X1 U13148 ( .A1(n10806), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10616) );
  OAI211_X1 U13149 ( .C1(n12199), .C2(n12499), .A(n10617), .B(n10616), .ZN(
        P3_U3172) );
  AND2_X1 U13150 ( .A1(n10618), .A2(n12903), .ZN(n10619) );
  OR2_X1 U13151 ( .A1(n12199), .A2(n10619), .ZN(n10621) );
  NAND2_X1 U13152 ( .A1(n12521), .A2(n12846), .ZN(n10620) );
  NAND2_X1 U13153 ( .A1(n10621), .A2(n10620), .ZN(n10809) );
  INV_X1 U13154 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10622) );
  OAI22_X1 U13155 ( .A1(n13053), .A2(n12219), .B1(n10622), .B2(n15004), .ZN(
        n10623) );
  AOI21_X1 U13156 ( .B1(n10809), .B2(n15004), .A(n10623), .ZN(n10624) );
  INV_X1 U13157 ( .A(n10624), .ZN(P3_U3390) );
  NAND2_X1 U13158 ( .A1(n12522), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n10625) );
  OAI21_X1 U13159 ( .B1(n12652), .B2(n12522), .A(n10625), .ZN(P3_U3519) );
  INV_X1 U13160 ( .A(n10626), .ZN(n10628) );
  AND2_X1 U13161 ( .A1(n12147), .A2(n13753), .ZN(n10631) );
  AOI21_X1 U13162 ( .B1(n10674), .B2(n10630), .A(n10631), .ZN(n10634) );
  INV_X1 U13163 ( .A(n10634), .ZN(n10632) );
  OAI22_X1 U13164 ( .A1(n14529), .A2(n12107), .B1(n14543), .B2(n12106), .ZN(
        n10633) );
  XNOR2_X1 U13165 ( .A(n10633), .B(n12141), .ZN(n10673) );
  NAND2_X1 U13166 ( .A1(n10692), .A2(n12146), .ZN(n10638) );
  NAND2_X1 U13167 ( .A1(n13752), .A2(n10630), .ZN(n10637) );
  NAND2_X1 U13168 ( .A1(n10638), .A2(n10637), .ZN(n10639) );
  XNOR2_X1 U13169 ( .A(n10639), .B(n12141), .ZN(n10643) );
  NAND2_X1 U13170 ( .A1(n10692), .A2(n10630), .ZN(n10641) );
  NAND2_X1 U13171 ( .A1(n12147), .A2(n13752), .ZN(n10640) );
  NAND2_X1 U13172 ( .A1(n10641), .A2(n10640), .ZN(n10642) );
  NAND2_X1 U13173 ( .A1(n10643), .A2(n10642), .ZN(n11012) );
  NAND2_X1 U13174 ( .A1(n6626), .A2(n11012), .ZN(n10644) );
  XNOR2_X1 U13175 ( .A(n6625), .B(n10644), .ZN(n10650) );
  NAND2_X1 U13176 ( .A1(n13729), .A2(n13751), .ZN(n10645) );
  NAND2_X1 U13177 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n13796) );
  OAI211_X1 U13178 ( .C1(n14543), .C2(n14419), .A(n10645), .B(n13796), .ZN(
        n10647) );
  NOR2_X1 U13179 ( .A1(n13737), .A2(n10685), .ZN(n10646) );
  AOI211_X1 U13180 ( .C1(n13733), .C2(n10648), .A(n10647), .B(n10646), .ZN(
        n10649) );
  OAI21_X1 U13181 ( .B1(n10650), .B2(n14426), .A(n10649), .ZN(P1_U3227) );
  NAND2_X1 U13182 ( .A1(n14815), .A2(n13198), .ZN(n10651) );
  OR2_X1 U13183 ( .A1(n10665), .A2(n13197), .ZN(n10653) );
  NAND2_X1 U13184 ( .A1(n10665), .A2(n13197), .ZN(n10654) );
  NAND2_X1 U13185 ( .A1(n10655), .A2(n10654), .ZN(n10724) );
  XNOR2_X1 U13186 ( .A(n10724), .B(n10723), .ZN(n10794) );
  INV_X1 U13187 ( .A(n13198), .ZN(n10656) );
  NAND2_X1 U13188 ( .A1(n14815), .A2(n10656), .ZN(n10657) );
  OR2_X1 U13189 ( .A1(n10665), .A2(n10660), .ZN(n10659) );
  NAND2_X1 U13190 ( .A1(n10665), .A2(n10660), .ZN(n10661) );
  NAND2_X1 U13191 ( .A1(n10662), .A2(n10661), .ZN(n10728) );
  INV_X1 U13192 ( .A(n10723), .ZN(n10727) );
  XNOR2_X1 U13193 ( .A(n10728), .B(n10727), .ZN(n10664) );
  AOI21_X1 U13194 ( .B1(n10664), .B2(n13437), .A(n10663), .ZN(n10797) );
  INV_X1 U13195 ( .A(n10665), .ZN(n14826) );
  NAND2_X1 U13196 ( .A1(n14826), .A2(n10769), .ZN(n10768) );
  NAND2_X1 U13197 ( .A1(n10768), .A2(n10790), .ZN(n10666) );
  NAND2_X1 U13198 ( .A1(n10666), .A2(n11850), .ZN(n10667) );
  NOR2_X1 U13199 ( .A1(n10734), .A2(n10667), .ZN(n10791) );
  AOI21_X1 U13200 ( .B1(n14816), .B2(n10790), .A(n10791), .ZN(n10668) );
  OAI211_X1 U13201 ( .C1(n10794), .C2(n14812), .A(n10797), .B(n10668), .ZN(
        n10670) );
  NAND2_X1 U13202 ( .A1(n10670), .A2(n14855), .ZN(n10669) );
  OAI21_X1 U13203 ( .B1(n14855), .B2(n9984), .A(n10669), .ZN(P2_U3507) );
  NAND2_X1 U13204 ( .A1(n10670), .A2(n14835), .ZN(n10671) );
  OAI21_X1 U13205 ( .B1(n14835), .B2(n7687), .A(n10671), .ZN(P2_U3454) );
  XOR2_X1 U13206 ( .A(n10673), .B(n10672), .Z(n10679) );
  NAND2_X1 U13207 ( .A1(n14432), .A2(n10674), .ZN(n10677) );
  AND2_X1 U13208 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14493) );
  AOI21_X1 U13209 ( .B1(n14414), .B2(n10675), .A(n14493), .ZN(n10676) );
  OAI211_X1 U13210 ( .C1(n14436), .C2(n14527), .A(n10677), .B(n10676), .ZN(
        n10678) );
  AOI21_X1 U13211 ( .B1(n10679), .B2(n14412), .A(n10678), .ZN(n10680) );
  INV_X1 U13212 ( .A(n10680), .ZN(P1_U3230) );
  INV_X1 U13213 ( .A(n13236), .ZN(n11766) );
  INV_X1 U13214 ( .A(n10681), .ZN(n10684) );
  OAI222_X1 U13215 ( .A1(P2_U3088), .A2(n11766), .B1(n13587), .B2(n10684), 
        .C1(n10682), .C2(n13593), .ZN(P2_U3311) );
  INV_X1 U13216 ( .A(n11145), .ZN(n11271) );
  OAI222_X1 U13217 ( .A1(P1_U3086), .A2(n11271), .B1(n14183), .B2(n10684), 
        .C1(n10683), .C2(n14180), .ZN(P1_U3339) );
  NAND2_X1 U13218 ( .A1(n10685), .A2(n13711), .ZN(n10686) );
  NAND2_X1 U13219 ( .A1(n10687), .A2(n10686), .ZN(n10688) );
  INV_X1 U13220 ( .A(n10902), .ZN(n10695) );
  NAND2_X1 U13221 ( .A1(n10688), .A2(n10695), .ZN(n10919) );
  OAI21_X1 U13222 ( .B1(n10688), .B2(n10695), .A(n10919), .ZN(n10696) );
  INV_X1 U13223 ( .A(n10696), .ZN(n14610) );
  INV_X1 U13224 ( .A(n14559), .ZN(n11010) );
  NAND2_X1 U13225 ( .A1(n10691), .A2(n10690), .ZN(n10694) );
  NAND2_X1 U13226 ( .A1(n10692), .A2(n13711), .ZN(n10693) );
  NAND2_X1 U13227 ( .A1(n10694), .A2(n10693), .ZN(n10903) );
  XNOR2_X1 U13228 ( .A(n10903), .B(n10695), .ZN(n10699) );
  NAND2_X1 U13229 ( .A1(n10696), .A2(n14593), .ZN(n10698) );
  AOI22_X1 U13230 ( .A1(n14033), .A2(n13752), .B1(n13750), .B2(n14055), .ZN(
        n10697) );
  OAI211_X1 U13231 ( .C1(n14580), .C2(n10699), .A(n10698), .B(n10697), .ZN(
        n14612) );
  MUX2_X1 U13232 ( .A(n14612), .B(P1_REG2_REG_6__SCAN_IN), .S(n14578), .Z(
        n10700) );
  INV_X1 U13233 ( .A(n10700), .ZN(n10705) );
  AOI211_X1 U13234 ( .C1(n14607), .C2(n10701), .A(n14058), .B(n10936), .ZN(
        n14605) );
  INV_X1 U13235 ( .A(n14607), .ZN(n10702) );
  OAI22_X1 U13236 ( .A1(n10702), .A2(n14530), .B1(n13713), .B2(n14526), .ZN(
        n10703) );
  AOI21_X1 U13237 ( .B1(n14605), .B2(n14558), .A(n10703), .ZN(n10704) );
  OAI211_X1 U13238 ( .C1(n14610), .C2(n11010), .A(n10705), .B(n10704), .ZN(
        P1_U3287) );
  NAND2_X1 U13239 ( .A1(n10707), .A2(n10706), .ZN(n10710) );
  NAND2_X1 U13240 ( .A1(n13054), .A2(n10708), .ZN(n10709) );
  NAND2_X1 U13241 ( .A1(n10710), .A2(n10709), .ZN(n10711) );
  NOR2_X1 U13242 ( .A1(n12941), .A2(n12359), .ZN(n10713) );
  MUX2_X1 U13243 ( .A(n10809), .B(P3_REG2_REG_0__SCAN_IN), .S(n12786), .Z(
        n10718) );
  OAI22_X1 U13244 ( .A1(n12870), .A2(n12219), .B1(n12910), .B2(n10716), .ZN(
        n10717) );
  OR2_X1 U13245 ( .A1(n10718), .A2(n10717), .ZN(P3_U3233) );
  NOR2_X1 U13246 ( .A1(n13059), .A2(SI_22_), .ZN(n10719) );
  AOI21_X1 U13247 ( .B1(n12218), .B2(P3_STATE_REG_SCAN_IN), .A(n10719), .ZN(
        n10720) );
  OAI21_X1 U13248 ( .B1(n10721), .B2(n13067), .A(n10720), .ZN(n10722) );
  INV_X1 U13249 ( .A(n10722), .ZN(P3_U3273) );
  NAND2_X1 U13250 ( .A1(n10724), .A2(n10723), .ZN(n10726) );
  NAND2_X1 U13251 ( .A1(n10790), .A2(n13196), .ZN(n10725) );
  NAND2_X1 U13252 ( .A1(n10726), .A2(n10725), .ZN(n10883) );
  XNOR2_X1 U13253 ( .A(n10883), .B(n10731), .ZN(n10836) );
  NAND2_X1 U13254 ( .A1(n10790), .A2(n10729), .ZN(n10730) );
  INV_X1 U13255 ( .A(n10731), .ZN(n10882) );
  XNOR2_X1 U13256 ( .A(n10889), .B(n10882), .ZN(n10732) );
  AOI22_X1 U13257 ( .A1(n13166), .A2(n13196), .B1(n13194), .B2(n13167), .ZN(
        n10762) );
  OAI21_X1 U13258 ( .B1(n10732), .B2(n13430), .A(n10762), .ZN(n10733) );
  AOI21_X1 U13259 ( .B1(n10836), .B2(n14823), .A(n10733), .ZN(n10838) );
  INV_X1 U13260 ( .A(n10734), .ZN(n10736) );
  INV_X1 U13261 ( .A(n10887), .ZN(n10737) );
  INV_X1 U13262 ( .A(n10894), .ZN(n10735) );
  AOI211_X1 U13263 ( .C1(n10887), .C2(n10736), .A(n13412), .B(n10735), .ZN(
        n10837) );
  NOR2_X1 U13264 ( .A1(n10737), .A2(n13443), .ZN(n10740) );
  OAI22_X1 U13265 ( .A1(n11334), .A2(n10738), .B1(n10761), .B2(n13385), .ZN(
        n10739) );
  AOI211_X1 U13266 ( .C1(n10837), .C2(n13455), .A(n10740), .B(n10739), .ZN(
        n10742) );
  NAND2_X1 U13267 ( .A1(n10836), .A2(n11197), .ZN(n10741) );
  OAI211_X1 U13268 ( .C1(n10838), .C2(n13453), .A(n10742), .B(n10741), .ZN(
        P2_U3256) );
  NAND2_X1 U13269 ( .A1(n10746), .A2(n10744), .ZN(n10802) );
  AOI211_X1 U13270 ( .C1(n10745), .C2(n12379), .A(n10872), .B(n10802), .ZN(
        n10800) );
  INV_X1 U13271 ( .A(n10746), .ZN(n10747) );
  NOR2_X1 U13272 ( .A1(n10800), .A2(n10747), .ZN(n10750) );
  XNOR2_X1 U13273 ( .A(n10748), .B(n12520), .ZN(n10749) );
  XNOR2_X1 U13274 ( .A(n10750), .B(n10749), .ZN(n10755) );
  AOI22_X1 U13275 ( .A1(n12493), .A2(n12521), .B1(n12468), .B2(n12519), .ZN(
        n10751) );
  OAI21_X1 U13276 ( .B1(n10752), .B2(n12485), .A(n10751), .ZN(n10753) );
  AOI21_X1 U13277 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10806), .A(n10753), .ZN(
        n10754) );
  OAI21_X1 U13278 ( .B1(n10755), .B2(n12499), .A(n10754), .ZN(P3_U3177) );
  INV_X1 U13279 ( .A(n10758), .ZN(n10759) );
  XNOR2_X1 U13280 ( .A(n10887), .B(n11963), .ZN(n10852) );
  NAND2_X1 U13281 ( .A1(n13195), .A2(n13412), .ZN(n10853) );
  XNOR2_X1 U13282 ( .A(n10852), .B(n10853), .ZN(n10850) );
  XOR2_X1 U13283 ( .A(n10851), .B(n10850), .Z(n10766) );
  NOR2_X1 U13284 ( .A1(n14672), .A2(n10761), .ZN(n10764) );
  INV_X1 U13285 ( .A(n14386), .ZN(n14660) );
  NAND2_X1 U13286 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14732) );
  OAI21_X1 U13287 ( .B1(n14660), .B2(n10762), .A(n14732), .ZN(n10763) );
  AOI211_X1 U13288 ( .C1(n10887), .C2(n14669), .A(n10764), .B(n10763), .ZN(
        n10765) );
  OAI21_X1 U13289 ( .B1(n10766), .B2(n14664), .A(n10765), .ZN(P2_U3203) );
  XNOR2_X1 U13290 ( .A(n10767), .B(n10773), .ZN(n14828) );
  INV_X1 U13291 ( .A(n13449), .ZN(n13457) );
  OAI211_X1 U13292 ( .C1(n14826), .C2(n10769), .A(n11850), .B(n10768), .ZN(
        n14824) );
  NOR2_X1 U13293 ( .A1(n14824), .A2(n13391), .ZN(n10772) );
  OAI22_X1 U13294 ( .A1(n14826), .A2(n13443), .B1(n13385), .B2(n10770), .ZN(
        n10771) );
  AOI211_X1 U13295 ( .C1(n14828), .C2(n13457), .A(n10772), .B(n10771), .ZN(
        n10779) );
  XNOR2_X1 U13296 ( .A(n10774), .B(n10773), .ZN(n10776) );
  AOI21_X1 U13297 ( .B1(n10776), .B2(n13437), .A(n10775), .ZN(n14825) );
  MUX2_X1 U13298 ( .A(n10777), .B(n14825), .S(n13432), .Z(n10778) );
  NAND2_X1 U13299 ( .A1(n10779), .A2(n10778), .ZN(P2_U3258) );
  AOI21_X1 U13300 ( .B1(n10781), .B2(n10780), .A(n12499), .ZN(n10782) );
  NAND2_X1 U13301 ( .A1(n10782), .A2(n11033), .ZN(n10786) );
  OAI22_X1 U13302 ( .A1(n12479), .A2(n10875), .B1(n10969), .B2(n12485), .ZN(
        n10783) );
  AOI211_X1 U13303 ( .C1(n12468), .C2(n12518), .A(n10784), .B(n10783), .ZN(
        n10785) );
  OAI211_X1 U13304 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12495), .A(n10786), .B(
        n10785), .ZN(P3_U3158) );
  OAI22_X1 U13305 ( .A1(n11334), .A2(n10788), .B1(n10787), .B2(n13385), .ZN(
        n10789) );
  AOI21_X1 U13306 ( .B1(n10790), .B2(n13460), .A(n10789), .ZN(n10793) );
  NAND2_X1 U13307 ( .A1(n10791), .A2(n13455), .ZN(n10792) );
  OAI211_X1 U13308 ( .C1(n10794), .C2(n13449), .A(n10793), .B(n10792), .ZN(
        n10795) );
  INV_X1 U13309 ( .A(n10795), .ZN(n10796) );
  OAI21_X1 U13310 ( .B1(n13453), .B2(n10797), .A(n10796), .ZN(P2_U3257) );
  INV_X1 U13311 ( .A(n12202), .ZN(n10799) );
  NOR3_X1 U13312 ( .A1(n10799), .A2(n12222), .A3(n10798), .ZN(n10801) );
  AOI211_X1 U13313 ( .C1(n10872), .C2(n10802), .A(n10801), .B(n10800), .ZN(
        n10808) );
  AOI22_X1 U13314 ( .A1(n12493), .A2(n12523), .B1(n12520), .B2(n12468), .ZN(
        n10803) );
  OAI21_X1 U13315 ( .B1(n10804), .B2(n12485), .A(n10803), .ZN(n10805) );
  AOI21_X1 U13316 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(n10806), .A(n10805), .ZN(
        n10807) );
  OAI21_X1 U13317 ( .B1(n10808), .B2(n12499), .A(n10807), .ZN(P3_U3162) );
  MUX2_X1 U13318 ( .A(n10809), .B(P3_REG1_REG_0__SCAN_IN), .S(n15014), .Z(
        n10810) );
  AOI21_X1 U13319 ( .B1(n8875), .B2(n10811), .A(n10810), .ZN(n10812) );
  INV_X1 U13320 ( .A(n10812), .ZN(P3_U3459) );
  INV_X1 U13321 ( .A(n10813), .ZN(n10816) );
  INV_X1 U13322 ( .A(n14777), .ZN(n11768) );
  OAI222_X1 U13323 ( .A1(n13593), .A2(n10814), .B1(n13587), .B2(n10816), .C1(
        n11768), .C2(P2_U3088), .ZN(P2_U3310) );
  OAI222_X1 U13324 ( .A1(P1_U3086), .A2(n13817), .B1(n14183), .B2(n10816), 
        .C1(n10815), .C2(n14180), .ZN(P1_U3338) );
  INV_X2 U13325 ( .A(n12786), .ZN(n12813) );
  AND2_X1 U13326 ( .A1(n12221), .A2(n11064), .ZN(n10817) );
  NAND2_X1 U13327 ( .A1(n12813), .A2(n10817), .ZN(n12656) );
  NAND2_X1 U13328 ( .A1(n12667), .A2(n12813), .ZN(n10819) );
  OAI21_X1 U13329 ( .B1(n10821), .B2(n12198), .A(n10820), .ZN(n10822) );
  INV_X1 U13330 ( .A(n10822), .ZN(n10965) );
  INV_X1 U13331 ( .A(n10823), .ZN(n10824) );
  AOI21_X1 U13332 ( .B1(n10824), .B2(n12198), .A(n12903), .ZN(n10828) );
  OAI22_X1 U13333 ( .A1(n10875), .A2(n12906), .B1(n10825), .B2(n12908), .ZN(
        n10826) );
  AOI21_X1 U13334 ( .B1(n10828), .B2(n10827), .A(n10826), .ZN(n10964) );
  MUX2_X1 U13335 ( .A(n10829), .B(n10964), .S(n12813), .Z(n10832) );
  INV_X1 U13336 ( .A(n12910), .ZN(n12868) );
  AOI22_X1 U13337 ( .A1(n12801), .A2(n10830), .B1(n12868), .B2(n8365), .ZN(
        n10831) );
  OAI211_X1 U13338 ( .C1(n12918), .C2(n10965), .A(n10832), .B(n10831), .ZN(
        P3_U3230) );
  INV_X1 U13339 ( .A(SI_23_), .ZN(n10835) );
  NAND2_X1 U13340 ( .A1(n10833), .A2(n13062), .ZN(n10834) );
  OAI211_X1 U13341 ( .C1(n10835), .C2(n13059), .A(n10834), .B(n12369), .ZN(
        P3_U3272) );
  INV_X1 U13342 ( .A(n10836), .ZN(n10840) );
  AOI21_X1 U13343 ( .B1(n14816), .B2(n10887), .A(n10837), .ZN(n10839) );
  OAI211_X1 U13344 ( .C1(n10840), .C2(n14819), .A(n10839), .B(n10838), .ZN(
        n10870) );
  NAND2_X1 U13345 ( .A1(n10870), .A2(n14855), .ZN(n10841) );
  OAI21_X1 U13346 ( .B1(n14855), .B2(n10097), .A(n10841), .ZN(P2_U3508) );
  MUX2_X1 U13347 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10842), .S(n13432), .Z(
        n10847) );
  AOI22_X1 U13348 ( .A1(n13460), .A2(n10843), .B1(n14694), .B2(n13458), .ZN(
        n10844) );
  OAI21_X1 U13349 ( .B1(n13391), .B2(n10845), .A(n10844), .ZN(n10846) );
  AOI211_X1 U13350 ( .C1(n11197), .C2(n10848), .A(n10847), .B(n10846), .ZN(
        n10849) );
  INV_X1 U13351 ( .A(n10849), .ZN(P2_U3262) );
  INV_X1 U13352 ( .A(n11072), .ZN(n14830) );
  INV_X1 U13353 ( .A(n10852), .ZN(n10854) );
  NAND2_X1 U13354 ( .A1(n10854), .A2(n10853), .ZN(n10855) );
  XNOR2_X1 U13355 ( .A(n11072), .B(n11963), .ZN(n10856) );
  AND2_X1 U13356 ( .A1(n13194), .A2(n13412), .ZN(n10857) );
  NAND2_X1 U13357 ( .A1(n10856), .A2(n10857), .ZN(n11241) );
  INV_X1 U13358 ( .A(n10856), .ZN(n10859) );
  INV_X1 U13359 ( .A(n10857), .ZN(n10858) );
  NAND2_X1 U13360 ( .A1(n10859), .A2(n10858), .ZN(n10860) );
  NAND2_X1 U13361 ( .A1(n11241), .A2(n10860), .ZN(n10862) );
  AOI21_X1 U13362 ( .B1(n10861), .B2(n10862), .A(n14664), .ZN(n10864) );
  NAND2_X1 U13363 ( .A1(n10864), .A2(n11245), .ZN(n10869) );
  INV_X1 U13364 ( .A(n10896), .ZN(n10867) );
  AOI22_X1 U13365 ( .A1(n13166), .A2(n13195), .B1(n13193), .B2(n13167), .ZN(
        n10892) );
  OAI21_X1 U13366 ( .B1(n14660), .B2(n10892), .A(n10865), .ZN(n10866) );
  AOI21_X1 U13367 ( .B1(n10867), .B2(n13159), .A(n10866), .ZN(n10868) );
  OAI211_X1 U13368 ( .C1(n14830), .C2(n13162), .A(n10869), .B(n10868), .ZN(
        P2_U3189) );
  NAND2_X1 U13369 ( .A1(n10870), .A2(n14835), .ZN(n10871) );
  OAI21_X1 U13370 ( .B1(n14835), .B2(n7720), .A(n10871), .ZN(P2_U3457) );
  XNOR2_X1 U13371 ( .A(n12222), .B(n12202), .ZN(n14978) );
  INV_X1 U13372 ( .A(n12523), .ZN(n10874) );
  XNOR2_X1 U13373 ( .A(n12202), .B(n10872), .ZN(n10873) );
  OAI222_X1 U13374 ( .A1(n12908), .A2(n10875), .B1(n12906), .B2(n10874), .C1(
        n12903), .C2(n10873), .ZN(n14980) );
  NAND2_X1 U13375 ( .A1(n10876), .A2(n12979), .ZN(n14976) );
  OAI22_X1 U13376 ( .A1(n14976), .A2(n11064), .B1(n12910), .B2(n10877), .ZN(
        n10878) );
  NOR2_X1 U13377 ( .A1(n14980), .A2(n10878), .ZN(n10879) );
  MUX2_X1 U13378 ( .A(n10880), .B(n10879), .S(n12813), .Z(n10881) );
  OAI21_X1 U13379 ( .B1(n12918), .B2(n14978), .A(n10881), .ZN(P3_U3232) );
  NAND2_X1 U13380 ( .A1(n10883), .A2(n10882), .ZN(n10885) );
  NAND2_X1 U13381 ( .A1(n10887), .A2(n13195), .ZN(n10884) );
  NAND2_X1 U13382 ( .A1(n10885), .A2(n10884), .ZN(n11071) );
  XOR2_X1 U13383 ( .A(n11071), .B(n11070), .Z(n14834) );
  INV_X1 U13384 ( .A(n14834), .ZN(n10901) );
  AND2_X1 U13385 ( .A1(n10887), .A2(n10886), .ZN(n10888) );
  INV_X1 U13386 ( .A(n11076), .ZN(n10890) );
  AOI21_X1 U13387 ( .B1(n11070), .B2(n10891), .A(n10890), .ZN(n10893) );
  OAI21_X1 U13388 ( .B1(n10893), .B2(n13430), .A(n10892), .ZN(n14831) );
  NAND2_X1 U13389 ( .A1(n11072), .A2(n10894), .ZN(n10895) );
  NAND3_X1 U13390 ( .A1(n11083), .A2(n11850), .A3(n10895), .ZN(n14829) );
  OAI22_X1 U13391 ( .A1(n11334), .A2(n7737), .B1(n10896), .B2(n13385), .ZN(
        n10897) );
  AOI21_X1 U13392 ( .B1(n11072), .B2(n13460), .A(n10897), .ZN(n10898) );
  OAI21_X1 U13393 ( .B1(n14829), .B2(n13391), .A(n10898), .ZN(n10899) );
  AOI21_X1 U13394 ( .B1(n14831), .B2(n13432), .A(n10899), .ZN(n10900) );
  OAI21_X1 U13395 ( .B1(n13449), .B2(n10901), .A(n10900), .ZN(P2_U3255) );
  NAND2_X1 U13396 ( .A1(n10903), .A2(n10902), .ZN(n10906) );
  INV_X1 U13397 ( .A(n13751), .ZN(n10904) );
  NAND2_X1 U13398 ( .A1(n14607), .A2(n10904), .ZN(n10905) );
  INV_X1 U13399 ( .A(n13750), .ZN(n10908) );
  AND2_X1 U13400 ( .A1(n11021), .A2(n10908), .ZN(n10907) );
  OR2_X1 U13401 ( .A1(n11021), .A2(n10908), .ZN(n10909) );
  INV_X1 U13402 ( .A(n10955), .ZN(n10911) );
  NOR2_X1 U13403 ( .A1(n11200), .A2(n10998), .ZN(n10910) );
  NAND2_X1 U13404 ( .A1(n10997), .A2(n10922), .ZN(n10914) );
  INV_X1 U13405 ( .A(n13748), .ZN(n10912) );
  NAND2_X1 U13406 ( .A1(n11466), .A2(n10912), .ZN(n10913) );
  NAND2_X1 U13407 ( .A1(n10914), .A2(n10913), .ZN(n10915) );
  AOI21_X1 U13408 ( .B1(n10915), .B2(n10924), .A(n14580), .ZN(n10917) );
  NAND2_X1 U13409 ( .A1(n13748), .A2(n14033), .ZN(n11610) );
  INV_X1 U13410 ( .A(n11610), .ZN(n10916) );
  AOI21_X1 U13411 ( .B1(n10917), .B2(n11110), .A(n10916), .ZN(n14639) );
  OR2_X1 U13412 ( .A1(n14607), .A2(n13751), .ZN(n10918) );
  NAND2_X1 U13413 ( .A1(n10919), .A2(n10918), .ZN(n10935) );
  INV_X1 U13414 ( .A(n10942), .ZN(n10934) );
  NAND2_X1 U13415 ( .A1(n10935), .A2(n10934), .ZN(n10933) );
  OR2_X1 U13416 ( .A1(n11021), .A2(n13750), .ZN(n10920) );
  OR2_X1 U13417 ( .A1(n11200), .A2(n13749), .ZN(n10921) );
  OR2_X1 U13418 ( .A1(n11466), .A2(n13748), .ZN(n10923) );
  NAND2_X1 U13419 ( .A1(n10925), .A2(n10924), .ZN(n11115) );
  OAI21_X1 U13420 ( .B1(n10925), .B2(n10924), .A(n11115), .ZN(n14643) );
  INV_X1 U13421 ( .A(n11021), .ZN(n10937) );
  NAND2_X1 U13422 ( .A1(n10937), .A2(n10936), .ZN(n10952) );
  INV_X1 U13423 ( .A(n11466), .ZN(n11004) );
  AOI21_X1 U13424 ( .B1(n11605), .B2(n11003), .A(n14058), .ZN(n10927) );
  NAND2_X1 U13425 ( .A1(n13746), .A2(n14055), .ZN(n11609) );
  INV_X1 U13426 ( .A(n11609), .ZN(n10926) );
  AOI21_X1 U13427 ( .B1(n10927), .B2(n11118), .A(n10926), .ZN(n14638) );
  OAI22_X1 U13428 ( .A1(n14576), .A2(n10928), .B1(n11608), .B2(n14526), .ZN(
        n10929) );
  AOI21_X1 U13429 ( .B1(n11605), .B2(n14550), .A(n10929), .ZN(n10930) );
  OAI21_X1 U13430 ( .B1(n14638), .B2(n13947), .A(n10930), .ZN(n10931) );
  AOI21_X1 U13431 ( .B1(n14643), .B2(n14571), .A(n10931), .ZN(n10932) );
  OAI21_X1 U13432 ( .B1(n14639), .B2(n14578), .A(n10932), .ZN(P1_U3283) );
  OAI21_X1 U13433 ( .B1(n10935), .B2(n10934), .A(n10933), .ZN(n14620) );
  OAI211_X1 U13434 ( .C1(n10937), .C2(n10936), .A(n14556), .B(n10952), .ZN(
        n14616) );
  INV_X1 U13435 ( .A(n14526), .ZN(n14574) );
  INV_X1 U13436 ( .A(n11025), .ZN(n10938) );
  AOI22_X1 U13437 ( .A1(n11021), .A2(n14550), .B1(n14574), .B2(n10938), .ZN(
        n10939) );
  OAI21_X1 U13438 ( .B1(n14616), .B2(n13947), .A(n10939), .ZN(n10948) );
  NAND2_X1 U13439 ( .A1(n14620), .A2(n14593), .ZN(n10945) );
  NAND2_X1 U13440 ( .A1(n13749), .A2(n14055), .ZN(n10941) );
  NAND2_X1 U13441 ( .A1(n13751), .A2(n14033), .ZN(n10940) );
  NAND2_X1 U13442 ( .A1(n10941), .A2(n10940), .ZN(n11028) );
  INV_X1 U13443 ( .A(n11028), .ZN(n14615) );
  XNOR2_X1 U13444 ( .A(n10943), .B(n10942), .ZN(n10944) );
  NAND2_X1 U13445 ( .A1(n10944), .A2(n14549), .ZN(n14617) );
  NAND3_X1 U13446 ( .A1(n10945), .A2(n14615), .A3(n14617), .ZN(n10946) );
  MUX2_X1 U13447 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10946), .S(n14576), .Z(
        n10947) );
  AOI211_X1 U13448 ( .C1(n14559), .C2(n14620), .A(n10948), .B(n10947), .ZN(
        n10949) );
  INV_X1 U13449 ( .A(n10949), .ZN(P1_U3286) );
  OAI21_X1 U13450 ( .B1(n6644), .B2(n10955), .A(n10950), .ZN(n14628) );
  INV_X1 U13451 ( .A(n11200), .ZN(n11209) );
  INV_X1 U13452 ( .A(n10952), .ZN(n10954) );
  INV_X1 U13453 ( .A(n11005), .ZN(n10953) );
  OAI211_X1 U13454 ( .C1(n11209), .C2(n10954), .A(n10953), .B(n14556), .ZN(
        n14624) );
  OAI22_X1 U13455 ( .A1(n14624), .A2(n13947), .B1(n11209), .B2(n14530), .ZN(
        n10962) );
  XNOR2_X1 U13456 ( .A(n10956), .B(n10955), .ZN(n10957) );
  NAND2_X1 U13457 ( .A1(n10957), .A2(n14549), .ZN(n14625) );
  NAND2_X1 U13458 ( .A1(n13748), .A2(n14055), .ZN(n10959) );
  NAND2_X1 U13459 ( .A1(n13750), .A2(n14033), .ZN(n10958) );
  NAND2_X1 U13460 ( .A1(n10959), .A2(n10958), .ZN(n11210) );
  INV_X1 U13461 ( .A(n11210), .ZN(n14623) );
  OAI211_X1 U13462 ( .C1(n14526), .C2(n11212), .A(n14625), .B(n14623), .ZN(
        n10960) );
  MUX2_X1 U13463 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10960), .S(n14576), .Z(
        n10961) );
  AOI211_X1 U13464 ( .C1(n14571), .C2(n14628), .A(n10962), .B(n10961), .ZN(
        n10963) );
  INV_X1 U13465 ( .A(n10963), .ZN(P1_U3285) );
  OAI21_X1 U13466 ( .B1(n14977), .B2(n10965), .A(n10964), .ZN(n10971) );
  INV_X1 U13467 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n10966) );
  OAI22_X1 U13468 ( .A1(n13053), .A2(n10969), .B1(n10966), .B2(n15004), .ZN(
        n10967) );
  AOI21_X1 U13469 ( .B1(n10971), .B2(n15004), .A(n10967), .ZN(n10968) );
  INV_X1 U13470 ( .A(n10968), .ZN(P3_U3399) );
  OAI22_X1 U13471 ( .A1(n12996), .A2(n10969), .B1(n15016), .B2(n10381), .ZN(
        n10970) );
  AOI21_X1 U13472 ( .B1(n10971), .B2(n15016), .A(n10970), .ZN(n10972) );
  INV_X1 U13473 ( .A(n10972), .ZN(P3_U3462) );
  INV_X1 U13474 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10979) );
  MUX2_X1 U13475 ( .A(n11300), .B(P2_REG2_REG_13__SCAN_IN), .S(n10987), .Z(
        n14759) );
  MUX2_X1 U13476 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11087), .S(n13228), .Z(
        n13219) );
  NAND2_X1 U13477 ( .A1(n13220), .A2(n13219), .ZN(n14742) );
  NAND2_X1 U13478 ( .A1(n10974), .A2(n11087), .ZN(n14740) );
  OR2_X1 U13479 ( .A1(n14749), .A2(n11193), .ZN(n10976) );
  NAND2_X1 U13480 ( .A1(n14749), .A2(n11193), .ZN(n10975) );
  AND2_X1 U13481 ( .A1(n10976), .A2(n10975), .ZN(n14741) );
  AOI21_X1 U13482 ( .B1(n14742), .B2(n14740), .A(n14741), .ZN(n14744) );
  AOI21_X1 U13483 ( .B1(n11193), .B2(n10986), .A(n14744), .ZN(n14760) );
  OAI21_X1 U13484 ( .B1(n11300), .B2(n10987), .A(n14758), .ZN(n11750) );
  NAND2_X1 U13485 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n10977), .ZN(n11752) );
  OAI211_X1 U13486 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n10977), .A(n14778), 
        .B(n11752), .ZN(n10978) );
  OAI21_X1 U13487 ( .B1(n10979), .B2(n14752), .A(n10978), .ZN(n10992) );
  NAND2_X1 U13488 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14378)
         );
  XNOR2_X1 U13489 ( .A(n11761), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n10989) );
  INV_X1 U13490 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n14397) );
  INV_X1 U13491 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14736) );
  NOR2_X1 U13492 ( .A1(n10986), .A2(n14736), .ZN(n10985) );
  NAND2_X1 U13493 ( .A1(n10980), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n13224) );
  NAND2_X1 U13494 ( .A1(n13225), .A2(n13224), .ZN(n10983) );
  INV_X1 U13495 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10981) );
  MUX2_X1 U13496 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10981), .S(n13228), .Z(
        n10982) );
  NAND2_X1 U13497 ( .A1(n10983), .A2(n10982), .ZN(n13227) );
  NAND2_X1 U13498 ( .A1(n13228), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10984) );
  NAND2_X1 U13499 ( .A1(n13227), .A2(n10984), .ZN(n14738) );
  AOI211_X1 U13500 ( .C1(n10986), .C2(n14736), .A(n10985), .B(n14738), .ZN(
        n14737) );
  AOI21_X1 U13501 ( .B1(n14736), .B2(n10986), .A(n14737), .ZN(n14757) );
  MUX2_X1 U13502 ( .A(n14397), .B(P2_REG1_REG_13__SCAN_IN), .S(n10987), .Z(
        n14756) );
  NAND2_X1 U13503 ( .A1(n14757), .A2(n14756), .ZN(n14755) );
  OAI21_X1 U13504 ( .B1(n10987), .B2(n14397), .A(n14755), .ZN(n10988) );
  NAND2_X1 U13505 ( .A1(n10989), .A2(n10988), .ZN(n11759) );
  OAI211_X1 U13506 ( .C1(n10989), .C2(n10988), .A(n14783), .B(n11759), .ZN(
        n10990) );
  NAND2_X1 U13507 ( .A1(n14378), .A2(n10990), .ZN(n10991) );
  AOI211_X1 U13508 ( .C1(n14776), .C2(n11751), .A(n10992), .B(n10991), .ZN(
        n10993) );
  INV_X1 U13509 ( .A(n10993), .ZN(P2_U3228) );
  OAI21_X1 U13510 ( .B1(n10995), .B2(n10996), .A(n10994), .ZN(n14635) );
  INV_X1 U13511 ( .A(n14635), .ZN(n11011) );
  XNOR2_X1 U13512 ( .A(n10997), .B(n10996), .ZN(n11001) );
  OAI22_X1 U13513 ( .A1(n14420), .A2(n14562), .B1(n10998), .B2(n14542), .ZN(
        n10999) );
  AOI21_X1 U13514 ( .B1(n14635), .B2(n14593), .A(n10999), .ZN(n11000) );
  OAI21_X1 U13515 ( .B1(n14580), .B2(n11001), .A(n11000), .ZN(n14633) );
  NAND2_X1 U13516 ( .A1(n14633), .A2(n14576), .ZN(n11009) );
  OAI22_X1 U13517 ( .A1(n14576), .A2(n11002), .B1(n11470), .B2(n14526), .ZN(
        n11007) );
  OAI211_X1 U13518 ( .C1(n11005), .C2(n11004), .A(n14556), .B(n11003), .ZN(
        n14632) );
  NOR2_X1 U13519 ( .A1(n14632), .A2(n13947), .ZN(n11006) );
  AOI211_X1 U13520 ( .C1(n14550), .C2(n11466), .A(n11007), .B(n11006), .ZN(
        n11008) );
  OAI211_X1 U13521 ( .C1(n11011), .C2(n11010), .A(n11009), .B(n11008), .ZN(
        P1_U3284) );
  INV_X1 U13522 ( .A(n11472), .ZN(n11031) );
  NAND2_X1 U13523 ( .A1(n11021), .A2(n14606), .ZN(n14614) );
  AND2_X1 U13524 ( .A1(n12147), .A2(n13751), .ZN(n11013) );
  AOI21_X1 U13525 ( .B1(n14607), .B2(n10630), .A(n11013), .ZN(n11016) );
  AOI22_X1 U13526 ( .A1(n14607), .A2(n12146), .B1(n10630), .B2(n13751), .ZN(
        n11014) );
  XNOR2_X1 U13527 ( .A(n11014), .B(n12141), .ZN(n11015) );
  XOR2_X1 U13528 ( .A(n11016), .B(n11015), .Z(n13707) );
  INV_X1 U13529 ( .A(n11015), .ZN(n11018) );
  INV_X1 U13530 ( .A(n11016), .ZN(n11017) );
  AND2_X1 U13531 ( .A1(n12147), .A2(n13750), .ZN(n11020) );
  AOI21_X1 U13532 ( .B1(n11021), .B2(n10630), .A(n11020), .ZN(n11202) );
  AOI22_X1 U13533 ( .A1(n11021), .A2(n12146), .B1(n10630), .B2(n13750), .ZN(
        n11022) );
  XNOR2_X1 U13534 ( .A(n11022), .B(n12141), .ZN(n11201) );
  XOR2_X1 U13535 ( .A(n11202), .B(n11201), .Z(n11023) );
  OAI211_X1 U13536 ( .C1(n11024), .C2(n11023), .A(n11206), .B(n14412), .ZN(
        n11030) );
  NOR2_X1 U13537 ( .A1(n14436), .A2(n11025), .ZN(n11026) );
  AOI211_X1 U13538 ( .C1(n14414), .C2(n11028), .A(n11027), .B(n11026), .ZN(
        n11029) );
  OAI211_X1 U13539 ( .C1(n11031), .C2(n14614), .A(n11030), .B(n11029), .ZN(
        P1_U3213) );
  NAND2_X1 U13540 ( .A1(n11093), .A2(n11034), .ZN(n11153) );
  OAI21_X1 U13541 ( .B1(n11034), .B2(n11093), .A(n11153), .ZN(n11035) );
  NAND2_X1 U13542 ( .A1(n11035), .A2(n12477), .ZN(n11041) );
  INV_X1 U13543 ( .A(n11036), .ZN(n11039) );
  INV_X1 U13544 ( .A(n12519), .ZN(n11057) );
  OAI22_X1 U13545 ( .A1(n12479), .A2(n11057), .B1(n11037), .B2(n12485), .ZN(
        n11038) );
  AOI211_X1 U13546 ( .C1(n12468), .C2(n12517), .A(n11039), .B(n11038), .ZN(
        n11040) );
  OAI211_X1 U13547 ( .C1(n11218), .C2(n12495), .A(n11041), .B(n11040), .ZN(
        P3_U3170) );
  INV_X1 U13548 ( .A(n11183), .ZN(n14838) );
  NAND2_X1 U13549 ( .A1(n11245), .A2(n11241), .ZN(n11048) );
  XNOR2_X1 U13550 ( .A(n11183), .B(n11963), .ZN(n11042) );
  AND2_X1 U13551 ( .A1(n13193), .A2(n13412), .ZN(n11043) );
  NAND2_X1 U13552 ( .A1(n11042), .A2(n11043), .ZN(n11240) );
  INV_X1 U13553 ( .A(n11042), .ZN(n11045) );
  INV_X1 U13554 ( .A(n11043), .ZN(n11044) );
  NAND2_X1 U13555 ( .A1(n11045), .A2(n11044), .ZN(n11242) );
  AND2_X1 U13556 ( .A1(n11240), .A2(n11242), .ZN(n11047) );
  NAND2_X1 U13557 ( .A1(n11048), .A2(n11047), .ZN(n11046) );
  OAI211_X1 U13558 ( .C1(n11048), .C2(n11047), .A(n11046), .B(n14384), .ZN(
        n11053) );
  NAND2_X1 U13559 ( .A1(n13192), .A2(n13167), .ZN(n11050) );
  NAND2_X1 U13560 ( .A1(n13194), .A2(n13166), .ZN(n11049) );
  NAND2_X1 U13561 ( .A1(n11050), .A2(n11049), .ZN(n11079) );
  AND2_X1 U13562 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n13222) );
  NOR2_X1 U13563 ( .A1(n14672), .A2(n11086), .ZN(n11051) );
  AOI211_X1 U13564 ( .C1(n14386), .C2(n11079), .A(n13222), .B(n11051), .ZN(
        n11052) );
  OAI211_X1 U13565 ( .C1(n14838), .C2(n13162), .A(n11053), .B(n11052), .ZN(
        P2_U3208) );
  OAI21_X1 U13566 ( .B1(n11055), .B2(n12224), .A(n11054), .ZN(n14985) );
  INV_X1 U13567 ( .A(n14985), .ZN(n11069) );
  INV_X1 U13568 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n11067) );
  XNOR2_X1 U13569 ( .A(n12224), .B(n11056), .ZN(n11061) );
  OAI22_X1 U13570 ( .A1(n11058), .A2(n12906), .B1(n11057), .B2(n12908), .ZN(
        n11059) );
  AOI21_X1 U13571 ( .B1(n14985), .B2(n12667), .A(n11059), .ZN(n11060) );
  OAI21_X1 U13572 ( .B1(n12903), .B2(n11061), .A(n11060), .ZN(n14983) );
  NAND2_X1 U13573 ( .A1(n11062), .A2(n12979), .ZN(n14982) );
  OAI22_X1 U13574 ( .A1(n14982), .A2(n11064), .B1(n12910), .B2(n11063), .ZN(
        n11065) );
  NOR2_X1 U13575 ( .A1(n14983), .A2(n11065), .ZN(n11066) );
  MUX2_X1 U13576 ( .A(n11067), .B(n11066), .S(n12813), .Z(n11068) );
  OAI21_X1 U13577 ( .B1(n11069), .B2(n12656), .A(n11068), .ZN(P3_U3231) );
  NAND2_X1 U13578 ( .A1(n11072), .A2(n13194), .ZN(n11073) );
  XNOR2_X1 U13579 ( .A(n11180), .B(n11077), .ZN(n14841) );
  NAND2_X1 U13580 ( .A1(n14841), .A2(n14823), .ZN(n11082) );
  OAI21_X1 U13581 ( .B1(n11078), .B2(n11077), .A(n11185), .ZN(n11080) );
  AOI21_X1 U13582 ( .B1(n11080), .B2(n13437), .A(n11079), .ZN(n11081) );
  AND2_X1 U13583 ( .A1(n11082), .A2(n11081), .ZN(n14843) );
  NAND2_X1 U13584 ( .A1(n11183), .A2(n11083), .ZN(n11084) );
  NAND2_X1 U13585 ( .A1(n11084), .A2(n11850), .ZN(n11085) );
  OR2_X1 U13586 ( .A1(n11192), .A2(n11085), .ZN(n14836) );
  OAI22_X1 U13587 ( .A1(n11334), .A2(n11087), .B1(n11086), .B2(n13385), .ZN(
        n11088) );
  AOI21_X1 U13588 ( .B1(n11183), .B2(n13460), .A(n11088), .ZN(n11089) );
  OAI21_X1 U13589 ( .B1(n14836), .B2(n13391), .A(n11089), .ZN(n11090) );
  AOI21_X1 U13590 ( .B1(n14841), .B2(n11197), .A(n11090), .ZN(n11091) );
  OAI21_X1 U13591 ( .B1(n14843), .B2(n13453), .A(n11091), .ZN(P2_U3254) );
  NAND2_X1 U13592 ( .A1(n11093), .A2(n11092), .ZN(n11098) );
  NAND2_X1 U13593 ( .A1(n11098), .A2(n11094), .ZN(n11096) );
  AOI21_X1 U13594 ( .B1(n11096), .B2(n11095), .A(n12499), .ZN(n11100) );
  NAND2_X1 U13595 ( .A1(n11098), .A2(n11097), .ZN(n11099) );
  NAND2_X1 U13596 ( .A1(n11100), .A2(n11099), .ZN(n11104) );
  NOR2_X1 U13597 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n6678), .ZN(n14885) );
  OAI22_X1 U13598 ( .A1(n11101), .A2(n12491), .B1(n11572), .B2(n12485), .ZN(
        n11102) );
  AOI211_X1 U13599 ( .C1(n12493), .C2(n12517), .A(n14885), .B(n11102), .ZN(
        n11103) );
  OAI211_X1 U13600 ( .C1(n11571), .C2(n12495), .A(n11104), .B(n11103), .ZN(
        P3_U3179) );
  INV_X1 U13601 ( .A(n11105), .ZN(n11108) );
  INV_X1 U13602 ( .A(n13249), .ZN(n11769) );
  OAI222_X1 U13603 ( .A1(n13593), .A2(n11106), .B1(n13587), .B2(n11108), .C1(
        n11769), .C2(P2_U3088), .ZN(P2_U3309) );
  INV_X1 U13604 ( .A(n13819), .ZN(n14520) );
  OAI222_X1 U13605 ( .A1(P1_U3086), .A2(n14520), .B1(n14183), .B2(n11108), 
        .C1(n11107), .C2(n14180), .ZN(P1_U3337) );
  XNOR2_X1 U13606 ( .A(n11311), .B(n11309), .ZN(n11113) );
  NAND2_X1 U13607 ( .A1(n13747), .A2(n14033), .ZN(n11111) );
  OAI21_X1 U13608 ( .B1(n14421), .B2(n14562), .A(n11111), .ZN(n11112) );
  AOI21_X1 U13609 ( .B1(n11113), .B2(n14549), .A(n11112), .ZN(n14451) );
  OR2_X1 U13610 ( .A1(n11605), .A2(n13747), .ZN(n11114) );
  NAND2_X1 U13611 ( .A1(n11115), .A2(n11114), .ZN(n11116) );
  NAND2_X1 U13612 ( .A1(n11116), .A2(n11309), .ZN(n11307) );
  OR2_X1 U13613 ( .A1(n11116), .A2(n11309), .ZN(n11117) );
  NAND2_X1 U13614 ( .A1(n11307), .A2(n11117), .ZN(n14450) );
  NAND2_X1 U13615 ( .A1(n14431), .A2(n11118), .ZN(n11119) );
  NAND2_X1 U13616 ( .A1(n11119), .A2(n14556), .ZN(n11120) );
  OR2_X1 U13617 ( .A1(n11318), .A2(n11120), .ZN(n14447) );
  OAI22_X1 U13618 ( .A1(n14576), .A2(n11121), .B1(n14435), .B2(n14526), .ZN(
        n11122) );
  AOI21_X1 U13619 ( .B1(n14431), .B2(n14550), .A(n11122), .ZN(n11123) );
  OAI21_X1 U13620 ( .B1(n14447), .B2(n13947), .A(n11123), .ZN(n11124) );
  AOI21_X1 U13621 ( .B1(n14450), .B2(n14571), .A(n11124), .ZN(n11125) );
  OAI21_X1 U13622 ( .B1(n14451), .B2(n14578), .A(n11125), .ZN(P1_U3282) );
  AND2_X1 U13623 ( .A1(n11127), .A2(n11126), .ZN(n11129) );
  OAI211_X1 U13624 ( .C1(n11129), .C2(n11128), .A(n11170), .B(n12477), .ZN(
        n11132) );
  INV_X1 U13625 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15149) );
  NOR2_X1 U13626 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15149), .ZN(n14904) );
  OAI22_X1 U13627 ( .A1(n11562), .A2(n12491), .B1(n11696), .B2(n12485), .ZN(
        n11130) );
  AOI211_X1 U13628 ( .C1(n12493), .C2(n12516), .A(n14904), .B(n11130), .ZN(
        n11131) );
  OAI211_X1 U13629 ( .C1(n11695), .C2(n12495), .A(n11132), .B(n11131), .ZN(
        P3_U3153) );
  NAND2_X1 U13630 ( .A1(n11133), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11135) );
  NAND2_X1 U13631 ( .A1(n11135), .A2(n11134), .ZN(n11136) );
  NOR2_X1 U13632 ( .A1(n11142), .A2(n11136), .ZN(n11137) );
  XOR2_X1 U13633 ( .A(n11136), .B(n14507), .Z(n14502) );
  NOR2_X1 U13634 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14502), .ZN(n14501) );
  NOR2_X1 U13635 ( .A1(n11137), .A2(n14501), .ZN(n11139) );
  XOR2_X1 U13636 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n11145), .Z(n11138) );
  NAND2_X1 U13637 ( .A1(n11138), .A2(n11139), .ZN(n11269) );
  OAI211_X1 U13638 ( .C1(n11139), .C2(n11138), .A(n14483), .B(n11269), .ZN(
        n11151) );
  NAND2_X1 U13639 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13643)
         );
  AOI21_X1 U13640 ( .B1(n11141), .B2(n9322), .A(n11140), .ZN(n11143) );
  NOR2_X1 U13641 ( .A1(n11142), .A2(n11143), .ZN(n11144) );
  XOR2_X1 U13642 ( .A(n14507), .B(n11143), .Z(n14504) );
  NOR2_X1 U13643 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14504), .ZN(n14503) );
  NOR2_X1 U13644 ( .A1(n11144), .A2(n14503), .ZN(n11147) );
  XOR2_X1 U13645 ( .A(n11145), .B(P1_REG1_REG_16__SCAN_IN), .Z(n11146) );
  NAND2_X1 U13646 ( .A1(n11146), .A2(n11147), .ZN(n11262) );
  OAI211_X1 U13647 ( .C1(n11147), .C2(n11146), .A(n14490), .B(n11262), .ZN(
        n11148) );
  NAND2_X1 U13648 ( .A1(n13643), .A2(n11148), .ZN(n11149) );
  AOI21_X1 U13649 ( .B1(n14494), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11149), 
        .ZN(n11150) );
  OAI211_X1 U13650 ( .C1(n14521), .C2(n11271), .A(n11151), .B(n11150), .ZN(
        P1_U3259) );
  NAND2_X1 U13651 ( .A1(n11153), .A2(n11152), .ZN(n11155) );
  XNOR2_X1 U13652 ( .A(n11155), .B(n11154), .ZN(n11156) );
  NAND2_X1 U13653 ( .A1(n11156), .A2(n12477), .ZN(n11160) );
  AND2_X1 U13654 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n14864) );
  OAI22_X1 U13655 ( .A1(n11516), .A2(n12491), .B1(n11157), .B2(n12485), .ZN(
        n11158) );
  AOI211_X1 U13656 ( .C1(n12493), .C2(n12518), .A(n14864), .B(n11158), .ZN(
        n11159) );
  OAI211_X1 U13657 ( .C1(n11283), .C2(n12495), .A(n11160), .B(n11159), .ZN(
        P3_U3167) );
  INV_X1 U13658 ( .A(n11161), .ZN(n11164) );
  OAI222_X1 U13659 ( .A1(n13593), .A2(n11162), .B1(n13587), .B2(n11164), .C1(
        n13257), .C2(P2_U3088), .ZN(P2_U3308) );
  OAI222_X1 U13660 ( .A1(n11165), .A2(P1_U3086), .B1(n14183), .B2(n11164), 
        .C1(n11163), .C2(n14180), .ZN(P1_U3336) );
  INV_X1 U13661 ( .A(n11166), .ZN(n11227) );
  OAI222_X1 U13662 ( .A1(P1_U3086), .A2(n11168), .B1(n14183), .B2(n11227), 
        .C1(n11167), .C2(n14180), .ZN(P1_U3335) );
  NAND2_X1 U13663 ( .A1(n11170), .A2(n11169), .ZN(n11172) );
  NAND2_X1 U13664 ( .A1(n11172), .A2(n11171), .ZN(n11230) );
  OAI211_X1 U13665 ( .C1(n11172), .C2(n11171), .A(n11230), .B(n12477), .ZN(
        n11177) );
  NOR2_X1 U13666 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n6680), .ZN(n14922) );
  OAI22_X1 U13667 ( .A1(n11174), .A2(n12491), .B1(n11173), .B2(n12485), .ZN(
        n11175) );
  AOI211_X1 U13668 ( .C1(n12493), .C2(n12515), .A(n14922), .B(n11175), .ZN(
        n11176) );
  OAI211_X1 U13669 ( .C1(n11638), .C2(n12495), .A(n11177), .B(n11176), .ZN(
        P3_U3161) );
  AND2_X1 U13670 ( .A1(n11183), .A2(n13193), .ZN(n11179) );
  OR2_X1 U13671 ( .A1(n11183), .A2(n13193), .ZN(n11178) );
  INV_X1 U13672 ( .A(n11186), .ZN(n11181) );
  XNOR2_X1 U13673 ( .A(n11296), .B(n11181), .ZN(n14401) );
  NAND2_X1 U13674 ( .A1(n14401), .A2(n14823), .ZN(n11191) );
  NAND2_X1 U13675 ( .A1(n11183), .A2(n11182), .ZN(n11184) );
  NAND2_X1 U13676 ( .A1(n11185), .A2(n11184), .ZN(n11288) );
  XNOR2_X1 U13677 ( .A(n11288), .B(n11186), .ZN(n11189) );
  NAND2_X1 U13678 ( .A1(n13191), .A2(n13167), .ZN(n11188) );
  NAND2_X1 U13679 ( .A1(n13193), .A2(n13166), .ZN(n11187) );
  NAND2_X1 U13680 ( .A1(n11188), .A2(n11187), .ZN(n11249) );
  AOI21_X1 U13681 ( .B1(n11189), .B2(n13437), .A(n11249), .ZN(n11190) );
  INV_X1 U13682 ( .A(n11290), .ZN(n14399) );
  NAND2_X1 U13683 ( .A1(n14399), .A2(n11192), .ZN(n11330) );
  OAI211_X1 U13684 ( .C1(n14399), .C2(n11192), .A(n11850), .B(n11330), .ZN(
        n14398) );
  OAI22_X1 U13685 ( .A1(n11334), .A2(n11193), .B1(n11251), .B2(n13385), .ZN(
        n11194) );
  AOI21_X1 U13686 ( .B1(n11290), .B2(n13460), .A(n11194), .ZN(n11195) );
  OAI21_X1 U13687 ( .B1(n14398), .B2(n13391), .A(n11195), .ZN(n11196) );
  AOI21_X1 U13688 ( .B1(n14401), .B2(n11197), .A(n11196), .ZN(n11198) );
  OAI21_X1 U13689 ( .B1(n14403), .B2(n13453), .A(n11198), .ZN(P2_U3253) );
  AOI22_X1 U13690 ( .A1(n11200), .A2(n12146), .B1(n10630), .B2(n13749), .ZN(
        n11199) );
  XNOR2_X1 U13691 ( .A(n11199), .B(n12141), .ZN(n11460) );
  AOI22_X1 U13692 ( .A1(n11200), .A2(n10630), .B1(n12147), .B2(n13749), .ZN(
        n11459) );
  XNOR2_X1 U13693 ( .A(n11460), .B(n11459), .ZN(n11208) );
  INV_X1 U13694 ( .A(n11202), .ZN(n11203) );
  NAND2_X1 U13695 ( .A1(n11204), .A2(n11203), .ZN(n11205) );
  AOI21_X1 U13696 ( .B1(n11208), .B2(n11207), .A(n6622), .ZN(n11215) );
  NOR2_X1 U13697 ( .A1(n11209), .A2(n14640), .ZN(n14621) );
  AOI22_X1 U13698 ( .A1(n14414), .A2(n11210), .B1(P1_REG3_REG_8__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11211) );
  OAI21_X1 U13699 ( .B1(n14436), .B2(n11212), .A(n11211), .ZN(n11213) );
  AOI21_X1 U13700 ( .B1(n14621), .B2(n11472), .A(n11213), .ZN(n11214) );
  OAI21_X1 U13701 ( .B1(n11215), .B2(n14426), .A(n11214), .ZN(P1_U3221) );
  XNOR2_X1 U13702 ( .A(n11216), .B(n12240), .ZN(n14989) );
  INV_X1 U13703 ( .A(n12914), .ZN(n11689) );
  NAND2_X1 U13704 ( .A1(n11217), .A2(n12979), .ZN(n14986) );
  OAI22_X1 U13705 ( .A1(n11689), .A2(n14986), .B1(n11218), .B2(n12910), .ZN(
        n11225) );
  OAI211_X1 U13706 ( .C1(n11221), .C2(n11220), .A(n11219), .B(n12878), .ZN(
        n11223) );
  AOI22_X1 U13707 ( .A1(n12517), .A2(n12846), .B1(n12847), .B2(n12519), .ZN(
        n11222) );
  NAND2_X1 U13708 ( .A1(n11223), .A2(n11222), .ZN(n14987) );
  MUX2_X1 U13709 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n14987), .S(n12813), .Z(
        n11224) );
  AOI211_X1 U13710 ( .C1(n14989), .C2(n12888), .A(n11225), .B(n11224), .ZN(
        n11226) );
  INV_X1 U13711 ( .A(n11226), .ZN(P3_U3229) );
  OAI222_X1 U13712 ( .A1(n13593), .A2(n6743), .B1(P2_U3088), .B2(n11228), .C1(
        n13587), .C2(n11227), .ZN(P2_U3307) );
  NAND2_X1 U13713 ( .A1(n11230), .A2(n11229), .ZN(n11233) );
  INV_X1 U13714 ( .A(n11231), .ZN(n11232) );
  AOI21_X1 U13715 ( .B1(n11234), .B2(n11233), .A(n11232), .ZN(n11239) );
  NOR2_X1 U13716 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8370), .ZN(n14942) );
  OAI22_X1 U13717 ( .A1(n12905), .A2(n12491), .B1(n12485), .B2(n12270), .ZN(
        n11235) );
  AOI211_X1 U13718 ( .C1(n12493), .C2(n12514), .A(n14942), .B(n11235), .ZN(
        n11238) );
  INV_X1 U13719 ( .A(n11566), .ZN(n11236) );
  NAND2_X1 U13720 ( .A1(n12482), .A2(n11236), .ZN(n11237) );
  OAI211_X1 U13721 ( .C1(n11239), .C2(n12499), .A(n11238), .B(n11237), .ZN(
        P3_U3171) );
  XNOR2_X1 U13722 ( .A(n11290), .B(n6488), .ZN(n11826) );
  NAND2_X1 U13723 ( .A1(n13192), .A2(n13412), .ZN(n11825) );
  XNOR2_X1 U13724 ( .A(n11826), .B(n11825), .ZN(n11248) );
  AND2_X1 U13725 ( .A1(n11241), .A2(n11240), .ZN(n11244) );
  AOI21_X1 U13726 ( .B1(n11245), .B2(n11244), .A(n11243), .ZN(n11247) );
  INV_X1 U13727 ( .A(n11829), .ZN(n11246) );
  AOI21_X1 U13728 ( .B1(n11248), .B2(n11247), .A(n11246), .ZN(n11254) );
  NAND2_X1 U13729 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14750)
         );
  NAND2_X1 U13730 ( .A1(n14386), .A2(n11249), .ZN(n11250) );
  OAI211_X1 U13731 ( .C1(n14672), .C2(n11251), .A(n14750), .B(n11250), .ZN(
        n11252) );
  AOI21_X1 U13732 ( .B1(n11290), .B2(n14669), .A(n11252), .ZN(n11253) );
  OAI21_X1 U13733 ( .B1(n11254), .B2(n14664), .A(n11253), .ZN(P2_U3196) );
  OAI222_X1 U13734 ( .A1(P3_U3151), .A2(n11255), .B1(n13059), .B2(n7155), .C1(
        n13067), .C2(n6623), .ZN(P3_U3271) );
  INV_X1 U13735 ( .A(n11256), .ZN(n11260) );
  OAI222_X1 U13736 ( .A1(n13593), .A2(n11258), .B1(n13587), .B2(n11260), .C1(
        n11257), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI222_X1 U13737 ( .A1(n11261), .A2(P1_U3086), .B1(n14183), .B2(n11260), 
        .C1(n11259), .C2(n14180), .ZN(P1_U3334) );
  NAND2_X1 U13738 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13653)
         );
  XNOR2_X1 U13739 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n13817), .ZN(n11265) );
  OAI21_X1 U13740 ( .B1(n11271), .B2(n11263), .A(n11262), .ZN(n11264) );
  NAND2_X1 U13741 ( .A1(n11265), .A2(n11264), .ZN(n13811) );
  OAI211_X1 U13742 ( .C1(n11265), .C2(n11264), .A(n13811), .B(n14490), .ZN(
        n11266) );
  NAND2_X1 U13743 ( .A1(n13653), .A2(n11266), .ZN(n11267) );
  AOI21_X1 U13744 ( .B1(n14494), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11267), 
        .ZN(n11275) );
  NOR2_X1 U13745 ( .A1(n13817), .A2(n14041), .ZN(n11268) );
  AOI21_X1 U13746 ( .B1(n14041), .B2(n13817), .A(n11268), .ZN(n11273) );
  INV_X1 U13747 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11270) );
  OAI21_X1 U13748 ( .B1(n11271), .B2(n11270), .A(n11269), .ZN(n11272) );
  NAND2_X1 U13749 ( .A1(n11273), .A2(n11272), .ZN(n13816) );
  OAI211_X1 U13750 ( .C1(n11273), .C2(n11272), .A(n14483), .B(n13816), .ZN(
        n11274) );
  OAI211_X1 U13751 ( .C1(n14521), .C2(n13817), .A(n11275), .B(n11274), .ZN(
        P1_U3260) );
  XOR2_X1 U13752 ( .A(n12245), .B(n11276), .Z(n14990) );
  INV_X1 U13753 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n14859) );
  INV_X1 U13754 ( .A(n11277), .ZN(n11280) );
  INV_X1 U13755 ( .A(n12245), .ZN(n11279) );
  OAI21_X1 U13756 ( .B1(n11280), .B2(n11279), .A(n11278), .ZN(n11281) );
  AOI222_X1 U13757 ( .A1(n12878), .A2(n11281), .B1(n12516), .B2(n12846), .C1(
        n12518), .C2(n12847), .ZN(n14991) );
  MUX2_X1 U13758 ( .A(n14859), .B(n14991), .S(n12813), .Z(n11286) );
  AND2_X1 U13759 ( .A1(n11282), .A2(n12979), .ZN(n14993) );
  INV_X1 U13760 ( .A(n11283), .ZN(n11284) );
  AOI22_X1 U13761 ( .A1(n12914), .A2(n14993), .B1(n12868), .B2(n11284), .ZN(
        n11285) );
  OAI211_X1 U13762 ( .C1(n12918), .C2(n14990), .A(n11286), .B(n11285), .ZN(
        P3_U3228) );
  INV_X1 U13763 ( .A(n13192), .ZN(n11289) );
  OR2_X1 U13764 ( .A1(n11290), .A2(n11289), .ZN(n11287) );
  NAND2_X1 U13765 ( .A1(n11288), .A2(n11287), .ZN(n11292) );
  NAND2_X1 U13766 ( .A1(n11290), .A2(n11289), .ZN(n11291) );
  NAND2_X1 U13767 ( .A1(n11292), .A2(n11291), .ZN(n11326) );
  XNOR2_X1 U13768 ( .A(n11326), .B(n11298), .ZN(n11293) );
  NAND2_X1 U13769 ( .A1(n11293), .A2(n13437), .ZN(n11294) );
  AOI22_X1 U13770 ( .A1(n13190), .A2(n13167), .B1(n13192), .B2(n13166), .ZN(
        n14659) );
  NAND2_X1 U13771 ( .A1(n11294), .A2(n14659), .ZN(n14394) );
  INV_X1 U13772 ( .A(n14394), .ZN(n11305) );
  XOR2_X1 U13773 ( .A(n11298), .B(n11339), .Z(n14396) );
  XOR2_X1 U13774 ( .A(n14670), .B(n11330), .Z(n11299) );
  NAND2_X1 U13775 ( .A1(n11299), .A2(n11850), .ZN(n14392) );
  OAI22_X1 U13776 ( .A1(n11334), .A2(n11300), .B1(n14673), .B2(n13385), .ZN(
        n11301) );
  AOI21_X1 U13777 ( .B1(n14670), .B2(n13460), .A(n11301), .ZN(n11302) );
  OAI21_X1 U13778 ( .B1(n14392), .B2(n13391), .A(n11302), .ZN(n11303) );
  AOI21_X1 U13779 ( .B1(n14396), .B2(n13457), .A(n11303), .ZN(n11304) );
  OAI21_X1 U13780 ( .B1(n13453), .B2(n11305), .A(n11304), .ZN(P2_U3252) );
  NAND2_X1 U13781 ( .A1(n11307), .A2(n11306), .ZN(n11308) );
  NAND2_X1 U13782 ( .A1(n11308), .A2(n11314), .ZN(n11367) );
  OAI21_X1 U13783 ( .B1(n11308), .B2(n11314), .A(n11367), .ZN(n11501) );
  OAI22_X1 U13784 ( .A1(n11312), .A2(n14542), .B1(n12038), .B2(n14562), .ZN(
        n11317) );
  INV_X1 U13785 ( .A(n11309), .ZN(n11310) );
  OR2_X1 U13786 ( .A1(n14431), .A2(n11312), .ZN(n11313) );
  INV_X1 U13787 ( .A(n11314), .ZN(n11361) );
  XNOR2_X1 U13788 ( .A(n11362), .B(n11361), .ZN(n11315) );
  NOR2_X1 U13789 ( .A1(n11315), .A2(n14580), .ZN(n11316) );
  AOI211_X1 U13790 ( .C1(n14593), .C2(n11501), .A(n11317), .B(n11316), .ZN(
        n11505) );
  INV_X1 U13791 ( .A(n11318), .ZN(n11319) );
  AND2_X1 U13792 ( .A1(n11816), .A2(n11318), .ZN(n11370) );
  AOI211_X1 U13793 ( .C1(n11503), .C2(n11319), .A(n14058), .B(n11370), .ZN(
        n11502) );
  NOR2_X1 U13794 ( .A1(n11816), .A2(n14530), .ZN(n11322) );
  OAI22_X1 U13795 ( .A1(n14576), .A2(n11320), .B1(n11810), .B2(n14526), .ZN(
        n11321) );
  AOI211_X1 U13796 ( .C1(n11502), .C2(n14558), .A(n11322), .B(n11321), .ZN(
        n11324) );
  NAND2_X1 U13797 ( .A1(n11501), .A2(n14559), .ZN(n11323) );
  OAI211_X1 U13798 ( .C1(n11505), .C2(n14578), .A(n11324), .B(n11323), .ZN(
        P1_U3281) );
  INV_X1 U13799 ( .A(n11340), .ZN(n11327) );
  INV_X1 U13800 ( .A(n13191), .ZN(n11328) );
  AND2_X1 U13801 ( .A1(n14670), .A2(n11328), .ZN(n11325) );
  OAI21_X1 U13802 ( .B1(n11327), .B2(n6613), .A(n11652), .ZN(n11329) );
  OAI22_X1 U13803 ( .A1(n11659), .A2(n13144), .B1(n11328), .B2(n13142), .ZN(
        n14376) );
  AOI21_X1 U13804 ( .B1(n11329), .B2(n13437), .A(n14376), .ZN(n13554) );
  NOR2_X2 U13805 ( .A1(n11331), .A2(n6677), .ZN(n11649) );
  AOI211_X1 U13806 ( .C1(n6677), .C2(n11331), .A(n13412), .B(n11649), .ZN(
        n13550) );
  INV_X1 U13807 ( .A(n6677), .ZN(n11332) );
  NOR2_X1 U13808 ( .A1(n11332), .A2(n13443), .ZN(n11336) );
  INV_X1 U13809 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11333) );
  OAI22_X1 U13810 ( .A1(n11334), .A2(n11333), .B1(n14380), .B2(n13385), .ZN(
        n11335) );
  AOI211_X1 U13811 ( .C1(n13550), .C2(n13455), .A(n11336), .B(n11335), .ZN(
        n11343) );
  NAND2_X1 U13812 ( .A1(n14670), .A2(n13191), .ZN(n11338) );
  NOR2_X1 U13813 ( .A1(n14670), .A2(n13191), .ZN(n11337) );
  OR2_X1 U13814 ( .A1(n11341), .A2(n11340), .ZN(n13552) );
  NAND2_X1 U13815 ( .A1(n11341), .A2(n11340), .ZN(n13551) );
  NAND3_X1 U13816 ( .A1(n13552), .A2(n13551), .A3(n13457), .ZN(n11342) );
  OAI211_X1 U13817 ( .C1(n13453), .C2(n13554), .A(n11343), .B(n11342), .ZN(
        P2_U3251) );
  OAI211_X1 U13818 ( .C1(n11346), .C2(n11345), .A(n11344), .B(n12477), .ZN(
        n11350) );
  INV_X1 U13819 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15134) );
  NOR2_X1 U13820 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15134), .ZN(n14953) );
  OAI22_X1 U13821 ( .A1(n12876), .A2(n12491), .B1(n11347), .B2(n12485), .ZN(
        n11348) );
  AOI211_X1 U13822 ( .C1(n12493), .C2(n12513), .A(n14953), .B(n11348), .ZN(
        n11349) );
  OAI211_X1 U13823 ( .C1(n11690), .C2(n12495), .A(n11350), .B(n11349), .ZN(
        P3_U3157) );
  OAI21_X1 U13824 ( .B1(n11352), .B2(n12197), .A(n11351), .ZN(n11576) );
  OAI211_X1 U13825 ( .C1(n8791), .C2(n8790), .A(n12878), .B(n11514), .ZN(
        n11354) );
  AOI22_X1 U13826 ( .A1(n12847), .A2(n12517), .B1(n12515), .B2(n12846), .ZN(
        n11353) );
  NAND2_X1 U13827 ( .A1(n11354), .A2(n11353), .ZN(n11573) );
  AOI21_X1 U13828 ( .B1(n8900), .B2(n11576), .A(n11573), .ZN(n11360) );
  INV_X1 U13829 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n11355) );
  OAI22_X1 U13830 ( .A1(n13053), .A2(n11572), .B1(n11355), .B2(n15004), .ZN(
        n11356) );
  INV_X1 U13831 ( .A(n11356), .ZN(n11357) );
  OAI21_X1 U13832 ( .B1(n11360), .B2(n15006), .A(n11357), .ZN(P3_U3408) );
  AOI22_X1 U13833 ( .A1(n8875), .A2(n11358), .B1(n15014), .B2(
        P3_REG1_REG_6__SCAN_IN), .ZN(n11359) );
  OAI21_X1 U13834 ( .B1(n11360), .B2(n15014), .A(n11359), .ZN(P3_U3465) );
  NAND2_X1 U13835 ( .A1(n11362), .A2(n11361), .ZN(n11364) );
  NAND2_X1 U13836 ( .A1(n11816), .A2(n13745), .ZN(n11363) );
  NAND2_X1 U13837 ( .A1(n11364), .A2(n11363), .ZN(n11665) );
  XNOR2_X1 U13838 ( .A(n11665), .B(n11664), .ZN(n11365) );
  OAI222_X1 U13839 ( .A1(n14562), .A2(n13731), .B1(n11365), .B2(n14580), .C1(
        n14542), .C2(n14421), .ZN(n14444) );
  INV_X1 U13840 ( .A(n14444), .ZN(n11375) );
  INV_X1 U13841 ( .A(n11664), .ZN(n11368) );
  OAI21_X1 U13842 ( .B1(n11369), .B2(n11368), .A(n11673), .ZN(n14446) );
  OAI211_X1 U13843 ( .C1(n14443), .C2(n11370), .A(n14556), .B(n11678), .ZN(
        n14442) );
  OAI22_X1 U13844 ( .A1(n14576), .A2(n9330), .B1(n13681), .B2(n14526), .ZN(
        n11371) );
  AOI21_X1 U13845 ( .B1(n11671), .B2(n14550), .A(n11371), .ZN(n11372) );
  OAI21_X1 U13846 ( .B1(n14442), .B2(n13947), .A(n11372), .ZN(n11373) );
  AOI21_X1 U13847 ( .B1(n14446), .B2(n14571), .A(n11373), .ZN(n11374) );
  OAI21_X1 U13848 ( .B1(n11375), .B2(n14578), .A(n11374), .ZN(P1_U3280) );
  INV_X1 U13849 ( .A(n14938), .ZN(n11435) );
  AOI21_X1 U13850 ( .B1(n14866), .B2(n11380), .A(n14857), .ZN(n14876) );
  NAND2_X1 U13851 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n14882), .ZN(n11381) );
  OAI21_X1 U13852 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n14882), .A(n11381), .ZN(
        n14875) );
  NOR2_X1 U13853 ( .A1(n14876), .A2(n14875), .ZN(n14874) );
  INV_X1 U13854 ( .A(n11381), .ZN(n11382) );
  NOR2_X1 U13855 ( .A1(n11422), .A2(n11383), .ZN(n11384) );
  NAND2_X1 U13856 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n14919), .ZN(n11385) );
  OAI21_X1 U13857 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n14919), .A(n11385), .ZN(
        n14912) );
  NOR2_X1 U13858 ( .A1(n11435), .A2(n11386), .ZN(n11387) );
  NAND2_X1 U13859 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n14969), .ZN(n11388) );
  OAI21_X1 U13860 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n14969), .A(n11388), 
        .ZN(n14957) );
  AOI21_X1 U13861 ( .B1(n12912), .B2(n11389), .A(n11480), .ZN(n11454) );
  INV_X1 U13862 ( .A(n11490), .ZN(n11479) );
  NAND2_X1 U13863 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n14969), .ZN(n11400) );
  AOI22_X1 U13864 ( .A1(n11441), .A2(n11440), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n14969), .ZN(n14952) );
  NAND2_X1 U13865 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n14919), .ZN(n11397) );
  AOI22_X1 U13866 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n14919), .B1(n11428), 
        .B2(n11427), .ZN(n14924) );
  NAND2_X1 U13867 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n14882), .ZN(n11394) );
  AOI22_X1 U13868 ( .A1(n11415), .A2(n11413), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n14882), .ZN(n14887) );
  OAI22_X1 U13869 ( .A1(n11391), .A2(n11390), .B1(n11406), .B2(n15009), .ZN(
        n11392) );
  XNOR2_X1 U13870 ( .A(n11392), .B(n14866), .ZN(n14869) );
  INV_X1 U13871 ( .A(n11392), .ZN(n11393) );
  NAND2_X1 U13872 ( .A1(n14887), .A2(n14888), .ZN(n14886) );
  NAND2_X1 U13873 ( .A1(n14901), .A2(n11395), .ZN(n11396) );
  NAND2_X1 U13874 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n14906), .ZN(n14905) );
  NAND2_X1 U13875 ( .A1(n11396), .A2(n14905), .ZN(n14925) );
  NAND2_X1 U13876 ( .A1(n14938), .A2(n11398), .ZN(n11399) );
  XNOR2_X1 U13877 ( .A(n11435), .B(n11398), .ZN(n14945) );
  NAND2_X1 U13878 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n14945), .ZN(n14944) );
  NAND2_X1 U13879 ( .A1(n11399), .A2(n14944), .ZN(n14951) );
  NAND2_X1 U13880 ( .A1(n14952), .A2(n14951), .ZN(n14950) );
  NAND2_X1 U13881 ( .A1(n11400), .A2(n14950), .ZN(n11484) );
  XNOR2_X1 U13882 ( .A(n11479), .B(n11484), .ZN(n11401) );
  NAND2_X1 U13883 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n11401), .ZN(n11485) );
  OAI21_X1 U13884 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n11401), .A(n11485), 
        .ZN(n11452) );
  NAND2_X1 U13885 ( .A1(n14343), .A2(n11479), .ZN(n11402) );
  INV_X1 U13886 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n15083) );
  OR2_X1 U13887 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15083), .ZN(n11591) );
  OAI211_X1 U13888 ( .C1(n14223), .C2(n14975), .A(n11402), .B(n11591), .ZN(
        n11451) );
  NAND2_X1 U13889 ( .A1(n11404), .A2(n11403), .ZN(n11409) );
  INV_X1 U13890 ( .A(n11405), .ZN(n11407) );
  NAND2_X1 U13891 ( .A1(n11407), .A2(n11406), .ZN(n11408) );
  NAND2_X1 U13892 ( .A1(n11409), .A2(n11408), .ZN(n14862) );
  MUX2_X1 U13893 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12601), .Z(n11410) );
  NAND2_X1 U13894 ( .A1(n11410), .A2(n14866), .ZN(n14860) );
  NAND2_X1 U13895 ( .A1(n14862), .A2(n14860), .ZN(n14880) );
  INV_X1 U13896 ( .A(n11410), .ZN(n11412) );
  NAND2_X1 U13897 ( .A1(n11412), .A2(n11411), .ZN(n14861) );
  NAND2_X1 U13898 ( .A1(n14880), .A2(n14861), .ZN(n11419) );
  MUX2_X1 U13899 ( .A(n11414), .B(n11413), .S(n12601), .Z(n11416) );
  NAND2_X1 U13900 ( .A1(n11416), .A2(n11415), .ZN(n14895) );
  INV_X1 U13901 ( .A(n11416), .ZN(n11417) );
  NAND2_X1 U13902 ( .A1(n11417), .A2(n14882), .ZN(n11418) );
  AND2_X1 U13903 ( .A1(n14895), .A2(n11418), .ZN(n14878) );
  NAND2_X1 U13904 ( .A1(n11419), .A2(n14878), .ZN(n14899) );
  NAND2_X1 U13905 ( .A1(n14899), .A2(n14895), .ZN(n11426) );
  MUX2_X1 U13906 ( .A(n11421), .B(n11420), .S(n12601), .Z(n11423) );
  NAND2_X1 U13907 ( .A1(n11423), .A2(n11422), .ZN(n14913) );
  INV_X1 U13908 ( .A(n11423), .ZN(n11424) );
  NAND2_X1 U13909 ( .A1(n11424), .A2(n14901), .ZN(n11425) );
  AND2_X1 U13910 ( .A1(n14913), .A2(n11425), .ZN(n14897) );
  NAND2_X1 U13911 ( .A1(n11426), .A2(n14897), .ZN(n14917) );
  NAND2_X1 U13912 ( .A1(n14917), .A2(n14913), .ZN(n11432) );
  MUX2_X1 U13913 ( .A(n11639), .B(n11427), .S(n12601), .Z(n11429) );
  NAND2_X1 U13914 ( .A1(n11429), .A2(n11428), .ZN(n14932) );
  INV_X1 U13915 ( .A(n11429), .ZN(n11430) );
  NAND2_X1 U13916 ( .A1(n11430), .A2(n14919), .ZN(n11431) );
  AND2_X1 U13917 ( .A1(n14932), .A2(n11431), .ZN(n14915) );
  NAND2_X1 U13918 ( .A1(n11432), .A2(n14915), .ZN(n14936) );
  NAND2_X1 U13919 ( .A1(n14936), .A2(n14932), .ZN(n11439) );
  MUX2_X1 U13920 ( .A(n11434), .B(n11433), .S(n12601), .Z(n11436) );
  NAND2_X1 U13921 ( .A1(n11436), .A2(n11435), .ZN(n14962) );
  INV_X1 U13922 ( .A(n11436), .ZN(n11437) );
  NAND2_X1 U13923 ( .A1(n11437), .A2(n14938), .ZN(n11438) );
  AND2_X1 U13924 ( .A1(n14962), .A2(n11438), .ZN(n14934) );
  NAND2_X1 U13925 ( .A1(n11439), .A2(n14934), .ZN(n14963) );
  MUX2_X1 U13926 ( .A(n11691), .B(n11440), .S(n12601), .Z(n11442) );
  NAND2_X1 U13927 ( .A1(n11442), .A2(n11441), .ZN(n11445) );
  INV_X1 U13928 ( .A(n11442), .ZN(n11443) );
  NAND2_X1 U13929 ( .A1(n11443), .A2(n14969), .ZN(n11444) );
  NAND2_X1 U13930 ( .A1(n11445), .A2(n11444), .ZN(n14961) );
  AOI21_X1 U13931 ( .B1(n14963), .B2(n14962), .A(n14961), .ZN(n14966) );
  INV_X1 U13932 ( .A(n11445), .ZN(n11446) );
  NOR2_X1 U13933 ( .A1(n14966), .A2(n11446), .ZN(n11448) );
  MUX2_X1 U13934 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12601), .Z(n11491) );
  XNOR2_X1 U13935 ( .A(n11491), .B(n11490), .ZN(n11447) );
  NOR2_X1 U13936 ( .A1(n11448), .A2(n11447), .ZN(n11493) );
  AOI21_X1 U13937 ( .B1(n11448), .B2(n11447), .A(n11493), .ZN(n11449) );
  NOR2_X1 U13938 ( .A1(n11449), .A2(n14939), .ZN(n11450) );
  AOI211_X1 U13939 ( .C1(n14954), .C2(n11452), .A(n11451), .B(n11450), .ZN(
        n11453) );
  OAI21_X1 U13940 ( .B1(n11454), .B2(n14959), .A(n11453), .ZN(P3_U3193) );
  INV_X1 U13941 ( .A(n11455), .ZN(n11457) );
  OAI222_X1 U13942 ( .A1(n13593), .A2(n11458), .B1(n13587), .B2(n11457), .C1(
        n11456), .C2(P2_U3088), .ZN(P2_U3305) );
  AOI22_X1 U13943 ( .A1(n11466), .A2(n10630), .B1(n12147), .B2(n13748), .ZN(
        n11598) );
  NAND2_X1 U13944 ( .A1(n11466), .A2(n12146), .ZN(n11462) );
  NAND2_X1 U13945 ( .A1(n13748), .A2(n10630), .ZN(n11461) );
  NAND2_X1 U13946 ( .A1(n11462), .A2(n11461), .ZN(n11463) );
  INV_X2 U13947 ( .A(n12042), .ZN(n12141) );
  XNOR2_X1 U13948 ( .A(n11463), .B(n12141), .ZN(n11597) );
  XOR2_X1 U13949 ( .A(n11598), .B(n11597), .Z(n11464) );
  AOI21_X1 U13950 ( .B1(n11465), .B2(n11464), .A(n11600), .ZN(n11474) );
  AND2_X1 U13951 ( .A1(n11466), .A2(n14606), .ZN(n14630) );
  INV_X1 U13952 ( .A(n14419), .ZN(n13685) );
  OAI22_X1 U13953 ( .A1(n14422), .A2(n14420), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11467), .ZN(n11468) );
  AOI21_X1 U13954 ( .B1(n13685), .B2(n13749), .A(n11468), .ZN(n11469) );
  OAI21_X1 U13955 ( .B1(n11470), .B2(n14436), .A(n11469), .ZN(n11471) );
  AOI21_X1 U13956 ( .B1(n14630), .B2(n11472), .A(n11471), .ZN(n11473) );
  OAI21_X1 U13957 ( .B1(n11474), .B2(n14426), .A(n11473), .ZN(P1_U3231) );
  INV_X1 U13958 ( .A(n11475), .ZN(n11476) );
  OAI222_X1 U13959 ( .A1(P3_U3151), .A2(n11477), .B1(n13059), .B2(n15169), 
        .C1(n13067), .C2(n11476), .ZN(P3_U3270) );
  NOR2_X1 U13960 ( .A1(n11479), .A2(n11478), .ZN(n11481) );
  AOI22_X1 U13961 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n11539), .B1(n11545), 
        .B2(n12882), .ZN(n11482) );
  AOI21_X1 U13962 ( .B1(n11483), .B2(n11482), .A(n11536), .ZN(n11500) );
  AOI22_X1 U13963 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n11545), .B1(n11539), 
        .B2(n8543), .ZN(n11488) );
  NAND2_X1 U13964 ( .A1(n11490), .A2(n11484), .ZN(n11486) );
  NAND2_X1 U13965 ( .A1(n11486), .A2(n11485), .ZN(n11487) );
  NAND2_X1 U13966 ( .A1(n11488), .A2(n11487), .ZN(n11538) );
  OAI21_X1 U13967 ( .B1(n11488), .B2(n11487), .A(n11538), .ZN(n11498) );
  INV_X1 U13968 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14225) );
  NAND2_X1 U13969 ( .A1(n14343), .A2(n11539), .ZN(n11489) );
  OR2_X1 U13970 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15111), .ZN(n11624) );
  OAI211_X1 U13971 ( .C1(n14225), .C2(n14975), .A(n11489), .B(n11624), .ZN(
        n11497) );
  MUX2_X1 U13972 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12601), .Z(n11546) );
  XNOR2_X1 U13973 ( .A(n11546), .B(n11545), .ZN(n11495) );
  NOR2_X1 U13974 ( .A1(n11491), .A2(n11490), .ZN(n11492) );
  OR2_X1 U13975 ( .A1(n11493), .A2(n11492), .ZN(n11494) );
  NOR3_X1 U13976 ( .A1(n11493), .A2(n11492), .A3(n11495), .ZN(n11544) );
  AOI211_X1 U13977 ( .C1(n11495), .C2(n11494), .A(n14939), .B(n11544), .ZN(
        n11496) );
  AOI211_X1 U13978 ( .C1(n14954), .C2(n11498), .A(n11497), .B(n11496), .ZN(
        n11499) );
  OAI21_X1 U13979 ( .B1(n11500), .B2(n14959), .A(n11499), .ZN(P3_U3194) );
  INV_X1 U13980 ( .A(n11501), .ZN(n11506) );
  AOI21_X1 U13981 ( .B1(n11503), .B2(n14606), .A(n11502), .ZN(n11504) );
  OAI211_X1 U13982 ( .C1(n11506), .C2(n14609), .A(n11505), .B(n11504), .ZN(
        n11508) );
  NAND2_X1 U13983 ( .A1(n11508), .A2(n14657), .ZN(n11507) );
  OAI21_X1 U13984 ( .B1(n14657), .B2(n9995), .A(n11507), .ZN(P1_U3540) );
  INV_X1 U13985 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11510) );
  NAND2_X1 U13986 ( .A1(n11508), .A2(n14646), .ZN(n11509) );
  OAI21_X1 U13987 ( .B1(n14646), .B2(n11510), .A(n11509), .ZN(P1_U3495) );
  OAI21_X1 U13988 ( .B1(n11512), .B2(n12258), .A(n11511), .ZN(n11700) );
  NAND2_X1 U13989 ( .A1(n11514), .A2(n11513), .ZN(n11557) );
  NAND2_X1 U13990 ( .A1(n11557), .A2(n11515), .ZN(n11632) );
  OAI211_X1 U13991 ( .C1(n11557), .C2(n11515), .A(n11632), .B(n12878), .ZN(
        n11519) );
  OAI22_X1 U13992 ( .A1(n11516), .A2(n12906), .B1(n11562), .B2(n12908), .ZN(
        n11517) );
  INV_X1 U13993 ( .A(n11517), .ZN(n11518) );
  NAND2_X1 U13994 ( .A1(n11519), .A2(n11518), .ZN(n11697) );
  AOI21_X1 U13995 ( .B1(n8900), .B2(n11700), .A(n11697), .ZN(n11525) );
  INV_X1 U13996 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n11520) );
  OAI22_X1 U13997 ( .A1(n13053), .A2(n11696), .B1(n11520), .B2(n15004), .ZN(
        n11521) );
  INV_X1 U13998 ( .A(n11521), .ZN(n11522) );
  OAI21_X1 U13999 ( .B1(n11525), .B2(n15006), .A(n11522), .ZN(P3_U3411) );
  OAI22_X1 U14000 ( .A1(n12996), .A2(n11696), .B1(n15016), .B2(n11420), .ZN(
        n11523) );
  INV_X1 U14001 ( .A(n11523), .ZN(n11524) );
  OAI21_X1 U14002 ( .B1(n11525), .B2(n15014), .A(n11524), .ZN(P3_U3466) );
  INV_X1 U14003 ( .A(n11529), .ZN(n11528) );
  NAND2_X1 U14004 ( .A1(n13585), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11527) );
  OAI211_X1 U14005 ( .C1(n11528), .C2(n13587), .A(n11527), .B(n11526), .ZN(
        P2_U3304) );
  NAND2_X1 U14006 ( .A1(n11529), .A2(n14178), .ZN(n11531) );
  OAI211_X1 U14007 ( .C1(n11532), .C2(n14180), .A(n11531), .B(n11530), .ZN(
        P1_U3332) );
  INV_X1 U14008 ( .A(n11533), .ZN(n11534) );
  OAI222_X1 U14009 ( .A1(P3_U3151), .A2(n11535), .B1(n13059), .B2(n15171), 
        .C1(n13067), .C2(n11534), .ZN(P3_U3269) );
  AOI21_X1 U14010 ( .B1(n8568), .B2(n11537), .A(n12525), .ZN(n11552) );
  OAI21_X1 U14011 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n11540), .A(n12530), 
        .ZN(n11543) );
  INV_X1 U14012 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14226) );
  NAND2_X1 U14013 ( .A1(n14343), .A2(n12538), .ZN(n11541) );
  INV_X1 U14014 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n15107) );
  OR2_X1 U14015 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15107), .ZN(n11727) );
  OAI211_X1 U14016 ( .C1(n14226), .C2(n14975), .A(n11541), .B(n11727), .ZN(
        n11542) );
  AOI21_X1 U14017 ( .B1(n11543), .B2(n14954), .A(n11542), .ZN(n11551) );
  AOI21_X1 U14018 ( .B1(n11546), .B2(n11545), .A(n11544), .ZN(n11548) );
  MUX2_X1 U14019 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12601), .Z(n12537) );
  XNOR2_X1 U14020 ( .A(n12537), .B(n12538), .ZN(n11547) );
  NAND2_X1 U14021 ( .A1(n11548), .A2(n11547), .ZN(n12545) );
  OAI21_X1 U14022 ( .B1(n11548), .B2(n11547), .A(n12545), .ZN(n11549) );
  NAND2_X1 U14023 ( .A1(n11549), .A2(n14964), .ZN(n11550) );
  OAI211_X1 U14024 ( .C1(n11552), .C2(n14959), .A(n11551), .B(n11550), .ZN(
        P3_U3195) );
  NAND2_X1 U14025 ( .A1(n11557), .A2(n11553), .ZN(n11555) );
  NAND2_X1 U14026 ( .A1(n11555), .A2(n11554), .ZN(n11561) );
  NAND2_X1 U14027 ( .A1(n11557), .A2(n11556), .ZN(n11559) );
  AND2_X1 U14028 ( .A1(n11559), .A2(n11558), .ZN(n11560) );
  OAI211_X1 U14029 ( .C1(n11561), .C2(n12200), .A(n11560), .B(n12878), .ZN(
        n11564) );
  OR2_X1 U14030 ( .A1(n11562), .A2(n12906), .ZN(n11563) );
  OAI211_X1 U14031 ( .C1(n12905), .C2(n12908), .A(n11564), .B(n11563), .ZN(
        n11578) );
  INV_X1 U14032 ( .A(n11578), .ZN(n11570) );
  XNOR2_X1 U14033 ( .A(n11565), .B(n12268), .ZN(n11579) );
  NOR2_X1 U14034 ( .A1(n12870), .A2(n12270), .ZN(n11568) );
  OAI22_X1 U14035 ( .A1(n12813), .A2(n11434), .B1(n11566), .B2(n12910), .ZN(
        n11567) );
  AOI211_X1 U14036 ( .C1(n11579), .C2(n12888), .A(n11568), .B(n11567), .ZN(
        n11569) );
  OAI21_X1 U14037 ( .B1(n11570), .B2(n12891), .A(n11569), .ZN(P3_U3224) );
  OAI22_X1 U14038 ( .A1(n12870), .A2(n11572), .B1(n11571), .B2(n12910), .ZN(
        n11575) );
  MUX2_X1 U14039 ( .A(n11573), .B(P3_REG2_REG_6__SCAN_IN), .S(n12786), .Z(
        n11574) );
  AOI211_X1 U14040 ( .C1(n12888), .C2(n11576), .A(n11575), .B(n11574), .ZN(
        n11577) );
  INV_X1 U14041 ( .A(n11577), .ZN(P3_U3227) );
  AOI21_X1 U14042 ( .B1(n11579), .B2(n8900), .A(n11578), .ZN(n11585) );
  INV_X1 U14043 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n11580) );
  OAI22_X1 U14044 ( .A1(n13053), .A2(n12270), .B1(n11580), .B2(n15004), .ZN(
        n11581) );
  INV_X1 U14045 ( .A(n11581), .ZN(n11582) );
  OAI21_X1 U14046 ( .B1(n11585), .B2(n15006), .A(n11582), .ZN(P3_U3417) );
  OAI22_X1 U14047 ( .A1(n12996), .A2(n12270), .B1(n15016), .B2(n11433), .ZN(
        n11583) );
  INV_X1 U14048 ( .A(n11583), .ZN(n11584) );
  OAI21_X1 U14049 ( .B1(n11585), .B2(n15014), .A(n11584), .ZN(P3_U3468) );
  INV_X1 U14050 ( .A(n11586), .ZN(n11588) );
  NAND2_X1 U14051 ( .A1(n11588), .A2(n11587), .ZN(n11589) );
  XNOR2_X1 U14052 ( .A(n11589), .B(n12876), .ZN(n11596) );
  INV_X1 U14053 ( .A(n12911), .ZN(n11594) );
  NOR2_X1 U14054 ( .A1(n12485), .A2(n12909), .ZN(n11593) );
  OR2_X1 U14055 ( .A1(n12491), .A2(n12907), .ZN(n11590) );
  OAI211_X1 U14056 ( .C1(n12479), .C2(n12905), .A(n11591), .B(n11590), .ZN(
        n11592) );
  AOI211_X1 U14057 ( .C1(n11594), .C2(n12482), .A(n11593), .B(n11592), .ZN(
        n11595) );
  OAI21_X1 U14058 ( .B1(n11596), .B2(n12499), .A(n11595), .ZN(P3_U3176) );
  INV_X1 U14059 ( .A(n11605), .ZN(n14641) );
  INV_X1 U14060 ( .A(n11597), .ZN(n11599) );
  NAND2_X1 U14061 ( .A1(n11605), .A2(n12146), .ZN(n11602) );
  NAND2_X1 U14062 ( .A1(n13747), .A2(n10630), .ZN(n11601) );
  NAND2_X1 U14063 ( .A1(n11602), .A2(n11601), .ZN(n11603) );
  XNOR2_X1 U14064 ( .A(n11603), .B(n12141), .ZN(n11798) );
  AND2_X1 U14065 ( .A1(n12147), .A2(n13747), .ZN(n11604) );
  AOI21_X1 U14066 ( .B1(n11605), .B2(n10630), .A(n11604), .ZN(n11796) );
  XNOR2_X1 U14067 ( .A(n11798), .B(n11796), .ZN(n11606) );
  OAI211_X1 U14068 ( .C1(n11607), .C2(n11606), .A(n11800), .B(n14412), .ZN(
        n11615) );
  INV_X1 U14069 ( .A(n11608), .ZN(n11613) );
  AOI21_X1 U14070 ( .B1(n11610), .B2(n11609), .A(n13672), .ZN(n11611) );
  AOI211_X1 U14071 ( .C1(n13733), .C2(n11613), .A(n11612), .B(n11611), .ZN(
        n11614) );
  OAI211_X1 U14072 ( .C1(n14641), .C2(n13737), .A(n11615), .B(n11614), .ZN(
        P1_U3217) );
  INV_X1 U14073 ( .A(n11616), .ZN(n11617) );
  INV_X1 U14074 ( .A(SI_27_), .ZN(n15059) );
  AOI21_X1 U14075 ( .B1(n11621), .B2(n11620), .A(n11619), .ZN(n11629) );
  INV_X1 U14076 ( .A(n12881), .ZN(n11627) );
  NOR2_X1 U14077 ( .A1(n11622), .A2(n12485), .ZN(n11626) );
  OR2_X1 U14078 ( .A1(n12491), .A2(n12875), .ZN(n11623) );
  OAI211_X1 U14079 ( .C1(n12479), .C2(n12876), .A(n11624), .B(n11623), .ZN(
        n11625) );
  AOI211_X1 U14080 ( .C1(n11627), .C2(n12482), .A(n11626), .B(n11625), .ZN(
        n11628) );
  OAI21_X1 U14081 ( .B1(n11629), .B2(n12499), .A(n11628), .ZN(P3_U3164) );
  XNOR2_X1 U14082 ( .A(n11630), .B(n12263), .ZN(n14998) );
  INV_X1 U14083 ( .A(n14998), .ZN(n11643) );
  NAND2_X1 U14084 ( .A1(n11632), .A2(n11631), .ZN(n11633) );
  AOI21_X1 U14085 ( .B1(n12263), .B2(n11633), .A(n6610), .ZN(n11636) );
  AOI22_X1 U14086 ( .A1(n12515), .A2(n12847), .B1(n12846), .B2(n12513), .ZN(
        n11635) );
  NAND2_X1 U14087 ( .A1(n14998), .A2(n12667), .ZN(n11634) );
  OAI211_X1 U14088 ( .C1(n11636), .C2(n12903), .A(n11635), .B(n11634), .ZN(
        n14995) );
  NAND2_X1 U14089 ( .A1(n14995), .A2(n12813), .ZN(n11642) );
  AND2_X1 U14090 ( .A1(n11637), .A2(n12979), .ZN(n14996) );
  OAI22_X1 U14091 ( .A1(n12813), .A2(n11639), .B1(n11638), .B2(n12910), .ZN(
        n11640) );
  AOI21_X1 U14092 ( .B1(n12914), .B2(n14996), .A(n11640), .ZN(n11641) );
  OAI211_X1 U14093 ( .C1(n11643), .C2(n12656), .A(n11642), .B(n11641), .ZN(
        P3_U3225) );
  NAND2_X1 U14094 ( .A1(n6677), .A2(n13190), .ZN(n11644) );
  NAND2_X1 U14095 ( .A1(n13551), .A2(n11644), .ZN(n11788) );
  INV_X1 U14096 ( .A(n11788), .ZN(n11646) );
  OR2_X1 U14097 ( .A1(n13546), .A2(n13189), .ZN(n11647) );
  OAI21_X1 U14098 ( .B1(n6617), .B2(n11656), .A(n11845), .ZN(n13544) );
  AOI211_X1 U14099 ( .C1(n14388), .C2(n11781), .A(n13412), .B(n11849), .ZN(
        n13541) );
  INV_X1 U14100 ( .A(n14388), .ZN(n11650) );
  INV_X1 U14101 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11756) );
  OAI22_X1 U14102 ( .A1(n11650), .A2(n13443), .B1(n11756), .B2(n13432), .ZN(
        n11651) );
  AOI21_X1 U14103 ( .B1(n13541), .B2(n13455), .A(n11651), .ZN(n11663) );
  NAND2_X1 U14104 ( .A1(n13546), .A2(n11659), .ZN(n11653) );
  NAND2_X1 U14105 ( .A1(n11654), .A2(n11653), .ZN(n11655) );
  AOI21_X1 U14106 ( .B1(n11655), .B2(n11656), .A(n13430), .ZN(n11660) );
  INV_X1 U14107 ( .A(n11655), .ZN(n11658) );
  INV_X1 U14108 ( .A(n13187), .ZN(n11974) );
  OAI22_X1 U14109 ( .A1(n11974), .A2(n13144), .B1(n11659), .B2(n13142), .ZN(
        n14387) );
  AOI21_X1 U14110 ( .B1(n11660), .B2(n11842), .A(n14387), .ZN(n13542) );
  OAI21_X1 U14111 ( .B1(n14391), .B2(n13385), .A(n13542), .ZN(n11661) );
  NAND2_X1 U14112 ( .A1(n11661), .A2(n13432), .ZN(n11662) );
  OAI211_X1 U14113 ( .C1(n13544), .C2(n13449), .A(n11663), .B(n11662), .ZN(
        P2_U3249) );
  NAND2_X1 U14114 ( .A1(n11665), .A2(n11664), .ZN(n11667) );
  NAND2_X1 U14115 ( .A1(n14443), .A2(n13744), .ZN(n11666) );
  NAND2_X1 U14116 ( .A1(n11667), .A2(n11666), .ZN(n11710) );
  XOR2_X1 U14117 ( .A(n11711), .B(n11710), .Z(n11670) );
  OR2_X1 U14118 ( .A1(n12057), .A2(n14562), .ZN(n11669) );
  OR2_X1 U14119 ( .A1(n12038), .A2(n14542), .ZN(n11668) );
  NAND2_X1 U14120 ( .A1(n11669), .A2(n11668), .ZN(n14415) );
  AOI21_X1 U14121 ( .B1(n11670), .B2(n14549), .A(n14415), .ZN(n11704) );
  AOI21_X1 U14122 ( .B1(n11711), .B2(n11674), .A(n11716), .ZN(n11675) );
  INV_X1 U14123 ( .A(n11675), .ZN(n11705) );
  OAI22_X1 U14124 ( .A1(n14576), .A2(n11676), .B1(n14418), .B2(n14526), .ZN(
        n11677) );
  AOI21_X1 U14125 ( .B1(n14411), .B2(n14550), .A(n11677), .ZN(n11681) );
  AOI21_X1 U14126 ( .B1(n14411), .B2(n11678), .A(n14058), .ZN(n11679) );
  AND2_X1 U14127 ( .A1(n11679), .A2(n11717), .ZN(n11702) );
  NAND2_X1 U14128 ( .A1(n11702), .A2(n14558), .ZN(n11680) );
  OAI211_X1 U14129 ( .C1(n11705), .C2(n14536), .A(n11681), .B(n11680), .ZN(
        n11682) );
  INV_X1 U14130 ( .A(n11682), .ZN(n11683) );
  OAI21_X1 U14131 ( .B1(n14578), .B2(n11704), .A(n11683), .ZN(P1_U3279) );
  OAI211_X1 U14132 ( .C1(n12274), .C2(n11685), .A(n11684), .B(n12878), .ZN(
        n11687) );
  AOI22_X1 U14133 ( .A1(n12511), .A2(n12846), .B1(n12847), .B2(n12513), .ZN(
        n11686) );
  INV_X1 U14134 ( .A(n12274), .ZN(n11688) );
  XNOR2_X1 U14135 ( .A(n12893), .B(n11688), .ZN(n15000) );
  NAND2_X1 U14136 ( .A1(n12275), .A2(n12979), .ZN(n15002) );
  NOR2_X1 U14137 ( .A1(n11689), .A2(n15002), .ZN(n11693) );
  OAI22_X1 U14138 ( .A1(n12813), .A2(n11691), .B1(n11690), .B2(n12910), .ZN(
        n11692) );
  AOI211_X1 U14139 ( .C1(n15000), .C2(n12888), .A(n11693), .B(n11692), .ZN(
        n11694) );
  OAI21_X1 U14140 ( .B1(n15003), .B2(n12891), .A(n11694), .ZN(P3_U3223) );
  OAI22_X1 U14141 ( .A1(n12870), .A2(n11696), .B1(n11695), .B2(n12910), .ZN(
        n11699) );
  MUX2_X1 U14142 ( .A(n11697), .B(P3_REG2_REG_7__SCAN_IN), .S(n12786), .Z(
        n11698) );
  AOI211_X1 U14143 ( .C1(n12888), .C2(n11700), .A(n11699), .B(n11698), .ZN(
        n11701) );
  INV_X1 U14144 ( .A(n11701), .ZN(P3_U3226) );
  AOI21_X1 U14145 ( .B1(n14411), .B2(n14606), .A(n11702), .ZN(n11703) );
  OAI211_X1 U14146 ( .C1(n11705), .C2(n14581), .A(n11704), .B(n11703), .ZN(
        n11707) );
  NAND2_X1 U14147 ( .A1(n11707), .A2(n14657), .ZN(n11706) );
  OAI21_X1 U14148 ( .B1(n14657), .B2(n9322), .A(n11706), .ZN(P1_U3542) );
  INV_X1 U14149 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11709) );
  NAND2_X1 U14150 ( .A1(n11707), .A2(n14646), .ZN(n11708) );
  OAI21_X1 U14151 ( .B1(n14646), .B2(n11709), .A(n11708), .ZN(P1_U3501) );
  NAND2_X1 U14152 ( .A1(n11711), .A2(n11710), .ZN(n11713) );
  NAND2_X1 U14153 ( .A1(n11713), .A2(n11712), .ZN(n11737) );
  XNOR2_X1 U14154 ( .A(n11733), .B(n11737), .ZN(n11714) );
  AOI222_X1 U14155 ( .A1(n14549), .A2(n11714), .B1(n14032), .B2(n14055), .C1(
        n13743), .C2(n14033), .ZN(n14438) );
  XNOR2_X1 U14156 ( .A(n11734), .B(n11733), .ZN(n14441) );
  INV_X1 U14157 ( .A(n11717), .ZN(n11718) );
  OAI211_X1 U14158 ( .C1(n14439), .C2(n11718), .A(n14556), .B(n11742), .ZN(
        n14437) );
  AOI22_X1 U14159 ( .A1(n14578), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n13734), 
        .B2(n14574), .ZN(n11720) );
  NAND2_X1 U14160 ( .A1(n12053), .A2(n14550), .ZN(n11719) );
  OAI211_X1 U14161 ( .C1(n14437), .C2(n13947), .A(n11720), .B(n11719), .ZN(
        n11721) );
  AOI21_X1 U14162 ( .B1(n14441), .B2(n14571), .A(n11721), .ZN(n11722) );
  OAI21_X1 U14163 ( .B1(n14578), .B2(n14438), .A(n11722), .ZN(P1_U3278) );
  XNOR2_X1 U14164 ( .A(n11723), .B(n12875), .ZN(n11724) );
  XNOR2_X1 U14165 ( .A(n6620), .B(n11724), .ZN(n11731) );
  INV_X1 U14166 ( .A(n11725), .ZN(n12867) );
  OR2_X1 U14167 ( .A1(n12491), .A2(n12862), .ZN(n11726) );
  OAI211_X1 U14168 ( .C1(n12479), .C2(n12907), .A(n11727), .B(n11726), .ZN(
        n11729) );
  NOR2_X1 U14169 ( .A1(n13052), .A2(n12485), .ZN(n11728) );
  AOI211_X1 U14170 ( .C1(n12867), .C2(n12482), .A(n11729), .B(n11728), .ZN(
        n11730) );
  OAI21_X1 U14171 ( .B1(n11731), .B2(n12499), .A(n11730), .ZN(P3_U3174) );
  INV_X1 U14172 ( .A(n12057), .ZN(n11732) );
  INV_X1 U14173 ( .A(n11740), .ZN(n11741) );
  AOI21_X1 U14174 ( .B1(n11735), .B2(n11741), .A(n11896), .ZN(n14156) );
  NAND2_X1 U14175 ( .A1(n11737), .A2(n11736), .ZN(n11739) );
  OAI21_X1 U14176 ( .B1(n6605), .B2(n11741), .A(n11883), .ZN(n14154) );
  NAND2_X1 U14177 ( .A1(n14152), .A2(n11743), .ZN(n14037) );
  OAI211_X1 U14178 ( .C1(n14152), .C2(n11743), .A(n14556), .B(n14037), .ZN(
        n14151) );
  INV_X1 U14179 ( .A(n14013), .ZN(n13700) );
  OAI22_X1 U14180 ( .A1(n13700), .A2(n14562), .B1(n12057), .B2(n14542), .ZN(
        n13641) );
  INV_X1 U14181 ( .A(n13641), .ZN(n14150) );
  OAI22_X1 U14182 ( .A1(n14578), .A2(n14150), .B1(n13644), .B2(n14526), .ZN(
        n11745) );
  NOR2_X1 U14183 ( .A1(n14152), .A2(n14530), .ZN(n11744) );
  AOI211_X1 U14184 ( .C1(n14578), .C2(P1_REG2_REG_16__SCAN_IN), .A(n11745), 
        .B(n11744), .ZN(n11746) );
  OAI21_X1 U14185 ( .B1(n13947), .B2(n14151), .A(n11746), .ZN(n11747) );
  AOI21_X1 U14186 ( .B1(n14570), .B2(n14154), .A(n11747), .ZN(n11748) );
  OAI21_X1 U14187 ( .B1(n14156), .B2(n14536), .A(n11748), .ZN(P1_U3277) );
  INV_X1 U14188 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11757) );
  NOR2_X1 U14189 ( .A1(n11768), .A2(n11757), .ZN(n11749) );
  AOI21_X1 U14190 ( .B1(n11757), .B2(n11768), .A(n11749), .ZN(n14781) );
  XNOR2_X1 U14191 ( .A(n13236), .B(n11756), .ZN(n13234) );
  NAND2_X1 U14192 ( .A1(n11751), .A2(n11750), .ZN(n11753) );
  NAND2_X1 U14193 ( .A1(n11753), .A2(n11752), .ZN(n11754) );
  NAND2_X1 U14194 ( .A1(n14765), .A2(n11754), .ZN(n11755) );
  XOR2_X1 U14195 ( .A(n14765), .B(n11754), .Z(n14767) );
  NAND2_X1 U14196 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14767), .ZN(n14766) );
  NAND2_X1 U14197 ( .A1(n11755), .A2(n14766), .ZN(n13235) );
  NAND2_X1 U14198 ( .A1(n13234), .A2(n13235), .ZN(n13233) );
  OAI21_X1 U14199 ( .B1(n11766), .B2(n11756), .A(n13233), .ZN(n14780) );
  NAND2_X1 U14200 ( .A1(n14781), .A2(n14780), .ZN(n14779) );
  XNOR2_X1 U14201 ( .A(n13249), .B(n13244), .ZN(n11758) );
  NOR2_X1 U14202 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n11758), .ZN(n13245) );
  AOI21_X1 U14203 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n11758), .A(n13245), 
        .ZN(n11774) );
  INV_X1 U14204 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n14305) );
  NAND2_X1 U14205 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13157)
         );
  XNOR2_X1 U14206 ( .A(n11768), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14785) );
  INV_X1 U14207 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11765) );
  XNOR2_X1 U14208 ( .A(n11766), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n13238) );
  OAI21_X1 U14209 ( .B1(n11761), .B2(n11760), .A(n11759), .ZN(n11762) );
  NAND2_X1 U14210 ( .A1(n14765), .A2(n11762), .ZN(n11764) );
  XNOR2_X1 U14211 ( .A(n11763), .B(n11762), .ZN(n14769) );
  NAND2_X1 U14212 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14769), .ZN(n14768) );
  NAND2_X1 U14213 ( .A1(n11764), .A2(n14768), .ZN(n13239) );
  NAND2_X1 U14214 ( .A1(n13238), .A2(n13239), .ZN(n13237) );
  OAI21_X1 U14215 ( .B1(n11766), .B2(n11765), .A(n13237), .ZN(n14784) );
  NAND2_X1 U14216 ( .A1(n14785), .A2(n14784), .ZN(n14782) );
  OAI21_X1 U14217 ( .B1(n11768), .B2(n11767), .A(n14782), .ZN(n13248) );
  XNOR2_X1 U14218 ( .A(n11769), .B(n13248), .ZN(n11770) );
  NAND2_X1 U14219 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n11770), .ZN(n13251) );
  OAI211_X1 U14220 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n11770), .A(n14783), 
        .B(n13251), .ZN(n11771) );
  OAI211_X1 U14221 ( .C1(n14305), .C2(n14752), .A(n13157), .B(n11771), .ZN(
        n11772) );
  AOI21_X1 U14222 ( .B1(n14776), .B2(n13249), .A(n11772), .ZN(n11773) );
  OAI21_X1 U14223 ( .B1(n11774), .B2(n14713), .A(n11773), .ZN(P2_U3232) );
  INV_X1 U14224 ( .A(n11775), .ZN(n11856) );
  OAI222_X1 U14225 ( .A1(n13593), .A2(n11777), .B1(n13587), .B2(n11856), .C1(
        n11776), .C2(P2_U3088), .ZN(P2_U3303) );
  XNOR2_X1 U14226 ( .A(n7079), .B(n11778), .ZN(n11780) );
  OAI22_X1 U14227 ( .A1(n11840), .A2(n13144), .B1(n11779), .B2(n13142), .ZN(
        n11817) );
  AOI21_X1 U14228 ( .B1(n11780), .B2(n13437), .A(n11817), .ZN(n13547) );
  INV_X1 U14229 ( .A(n11781), .ZN(n11782) );
  AOI211_X1 U14230 ( .C1(n13546), .C2(n11783), .A(n13412), .B(n11782), .ZN(
        n13545) );
  INV_X1 U14231 ( .A(n11819), .ZN(n11784) );
  AOI22_X1 U14232 ( .A1(n13453), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11784), 
        .B2(n13458), .ZN(n11785) );
  OAI21_X1 U14233 ( .B1(n11648), .B2(n13443), .A(n11785), .ZN(n11790) );
  INV_X1 U14234 ( .A(n11786), .ZN(n11787) );
  AOI21_X1 U14235 ( .B1(n7079), .B2(n11788), .A(n11787), .ZN(n13549) );
  NOR2_X1 U14236 ( .A1(n13549), .A2(n13449), .ZN(n11789) );
  AOI211_X1 U14237 ( .C1(n13545), .C2(n13455), .A(n11790), .B(n11789), .ZN(
        n11791) );
  OAI21_X1 U14238 ( .B1(n13453), .B2(n13547), .A(n11791), .ZN(P2_U3250) );
  NAND2_X1 U14239 ( .A1(n14431), .A2(n12146), .ZN(n11793) );
  NAND2_X1 U14240 ( .A1(n13746), .A2(n10630), .ZN(n11792) );
  NAND2_X1 U14241 ( .A1(n11793), .A2(n11792), .ZN(n11794) );
  XNOR2_X1 U14242 ( .A(n11794), .B(n12141), .ZN(n11801) );
  AND2_X1 U14243 ( .A1(n12147), .A2(n13746), .ZN(n11795) );
  AOI21_X1 U14244 ( .B1(n14431), .B2(n10630), .A(n11795), .ZN(n11802) );
  XNOR2_X1 U14245 ( .A(n11801), .B(n11802), .ZN(n14423) );
  INV_X1 U14246 ( .A(n11796), .ZN(n11797) );
  NAND2_X1 U14247 ( .A1(n11798), .A2(n11797), .ZN(n14424) );
  AND2_X1 U14248 ( .A1(n14423), .A2(n14424), .ZN(n11799) );
  INV_X1 U14249 ( .A(n11801), .ZN(n11803) );
  NAND2_X1 U14250 ( .A1(n11803), .A2(n11802), .ZN(n11804) );
  OAI22_X1 U14251 ( .A1(n11816), .A2(n12107), .B1(n14421), .B2(n12106), .ZN(
        n11805) );
  XNOR2_X1 U14252 ( .A(n11805), .B(n12141), .ZN(n12035) );
  OAI22_X1 U14253 ( .A1(n11816), .A2(n12106), .B1(n14421), .B2(n12105), .ZN(
        n12034) );
  XNOR2_X1 U14254 ( .A(n12035), .B(n12034), .ZN(n11807) );
  AOI21_X1 U14255 ( .B1(n11806), .B2(n11807), .A(n14426), .ZN(n11809) );
  INV_X1 U14256 ( .A(n11807), .ZN(n11808) );
  NAND2_X1 U14257 ( .A1(n11809), .A2(n12037), .ZN(n11815) );
  NOR2_X1 U14258 ( .A1(n14436), .A2(n11810), .ZN(n11813) );
  OAI22_X1 U14259 ( .A1(n14422), .A2(n12038), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11811), .ZN(n11812) );
  AOI211_X1 U14260 ( .C1(n13685), .C2(n13746), .A(n11813), .B(n11812), .ZN(
        n11814) );
  OAI211_X1 U14261 ( .C1(n11816), .C2(n13737), .A(n11815), .B(n11814), .ZN(
        P1_U3224) );
  AOI22_X1 U14262 ( .A1(n14386), .A2(n11817), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11818) );
  OAI21_X1 U14263 ( .B1(n14672), .B2(n11819), .A(n11818), .ZN(n11837) );
  XNOR2_X1 U14264 ( .A(n14670), .B(n11963), .ZN(n11820) );
  AND2_X1 U14265 ( .A1(n13191), .A2(n13412), .ZN(n11821) );
  NAND2_X1 U14266 ( .A1(n11820), .A2(n11821), .ZN(n11830) );
  INV_X1 U14267 ( .A(n11820), .ZN(n11823) );
  INV_X1 U14268 ( .A(n11821), .ZN(n11822) );
  NAND2_X1 U14269 ( .A1(n11823), .A2(n11822), .ZN(n11824) );
  NAND2_X1 U14270 ( .A1(n11830), .A2(n11824), .ZN(n14666) );
  INV_X1 U14271 ( .A(n14666), .ZN(n11827) );
  NAND2_X1 U14272 ( .A1(n11826), .A2(n11825), .ZN(n14661) );
  AND2_X1 U14273 ( .A1(n11827), .A2(n14661), .ZN(n11828) );
  XNOR2_X1 U14274 ( .A(n14377), .B(n11963), .ZN(n11831) );
  NAND2_X1 U14275 ( .A1(n13190), .A2(n13412), .ZN(n11832) );
  XNOR2_X1 U14276 ( .A(n11831), .B(n11832), .ZN(n14373) );
  INV_X1 U14277 ( .A(n11831), .ZN(n11833) );
  XOR2_X1 U14278 ( .A(n11963), .B(n13546), .Z(n11924) );
  NAND2_X1 U14279 ( .A1(n13189), .A2(n13412), .ZN(n11834) );
  AOI211_X1 U14280 ( .C1(n11835), .C2(n11834), .A(n14664), .B(n11925), .ZN(
        n11836) );
  AOI211_X1 U14281 ( .C1(n13546), .C2(n14669), .A(n11837), .B(n11836), .ZN(
        n11838) );
  INV_X1 U14282 ( .A(n11838), .ZN(P2_U3213) );
  OR2_X1 U14283 ( .A1(n14388), .A2(n11840), .ZN(n11841) );
  XNOR2_X1 U14284 ( .A(n11846), .B(n11976), .ZN(n11844) );
  AOI22_X1 U14285 ( .A1(n13186), .A2(n13167), .B1(n13166), .B2(n13188), .ZN(
        n13118) );
  INV_X1 U14286 ( .A(n13118), .ZN(n11843) );
  AOI21_X1 U14287 ( .B1(n11844), .B2(n13437), .A(n11843), .ZN(n13539) );
  NAND2_X1 U14288 ( .A1(n11847), .A2(n11846), .ZN(n11997) );
  OAI21_X1 U14289 ( .B1(n11847), .B2(n11846), .A(n11997), .ZN(n13540) );
  OAI22_X1 U14290 ( .A1(n13432), .A2(n11757), .B1(n13116), .B2(n13385), .ZN(
        n11848) );
  AOI21_X1 U14291 ( .B1(n13537), .B2(n13460), .A(n11848), .ZN(n11853) );
  INV_X1 U14292 ( .A(n13537), .ZN(n13123) );
  OR2_X1 U14293 ( .A1(n13123), .A2(n11849), .ZN(n11851) );
  AND3_X1 U14294 ( .A1(n13440), .A2(n11851), .A3(n11850), .ZN(n13536) );
  NAND2_X1 U14295 ( .A1(n13536), .A2(n13455), .ZN(n11852) );
  OAI211_X1 U14296 ( .C1(n13540), .C2(n13449), .A(n11853), .B(n11852), .ZN(
        n11854) );
  INV_X1 U14297 ( .A(n11854), .ZN(n11855) );
  OAI21_X1 U14298 ( .B1(n13453), .B2(n13539), .A(n11855), .ZN(P2_U3248) );
  OAI222_X1 U14299 ( .A1(P1_U3086), .A2(n11857), .B1(n14183), .B2(n11856), 
        .C1(n7163), .C2(n14180), .ZN(P1_U3331) );
  INV_X1 U14300 ( .A(n11858), .ZN(n11862) );
  OAI222_X1 U14301 ( .A1(P1_U3086), .A2(n11860), .B1(n14183), .B2(n11862), 
        .C1(n11859), .C2(n14180), .ZN(P1_U3330) );
  OAI222_X1 U14302 ( .A1(n13593), .A2(n11863), .B1(n13587), .B2(n11862), .C1(
        n11861), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U14303 ( .A(n11864), .ZN(n13583) );
  OAI222_X1 U14304 ( .A1(P1_U3086), .A2(n11865), .B1(n14183), .B2(n13583), 
        .C1(n12163), .C2(n14180), .ZN(P1_U3326) );
  INV_X1 U14305 ( .A(n11866), .ZN(n11868) );
  OAI222_X1 U14306 ( .A1(n13070), .A2(n11869), .B1(n13067), .B2(n11868), .C1(
        n11867), .C2(P3_U3151), .ZN(P3_U3266) );
  AOI21_X1 U14307 ( .B1(n11871), .B2(n11870), .A(n14519), .ZN(n11873) );
  NAND2_X1 U14308 ( .A1(n11873), .A2(n11872), .ZN(n11880) );
  NAND2_X1 U14309 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n13682)
         );
  OAI211_X1 U14310 ( .C1(n11876), .C2(n11875), .A(n14490), .B(n11874), .ZN(
        n11877) );
  NAND2_X1 U14311 ( .A1(n13682), .A2(n11877), .ZN(n11878) );
  AOI21_X1 U14312 ( .B1(n14494), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11878), 
        .ZN(n11879) );
  OAI211_X1 U14313 ( .C1(n14521), .C2(n11881), .A(n11880), .B(n11879), .ZN(
        P1_U3256) );
  INV_X1 U14314 ( .A(n13741), .ZN(n11887) );
  INV_X1 U14315 ( .A(n13954), .ZN(n11886) );
  OR2_X1 U14316 ( .A1(n14152), .A2(n14032), .ZN(n11882) );
  INV_X1 U14317 ( .A(n14028), .ZN(n14031) );
  OR2_X1 U14318 ( .A1(n14147), .A2(n13700), .ZN(n11884) );
  INV_X1 U14319 ( .A(n14141), .ZN(n11899) );
  INV_X1 U14320 ( .A(n13982), .ZN(n13980) );
  INV_X1 U14321 ( .A(n13975), .ZN(n11902) );
  INV_X1 U14322 ( .A(n13963), .ZN(n14115) );
  INV_X1 U14323 ( .A(n13935), .ZN(n13936) );
  OAI21_X1 U14324 ( .B1(n11887), .B2(n14102), .A(n13917), .ZN(n13911) );
  INV_X1 U14325 ( .A(n14095), .ZN(n11904) );
  INV_X1 U14326 ( .A(n13883), .ZN(n13886) );
  OR2_X1 U14327 ( .A1(n11890), .A2(n11906), .ZN(n11891) );
  NAND2_X1 U14328 ( .A1(n13739), .A2(n14055), .ZN(n11893) );
  NAND2_X1 U14329 ( .A1(n13740), .A2(n14033), .ZN(n11892) );
  AOI21_X2 U14330 ( .B1(n11895), .B2(n14549), .A(n11894), .ZN(n14081) );
  INV_X1 U14331 ( .A(n14034), .ZN(n13654) );
  NAND2_X1 U14332 ( .A1(n14008), .A2(n11900), .ZN(n11901) );
  INV_X1 U14333 ( .A(n14130), .ZN(n13677) );
  OAI22_X2 U14334 ( .A1(n13966), .A2(n11902), .B1(n13953), .B2(n14121), .ZN(
        n13957) );
  INV_X1 U14335 ( .A(n13918), .ZN(n13915) );
  AND2_X2 U14336 ( .A1(n13914), .A2(n11903), .ZN(n13900) );
  INV_X1 U14337 ( .A(n13920), .ZN(n13720) );
  NAND2_X1 U14338 ( .A1(n11907), .A2(n7190), .ZN(n13850) );
  OAI21_X1 U14339 ( .B1(n11907), .B2(n7190), .A(n13850), .ZN(n14082) );
  INV_X1 U14340 ( .A(n14082), .ZN(n11913) );
  AND2_X2 U14341 ( .A1(n13986), .A2(n13973), .ZN(n13967) );
  AND2_X2 U14342 ( .A1(n13967), .A2(n13963), .ZN(n13958) );
  INV_X1 U14343 ( .A(n14108), .ZN(n13942) );
  INV_X1 U14344 ( .A(n14089), .ZN(n13892) );
  OR2_X2 U14345 ( .A1(n13894), .A2(n14084), .ZN(n13876) );
  NOR2_X2 U14346 ( .A1(n14079), .A2(n13876), .ZN(n13854) );
  AND2_X1 U14347 ( .A1(n14079), .A2(n13876), .ZN(n11908) );
  OAI22_X1 U14348 ( .A1(n14576), .A2(n11909), .B1(n12155), .B2(n14526), .ZN(
        n11910) );
  AOI21_X1 U14349 ( .B1(n14079), .B2(n14550), .A(n11910), .ZN(n11911) );
  OAI21_X1 U14350 ( .B1(n14077), .B2(n13947), .A(n11911), .ZN(n11912) );
  AOI21_X1 U14351 ( .B1(n11913), .B2(n14571), .A(n11912), .ZN(n11914) );
  OAI21_X1 U14352 ( .B1(n14578), .B2(n14081), .A(n11914), .ZN(P1_U3265) );
  AOI22_X1 U14353 ( .A1(n14386), .A2(n11916), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n11915), .ZN(n11922) );
  OAI21_X1 U14354 ( .B1(n11919), .B2(n11918), .A(n11917), .ZN(n11920) );
  NAND2_X1 U14355 ( .A1(n14384), .A2(n11920), .ZN(n11921) );
  OAI211_X1 U14356 ( .C1(n13162), .C2(n7048), .A(n11922), .B(n11921), .ZN(
        P2_U3209) );
  XNOR2_X1 U14357 ( .A(n13532), .B(n11963), .ZN(n11933) );
  NAND2_X1 U14358 ( .A1(n13186), .A2(n13412), .ZN(n11934) );
  INV_X1 U14359 ( .A(n11923), .ZN(n11927) );
  INV_X1 U14360 ( .A(n11924), .ZN(n11926) );
  XNOR2_X1 U14361 ( .A(n14388), .B(n11963), .ZN(n11928) );
  NAND2_X1 U14362 ( .A1(n13188), .A2(n13412), .ZN(n11929) );
  XNOR2_X1 U14363 ( .A(n11928), .B(n11929), .ZN(n14382) );
  INV_X1 U14364 ( .A(n11928), .ZN(n11930) );
  NAND2_X1 U14365 ( .A1(n11930), .A2(n11929), .ZN(n13112) );
  XNOR2_X1 U14366 ( .A(n13537), .B(n6487), .ZN(n11932) );
  NAND2_X1 U14367 ( .A1(n13187), .A2(n13412), .ZN(n11931) );
  XNOR2_X1 U14368 ( .A(n11932), .B(n11931), .ZN(n13113) );
  XNOR2_X1 U14369 ( .A(n11933), .B(n11934), .ZN(n13154) );
  XNOR2_X1 U14370 ( .A(n13528), .B(n6488), .ZN(n11936) );
  NAND2_X1 U14371 ( .A1(n13185), .A2(n13412), .ZN(n11935) );
  NAND2_X1 U14372 ( .A1(n11936), .A2(n11935), .ZN(n13087) );
  NOR2_X1 U14373 ( .A1(n11936), .A2(n11935), .ZN(n13089) );
  XNOR2_X1 U14374 ( .A(n13523), .B(n11963), .ZN(n11938) );
  AND2_X1 U14375 ( .A1(n13184), .A2(n13412), .ZN(n11937) );
  NAND2_X1 U14376 ( .A1(n11938), .A2(n11937), .ZN(n13134) );
  XNOR2_X1 U14377 ( .A(n13518), .B(n11963), .ZN(n11939) );
  NAND2_X1 U14378 ( .A1(n13183), .A2(n13412), .ZN(n11940) );
  XNOR2_X1 U14379 ( .A(n11939), .B(n11940), .ZN(n13097) );
  INV_X1 U14380 ( .A(n11940), .ZN(n11941) );
  NAND2_X1 U14381 ( .A1(n11939), .A2(n11941), .ZN(n11942) );
  XNOR2_X1 U14382 ( .A(n13511), .B(n11963), .ZN(n11943) );
  NAND2_X1 U14383 ( .A1(n13182), .A2(n13412), .ZN(n13148) );
  NOR2_X1 U14384 ( .A1(n13147), .A2(n7425), .ZN(n11947) );
  XNOR2_X1 U14385 ( .A(n13505), .B(n11963), .ZN(n11945) );
  XNOR2_X1 U14386 ( .A(n11947), .B(n11945), .ZN(n13079) );
  NAND2_X1 U14387 ( .A1(n13181), .A2(n13412), .ZN(n13080) );
  INV_X1 U14388 ( .A(n11945), .ZN(n11946) );
  XNOR2_X1 U14389 ( .A(n13496), .B(n6487), .ZN(n11949) );
  NAND2_X1 U14390 ( .A1(n13180), .A2(n13412), .ZN(n11948) );
  NOR2_X1 U14391 ( .A1(n11949), .A2(n11948), .ZN(n11950) );
  AOI21_X1 U14392 ( .B1(n11949), .B2(n11948), .A(n11950), .ZN(n13125) );
  INV_X1 U14393 ( .A(n11950), .ZN(n11951) );
  XNOR2_X1 U14394 ( .A(n13335), .B(n6488), .ZN(n11953) );
  NAND2_X1 U14395 ( .A1(n13179), .A2(n13412), .ZN(n11952) );
  NOR2_X1 U14396 ( .A1(n11953), .A2(n11952), .ZN(n11954) );
  AOI21_X1 U14397 ( .B1(n11953), .B2(n11952), .A(n11954), .ZN(n13105) );
  INV_X1 U14398 ( .A(n11954), .ZN(n11955) );
  NAND2_X1 U14399 ( .A1(n13178), .A2(n13412), .ZN(n11956) );
  XNOR2_X1 U14400 ( .A(n13487), .B(n11963), .ZN(n11958) );
  XOR2_X1 U14401 ( .A(n11956), .B(n11958), .Z(n13165) );
  INV_X1 U14402 ( .A(n11956), .ZN(n11957) );
  NOR2_X1 U14403 ( .A1(n11958), .A2(n11957), .ZN(n11959) );
  XNOR2_X1 U14404 ( .A(n13304), .B(n6487), .ZN(n11961) );
  NAND2_X1 U14405 ( .A1(n13177), .A2(n13412), .ZN(n11960) );
  NOR2_X1 U14406 ( .A1(n11961), .A2(n11960), .ZN(n11962) );
  AOI21_X1 U14407 ( .B1(n11961), .B2(n11960), .A(n11962), .ZN(n13072) );
  NAND2_X1 U14408 ( .A1(n13176), .A2(n13412), .ZN(n11964) );
  XNOR2_X1 U14409 ( .A(n11964), .B(n11963), .ZN(n11965) );
  XNOR2_X1 U14410 ( .A(n13475), .B(n11965), .ZN(n11966) );
  XNOR2_X1 U14411 ( .A(n11967), .B(n11966), .ZN(n11973) );
  NAND2_X1 U14412 ( .A1(n13175), .A2(n13167), .ZN(n11969) );
  NAND2_X1 U14413 ( .A1(n13177), .A2(n13166), .ZN(n11968) );
  NAND2_X1 U14414 ( .A1(n11969), .A2(n11968), .ZN(n13279) );
  AOI22_X1 U14415 ( .A1(n14386), .A2(n13279), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11970) );
  OAI21_X1 U14416 ( .B1(n14672), .B2(n13285), .A(n11970), .ZN(n11971) );
  AOI21_X1 U14417 ( .B1(n13475), .B2(n14669), .A(n11971), .ZN(n11972) );
  OAI21_X1 U14418 ( .B1(n11973), .B2(n14664), .A(n11972), .ZN(P2_U3192) );
  INV_X1 U14419 ( .A(n13496), .ZN(n13133) );
  NAND2_X1 U14420 ( .A1(n13537), .A2(n11974), .ZN(n11975) );
  INV_X1 U14421 ( .A(n13186), .ZN(n11978) );
  OR2_X1 U14422 ( .A1(n13532), .A2(n11978), .ZN(n11977) );
  NAND2_X1 U14423 ( .A1(n13532), .A2(n11978), .ZN(n11979) );
  NAND2_X1 U14424 ( .A1(n11980), .A2(n11979), .ZN(n13428) );
  NAND2_X1 U14425 ( .A1(n13428), .A2(n13427), .ZN(n11982) );
  INV_X1 U14426 ( .A(n13185), .ZN(n11999) );
  NAND2_X1 U14427 ( .A1(n13528), .A2(n11999), .ZN(n11981) );
  AND2_X1 U14428 ( .A1(n13523), .A2(n11983), .ZN(n11984) );
  NAND2_X1 U14429 ( .A1(n13378), .A2(n13383), .ZN(n11987) );
  NAND2_X1 U14430 ( .A1(n13511), .A2(n13082), .ZN(n11986) );
  OR2_X1 U14431 ( .A1(n13505), .A2(n13145), .ZN(n11988) );
  INV_X1 U14432 ( .A(n13340), .ZN(n13344) );
  INV_X1 U14433 ( .A(n13179), .ZN(n11989) );
  NOR2_X1 U14434 ( .A1(n13483), .A2(n13177), .ZN(n13278) );
  NAND2_X1 U14435 ( .A1(n13176), .A2(n13166), .ZN(n11993) );
  AOI21_X1 U14436 ( .B1(n11991), .B2(P2_B_REG_SCAN_IN), .A(n13144), .ZN(n13266) );
  NAND2_X1 U14437 ( .A1(n13266), .A2(n13174), .ZN(n11992) );
  INV_X1 U14438 ( .A(n13177), .ZN(n12009) );
  NAND2_X1 U14439 ( .A1(n13537), .A2(n13187), .ZN(n11996) );
  NAND2_X1 U14440 ( .A1(n11997), .A2(n11996), .ZN(n13447) );
  OR2_X1 U14441 ( .A1(n13532), .A2(n13186), .ZN(n11998) );
  INV_X1 U14442 ( .A(n13528), .ZN(n13425) );
  AND2_X1 U14443 ( .A1(n13523), .A2(n13184), .ZN(n12000) );
  OR2_X1 U14444 ( .A1(n13523), .A2(n13184), .ZN(n12001) );
  NAND2_X1 U14445 ( .A1(n12002), .A2(n12001), .ZN(n13394) );
  OR2_X1 U14446 ( .A1(n13183), .A2(n13518), .ZN(n12003) );
  NAND2_X1 U14447 ( .A1(n13511), .A2(n13182), .ZN(n12004) );
  NAND2_X1 U14448 ( .A1(n13367), .A2(n6976), .ZN(n13366) );
  OR2_X1 U14449 ( .A1(n13505), .A2(n13181), .ZN(n12005) );
  OAI21_X1 U14450 ( .B1(n13179), .B2(n13335), .A(n13328), .ZN(n13309) );
  INV_X1 U14451 ( .A(n13487), .ZN(n13312) );
  NAND2_X1 U14452 ( .A1(n13282), .A2(n12010), .ZN(n12011) );
  INV_X1 U14453 ( .A(n13511), .ZN(n13382) );
  NAND2_X1 U14454 ( .A1(n13399), .A2(n13382), .ZN(n13381) );
  OR2_X1 U14455 ( .A1(n13381), .A2(n13505), .ZN(n13372) );
  OR2_X2 U14456 ( .A1(n13288), .A2(n13471), .ZN(n13270) );
  AOI21_X1 U14457 ( .B1(n13471), .B2(n13288), .A(n13412), .ZN(n12015) );
  INV_X1 U14458 ( .A(n13471), .ZN(n12019) );
  INV_X1 U14459 ( .A(n12016), .ZN(n12017) );
  AOI22_X1 U14460 ( .A1(n13453), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n12017), 
        .B2(n13458), .ZN(n12018) );
  OAI21_X1 U14461 ( .B1(n12019), .B2(n13443), .A(n12018), .ZN(n12020) );
  OAI21_X1 U14462 ( .B1(n13472), .B2(n13453), .A(n12023), .ZN(P2_U3236) );
  OAI21_X1 U14463 ( .B1(n12026), .B2(n12025), .A(n12024), .ZN(n12027) );
  NAND2_X1 U14464 ( .A1(n12027), .A2(n14412), .ZN(n12031) );
  AOI22_X1 U14465 ( .A1(n12029), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n14414), 
        .B2(n12028), .ZN(n12030) );
  OAI211_X1 U14466 ( .C1(n14595), .C2(n13737), .A(n12031), .B(n12030), .ZN(
        P1_U3237) );
  INV_X1 U14467 ( .A(n12032), .ZN(n13588) );
  OAI222_X1 U14468 ( .A1(n9665), .A2(P1_U3086), .B1(n14183), .B2(n13588), .C1(
        n12033), .C2(n14180), .ZN(P1_U3327) );
  NAND2_X1 U14469 ( .A1(n12035), .A2(n12034), .ZN(n12036) );
  OAI22_X1 U14470 ( .A1(n14443), .A2(n12106), .B1(n12038), .B2(n12105), .ZN(
        n12046) );
  OAI22_X1 U14471 ( .A1(n14443), .A2(n12107), .B1(n12038), .B2(n12106), .ZN(
        n12039) );
  XNOR2_X1 U14472 ( .A(n12039), .B(n12141), .ZN(n12045) );
  XOR2_X1 U14473 ( .A(n12046), .B(n12045), .Z(n13680) );
  NAND2_X1 U14474 ( .A1(n14411), .A2(n12146), .ZN(n12041) );
  NAND2_X1 U14475 ( .A1(n13743), .A2(n10630), .ZN(n12040) );
  NAND2_X1 U14476 ( .A1(n12041), .A2(n12040), .ZN(n12043) );
  XNOR2_X1 U14477 ( .A(n12043), .B(n12042), .ZN(n12051) );
  AND2_X1 U14478 ( .A1(n12147), .A2(n13743), .ZN(n12044) );
  AOI21_X1 U14479 ( .B1(n14411), .B2(n10630), .A(n12044), .ZN(n12050) );
  XNOR2_X1 U14480 ( .A(n12051), .B(n12050), .ZN(n14406) );
  INV_X1 U14481 ( .A(n12045), .ZN(n12048) );
  INV_X1 U14482 ( .A(n12046), .ZN(n12047) );
  NOR2_X1 U14483 ( .A1(n12048), .A2(n12047), .ZN(n14407) );
  NOR2_X1 U14484 ( .A1(n14406), .A2(n14407), .ZN(n12049) );
  NAND2_X1 U14485 ( .A1(n12051), .A2(n12050), .ZN(n12052) );
  NAND2_X1 U14486 ( .A1(n14409), .A2(n12052), .ZN(n12058) );
  NAND2_X1 U14487 ( .A1(n12053), .A2(n12146), .ZN(n12055) );
  OR2_X1 U14488 ( .A1(n12057), .A2(n12106), .ZN(n12054) );
  NAND2_X1 U14489 ( .A1(n12055), .A2(n12054), .ZN(n12056) );
  XNOR2_X1 U14490 ( .A(n12056), .B(n12141), .ZN(n12059) );
  XNOR2_X1 U14491 ( .A(n12058), .B(n12059), .ZN(n13728) );
  OAI22_X1 U14492 ( .A1(n14439), .A2(n12106), .B1(n12057), .B2(n12105), .ZN(
        n13727) );
  INV_X1 U14493 ( .A(n12058), .ZN(n12060) );
  NAND2_X1 U14494 ( .A1(n12060), .A2(n12059), .ZN(n12061) );
  OAI22_X1 U14495 ( .A1(n14152), .A2(n12107), .B1(n12062), .B2(n12106), .ZN(
        n12063) );
  XNOR2_X1 U14496 ( .A(n12063), .B(n12141), .ZN(n12066) );
  OR2_X1 U14497 ( .A1(n14152), .A2(n12106), .ZN(n12065) );
  NAND2_X1 U14498 ( .A1(n12147), .A2(n14032), .ZN(n12064) );
  NAND2_X1 U14499 ( .A1(n12065), .A2(n12064), .ZN(n12067) );
  XNOR2_X1 U14500 ( .A(n12066), .B(n12067), .ZN(n13640) );
  INV_X1 U14501 ( .A(n12066), .ZN(n12069) );
  INV_X1 U14502 ( .A(n12067), .ZN(n12068) );
  NAND2_X1 U14503 ( .A1(n12069), .A2(n12068), .ZN(n12070) );
  NAND2_X1 U14504 ( .A1(n14147), .A2(n12146), .ZN(n12072) );
  NAND2_X1 U14505 ( .A1(n14013), .A2(n10630), .ZN(n12071) );
  NAND2_X1 U14506 ( .A1(n12072), .A2(n12071), .ZN(n12073) );
  XNOR2_X1 U14507 ( .A(n12073), .B(n12141), .ZN(n12074) );
  AOI22_X1 U14508 ( .A1(n14147), .A2(n10630), .B1(n12147), .B2(n14013), .ZN(
        n12075) );
  XNOR2_X1 U14509 ( .A(n12074), .B(n12075), .ZN(n13651) );
  INV_X1 U14510 ( .A(n12074), .ZN(n12076) );
  NAND2_X1 U14511 ( .A1(n12076), .A2(n12075), .ZN(n12077) );
  NAND2_X1 U14512 ( .A1(n14141), .A2(n12146), .ZN(n12079) );
  NAND2_X1 U14513 ( .A1(n14034), .A2(n10630), .ZN(n12078) );
  NAND2_X1 U14514 ( .A1(n12079), .A2(n12078), .ZN(n12080) );
  XNOR2_X1 U14515 ( .A(n12080), .B(n12141), .ZN(n12081) );
  AOI22_X1 U14516 ( .A1(n14141), .A2(n10630), .B1(n12147), .B2(n14034), .ZN(
        n12082) );
  XNOR2_X1 U14517 ( .A(n12081), .B(n12082), .ZN(n13699) );
  INV_X1 U14518 ( .A(n12081), .ZN(n12083) );
  NAND2_X1 U14519 ( .A1(n12083), .A2(n12082), .ZN(n12084) );
  AND2_X1 U14520 ( .A1(n14021), .A2(n12147), .ZN(n12085) );
  AOI21_X1 U14521 ( .B1(n14136), .B2(n10630), .A(n12085), .ZN(n12090) );
  NAND2_X1 U14522 ( .A1(n14136), .A2(n12146), .ZN(n12087) );
  NAND2_X1 U14523 ( .A1(n14021), .A2(n10630), .ZN(n12086) );
  NAND2_X1 U14524 ( .A1(n12087), .A2(n12086), .ZN(n12088) );
  XNOR2_X1 U14525 ( .A(n12088), .B(n12141), .ZN(n12092) );
  XOR2_X1 U14526 ( .A(n12090), .B(n12092), .Z(n13611) );
  INV_X1 U14527 ( .A(n12090), .ZN(n12091) );
  NAND2_X1 U14528 ( .A1(n12092), .A2(n12091), .ZN(n12093) );
  AND2_X1 U14529 ( .A1(n13998), .A2(n12147), .ZN(n12094) );
  AOI21_X1 U14530 ( .B1(n14130), .B2(n10630), .A(n12094), .ZN(n12097) );
  AOI22_X1 U14531 ( .A1(n14130), .A2(n12146), .B1(n10630), .B2(n13998), .ZN(
        n12095) );
  XNOR2_X1 U14532 ( .A(n12095), .B(n12141), .ZN(n12096) );
  XOR2_X1 U14533 ( .A(n12097), .B(n12096), .Z(n13668) );
  INV_X1 U14534 ( .A(n12096), .ZN(n12099) );
  INV_X1 U14535 ( .A(n12097), .ZN(n12098) );
  NAND2_X1 U14536 ( .A1(n12099), .A2(n12098), .ZN(n12100) );
  AOI22_X1 U14537 ( .A1(n14121), .A2(n12146), .B1(n10630), .B2(n13953), .ZN(
        n12101) );
  XNOR2_X1 U14538 ( .A(n12101), .B(n12141), .ZN(n12103) );
  AOI22_X1 U14539 ( .A1(n14121), .A2(n10630), .B1(n12147), .B2(n13953), .ZN(
        n12102) );
  XNOR2_X1 U14540 ( .A(n12103), .B(n12102), .ZN(n13621) );
  NAND2_X1 U14541 ( .A1(n12103), .A2(n12102), .ZN(n12104) );
  NAND2_X1 U14542 ( .A1(n13619), .A2(n12104), .ZN(n13689) );
  OAI22_X1 U14543 ( .A1(n13963), .A2(n12106), .B1(n13622), .B2(n12105), .ZN(
        n12109) );
  OAI22_X1 U14544 ( .A1(n13963), .A2(n12107), .B1(n13622), .B2(n12106), .ZN(
        n12108) );
  XNOR2_X1 U14545 ( .A(n12108), .B(n12141), .ZN(n12110) );
  XOR2_X1 U14546 ( .A(n12109), .B(n12110), .Z(n13690) );
  OR2_X1 U14547 ( .A1(n12110), .A2(n12109), .ZN(n12111) );
  NAND2_X1 U14548 ( .A1(n14108), .A2(n12146), .ZN(n12113) );
  NAND2_X1 U14549 ( .A1(n13954), .A2(n10630), .ZN(n12112) );
  NAND2_X1 U14550 ( .A1(n12113), .A2(n12112), .ZN(n12114) );
  XNOR2_X1 U14551 ( .A(n12114), .B(n12141), .ZN(n12115) );
  AOI22_X1 U14552 ( .A1(n14108), .A2(n10630), .B1(n12147), .B2(n13954), .ZN(
        n12116) );
  XNOR2_X1 U14553 ( .A(n12115), .B(n12116), .ZN(n13603) );
  INV_X1 U14554 ( .A(n12115), .ZN(n12117) );
  NAND2_X1 U14555 ( .A1(n14102), .A2(n12146), .ZN(n12119) );
  NAND2_X1 U14556 ( .A1(n13741), .A2(n10630), .ZN(n12118) );
  NAND2_X1 U14557 ( .A1(n12119), .A2(n12118), .ZN(n12120) );
  XNOR2_X1 U14558 ( .A(n12120), .B(n12141), .ZN(n12121) );
  AOI22_X1 U14559 ( .A1(n14102), .A2(n10630), .B1(n12147), .B2(n13741), .ZN(
        n12122) );
  XNOR2_X1 U14560 ( .A(n12121), .B(n12122), .ZN(n13661) );
  INV_X1 U14561 ( .A(n12121), .ZN(n12123) );
  NAND2_X1 U14562 ( .A1(n14095), .A2(n12146), .ZN(n12125) );
  NAND2_X1 U14563 ( .A1(n13920), .A2(n10630), .ZN(n12124) );
  NAND2_X1 U14564 ( .A1(n12125), .A2(n12124), .ZN(n12126) );
  XNOR2_X1 U14565 ( .A(n12126), .B(n12141), .ZN(n12127) );
  AOI22_X1 U14566 ( .A1(n14095), .A2(n10630), .B1(n12147), .B2(n13920), .ZN(
        n12128) );
  XNOR2_X1 U14567 ( .A(n12127), .B(n12128), .ZN(n13630) );
  NAND2_X1 U14568 ( .A1(n13629), .A2(n13630), .ZN(n12131) );
  INV_X1 U14569 ( .A(n12127), .ZN(n12129) );
  NAND2_X1 U14570 ( .A1(n12129), .A2(n12128), .ZN(n12130) );
  NAND2_X1 U14571 ( .A1(n14089), .A2(n12146), .ZN(n12133) );
  NAND2_X1 U14572 ( .A1(n13871), .A2(n10630), .ZN(n12132) );
  NAND2_X1 U14573 ( .A1(n12133), .A2(n12132), .ZN(n12134) );
  XNOR2_X1 U14574 ( .A(n12134), .B(n12141), .ZN(n12135) );
  AOI22_X1 U14575 ( .A1(n14089), .A2(n10630), .B1(n12147), .B2(n13871), .ZN(
        n12136) );
  XNOR2_X1 U14576 ( .A(n12135), .B(n12136), .ZN(n13719) );
  INV_X1 U14577 ( .A(n12135), .ZN(n12137) );
  NAND2_X1 U14578 ( .A1(n12137), .A2(n12136), .ZN(n12138) );
  NAND2_X1 U14579 ( .A1(n14084), .A2(n12146), .ZN(n12140) );
  NAND2_X1 U14580 ( .A1(n13740), .A2(n10630), .ZN(n12139) );
  NAND2_X1 U14581 ( .A1(n12140), .A2(n12139), .ZN(n12142) );
  XNOR2_X1 U14582 ( .A(n12142), .B(n12141), .ZN(n12143) );
  AOI22_X1 U14583 ( .A1(n14084), .A2(n10630), .B1(n12147), .B2(n13740), .ZN(
        n12144) );
  XNOR2_X1 U14584 ( .A(n12143), .B(n12144), .ZN(n13596) );
  INV_X1 U14585 ( .A(n12143), .ZN(n12145) );
  AOI22_X1 U14586 ( .A1(n14079), .A2(n12146), .B1(n10630), .B2(n13872), .ZN(
        n12150) );
  AOI22_X1 U14587 ( .A1(n14079), .A2(n10630), .B1(n12147), .B2(n13872), .ZN(
        n12148) );
  XNOR2_X1 U14588 ( .A(n12148), .B(n12141), .ZN(n12149) );
  XOR2_X1 U14589 ( .A(n12150), .B(n12149), .Z(n12151) );
  OAI22_X1 U14590 ( .A1(n14419), .A2(n13721), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12152), .ZN(n12153) );
  AOI21_X1 U14591 ( .B1(n13729), .B2(n13739), .A(n12153), .ZN(n12154) );
  OAI21_X1 U14592 ( .B1(n12155), .B2(n14436), .A(n12154), .ZN(n12156) );
  AOI21_X1 U14593 ( .B1(n14079), .B2(n14432), .A(n12156), .ZN(n12157) );
  OAI21_X1 U14594 ( .B1(n12158), .B2(n14426), .A(n12157), .ZN(P1_U3220) );
  INV_X1 U14595 ( .A(n12159), .ZN(n14182) );
  INV_X1 U14596 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12165) );
  INV_X1 U14597 ( .A(n12160), .ZN(n12161) );
  NAND2_X1 U14598 ( .A1(n12163), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12164) );
  NAND2_X1 U14599 ( .A1(n12165), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12167) );
  NAND2_X1 U14600 ( .A1(n14181), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12166) );
  NAND2_X1 U14601 ( .A1(n12167), .A2(n12166), .ZN(n12179) );
  OAI21_X1 U14602 ( .B1(n12180), .B2(n12179), .A(n12167), .ZN(n12169) );
  XNOR2_X1 U14603 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12168) );
  XNOR2_X1 U14604 ( .A(n12169), .B(n12168), .ZN(n13063) );
  NAND2_X1 U14605 ( .A1(n13063), .A2(n12181), .ZN(n12171) );
  NAND2_X1 U14606 ( .A1(n12182), .A2(SI_31_), .ZN(n12170) );
  INV_X1 U14607 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12635) );
  NAND2_X1 U14608 ( .A1(n12172), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12175) );
  NAND2_X1 U14609 ( .A1(n12173), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12174) );
  OAI211_X1 U14610 ( .C1(n8420), .C2(n12635), .A(n12175), .B(n12174), .ZN(
        n12176) );
  INV_X1 U14611 ( .A(n12176), .ZN(n12177) );
  XNOR2_X1 U14612 ( .A(n12180), .B(n12179), .ZN(n12371) );
  NAND2_X1 U14613 ( .A1(n12371), .A2(n12181), .ZN(n12184) );
  NAND2_X1 U14614 ( .A1(n12182), .A2(SI_30_), .ZN(n12183) );
  NAND2_X1 U14615 ( .A1(n13001), .A2(n12188), .ZN(n12185) );
  INV_X1 U14616 ( .A(n12632), .ZN(n12501) );
  OAI21_X1 U14617 ( .B1(n12638), .B2(n12501), .A(n12350), .ZN(n12186) );
  AOI211_X1 U14618 ( .C1(n12187), .C2(n12354), .A(n12356), .B(n12186), .ZN(
        n12192) );
  INV_X1 U14619 ( .A(n12188), .ZN(n12502) );
  INV_X1 U14620 ( .A(n12196), .ZN(n12215) );
  INV_X1 U14621 ( .A(n12380), .ZN(n12347) );
  INV_X1 U14622 ( .A(n12743), .ZN(n12746) );
  INV_X1 U14623 ( .A(n12833), .ZN(n12830) );
  NAND4_X1 U14624 ( .A1(n12199), .A2(n12198), .A3(n12197), .A4(n12263), .ZN(
        n12201) );
  NOR2_X1 U14625 ( .A1(n12201), .A2(n12200), .ZN(n12205) );
  NOR2_X1 U14626 ( .A1(n12274), .A2(n12202), .ZN(n12204) );
  AND4_X1 U14627 ( .A1(n12258), .A2(n12224), .A3(n12240), .A4(n12245), .ZN(
        n12203) );
  NAND4_X1 U14628 ( .A1(n12205), .A2(n12899), .A3(n12204), .A4(n12203), .ZN(
        n12208) );
  INV_X1 U14629 ( .A(n12850), .ZN(n12206) );
  NOR4_X1 U14630 ( .A1(n12830), .A2(n12208), .A3(n12207), .A4(n12866), .ZN(
        n12209) );
  NAND4_X1 U14631 ( .A1(n12789), .A2(n12852), .A3(n12821), .A4(n12209), .ZN(
        n12210) );
  NOR4_X1 U14632 ( .A1(n12746), .A2(n12211), .A3(n12779), .A4(n12210), .ZN(
        n12212) );
  INV_X1 U14633 ( .A(n12763), .ZN(n12319) );
  NAND4_X1 U14634 ( .A1(n12716), .A2(n12729), .A3(n12212), .A4(n12319), .ZN(
        n12213) );
  NOR4_X1 U14635 ( .A1(n12663), .A2(n12329), .A3(n12677), .A4(n12213), .ZN(
        n12214) );
  NAND4_X1 U14636 ( .A1(n12215), .A2(n12347), .A3(n12214), .A4(n12649), .ZN(
        n12216) );
  XNOR2_X1 U14637 ( .A(n12217), .B(n12609), .ZN(n12361) );
  NAND3_X1 U14638 ( .A1(n12523), .A2(n12219), .A3(n12218), .ZN(n12220) );
  OAI21_X1 U14639 ( .B1(n12222), .B2(n12221), .A(n12220), .ZN(n12223) );
  NAND2_X1 U14640 ( .A1(n12225), .A2(n12224), .ZN(n12235) );
  NAND2_X1 U14641 ( .A1(n12229), .A2(n12227), .ZN(n12228) );
  INV_X1 U14642 ( .A(n12229), .ZN(n12230) );
  MUX2_X1 U14643 ( .A(n12231), .B(n12230), .S(n12312), .Z(n12234) );
  AND2_X1 U14644 ( .A1(n12241), .A2(n12232), .ZN(n12233) );
  OAI22_X1 U14645 ( .A1(n12235), .A2(n12234), .B1(n12346), .B2(n12233), .ZN(
        n12239) );
  AOI21_X1 U14646 ( .B1(n12238), .B2(n12236), .A(n12312), .ZN(n12237) );
  AOI21_X1 U14647 ( .B1(n12239), .B2(n12238), .A(n12237), .ZN(n12247) );
  OAI21_X1 U14648 ( .B1(n12241), .B2(n12312), .A(n12240), .ZN(n12246) );
  MUX2_X1 U14649 ( .A(n12243), .B(n12242), .S(n12312), .Z(n12244) );
  OAI211_X1 U14650 ( .C1(n12247), .C2(n12246), .A(n12245), .B(n12244), .ZN(
        n12254) );
  NAND2_X1 U14651 ( .A1(n12256), .A2(n12248), .ZN(n12251) );
  NAND2_X1 U14652 ( .A1(n12255), .A2(n12249), .ZN(n12250) );
  MUX2_X1 U14653 ( .A(n12251), .B(n12250), .S(n12346), .Z(n12252) );
  INV_X1 U14654 ( .A(n12252), .ZN(n12253) );
  NAND2_X1 U14655 ( .A1(n12254), .A2(n12253), .ZN(n12259) );
  MUX2_X1 U14656 ( .A(n12256), .B(n12255), .S(n12312), .Z(n12257) );
  NAND3_X1 U14657 ( .A1(n12259), .A2(n12258), .A3(n12257), .ZN(n12264) );
  MUX2_X1 U14658 ( .A(n12261), .B(n12260), .S(n12346), .Z(n12262) );
  NAND3_X1 U14659 ( .A1(n12264), .A2(n12263), .A3(n12262), .ZN(n12269) );
  MUX2_X1 U14660 ( .A(n12266), .B(n12265), .S(n12312), .Z(n12267) );
  NAND3_X1 U14661 ( .A1(n12269), .A2(n12268), .A3(n12267), .ZN(n12278) );
  AND2_X1 U14662 ( .A1(n12513), .A2(n12270), .ZN(n12272) );
  NOR2_X1 U14663 ( .A1(n12513), .A2(n12270), .ZN(n12271) );
  MUX2_X1 U14664 ( .A(n12272), .B(n12271), .S(n12346), .Z(n12273) );
  NOR2_X1 U14665 ( .A1(n12274), .A2(n12273), .ZN(n12277) );
  NOR3_X1 U14666 ( .A1(n12905), .A2(n12275), .A3(n12312), .ZN(n12276) );
  AOI21_X1 U14667 ( .B1(n12278), .B2(n12277), .A(n12276), .ZN(n12283) );
  INV_X1 U14668 ( .A(n12894), .ZN(n12281) );
  NAND2_X1 U14669 ( .A1(n12863), .A2(n12279), .ZN(n12280) );
  AOI21_X1 U14670 ( .B1(n12899), .B2(n12281), .A(n12280), .ZN(n12282) );
  AOI21_X1 U14671 ( .B1(n12286), .B2(n12284), .A(n12312), .ZN(n12285) );
  NOR2_X1 U14672 ( .A1(n12863), .A2(n12312), .ZN(n12287) );
  NAND2_X1 U14673 ( .A1(n12288), .A2(n12312), .ZN(n12289) );
  AND2_X1 U14674 ( .A1(n12852), .A2(n12289), .ZN(n12293) );
  OAI211_X1 U14675 ( .C1(n12292), .C2(n12830), .A(n12291), .B(n12290), .ZN(
        n12298) );
  NAND3_X1 U14676 ( .A1(n12294), .A2(n12293), .A3(n12850), .ZN(n12296) );
  OR3_X1 U14677 ( .A1(n13046), .A2(n12509), .A3(n12312), .ZN(n12295) );
  AOI21_X1 U14678 ( .B1(n12296), .B2(n12295), .A(n12830), .ZN(n12297) );
  AOI21_X1 U14679 ( .B1(n12298), .B2(n12312), .A(n12297), .ZN(n12303) );
  INV_X1 U14680 ( .A(n12300), .ZN(n12302) );
  AND2_X1 U14681 ( .A1(n12300), .A2(n12299), .ZN(n12301) );
  OAI22_X1 U14682 ( .A1(n12303), .A2(n12302), .B1(n12301), .B2(n12312), .ZN(
        n12305) );
  OR3_X1 U14683 ( .A1(n12978), .A2(n12832), .A3(n12312), .ZN(n12304) );
  NAND2_X1 U14684 ( .A1(n12305), .A2(n12304), .ZN(n12311) );
  INV_X1 U14685 ( .A(n12794), .ZN(n12310) );
  INV_X1 U14686 ( .A(n12313), .ZN(n12309) );
  AND2_X1 U14687 ( .A1(n12306), .A2(n12346), .ZN(n12307) );
  OAI211_X1 U14688 ( .C1(n12309), .C2(n12308), .A(n12317), .B(n12307), .ZN(
        n12315) );
  NAND3_X1 U14689 ( .A1(n12316), .A2(n12313), .A3(n12312), .ZN(n12314) );
  MUX2_X1 U14690 ( .A(n12317), .B(n12316), .S(n12346), .Z(n12318) );
  NAND2_X1 U14691 ( .A1(n12954), .A2(n12774), .ZN(n12321) );
  MUX2_X1 U14692 ( .A(n12321), .B(n12320), .S(n12346), .Z(n12322) );
  MUX2_X1 U14693 ( .A(n12324), .B(n12323), .S(n12346), .Z(n12325) );
  NAND3_X1 U14694 ( .A1(n12326), .A2(n12729), .A3(n12325), .ZN(n12328) );
  MUX2_X1 U14695 ( .A(n12713), .B(n12714), .S(n12346), .Z(n12327) );
  XNOR2_X1 U14696 ( .A(n12330), .B(n12346), .ZN(n12331) );
  NOR2_X1 U14697 ( .A1(n12663), .A2(n12333), .ZN(n12335) );
  INV_X1 U14698 ( .A(n12336), .ZN(n12337) );
  NOR2_X1 U14699 ( .A1(n12663), .A2(n12337), .ZN(n12338) );
  OAI21_X1 U14700 ( .B1(n12665), .B2(n12339), .A(n12345), .ZN(n12340) );
  NAND2_X1 U14701 ( .A1(n12340), .A2(n12347), .ZN(n12344) );
  AOI21_X1 U14702 ( .B1(n12342), .B2(n12346), .A(n12341), .ZN(n12343) );
  NAND2_X1 U14703 ( .A1(n12344), .A2(n12343), .ZN(n12351) );
  INV_X1 U14704 ( .A(n12345), .ZN(n12348) );
  NAND3_X1 U14705 ( .A1(n12348), .A2(n12347), .A3(n12346), .ZN(n12349) );
  NAND3_X1 U14706 ( .A1(n12351), .A2(n12350), .A3(n12349), .ZN(n12355) );
  INV_X1 U14707 ( .A(n12352), .ZN(n12353) );
  NAND3_X1 U14708 ( .A1(n12355), .A2(n12354), .A3(n12353), .ZN(n12358) );
  AOI21_X1 U14709 ( .B1(n12358), .B2(n6755), .A(n12357), .ZN(n12363) );
  NAND2_X1 U14710 ( .A1(n12365), .A2(n12364), .ZN(n12366) );
  OAI211_X1 U14711 ( .C1(n12367), .C2(n12369), .A(n12366), .B(P3_B_REG_SCAN_IN), .ZN(n12368) );
  INV_X1 U14712 ( .A(n12371), .ZN(n12372) );
  NOR2_X1 U14713 ( .A1(n12373), .A2(n12910), .ZN(n12633) );
  AOI21_X1 U14714 ( .B1(n12786), .B2(P3_REG2_REG_29__SCAN_IN), .A(n12633), 
        .ZN(n12374) );
  OAI21_X1 U14715 ( .B1(n12375), .B2(n12870), .A(n12374), .ZN(n12376) );
  AOI21_X1 U14716 ( .B1(n7420), .B2(n12888), .A(n12376), .ZN(n12377) );
  OAI21_X1 U14717 ( .B1(n12378), .B2(n12891), .A(n12377), .ZN(P3_U3204) );
  XNOR2_X1 U14718 ( .A(n12380), .B(n12379), .ZN(n12388) );
  INV_X1 U14719 ( .A(n12388), .ZN(n12381) );
  NAND2_X1 U14720 ( .A1(n12381), .A2(n12477), .ZN(n12395) );
  INV_X1 U14721 ( .A(n12382), .ZN(n12383) );
  NAND4_X1 U14722 ( .A1(n12394), .A2(n12477), .A3(n12383), .A4(n12388), .ZN(
        n12393) );
  AOI22_X1 U14723 ( .A1(n7132), .A2(n12468), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12386) );
  NAND2_X1 U14724 ( .A1(n12640), .A2(n12482), .ZN(n12385) );
  OAI211_X1 U14725 ( .C1(n12665), .C2(n12479), .A(n12386), .B(n12385), .ZN(
        n12390) );
  NOR4_X1 U14726 ( .A1(n12388), .A2(n12387), .A3(n12499), .A4(n12503), .ZN(
        n12389) );
  AOI211_X1 U14727 ( .C1(n12497), .C2(n12391), .A(n12390), .B(n12389), .ZN(
        n12392) );
  OAI211_X1 U14728 ( .C1(n12395), .C2(n12394), .A(n12393), .B(n12392), .ZN(
        P3_U3160) );
  XNOR2_X1 U14729 ( .A(n12397), .B(n12396), .ZN(n12404) );
  INV_X1 U14730 ( .A(n13046), .ZN(n12402) );
  INV_X1 U14731 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n15151) );
  NOR2_X1 U14732 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15151), .ZN(n12533) );
  NOR2_X1 U14733 ( .A1(n12398), .A2(n12491), .ZN(n12399) );
  AOI211_X1 U14734 ( .C1(n12493), .C2(n8969), .A(n12533), .B(n12399), .ZN(
        n12400) );
  OAI21_X1 U14735 ( .B1(n12855), .B2(n12495), .A(n12400), .ZN(n12401) );
  AOI21_X1 U14736 ( .B1(n12402), .B2(n12497), .A(n12401), .ZN(n12403) );
  OAI21_X1 U14737 ( .B1(n12404), .B2(n12499), .A(n12403), .ZN(P3_U3155) );
  AOI21_X1 U14738 ( .B1(n12505), .B2(n12405), .A(n6502), .ZN(n12411) );
  AOI22_X1 U14739 ( .A1(n12493), .A2(n12708), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12407) );
  NAND2_X1 U14740 ( .A1(n12482), .A2(n12720), .ZN(n12406) );
  OAI211_X1 U14741 ( .C1(n12408), .C2(n12491), .A(n12407), .B(n12406), .ZN(
        n12409) );
  AOI21_X1 U14742 ( .B1(n12721), .B2(n12497), .A(n12409), .ZN(n12410) );
  OAI21_X1 U14743 ( .B1(n12411), .B2(n12499), .A(n12410), .ZN(P3_U3156) );
  XOR2_X1 U14744 ( .A(n12412), .B(n12413), .Z(n12414) );
  NAND2_X1 U14745 ( .A1(n12414), .A2(n12477), .ZN(n12418) );
  NAND2_X1 U14746 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12626)
         );
  OAI21_X1 U14747 ( .B1(n12774), .B2(n12491), .A(n12626), .ZN(n12416) );
  NOR2_X1 U14748 ( .A1(n12495), .A2(n12781), .ZN(n12415) );
  AOI211_X1 U14749 ( .C1(n12493), .C2(n12806), .A(n12416), .B(n12415), .ZN(
        n12417) );
  OAI211_X1 U14750 ( .C1(n12485), .C2(n13034), .A(n12418), .B(n12417), .ZN(
        P3_U3159) );
  AOI21_X1 U14751 ( .B1(n12420), .B2(n12419), .A(n6549), .ZN(n12425) );
  AOI22_X1 U14752 ( .A1(n12493), .A2(n12507), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12422) );
  NAND2_X1 U14753 ( .A1(n12482), .A2(n12749), .ZN(n12421) );
  OAI211_X1 U14754 ( .C1(n12745), .C2(n12491), .A(n12422), .B(n12421), .ZN(
        n12423) );
  AOI21_X1 U14755 ( .B1(n12748), .B2(n12497), .A(n12423), .ZN(n12424) );
  OAI21_X1 U14756 ( .B1(n12425), .B2(n12499), .A(n12424), .ZN(P3_U3163) );
  INV_X1 U14757 ( .A(n12978), .ZN(n12823) );
  OAI211_X1 U14758 ( .C1(n12428), .C2(n12427), .A(n12426), .B(n12477), .ZN(
        n12432) );
  NAND2_X1 U14759 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12582)
         );
  OAI21_X1 U14760 ( .B1(n12791), .B2(n12491), .A(n12582), .ZN(n12430) );
  NOR2_X1 U14761 ( .A1(n12495), .A2(n12824), .ZN(n12429) );
  AOI211_X1 U14762 ( .C1(n12493), .C2(n12845), .A(n12430), .B(n12429), .ZN(
        n12431) );
  OAI211_X1 U14763 ( .C1(n12823), .C2(n12485), .A(n12432), .B(n12431), .ZN(
        P3_U3166) );
  INV_X1 U14764 ( .A(n12974), .ZN(n12810) );
  OAI211_X1 U14765 ( .C1(n12435), .C2(n12434), .A(n12433), .B(n12477), .ZN(
        n12439) );
  NOR2_X1 U14766 ( .A1(n12495), .A2(n12811), .ZN(n12437) );
  NAND2_X1 U14767 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14331)
         );
  OAI21_X1 U14768 ( .B1(n12479), .B2(n12832), .A(n14331), .ZN(n12436) );
  AOI211_X1 U14769 ( .C1(n12468), .C2(n12806), .A(n12437), .B(n12436), .ZN(
        n12438) );
  OAI211_X1 U14770 ( .C1(n12810), .C2(n12485), .A(n12439), .B(n12438), .ZN(
        P3_U3168) );
  NOR3_X1 U14771 ( .A1(n6502), .A2(n7254), .A3(n12441), .ZN(n12444) );
  INV_X1 U14772 ( .A(n12442), .ZN(n12443) );
  OAI21_X1 U14773 ( .B1(n12444), .B2(n12443), .A(n12477), .ZN(n12448) );
  AOI22_X1 U14774 ( .A1(n12505), .A2(n12493), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12445) );
  OAI21_X1 U14775 ( .B1(n12690), .B2(n12491), .A(n12445), .ZN(n12446) );
  AOI21_X1 U14776 ( .B1(n12700), .B2(n12482), .A(n12446), .ZN(n12447) );
  OAI211_X1 U14777 ( .C1(n12485), .C2(n12702), .A(n12448), .B(n12447), .ZN(
        P3_U3169) );
  XNOR2_X1 U14778 ( .A(n12449), .B(n12450), .ZN(n12455) );
  AOI22_X1 U14779 ( .A1(n12493), .A2(n12508), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12452) );
  NAND2_X1 U14780 ( .A1(n12482), .A2(n12760), .ZN(n12451) );
  OAI211_X1 U14781 ( .C1(n12759), .C2(n12491), .A(n12452), .B(n12451), .ZN(
        n12453) );
  AOI21_X1 U14782 ( .B1(n12954), .B2(n12497), .A(n12453), .ZN(n12454) );
  OAI21_X1 U14783 ( .B1(n12455), .B2(n12499), .A(n12454), .ZN(P3_U3173) );
  INV_X1 U14784 ( .A(n12456), .ZN(n12457) );
  AOI21_X1 U14785 ( .B1(n12708), .B2(n12458), .A(n12457), .ZN(n12463) );
  NOR2_X1 U14786 ( .A1(n12479), .A2(n12759), .ZN(n12460) );
  INV_X1 U14787 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n15057) );
  OAI22_X1 U14788 ( .A1(n12728), .A2(n12491), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15057), .ZN(n12459) );
  AOI211_X1 U14789 ( .C1(n12731), .C2(n12482), .A(n12460), .B(n12459), .ZN(
        n12462) );
  NAND2_X1 U14790 ( .A1(n12730), .A2(n12497), .ZN(n12461) );
  OAI211_X1 U14791 ( .C1(n12463), .C2(n12499), .A(n12462), .B(n12461), .ZN(
        P3_U3175) );
  XNOR2_X1 U14792 ( .A(n12464), .B(n12775), .ZN(n12465) );
  XNOR2_X1 U14793 ( .A(n12466), .B(n12465), .ZN(n12472) );
  NAND2_X1 U14794 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n14358)
         );
  OAI21_X1 U14795 ( .B1(n12479), .B2(n12791), .A(n14358), .ZN(n12467) );
  AOI21_X1 U14796 ( .B1(n12468), .B2(n12508), .A(n12467), .ZN(n12469) );
  OAI21_X1 U14797 ( .B1(n12793), .B2(n12495), .A(n12469), .ZN(n12470) );
  AOI21_X1 U14798 ( .B1(n12967), .B2(n12497), .A(n12470), .ZN(n12471) );
  OAI21_X1 U14799 ( .B1(n12472), .B2(n12499), .A(n12471), .ZN(P3_U3178) );
  NAND2_X1 U14800 ( .A1(n12474), .A2(n12473), .ZN(n12476) );
  XNOR2_X1 U14801 ( .A(n12476), .B(n12475), .ZN(n12478) );
  NAND2_X1 U14802 ( .A1(n12478), .A2(n12477), .ZN(n12484) );
  INV_X1 U14803 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n15093) );
  OAI22_X1 U14804 ( .A1(n12690), .A2(n12479), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15093), .ZN(n12481) );
  NOR2_X1 U14805 ( .A1(n12665), .A2(n12491), .ZN(n12480) );
  AOI211_X1 U14806 ( .C1(n12671), .C2(n12482), .A(n12481), .B(n12480), .ZN(
        n12483) );
  OAI211_X1 U14807 ( .C1(n13015), .C2(n12485), .A(n12484), .B(n12483), .ZN(
        P3_U3180) );
  INV_X1 U14808 ( .A(n12486), .ZN(n12488) );
  NAND2_X1 U14809 ( .A1(n12488), .A2(n12487), .ZN(n12489) );
  XNOR2_X1 U14810 ( .A(n12490), .B(n12489), .ZN(n12500) );
  NOR2_X1 U14811 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8373), .ZN(n12556) );
  NOR2_X1 U14812 ( .A1(n12832), .A2(n12491), .ZN(n12492) );
  AOI211_X1 U14813 ( .C1(n12493), .C2(n12509), .A(n12556), .B(n12492), .ZN(
        n12494) );
  OAI21_X1 U14814 ( .B1(n12836), .B2(n12495), .A(n12494), .ZN(n12496) );
  AOI21_X1 U14815 ( .B1(n12497), .B2(n12835), .A(n12496), .ZN(n12498) );
  OAI21_X1 U14816 ( .B1(n12500), .B2(n12499), .A(n12498), .ZN(P3_U3181) );
  MUX2_X1 U14817 ( .A(n12501), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12522), .Z(
        P3_U3522) );
  MUX2_X1 U14818 ( .A(n12502), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12522), .Z(
        P3_U3521) );
  MUX2_X1 U14819 ( .A(n7132), .B(P3_DATAO_REG_29__SCAN_IN), .S(n12522), .Z(
        P3_U3520) );
  MUX2_X1 U14820 ( .A(n12503), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12522), .Z(
        P3_U3518) );
  MUX2_X1 U14821 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12679), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14822 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12504), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14823 ( .A(n12709), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12522), .Z(
        P3_U3515) );
  MUX2_X1 U14824 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12505), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14825 ( .A(n12708), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12522), .Z(
        P3_U3513) );
  MUX2_X1 U14826 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12506), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14827 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12507), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14828 ( .A(n12508), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12522), .Z(
        P3_U3510) );
  MUX2_X1 U14829 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12806), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14830 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12818), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14831 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12805), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14832 ( .A(n12845), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12522), .Z(
        P3_U3506) );
  MUX2_X1 U14833 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12509), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14834 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n8969), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14835 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12510), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14836 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12511), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14837 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12512), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14838 ( .A(n12513), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12522), .Z(
        P3_U3500) );
  MUX2_X1 U14839 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12514), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14840 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12515), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14841 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12516), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14842 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12517), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14843 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12518), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14844 ( .A(n12519), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12522), .Z(
        P3_U3494) );
  MUX2_X1 U14845 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12520), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14846 ( .A(n12521), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12522), .Z(
        P3_U3492) );
  MUX2_X1 U14847 ( .A(n12523), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12522), .Z(
        P3_U3491) );
  NOR2_X1 U14848 ( .A1(n12538), .A2(n12524), .ZN(n12526) );
  XNOR2_X1 U14849 ( .A(n12558), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n12540) );
  AOI21_X1 U14850 ( .B1(n6609), .B2(n12540), .A(n12551), .ZN(n12550) );
  NOR2_X1 U14851 ( .A1(n12558), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12527) );
  AOI21_X1 U14852 ( .B1(P3_REG1_REG_14__SCAN_IN), .B2(n12558), .A(n12527), 
        .ZN(n12543) );
  NAND2_X1 U14853 ( .A1(n12529), .A2(n12528), .ZN(n12531) );
  NAND2_X1 U14854 ( .A1(n12531), .A2(n12530), .ZN(n12532) );
  NAND2_X1 U14855 ( .A1(n12543), .A2(n12532), .ZN(n12554) );
  OAI21_X1 U14856 ( .B1(n12543), .B2(n12532), .A(n12554), .ZN(n12536) );
  AOI21_X1 U14857 ( .B1(n14943), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12533), 
        .ZN(n12534) );
  OAI21_X1 U14858 ( .B1(n14970), .B2(n12558), .A(n12534), .ZN(n12535) );
  AOI21_X1 U14859 ( .B1(n12536), .B2(n14954), .A(n12535), .ZN(n12549) );
  INV_X1 U14860 ( .A(n12537), .ZN(n12539) );
  NAND2_X1 U14861 ( .A1(n12539), .A2(n12538), .ZN(n12544) );
  AND2_X1 U14862 ( .A1(n12545), .A2(n12544), .ZN(n12547) );
  INV_X1 U14863 ( .A(n12540), .ZN(n12542) );
  MUX2_X1 U14864 ( .A(n12543), .B(n12542), .S(n12541), .Z(n12546) );
  NAND3_X1 U14865 ( .A1(n12545), .A2(n12544), .A3(n12546), .ZN(n12562) );
  OAI211_X1 U14866 ( .C1(n12547), .C2(n12546), .A(n14964), .B(n12562), .ZN(
        n12548) );
  OAI211_X1 U14867 ( .C1(n12550), .C2(n14959), .A(n12549), .B(n12548), .ZN(
        P3_U3196) );
  AOI21_X1 U14868 ( .B1(n12553), .B2(n12552), .A(n12572), .ZN(n12570) );
  NAND2_X1 U14869 ( .A1(n12558), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12559) );
  NAND2_X1 U14870 ( .A1(n12559), .A2(n12554), .ZN(n12576) );
  XNOR2_X1 U14871 ( .A(n12588), .B(n12576), .ZN(n12555) );
  NAND2_X1 U14872 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12555), .ZN(n12578) );
  OAI21_X1 U14873 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12555), .A(n12578), 
        .ZN(n12568) );
  AOI21_X1 U14874 ( .B1(n14943), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n12556), 
        .ZN(n12557) );
  OAI21_X1 U14875 ( .B1(n14970), .B2(n12577), .A(n12557), .ZN(n12567) );
  MUX2_X1 U14876 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12601), .Z(n12564) );
  NAND2_X1 U14877 ( .A1(n12558), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12560) );
  MUX2_X1 U14878 ( .A(n12560), .B(n12559), .S(n12601), .Z(n12561) );
  NAND2_X1 U14879 ( .A1(n12562), .A2(n12561), .ZN(n12586) );
  XNOR2_X1 U14880 ( .A(n12586), .B(n12577), .ZN(n12563) );
  NOR2_X1 U14881 ( .A1(n12563), .A2(n12564), .ZN(n12587) );
  AOI21_X1 U14882 ( .B1(n12564), .B2(n12563), .A(n12587), .ZN(n12565) );
  NOR2_X1 U14883 ( .A1(n12565), .A2(n14939), .ZN(n12566) );
  AOI211_X1 U14884 ( .C1(n14954), .C2(n12568), .A(n12567), .B(n12566), .ZN(
        n12569) );
  OAI21_X1 U14885 ( .B1(n12570), .B2(n14959), .A(n12569), .ZN(P3_U3197) );
  NOR2_X1 U14886 ( .A1(n12588), .A2(n12571), .ZN(n12573) );
  AOI22_X1 U14887 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12617), .B1(n12598), 
        .B2(n12825), .ZN(n12574) );
  AOI21_X1 U14888 ( .B1(n12575), .B2(n12574), .A(n12597), .ZN(n12596) );
  AOI22_X1 U14889 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12598), .B1(n12617), 
        .B2(n12616), .ZN(n12581) );
  NAND2_X1 U14890 ( .A1(n12577), .A2(n12576), .ZN(n12579) );
  NAND2_X1 U14891 ( .A1(n12579), .A2(n12578), .ZN(n12580) );
  NAND2_X1 U14892 ( .A1(n12581), .A2(n12580), .ZN(n12615) );
  OAI21_X1 U14893 ( .B1(n12581), .B2(n12580), .A(n12615), .ZN(n12585) );
  NOR2_X1 U14894 ( .A1(n14970), .A2(n12598), .ZN(n12584) );
  INV_X1 U14895 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14233) );
  OAI21_X1 U14896 ( .B1(n14975), .B2(n14233), .A(n12582), .ZN(n12583) );
  AOI211_X1 U14897 ( .C1(n12585), .C2(n14954), .A(n12584), .B(n12583), .ZN(
        n12595) );
  INV_X1 U14898 ( .A(n12586), .ZN(n12589) );
  AOI21_X1 U14899 ( .B1(n12589), .B2(n12588), .A(n12587), .ZN(n12604) );
  MUX2_X1 U14900 ( .A(n12825), .B(n12616), .S(n12601), .Z(n12590) );
  NOR2_X1 U14901 ( .A1(n12590), .A2(n12617), .ZN(n12603) );
  INV_X1 U14902 ( .A(n12603), .ZN(n12591) );
  NAND2_X1 U14903 ( .A1(n12590), .A2(n12617), .ZN(n12602) );
  NAND2_X1 U14904 ( .A1(n12591), .A2(n12602), .ZN(n12592) );
  XNOR2_X1 U14905 ( .A(n12604), .B(n12592), .ZN(n12593) );
  NAND2_X1 U14906 ( .A1(n12593), .A2(n14964), .ZN(n12594) );
  OAI211_X1 U14907 ( .C1(n12596), .C2(n14959), .A(n12595), .B(n12594), .ZN(
        P3_U3198) );
  INV_X1 U14908 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12600) );
  AOI22_X1 U14909 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n14342), .B1(n12614), 
        .B2(n12600), .ZN(n14354) );
  XNOR2_X1 U14910 ( .A(n12609), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12608) );
  MUX2_X1 U14911 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12601), .Z(n12605) );
  OAI21_X1 U14912 ( .B1(n12604), .B2(n12603), .A(n12602), .ZN(n14335) );
  XNOR2_X1 U14913 ( .A(n12605), .B(n12618), .ZN(n14336) );
  NOR2_X1 U14914 ( .A1(n14335), .A2(n14336), .ZN(n14334) );
  AOI21_X1 U14915 ( .B1(n12605), .B2(n12618), .A(n14334), .ZN(n12607) );
  INV_X1 U14916 ( .A(n12607), .ZN(n12606) );
  XNOR2_X1 U14917 ( .A(n12606), .B(n12614), .ZN(n14348) );
  MUX2_X1 U14918 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12601), .Z(n14349) );
  NOR2_X1 U14919 ( .A1(n14348), .A2(n14349), .ZN(n14347) );
  AOI21_X1 U14920 ( .B1(n12607), .B2(n14342), .A(n14347), .ZN(n12613) );
  INV_X1 U14921 ( .A(n12608), .ZN(n12611) );
  XNOR2_X1 U14922 ( .A(n12609), .B(n12964), .ZN(n12621) );
  MUX2_X1 U14923 ( .A(n12611), .B(n12621), .S(n12601), .Z(n12612) );
  XNOR2_X1 U14924 ( .A(n12613), .B(n12612), .ZN(n12629) );
  AOI22_X1 U14925 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n12614), .B1(n14342), 
        .B2(n12972), .ZN(n14346) );
  NAND2_X1 U14926 ( .A1(n12618), .A2(n12619), .ZN(n12620) );
  XNOR2_X1 U14927 ( .A(n12619), .B(n14330), .ZN(n14329) );
  NAND2_X1 U14928 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14329), .ZN(n14328) );
  NAND2_X1 U14929 ( .A1(n12620), .A2(n14328), .ZN(n14345) );
  XNOR2_X1 U14930 ( .A(n12622), .B(n12621), .ZN(n12624) );
  NOR2_X1 U14931 ( .A1(n12624), .A2(n12623), .ZN(n12628) );
  NAND2_X1 U14932 ( .A1(n14943), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12625) );
  OAI211_X1 U14933 ( .C1(n14970), .C2(n12193), .A(n12626), .B(n12625), .ZN(
        n12627) );
  NAND2_X1 U14934 ( .A1(n12997), .A2(n12801), .ZN(n12634) );
  NOR2_X1 U14935 ( .A1(n12632), .A2(n12631), .ZN(n12998) );
  AOI21_X1 U14936 ( .B1(n12998), .B2(n12813), .A(n12633), .ZN(n12637) );
  OAI211_X1 U14937 ( .C1(n12635), .C2(n12813), .A(n12634), .B(n12637), .ZN(
        P3_U3202) );
  NAND2_X1 U14938 ( .A1(n12891), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n12636) );
  OAI211_X1 U14939 ( .C1(n12638), .C2(n12870), .A(n12637), .B(n12636), .ZN(
        P3_U3203) );
  INV_X1 U14940 ( .A(n12639), .ZN(n12645) );
  AOI22_X1 U14941 ( .A1(n12640), .A2(n12868), .B1(n12891), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12641) );
  OAI21_X1 U14942 ( .B1(n13007), .B2(n12870), .A(n12641), .ZN(n12642) );
  AOI21_X1 U14943 ( .B1(n12643), .B2(n12888), .A(n12642), .ZN(n12644) );
  OAI21_X1 U14944 ( .B1(n12645), .B2(n12891), .A(n12644), .ZN(P3_U3205) );
  AOI21_X1 U14945 ( .B1(n12649), .B2(n12647), .A(n12646), .ZN(n12655) );
  OAI21_X1 U14946 ( .B1(n12650), .B2(n12649), .A(n12648), .ZN(n12926) );
  OAI22_X1 U14947 ( .A1(n12652), .A2(n12908), .B1(n12651), .B2(n12906), .ZN(
        n12653) );
  AOI21_X1 U14948 ( .B1(n12926), .B2(n12667), .A(n12653), .ZN(n12654) );
  INV_X1 U14949 ( .A(n12925), .ZN(n12661) );
  INV_X1 U14950 ( .A(n12656), .ZN(n12670) );
  AOI22_X1 U14951 ( .A1(n12657), .A2(n12868), .B1(n12786), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12658) );
  OAI21_X1 U14952 ( .B1(n13011), .B2(n12870), .A(n12658), .ZN(n12659) );
  AOI21_X1 U14953 ( .B1(n12926), .B2(n12670), .A(n12659), .ZN(n12660) );
  OAI21_X1 U14954 ( .B1(n12661), .B2(n12786), .A(n12660), .ZN(P3_U3206) );
  XNOR2_X1 U14955 ( .A(n12662), .B(n12663), .ZN(n12669) );
  XNOR2_X1 U14956 ( .A(n12664), .B(n12663), .ZN(n12930) );
  OAI22_X1 U14957 ( .A1(n12665), .A2(n12908), .B1(n12690), .B2(n12906), .ZN(
        n12666) );
  AOI21_X1 U14958 ( .B1(n12930), .B2(n12667), .A(n12666), .ZN(n12668) );
  OAI21_X1 U14959 ( .B1(n12669), .B2(n12903), .A(n12668), .ZN(n12929) );
  NAND2_X1 U14960 ( .A1(n12930), .A2(n12670), .ZN(n12673) );
  AOI22_X1 U14961 ( .A1(n12671), .A2(n12868), .B1(P3_REG2_REG_26__SCAN_IN), 
        .B2(n12891), .ZN(n12672) );
  OAI211_X1 U14962 ( .C1(n13015), .C2(n12870), .A(n12673), .B(n12672), .ZN(
        n12674) );
  AOI21_X1 U14963 ( .B1(n12929), .B2(n12813), .A(n12674), .ZN(n12675) );
  INV_X1 U14964 ( .A(n12675), .ZN(P3_U3207) );
  OAI211_X1 U14965 ( .C1(n12678), .C2(n12677), .A(n12676), .B(n12878), .ZN(
        n12681) );
  AOI22_X1 U14966 ( .A1(n12679), .A2(n12846), .B1(n12847), .B2(n12709), .ZN(
        n12680) );
  AND2_X1 U14967 ( .A1(n12681), .A2(n12680), .ZN(n12936) );
  XNOR2_X1 U14968 ( .A(n12682), .B(n6704), .ZN(n12934) );
  NAND2_X1 U14969 ( .A1(n12933), .A2(n12801), .ZN(n12685) );
  AOI22_X1 U14970 ( .A1(n12683), .A2(n12868), .B1(n12891), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12684) );
  NAND2_X1 U14971 ( .A1(n12685), .A2(n12684), .ZN(n12686) );
  AOI21_X1 U14972 ( .B1(n12934), .B2(n12888), .A(n12686), .ZN(n12687) );
  OAI21_X1 U14973 ( .B1(n12936), .B2(n12786), .A(n12687), .ZN(P3_U3208) );
  INV_X1 U14974 ( .A(n12688), .ZN(n12689) );
  AOI21_X1 U14975 ( .B1(n12689), .B2(n12698), .A(n12903), .ZN(n12693) );
  OAI22_X1 U14976 ( .A1(n12690), .A2(n12908), .B1(n12728), .B2(n12906), .ZN(
        n12691) );
  AOI21_X1 U14977 ( .B1(n12693), .B2(n12692), .A(n12691), .ZN(n12940) );
  AND2_X1 U14978 ( .A1(n12695), .A2(n12694), .ZN(n12719) );
  AND2_X1 U14979 ( .A1(n12719), .A2(n12696), .ZN(n12699) );
  OAI21_X1 U14980 ( .B1(n12699), .B2(n12698), .A(n12697), .ZN(n12938) );
  AOI22_X1 U14981 ( .A1(n12700), .A2(n12868), .B1(n12891), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12701) );
  OAI21_X1 U14982 ( .B1(n12702), .B2(n12870), .A(n12701), .ZN(n12703) );
  AOI21_X1 U14983 ( .B1(n12938), .B2(n12888), .A(n12703), .ZN(n12704) );
  OAI21_X1 U14984 ( .B1(n12940), .B2(n12891), .A(n12704), .ZN(P3_U3209) );
  OAI211_X1 U14985 ( .C1(n12707), .C2(n12706), .A(n12705), .B(n12878), .ZN(
        n12711) );
  AOI22_X1 U14986 ( .A1(n12709), .A2(n12846), .B1(n12847), .B2(n12708), .ZN(
        n12710) );
  NAND2_X1 U14987 ( .A1(n12711), .A2(n12710), .ZN(n12945) );
  NAND2_X1 U14988 ( .A1(n12712), .A2(n12713), .ZN(n12715) );
  NAND2_X1 U14989 ( .A1(n12715), .A2(n12714), .ZN(n12717) );
  OR2_X1 U14990 ( .A1(n12717), .A2(n12716), .ZN(n12718) );
  NAND2_X1 U14991 ( .A1(n12719), .A2(n12718), .ZN(n12943) );
  AOI22_X1 U14992 ( .A1(n12891), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n12720), 
        .B2(n12868), .ZN(n12723) );
  NAND2_X1 U14993 ( .A1(n12721), .A2(n12801), .ZN(n12722) );
  OAI211_X1 U14994 ( .C1(n12943), .C2(n12918), .A(n12723), .B(n12722), .ZN(
        n12724) );
  AOI21_X1 U14995 ( .B1(n12945), .B2(n12813), .A(n12724), .ZN(n12725) );
  INV_X1 U14996 ( .A(n12725), .ZN(P3_U3210) );
  XNOR2_X1 U14997 ( .A(n12726), .B(n12729), .ZN(n12727) );
  OAI222_X1 U14998 ( .A1(n12906), .A2(n12759), .B1(n12908), .B2(n12728), .C1(
        n12903), .C2(n12727), .ZN(n12946) );
  INV_X1 U14999 ( .A(n12946), .ZN(n12735) );
  XOR2_X1 U15000 ( .A(n12729), .B(n12712), .Z(n12947) );
  INV_X1 U15001 ( .A(n12730), .ZN(n13022) );
  AOI22_X1 U15002 ( .A1(n12891), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n12868), 
        .B2(n12731), .ZN(n12732) );
  OAI21_X1 U15003 ( .B1(n13022), .B2(n12870), .A(n12732), .ZN(n12733) );
  AOI21_X1 U15004 ( .B1(n12947), .B2(n12888), .A(n12733), .ZN(n12734) );
  OAI21_X1 U15005 ( .B1(n12735), .B2(n12891), .A(n12734), .ZN(P3_U3211) );
  OR2_X1 U15006 ( .A1(n12736), .A2(n12737), .ZN(n12739) );
  AND2_X1 U15007 ( .A1(n12739), .A2(n12738), .ZN(n12742) );
  AOI21_X1 U15008 ( .B1(n12743), .B2(n12742), .A(n6558), .ZN(n12744) );
  OAI222_X1 U15009 ( .A1(n12908), .A2(n12745), .B1(n12906), .B2(n12774), .C1(
        n12903), .C2(n12744), .ZN(n12950) );
  INV_X1 U15010 ( .A(n12950), .ZN(n12753) );
  XNOR2_X1 U15011 ( .A(n12747), .B(n12746), .ZN(n12951) );
  INV_X1 U15012 ( .A(n12748), .ZN(n13026) );
  AOI22_X1 U15013 ( .A1(n12891), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n12749), 
        .B2(n12868), .ZN(n12750) );
  OAI21_X1 U15014 ( .B1(n13026), .B2(n12870), .A(n12750), .ZN(n12751) );
  AOI21_X1 U15015 ( .B1(n12951), .B2(n12888), .A(n12751), .ZN(n12752) );
  OAI21_X1 U15016 ( .B1(n12753), .B2(n12786), .A(n12752), .ZN(P3_U3212) );
  OR2_X1 U15017 ( .A1(n12736), .A2(n12754), .ZN(n12756) );
  AND2_X1 U15018 ( .A1(n12756), .A2(n12755), .ZN(n12757) );
  XNOR2_X1 U15019 ( .A(n12757), .B(n12763), .ZN(n12758) );
  OAI222_X1 U15020 ( .A1(n12908), .A2(n12759), .B1(n12906), .B2(n12792), .C1(
        n12903), .C2(n12758), .ZN(n12956) );
  INV_X1 U15021 ( .A(n12956), .ZN(n12769) );
  INV_X1 U15022 ( .A(n12760), .ZN(n12761) );
  OAI22_X1 U15023 ( .A1(n12813), .A2(n12762), .B1(n12761), .B2(n12910), .ZN(
        n12767) );
  INV_X1 U15024 ( .A(n12957), .ZN(n12765) );
  AND2_X1 U15025 ( .A1(n12764), .A2(n12763), .ZN(n12955) );
  NOR3_X1 U15026 ( .A1(n12765), .A2(n12955), .A3(n12918), .ZN(n12766) );
  AOI211_X1 U15027 ( .C1(n12801), .C2(n12954), .A(n12767), .B(n12766), .ZN(
        n12768) );
  OAI21_X1 U15028 ( .B1(n12769), .B2(n12786), .A(n12768), .ZN(P3_U3213) );
  AND2_X1 U15029 ( .A1(n12787), .A2(n12770), .ZN(n12773) );
  NAND2_X1 U15030 ( .A1(n12787), .A2(n12771), .ZN(n12772) );
  OAI211_X1 U15031 ( .C1(n12773), .C2(n12779), .A(n12772), .B(n12878), .ZN(
        n12778) );
  OAI22_X1 U15032 ( .A1(n12775), .A2(n12906), .B1(n12774), .B2(n12908), .ZN(
        n12776) );
  INV_X1 U15033 ( .A(n12776), .ZN(n12777) );
  XNOR2_X1 U15034 ( .A(n12780), .B(n12779), .ZN(n12961) );
  NOR2_X1 U15035 ( .A1(n13034), .A2(n12870), .ZN(n12784) );
  OAI22_X1 U15036 ( .A1(n12813), .A2(n12782), .B1(n12781), .B2(n12910), .ZN(
        n12783) );
  AOI211_X1 U15037 ( .C1(n12961), .C2(n12888), .A(n12784), .B(n12783), .ZN(
        n12785) );
  OAI21_X1 U15038 ( .B1(n12963), .B2(n12786), .A(n12785), .ZN(P3_U3214) );
  INV_X1 U15039 ( .A(n12787), .ZN(n12788) );
  AOI21_X1 U15040 ( .B1(n12789), .B2(n12736), .A(n12788), .ZN(n12790) );
  OAI222_X1 U15041 ( .A1(n12908), .A2(n12792), .B1(n12906), .B2(n12791), .C1(
        n12903), .C2(n12790), .ZN(n12969) );
  INV_X1 U15042 ( .A(n12969), .ZN(n12803) );
  OAI22_X1 U15043 ( .A1(n12813), .A2(n12600), .B1(n12793), .B2(n12910), .ZN(
        n12800) );
  INV_X1 U15044 ( .A(n12970), .ZN(n12798) );
  NAND2_X1 U15045 ( .A1(n12795), .A2(n12794), .ZN(n12797) );
  NOR3_X1 U15046 ( .A1(n12798), .A2(n12968), .A3(n12918), .ZN(n12799) );
  AOI211_X1 U15047 ( .C1(n12801), .C2(n12967), .A(n12800), .B(n12799), .ZN(
        n12802) );
  OAI21_X1 U15048 ( .B1(n12803), .B2(n12891), .A(n12802), .ZN(P3_U3215) );
  XNOR2_X1 U15049 ( .A(n12804), .B(n12808), .ZN(n12807) );
  AOI222_X1 U15050 ( .A1(n12878), .A2(n12807), .B1(n12806), .B2(n12846), .C1(
        n12805), .C2(n12847), .ZN(n12977) );
  XNOR2_X1 U15051 ( .A(n12809), .B(n12808), .ZN(n12975) );
  NOR2_X1 U15052 ( .A1(n12810), .A2(n12870), .ZN(n12815) );
  OAI22_X1 U15053 ( .A1(n12813), .A2(n12812), .B1(n12811), .B2(n12910), .ZN(
        n12814) );
  AOI211_X1 U15054 ( .C1(n12975), .C2(n12888), .A(n12815), .B(n12814), .ZN(
        n12816) );
  OAI21_X1 U15055 ( .B1(n12977), .B2(n12891), .A(n12816), .ZN(P3_U3216) );
  XNOR2_X1 U15056 ( .A(n12817), .B(n12821), .ZN(n12819) );
  AOI222_X1 U15057 ( .A1(n12878), .A2(n12819), .B1(n12818), .B2(n12846), .C1(
        n12845), .C2(n12847), .ZN(n12982) );
  OAI21_X1 U15058 ( .B1(n12822), .B2(n12821), .A(n12820), .ZN(n12980) );
  NOR2_X1 U15059 ( .A1(n12823), .A2(n12870), .ZN(n12827) );
  OAI22_X1 U15060 ( .A1(n12813), .A2(n12825), .B1(n12824), .B2(n12910), .ZN(
        n12826) );
  AOI211_X1 U15061 ( .C1(n12980), .C2(n12888), .A(n12827), .B(n12826), .ZN(
        n12828) );
  OAI21_X1 U15062 ( .B1(n12982), .B2(n12891), .A(n12828), .ZN(P3_U3217) );
  XNOR2_X1 U15063 ( .A(n12829), .B(n12830), .ZN(n12831) );
  OAI222_X1 U15064 ( .A1(n12908), .A2(n12832), .B1(n12906), .B2(n12862), .C1(
        n12831), .C2(n12903), .ZN(n12983) );
  INV_X1 U15065 ( .A(n12983), .ZN(n12841) );
  XNOR2_X1 U15066 ( .A(n12834), .B(n12833), .ZN(n12984) );
  INV_X1 U15067 ( .A(n12835), .ZN(n13044) );
  INV_X1 U15068 ( .A(n12836), .ZN(n12837) );
  AOI22_X1 U15069 ( .A1(n12891), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n12868), 
        .B2(n12837), .ZN(n12838) );
  OAI21_X1 U15070 ( .B1(n13044), .B2(n12870), .A(n12838), .ZN(n12839) );
  AOI21_X1 U15071 ( .B1(n12984), .B2(n12888), .A(n12839), .ZN(n12840) );
  OAI21_X1 U15072 ( .B1(n12841), .B2(n12891), .A(n12840), .ZN(P3_U3218) );
  NAND2_X1 U15073 ( .A1(n12842), .A2(n12852), .ZN(n12843) );
  NAND3_X1 U15074 ( .A1(n12844), .A2(n12878), .A3(n12843), .ZN(n12849) );
  AOI22_X1 U15075 ( .A1(n8969), .A2(n12847), .B1(n12846), .B2(n12845), .ZN(
        n12848) );
  AND2_X1 U15076 ( .A1(n12849), .A2(n12848), .ZN(n12989) );
  NAND2_X1 U15077 ( .A1(n12851), .A2(n12850), .ZN(n12854) );
  INV_X1 U15078 ( .A(n12852), .ZN(n12853) );
  XNOR2_X1 U15079 ( .A(n12854), .B(n12853), .ZN(n12987) );
  NOR2_X1 U15080 ( .A1(n13046), .A2(n12870), .ZN(n12858) );
  OAI22_X1 U15081 ( .A1(n12813), .A2(n12856), .B1(n12855), .B2(n12910), .ZN(
        n12857) );
  AOI211_X1 U15082 ( .C1(n12987), .C2(n12888), .A(n12858), .B(n12857), .ZN(
        n12859) );
  OAI21_X1 U15083 ( .B1(n12989), .B2(n12891), .A(n12859), .ZN(P3_U3219) );
  XNOR2_X1 U15084 ( .A(n12860), .B(n12866), .ZN(n12861) );
  OAI222_X1 U15085 ( .A1(n12908), .A2(n12862), .B1(n12906), .B2(n12907), .C1(
        n12861), .C2(n12903), .ZN(n12992) );
  INV_X1 U15086 ( .A(n12992), .ZN(n12873) );
  NAND2_X1 U15087 ( .A1(n12864), .A2(n12863), .ZN(n12865) );
  XOR2_X1 U15088 ( .A(n12866), .B(n12865), .Z(n12993) );
  AOI22_X1 U15089 ( .A1(n12891), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n12868), 
        .B2(n12867), .ZN(n12869) );
  OAI21_X1 U15090 ( .B1(n13052), .B2(n12870), .A(n12869), .ZN(n12871) );
  AOI21_X1 U15091 ( .B1(n12993), .B2(n12888), .A(n12871), .ZN(n12872) );
  OAI21_X1 U15092 ( .B1(n12873), .B2(n12891), .A(n12872), .ZN(P3_U3220) );
  XNOR2_X1 U15093 ( .A(n12874), .B(n12886), .ZN(n12879) );
  OAI22_X1 U15094 ( .A1(n12876), .A2(n12906), .B1(n12875), .B2(n12908), .ZN(
        n12877) );
  AOI21_X1 U15095 ( .B1(n12879), .B2(n12878), .A(n12877), .ZN(n14364) );
  AND2_X1 U15096 ( .A1(n12880), .A2(n12979), .ZN(n14361) );
  OAI22_X1 U15097 ( .A1(n12813), .A2(n12882), .B1(n12881), .B2(n12910), .ZN(
        n12883) );
  AOI21_X1 U15098 ( .B1(n12914), .B2(n14361), .A(n12883), .ZN(n12890) );
  NAND2_X1 U15099 ( .A1(n12893), .A2(n12884), .ZN(n12897) );
  NAND2_X1 U15100 ( .A1(n12897), .A2(n12885), .ZN(n12887) );
  XNOR2_X1 U15101 ( .A(n12887), .B(n12886), .ZN(n14362) );
  NAND2_X1 U15102 ( .A1(n14362), .A2(n12888), .ZN(n12889) );
  OAI211_X1 U15103 ( .C1(n14364), .C2(n12891), .A(n12890), .B(n12889), .ZN(
        P3_U3221) );
  NAND2_X1 U15104 ( .A1(n12893), .A2(n12892), .ZN(n12895) );
  NAND2_X1 U15105 ( .A1(n12895), .A2(n12894), .ZN(n12900) );
  AND2_X1 U15106 ( .A1(n12897), .A2(n12896), .ZN(n12898) );
  OAI21_X1 U15107 ( .B1(n12900), .B2(n12899), .A(n12898), .ZN(n14367) );
  INV_X1 U15108 ( .A(n14367), .ZN(n12917) );
  XNOR2_X1 U15109 ( .A(n12902), .B(n12901), .ZN(n12904) );
  OAI222_X1 U15110 ( .A1(n12908), .A2(n12907), .B1(n12906), .B2(n12905), .C1(
        n12904), .C2(n12903), .ZN(n14365) );
  NAND2_X1 U15111 ( .A1(n14365), .A2(n12813), .ZN(n12916) );
  NOR2_X1 U15112 ( .A1(n12909), .A2(n12941), .ZN(n14366) );
  OAI22_X1 U15113 ( .A1(n12813), .A2(n12912), .B1(n12911), .B2(n12910), .ZN(
        n12913) );
  AOI21_X1 U15114 ( .B1(n12914), .B2(n14366), .A(n12913), .ZN(n12915) );
  OAI211_X1 U15115 ( .C1(n12918), .C2(n12917), .A(n12916), .B(n12915), .ZN(
        P3_U3222) );
  INV_X1 U15116 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12920) );
  NAND2_X1 U15117 ( .A1(n12997), .A2(n8875), .ZN(n12919) );
  NAND2_X1 U15118 ( .A1(n12998), .A2(n15016), .ZN(n12921) );
  OAI211_X1 U15119 ( .C1(n15016), .C2(n12920), .A(n12919), .B(n12921), .ZN(
        P3_U3490) );
  INV_X1 U15120 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n12923) );
  NAND2_X1 U15121 ( .A1(n13001), .A2(n8875), .ZN(n12922) );
  OAI211_X1 U15122 ( .C1(n15016), .C2(n12923), .A(n12922), .B(n12921), .ZN(
        P3_U3489) );
  INV_X1 U15123 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12927) );
  INV_X1 U15124 ( .A(n12924), .ZN(n14997) );
  AOI21_X1 U15125 ( .B1(n14997), .B2(n12926), .A(n12925), .ZN(n13008) );
  MUX2_X1 U15126 ( .A(n12927), .B(n13008), .S(n15016), .Z(n12928) );
  OAI21_X1 U15127 ( .B1(n13011), .B2(n12996), .A(n12928), .ZN(P3_U3486) );
  INV_X1 U15128 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12931) );
  AOI21_X1 U15129 ( .B1(n14997), .B2(n12930), .A(n12929), .ZN(n13012) );
  MUX2_X1 U15130 ( .A(n12931), .B(n13012), .S(n15016), .Z(n12932) );
  OAI21_X1 U15131 ( .B1(n13015), .B2(n12996), .A(n12932), .ZN(P3_U3485) );
  AOI22_X1 U15132 ( .A1(n12934), .A2(n8900), .B1(n12979), .B2(n12933), .ZN(
        n12935) );
  NAND2_X1 U15133 ( .A1(n12936), .A2(n12935), .ZN(n13016) );
  MUX2_X1 U15134 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13016), .S(n15016), .Z(
        P3_U3484) );
  AOI22_X1 U15135 ( .A1(n12938), .A2(n8900), .B1(n12979), .B2(n12937), .ZN(
        n12939) );
  NAND2_X1 U15136 ( .A1(n12940), .A2(n12939), .ZN(n13017) );
  MUX2_X1 U15137 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13017), .S(n15016), .Z(
        P3_U3483) );
  OAI22_X1 U15138 ( .A1(n12943), .A2(n14977), .B1(n12942), .B2(n12941), .ZN(
        n12944) );
  MUX2_X1 U15139 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n13018), .S(n15016), .Z(
        P3_U3482) );
  INV_X1 U15140 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12948) );
  AOI21_X1 U15141 ( .B1(n8900), .B2(n12947), .A(n12946), .ZN(n13019) );
  MUX2_X1 U15142 ( .A(n12948), .B(n13019), .S(n15016), .Z(n12949) );
  OAI21_X1 U15143 ( .B1(n13022), .B2(n12996), .A(n12949), .ZN(P3_U3481) );
  INV_X1 U15144 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12952) );
  AOI21_X1 U15145 ( .B1(n8900), .B2(n12951), .A(n12950), .ZN(n13023) );
  MUX2_X1 U15146 ( .A(n12952), .B(n13023), .S(n15016), .Z(n12953) );
  OAI21_X1 U15147 ( .B1(n13026), .B2(n12996), .A(n12953), .ZN(P3_U3480) );
  INV_X1 U15148 ( .A(n12954), .ZN(n13030) );
  NOR2_X1 U15149 ( .A1(n12955), .A2(n14977), .ZN(n12958) );
  AOI21_X1 U15150 ( .B1(n12958), .B2(n12957), .A(n12956), .ZN(n13027) );
  MUX2_X1 U15151 ( .A(n12959), .B(n13027), .S(n15016), .Z(n12960) );
  OAI21_X1 U15152 ( .B1(n13030), .B2(n12996), .A(n12960), .ZN(P3_U3479) );
  NAND2_X1 U15153 ( .A1(n12961), .A2(n8900), .ZN(n12962) );
  NAND2_X1 U15154 ( .A1(n12963), .A2(n12962), .ZN(n13031) );
  INV_X1 U15155 ( .A(n13031), .ZN(n12965) );
  MUX2_X1 U15156 ( .A(n12965), .B(n12964), .S(n15014), .Z(n12966) );
  OAI21_X1 U15157 ( .B1(n12996), .B2(n13034), .A(n12966), .ZN(P3_U3478) );
  INV_X1 U15158 ( .A(n12967), .ZN(n13038) );
  NOR2_X1 U15159 ( .A1(n12968), .A2(n14977), .ZN(n12971) );
  AOI21_X1 U15160 ( .B1(n12971), .B2(n12970), .A(n12969), .ZN(n13035) );
  MUX2_X1 U15161 ( .A(n12972), .B(n13035), .S(n15016), .Z(n12973) );
  OAI21_X1 U15162 ( .B1(n13038), .B2(n12996), .A(n12973), .ZN(P3_U3477) );
  AOI22_X1 U15163 ( .A1(n12975), .A2(n8900), .B1(n12979), .B2(n12974), .ZN(
        n12976) );
  NAND2_X1 U15164 ( .A1(n12977), .A2(n12976), .ZN(n13039) );
  MUX2_X1 U15165 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13039), .S(n15016), .Z(
        P3_U3476) );
  AOI22_X1 U15166 ( .A1(n12980), .A2(n8900), .B1(n12979), .B2(n12978), .ZN(
        n12981) );
  NAND2_X1 U15167 ( .A1(n12982), .A2(n12981), .ZN(n13040) );
  MUX2_X1 U15168 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n13040), .S(n15016), .Z(
        P3_U3475) );
  AOI21_X1 U15169 ( .B1(n12984), .B2(n8900), .A(n12983), .ZN(n13041) );
  MUX2_X1 U15170 ( .A(n12985), .B(n13041), .S(n15016), .Z(n12986) );
  OAI21_X1 U15171 ( .B1(n13044), .B2(n12996), .A(n12986), .ZN(P3_U3474) );
  NAND2_X1 U15172 ( .A1(n12987), .A2(n8900), .ZN(n12988) );
  NAND2_X1 U15173 ( .A1(n12989), .A2(n12988), .ZN(n13045) );
  MUX2_X1 U15174 ( .A(n13045), .B(P3_REG1_REG_14__SCAN_IN), .S(n15014), .Z(
        n12991) );
  NOR2_X1 U15175 ( .A1(n13046), .A2(n12996), .ZN(n12990) );
  AOI21_X1 U15176 ( .B1(n12993), .B2(n8900), .A(n12992), .ZN(n13049) );
  MUX2_X1 U15177 ( .A(n12994), .B(n13049), .S(n15016), .Z(n12995) );
  OAI21_X1 U15178 ( .B1(n12996), .B2(n13052), .A(n12995), .ZN(P3_U3472) );
  INV_X1 U15179 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n13000) );
  NAND2_X1 U15180 ( .A1(n12997), .A2(n8912), .ZN(n12999) );
  NAND2_X1 U15181 ( .A1(n12998), .A2(n15004), .ZN(n13002) );
  OAI211_X1 U15182 ( .C1(n13000), .C2(n15004), .A(n12999), .B(n13002), .ZN(
        P3_U3458) );
  NAND2_X1 U15183 ( .A1(n13001), .A2(n8912), .ZN(n13003) );
  OAI211_X1 U15184 ( .C1(n8891), .C2(n15004), .A(n13003), .B(n13002), .ZN(
        P3_U3457) );
  MUX2_X1 U15185 ( .A(n13005), .B(n13004), .S(n15004), .Z(n13006) );
  OAI21_X1 U15186 ( .B1(n13007), .B2(n13053), .A(n13006), .ZN(P3_U3455) );
  MUX2_X1 U15187 ( .A(n13009), .B(n13008), .S(n15004), .Z(n13010) );
  OAI21_X1 U15188 ( .B1(n13011), .B2(n13053), .A(n13010), .ZN(P3_U3454) );
  MUX2_X1 U15189 ( .A(n13013), .B(n13012), .S(n15004), .Z(n13014) );
  OAI21_X1 U15190 ( .B1(n13015), .B2(n13053), .A(n13014), .ZN(P3_U3453) );
  MUX2_X1 U15191 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n13016), .S(n15004), .Z(
        P3_U3452) );
  MUX2_X1 U15192 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n13017), .S(n15004), .Z(
        P3_U3451) );
  MUX2_X1 U15193 ( .A(n13018), .B(P3_REG0_REG_23__SCAN_IN), .S(n15006), .Z(
        P3_U3450) );
  MUX2_X1 U15194 ( .A(n13020), .B(n13019), .S(n15004), .Z(n13021) );
  OAI21_X1 U15195 ( .B1(n13022), .B2(n13053), .A(n13021), .ZN(P3_U3449) );
  INV_X1 U15196 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13024) );
  MUX2_X1 U15197 ( .A(n13024), .B(n13023), .S(n15004), .Z(n13025) );
  OAI21_X1 U15198 ( .B1(n13026), .B2(n13053), .A(n13025), .ZN(P3_U3448) );
  MUX2_X1 U15199 ( .A(n13028), .B(n13027), .S(n15004), .Z(n13029) );
  OAI21_X1 U15200 ( .B1(n13030), .B2(n13053), .A(n13029), .ZN(P3_U3447) );
  MUX2_X1 U15201 ( .A(n13031), .B(P3_REG0_REG_19__SCAN_IN), .S(n15006), .Z(
        n13032) );
  INV_X1 U15202 ( .A(n13032), .ZN(n13033) );
  OAI21_X1 U15203 ( .B1(n13053), .B2(n13034), .A(n13033), .ZN(P3_U3446) );
  MUX2_X1 U15204 ( .A(n13036), .B(n13035), .S(n15004), .Z(n13037) );
  OAI21_X1 U15205 ( .B1(n13038), .B2(n13053), .A(n13037), .ZN(P3_U3444) );
  MUX2_X1 U15206 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13039), .S(n15004), .Z(
        P3_U3441) );
  MUX2_X1 U15207 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n13040), .S(n15004), .Z(
        P3_U3438) );
  INV_X1 U15208 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13042) );
  MUX2_X1 U15209 ( .A(n13042), .B(n13041), .S(n15004), .Z(n13043) );
  OAI21_X1 U15210 ( .B1(n13044), .B2(n13053), .A(n13043), .ZN(P3_U3435) );
  MUX2_X1 U15211 ( .A(n13045), .B(P3_REG0_REG_14__SCAN_IN), .S(n15006), .Z(
        n13048) );
  NOR2_X1 U15212 ( .A1(n13046), .A2(n13053), .ZN(n13047) );
  INV_X1 U15213 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n13050) );
  MUX2_X1 U15214 ( .A(n13050), .B(n13049), .S(n15004), .Z(n13051) );
  OAI21_X1 U15215 ( .B1(n13053), .B2(n13052), .A(n13051), .ZN(P3_U3429) );
  MUX2_X1 U15216 ( .A(P3_D_REG_1__SCAN_IN), .B(n13054), .S(n13055), .Z(
        P3_U3377) );
  MUX2_X1 U15217 ( .A(P3_D_REG_0__SCAN_IN), .B(n13056), .S(n13055), .Z(
        P3_U3376) );
  NAND3_X1 U15218 ( .A1(n13058), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n13060) );
  INV_X1 U15219 ( .A(SI_31_), .ZN(n15112) );
  OAI22_X1 U15220 ( .A1(n13057), .A2(n13060), .B1(n15112), .B2(n13059), .ZN(
        n13061) );
  AOI21_X1 U15221 ( .B1(n13063), .B2(n13062), .A(n13061), .ZN(n13064) );
  INV_X1 U15222 ( .A(n13064), .ZN(P3_U3264) );
  INV_X1 U15223 ( .A(n13065), .ZN(n13066) );
  OAI222_X1 U15224 ( .A1(n13070), .A2(n13069), .B1(P3_U3151), .B2(n13068), 
        .C1(n13067), .C2(n13066), .ZN(P3_U3267) );
  OAI211_X1 U15225 ( .C1(n13073), .C2(n13072), .A(n13071), .B(n14384), .ZN(
        n13078) );
  INV_X1 U15226 ( .A(n13301), .ZN(n13076) );
  AOI22_X1 U15227 ( .A1(n13167), .A2(n13176), .B1(n13178), .B2(n13166), .ZN(
        n13296) );
  OAI22_X1 U15228 ( .A1(n14660), .A2(n13296), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13074), .ZN(n13075) );
  AOI21_X1 U15229 ( .B1(n13076), .B2(n13159), .A(n13075), .ZN(n13077) );
  OAI211_X1 U15230 ( .C1(n13483), .C2(n13162), .A(n13078), .B(n13077), .ZN(
        P2_U3186) );
  XOR2_X1 U15231 ( .A(n13080), .B(n13079), .Z(n13086) );
  INV_X1 U15232 ( .A(n13180), .ZN(n13081) );
  OAI22_X1 U15233 ( .A1(n13082), .A2(n13142), .B1(n13081), .B2(n13144), .ZN(
        n13364) );
  AOI22_X1 U15234 ( .A1(n13364), .A2(n14386), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13083) );
  OAI21_X1 U15235 ( .B1(n13370), .B2(n14672), .A(n13083), .ZN(n13084) );
  AOI21_X1 U15236 ( .B1(n13505), .B2(n14669), .A(n13084), .ZN(n13085) );
  OAI21_X1 U15237 ( .B1(n13086), .B2(n14664), .A(n13085), .ZN(P2_U3188) );
  INV_X1 U15238 ( .A(n13087), .ZN(n13088) );
  NOR2_X1 U15239 ( .A1(n13089), .A2(n13088), .ZN(n13090) );
  XNOR2_X1 U15240 ( .A(n13091), .B(n13090), .ZN(n13095) );
  AOI22_X1 U15241 ( .A1(n13184), .A2(n13167), .B1(n13166), .B2(n13186), .ZN(
        n13429) );
  NAND2_X1 U15242 ( .A1(n13159), .A2(n13423), .ZN(n13092) );
  NAND2_X1 U15243 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13260)
         );
  OAI211_X1 U15244 ( .C1(n13429), .C2(n14660), .A(n13092), .B(n13260), .ZN(
        n13093) );
  AOI21_X1 U15245 ( .B1(n13528), .B2(n14669), .A(n13093), .ZN(n13094) );
  OAI21_X1 U15246 ( .B1(n13095), .B2(n14664), .A(n13094), .ZN(P2_U3191) );
  INV_X1 U15247 ( .A(n13518), .ZN(n13402) );
  OAI211_X1 U15248 ( .C1(n13098), .C2(n13097), .A(n13096), .B(n14384), .ZN(
        n13103) );
  INV_X1 U15249 ( .A(n13099), .ZN(n13400) );
  AOI22_X1 U15250 ( .A1(n13182), .A2(n13167), .B1(n13166), .B2(n13184), .ZN(
        n13397) );
  OAI22_X1 U15251 ( .A1(n13397), .A2(n14660), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13100), .ZN(n13101) );
  AOI21_X1 U15252 ( .B1(n13400), .B2(n13159), .A(n13101), .ZN(n13102) );
  OAI211_X1 U15253 ( .C1(n13402), .C2(n13162), .A(n13103), .B(n13102), .ZN(
        P2_U3195) );
  OAI211_X1 U15254 ( .C1(n13106), .C2(n13105), .A(n13104), .B(n14384), .ZN(
        n13111) );
  INV_X1 U15255 ( .A(n13332), .ZN(n13109) );
  AOI22_X1 U15256 ( .A1(n13166), .A2(n13180), .B1(n13178), .B2(n13167), .ZN(
        n13326) );
  OAI22_X1 U15257 ( .A1(n14660), .A2(n13326), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13107), .ZN(n13108) );
  AOI21_X1 U15258 ( .B1(n13109), .B2(n13159), .A(n13108), .ZN(n13110) );
  OAI211_X1 U15259 ( .C1(n13491), .C2(n13162), .A(n13111), .B(n13110), .ZN(
        P2_U3197) );
  AND3_X1 U15260 ( .A1(n14381), .A2(n13113), .A3(n13112), .ZN(n13114) );
  OAI21_X1 U15261 ( .B1(n13115), .B2(n13114), .A(n14384), .ZN(n13122) );
  INV_X1 U15262 ( .A(n13116), .ZN(n13120) );
  OAI22_X1 U15263 ( .A1(n13118), .A2(n14660), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13117), .ZN(n13119) );
  AOI21_X1 U15264 ( .B1(n13120), .B2(n13159), .A(n13119), .ZN(n13121) );
  OAI211_X1 U15265 ( .C1(n13123), .C2(n13162), .A(n13122), .B(n13121), .ZN(
        P2_U3200) );
  OAI211_X1 U15266 ( .C1(n13126), .C2(n13125), .A(n13124), .B(n14384), .ZN(
        n13132) );
  INV_X1 U15267 ( .A(n13352), .ZN(n13130) );
  AND2_X1 U15268 ( .A1(n13179), .A2(n13167), .ZN(n13127) );
  AOI21_X1 U15269 ( .B1(n13181), .B2(n13166), .A(n13127), .ZN(n13348) );
  INV_X1 U15270 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13128) );
  OAI22_X1 U15271 ( .A1(n13348), .A2(n14660), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13128), .ZN(n13129) );
  AOI21_X1 U15272 ( .B1(n13130), .B2(n13159), .A(n13129), .ZN(n13131) );
  OAI211_X1 U15273 ( .C1(n13133), .C2(n13162), .A(n13132), .B(n13131), .ZN(
        P2_U3201) );
  NAND2_X1 U15274 ( .A1(n6515), .A2(n13134), .ZN(n13135) );
  XNOR2_X1 U15275 ( .A(n13136), .B(n13135), .ZN(n13141) );
  AOI22_X1 U15276 ( .A1(n13183), .A2(n13167), .B1(n13166), .B2(n13185), .ZN(
        n13409) );
  OAI22_X1 U15277 ( .A1(n13409), .A2(n14660), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13137), .ZN(n13138) );
  AOI21_X1 U15278 ( .B1(n13415), .B2(n13159), .A(n13138), .ZN(n13140) );
  NAND2_X1 U15279 ( .A1(n13523), .A2(n14669), .ZN(n13139) );
  OAI211_X1 U15280 ( .C1(n13141), .C2(n14664), .A(n13140), .B(n13139), .ZN(
        P2_U3205) );
  OAI22_X1 U15281 ( .A1(n13145), .A2(n13144), .B1(n13143), .B2(n13142), .ZN(
        n13379) );
  AOI22_X1 U15282 ( .A1(n13379), .A2(n14386), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13146) );
  OAI21_X1 U15283 ( .B1(n13386), .B2(n14672), .A(n13146), .ZN(n13151) );
  AOI211_X1 U15284 ( .C1(n13149), .C2(n13148), .A(n14664), .B(n13147), .ZN(
        n13150) );
  AOI211_X1 U15285 ( .C1(n13511), .C2(n14669), .A(n13151), .B(n13150), .ZN(
        n13152) );
  INV_X1 U15286 ( .A(n13152), .ZN(P2_U3207) );
  INV_X1 U15287 ( .A(n13532), .ZN(n13444) );
  OAI211_X1 U15288 ( .C1(n13155), .C2(n13154), .A(n13153), .B(n14384), .ZN(
        n13161) );
  INV_X1 U15289 ( .A(n13156), .ZN(n13441) );
  AOI22_X1 U15290 ( .A1(n13185), .A2(n13167), .B1(n13166), .B2(n13187), .ZN(
        n13435) );
  OAI21_X1 U15291 ( .B1(n13435), .B2(n14660), .A(n13157), .ZN(n13158) );
  AOI21_X1 U15292 ( .B1(n13441), .B2(n13159), .A(n13158), .ZN(n13160) );
  OAI211_X1 U15293 ( .C1(n13444), .C2(n13162), .A(n13161), .B(n13160), .ZN(
        P2_U3210) );
  AOI21_X1 U15294 ( .B1(n13165), .B2(n13164), .A(n13163), .ZN(n13173) );
  NAND2_X1 U15295 ( .A1(n13179), .A2(n13166), .ZN(n13169) );
  NAND2_X1 U15296 ( .A1(n13177), .A2(n13167), .ZN(n13168) );
  NAND2_X1 U15297 ( .A1(n13169), .A2(n13168), .ZN(n13320) );
  AOI22_X1 U15298 ( .A1(n14386), .A2(n13320), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13170) );
  OAI21_X1 U15299 ( .B1(n14672), .B2(n13313), .A(n13170), .ZN(n13171) );
  AOI21_X1 U15300 ( .B1(n13487), .B2(n14669), .A(n13171), .ZN(n13172) );
  OAI21_X1 U15301 ( .B1(n13173), .B2(n14664), .A(n13172), .ZN(P2_U3212) );
  MUX2_X1 U15302 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13265), .S(n6480), .Z(
        P2_U3562) );
  MUX2_X1 U15303 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13174), .S(n6480), .Z(
        P2_U3561) );
  MUX2_X1 U15304 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13175), .S(n6480), .Z(
        P2_U3560) );
  MUX2_X1 U15305 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13176), .S(n6480), .Z(
        P2_U3559) );
  MUX2_X1 U15306 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13177), .S(n6480), .Z(
        P2_U3558) );
  MUX2_X1 U15307 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13178), .S(n6480), .Z(
        P2_U3557) );
  MUX2_X1 U15308 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13179), .S(n6480), .Z(
        P2_U3556) );
  MUX2_X1 U15309 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13180), .S(n6480), .Z(
        P2_U3555) );
  MUX2_X1 U15310 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13181), .S(n6480), .Z(
        P2_U3554) );
  MUX2_X1 U15311 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13182), .S(n6480), .Z(
        P2_U3553) );
  MUX2_X1 U15312 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13183), .S(n6480), .Z(
        P2_U3552) );
  MUX2_X1 U15313 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13184), .S(n6480), .Z(
        P2_U3551) );
  MUX2_X1 U15314 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13185), .S(n6480), .Z(
        P2_U3550) );
  MUX2_X1 U15315 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13186), .S(n6480), .Z(
        P2_U3549) );
  MUX2_X1 U15316 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13187), .S(n6480), .Z(
        P2_U3548) );
  MUX2_X1 U15317 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13188), .S(n6480), .Z(
        P2_U3547) );
  MUX2_X1 U15318 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13189), .S(n6480), .Z(
        P2_U3546) );
  MUX2_X1 U15319 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13190), .S(n6480), .Z(
        P2_U3545) );
  MUX2_X1 U15320 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13191), .S(n6480), .Z(
        P2_U3544) );
  MUX2_X1 U15321 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13192), .S(n6480), .Z(
        P2_U3543) );
  MUX2_X1 U15322 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13193), .S(n6480), .Z(
        P2_U3542) );
  MUX2_X1 U15323 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13194), .S(n6480), .Z(
        P2_U3541) );
  MUX2_X1 U15324 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13195), .S(n6480), .Z(
        P2_U3540) );
  MUX2_X1 U15325 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13196), .S(n6480), .Z(
        P2_U3539) );
  MUX2_X1 U15326 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13197), .S(n6480), .Z(
        P2_U3538) );
  MUX2_X1 U15327 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13198), .S(n6480), .Z(
        P2_U3537) );
  MUX2_X1 U15328 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13199), .S(n6480), .Z(
        P2_U3536) );
  MUX2_X1 U15329 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13200), .S(n6480), .Z(
        P2_U3535) );
  MUX2_X1 U15330 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13201), .S(n6480), .Z(
        P2_U3534) );
  MUX2_X1 U15331 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n10068), .S(n6480), .Z(
        P2_U3533) );
  MUX2_X1 U15332 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n13202), .S(n6480), .Z(
        P2_U3532) );
  MUX2_X1 U15333 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n13203), .S(n6480), .Z(
        P2_U3531) );
  AND3_X1 U15334 ( .A1(n14697), .A2(n13205), .A3(n13204), .ZN(n13206) );
  NOR3_X1 U15335 ( .A1(n14713), .A2(n13207), .A3(n13206), .ZN(n13208) );
  AOI21_X1 U15336 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(n14775), .A(n13208), .ZN(
        n13218) );
  INV_X1 U15337 ( .A(n13209), .ZN(n13217) );
  NAND2_X1 U15338 ( .A1(n14776), .A2(n13210), .ZN(n13216) );
  MUX2_X1 U15339 ( .A(n9832), .B(P2_REG1_REG_4__SCAN_IN), .S(n13210), .Z(
        n13211) );
  NAND3_X1 U15340 ( .A1(n14700), .A2(n13212), .A3(n13211), .ZN(n13213) );
  NAND3_X1 U15341 ( .A1(n14783), .A2(n13214), .A3(n13213), .ZN(n13215) );
  NAND4_X1 U15342 ( .A1(n13218), .A2(n13217), .A3(n13216), .A4(n13215), .ZN(
        P2_U3218) );
  OAI21_X1 U15343 ( .B1(n13220), .B2(n13219), .A(n14742), .ZN(n13221) );
  NAND2_X1 U15344 ( .A1(n13221), .A2(n14778), .ZN(n13232) );
  AOI21_X1 U15345 ( .B1(n14775), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n13222), 
        .ZN(n13231) );
  MUX2_X1 U15346 ( .A(n10981), .B(P2_REG1_REG_11__SCAN_IN), .S(n13228), .Z(
        n13223) );
  NAND3_X1 U15347 ( .A1(n13225), .A2(n13224), .A3(n13223), .ZN(n13226) );
  NAND3_X1 U15348 ( .A1(n13227), .A2(n14783), .A3(n13226), .ZN(n13230) );
  NAND2_X1 U15349 ( .A1(n14776), .A2(n13228), .ZN(n13229) );
  NAND4_X1 U15350 ( .A1(n13232), .A2(n13231), .A3(n13230), .A4(n13229), .ZN(
        P2_U3225) );
  OAI211_X1 U15351 ( .C1(n13235), .C2(n13234), .A(n14778), .B(n13233), .ZN(
        n13243) );
  AOI22_X1 U15352 ( .A1(n14776), .A2(n13236), .B1(n14775), .B2(
        P2_ADDR_REG_16__SCAN_IN), .ZN(n13242) );
  NAND2_X1 U15353 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n14389)
         );
  OAI211_X1 U15354 ( .C1(n13239), .C2(n13238), .A(n14783), .B(n13237), .ZN(
        n13240) );
  AND2_X1 U15355 ( .A1(n14389), .A2(n13240), .ZN(n13241) );
  NAND3_X1 U15356 ( .A1(n13243), .A2(n13242), .A3(n13241), .ZN(P2_U3230) );
  NOR2_X1 U15357 ( .A1(n13249), .A2(n13244), .ZN(n13246) );
  NOR2_X1 U15358 ( .A1(n13246), .A2(n13245), .ZN(n13247) );
  NAND2_X1 U15359 ( .A1(n13249), .A2(n13248), .ZN(n13250) );
  NAND2_X1 U15360 ( .A1(n13251), .A2(n13250), .ZN(n13252) );
  XOR2_X1 U15361 ( .A(n13252), .B(P2_REG1_REG_19__SCAN_IN), .Z(n13255) );
  NOR2_X1 U15362 ( .A1(n13255), .A2(n14746), .ZN(n13253) );
  AOI211_X1 U15363 ( .C1(n13254), .C2(n14778), .A(n14776), .B(n13253), .ZN(
        n13259) );
  AOI22_X1 U15364 ( .A1(n13256), .A2(n14778), .B1(n14783), .B2(n13255), .ZN(
        n13258) );
  MUX2_X1 U15365 ( .A(n13259), .B(n13258), .S(n13257), .Z(n13261) );
  OAI211_X1 U15366 ( .C1(n13262), .C2(n14752), .A(n13261), .B(n13260), .ZN(
        P2_U3233) );
  NOR2_X2 U15367 ( .A1(n13270), .A2(n13269), .ZN(n13271) );
  XNOR2_X1 U15368 ( .A(n13263), .B(n13271), .ZN(n13264) );
  NAND2_X1 U15369 ( .A1(n13264), .A2(n11850), .ZN(n13466) );
  NAND2_X1 U15370 ( .A1(n13266), .A2(n13265), .ZN(n13467) );
  NOR2_X1 U15371 ( .A1(n13453), .A2(n13467), .ZN(n13275) );
  NOR2_X1 U15372 ( .A1(n8141), .A2(n13443), .ZN(n13267) );
  AOI211_X1 U15373 ( .C1(n13453), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13275), 
        .B(n13267), .ZN(n13268) );
  OAI21_X1 U15374 ( .B1(n13466), .B2(n13391), .A(n13268), .ZN(P2_U3234) );
  INV_X1 U15375 ( .A(n13270), .ZN(n13273) );
  INV_X1 U15376 ( .A(n13271), .ZN(n13272) );
  OAI211_X1 U15377 ( .C1(n13469), .C2(n13273), .A(n13272), .B(n11850), .ZN(
        n13468) );
  NOR2_X1 U15378 ( .A1(n13469), .A2(n13443), .ZN(n13274) );
  AOI211_X1 U15379 ( .C1(n13453), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13275), 
        .B(n13274), .ZN(n13276) );
  OAI21_X1 U15380 ( .B1(n13391), .B2(n13468), .A(n13276), .ZN(P2_U3235) );
  NOR2_X1 U15381 ( .A1(n13277), .A2(n13430), .ZN(n13281) );
  OAI21_X1 U15382 ( .B1(n13294), .B2(n13278), .A(n13283), .ZN(n13280) );
  OAI21_X1 U15383 ( .B1(n13284), .B2(n13283), .A(n13282), .ZN(n13478) );
  OAI22_X1 U15384 ( .A1(n13432), .A2(n13286), .B1(n13285), .B2(n13385), .ZN(
        n13287) );
  AOI21_X1 U15385 ( .B1(n13475), .B2(n13460), .A(n13287), .ZN(n13291) );
  AOI21_X1 U15386 ( .B1(n13475), .B2(n6538), .A(n13412), .ZN(n13289) );
  AND2_X1 U15387 ( .A1(n13289), .A2(n13288), .ZN(n13474) );
  NAND2_X1 U15388 ( .A1(n13474), .A2(n13455), .ZN(n13290) );
  OAI211_X1 U15389 ( .C1(n13478), .C2(n13449), .A(n13291), .B(n13290), .ZN(
        n13292) );
  INV_X1 U15390 ( .A(n13292), .ZN(n13293) );
  OAI21_X1 U15391 ( .B1(n13453), .B2(n13477), .A(n13293), .ZN(P2_U3237) );
  AOI21_X1 U15392 ( .B1(n13299), .B2(n13295), .A(n13294), .ZN(n13297) );
  OAI21_X1 U15393 ( .B1(n13297), .B2(n13430), .A(n13296), .ZN(n13484) );
  AOI21_X1 U15394 ( .B1(n13304), .B2(n13310), .A(n13412), .ZN(n13298) );
  NAND2_X1 U15395 ( .A1(n13298), .A2(n6538), .ZN(n13481) );
  OR2_X1 U15396 ( .A1(n13300), .A2(n13299), .ZN(n13480) );
  NAND3_X1 U15397 ( .A1(n13480), .A2(n13479), .A3(n13457), .ZN(n13306) );
  OAI22_X1 U15398 ( .A1(n13432), .A2(n13302), .B1(n13301), .B2(n13385), .ZN(
        n13303) );
  AOI21_X1 U15399 ( .B1(n13304), .B2(n13460), .A(n13303), .ZN(n13305) );
  OAI211_X1 U15400 ( .C1(n13481), .C2(n13391), .A(n13306), .B(n13305), .ZN(
        n13307) );
  AOI21_X1 U15401 ( .B1(n13432), .B2(n13484), .A(n13307), .ZN(n13308) );
  INV_X1 U15402 ( .A(n13308), .ZN(P2_U3238) );
  XNOR2_X1 U15403 ( .A(n13309), .B(n13318), .ZN(n13489) );
  INV_X1 U15404 ( .A(n13310), .ZN(n13311) );
  AOI211_X1 U15405 ( .C1(n13487), .C2(n13331), .A(n13412), .B(n13311), .ZN(
        n13486) );
  NOR2_X1 U15406 ( .A1(n13312), .A2(n13443), .ZN(n13316) );
  OAI22_X1 U15407 ( .A1(n13432), .A2(n13314), .B1(n13313), .B2(n13385), .ZN(
        n13315) );
  AOI211_X1 U15408 ( .C1(n13486), .C2(n13455), .A(n13316), .B(n13315), .ZN(
        n13324) );
  OAI211_X1 U15409 ( .C1(n13319), .C2(n13318), .A(n13317), .B(n13437), .ZN(
        n13322) );
  INV_X1 U15410 ( .A(n13320), .ZN(n13321) );
  NAND2_X1 U15411 ( .A1(n13322), .A2(n13321), .ZN(n13485) );
  NAND2_X1 U15412 ( .A1(n13485), .A2(n13432), .ZN(n13323) );
  OAI211_X1 U15413 ( .C1(n13489), .C2(n13449), .A(n13324), .B(n13323), .ZN(
        P2_U3239) );
  XNOR2_X1 U15414 ( .A(n13325), .B(n13329), .ZN(n13327) );
  OAI21_X1 U15415 ( .B1(n13327), .B2(n13430), .A(n13326), .ZN(n13493) );
  INV_X1 U15416 ( .A(n13493), .ZN(n13339) );
  OAI21_X1 U15417 ( .B1(n13330), .B2(n13329), .A(n13328), .ZN(n13494) );
  OAI211_X1 U15418 ( .C1(n13491), .C2(n13356), .A(n11850), .B(n13331), .ZN(
        n13490) );
  OAI22_X1 U15419 ( .A1(n13432), .A2(n13333), .B1(n13332), .B2(n13385), .ZN(
        n13334) );
  AOI21_X1 U15420 ( .B1(n13335), .B2(n13460), .A(n13334), .ZN(n13336) );
  OAI21_X1 U15421 ( .B1(n13490), .B2(n13391), .A(n13336), .ZN(n13337) );
  AOI21_X1 U15422 ( .B1(n13494), .B2(n13457), .A(n13337), .ZN(n13338) );
  OAI21_X1 U15423 ( .B1(n13453), .B2(n13339), .A(n13338), .ZN(P2_U3240) );
  AND2_X1 U15424 ( .A1(n13341), .A2(n13340), .ZN(n13343) );
  NAND2_X1 U15425 ( .A1(n13345), .A2(n13344), .ZN(n13346) );
  NAND2_X1 U15426 ( .A1(n13347), .A2(n13346), .ZN(n13350) );
  INV_X1 U15427 ( .A(n13348), .ZN(n13349) );
  AOI21_X1 U15428 ( .B1(n13350), .B2(n13437), .A(n13349), .ZN(n13351) );
  OAI21_X1 U15429 ( .B1(n13499), .B2(n10179), .A(n13351), .ZN(n13501) );
  NAND2_X1 U15430 ( .A1(n13501), .A2(n13432), .ZN(n13360) );
  OAI22_X1 U15431 ( .A1(n13432), .A2(n13353), .B1(n13352), .B2(n13385), .ZN(
        n13358) );
  NAND2_X1 U15432 ( .A1(n13496), .A2(n13372), .ZN(n13354) );
  NAND2_X1 U15433 ( .A1(n13354), .A2(n11850), .ZN(n13355) );
  OR2_X1 U15434 ( .A1(n13356), .A2(n13355), .ZN(n13497) );
  NOR2_X1 U15435 ( .A1(n13497), .A2(n13391), .ZN(n13357) );
  AOI211_X1 U15436 ( .C1(n13460), .C2(n13496), .A(n13358), .B(n13357), .ZN(
        n13359) );
  OAI211_X1 U15437 ( .C1(n13499), .C2(n13361), .A(n13360), .B(n13359), .ZN(
        P2_U3241) );
  XNOR2_X1 U15438 ( .A(n13363), .B(n13362), .ZN(n13365) );
  AOI21_X1 U15439 ( .B1(n13365), .B2(n13437), .A(n13364), .ZN(n13507) );
  OAI21_X1 U15440 ( .B1(n6976), .B2(n13367), .A(n13366), .ZN(n13368) );
  INV_X1 U15441 ( .A(n13368), .ZN(n13508) );
  INV_X1 U15442 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13369) );
  OAI22_X1 U15443 ( .A1(n13370), .A2(n13385), .B1(n13432), .B2(n13369), .ZN(
        n13371) );
  AOI21_X1 U15444 ( .B1(n13505), .B2(n13460), .A(n13371), .ZN(n13375) );
  AOI21_X1 U15445 ( .B1(n13381), .B2(n13505), .A(n13412), .ZN(n13373) );
  AND2_X1 U15446 ( .A1(n13373), .A2(n13372), .ZN(n13504) );
  NAND2_X1 U15447 ( .A1(n13504), .A2(n13455), .ZN(n13374) );
  OAI211_X1 U15448 ( .C1(n13508), .C2(n13449), .A(n13375), .B(n13374), .ZN(
        n13376) );
  INV_X1 U15449 ( .A(n13376), .ZN(n13377) );
  OAI21_X1 U15450 ( .B1(n13453), .B2(n13507), .A(n13377), .ZN(P2_U3242) );
  XNOR2_X1 U15451 ( .A(n13378), .B(n13383), .ZN(n13380) );
  AOI21_X1 U15452 ( .B1(n13380), .B2(n13437), .A(n13379), .ZN(n13514) );
  OAI211_X1 U15453 ( .C1(n13399), .C2(n13382), .A(n11850), .B(n13381), .ZN(
        n13513) );
  NAND2_X1 U15454 ( .A1(n13384), .A2(n13383), .ZN(n13509) );
  NAND3_X1 U15455 ( .A1(n13510), .A2(n13509), .A3(n13457), .ZN(n13390) );
  INV_X1 U15456 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13387) );
  OAI22_X1 U15457 ( .A1(n13432), .A2(n13387), .B1(n13386), .B2(n13385), .ZN(
        n13388) );
  AOI21_X1 U15458 ( .B1(n13511), .B2(n13460), .A(n13388), .ZN(n13389) );
  OAI211_X1 U15459 ( .C1(n13513), .C2(n13391), .A(n13390), .B(n13389), .ZN(
        n13392) );
  INV_X1 U15460 ( .A(n13392), .ZN(n13393) );
  OAI21_X1 U15461 ( .B1(n13514), .B2(n13453), .A(n13393), .ZN(P2_U3243) );
  XOR2_X1 U15462 ( .A(n13394), .B(n13395), .Z(n13520) );
  XOR2_X1 U15463 ( .A(n13396), .B(n13395), .Z(n13398) );
  OAI21_X1 U15464 ( .B1(n13398), .B2(n13430), .A(n13397), .ZN(n13516) );
  NAND2_X1 U15465 ( .A1(n13516), .A2(n13432), .ZN(n13405) );
  AOI211_X1 U15466 ( .C1(n13518), .C2(n13413), .A(n13412), .B(n13399), .ZN(
        n13517) );
  AOI22_X1 U15467 ( .A1(n13453), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13400), 
        .B2(n13458), .ZN(n13401) );
  OAI21_X1 U15468 ( .B1(n13402), .B2(n13443), .A(n13401), .ZN(n13403) );
  AOI21_X1 U15469 ( .B1(n13517), .B2(n13455), .A(n13403), .ZN(n13404) );
  OAI211_X1 U15470 ( .C1(n13520), .C2(n13449), .A(n13405), .B(n13404), .ZN(
        P2_U3244) );
  XNOR2_X1 U15471 ( .A(n13406), .B(n13408), .ZN(n13525) );
  XNOR2_X1 U15472 ( .A(n13407), .B(n13408), .ZN(n13410) );
  OAI21_X1 U15473 ( .B1(n13410), .B2(n13430), .A(n13409), .ZN(n13521) );
  NAND2_X1 U15474 ( .A1(n13521), .A2(n13432), .ZN(n13420) );
  AOI21_X1 U15475 ( .B1(n13422), .B2(n13523), .A(n13412), .ZN(n13414) );
  AND2_X1 U15476 ( .A1(n13414), .A2(n13413), .ZN(n13522) );
  NAND2_X1 U15477 ( .A1(n13523), .A2(n13460), .ZN(n13417) );
  AOI22_X1 U15478 ( .A1(n13453), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13415), 
        .B2(n13458), .ZN(n13416) );
  NAND2_X1 U15479 ( .A1(n13417), .A2(n13416), .ZN(n13418) );
  AOI21_X1 U15480 ( .B1(n13522), .B2(n13455), .A(n13418), .ZN(n13419) );
  OAI211_X1 U15481 ( .C1(n13525), .C2(n13449), .A(n13420), .B(n13419), .ZN(
        P2_U3245) );
  XNOR2_X1 U15482 ( .A(n13421), .B(n13427), .ZN(n13530) );
  AOI211_X1 U15483 ( .C1(n13528), .C2(n13439), .A(n13412), .B(n13411), .ZN(
        n13527) );
  AOI22_X1 U15484 ( .A1(n13453), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13423), 
        .B2(n13458), .ZN(n13424) );
  OAI21_X1 U15485 ( .B1(n13425), .B2(n13443), .A(n13424), .ZN(n13426) );
  AOI21_X1 U15486 ( .B1(n13527), .B2(n13455), .A(n13426), .ZN(n13434) );
  XOR2_X1 U15487 ( .A(n13428), .B(n13427), .Z(n13431) );
  OAI21_X1 U15488 ( .B1(n13431), .B2(n13430), .A(n13429), .ZN(n13526) );
  NAND2_X1 U15489 ( .A1(n13526), .A2(n13432), .ZN(n13433) );
  OAI211_X1 U15490 ( .C1(n13530), .C2(n13449), .A(n13434), .B(n13433), .ZN(
        P2_U3246) );
  XNOR2_X1 U15491 ( .A(n13448), .B(n6615), .ZN(n13438) );
  INV_X1 U15492 ( .A(n13435), .ZN(n13436) );
  AOI21_X1 U15493 ( .B1(n13438), .B2(n13437), .A(n13436), .ZN(n13533) );
  AOI211_X1 U15494 ( .C1(n13532), .C2(n13440), .A(n13412), .B(n6958), .ZN(
        n13531) );
  AOI22_X1 U15495 ( .A1(n13453), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13441), 
        .B2(n13458), .ZN(n13442) );
  OAI21_X1 U15496 ( .B1(n13444), .B2(n13443), .A(n13442), .ZN(n13451) );
  INV_X1 U15497 ( .A(n13445), .ZN(n13446) );
  AOI21_X1 U15498 ( .B1(n13448), .B2(n13447), .A(n13446), .ZN(n13535) );
  NOR2_X1 U15499 ( .A1(n13535), .A2(n13449), .ZN(n13450) );
  AOI211_X1 U15500 ( .C1(n13531), .C2(n13455), .A(n13451), .B(n13450), .ZN(
        n13452) );
  OAI21_X1 U15501 ( .B1(n13453), .B2(n13533), .A(n13452), .ZN(P2_U3247) );
  AOI22_X1 U15502 ( .A1(n13457), .A2(n13456), .B1(n13455), .B2(n13454), .ZN(
        n13465) );
  AOI22_X1 U15503 ( .A1(n13460), .A2(n13459), .B1(n13458), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n13464) );
  MUX2_X1 U15504 ( .A(n13462), .B(n13461), .S(n13432), .Z(n13463) );
  NAND3_X1 U15505 ( .A1(n13465), .A2(n13464), .A3(n13463), .ZN(P2_U3263) );
  OAI211_X1 U15506 ( .C1(n8141), .C2(n14837), .A(n13466), .B(n13467), .ZN(
        n13557) );
  MUX2_X1 U15507 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13557), .S(n14855), .Z(
        P2_U3530) );
  OAI211_X1 U15508 ( .C1(n13469), .C2(n14837), .A(n13468), .B(n13467), .ZN(
        n13558) );
  MUX2_X1 U15509 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13558), .S(n14855), .Z(
        P2_U3529) );
  AOI21_X1 U15510 ( .B1(n14816), .B2(n13475), .A(n13474), .ZN(n13476) );
  OAI211_X1 U15511 ( .C1(n13478), .C2(n14812), .A(n13477), .B(n13476), .ZN(
        n13560) );
  MUX2_X1 U15512 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13560), .S(n14855), .Z(
        P2_U3527) );
  NAND3_X1 U15513 ( .A1(n13480), .A2(n13479), .A3(n14833), .ZN(n13482) );
  MUX2_X1 U15514 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13561), .S(n14855), .Z(
        P2_U3526) );
  AOI211_X1 U15515 ( .C1(n14816), .C2(n13487), .A(n13486), .B(n13485), .ZN(
        n13488) );
  OAI21_X1 U15516 ( .B1(n13489), .B2(n14812), .A(n13488), .ZN(n13562) );
  MUX2_X1 U15517 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13562), .S(n14855), .Z(
        P2_U3525) );
  OAI21_X1 U15518 ( .B1(n13491), .B2(n14837), .A(n13490), .ZN(n13492) );
  AOI211_X1 U15519 ( .C1(n13494), .C2(n14833), .A(n13493), .B(n13492), .ZN(
        n13495) );
  INV_X1 U15520 ( .A(n13495), .ZN(n13563) );
  MUX2_X1 U15521 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13563), .S(n14855), .Z(
        P2_U3524) );
  INV_X1 U15522 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n13502) );
  NAND2_X1 U15523 ( .A1(n13496), .A2(n14816), .ZN(n13498) );
  OAI211_X1 U15524 ( .C1(n13499), .C2(n14819), .A(n13498), .B(n13497), .ZN(
        n13500) );
  NOR2_X1 U15525 ( .A1(n13501), .A2(n13500), .ZN(n13564) );
  MUX2_X1 U15526 ( .A(n13502), .B(n13564), .S(n14855), .Z(n13503) );
  INV_X1 U15527 ( .A(n13503), .ZN(P2_U3523) );
  AOI21_X1 U15528 ( .B1(n14816), .B2(n13505), .A(n13504), .ZN(n13506) );
  OAI211_X1 U15529 ( .C1(n13508), .C2(n14812), .A(n13507), .B(n13506), .ZN(
        n13567) );
  MUX2_X1 U15530 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13567), .S(n14855), .Z(
        P2_U3522) );
  NAND3_X1 U15531 ( .A1(n13510), .A2(n14833), .A3(n13509), .ZN(n13515) );
  NAND2_X1 U15532 ( .A1(n13511), .A2(n14816), .ZN(n13512) );
  NAND4_X1 U15533 ( .A1(n13515), .A2(n13514), .A3(n13513), .A4(n13512), .ZN(
        n13568) );
  MUX2_X1 U15534 ( .A(n13568), .B(P2_REG1_REG_22__SCAN_IN), .S(n14853), .Z(
        P2_U3521) );
  AOI211_X1 U15535 ( .C1(n14816), .C2(n13518), .A(n13517), .B(n13516), .ZN(
        n13519) );
  OAI21_X1 U15536 ( .B1(n14812), .B2(n13520), .A(n13519), .ZN(n13569) );
  MUX2_X1 U15537 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13569), .S(n14855), .Z(
        P2_U3520) );
  AOI211_X1 U15538 ( .C1(n14816), .C2(n13523), .A(n13522), .B(n13521), .ZN(
        n13524) );
  OAI21_X1 U15539 ( .B1(n14812), .B2(n13525), .A(n13524), .ZN(n13570) );
  MUX2_X1 U15540 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13570), .S(n14855), .Z(
        P2_U3519) );
  AOI211_X1 U15541 ( .C1(n14816), .C2(n13528), .A(n13527), .B(n13526), .ZN(
        n13529) );
  OAI21_X1 U15542 ( .B1(n14812), .B2(n13530), .A(n13529), .ZN(n13571) );
  MUX2_X1 U15543 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13571), .S(n14855), .Z(
        P2_U3518) );
  AOI21_X1 U15544 ( .B1(n14816), .B2(n13532), .A(n13531), .ZN(n13534) );
  OAI211_X1 U15545 ( .C1(n14812), .C2(n13535), .A(n13534), .B(n13533), .ZN(
        n13572) );
  MUX2_X1 U15546 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13572), .S(n14855), .Z(
        P2_U3517) );
  AOI21_X1 U15547 ( .B1(n14816), .B2(n13537), .A(n13536), .ZN(n13538) );
  OAI211_X1 U15548 ( .C1(n13540), .C2(n14812), .A(n13539), .B(n13538), .ZN(
        n13573) );
  MUX2_X1 U15549 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13573), .S(n14855), .Z(
        P2_U3516) );
  AOI21_X1 U15550 ( .B1(n14816), .B2(n14388), .A(n13541), .ZN(n13543) );
  OAI211_X1 U15551 ( .C1(n14812), .C2(n13544), .A(n13543), .B(n13542), .ZN(
        n13574) );
  MUX2_X1 U15552 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13574), .S(n14855), .Z(
        P2_U3515) );
  AOI21_X1 U15553 ( .B1(n14816), .B2(n13546), .A(n13545), .ZN(n13548) );
  OAI211_X1 U15554 ( .C1(n13549), .C2(n14812), .A(n13548), .B(n13547), .ZN(
        n13575) );
  MUX2_X1 U15555 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13575), .S(n14855), .Z(
        P2_U3514) );
  AOI21_X1 U15556 ( .B1(n14816), .B2(n6677), .A(n13550), .ZN(n13555) );
  NAND3_X1 U15557 ( .A1(n13552), .A2(n13551), .A3(n14833), .ZN(n13553) );
  NAND3_X1 U15558 ( .A1(n13555), .A2(n13554), .A3(n13553), .ZN(n13576) );
  MUX2_X1 U15559 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13576), .S(n14855), .Z(
        P2_U3513) );
  MUX2_X1 U15560 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n13556), .S(n14855), .Z(
        P2_U3501) );
  MUX2_X1 U15561 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13557), .S(n14835), .Z(
        P2_U3498) );
  MUX2_X1 U15562 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13558), .S(n14835), .Z(
        P2_U3497) );
  MUX2_X1 U15563 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13560), .S(n14835), .Z(
        P2_U3495) );
  MUX2_X1 U15564 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13561), .S(n14835), .Z(
        P2_U3494) );
  MUX2_X1 U15565 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13562), .S(n14835), .Z(
        P2_U3493) );
  MUX2_X1 U15566 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13563), .S(n14835), .Z(
        P2_U3492) );
  MUX2_X1 U15567 ( .A(n13565), .B(n13564), .S(n14835), .Z(n13566) );
  INV_X1 U15568 ( .A(n13566), .ZN(P2_U3491) );
  MUX2_X1 U15569 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13567), .S(n14835), .Z(
        P2_U3490) );
  MUX2_X1 U15570 ( .A(n13568), .B(P2_REG0_REG_22__SCAN_IN), .S(n14844), .Z(
        P2_U3489) );
  MUX2_X1 U15571 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13569), .S(n14835), .Z(
        P2_U3488) );
  MUX2_X1 U15572 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13570), .S(n14835), .Z(
        P2_U3487) );
  MUX2_X1 U15573 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13571), .S(n14835), .Z(
        P2_U3486) );
  MUX2_X1 U15574 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13572), .S(n14835), .Z(
        P2_U3484) );
  MUX2_X1 U15575 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13573), .S(n14835), .Z(
        P2_U3481) );
  MUX2_X1 U15576 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13574), .S(n14835), .Z(
        P2_U3478) );
  MUX2_X1 U15577 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13575), .S(n14835), .Z(
        P2_U3475) );
  MUX2_X1 U15578 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13576), .S(n14835), .Z(
        P2_U3472) );
  INV_X1 U15579 ( .A(n9563), .ZN(n13580) );
  NOR4_X1 U15580 ( .A1(n13577), .A2(P2_IR_REG_30__SCAN_IN), .A3(n7445), .A4(
        P2_U3088), .ZN(n13578) );
  AOI21_X1 U15581 ( .B1(n13585), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13578), 
        .ZN(n13579) );
  OAI21_X1 U15582 ( .B1(n13580), .B2(n13587), .A(n13579), .ZN(P2_U3296) );
  INV_X1 U15583 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13581) );
  OAI222_X1 U15584 ( .A1(n13587), .A2(n13583), .B1(P2_U3088), .B2(n13582), 
        .C1(n13581), .C2(n13593), .ZN(P2_U3298) );
  AOI21_X1 U15585 ( .B1(n13585), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13584), 
        .ZN(n13586) );
  OAI21_X1 U15586 ( .B1(n13588), .B2(n13587), .A(n13586), .ZN(P2_U3299) );
  INV_X1 U15587 ( .A(n13589), .ZN(n14185) );
  OAI222_X1 U15588 ( .A1(n13593), .A2(n13591), .B1(n13587), .B2(n14185), .C1(
        n13590), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U15589 ( .A(n13592), .ZN(n14187) );
  OAI222_X1 U15590 ( .A1(n13595), .A2(P2_U3088), .B1(n13587), .B2(n14187), 
        .C1(n13594), .C2(n13593), .ZN(P2_U3301) );
  MUX2_X1 U15591 ( .A(n6499), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  AOI22_X1 U15592 ( .A1(n13685), .A2(n13871), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13598) );
  NAND2_X1 U15593 ( .A1(n13729), .A2(n13872), .ZN(n13597) );
  OAI211_X1 U15594 ( .C1(n14436), .C2(n13873), .A(n13598), .B(n13597), .ZN(
        n13599) );
  AOI21_X1 U15595 ( .B1(n14084), .B2(n14432), .A(n13599), .ZN(n13600) );
  OAI21_X1 U15596 ( .B1(n13601), .B2(n14426), .A(n13600), .ZN(P1_U3214) );
  XOR2_X1 U15597 ( .A(n13603), .B(n13602), .Z(n13609) );
  OR2_X1 U15598 ( .A1(n13622), .A2(n14542), .ZN(n13605) );
  NAND2_X1 U15599 ( .A1(n13741), .A2(n14055), .ZN(n13604) );
  NAND2_X1 U15600 ( .A1(n13605), .A2(n13604), .ZN(n14107) );
  AOI22_X1 U15601 ( .A1(n14414), .A2(n14107), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13606) );
  OAI21_X1 U15602 ( .B1(n14436), .B2(n13943), .A(n13606), .ZN(n13607) );
  AOI21_X1 U15603 ( .B1(n14108), .B2(n14432), .A(n13607), .ZN(n13608) );
  OAI21_X1 U15604 ( .B1(n13609), .B2(n14426), .A(n13608), .ZN(P1_U3216) );
  INV_X1 U15605 ( .A(n14136), .ZN(n14008) );
  AOI21_X1 U15606 ( .B1(n13610), .B2(n13611), .A(n14426), .ZN(n13613) );
  NAND2_X1 U15607 ( .A1(n13613), .A2(n13612), .ZN(n13617) );
  NOR2_X1 U15608 ( .A1(n14436), .A2(n14004), .ZN(n13615) );
  NAND2_X1 U15609 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13829)
         );
  OAI21_X1 U15610 ( .B1(n14422), .B2(n13623), .A(n13829), .ZN(n13614) );
  AOI211_X1 U15611 ( .C1(n13685), .C2(n14034), .A(n13615), .B(n13614), .ZN(
        n13616) );
  OAI211_X1 U15612 ( .C1(n14008), .C2(n13737), .A(n13617), .B(n13616), .ZN(
        P1_U3219) );
  INV_X1 U15613 ( .A(n13619), .ZN(n13620) );
  AOI21_X1 U15614 ( .B1(n13621), .B2(n13618), .A(n13620), .ZN(n13628) );
  INV_X1 U15615 ( .A(n13969), .ZN(n13625) );
  OAI22_X1 U15616 ( .A1(n13623), .A2(n14542), .B1(n13622), .B2(n14562), .ZN(
        n14120) );
  AOI22_X1 U15617 ( .A1(n14120), .A2(n14414), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13624) );
  OAI21_X1 U15618 ( .B1(n13625), .B2(n14436), .A(n13624), .ZN(n13626) );
  AOI21_X1 U15619 ( .B1(n14121), .B2(n14432), .A(n13626), .ZN(n13627) );
  OAI21_X1 U15620 ( .B1(n13628), .B2(n14426), .A(n13627), .ZN(P1_U3223) );
  XOR2_X1 U15621 ( .A(n13630), .B(n13629), .Z(n13636) );
  NAND2_X1 U15622 ( .A1(n13741), .A2(n14033), .ZN(n13632) );
  NAND2_X1 U15623 ( .A1(n13871), .A2(n14055), .ZN(n13631) );
  NAND2_X1 U15624 ( .A1(n13632), .A2(n13631), .ZN(n14094) );
  AOI22_X1 U15625 ( .A1(n14414), .A2(n14094), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13633) );
  OAI21_X1 U15626 ( .B1(n14436), .B2(n13904), .A(n13633), .ZN(n13634) );
  AOI21_X1 U15627 ( .B1(n14095), .B2(n14432), .A(n13634), .ZN(n13635) );
  OAI21_X1 U15628 ( .B1(n13636), .B2(n14426), .A(n13635), .ZN(P1_U3225) );
  INV_X1 U15629 ( .A(n13638), .ZN(n13639) );
  AOI21_X1 U15630 ( .B1(n13640), .B2(n13637), .A(n13639), .ZN(n13648) );
  NAND2_X1 U15631 ( .A1(n14414), .A2(n13641), .ZN(n13642) );
  OAI211_X1 U15632 ( .C1(n14436), .C2(n13644), .A(n13643), .B(n13642), .ZN(
        n13645) );
  AOI21_X1 U15633 ( .B1(n13646), .B2(n14432), .A(n13645), .ZN(n13647) );
  OAI21_X1 U15634 ( .B1(n13648), .B2(n14426), .A(n13647), .ZN(P1_U3226) );
  INV_X1 U15635 ( .A(n14147), .ZN(n13659) );
  OAI21_X1 U15636 ( .B1(n13651), .B2(n13649), .A(n13650), .ZN(n13652) );
  NAND2_X1 U15637 ( .A1(n13652), .A2(n14412), .ZN(n13658) );
  NOR2_X1 U15638 ( .A1(n14436), .A2(n14040), .ZN(n13656) );
  OAI21_X1 U15639 ( .B1(n14422), .B2(n13654), .A(n13653), .ZN(n13655) );
  AOI211_X1 U15640 ( .C1(n13685), .C2(n14032), .A(n13656), .B(n13655), .ZN(
        n13657) );
  OAI211_X1 U15641 ( .C1(n13659), .C2(n13737), .A(n13658), .B(n13657), .ZN(
        P1_U3228) );
  XOR2_X1 U15642 ( .A(n13661), .B(n13660), .Z(n13666) );
  AOI22_X1 U15643 ( .A1(n13685), .A2(n13954), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13663) );
  NAND2_X1 U15644 ( .A1(n13729), .A2(n13920), .ZN(n13662) );
  OAI211_X1 U15645 ( .C1(n14436), .C2(n13927), .A(n13663), .B(n13662), .ZN(
        n13664) );
  AOI21_X1 U15646 ( .B1(n14102), .B2(n14432), .A(n13664), .ZN(n13665) );
  OAI21_X1 U15647 ( .B1(n13666), .B2(n14426), .A(n13665), .ZN(P1_U3229) );
  OAI211_X1 U15648 ( .C1(n13669), .C2(n13668), .A(n13667), .B(n14412), .ZN(
        n13676) );
  INV_X1 U15649 ( .A(n13987), .ZN(n13674) );
  AND2_X1 U15650 ( .A1(n14021), .A2(n14033), .ZN(n13670) );
  AOI21_X1 U15651 ( .B1(n13953), .B2(n14055), .A(n13670), .ZN(n14127) );
  OAI22_X1 U15652 ( .A1(n14127), .A2(n13672), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13671), .ZN(n13673) );
  AOI21_X1 U15653 ( .B1(n13674), .B2(n13733), .A(n13673), .ZN(n13675) );
  OAI211_X1 U15654 ( .C1(n13677), .C2(n13737), .A(n13676), .B(n13675), .ZN(
        P1_U3233) );
  OAI211_X1 U15655 ( .C1(n13680), .C2(n13679), .A(n13678), .B(n14412), .ZN(
        n13687) );
  NOR2_X1 U15656 ( .A1(n14436), .A2(n13681), .ZN(n13684) );
  OAI21_X1 U15657 ( .B1(n14422), .B2(n13731), .A(n13682), .ZN(n13683) );
  AOI211_X1 U15658 ( .C1(n13685), .C2(n13745), .A(n13684), .B(n13683), .ZN(
        n13686) );
  OAI211_X1 U15659 ( .C1(n14443), .C2(n13737), .A(n13687), .B(n13686), .ZN(
        P1_U3234) );
  OAI21_X1 U15660 ( .B1(n13690), .B2(n13689), .A(n13688), .ZN(n13691) );
  NAND2_X1 U15661 ( .A1(n13691), .A2(n14412), .ZN(n13697) );
  INV_X1 U15662 ( .A(n13692), .ZN(n13960) );
  AOI22_X1 U15663 ( .A1(n13729), .A2(n13954), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13693) );
  OAI21_X1 U15664 ( .B1(n13694), .B2(n14419), .A(n13693), .ZN(n13695) );
  AOI21_X1 U15665 ( .B1(n13960), .B2(n13733), .A(n13695), .ZN(n13696) );
  OAI211_X1 U15666 ( .C1(n13737), .C2(n13963), .A(n13697), .B(n13696), .ZN(
        P1_U3235) );
  XOR2_X1 U15667 ( .A(n13698), .B(n13699), .Z(n13705) );
  NAND2_X1 U15668 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14523)
         );
  OAI21_X1 U15669 ( .B1(n14419), .B2(n13700), .A(n14523), .ZN(n13701) );
  AOI21_X1 U15670 ( .B1(n13729), .B2(n14021), .A(n13701), .ZN(n13702) );
  OAI21_X1 U15671 ( .B1(n14017), .B2(n14436), .A(n13702), .ZN(n13703) );
  AOI21_X1 U15672 ( .B1(n14141), .B2(n14432), .A(n13703), .ZN(n13704) );
  OAI21_X1 U15673 ( .B1(n13705), .B2(n14426), .A(n13704), .ZN(P1_U3238) );
  OAI211_X1 U15674 ( .C1(n13708), .C2(n13707), .A(n13706), .B(n14412), .ZN(
        n13717) );
  NAND2_X1 U15675 ( .A1(n13729), .A2(n13750), .ZN(n13710) );
  OAI211_X1 U15676 ( .C1(n13711), .C2(n14419), .A(n13710), .B(n13709), .ZN(
        n13712) );
  INV_X1 U15677 ( .A(n13712), .ZN(n13716) );
  NAND2_X1 U15678 ( .A1(n14432), .A2(n14607), .ZN(n13715) );
  OR2_X1 U15679 ( .A1(n14436), .A2(n13713), .ZN(n13714) );
  NAND4_X1 U15680 ( .A1(n13717), .A2(n13716), .A3(n13715), .A4(n13714), .ZN(
        P1_U3239) );
  XOR2_X1 U15681 ( .A(n13719), .B(n13718), .Z(n13725) );
  OAI22_X1 U15682 ( .A1(n13721), .A2(n14562), .B1(n13720), .B2(n14542), .ZN(
        n13887) );
  AOI22_X1 U15683 ( .A1(n14414), .A2(n13887), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13722) );
  OAI21_X1 U15684 ( .B1(n14436), .B2(n13889), .A(n13722), .ZN(n13723) );
  AOI21_X1 U15685 ( .B1(n14089), .B2(n14432), .A(n13723), .ZN(n13724) );
  OAI21_X1 U15686 ( .B1(n13725), .B2(n14426), .A(n13724), .ZN(P1_U3240) );
  OAI211_X1 U15687 ( .C1(n13728), .C2(n13727), .A(n13726), .B(n14412), .ZN(
        n13736) );
  NAND2_X1 U15688 ( .A1(n13729), .A2(n14032), .ZN(n13730) );
  NAND2_X1 U15689 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14509)
         );
  OAI211_X1 U15690 ( .C1(n13731), .C2(n14419), .A(n13730), .B(n14509), .ZN(
        n13732) );
  AOI21_X1 U15691 ( .B1(n13734), .B2(n13733), .A(n13732), .ZN(n13735) );
  OAI211_X1 U15692 ( .C1(n14439), .C2(n13737), .A(n13736), .B(n13735), .ZN(
        P1_U3241) );
  MUX2_X1 U15693 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13836), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15694 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13857), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15695 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13739), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15696 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13872), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15697 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13740), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15698 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13871), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15699 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13920), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15700 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13741), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15701 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13954), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15702 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13742), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15703 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13953), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15704 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13998), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15705 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14021), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15706 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14034), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15707 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14013), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15708 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14032), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15709 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13743), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15710 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13744), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15711 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13745), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15712 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13746), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15713 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13747), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15714 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13748), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15715 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13749), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U15716 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13750), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15717 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13751), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15718 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13752), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15719 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13753), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15720 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13754), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15721 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14054), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15722 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13755), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15723 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14049), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U15724 ( .C1(n13766), .C2(n13757), .A(n14483), .B(n13756), .ZN(
        n13765) );
  MUX2_X1 U15725 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9766), .S(n13761), .Z(
        n13758) );
  OAI21_X1 U15726 ( .B1(n9738), .B2(n13769), .A(n13758), .ZN(n13759) );
  NAND3_X1 U15727 ( .A1(n14490), .A2(n13760), .A3(n13759), .ZN(n13764) );
  NAND2_X1 U15728 ( .A1(n14492), .A2(n7237), .ZN(n13763) );
  AOI22_X1 U15729 ( .A1(n14494), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13762) );
  NAND4_X1 U15730 ( .A1(n13765), .A2(n13764), .A3(n13763), .A4(n13762), .ZN(
        P1_U3244) );
  INV_X1 U15731 ( .A(n13766), .ZN(n13768) );
  MUX2_X1 U15732 ( .A(n13768), .B(n13767), .S(n9666), .Z(n13772) );
  NAND2_X1 U15733 ( .A1(n13770), .A2(n13769), .ZN(n13771) );
  OAI211_X1 U15734 ( .C1(n13772), .C2(n9665), .A(P1_U4016), .B(n13771), .ZN(
        n14499) );
  AOI22_X1 U15735 ( .A1(n14494), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13782) );
  OAI211_X1 U15736 ( .C1(n13774), .C2(n13773), .A(n14483), .B(n13790), .ZN(
        n13777) );
  NAND2_X1 U15737 ( .A1(n14492), .A2(n13775), .ZN(n13776) );
  AND2_X1 U15738 ( .A1(n13777), .A2(n13776), .ZN(n13781) );
  OAI211_X1 U15739 ( .C1(n13779), .C2(n13778), .A(n14490), .B(n13785), .ZN(
        n13780) );
  NAND4_X1 U15740 ( .A1(n14499), .A2(n13782), .A3(n13781), .A4(n13780), .ZN(
        P1_U3245) );
  OAI22_X1 U15741 ( .A1(n14525), .A2(n14198), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14551), .ZN(n13783) );
  AOI21_X1 U15742 ( .B1(n13788), .B2(n14492), .A(n13783), .ZN(n13795) );
  MUX2_X1 U15743 ( .A(n9770), .B(P1_REG1_REG_3__SCAN_IN), .S(n13788), .Z(
        n13786) );
  NAND3_X1 U15744 ( .A1(n13786), .A2(n13785), .A3(n13784), .ZN(n13787) );
  NAND3_X1 U15745 ( .A1(n14490), .A2(n14487), .A3(n13787), .ZN(n13794) );
  MUX2_X1 U15746 ( .A(n9780), .B(P1_REG2_REG_3__SCAN_IN), .S(n13788), .Z(
        n13791) );
  NAND3_X1 U15747 ( .A1(n13791), .A2(n13790), .A3(n13789), .ZN(n13792) );
  NAND3_X1 U15748 ( .A1(n14483), .A2(n14480), .A3(n13792), .ZN(n13793) );
  NAND3_X1 U15749 ( .A1(n13795), .A2(n13794), .A3(n13793), .ZN(P1_U3246) );
  INV_X1 U15750 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14205) );
  OAI21_X1 U15751 ( .B1(n14525), .B2(n14205), .A(n13796), .ZN(n13797) );
  AOI21_X1 U15752 ( .B1(n13798), .B2(n14492), .A(n13797), .ZN(n13810) );
  OAI21_X1 U15753 ( .B1(n13801), .B2(n13800), .A(n13799), .ZN(n13802) );
  NAND2_X1 U15754 ( .A1(n14490), .A2(n13802), .ZN(n13809) );
  INV_X1 U15755 ( .A(n13803), .ZN(n13807) );
  NAND3_X1 U15756 ( .A1(n14482), .A2(n13805), .A3(n13804), .ZN(n13806) );
  NAND3_X1 U15757 ( .A1(n14483), .A2(n13807), .A3(n13806), .ZN(n13808) );
  NAND3_X1 U15758 ( .A1(n13810), .A2(n13809), .A3(n13808), .ZN(P1_U3248) );
  OAI21_X1 U15759 ( .B1(n13812), .B2(n13817), .A(n13811), .ZN(n13813) );
  XNOR2_X1 U15760 ( .A(n14520), .B(n13813), .ZN(n14515) );
  NAND2_X1 U15761 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n14515), .ZN(n14514) );
  NAND2_X1 U15762 ( .A1(n13819), .A2(n13813), .ZN(n13814) );
  NAND2_X1 U15763 ( .A1(n14514), .A2(n13814), .ZN(n13815) );
  XOR2_X1 U15764 ( .A(n13815), .B(P1_REG1_REG_19__SCAN_IN), .Z(n13823) );
  OAI21_X1 U15765 ( .B1(n14041), .B2(n13817), .A(n13816), .ZN(n13818) );
  NAND2_X1 U15766 ( .A1(n13819), .A2(n13818), .ZN(n13820) );
  XOR2_X1 U15767 ( .A(n13819), .B(n13818), .Z(n14513) );
  NAND2_X1 U15768 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14513), .ZN(n14512) );
  NAND2_X1 U15769 ( .A1(n13820), .A2(n14512), .ZN(n13821) );
  XOR2_X1 U15770 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13821), .Z(n13822) );
  AOI22_X1 U15771 ( .A1(n13823), .A2(n14490), .B1(n14483), .B2(n13822), .ZN(
        n13828) );
  INV_X1 U15772 ( .A(n13822), .ZN(n13825) );
  NOR2_X1 U15773 ( .A1(n13823), .A2(n14517), .ZN(n13824) );
  AOI211_X1 U15774 ( .C1(n14483), .C2(n13825), .A(n14492), .B(n13824), .ZN(
        n13827) );
  MUX2_X1 U15775 ( .A(n13828), .B(n13827), .S(n13826), .Z(n13830) );
  OAI211_X1 U15776 ( .C1(n7462), .C2(n14525), .A(n13830), .B(n13829), .ZN(
        P1_U3262) );
  NAND2_X1 U15777 ( .A1(n13855), .A2(n13854), .ZN(n13853) );
  NOR2_X1 U15778 ( .A1(n13842), .A2(n13853), .ZN(n13831) );
  XNOR2_X1 U15779 ( .A(n13831), .B(n13838), .ZN(n13832) );
  NAND2_X1 U15780 ( .A1(n13832), .A2(n14556), .ZN(n14064) );
  NOR2_X1 U15781 ( .A1(n14576), .A2(n13833), .ZN(n13837) );
  INV_X1 U15782 ( .A(P1_B_REG_SCAN_IN), .ZN(n13834) );
  NOR2_X1 U15783 ( .A1(n9666), .A2(n13834), .ZN(n13835) );
  NOR2_X1 U15784 ( .A1(n14562), .A2(n13835), .ZN(n13856) );
  NAND2_X1 U15785 ( .A1(n13836), .A2(n13856), .ZN(n14066) );
  NOR2_X1 U15786 ( .A1(n14578), .A2(n14066), .ZN(n13841) );
  AOI211_X1 U15787 ( .C1(n13838), .C2(n14550), .A(n13837), .B(n13841), .ZN(
        n13839) );
  OAI21_X1 U15788 ( .B1(n14064), .B2(n13947), .A(n13839), .ZN(P1_U3263) );
  XNOR2_X1 U15789 ( .A(n14068), .B(n13853), .ZN(n13840) );
  NAND2_X1 U15790 ( .A1(n13840), .A2(n14556), .ZN(n14067) );
  AOI21_X1 U15791 ( .B1(n14578), .B2(P1_REG2_REG_30__SCAN_IN), .A(n13841), 
        .ZN(n13844) );
  NAND2_X1 U15792 ( .A1(n13842), .A2(n14550), .ZN(n13843) );
  OAI211_X1 U15793 ( .C1(n14067), .C2(n13947), .A(n13844), .B(n13843), .ZN(
        P1_U3264) );
  NAND2_X1 U15794 ( .A1(n14079), .A2(n13872), .ZN(n13849) );
  NAND2_X1 U15795 ( .A1(n13850), .A2(n13849), .ZN(n13852) );
  XNOR2_X1 U15796 ( .A(n13852), .B(n13851), .ZN(n14069) );
  OAI211_X1 U15797 ( .C1(n13855), .C2(n13854), .A(n14556), .B(n13853), .ZN(
        n14073) );
  INV_X1 U15798 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n13864) );
  AND2_X1 U15799 ( .A1(n13857), .A2(n13856), .ZN(n14070) );
  INV_X1 U15800 ( .A(n14070), .ZN(n13859) );
  NOR2_X1 U15801 ( .A1(n13859), .A2(n13858), .ZN(n13861) );
  AOI22_X1 U15802 ( .A1(n13862), .A2(n13861), .B1(n13860), .B2(n14574), .ZN(
        n13863) );
  OAI21_X1 U15803 ( .B1(n14576), .B2(n13864), .A(n13863), .ZN(n13865) );
  AOI21_X1 U15804 ( .B1(n14071), .B2(n14550), .A(n13865), .ZN(n13866) );
  OAI21_X1 U15805 ( .B1(n14073), .B2(n13947), .A(n13866), .ZN(n13867) );
  AOI21_X1 U15806 ( .B1(n14069), .B2(n14571), .A(n13867), .ZN(n13868) );
  OAI21_X1 U15807 ( .B1(n14075), .B2(n14578), .A(n13868), .ZN(P1_U3356) );
  XNOR2_X1 U15808 ( .A(n13869), .B(n7218), .ZN(n14087) );
  INV_X1 U15809 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n13874) );
  OAI22_X1 U15810 ( .A1(n14576), .A2(n13874), .B1(n13873), .B2(n14526), .ZN(
        n13875) );
  AOI21_X1 U15811 ( .B1(n14084), .B2(n14550), .A(n13875), .ZN(n13879) );
  AOI21_X1 U15812 ( .B1(n14084), .B2(n13894), .A(n14058), .ZN(n13877) );
  NAND2_X1 U15813 ( .A1(n14083), .A2(n14558), .ZN(n13878) );
  OAI211_X1 U15814 ( .C1(n14086), .C2(n14578), .A(n13879), .B(n13878), .ZN(
        n13880) );
  INV_X1 U15815 ( .A(n13880), .ZN(n13881) );
  OAI21_X1 U15816 ( .B1(n14087), .B2(n14536), .A(n13881), .ZN(P1_U3266) );
  XNOR2_X1 U15817 ( .A(n13882), .B(n13883), .ZN(n14092) );
  OAI21_X1 U15818 ( .B1(n13886), .B2(n13885), .A(n13884), .ZN(n13888) );
  AOI21_X1 U15819 ( .B1(n13888), .B2(n14549), .A(n13887), .ZN(n14091) );
  OAI22_X1 U15820 ( .A1(n14576), .A2(n13890), .B1(n13889), .B2(n14526), .ZN(
        n13891) );
  AOI21_X1 U15821 ( .B1(n14089), .B2(n14550), .A(n13891), .ZN(n13896) );
  OR2_X1 U15822 ( .A1(n13892), .A2(n6524), .ZN(n13893) );
  AND3_X1 U15823 ( .A1(n13894), .A2(n13893), .A3(n14556), .ZN(n14088) );
  NAND2_X1 U15824 ( .A1(n14088), .A2(n14558), .ZN(n13895) );
  OAI211_X1 U15825 ( .C1(n14091), .C2(n14578), .A(n13896), .B(n13895), .ZN(
        n13897) );
  INV_X1 U15826 ( .A(n13897), .ZN(n13898) );
  OAI21_X1 U15827 ( .B1(n14092), .B2(n14536), .A(n13898), .ZN(P1_U3267) );
  OAI21_X1 U15828 ( .B1(n13900), .B2(n13910), .A(n13899), .ZN(n14099) );
  NAND2_X1 U15829 ( .A1(n14095), .A2(n13924), .ZN(n13901) );
  NAND2_X1 U15830 ( .A1(n13901), .A2(n14556), .ZN(n13902) );
  NOR2_X1 U15831 ( .A1(n6524), .A2(n13902), .ZN(n14093) );
  INV_X1 U15832 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n13908) );
  NAND2_X1 U15833 ( .A1(n14095), .A2(n14550), .ZN(n13907) );
  INV_X1 U15834 ( .A(n14094), .ZN(n13903) );
  OAI21_X1 U15835 ( .B1(n13904), .B2(n14526), .A(n13903), .ZN(n13905) );
  NAND2_X1 U15836 ( .A1(n14576), .A2(n13905), .ZN(n13906) );
  OAI211_X1 U15837 ( .C1(n14576), .C2(n13908), .A(n13907), .B(n13906), .ZN(
        n13909) );
  AOI21_X1 U15838 ( .B1(n14093), .B2(n14558), .A(n13909), .ZN(n13913) );
  XNOR2_X1 U15839 ( .A(n13911), .B(n13910), .ZN(n14096) );
  NAND2_X1 U15840 ( .A1(n14096), .A2(n14570), .ZN(n13912) );
  OAI211_X1 U15841 ( .C1(n14099), .C2(n14536), .A(n13913), .B(n13912), .ZN(
        P1_U3268) );
  OAI21_X1 U15842 ( .B1(n13916), .B2(n13915), .A(n13914), .ZN(n14100) );
  OAI211_X1 U15843 ( .C1(n13919), .C2(n13918), .A(n13917), .B(n14549), .ZN(
        n13922) );
  AOI22_X1 U15844 ( .A1(n14033), .A2(n13954), .B1(n13920), .B2(n14055), .ZN(
        n13921) );
  NAND2_X1 U15845 ( .A1(n13922), .A2(n13921), .ZN(n13923) );
  AOI21_X1 U15846 ( .B1(n14100), .B2(n14593), .A(n13923), .ZN(n14104) );
  INV_X1 U15847 ( .A(n13924), .ZN(n13925) );
  AOI211_X1 U15848 ( .C1(n14102), .C2(n13941), .A(n14058), .B(n13925), .ZN(
        n14101) );
  INV_X1 U15849 ( .A(n14102), .ZN(n13926) );
  NOR2_X1 U15850 ( .A1(n13926), .A2(n14530), .ZN(n13930) );
  OAI22_X1 U15851 ( .A1(n14576), .A2(n13928), .B1(n13927), .B2(n14526), .ZN(
        n13929) );
  AOI211_X1 U15852 ( .C1(n14101), .C2(n14558), .A(n13930), .B(n13929), .ZN(
        n13932) );
  NAND2_X1 U15853 ( .A1(n14100), .A2(n14559), .ZN(n13931) );
  OAI211_X1 U15854 ( .C1(n14104), .C2(n14578), .A(n13932), .B(n13931), .ZN(
        P1_U3269) );
  AOI21_X1 U15855 ( .B1(n13935), .B2(n13934), .A(n13933), .ZN(n14106) );
  AND2_X1 U15856 ( .A1(n13937), .A2(n13936), .ZN(n13938) );
  OAI21_X1 U15857 ( .B1(n13939), .B2(n13938), .A(n14549), .ZN(n14110) );
  INV_X1 U15858 ( .A(n14107), .ZN(n13940) );
  AOI21_X1 U15859 ( .B1(n14110), .B2(n13940), .A(n14578), .ZN(n13949) );
  OAI211_X1 U15860 ( .C1(n13958), .C2(n13942), .A(n14556), .B(n13941), .ZN(
        n14109) );
  INV_X1 U15861 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n13944) );
  OAI22_X1 U15862 ( .A1(n14576), .A2(n13944), .B1(n13943), .B2(n14526), .ZN(
        n13945) );
  AOI21_X1 U15863 ( .B1(n14108), .B2(n14550), .A(n13945), .ZN(n13946) );
  OAI21_X1 U15864 ( .B1(n14109), .B2(n13947), .A(n13946), .ZN(n13948) );
  AOI211_X1 U15865 ( .C1(n14106), .C2(n14571), .A(n13949), .B(n13948), .ZN(
        n13950) );
  INV_X1 U15866 ( .A(n13950), .ZN(P1_U3270) );
  XNOR2_X1 U15867 ( .A(n13952), .B(n13951), .ZN(n13955) );
  AOI222_X1 U15868 ( .A1(n14549), .A2(n13955), .B1(n13954), .B2(n14055), .C1(
        n13953), .C2(n14033), .ZN(n14117) );
  OAI21_X1 U15869 ( .B1(n13957), .B2(n7199), .A(n13956), .ZN(n14113) );
  INV_X1 U15870 ( .A(n13967), .ZN(n13959) );
  AOI211_X1 U15871 ( .C1(n14115), .C2(n13959), .A(n14058), .B(n13958), .ZN(
        n14114) );
  NAND2_X1 U15872 ( .A1(n14114), .A2(n14558), .ZN(n13962) );
  AOI22_X1 U15873 ( .A1(n14578), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n13960), 
        .B2(n14574), .ZN(n13961) );
  OAI211_X1 U15874 ( .C1(n14530), .C2(n13963), .A(n13962), .B(n13961), .ZN(
        n13964) );
  AOI21_X1 U15875 ( .B1(n14113), .B2(n14571), .A(n13964), .ZN(n13965) );
  OAI21_X1 U15876 ( .B1(n14578), .B2(n14117), .A(n13965), .ZN(P1_U3271) );
  XNOR2_X1 U15877 ( .A(n13966), .B(n13975), .ZN(n14125) );
  OAI21_X1 U15878 ( .B1(n13986), .B2(n13973), .A(n14556), .ZN(n13968) );
  NOR2_X1 U15879 ( .A1(n13968), .A2(n13967), .ZN(n14119) );
  AOI21_X1 U15880 ( .B1(n13969), .B2(n14574), .A(n14120), .ZN(n13970) );
  NOR2_X1 U15881 ( .A1(n13970), .A2(n14578), .ZN(n13971) );
  AOI21_X1 U15882 ( .B1(n14578), .B2(P1_REG2_REG_21__SCAN_IN), .A(n13971), 
        .ZN(n13972) );
  OAI21_X1 U15883 ( .B1(n13973), .B2(n14530), .A(n13972), .ZN(n13974) );
  AOI21_X1 U15884 ( .B1(n14119), .B2(n14558), .A(n13974), .ZN(n13978) );
  XNOR2_X1 U15885 ( .A(n13976), .B(n13975), .ZN(n14122) );
  NAND2_X1 U15886 ( .A1(n14122), .A2(n14570), .ZN(n13977) );
  OAI211_X1 U15887 ( .C1(n14125), .C2(n14536), .A(n13978), .B(n13977), .ZN(
        P1_U3272) );
  OAI21_X1 U15888 ( .B1(n13981), .B2(n13980), .A(n13979), .ZN(n14133) );
  XNOR2_X1 U15889 ( .A(n13983), .B(n13982), .ZN(n14126) );
  NAND2_X1 U15890 ( .A1(n14126), .A2(n14571), .ZN(n13994) );
  NAND2_X1 U15891 ( .A1(n14002), .A2(n14130), .ZN(n13984) );
  NAND2_X1 U15892 ( .A1(n13984), .A2(n14556), .ZN(n13985) );
  NOR2_X1 U15893 ( .A1(n13986), .A2(n13985), .ZN(n14128) );
  INV_X1 U15894 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n13991) );
  NAND2_X1 U15895 ( .A1(n14130), .A2(n14550), .ZN(n13990) );
  OAI22_X1 U15896 ( .A1(n14127), .A2(n14578), .B1(n13987), .B2(n14526), .ZN(
        n13988) );
  INV_X1 U15897 ( .A(n13988), .ZN(n13989) );
  OAI211_X1 U15898 ( .C1(n14576), .C2(n13991), .A(n13990), .B(n13989), .ZN(
        n13992) );
  AOI21_X1 U15899 ( .B1(n14128), .B2(n14558), .A(n13992), .ZN(n13993) );
  OAI211_X1 U15900 ( .C1(n14133), .C2(n13995), .A(n13994), .B(n13993), .ZN(
        P1_U3273) );
  XNOR2_X1 U15901 ( .A(n13997), .B(n13996), .ZN(n13999) );
  AOI222_X1 U15902 ( .A1(n14549), .A2(n13999), .B1(n13998), .B2(n14055), .C1(
        n14034), .C2(n14033), .ZN(n14138) );
  OAI21_X1 U15903 ( .B1(n14001), .B2(n7168), .A(n14000), .ZN(n14134) );
  AOI211_X1 U15904 ( .C1(n14136), .C2(n14003), .A(n14058), .B(n6939), .ZN(
        n14135) );
  NAND2_X1 U15905 ( .A1(n14135), .A2(n14558), .ZN(n14007) );
  INV_X1 U15906 ( .A(n14004), .ZN(n14005) );
  AOI22_X1 U15907 ( .A1(n14578), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14005), 
        .B2(n14574), .ZN(n14006) );
  OAI211_X1 U15908 ( .C1(n14008), .C2(n14530), .A(n14007), .B(n14006), .ZN(
        n14009) );
  AOI21_X1 U15909 ( .B1(n14134), .B2(n14571), .A(n14009), .ZN(n14010) );
  OAI21_X1 U15910 ( .B1(n14578), .B2(n14138), .A(n14010), .ZN(P1_U3274) );
  XNOR2_X1 U15911 ( .A(n14012), .B(n14011), .ZN(n14014) );
  AOI22_X1 U15912 ( .A1(n14014), .A2(n14549), .B1(n14033), .B2(n14013), .ZN(
        n14143) );
  XNOR2_X1 U15913 ( .A(n14016), .B(n14015), .ZN(n14144) );
  OAI22_X1 U15914 ( .A1(n14576), .A2(n14018), .B1(n14017), .B2(n14526), .ZN(
        n14019) );
  AOI21_X1 U15915 ( .B1(n14141), .B2(n14550), .A(n14019), .ZN(n14025) );
  XNOR2_X1 U15916 ( .A(n14141), .B(n6940), .ZN(n14020) );
  NAND2_X1 U15917 ( .A1(n14020), .A2(n14556), .ZN(n14023) );
  NAND2_X1 U15918 ( .A1(n14021), .A2(n14055), .ZN(n14022) );
  NAND2_X1 U15919 ( .A1(n14023), .A2(n14022), .ZN(n14140) );
  NAND2_X1 U15920 ( .A1(n14140), .A2(n14558), .ZN(n14024) );
  OAI211_X1 U15921 ( .C1(n14144), .C2(n14536), .A(n14025), .B(n14024), .ZN(
        n14026) );
  INV_X1 U15922 ( .A(n14026), .ZN(n14027) );
  OAI21_X1 U15923 ( .B1(n14578), .B2(n14143), .A(n14027), .ZN(P1_U3275) );
  XNOR2_X1 U15924 ( .A(n14029), .B(n14028), .ZN(n14149) );
  OAI211_X1 U15925 ( .C1(n6517), .C2(n14031), .A(n14030), .B(n14549), .ZN(
        n14036) );
  AOI22_X1 U15926 ( .A1(n14034), .A2(n14055), .B1(n14033), .B2(n14032), .ZN(
        n14035) );
  NAND2_X1 U15927 ( .A1(n14036), .A2(n14035), .ZN(n14145) );
  AOI21_X1 U15928 ( .B1(n14147), .B2(n14037), .A(n14058), .ZN(n14039) );
  AND2_X1 U15929 ( .A1(n14039), .A2(n14038), .ZN(n14146) );
  NAND2_X1 U15930 ( .A1(n14146), .A2(n14558), .ZN(n14044) );
  OAI22_X1 U15931 ( .A1(n14576), .A2(n14041), .B1(n14040), .B2(n14526), .ZN(
        n14042) );
  AOI21_X1 U15932 ( .B1(n14147), .B2(n14550), .A(n14042), .ZN(n14043) );
  NAND2_X1 U15933 ( .A1(n14044), .A2(n14043), .ZN(n14045) );
  AOI21_X1 U15934 ( .B1(n14145), .B2(n14576), .A(n14045), .ZN(n14046) );
  OAI21_X1 U15935 ( .B1(n14149), .B2(n14536), .A(n14046), .ZN(P1_U3276) );
  OAI21_X1 U15936 ( .B1(n10219), .B2(n14047), .A(n14549), .ZN(n14052) );
  AOI21_X1 U15937 ( .B1(n14565), .B2(n14586), .A(n6491), .ZN(n14057) );
  XNOR2_X1 U15938 ( .A(n14057), .B(n14563), .ZN(n14050) );
  AOI21_X1 U15939 ( .B1(n14050), .B2(n14549), .A(n14049), .ZN(n14051) );
  AOI21_X1 U15940 ( .B1(n14542), .B2(n14052), .A(n14051), .ZN(n14053) );
  AOI21_X1 U15941 ( .B1(n14055), .B2(n14054), .A(n14053), .ZN(n14589) );
  MUX2_X1 U15942 ( .A(n14056), .B(n14589), .S(n14576), .Z(n14063) );
  AOI22_X1 U15943 ( .A1(n14550), .A2(n14586), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n14574), .ZN(n14062) );
  INV_X1 U15944 ( .A(n14057), .ZN(n14059) );
  NOR2_X1 U15945 ( .A1(n14059), .A2(n14058), .ZN(n14585) );
  XNOR2_X1 U15946 ( .A(n10219), .B(n14060), .ZN(n14592) );
  AOI22_X1 U15947 ( .A1(n14558), .A2(n14585), .B1(n14571), .B2(n14592), .ZN(
        n14061) );
  NAND3_X1 U15948 ( .A1(n14063), .A2(n14062), .A3(n14061), .ZN(P1_U3292) );
  OAI211_X1 U15949 ( .C1(n14065), .C2(n14640), .A(n14064), .B(n14066), .ZN(
        n14157) );
  MUX2_X1 U15950 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14157), .S(n14657), .Z(
        P1_U3559) );
  OAI211_X1 U15951 ( .C1(n14068), .C2(n14640), .A(n14067), .B(n14066), .ZN(
        n14158) );
  MUX2_X1 U15952 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14158), .S(n14657), .Z(
        P1_U3558) );
  NAND2_X1 U15953 ( .A1(n14069), .A2(n14644), .ZN(n14076) );
  AOI21_X1 U15954 ( .B1(n14071), .B2(n14606), .A(n14070), .ZN(n14072) );
  NAND2_X1 U15955 ( .A1(n14076), .A2(n7429), .ZN(n14159) );
  MUX2_X1 U15956 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14159), .S(n14657), .Z(
        P1_U3557) );
  INV_X1 U15957 ( .A(n14077), .ZN(n14078) );
  AOI21_X1 U15958 ( .B1(n14079), .B2(n14606), .A(n14078), .ZN(n14080) );
  OAI211_X1 U15959 ( .C1(n14082), .C2(n14581), .A(n14081), .B(n14080), .ZN(
        n14160) );
  MUX2_X1 U15960 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14160), .S(n14657), .Z(
        P1_U3556) );
  AOI21_X1 U15961 ( .B1(n14084), .B2(n14606), .A(n14083), .ZN(n14085) );
  OAI211_X1 U15962 ( .C1(n14087), .C2(n14581), .A(n14086), .B(n14085), .ZN(
        n14161) );
  MUX2_X1 U15963 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14161), .S(n14657), .Z(
        P1_U3555) );
  AOI21_X1 U15964 ( .B1(n14089), .B2(n14606), .A(n14088), .ZN(n14090) );
  OAI211_X1 U15965 ( .C1(n14092), .C2(n14581), .A(n14091), .B(n14090), .ZN(
        n14162) );
  MUX2_X1 U15966 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14162), .S(n14657), .Z(
        P1_U3554) );
  AOI211_X1 U15967 ( .C1(n14095), .C2(n14606), .A(n14094), .B(n14093), .ZN(
        n14098) );
  NAND2_X1 U15968 ( .A1(n14096), .A2(n14549), .ZN(n14097) );
  OAI211_X1 U15969 ( .C1(n14099), .C2(n14581), .A(n14098), .B(n14097), .ZN(
        n14163) );
  MUX2_X1 U15970 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14163), .S(n14657), .Z(
        P1_U3553) );
  INV_X1 U15971 ( .A(n14100), .ZN(n14105) );
  AOI21_X1 U15972 ( .B1(n14102), .B2(n14606), .A(n14101), .ZN(n14103) );
  OAI211_X1 U15973 ( .C1(n14105), .C2(n14609), .A(n14104), .B(n14103), .ZN(
        n14164) );
  MUX2_X1 U15974 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14164), .S(n14657), .Z(
        P1_U3552) );
  NAND2_X1 U15975 ( .A1(n14106), .A2(n14644), .ZN(n14112) );
  AOI21_X1 U15976 ( .B1(n14108), .B2(n14606), .A(n14107), .ZN(n14111) );
  NAND4_X1 U15977 ( .A1(n14112), .A2(n14111), .A3(n14110), .A4(n14109), .ZN(
        n14165) );
  MUX2_X1 U15978 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14165), .S(n14657), .Z(
        P1_U3551) );
  INV_X1 U15979 ( .A(n14113), .ZN(n14118) );
  AOI21_X1 U15980 ( .B1(n14115), .B2(n14606), .A(n14114), .ZN(n14116) );
  OAI211_X1 U15981 ( .C1(n14118), .C2(n14581), .A(n14117), .B(n14116), .ZN(
        n14166) );
  MUX2_X1 U15982 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14166), .S(n14657), .Z(
        P1_U3550) );
  AOI211_X1 U15983 ( .C1(n14121), .C2(n14606), .A(n14120), .B(n14119), .ZN(
        n14124) );
  NAND2_X1 U15984 ( .A1(n14122), .A2(n14549), .ZN(n14123) );
  OAI211_X1 U15985 ( .C1(n14125), .C2(n14581), .A(n14124), .B(n14123), .ZN(
        n14167) );
  MUX2_X1 U15986 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14167), .S(n14657), .Z(
        P1_U3549) );
  NAND2_X1 U15987 ( .A1(n14126), .A2(n14644), .ZN(n14132) );
  INV_X1 U15988 ( .A(n14127), .ZN(n14129) );
  AOI211_X1 U15989 ( .C1(n14130), .C2(n14606), .A(n14129), .B(n14128), .ZN(
        n14131) );
  OAI211_X1 U15990 ( .C1(n14580), .C2(n14133), .A(n14132), .B(n14131), .ZN(
        n14168) );
  MUX2_X1 U15991 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14168), .S(n14657), .Z(
        P1_U3548) );
  INV_X1 U15992 ( .A(n14134), .ZN(n14139) );
  AOI21_X1 U15993 ( .B1(n14136), .B2(n14606), .A(n14135), .ZN(n14137) );
  OAI211_X1 U15994 ( .C1(n14139), .C2(n14581), .A(n14138), .B(n14137), .ZN(
        n14169) );
  MUX2_X1 U15995 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14169), .S(n14657), .Z(
        P1_U3547) );
  AOI21_X1 U15996 ( .B1(n14141), .B2(n14606), .A(n14140), .ZN(n14142) );
  OAI211_X1 U15997 ( .C1(n14144), .C2(n14581), .A(n14143), .B(n14142), .ZN(
        n14170) );
  MUX2_X1 U15998 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14170), .S(n14657), .Z(
        P1_U3546) );
  AOI211_X1 U15999 ( .C1(n14147), .C2(n14606), .A(n14146), .B(n14145), .ZN(
        n14148) );
  OAI21_X1 U16000 ( .B1(n14149), .B2(n14581), .A(n14148), .ZN(n14171) );
  MUX2_X1 U16001 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14171), .S(n14657), .Z(
        P1_U3545) );
  OAI211_X1 U16002 ( .C1(n14152), .C2(n14640), .A(n14151), .B(n14150), .ZN(
        n14153) );
  AOI21_X1 U16003 ( .B1(n14154), .B2(n14549), .A(n14153), .ZN(n14155) );
  OAI21_X1 U16004 ( .B1(n14156), .B2(n14581), .A(n14155), .ZN(n14172) );
  MUX2_X1 U16005 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14172), .S(n14657), .Z(
        P1_U3544) );
  MUX2_X1 U16006 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14157), .S(n14646), .Z(
        P1_U3527) );
  MUX2_X1 U16007 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14158), .S(n14646), .Z(
        P1_U3526) );
  MUX2_X1 U16008 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14159), .S(n14646), .Z(
        P1_U3525) );
  MUX2_X1 U16009 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14160), .S(n14646), .Z(
        P1_U3524) );
  MUX2_X1 U16010 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14161), .S(n14646), .Z(
        P1_U3523) );
  MUX2_X1 U16011 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14162), .S(n14646), .Z(
        P1_U3522) );
  MUX2_X1 U16012 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14163), .S(n14646), .Z(
        P1_U3521) );
  MUX2_X1 U16013 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14164), .S(n14646), .Z(
        P1_U3520) );
  MUX2_X1 U16014 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14165), .S(n14646), .Z(
        P1_U3519) );
  MUX2_X1 U16015 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14166), .S(n14646), .Z(
        P1_U3518) );
  MUX2_X1 U16016 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14167), .S(n14646), .Z(
        P1_U3517) );
  MUX2_X1 U16017 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14168), .S(n14646), .Z(
        P1_U3516) );
  MUX2_X1 U16018 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14169), .S(n14646), .Z(
        P1_U3515) );
  MUX2_X1 U16019 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14170), .S(n14646), .Z(
        P1_U3513) );
  MUX2_X1 U16020 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14171), .S(n14646), .Z(
        P1_U3510) );
  MUX2_X1 U16021 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14172), .S(n14646), .Z(
        P1_U3507) );
  NAND3_X1 U16022 ( .A1(n14174), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n14176) );
  OAI22_X1 U16023 ( .A1(n14173), .A2(n14176), .B1(n14175), .B2(n14180), .ZN(
        n14177) );
  AOI21_X1 U16024 ( .B1(n9563), .B2(n14178), .A(n14177), .ZN(n14179) );
  INV_X1 U16025 ( .A(n14179), .ZN(P1_U3324) );
  OAI222_X1 U16026 ( .A1(P1_U3086), .A2(n9666), .B1(n14183), .B2(n14185), .C1(
        n14184), .C2(n14180), .ZN(P1_U3328) );
  OAI222_X1 U16027 ( .A1(n14188), .A2(P1_U3086), .B1(n14183), .B2(n14187), 
        .C1(n14186), .C2(n14180), .ZN(P1_U3329) );
  MUX2_X1 U16028 ( .A(n14190), .B(n14189), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U16029 ( .A(n14191), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16030 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14333) );
  NAND2_X1 U16031 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14233), .ZN(n14192) );
  OAI21_X1 U16032 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n14233), .A(n14192), 
        .ZN(n14295) );
  INV_X1 U16033 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14511) );
  NOR2_X1 U16034 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14511), .ZN(n14231) );
  INV_X1 U16035 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14193) );
  XOR2_X1 U16036 ( .A(n14193), .B(P1_ADDR_REG_14__SCAN_IN), .Z(n14238) );
  INV_X1 U16037 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14289) );
  XOR2_X1 U16038 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(n14225), .Z(n14285) );
  XNOR2_X1 U16039 ( .A(n14194), .B(n14223), .ZN(n14279) );
  XOR2_X1 U16040 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n14217), .Z(n14273) );
  INV_X1 U16041 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14215) );
  XOR2_X1 U16042 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n14215), .Z(n14268) );
  XOR2_X1 U16043 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n14209), .Z(n14261) );
  NAND2_X1 U16044 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14197), .ZN(n14200) );
  NAND2_X1 U16045 ( .A1(n14252), .A2(n14198), .ZN(n14199) );
  NAND2_X1 U16046 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14202), .ZN(n14203) );
  NAND2_X1 U16047 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14204), .ZN(n14207) );
  NAND2_X1 U16048 ( .A1(n14255), .A2(n14205), .ZN(n14206) );
  NAND2_X1 U16049 ( .A1(n14207), .A2(n14206), .ZN(n14262) );
  NAND2_X1 U16050 ( .A1(n14261), .A2(n14262), .ZN(n14208) );
  NAND2_X1 U16051 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14210), .ZN(n14213) );
  XOR2_X1 U16052 ( .A(n14210), .B(P3_ADDR_REG_7__SCAN_IN), .Z(n14265) );
  INV_X1 U16053 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14211) );
  NAND2_X1 U16054 ( .A1(n14265), .A2(n14211), .ZN(n14212) );
  NAND2_X1 U16055 ( .A1(n14213), .A2(n14212), .ZN(n14269) );
  NAND2_X1 U16056 ( .A1(n14268), .A2(n14269), .ZN(n14214) );
  NAND2_X1 U16057 ( .A1(n14273), .A2(n14274), .ZN(n14216) );
  NAND2_X1 U16058 ( .A1(n14219), .A2(n14218), .ZN(n14221) );
  XOR2_X1 U16059 ( .A(n14219), .B(n14218), .Z(n14275) );
  NAND2_X1 U16060 ( .A1(n14275), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n14220) );
  NAND2_X1 U16061 ( .A1(n14221), .A2(n14220), .ZN(n14280) );
  NAND2_X1 U16062 ( .A1(n14279), .A2(n14280), .ZN(n14222) );
  NAND2_X1 U16063 ( .A1(n14285), .A2(n14286), .ZN(n14224) );
  NAND2_X1 U16064 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14226), .ZN(n14227) );
  NAND2_X1 U16065 ( .A1(n14238), .A2(n14237), .ZN(n14228) );
  INV_X1 U16066 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14230) );
  OAI22_X1 U16067 ( .A1(n14231), .A2(n14235), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n14230), .ZN(n14296) );
  NOR2_X1 U16068 ( .A1(n14295), .A2(n14296), .ZN(n14232) );
  AOI21_X1 U16069 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n14233), .A(n14232), 
        .ZN(n14234) );
  INV_X1 U16070 ( .A(n14234), .ZN(n14300) );
  XNOR2_X1 U16071 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14300), .ZN(n14301) );
  XOR2_X1 U16072 ( .A(n14333), .B(n14301), .Z(n14323) );
  INV_X1 U16073 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14477) );
  INV_X1 U16074 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14294) );
  XOR2_X1 U16075 ( .A(n14511), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n14236) );
  XOR2_X1 U16076 ( .A(n14236), .B(n14235), .Z(n14470) );
  XOR2_X1 U16077 ( .A(n14238), .B(n14237), .Z(n14466) );
  NAND2_X1 U16078 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14241), .ZN(n14254) );
  INV_X1 U16079 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14251) );
  XNOR2_X1 U16080 ( .A(n14243), .B(n14242), .ZN(n14309) );
  XNOR2_X1 U16081 ( .A(n14244), .B(n14245), .ZN(n14247) );
  NAND2_X1 U16082 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14247), .ZN(n14249) );
  AOI21_X1 U16083 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14246), .A(n14245), .ZN(
        n15216) );
  INV_X1 U16084 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15215) );
  NOR2_X1 U16085 ( .A1(n15216), .A2(n15215), .ZN(n15225) );
  XOR2_X1 U16086 ( .A(n14247), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15224) );
  NAND2_X1 U16087 ( .A1(n15225), .A2(n15224), .ZN(n14248) );
  NAND2_X1 U16088 ( .A1(n14309), .A2(n14310), .ZN(n14250) );
  NOR2_X1 U16089 ( .A1(n14309), .A2(n14310), .ZN(n14308) );
  XOR2_X1 U16090 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14252), .Z(n15221) );
  NOR2_X1 U16091 ( .A1(n15220), .A2(n15221), .ZN(n14253) );
  INV_X1 U16092 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15222) );
  NAND2_X1 U16093 ( .A1(n15220), .A2(n15221), .ZN(n15219) );
  NOR2_X1 U16094 ( .A1(n14257), .A2(n14256), .ZN(n14259) );
  XNOR2_X1 U16095 ( .A(n14256), .B(n14257), .ZN(n15214) );
  NOR2_X1 U16096 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n15214), .ZN(n14258) );
  NAND2_X1 U16097 ( .A1(n14260), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14263) );
  XNOR2_X1 U16098 ( .A(n14262), .B(n14261), .ZN(n14312) );
  NOR2_X1 U16099 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14264), .ZN(n14267) );
  XOR2_X1 U16100 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14265), .Z(n15217) );
  NOR2_X1 U16101 ( .A1(n15218), .A2(n15217), .ZN(n14266) );
  XNOR2_X1 U16102 ( .A(n14269), .B(n14268), .ZN(n14271) );
  NAND2_X1 U16103 ( .A1(n14270), .A2(n14271), .ZN(n14272) );
  XNOR2_X1 U16104 ( .A(n14274), .B(n14273), .ZN(n14316) );
  INV_X1 U16105 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14734) );
  NAND2_X1 U16106 ( .A1(n14317), .A2(n14316), .ZN(n14315) );
  INV_X1 U16107 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14974) );
  XOR2_X1 U16108 ( .A(n14275), .B(n14974), .Z(n14276) );
  NOR2_X1 U16109 ( .A1(n14277), .A2(n14276), .ZN(n14320) );
  XNOR2_X1 U16110 ( .A(n14280), .B(n14279), .ZN(n14281) );
  NOR2_X1 U16111 ( .A1(n14282), .A2(n14281), .ZN(n14284) );
  NOR2_X1 U16112 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n14458), .ZN(n14283) );
  XNOR2_X1 U16113 ( .A(n14286), .B(n14285), .ZN(n14287) );
  XOR2_X1 U16114 ( .A(n14289), .B(P3_ADDR_REG_13__SCAN_IN), .Z(n14291) );
  XNOR2_X1 U16115 ( .A(n14291), .B(n14290), .ZN(n14461) );
  INV_X1 U16116 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14463) );
  NAND2_X1 U16117 ( .A1(n14470), .A2(n14471), .ZN(n14293) );
  XOR2_X1 U16118 ( .A(n14296), .B(n14295), .Z(n14297) );
  NAND2_X1 U16119 ( .A1(n14323), .A2(n14324), .ZN(n14322) );
  INV_X1 U16120 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15210) );
  XOR2_X1 U16121 ( .A(n15210), .B(P1_ADDR_REG_18__SCAN_IN), .Z(n14304) );
  NOR2_X1 U16122 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14300), .ZN(n14303) );
  NOR2_X1 U16123 ( .A1(n14333), .A2(n14301), .ZN(n14302) );
  NOR2_X1 U16124 ( .A1(n14303), .A2(n14302), .ZN(n15209) );
  XNOR2_X1 U16125 ( .A(n14304), .B(n15209), .ZN(n15017) );
  AOI21_X1 U16126 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14306) );
  OAI21_X1 U16127 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14306), 
        .ZN(U28) );
  INV_X1 U16128 ( .A(P3_RD_REG_SCAN_IN), .ZN(n15152) );
  OAI221_X1 U16129 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(n7464), .C2(n7461), .A(n15152), .ZN(U29) );
  AOI21_X1 U16130 ( .B1(n14310), .B2(n14309), .A(n14308), .ZN(n14311) );
  XOR2_X1 U16131 ( .A(n14311), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  XOR2_X1 U16132 ( .A(n14313), .B(n14312), .Z(SUB_1596_U57) );
  XOR2_X1 U16133 ( .A(n14314), .B(P2_ADDR_REG_8__SCAN_IN), .Z(SUB_1596_U55) );
  OAI21_X1 U16134 ( .B1(n14317), .B2(n14316), .A(n14315), .ZN(n14318) );
  XOR2_X1 U16135 ( .A(n14318), .B(n14734), .Z(SUB_1596_U54) );
  NOR2_X1 U16136 ( .A1(n14320), .A2(n14319), .ZN(n14321) );
  XOR2_X1 U16137 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14321), .Z(SUB_1596_U70)
         );
  OAI21_X1 U16138 ( .B1(n14324), .B2(n14323), .A(n14322), .ZN(n14325) );
  XNOR2_X1 U16139 ( .A(n14325), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  AOI21_X1 U16140 ( .B1(n12812), .B2(n14327), .A(n14326), .ZN(n14341) );
  OAI21_X1 U16141 ( .B1(n14329), .B2(P3_REG1_REG_17__SCAN_IN), .A(n14328), 
        .ZN(n14339) );
  NAND2_X1 U16142 ( .A1(n14343), .A2(n14330), .ZN(n14332) );
  OAI211_X1 U16143 ( .C1(n14333), .C2(n14975), .A(n14332), .B(n14331), .ZN(
        n14338) );
  AOI211_X1 U16144 ( .C1(n14336), .C2(n14335), .A(n14939), .B(n14334), .ZN(
        n14337) );
  AOI211_X1 U16145 ( .C1(n14954), .C2(n14339), .A(n14338), .B(n14337), .ZN(
        n14340) );
  OAI21_X1 U16146 ( .B1(n14341), .B2(n14959), .A(n14340), .ZN(P3_U3199) );
  AOI22_X1 U16147 ( .A1(n14343), .A2(n14342), .B1(n14943), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n14360) );
  OAI21_X1 U16148 ( .B1(n14346), .B2(n14345), .A(n14344), .ZN(n14352) );
  AOI21_X1 U16149 ( .B1(n14349), .B2(n14348), .A(n14347), .ZN(n14350) );
  NOR2_X1 U16150 ( .A1(n14350), .A2(n14939), .ZN(n14351) );
  AOI21_X1 U16151 ( .B1(n14954), .B2(n14352), .A(n14351), .ZN(n14359) );
  OAI221_X1 U16152 ( .B1(n14356), .B2(n14355), .C1(n14356), .C2(n14354), .A(
        n14353), .ZN(n14357) );
  NAND4_X1 U16153 ( .A1(n14360), .A2(n14359), .A3(n14358), .A4(n14357), .ZN(
        P3_U3200) );
  AOI21_X1 U16154 ( .B1(n14362), .B2(n8900), .A(n14361), .ZN(n14363) );
  AND2_X1 U16155 ( .A1(n14364), .A2(n14363), .ZN(n14368) );
  AOI22_X1 U16156 ( .A1(n15016), .A2(n14368), .B1(n8543), .B2(n15014), .ZN(
        P3_U3471) );
  AOI211_X1 U16157 ( .C1(n8900), .C2(n14367), .A(n14366), .B(n14365), .ZN(
        n14370) );
  AOI22_X1 U16158 ( .A1(n15016), .A2(n14370), .B1(n8531), .B2(n15014), .ZN(
        P3_U3470) );
  INV_X1 U16159 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14369) );
  AOI22_X1 U16160 ( .A1(n15006), .A2(n14369), .B1(n14368), .B2(n15004), .ZN(
        P3_U3426) );
  INV_X1 U16161 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14371) );
  AOI22_X1 U16162 ( .A1(n15006), .A2(n14371), .B1(n14370), .B2(n15004), .ZN(
        P3_U3423) );
  OAI21_X1 U16163 ( .B1(n14374), .B2(n14373), .A(n14372), .ZN(n14375) );
  AOI222_X1 U16164 ( .A1(n14669), .A2(n6677), .B1(n14376), .B2(n14386), .C1(
        n14375), .C2(n14384), .ZN(n14379) );
  OAI211_X1 U16165 ( .C1(n14672), .C2(n14380), .A(n14379), .B(n14378), .ZN(
        P2_U3187) );
  OAI21_X1 U16166 ( .B1(n14383), .B2(n14382), .A(n14381), .ZN(n14385) );
  AOI222_X1 U16167 ( .A1(n14669), .A2(n14388), .B1(n14387), .B2(n14386), .C1(
        n14385), .C2(n14384), .ZN(n14390) );
  OAI211_X1 U16168 ( .C1(n14672), .C2(n14391), .A(n14390), .B(n14389), .ZN(
        P2_U3198) );
  INV_X1 U16169 ( .A(n14670), .ZN(n14393) );
  OAI21_X1 U16170 ( .B1(n14393), .B2(n14837), .A(n14392), .ZN(n14395) );
  AOI211_X1 U16171 ( .C1(n14396), .C2(n14833), .A(n14395), .B(n14394), .ZN(
        n14404) );
  AOI22_X1 U16172 ( .A1(n14855), .A2(n14404), .B1(n14397), .B2(n14853), .ZN(
        P2_U3512) );
  OAI21_X1 U16173 ( .B1(n14399), .B2(n14837), .A(n14398), .ZN(n14400) );
  AOI21_X1 U16174 ( .B1(n14401), .B2(n14840), .A(n14400), .ZN(n14402) );
  AOI22_X1 U16175 ( .A1(n14855), .A2(n14405), .B1(n14736), .B2(n14853), .ZN(
        P2_U3511) );
  AOI22_X1 U16176 ( .A1(n14835), .A2(n14404), .B1(n7811), .B2(n14844), .ZN(
        P2_U3469) );
  AOI22_X1 U16177 ( .A1(n14835), .A2(n14405), .B1(n7789), .B2(n14844), .ZN(
        P2_U3466) );
  INV_X1 U16178 ( .A(n13678), .ZN(n14408) );
  OAI21_X1 U16179 ( .B1(n14408), .B2(n14407), .A(n14406), .ZN(n14410) );
  NAND2_X1 U16180 ( .A1(n14410), .A2(n14409), .ZN(n14413) );
  AOI222_X1 U16181 ( .A1(n14415), .A2(n14414), .B1(n14413), .B2(n14412), .C1(
        n14411), .C2(n14432), .ZN(n14417) );
  OAI211_X1 U16182 ( .C1(n14436), .C2(n14418), .A(n14417), .B(n14416), .ZN(
        P1_U3215) );
  OAI22_X1 U16183 ( .A1(n14422), .A2(n14421), .B1(n14420), .B2(n14419), .ZN(
        n14430) );
  AOI21_X1 U16184 ( .B1(n11800), .B2(n14424), .A(n14423), .ZN(n14425) );
  INV_X1 U16185 ( .A(n14425), .ZN(n14428) );
  AOI21_X1 U16186 ( .B1(n14428), .B2(n14427), .A(n14426), .ZN(n14429) );
  AOI211_X1 U16187 ( .C1(n14432), .C2(n14431), .A(n14430), .B(n14429), .ZN(
        n14434) );
  OAI211_X1 U16188 ( .C1(n14436), .C2(n14435), .A(n14434), .B(n14433), .ZN(
        P1_U3236) );
  OAI211_X1 U16189 ( .C1(n14439), .C2(n14640), .A(n14438), .B(n14437), .ZN(
        n14440) );
  AOI21_X1 U16190 ( .B1(n14441), .B2(n14644), .A(n14440), .ZN(n14453) );
  AOI22_X1 U16191 ( .A1(n14657), .A2(n14453), .B1(n9360), .B2(n14655), .ZN(
        P1_U3543) );
  OAI21_X1 U16192 ( .B1(n14443), .B2(n14640), .A(n14442), .ZN(n14445) );
  AOI211_X1 U16193 ( .C1(n14644), .C2(n14446), .A(n14445), .B(n14444), .ZN(
        n14455) );
  AOI22_X1 U16194 ( .A1(n14657), .A2(n14455), .B1(n10269), .B2(n14655), .ZN(
        P1_U3541) );
  OAI21_X1 U16195 ( .B1(n14448), .B2(n14640), .A(n14447), .ZN(n14449) );
  AOI21_X1 U16196 ( .B1(n14450), .B2(n14644), .A(n14449), .ZN(n14452) );
  AND2_X1 U16197 ( .A1(n14452), .A2(n14451), .ZN(n14457) );
  AOI22_X1 U16198 ( .A1(n14657), .A2(n14457), .B1(n9276), .B2(n14655), .ZN(
        P1_U3539) );
  AOI22_X1 U16199 ( .A1(n14646), .A2(n14453), .B1(n9361), .B2(n14645), .ZN(
        P1_U3504) );
  INV_X1 U16200 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14454) );
  AOI22_X1 U16201 ( .A1(n14646), .A2(n14455), .B1(n14454), .B2(n14645), .ZN(
        P1_U3498) );
  INV_X1 U16202 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14456) );
  AOI22_X1 U16203 ( .A1(n14646), .A2(n14457), .B1(n14456), .B2(n14645), .ZN(
        P1_U3492) );
  XNOR2_X1 U16204 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n14458), .ZN(SUB_1596_U69)
         );
  INV_X1 U16205 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14753) );
  XOR2_X1 U16206 ( .A(n14753), .B(n14459), .Z(SUB_1596_U68) );
  OAI21_X1 U16207 ( .B1(n14462), .B2(n14461), .A(n14460), .ZN(n14464) );
  XOR2_X1 U16208 ( .A(n14464), .B(n14463), .Z(SUB_1596_U67) );
  OAI21_X1 U16209 ( .B1(n14467), .B2(n14466), .A(n14465), .ZN(n14468) );
  XOR2_X1 U16210 ( .A(n14468), .B(n10979), .Z(SUB_1596_U66) );
  AOI21_X1 U16211 ( .B1(n14471), .B2(n14470), .A(n14469), .ZN(n14472) );
  XOR2_X1 U16212 ( .A(n14472), .B(P2_ADDR_REG_15__SCAN_IN), .Z(SUB_1596_U65)
         );
  OAI222_X1 U16213 ( .A1(n14477), .A2(n14476), .B1(n14477), .B2(n14475), .C1(
        n14474), .C2(n14473), .ZN(SUB_1596_U64) );
  MUX2_X1 U16214 ( .A(n14528), .B(P1_REG2_REG_4__SCAN_IN), .S(n14491), .Z(
        n14478) );
  NAND3_X1 U16215 ( .A1(n14480), .A2(n14479), .A3(n14478), .ZN(n14481) );
  NAND3_X1 U16216 ( .A1(n14483), .A2(n14482), .A3(n14481), .ZN(n14498) );
  INV_X1 U16217 ( .A(n14484), .ZN(n14489) );
  NAND3_X1 U16218 ( .A1(n14487), .A2(n14486), .A3(n14485), .ZN(n14488) );
  NAND3_X1 U16219 ( .A1(n14490), .A2(n14489), .A3(n14488), .ZN(n14497) );
  NAND2_X1 U16220 ( .A1(n14492), .A2(n14491), .ZN(n14496) );
  AOI21_X1 U16221 ( .B1(n14494), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n14493), .ZN(
        n14495) );
  AND4_X1 U16222 ( .A1(n14498), .A2(n14497), .A3(n14496), .A4(n14495), .ZN(
        n14500) );
  NAND2_X1 U16223 ( .A1(n14500), .A2(n14499), .ZN(P1_U3247) );
  AOI21_X1 U16224 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14502), .A(n14501), 
        .ZN(n14506) );
  AOI21_X1 U16225 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n14504), .A(n14503), 
        .ZN(n14505) );
  OAI222_X1 U16226 ( .A1(n14521), .A2(n14507), .B1(n14519), .B2(n14506), .C1(
        n14517), .C2(n14505), .ZN(n14508) );
  INV_X1 U16227 ( .A(n14508), .ZN(n14510) );
  OAI211_X1 U16228 ( .C1(n14511), .C2(n14525), .A(n14510), .B(n14509), .ZN(
        P1_U3258) );
  INV_X1 U16229 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15207) );
  OAI21_X1 U16230 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n14513), .A(n14512), 
        .ZN(n14518) );
  OAI21_X1 U16231 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n14515), .A(n14514), 
        .ZN(n14516) );
  OAI222_X1 U16232 ( .A1(n14521), .A2(n14520), .B1(n14519), .B2(n14518), .C1(
        n14517), .C2(n14516), .ZN(n14522) );
  INV_X1 U16233 ( .A(n14522), .ZN(n14524) );
  OAI211_X1 U16234 ( .C1(n15207), .C2(n14525), .A(n14524), .B(n14523), .ZN(
        P1_U3261) );
  OAI22_X1 U16235 ( .A1(n14576), .A2(n14528), .B1(n14527), .B2(n14526), .ZN(
        n14532) );
  NOR2_X1 U16236 ( .A1(n14530), .A2(n14529), .ZN(n14531) );
  AOI211_X1 U16237 ( .C1(n14533), .C2(n14558), .A(n14532), .B(n14531), .ZN(
        n14534) );
  OAI21_X1 U16238 ( .B1(n14536), .B2(n14535), .A(n14534), .ZN(n14537) );
  INV_X1 U16239 ( .A(n14537), .ZN(n14538) );
  OAI21_X1 U16240 ( .B1(n14578), .B2(n14539), .A(n14538), .ZN(P1_U3289) );
  OAI21_X1 U16241 ( .B1(n14541), .B2(n10226), .A(n14540), .ZN(n14548) );
  OAI22_X1 U16242 ( .A1(n14543), .A2(n14562), .B1(n7406), .B2(n14542), .ZN(
        n14547) );
  XNOR2_X1 U16243 ( .A(n14544), .B(n10226), .ZN(n14552) );
  NOR2_X1 U16244 ( .A1(n14552), .A2(n14545), .ZN(n14546) );
  AOI211_X1 U16245 ( .C1(n14549), .C2(n14548), .A(n14547), .B(n14546), .ZN(
        n14601) );
  AOI222_X1 U16246 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n14578), .B1(n14574), 
        .B2(n14551), .C1(n14554), .C2(n14550), .ZN(n14561) );
  INV_X1 U16247 ( .A(n14552), .ZN(n14604) );
  OAI211_X1 U16248 ( .C1(n6938), .C2(n6937), .A(n14556), .B(n14555), .ZN(
        n14600) );
  INV_X1 U16249 ( .A(n14600), .ZN(n14557) );
  AOI22_X1 U16250 ( .A1(n14604), .A2(n14559), .B1(n14558), .B2(n14557), .ZN(
        n14560) );
  OAI211_X1 U16251 ( .C1(n14578), .C2(n14601), .A(n14561), .B(n14560), .ZN(
        P1_U3290) );
  OR2_X1 U16252 ( .A1(n14563), .A2(n14562), .ZN(n14567) );
  NAND2_X1 U16253 ( .A1(n14565), .A2(n14564), .ZN(n14566) );
  NAND2_X1 U16254 ( .A1(n14567), .A2(n14566), .ZN(n14582) );
  INV_X1 U16255 ( .A(n14568), .ZN(n14569) );
  NAND2_X1 U16256 ( .A1(n14582), .A2(n14569), .ZN(n14577) );
  OAI21_X1 U16257 ( .B1(n14571), .B2(n14570), .A(n14584), .ZN(n14572) );
  INV_X1 U16258 ( .A(n14572), .ZN(n14573) );
  AOI21_X1 U16259 ( .B1(n14574), .B2(P1_REG3_REG_0__SCAN_IN), .A(n14573), .ZN(
        n14575) );
  OAI221_X1 U16260 ( .B1(n14578), .B2(n14577), .C1(n14576), .C2(n9115), .A(
        n14575), .ZN(P1_U3293) );
  AND2_X1 U16261 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14579), .ZN(P1_U3294) );
  AND2_X1 U16262 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14579), .ZN(P1_U3295) );
  AND2_X1 U16263 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14579), .ZN(P1_U3296) );
  AND2_X1 U16264 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14579), .ZN(P1_U3297) );
  AND2_X1 U16265 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14579), .ZN(P1_U3298) );
  AND2_X1 U16266 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14579), .ZN(P1_U3299) );
  AND2_X1 U16267 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14579), .ZN(P1_U3300) );
  AND2_X1 U16268 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14579), .ZN(P1_U3301) );
  AND2_X1 U16269 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14579), .ZN(P1_U3302) );
  AND2_X1 U16270 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14579), .ZN(P1_U3303) );
  AND2_X1 U16271 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14579), .ZN(P1_U3304) );
  AND2_X1 U16272 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14579), .ZN(P1_U3305) );
  AND2_X1 U16273 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14579), .ZN(P1_U3306) );
  AND2_X1 U16274 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14579), .ZN(P1_U3307) );
  AND2_X1 U16275 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14579), .ZN(P1_U3308) );
  AND2_X1 U16276 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14579), .ZN(P1_U3309) );
  AND2_X1 U16277 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14579), .ZN(P1_U3310) );
  AND2_X1 U16278 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14579), .ZN(P1_U3311) );
  AND2_X1 U16279 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14579), .ZN(P1_U3312) );
  AND2_X1 U16280 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14579), .ZN(P1_U3313) );
  AND2_X1 U16281 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14579), .ZN(P1_U3314) );
  AND2_X1 U16282 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14579), .ZN(P1_U3315) );
  AND2_X1 U16283 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14579), .ZN(P1_U3316) );
  AND2_X1 U16284 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14579), .ZN(P1_U3317) );
  AND2_X1 U16285 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14579), .ZN(P1_U3318) );
  AND2_X1 U16286 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14579), .ZN(P1_U3319) );
  AND2_X1 U16287 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14579), .ZN(P1_U3320) );
  AND2_X1 U16288 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14579), .ZN(P1_U3321) );
  AND2_X1 U16289 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14579), .ZN(P1_U3322) );
  AND2_X1 U16290 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14579), .ZN(P1_U3323) );
  NAND2_X1 U16291 ( .A1(n14581), .A2(n14580), .ZN(n14583) );
  AOI21_X1 U16292 ( .B1(n14584), .B2(n14583), .A(n14582), .ZN(n14647) );
  AOI22_X1 U16293 ( .A1(n14646), .A2(n14647), .B1(n9113), .B2(n14645), .ZN(
        P1_U3459) );
  INV_X1 U16294 ( .A(n14592), .ZN(n14588) );
  AOI21_X1 U16295 ( .B1(n14586), .B2(n14606), .A(n14585), .ZN(n14587) );
  OAI21_X1 U16296 ( .B1(n14588), .B2(n14609), .A(n14587), .ZN(n14591) );
  INV_X1 U16297 ( .A(n14589), .ZN(n14590) );
  AOI211_X1 U16298 ( .C1(n14593), .C2(n14592), .A(n14591), .B(n14590), .ZN(
        n14648) );
  AOI22_X1 U16299 ( .A1(n14646), .A2(n14648), .B1(n9103), .B2(n14645), .ZN(
        P1_U3462) );
  OAI21_X1 U16300 ( .B1(n14595), .B2(n14640), .A(n14594), .ZN(n14596) );
  AOI21_X1 U16301 ( .B1(n14597), .B2(n14636), .A(n14596), .ZN(n14598) );
  AND2_X1 U16302 ( .A1(n14599), .A2(n14598), .ZN(n14649) );
  AOI22_X1 U16303 ( .A1(n14646), .A2(n14649), .B1(n9135), .B2(n14645), .ZN(
        P1_U3465) );
  OAI21_X1 U16304 ( .B1(n6937), .B2(n14640), .A(n14600), .ZN(n14603) );
  INV_X1 U16305 ( .A(n14601), .ZN(n14602) );
  AOI211_X1 U16306 ( .C1(n14636), .C2(n14604), .A(n14603), .B(n14602), .ZN(
        n14650) );
  AOI22_X1 U16307 ( .A1(n14646), .A2(n14650), .B1(n6649), .B2(n14645), .ZN(
        P1_U3468) );
  AOI21_X1 U16308 ( .B1(n14607), .B2(n14606), .A(n14605), .ZN(n14608) );
  OAI21_X1 U16309 ( .B1(n14610), .B2(n14609), .A(n14608), .ZN(n14611) );
  NOR2_X1 U16310 ( .A1(n14612), .A2(n14611), .ZN(n14651) );
  INV_X1 U16311 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14613) );
  AOI22_X1 U16312 ( .A1(n14646), .A2(n14651), .B1(n14613), .B2(n14645), .ZN(
        P1_U3477) );
  NAND3_X1 U16313 ( .A1(n14616), .A2(n14615), .A3(n14614), .ZN(n14619) );
  INV_X1 U16314 ( .A(n14617), .ZN(n14618) );
  AOI211_X1 U16315 ( .C1(n14644), .C2(n14620), .A(n14619), .B(n14618), .ZN(
        n14652) );
  AOI22_X1 U16316 ( .A1(n14646), .A2(n14652), .B1(n9211), .B2(n14645), .ZN(
        P1_U3480) );
  INV_X1 U16317 ( .A(n14621), .ZN(n14622) );
  NAND3_X1 U16318 ( .A1(n14624), .A2(n14623), .A3(n14622), .ZN(n14627) );
  INV_X1 U16319 ( .A(n14625), .ZN(n14626) );
  AOI211_X1 U16320 ( .C1(n14644), .C2(n14628), .A(n14627), .B(n14626), .ZN(
        n14653) );
  INV_X1 U16321 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14629) );
  AOI22_X1 U16322 ( .A1(n14646), .A2(n14653), .B1(n14629), .B2(n14645), .ZN(
        P1_U3483) );
  INV_X1 U16323 ( .A(n14630), .ZN(n14631) );
  NAND2_X1 U16324 ( .A1(n14632), .A2(n14631), .ZN(n14634) );
  AOI211_X1 U16325 ( .C1(n14636), .C2(n14635), .A(n14634), .B(n14633), .ZN(
        n14654) );
  INV_X1 U16326 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14637) );
  AOI22_X1 U16327 ( .A1(n14646), .A2(n14654), .B1(n14637), .B2(n14645), .ZN(
        P1_U3486) );
  OAI211_X1 U16328 ( .C1(n14641), .C2(n14640), .A(n14639), .B(n14638), .ZN(
        n14642) );
  AOI21_X1 U16329 ( .B1(n14644), .B2(n14643), .A(n14642), .ZN(n14656) );
  AOI22_X1 U16330 ( .A1(n14646), .A2(n14656), .B1(n9266), .B2(n14645), .ZN(
        P1_U3489) );
  AOI22_X1 U16331 ( .A1(n14657), .A2(n14647), .B1(n9738), .B2(n14655), .ZN(
        P1_U3528) );
  AOI22_X1 U16332 ( .A1(n14657), .A2(n14648), .B1(n9766), .B2(n14655), .ZN(
        P1_U3529) );
  AOI22_X1 U16333 ( .A1(n14657), .A2(n14649), .B1(n9765), .B2(n14655), .ZN(
        P1_U3530) );
  AOI22_X1 U16334 ( .A1(n14657), .A2(n14650), .B1(n9770), .B2(n14655), .ZN(
        P1_U3531) );
  AOI22_X1 U16335 ( .A1(n14657), .A2(n14651), .B1(n9803), .B2(n14655), .ZN(
        P1_U3534) );
  AOI22_X1 U16336 ( .A1(n14657), .A2(n14652), .B1(n9806), .B2(n14655), .ZN(
        P1_U3535) );
  AOI22_X1 U16337 ( .A1(n14657), .A2(n14653), .B1(n9807), .B2(n14655), .ZN(
        P1_U3536) );
  AOI22_X1 U16338 ( .A1(n14657), .A2(n14654), .B1(n9249), .B2(n14655), .ZN(
        P1_U3537) );
  AOI22_X1 U16339 ( .A1(n14657), .A2(n14656), .B1(n9265), .B2(n14655), .ZN(
        P1_U3538) );
  NOR2_X1 U16340 ( .A1(n14775), .A2(P2_U3947), .ZN(P2_U3087) );
  OAI22_X1 U16341 ( .A1(n14660), .A2(n14659), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14658), .ZN(n14668) );
  NAND2_X1 U16342 ( .A1(n11829), .A2(n14661), .ZN(n14665) );
  INV_X1 U16343 ( .A(n14662), .ZN(n14663) );
  AOI211_X1 U16344 ( .C1(n14666), .C2(n14665), .A(n14664), .B(n14663), .ZN(
        n14667) );
  AOI211_X1 U16345 ( .C1(n14670), .C2(n14669), .A(n14668), .B(n14667), .ZN(
        n14671) );
  OAI21_X1 U16346 ( .B1(n14673), .B2(n14672), .A(n14671), .ZN(P2_U3206) );
  AOI21_X1 U16347 ( .B1(n14783), .B2(P2_REG1_REG_0__SCAN_IN), .A(n14674), .ZN(
        n14678) );
  AOI22_X1 U16348 ( .A1(n14775), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14677) );
  OAI22_X1 U16349 ( .A1(n14713), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n14746), .ZN(n14675) );
  OAI21_X1 U16350 ( .B1(n14776), .B2(n14675), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n14676) );
  OAI211_X1 U16351 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n14678), .A(n14677), .B(
        n14676), .ZN(P2_U3214) );
  INV_X1 U16352 ( .A(n14680), .ZN(n14682) );
  OAI21_X1 U16353 ( .B1(n14682), .B2(n14681), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14683) );
  OAI21_X1 U16354 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n14683), .ZN(n14693) );
  OAI211_X1 U16355 ( .C1(n14686), .C2(n14685), .A(n14778), .B(n14684), .ZN(
        n14692) );
  NAND2_X1 U16356 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(n14775), .ZN(n14691) );
  OAI211_X1 U16357 ( .C1(n14689), .C2(n14688), .A(n14783), .B(n14687), .ZN(
        n14690) );
  NAND4_X1 U16358 ( .A1(n14693), .A2(n14692), .A3(n14691), .A4(n14690), .ZN(
        P2_U3216) );
  OAI22_X1 U16359 ( .A1(n14707), .A2(n14695), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14694), .ZN(n14696) );
  AOI21_X1 U16360 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n14775), .A(n14696), .ZN(
        n14705) );
  OAI211_X1 U16361 ( .C1(n14699), .C2(n14698), .A(n14778), .B(n14697), .ZN(
        n14704) );
  OAI211_X1 U16362 ( .C1(n14702), .C2(n14701), .A(n14783), .B(n14700), .ZN(
        n14703) );
  NAND3_X1 U16363 ( .A1(n14705), .A2(n14704), .A3(n14703), .ZN(P2_U3217) );
  NOR2_X1 U16364 ( .A1(n14707), .A2(n14706), .ZN(n14708) );
  AOI211_X1 U16365 ( .C1(n14775), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n14709), .B(
        n14708), .ZN(n14720) );
  OAI211_X1 U16366 ( .C1(n14712), .C2(n14711), .A(n14783), .B(n14710), .ZN(
        n14719) );
  AOI211_X1 U16367 ( .C1(n14716), .C2(n14715), .A(n14714), .B(n14713), .ZN(
        n14717) );
  INV_X1 U16368 ( .A(n14717), .ZN(n14718) );
  NAND3_X1 U16369 ( .A1(n14720), .A2(n14719), .A3(n14718), .ZN(P2_U3219) );
  INV_X1 U16370 ( .A(n14721), .ZN(n14725) );
  MUX2_X1 U16371 ( .A(n10097), .B(P2_REG1_REG_9__SCAN_IN), .S(n14722), .Z(
        n14724) );
  OAI21_X1 U16372 ( .B1(n14725), .B2(n14724), .A(n14723), .ZN(n14731) );
  OAI21_X1 U16373 ( .B1(n14728), .B2(n14727), .A(n14726), .ZN(n14729) );
  AOI222_X1 U16374 ( .A1(n14731), .A2(n14783), .B1(n14730), .B2(n14776), .C1(
        n14729), .C2(n14778), .ZN(n14733) );
  OAI211_X1 U16375 ( .C1(n14734), .C2(n14752), .A(n14733), .B(n14732), .ZN(
        P2_U3223) );
  NOR2_X1 U16376 ( .A1(n14749), .A2(n14736), .ZN(n14735) );
  AOI21_X1 U16377 ( .B1(n14736), .B2(n14749), .A(n14735), .ZN(n14739) );
  AOI21_X1 U16378 ( .B1(n14739), .B2(n14738), .A(n14737), .ZN(n14747) );
  AND3_X1 U16379 ( .A1(n14742), .A2(n14741), .A3(n14740), .ZN(n14743) );
  OAI21_X1 U16380 ( .B1(n14744), .B2(n14743), .A(n14778), .ZN(n14745) );
  OAI21_X1 U16381 ( .B1(n14747), .B2(n14746), .A(n14745), .ZN(n14748) );
  AOI21_X1 U16382 ( .B1(n14749), .B2(n14776), .A(n14748), .ZN(n14751) );
  OAI211_X1 U16383 ( .C1(n14753), .C2(n14752), .A(n14751), .B(n14750), .ZN(
        P2_U3226) );
  AOI22_X1 U16384 ( .A1(n14775), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n14764) );
  NAND2_X1 U16385 ( .A1(n14776), .A2(n14754), .ZN(n14763) );
  OAI211_X1 U16386 ( .C1(n14757), .C2(n14756), .A(n14783), .B(n14755), .ZN(
        n14762) );
  OAI211_X1 U16387 ( .C1(n14760), .C2(n14759), .A(n14778), .B(n14758), .ZN(
        n14761) );
  NAND4_X1 U16388 ( .A1(n14764), .A2(n14763), .A3(n14762), .A4(n14761), .ZN(
        P2_U3227) );
  AOI22_X1 U16389 ( .A1(n14775), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14773) );
  NAND2_X1 U16390 ( .A1(n14776), .A2(n14765), .ZN(n14772) );
  OAI211_X1 U16391 ( .C1(n14767), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14778), 
        .B(n14766), .ZN(n14771) );
  OAI211_X1 U16392 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n14769), .A(n14783), 
        .B(n14768), .ZN(n14770) );
  NAND4_X1 U16393 ( .A1(n14773), .A2(n14772), .A3(n14771), .A4(n14770), .ZN(
        P2_U3229) );
  AOI22_X1 U16394 ( .A1(n14775), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n14789) );
  NAND2_X1 U16395 ( .A1(n14777), .A2(n14776), .ZN(n14788) );
  OAI211_X1 U16396 ( .C1(n14781), .C2(n14780), .A(n14779), .B(n14778), .ZN(
        n14787) );
  OAI211_X1 U16397 ( .C1(n14785), .C2(n14784), .A(n14783), .B(n14782), .ZN(
        n14786) );
  NAND4_X1 U16398 ( .A1(n14789), .A2(n14788), .A3(n14787), .A4(n14786), .ZN(
        P2_U3231) );
  NAND2_X1 U16399 ( .A1(n14795), .A2(n14790), .ZN(n14791) );
  AND2_X1 U16400 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14791), .ZN(P2_U3266) );
  AND2_X1 U16401 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14791), .ZN(P2_U3267) );
  AND2_X1 U16402 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14791), .ZN(P2_U3268) );
  AND2_X1 U16403 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14791), .ZN(P2_U3269) );
  AND2_X1 U16404 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14791), .ZN(P2_U3270) );
  AND2_X1 U16405 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14791), .ZN(P2_U3271) );
  AND2_X1 U16406 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14791), .ZN(P2_U3272) );
  AND2_X1 U16407 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14791), .ZN(P2_U3273) );
  AND2_X1 U16408 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14791), .ZN(P2_U3274) );
  AND2_X1 U16409 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14791), .ZN(P2_U3275) );
  AND2_X1 U16410 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14791), .ZN(P2_U3276) );
  AND2_X1 U16411 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14791), .ZN(P2_U3277) );
  AND2_X1 U16412 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14791), .ZN(P2_U3278) );
  AND2_X1 U16413 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14791), .ZN(P2_U3279) );
  AND2_X1 U16414 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14791), .ZN(P2_U3280) );
  AND2_X1 U16415 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14791), .ZN(P2_U3281) );
  AND2_X1 U16416 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14791), .ZN(P2_U3282) );
  AND2_X1 U16417 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14791), .ZN(P2_U3283) );
  AND2_X1 U16418 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14791), .ZN(P2_U3284) );
  AND2_X1 U16419 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14791), .ZN(P2_U3285) );
  AND2_X1 U16420 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14791), .ZN(P2_U3286) );
  AND2_X1 U16421 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14791), .ZN(P2_U3287) );
  AND2_X1 U16422 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14791), .ZN(P2_U3288) );
  AND2_X1 U16423 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14791), .ZN(P2_U3289) );
  AND2_X1 U16424 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14791), .ZN(P2_U3290) );
  AND2_X1 U16425 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14791), .ZN(P2_U3291) );
  AND2_X1 U16426 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14791), .ZN(P2_U3292) );
  AND2_X1 U16427 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14791), .ZN(P2_U3293) );
  AND2_X1 U16428 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14791), .ZN(P2_U3294) );
  AND2_X1 U16429 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14791), .ZN(P2_U3295) );
  MUX2_X1 U16430 ( .A(n14792), .B(P2_D_REG_0__SCAN_IN), .S(n14791), .Z(
        P2_U3416) );
  INV_X1 U16431 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14794) );
  OAI21_X1 U16432 ( .B1(n14795), .B2(n14794), .A(n14793), .ZN(P2_U3417) );
  OAI211_X1 U16433 ( .C1(n14798), .C2(n14819), .A(n14797), .B(n14796), .ZN(
        n14799) );
  INV_X1 U16434 ( .A(n14799), .ZN(n14846) );
  INV_X1 U16435 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14800) );
  AOI22_X1 U16436 ( .A1(n14835), .A2(n14846), .B1(n14800), .B2(n14844), .ZN(
        P2_U3430) );
  AOI21_X1 U16437 ( .B1(n14816), .B2(n14802), .A(n14801), .ZN(n14803) );
  OAI211_X1 U16438 ( .C1(n14805), .C2(n14812), .A(n14804), .B(n14803), .ZN(
        n14806) );
  INV_X1 U16439 ( .A(n14806), .ZN(n14847) );
  AOI22_X1 U16440 ( .A1(n14835), .A2(n14847), .B1(n7594), .B2(n14844), .ZN(
        P2_U3442) );
  AOI21_X1 U16441 ( .B1(n14816), .B2(n14808), .A(n14807), .ZN(n14810) );
  OAI211_X1 U16442 ( .C1(n14812), .C2(n14811), .A(n14810), .B(n14809), .ZN(
        n14813) );
  INV_X1 U16443 ( .A(n14813), .ZN(n14848) );
  AOI22_X1 U16444 ( .A1(n14835), .A2(n14848), .B1(n7620), .B2(n14844), .ZN(
        P2_U3445) );
  INV_X1 U16445 ( .A(n14818), .ZN(n14822) );
  AOI21_X1 U16446 ( .B1(n14816), .B2(n14815), .A(n14814), .ZN(n14817) );
  OAI21_X1 U16447 ( .B1(n14819), .B2(n14818), .A(n14817), .ZN(n14820) );
  AOI211_X1 U16448 ( .C1(n14823), .C2(n14822), .A(n14821), .B(n14820), .ZN(
        n14849) );
  AOI22_X1 U16449 ( .A1(n14835), .A2(n14849), .B1(n7643), .B2(n14844), .ZN(
        P2_U3448) );
  OAI211_X1 U16450 ( .C1(n14826), .C2(n14837), .A(n14825), .B(n14824), .ZN(
        n14827) );
  AOI21_X1 U16451 ( .B1(n14833), .B2(n14828), .A(n14827), .ZN(n14850) );
  AOI22_X1 U16452 ( .A1(n14835), .A2(n14850), .B1(n7667), .B2(n14844), .ZN(
        P2_U3451) );
  OAI21_X1 U16453 ( .B1(n14830), .B2(n14837), .A(n14829), .ZN(n14832) );
  AOI211_X1 U16454 ( .C1(n14834), .C2(n14833), .A(n14832), .B(n14831), .ZN(
        n14852) );
  AOI22_X1 U16455 ( .A1(n14835), .A2(n14852), .B1(n7738), .B2(n14844), .ZN(
        P2_U3460) );
  OAI21_X1 U16456 ( .B1(n14838), .B2(n14837), .A(n14836), .ZN(n14839) );
  AOI21_X1 U16457 ( .B1(n14841), .B2(n14840), .A(n14839), .ZN(n14842) );
  AOI22_X1 U16458 ( .A1(n14835), .A2(n14854), .B1(n7767), .B2(n14844), .ZN(
        P2_U3463) );
  AOI22_X1 U16459 ( .A1(n14855), .A2(n14846), .B1(n14845), .B2(n14853), .ZN(
        P2_U3499) );
  AOI22_X1 U16460 ( .A1(n14855), .A2(n14847), .B1(n9832), .B2(n14853), .ZN(
        P2_U3503) );
  AOI22_X1 U16461 ( .A1(n14855), .A2(n14848), .B1(n9836), .B2(n14853), .ZN(
        P2_U3504) );
  AOI22_X1 U16462 ( .A1(n14855), .A2(n14849), .B1(n9837), .B2(n14853), .ZN(
        P2_U3505) );
  AOI22_X1 U16463 ( .A1(n14855), .A2(n14850), .B1(n9840), .B2(n14853), .ZN(
        P2_U3506) );
  AOI22_X1 U16464 ( .A1(n14855), .A2(n14852), .B1(n14851), .B2(n14853), .ZN(
        P2_U3509) );
  AOI22_X1 U16465 ( .A1(n14855), .A2(n14854), .B1(n10981), .B2(n14853), .ZN(
        P2_U3510) );
  NOR2_X1 U16466 ( .A1(P3_U3897), .A2(n14943), .ZN(P3_U3150) );
  INV_X1 U16467 ( .A(n14856), .ZN(n14858) );
  AOI21_X1 U16468 ( .B1(n14859), .B2(n14858), .A(n14857), .ZN(n14873) );
  INV_X1 U16469 ( .A(n14861), .ZN(n14877) );
  AND2_X1 U16470 ( .A1(n14861), .A2(n14860), .ZN(n14863) );
  OAI22_X1 U16471 ( .A1(n14880), .A2(n14877), .B1(n14863), .B2(n14862), .ZN(
        n14868) );
  AOI21_X1 U16472 ( .B1(n14943), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n14864), .ZN(
        n14865) );
  OAI21_X1 U16473 ( .B1(n14970), .B2(n14866), .A(n14865), .ZN(n14867) );
  AOI21_X1 U16474 ( .B1(n14868), .B2(n14964), .A(n14867), .ZN(n14872) );
  XOR2_X1 U16475 ( .A(P3_REG1_REG_5__SCAN_IN), .B(n14869), .Z(n14870) );
  NAND2_X1 U16476 ( .A1(n14954), .A2(n14870), .ZN(n14871) );
  OAI211_X1 U16477 ( .C1(n14873), .C2(n14959), .A(n14872), .B(n14871), .ZN(
        P3_U3187) );
  AOI21_X1 U16478 ( .B1(n14876), .B2(n14875), .A(n14874), .ZN(n14892) );
  NOR2_X1 U16479 ( .A1(n14878), .A2(n14877), .ZN(n14881) );
  INV_X1 U16480 ( .A(n14899), .ZN(n14879) );
  AOI21_X1 U16481 ( .B1(n14881), .B2(n14880), .A(n14879), .ZN(n14883) );
  OAI22_X1 U16482 ( .A1(n14883), .A2(n14939), .B1(n14882), .B2(n14970), .ZN(
        n14884) );
  AOI211_X1 U16483 ( .C1(P3_ADDR_REG_6__SCAN_IN), .C2(n14943), .A(n14885), .B(
        n14884), .ZN(n14891) );
  OAI21_X1 U16484 ( .B1(n14888), .B2(n14887), .A(n14886), .ZN(n14889) );
  NAND2_X1 U16485 ( .A1(n14954), .A2(n14889), .ZN(n14890) );
  OAI211_X1 U16486 ( .C1(n14892), .C2(n14959), .A(n14891), .B(n14890), .ZN(
        P3_U3188) );
  AOI21_X1 U16487 ( .B1(n11421), .B2(n14894), .A(n14893), .ZN(n14910) );
  INV_X1 U16488 ( .A(n14895), .ZN(n14896) );
  NOR2_X1 U16489 ( .A1(n14897), .A2(n14896), .ZN(n14900) );
  INV_X1 U16490 ( .A(n14917), .ZN(n14898) );
  AOI21_X1 U16491 ( .B1(n14900), .B2(n14899), .A(n14898), .ZN(n14902) );
  OAI22_X1 U16492 ( .A1(n14902), .A2(n14939), .B1(n14901), .B2(n14970), .ZN(
        n14903) );
  AOI211_X1 U16493 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n14943), .A(n14904), .B(
        n14903), .ZN(n14909) );
  OAI21_X1 U16494 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n14906), .A(n14905), .ZN(
        n14907) );
  NAND2_X1 U16495 ( .A1(n14907), .A2(n14954), .ZN(n14908) );
  OAI211_X1 U16496 ( .C1(n14910), .C2(n14959), .A(n14909), .B(n14908), .ZN(
        P3_U3189) );
  AOI21_X1 U16497 ( .B1(n6627), .B2(n14912), .A(n14911), .ZN(n14929) );
  INV_X1 U16498 ( .A(n14913), .ZN(n14914) );
  NOR2_X1 U16499 ( .A1(n14915), .A2(n14914), .ZN(n14918) );
  INV_X1 U16500 ( .A(n14936), .ZN(n14916) );
  AOI21_X1 U16501 ( .B1(n14918), .B2(n14917), .A(n14916), .ZN(n14920) );
  OAI22_X1 U16502 ( .A1(n14920), .A2(n14939), .B1(n14919), .B2(n14970), .ZN(
        n14921) );
  AOI211_X1 U16503 ( .C1(P3_ADDR_REG_8__SCAN_IN), .C2(n14943), .A(n14922), .B(
        n14921), .ZN(n14928) );
  OAI21_X1 U16504 ( .B1(n14925), .B2(n14924), .A(n14923), .ZN(n14926) );
  NAND2_X1 U16505 ( .A1(n14926), .A2(n14954), .ZN(n14927) );
  OAI211_X1 U16506 ( .C1(n14929), .C2(n14959), .A(n14928), .B(n14927), .ZN(
        P3_U3190) );
  AOI21_X1 U16507 ( .B1(n11434), .B2(n14931), .A(n14930), .ZN(n14949) );
  INV_X1 U16508 ( .A(n14932), .ZN(n14933) );
  NOR2_X1 U16509 ( .A1(n14934), .A2(n14933), .ZN(n14937) );
  INV_X1 U16510 ( .A(n14963), .ZN(n14935) );
  AOI21_X1 U16511 ( .B1(n14937), .B2(n14936), .A(n14935), .ZN(n14940) );
  OAI22_X1 U16512 ( .A1(n14940), .A2(n14939), .B1(n14938), .B2(n14970), .ZN(
        n14941) );
  AOI211_X1 U16513 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n14943), .A(n14942), .B(
        n14941), .ZN(n14948) );
  OAI21_X1 U16514 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n14945), .A(n14944), .ZN(
        n14946) );
  NAND2_X1 U16515 ( .A1(n14946), .A2(n14954), .ZN(n14947) );
  OAI211_X1 U16516 ( .C1(n14949), .C2(n14959), .A(n14948), .B(n14947), .ZN(
        P3_U3191) );
  OAI21_X1 U16517 ( .B1(n14952), .B2(n14951), .A(n14950), .ZN(n14955) );
  AOI21_X1 U16518 ( .B1(n14955), .B2(n14954), .A(n14953), .ZN(n14973) );
  AOI21_X1 U16519 ( .B1(n14958), .B2(n14957), .A(n14956), .ZN(n14960) );
  OR2_X1 U16520 ( .A1(n14960), .A2(n14959), .ZN(n14968) );
  AND3_X1 U16521 ( .A1(n14963), .A2(n14962), .A3(n14961), .ZN(n14965) );
  OAI21_X1 U16522 ( .B1(n14966), .B2(n14965), .A(n14964), .ZN(n14967) );
  OAI211_X1 U16523 ( .C1(n14970), .C2(n14969), .A(n14968), .B(n14967), .ZN(
        n14971) );
  INV_X1 U16524 ( .A(n14971), .ZN(n14972) );
  OAI211_X1 U16525 ( .C1(n14975), .C2(n14974), .A(n14973), .B(n14972), .ZN(
        P3_U3192) );
  INV_X1 U16526 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n14981) );
  OAI21_X1 U16527 ( .B1(n14978), .B2(n14977), .A(n14976), .ZN(n14979) );
  NOR2_X1 U16528 ( .A1(n14980), .A2(n14979), .ZN(n15007) );
  AOI22_X1 U16529 ( .A1(n15006), .A2(n14981), .B1(n15007), .B2(n15004), .ZN(
        P3_U3393) );
  INV_X1 U16530 ( .A(n14982), .ZN(n14984) );
  AOI211_X1 U16531 ( .C1(n14997), .C2(n14985), .A(n14984), .B(n14983), .ZN(
        n15008) );
  AOI22_X1 U16532 ( .A1(n15006), .A2(n8409), .B1(n15008), .B2(n15004), .ZN(
        P3_U3396) );
  INV_X1 U16533 ( .A(n14986), .ZN(n14988) );
  AOI211_X1 U16534 ( .C1(n14989), .C2(n8900), .A(n14988), .B(n14987), .ZN(
        n15010) );
  AOI22_X1 U16535 ( .A1(n15006), .A2(n8432), .B1(n15010), .B2(n15004), .ZN(
        P3_U3402) );
  INV_X1 U16536 ( .A(n14990), .ZN(n14994) );
  INV_X1 U16537 ( .A(n14991), .ZN(n14992) );
  AOI211_X1 U16538 ( .C1(n14994), .C2(n8900), .A(n14993), .B(n14992), .ZN(
        n15012) );
  AOI22_X1 U16539 ( .A1(n15006), .A2(n8445), .B1(n15012), .B2(n15004), .ZN(
        P3_U3405) );
  INV_X1 U16540 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n14999) );
  AOI211_X1 U16541 ( .C1(n14998), .C2(n14997), .A(n14996), .B(n14995), .ZN(
        n15013) );
  AOI22_X1 U16542 ( .A1(n15006), .A2(n14999), .B1(n15013), .B2(n15004), .ZN(
        P3_U3414) );
  INV_X1 U16543 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15005) );
  NAND2_X1 U16544 ( .A1(n15000), .A2(n8900), .ZN(n15001) );
  AND3_X1 U16545 ( .A1(n15003), .A2(n15002), .A3(n15001), .ZN(n15015) );
  AOI22_X1 U16546 ( .A1(n15006), .A2(n15005), .B1(n15015), .B2(n15004), .ZN(
        P3_U3420) );
  AOI22_X1 U16547 ( .A1(n15016), .A2(n15007), .B1(n10408), .B2(n15014), .ZN(
        P3_U3460) );
  AOI22_X1 U16548 ( .A1(n15016), .A2(n15008), .B1(n10350), .B2(n15014), .ZN(
        P3_U3461) );
  AOI22_X1 U16549 ( .A1(n15016), .A2(n15010), .B1(n15009), .B2(n15014), .ZN(
        P3_U3463) );
  AOI22_X1 U16550 ( .A1(n15016), .A2(n15012), .B1(n15011), .B2(n15014), .ZN(
        P3_U3464) );
  AOI22_X1 U16551 ( .A1(n15016), .A2(n15013), .B1(n11427), .B2(n15014), .ZN(
        P3_U3467) );
  AOI22_X1 U16552 ( .A1(n15016), .A2(n15015), .B1(n11440), .B2(n15014), .ZN(
        P3_U3469) );
  AOI22_X1 U16553 ( .A1(SI_25_), .A2(keyinput_f7), .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .ZN(n15020) );
  OAI221_X1 U16554 ( .B1(SI_25_), .B2(keyinput_f7), .C1(
        P3_REG3_REG_19__SCAN_IN), .C2(keyinput_f41), .A(n15020), .ZN(n15027)
         );
  AOI22_X1 U16555 ( .A1(SI_12_), .A2(keyinput_f20), .B1(
        P3_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .ZN(n15021) );
  OAI221_X1 U16556 ( .B1(SI_12_), .B2(keyinput_f20), .C1(
        P3_REG3_REG_21__SCAN_IN), .C2(keyinput_f45), .A(n15021), .ZN(n15026)
         );
  AOI22_X1 U16557 ( .A1(SI_29_), .A2(keyinput_f3), .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .ZN(n15022) );
  OAI221_X1 U16558 ( .B1(SI_29_), .B2(keyinput_f3), .C1(
        P3_REG3_REG_17__SCAN_IN), .C2(keyinput_f50), .A(n15022), .ZN(n15025)
         );
  AOI22_X1 U16559 ( .A1(SI_10_), .A2(keyinput_f22), .B1(SI_28_), .B2(
        keyinput_f4), .ZN(n15023) );
  OAI221_X1 U16560 ( .B1(SI_10_), .B2(keyinput_f22), .C1(SI_28_), .C2(
        keyinput_f4), .A(n15023), .ZN(n15024) );
  NOR4_X1 U16561 ( .A1(n15027), .A2(n15026), .A3(n15025), .A4(n15024), .ZN(
        n15054) );
  XNOR2_X1 U16562 ( .A(n15134), .B(keyinput_f39), .ZN(n15034) );
  AOI22_X1 U16563 ( .A1(SI_31_), .A2(keyinput_f1), .B1(P3_REG3_REG_5__SCAN_IN), 
        .B2(keyinput_f49), .ZN(n15028) );
  OAI221_X1 U16564 ( .B1(SI_31_), .B2(keyinput_f1), .C1(P3_REG3_REG_5__SCAN_IN), .C2(keyinput_f49), .A(n15028), .ZN(n15033) );
  AOI22_X1 U16565 ( .A1(SI_22_), .A2(keyinput_f10), .B1(
        P3_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .ZN(n15029) );
  OAI221_X1 U16566 ( .B1(SI_22_), .B2(keyinput_f10), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_f60), .A(n15029), .ZN(n15032)
         );
  AOI22_X1 U16567 ( .A1(SI_8_), .A2(keyinput_f24), .B1(P3_REG3_REG_4__SCAN_IN), 
        .B2(keyinput_f52), .ZN(n15030) );
  OAI221_X1 U16568 ( .B1(SI_8_), .B2(keyinput_f24), .C1(P3_REG3_REG_4__SCAN_IN), .C2(keyinput_f52), .A(n15030), .ZN(n15031) );
  NOR4_X1 U16569 ( .A1(n15034), .A2(n15033), .A3(n15032), .A4(n15031), .ZN(
        n15053) );
  AOI22_X1 U16570 ( .A1(SI_17_), .A2(keyinput_f15), .B1(SI_19_), .B2(
        keyinput_f13), .ZN(n15035) );
  OAI221_X1 U16571 ( .B1(SI_17_), .B2(keyinput_f15), .C1(SI_19_), .C2(
        keyinput_f13), .A(n15035), .ZN(n15042) );
  AOI22_X1 U16572 ( .A1(SI_4_), .A2(keyinput_f28), .B1(P3_STATE_REG_SCAN_IN), 
        .B2(keyinput_f34), .ZN(n15036) );
  OAI221_X1 U16573 ( .B1(SI_4_), .B2(keyinput_f28), .C1(P3_STATE_REG_SCAN_IN), 
        .C2(keyinput_f34), .A(n15036), .ZN(n15041) );
  AOI22_X1 U16574 ( .A1(SI_6_), .A2(keyinput_f26), .B1(P3_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .ZN(n15037) );
  OAI221_X1 U16575 ( .B1(SI_6_), .B2(keyinput_f26), .C1(
        P3_REG3_REG_25__SCAN_IN), .C2(keyinput_f47), .A(n15037), .ZN(n15040)
         );
  AOI22_X1 U16576 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput_f59), .B1(
        P3_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .ZN(n15038) );
  OAI221_X1 U16577 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_f59), .C1(
        P3_REG3_REG_20__SCAN_IN), .C2(keyinput_f55), .A(n15038), .ZN(n15039)
         );
  NOR4_X1 U16578 ( .A1(n15042), .A2(n15041), .A3(n15040), .A4(n15039), .ZN(
        n15052) );
  AOI22_X1 U16579 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(
        P3_REG3_REG_16__SCAN_IN), .B2(keyinput_f48), .ZN(n15043) );
  OAI221_X1 U16580 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(
        P3_REG3_REG_16__SCAN_IN), .C2(keyinput_f48), .A(n15043), .ZN(n15050)
         );
  AOI22_X1 U16581 ( .A1(SI_23_), .A2(keyinput_f9), .B1(P3_REG3_REG_9__SCAN_IN), 
        .B2(keyinput_f53), .ZN(n15044) );
  OAI221_X1 U16582 ( .B1(SI_23_), .B2(keyinput_f9), .C1(P3_REG3_REG_9__SCAN_IN), .C2(keyinput_f53), .A(n15044), .ZN(n15049) );
  AOI22_X1 U16583 ( .A1(SI_21_), .A2(keyinput_f11), .B1(SI_24_), .B2(
        keyinput_f8), .ZN(n15045) );
  OAI221_X1 U16584 ( .B1(SI_21_), .B2(keyinput_f11), .C1(SI_24_), .C2(
        keyinput_f8), .A(n15045), .ZN(n15048) );
  AOI22_X1 U16585 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(
        P3_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .ZN(n15046) );
  OAI221_X1 U16586 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        P3_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(n15046), .ZN(n15047)
         );
  NOR4_X1 U16587 ( .A1(n15050), .A2(n15049), .A3(n15048), .A4(n15047), .ZN(
        n15051) );
  NAND4_X1 U16588 ( .A1(n15054), .A2(n15053), .A3(n15052), .A4(n15051), .ZN(
        n15104) );
  INV_X1 U16589 ( .A(P3_WR_REG_SCAN_IN), .ZN(n15056) );
  AOI22_X1 U16590 ( .A1(n15057), .A2(keyinput_f57), .B1(keyinput_f0), .B2(
        n15056), .ZN(n15055) );
  OAI221_X1 U16591 ( .B1(n15057), .B2(keyinput_f57), .C1(n15056), .C2(
        keyinput_f0), .A(n15055), .ZN(n15066) );
  AOI22_X1 U16592 ( .A1(n15126), .A2(keyinput_f14), .B1(n15059), .B2(
        keyinput_f5), .ZN(n15058) );
  OAI221_X1 U16593 ( .B1(n15126), .B2(keyinput_f14), .C1(n15059), .C2(
        keyinput_f5), .A(n15058), .ZN(n15065) );
  XOR2_X1 U16594 ( .A(n10877), .B(keyinput_f44), .Z(n15063) );
  INV_X1 U16595 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n15132) );
  XOR2_X1 U16596 ( .A(n15132), .B(keyinput_f38), .Z(n15062) );
  XNOR2_X1 U16597 ( .A(SI_7_), .B(keyinput_f25), .ZN(n15061) );
  XNOR2_X1 U16598 ( .A(SI_0_), .B(keyinput_f32), .ZN(n15060) );
  NAND4_X1 U16599 ( .A1(n15063), .A2(n15062), .A3(n15061), .A4(n15060), .ZN(
        n15064) );
  NOR3_X1 U16600 ( .A1(n15066), .A2(n15065), .A3(n15064), .ZN(n15102) );
  AOI22_X1 U16601 ( .A1(n15068), .A2(keyinput_f17), .B1(n8373), .B2(
        keyinput_f63), .ZN(n15067) );
  OAI221_X1 U16602 ( .B1(n15068), .B2(keyinput_f17), .C1(n8373), .C2(
        keyinput_f63), .A(n15067), .ZN(n15076) );
  AOI22_X1 U16603 ( .A1(n15149), .A2(keyinput_f35), .B1(keyinput_f18), .B2(
        n7301), .ZN(n15069) );
  OAI221_X1 U16604 ( .B1(n15149), .B2(keyinput_f35), .C1(n7301), .C2(
        keyinput_f18), .A(n15069), .ZN(n15075) );
  AOI22_X1 U16605 ( .A1(n15107), .A2(keyinput_f56), .B1(keyinput_f2), .B2(
        n15145), .ZN(n15070) );
  OAI221_X1 U16606 ( .B1(n15107), .B2(keyinput_f56), .C1(n15145), .C2(
        keyinput_f2), .A(n15070), .ZN(n15074) );
  XOR2_X1 U16607 ( .A(SI_1_), .B(keyinput_f31), .Z(n15072) );
  XNOR2_X1 U16608 ( .A(SI_2_), .B(keyinput_f30), .ZN(n15071) );
  NAND2_X1 U16609 ( .A1(n15072), .A2(n15071), .ZN(n15073) );
  NOR4_X1 U16610 ( .A1(n15076), .A2(n15075), .A3(n15074), .A4(n15073), .ZN(
        n15101) );
  AOI22_X1 U16611 ( .A1(n15078), .A2(keyinput_f36), .B1(keyinput_f19), .B2(
        n15144), .ZN(n15077) );
  OAI221_X1 U16612 ( .B1(n15078), .B2(keyinput_f36), .C1(n15144), .C2(
        keyinput_f19), .A(n15077), .ZN(n15087) );
  XNOR2_X1 U16613 ( .A(P3_REG3_REG_14__SCAN_IN), .B(keyinput_f37), .ZN(n15082)
         );
  XNOR2_X1 U16614 ( .A(SI_3_), .B(keyinput_f29), .ZN(n15081) );
  XNOR2_X1 U16615 ( .A(SI_5_), .B(keyinput_f27), .ZN(n15080) );
  XNOR2_X1 U16616 ( .A(SI_9_), .B(keyinput_f23), .ZN(n15079) );
  NAND4_X1 U16617 ( .A1(n15082), .A2(n15081), .A3(n15080), .A4(n15079), .ZN(
        n15086) );
  XNOR2_X1 U16618 ( .A(keyinput_f58), .B(n15083), .ZN(n15085) );
  XNOR2_X1 U16619 ( .A(keyinput_f40), .B(n8365), .ZN(n15084) );
  NOR4_X1 U16620 ( .A1(n15087), .A2(n15086), .A3(n15085), .A4(n15084), .ZN(
        n15100) );
  AOI22_X1 U16621 ( .A1(n15152), .A2(keyinput_f33), .B1(n6678), .B2(
        keyinput_f61), .ZN(n15088) );
  OAI221_X1 U16622 ( .B1(n15152), .B2(keyinput_f33), .C1(n6678), .C2(
        keyinput_f61), .A(n15088), .ZN(n15098) );
  AOI22_X1 U16623 ( .A1(n15090), .A2(keyinput_f12), .B1(n6680), .B2(
        keyinput_f43), .ZN(n15089) );
  OAI221_X1 U16624 ( .B1(n15090), .B2(keyinput_f12), .C1(n6680), .C2(
        keyinput_f43), .A(n15089), .ZN(n15097) );
  INV_X1 U16625 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n15109) );
  AOI22_X1 U16626 ( .A1(n15109), .A2(keyinput_f42), .B1(keyinput_f6), .B2(
        n15171), .ZN(n15091) );
  OAI221_X1 U16627 ( .B1(n15109), .B2(keyinput_f42), .C1(n15171), .C2(
        keyinput_f6), .A(n15091), .ZN(n15096) );
  AOI22_X1 U16628 ( .A1(n15094), .A2(keyinput_f16), .B1(n15093), .B2(
        keyinput_f62), .ZN(n15092) );
  OAI221_X1 U16629 ( .B1(n15094), .B2(keyinput_f16), .C1(n15093), .C2(
        keyinput_f62), .A(n15092), .ZN(n15095) );
  NOR4_X1 U16630 ( .A1(n15098), .A2(n15097), .A3(n15096), .A4(n15095), .ZN(
        n15099) );
  NAND4_X1 U16631 ( .A1(n15102), .A2(n15101), .A3(n15100), .A4(n15099), .ZN(
        n15103) );
  OAI22_X1 U16632 ( .A1(keyinput_f21), .A2(n15202), .B1(n15104), .B2(n15103), 
        .ZN(n15105) );
  AOI21_X1 U16633 ( .B1(keyinput_f21), .B2(n15202), .A(n15105), .ZN(n15201) );
  AOI22_X1 U16634 ( .A1(n6678), .A2(keyinput_g61), .B1(n15107), .B2(
        keyinput_g56), .ZN(n15106) );
  OAI221_X1 U16635 ( .B1(n6678), .B2(keyinput_g61), .C1(n15107), .C2(
        keyinput_g56), .A(n15106), .ZN(n15118) );
  AOI22_X1 U16636 ( .A1(n7155), .A2(keyinput_g8), .B1(n15109), .B2(
        keyinput_g42), .ZN(n15108) );
  OAI221_X1 U16637 ( .B1(n7155), .B2(keyinput_g8), .C1(n15109), .C2(
        keyinput_g42), .A(n15108), .ZN(n15117) );
  AOI22_X1 U16638 ( .A1(n15112), .A2(keyinput_g1), .B1(n15111), .B2(
        keyinput_g46), .ZN(n15110) );
  OAI221_X1 U16639 ( .B1(n15112), .B2(keyinput_g1), .C1(n15111), .C2(
        keyinput_g46), .A(n15110), .ZN(n15116) );
  XNOR2_X1 U16640 ( .A(SI_1_), .B(keyinput_g31), .ZN(n15114) );
  XNOR2_X1 U16641 ( .A(SI_10_), .B(keyinput_g22), .ZN(n15113) );
  NAND2_X1 U16642 ( .A1(n15114), .A2(n15113), .ZN(n15115) );
  NOR4_X1 U16643 ( .A1(n15118), .A2(n15117), .A3(n15116), .A4(n15115), .ZN(
        n15160) );
  INV_X1 U16644 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n15120) );
  AOI22_X1 U16645 ( .A1(n6680), .A2(keyinput_g43), .B1(n15120), .B2(
        keyinput_g60), .ZN(n15119) );
  OAI221_X1 U16646 ( .B1(n6680), .B2(keyinput_g43), .C1(n15120), .C2(
        keyinput_g60), .A(n15119), .ZN(n15130) );
  AOI22_X1 U16647 ( .A1(SI_27_), .A2(keyinput_g5), .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .ZN(n15121) );
  OAI221_X1 U16648 ( .B1(SI_27_), .B2(keyinput_g5), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput_g57), .A(n15121), .ZN(n15129)
         );
  INV_X1 U16649 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n15123) );
  AOI22_X1 U16650 ( .A1(n15124), .A2(keyinput_g11), .B1(n15123), .B2(
        keyinput_g51), .ZN(n15122) );
  OAI221_X1 U16651 ( .B1(n15124), .B2(keyinput_g11), .C1(n15123), .C2(
        keyinput_g51), .A(n15122), .ZN(n15128) );
  AOI22_X1 U16652 ( .A1(n8370), .A2(keyinput_g53), .B1(keyinput_g14), .B2(
        n15126), .ZN(n15125) );
  OAI221_X1 U16653 ( .B1(n8370), .B2(keyinput_g53), .C1(n15126), .C2(
        keyinput_g14), .A(n15125), .ZN(n15127) );
  NOR4_X1 U16654 ( .A1(n15130), .A2(n15129), .A3(n15128), .A4(n15127), .ZN(
        n15159) );
  AOI22_X1 U16655 ( .A1(n10877), .A2(keyinput_g44), .B1(n15132), .B2(
        keyinput_g38), .ZN(n15131) );
  OAI221_X1 U16656 ( .B1(n10877), .B2(keyinput_g44), .C1(n15132), .C2(
        keyinput_g38), .A(n15131), .ZN(n15142) );
  AOI22_X1 U16657 ( .A1(P3_U3151), .A2(keyinput_g34), .B1(keyinput_g39), .B2(
        n15134), .ZN(n15133) );
  OAI221_X1 U16658 ( .B1(P3_U3151), .B2(keyinput_g34), .C1(n15134), .C2(
        keyinput_g39), .A(n15133), .ZN(n15141) );
  AOI22_X1 U16659 ( .A1(n7301), .A2(keyinput_g18), .B1(n15136), .B2(
        keyinput_g50), .ZN(n15135) );
  OAI221_X1 U16660 ( .B1(n7301), .B2(keyinput_g18), .C1(n15136), .C2(
        keyinput_g50), .A(n15135), .ZN(n15140) );
  XNOR2_X1 U16661 ( .A(SI_5_), .B(keyinput_g27), .ZN(n15138) );
  XNOR2_X1 U16662 ( .A(SI_16_), .B(keyinput_g16), .ZN(n15137) );
  NAND2_X1 U16663 ( .A1(n15138), .A2(n15137), .ZN(n15139) );
  NOR4_X1 U16664 ( .A1(n15142), .A2(n15141), .A3(n15140), .A4(n15139), .ZN(
        n15158) );
  AOI22_X1 U16665 ( .A1(n15145), .A2(keyinput_g2), .B1(n15144), .B2(
        keyinput_g19), .ZN(n15143) );
  OAI221_X1 U16666 ( .B1(n15145), .B2(keyinput_g2), .C1(n15144), .C2(
        keyinput_g19), .A(n15143), .ZN(n15156) );
  AOI22_X1 U16667 ( .A1(n8379), .A2(keyinput_g47), .B1(keyinput_g54), .B2(
        n10716), .ZN(n15146) );
  OAI221_X1 U16668 ( .B1(n8379), .B2(keyinput_g47), .C1(n10716), .C2(
        keyinput_g54), .A(n15146), .ZN(n15155) );
  INV_X1 U16669 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n15148) );
  AOI22_X1 U16670 ( .A1(n15149), .A2(keyinput_g35), .B1(n15148), .B2(
        keyinput_g45), .ZN(n15147) );
  OAI221_X1 U16671 ( .B1(n15149), .B2(keyinput_g35), .C1(n15148), .C2(
        keyinput_g45), .A(n15147), .ZN(n15154) );
  AOI22_X1 U16672 ( .A1(n15152), .A2(keyinput_g33), .B1(n15151), .B2(
        keyinput_g37), .ZN(n15150) );
  OAI221_X1 U16673 ( .B1(n15152), .B2(keyinput_g33), .C1(n15151), .C2(
        keyinput_g37), .A(n15150), .ZN(n15153) );
  NOR4_X1 U16674 ( .A1(n15156), .A2(n15155), .A3(n15154), .A4(n15153), .ZN(
        n15157) );
  NAND4_X1 U16675 ( .A1(n15160), .A2(n15159), .A3(n15158), .A4(n15157), .ZN(
        n15199) );
  AOI22_X1 U16676 ( .A1(SI_6_), .A2(keyinput_g26), .B1(SI_19_), .B2(
        keyinput_g13), .ZN(n15161) );
  OAI221_X1 U16677 ( .B1(SI_6_), .B2(keyinput_g26), .C1(SI_19_), .C2(
        keyinput_g13), .A(n15161), .ZN(n15168) );
  AOI22_X1 U16678 ( .A1(SI_9_), .A2(keyinput_g23), .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .ZN(n15162) );
  OAI221_X1 U16679 ( .B1(SI_9_), .B2(keyinput_g23), .C1(
        P3_REG3_REG_27__SCAN_IN), .C2(keyinput_g36), .A(n15162), .ZN(n15167)
         );
  AOI22_X1 U16680 ( .A1(SI_12_), .A2(keyinput_g20), .B1(SI_22_), .B2(
        keyinput_g10), .ZN(n15163) );
  OAI221_X1 U16681 ( .B1(SI_12_), .B2(keyinput_g20), .C1(SI_22_), .C2(
        keyinput_g10), .A(n15163), .ZN(n15166) );
  AOI22_X1 U16682 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(SI_4_), 
        .B2(keyinput_g28), .ZN(n15164) );
  OAI221_X1 U16683 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(SI_4_), .C2(keyinput_g28), .A(n15164), .ZN(n15165) );
  NOR4_X1 U16684 ( .A1(n15168), .A2(n15167), .A3(n15166), .A4(n15165), .ZN(
        n15197) );
  XOR2_X1 U16685 ( .A(n15169), .B(keyinput_g7), .Z(n15177) );
  AOI22_X1 U16686 ( .A1(SI_20_), .A2(keyinput_g12), .B1(n15171), .B2(
        keyinput_g6), .ZN(n15170) );
  OAI221_X1 U16687 ( .B1(SI_20_), .B2(keyinput_g12), .C1(n15171), .C2(
        keyinput_g6), .A(n15170), .ZN(n15176) );
  AOI22_X1 U16688 ( .A1(SI_2_), .A2(keyinput_g30), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(keyinput_g40), .ZN(n15172) );
  OAI221_X1 U16689 ( .B1(SI_2_), .B2(keyinput_g30), .C1(P3_REG3_REG_3__SCAN_IN), .C2(keyinput_g40), .A(n15172), .ZN(n15175) );
  AOI22_X1 U16690 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        P3_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .ZN(n15173) );
  OAI221_X1 U16691 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        P3_REG3_REG_20__SCAN_IN), .C2(keyinput_g55), .A(n15173), .ZN(n15174)
         );
  NOR4_X1 U16692 ( .A1(n15177), .A2(n15176), .A3(n15175), .A4(n15174), .ZN(
        n15196) );
  AOI22_X1 U16693 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(keyinput_g48), .B1(
        P3_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n15178) );
  OAI221_X1 U16694 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .C1(
        P3_REG3_REG_19__SCAN_IN), .C2(keyinput_g41), .A(n15178), .ZN(n15185)
         );
  AOI22_X1 U16695 ( .A1(SI_17_), .A2(keyinput_g15), .B1(SI_28_), .B2(
        keyinput_g4), .ZN(n15179) );
  OAI221_X1 U16696 ( .B1(SI_17_), .B2(keyinput_g15), .C1(SI_28_), .C2(
        keyinput_g4), .A(n15179), .ZN(n15184) );
  AOI22_X1 U16697 ( .A1(SI_15_), .A2(keyinput_g17), .B1(
        P3_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .ZN(n15180) );
  OAI221_X1 U16698 ( .B1(SI_15_), .B2(keyinput_g17), .C1(
        P3_REG3_REG_11__SCAN_IN), .C2(keyinput_g58), .A(n15180), .ZN(n15183)
         );
  AOI22_X1 U16699 ( .A1(SI_0_), .A2(keyinput_g32), .B1(SI_29_), .B2(
        keyinput_g3), .ZN(n15181) );
  OAI221_X1 U16700 ( .B1(SI_0_), .B2(keyinput_g32), .C1(SI_29_), .C2(
        keyinput_g3), .A(n15181), .ZN(n15182) );
  NOR4_X1 U16701 ( .A1(n15185), .A2(n15184), .A3(n15183), .A4(n15182), .ZN(
        n15195) );
  AOI22_X1 U16702 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(keyinput_g63), .B1(
        P3_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .ZN(n15186) );
  OAI221_X1 U16703 ( .B1(P3_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput_g62), .A(n15186), .ZN(n15193)
         );
  AOI22_X1 U16704 ( .A1(SI_8_), .A2(keyinput_g24), .B1(SI_23_), .B2(
        keyinput_g9), .ZN(n15187) );
  OAI221_X1 U16705 ( .B1(SI_8_), .B2(keyinput_g24), .C1(SI_23_), .C2(
        keyinput_g9), .A(n15187), .ZN(n15192) );
  AOI22_X1 U16706 ( .A1(SI_7_), .A2(keyinput_g25), .B1(P3_REG3_REG_4__SCAN_IN), 
        .B2(keyinput_g52), .ZN(n15188) );
  OAI221_X1 U16707 ( .B1(SI_7_), .B2(keyinput_g25), .C1(P3_REG3_REG_4__SCAN_IN), .C2(keyinput_g52), .A(n15188), .ZN(n15191) );
  AOI22_X1 U16708 ( .A1(SI_3_), .A2(keyinput_g29), .B1(P3_REG3_REG_5__SCAN_IN), 
        .B2(keyinput_g49), .ZN(n15189) );
  OAI221_X1 U16709 ( .B1(SI_3_), .B2(keyinput_g29), .C1(P3_REG3_REG_5__SCAN_IN), .C2(keyinput_g49), .A(n15189), .ZN(n15190) );
  NOR4_X1 U16710 ( .A1(n15193), .A2(n15192), .A3(n15191), .A4(n15190), .ZN(
        n15194) );
  NAND4_X1 U16711 ( .A1(n15197), .A2(n15196), .A3(n15195), .A4(n15194), .ZN(
        n15198) );
  OAI22_X1 U16712 ( .A1(keyinput_g21), .A2(n15202), .B1(n15199), .B2(n15198), 
        .ZN(n15200) );
  AOI211_X1 U16713 ( .C1(keyinput_g21), .C2(n15202), .A(n15201), .B(n15200), 
        .ZN(n15205) );
  XNOR2_X1 U16714 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n15203) );
  XNOR2_X1 U16715 ( .A(n15203), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n15204) );
  NOR2_X1 U16716 ( .A1(P3_ADDR_REG_18__SCAN_IN), .A2(n15207), .ZN(n15208) );
  OAI22_X1 U16717 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n15210), .B1(n15209), 
        .B2(n15208), .ZN(n15211) );
  XOR2_X1 U16718 ( .A(n15213), .B(n15212), .Z(SUB_1596_U59) );
  XNOR2_X1 U16719 ( .A(n15214), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16720 ( .B1(n15216), .B2(n15215), .A(n15225), .ZN(SUB_1596_U53) );
  XNOR2_X1 U16721 ( .A(n15218), .B(n15217), .ZN(SUB_1596_U56) );
  OAI21_X1 U16722 ( .B1(n15221), .B2(n15220), .A(n15219), .ZN(n15223) );
  XOR2_X1 U16723 ( .A(n15223), .B(n15222), .Z(SUB_1596_U60) );
  XOR2_X1 U16724 ( .A(n15225), .B(n15224), .Z(SUB_1596_U5) );
  NAND2_X1 U7279 ( .A1(n8214), .A2(n11228), .ZN(n10178) );
  CLKBUF_X1 U7220 ( .A(n7557), .Z(n8211) );
  CLKBUF_X1 U7453 ( .A(n9350), .Z(n9351) );
  CLKBUF_X1 U9106 ( .A(n10254), .Z(n6653) );
endmodule

