

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4373, n4374, n4376, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10240;

  NAND2_X1 U4878 ( .A1(n8490), .A2(n8491), .ZN(n8489) );
  INV_X1 U4879 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n10240) );
  CLKBUF_X2 U4880 ( .A(n5240), .Z(n5569) );
  INV_X1 U4881 ( .A(n5200), .ZN(n6304) );
  BUF_X2 U4882 ( .A(n6356), .Z(n8925) );
  INV_X1 U4883 ( .A(n5638), .ZN(n8615) );
  CLKBUF_X1 U4884 ( .A(n6722), .Z(n6723) );
  CLKBUF_X2 U4885 ( .A(n6280), .Z(n7703) );
  NAND2_X1 U4886 ( .A1(n5605), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5606) );
  NAND2_X2 U4887 ( .A1(n6177), .A2(n7883), .ZN(n6737) );
  NOR3_X1 U4888 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .A3(
        P2_IR_REG_6__SCAN_IN), .ZN(n5144) );
  INV_X1 U4889 ( .A(n10240), .ZN(n4373) );
  INV_X1 U4890 ( .A(n4373), .ZN(n4374) );
  INV_X1 U4891 ( .A(n4373), .ZN(P2_U3152) );
  NAND2_X1 U4892 ( .A1(n8489), .A2(n5022), .ZN(n8466) );
  CLKBUF_X2 U4893 ( .A(n6226), .Z(n8918) );
  NAND2_X1 U4894 ( .A1(n7533), .A2(n5639), .ZN(n4399) );
  INV_X1 U4896 ( .A(n4504), .ZN(n5819) );
  OR2_X1 U4897 ( .A1(n5650), .A2(n8024), .ZN(n6402) );
  OR2_X1 U4898 ( .A1(n9524), .A2(n4854), .ZN(n4853) );
  INV_X2 U4899 ( .A(n6476), .ZN(n7748) );
  NAND2_X1 U4900 ( .A1(n8318), .A2(n5804), .ZN(n5806) );
  OAI21_X2 U4901 ( .B1(n5689), .B2(n8179), .A(n6402), .ZN(n4504) );
  AOI211_X1 U4902 ( .C1(n4491), .C2(n8296), .A(n8294), .B(n8260), .ZN(n5811)
         );
  NAND2_X1 U4903 ( .A1(n7114), .A2(n7113), .ZN(n7112) );
  INV_X1 U4904 ( .A(n8023), .ZN(n8232) );
  INV_X1 U4905 ( .A(n5205), .ZN(n5206) );
  AND3_X1 U4906 ( .A1(n5217), .A2(n5216), .A3(n5215), .ZN(n10105) );
  NOR2_X1 U4907 ( .A1(n5607), .A2(n4715), .ZN(n5658) );
  INV_X2 U4908 ( .A(n8922), .ZN(n6247) );
  NAND2_X1 U4909 ( .A1(n5571), .A2(n5570), .ZN(n8654) );
  NAND2_X1 U4910 ( .A1(n5728), .A2(n5727), .ZN(n7021) );
  INV_X1 U4911 ( .A(n5323), .ZN(n6186) );
  CLKBUF_X2 U4912 ( .A(n6250), .Z(n7279) );
  NAND2_X1 U4913 ( .A1(n7631), .A2(n7630), .ZN(n9631) );
  NAND2_X1 U4914 ( .A1(n7607), .A2(n7606), .ZN(n9640) );
  AOI22_X1 U4915 ( .A1(n9599), .A2(n10005), .B1(n10004), .B2(n9598), .ZN(n9600) );
  INV_X2 U4916 ( .A(n6401), .ZN(n8646) );
  AOI211_X1 U4917 ( .C1(n9599), .C2(n9909), .A(n7733), .B(n7732), .ZN(n7734)
         );
  OR2_X1 U4918 ( .A1(n4399), .A2(n10059), .ZN(n4376) );
  INV_X1 U4920 ( .A(n4504), .ZN(n4378) );
  NAND2_X1 U4921 ( .A1(n6628), .A2(n7743), .ZN(n6813) );
  XNOR2_X2 U4922 ( .A(n6095), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6099) );
  NOR2_X2 U4923 ( .A1(n6445), .A2(n4478), .ZN(n5946) );
  OAI21_X2 U4924 ( .B1(n7517), .B2(n7516), .A(n5780), .ZN(n7548) );
  XNOR2_X1 U4925 ( .A(n10105), .B(n4504), .ZN(n5697) );
  NAND2_X1 U4926 ( .A1(n5178), .A2(n8763), .ZN(n4379) );
  NAND2_X1 U4927 ( .A1(n5178), .A2(n8763), .ZN(n4380) );
  OAI21_X2 U4928 ( .B1(n5360), .B2(n5091), .A(n5090), .ZN(n5385) );
  OAI21_X2 U4929 ( .B1(n5344), .B2(n5076), .A(n5075), .ZN(n5360) );
  NAND2_X1 U4930 ( .A1(n6304), .A2(n8023), .ZN(n5691) );
  NAND2_X4 U4931 ( .A1(n6099), .A2(n9696), .ZN(n7679) );
  AOI21_X2 U4933 ( .B1(n8503), .B2(n4491), .A(n8499), .ZN(n8481) );
  OR2_X1 U4934 ( .A1(n8931), .A2(n4595), .ZN(n4594) );
  NOR2_X1 U4935 ( .A1(n8915), .A2(n8914), .ZN(n8931) );
  NAND2_X2 U4936 ( .A1(n9017), .A2(n9014), .ZN(n8909) );
  INV_X1 U4937 ( .A(n8607), .ZN(n4381) );
  NAND2_X1 U4938 ( .A1(n5014), .A2(n5621), .ZN(n6760) );
  AND2_X1 U4939 ( .A1(n7091), .A2(n7094), .ZN(n7153) );
  NAND2_X1 U4940 ( .A1(n4388), .A2(n4384), .ZN(n6585) );
  NAND2_X1 U4941 ( .A1(n4386), .A2(n4388), .ZN(n6767) );
  AND2_X1 U4942 ( .A1(n5648), .A2(n4384), .ZN(n4386) );
  NAND4_X2 U4943 ( .A1(n5210), .A2(n5209), .A3(n5208), .A4(n5207), .ZN(n10064)
         );
  INV_X1 U4944 ( .A(n6865), .ZN(n9982) );
  NAND2_X2 U4945 ( .A1(n8218), .A2(n8615), .ZN(n8224) );
  INV_X1 U4946 ( .A(n6433), .ZN(n4384) );
  INV_X2 U4948 ( .A(n5203), .ZN(n5599) );
  INV_X1 U4949 ( .A(n6349), .ZN(n7700) );
  INV_X2 U4950 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  AND2_X1 U4951 ( .A1(n9605), .A2(n4838), .ZN(n4837) );
  NAND2_X1 U4952 ( .A1(n4497), .A2(n4433), .ZN(n7848) );
  NAND2_X1 U4953 ( .A1(n8899), .A2(n8898), .ZN(n8981) );
  NAND2_X1 U4954 ( .A1(n8853), .A2(n8857), .ZN(n8980) );
  AOI21_X1 U4955 ( .B1(n7727), .B2(n9916), .A(n7726), .ZN(n9601) );
  AND2_X1 U4956 ( .A1(n4518), .A2(n4517), .ZN(n9761) );
  OR2_X1 U4957 ( .A1(n9757), .A2(n10155), .ZN(n4518) );
  OAI21_X1 U4958 ( .B1(n4687), .B2(n4689), .A(n7831), .ZN(n4686) );
  OR2_X1 U4959 ( .A1(n9476), .A2(n7850), .ZN(n4884) );
  NAND2_X1 U4960 ( .A1(n8808), .A2(n8807), .ZN(n9014) );
  NOR2_X2 U4961 ( .A1(n8432), .A2(n8240), .ZN(n8424) );
  AND2_X1 U4962 ( .A1(n4943), .A2(n4939), .ZN(n7838) );
  NAND2_X1 U4963 ( .A1(n4798), .A2(n4492), .ZN(n8490) );
  NAND2_X1 U4964 ( .A1(n5597), .A2(n5596), .ZN(n8240) );
  NAND2_X1 U4965 ( .A1(n7698), .A2(n7697), .ZN(n9598) );
  NOR2_X1 U4966 ( .A1(n8486), .A2(n8661), .ZN(n4389) );
  NAND2_X1 U4967 ( .A1(n8485), .A2(n4747), .ZN(n8486) );
  XNOR2_X1 U4968 ( .A(n5595), .B(n5594), .ZN(n8760) );
  NAND2_X1 U4969 ( .A1(n8888), .A2(n8890), .ZN(n4603) );
  NOR2_X2 U4970 ( .A1(n8518), .A2(n8669), .ZN(n8485) );
  INV_X1 U4971 ( .A(n8339), .ZN(n8661) );
  NAND2_X1 U4972 ( .A1(n4493), .A2(n7676), .ZN(n9609) );
  NAND2_X2 U4973 ( .A1(n7665), .A2(n7664), .ZN(n9614) );
  XNOR2_X1 U4974 ( .A(n7562), .B(n7554), .ZN(n8010) );
  NAND2_X1 U4975 ( .A1(n7651), .A2(n7747), .ZN(n7653) );
  NAND2_X1 U4976 ( .A1(n8559), .A2(n8544), .ZN(n8531) );
  XNOR2_X1 U4977 ( .A(n5559), .B(n5558), .ZN(n7663) );
  XNOR2_X1 U4978 ( .A(n5545), .B(n5544), .ZN(n7651) );
  XNOR2_X1 U4979 ( .A(n5531), .B(n5528), .ZN(n7642) );
  NAND2_X1 U4980 ( .A1(n4381), .A2(n8592), .ZN(n4413) );
  NAND2_X1 U4981 ( .A1(n5517), .A2(n5141), .ZN(n5531) );
  OAI21_X1 U4982 ( .B1(n7189), .B2(n9785), .A(n7776), .ZN(n7324) );
  OAI21_X1 U4983 ( .B1(n5503), .B2(n5502), .A(n5136), .ZN(n5515) );
  NAND2_X1 U4984 ( .A1(n5471), .A2(n5470), .ZN(n8698) );
  NOR2_X2 U4985 ( .A1(n7451), .A2(n8718), .ZN(n8634) );
  OR2_X2 U4986 ( .A1(n7468), .A2(n8723), .ZN(n7451) );
  NAND2_X1 U4987 ( .A1(n4489), .A2(n4488), .ZN(n6961) );
  AND2_X1 U4988 ( .A1(n5620), .A2(n8028), .ZN(n5014) );
  NAND2_X1 U4989 ( .A1(n4514), .A2(n4513), .ZN(n6845) );
  INV_X1 U4990 ( .A(n6767), .ZN(n4514) );
  INV_X1 U4991 ( .A(n6585), .ZN(n4387) );
  CLKBUF_X1 U4992 ( .A(n8237), .Z(n8314) );
  XNOR2_X1 U4993 ( .A(n5344), .B(n5343), .ZN(n7033) );
  INV_X2 U4994 ( .A(n9926), .ZN(n4382) );
  INV_X1 U4995 ( .A(n6460), .ZN(n4388) );
  INV_X1 U4996 ( .A(n10073), .ZN(n5647) );
  AND4_X1 U4997 ( .A1(n5254), .A2(n5253), .A3(n5252), .A4(n5251), .ZN(n6762)
         );
  BUF_X2 U4998 ( .A(n6356), .Z(n8919) );
  INV_X1 U4999 ( .A(n10116), .ZN(n4383) );
  INV_X1 U5000 ( .A(n4505), .ZN(n10096) );
  AND4_X1 U5001 ( .A1(n5184), .A2(n5183), .A3(n5182), .A4(n5181), .ZN(n5200)
         );
  INV_X2 U5002 ( .A(n4503), .ZN(n8015) );
  NAND4_X1 U5003 ( .A1(n6284), .A2(n6283), .A3(n6282), .A4(n6281), .ZN(n6866)
         );
  NAND3_X1 U5004 ( .A1(n4646), .A2(n6104), .A3(n6106), .ZN(n8942) );
  NAND4_X1 U5005 ( .A1(n6372), .A2(n6371), .A3(n6370), .A4(n6369), .ZN(n9068)
         );
  AND2_X1 U5006 ( .A1(n4390), .A2(n4376), .ZN(n4505) );
  OR2_X1 U5007 ( .A1(n4395), .A2(n6073), .ZN(n4485) );
  NAND2_X1 U5008 ( .A1(n4398), .A2(n7743), .ZN(n4395) );
  CLKBUF_X1 U5009 ( .A(n6172), .Z(n7719) );
  NAND2_X1 U5010 ( .A1(n4613), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4612) );
  NAND2_X1 U5011 ( .A1(n7533), .A2(n5639), .ZN(n4398) );
  INV_X1 U5012 ( .A(n6250), .ZN(n6628) );
  INV_X1 U5013 ( .A(n6099), .ZN(n7563) );
  NAND2_X1 U5014 ( .A1(n5465), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5467) );
  INV_X1 U5015 ( .A(n6101), .ZN(n9696) );
  OR2_X1 U5016 ( .A1(n8755), .A2(n5657), .ZN(n5172) );
  NAND2_X1 U5017 ( .A1(n5664), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4392) );
  OR2_X1 U5018 ( .A1(n5170), .A2(n5657), .ZN(n4391) );
  AOI21_X1 U5019 ( .B1(n5438), .B2(P2_IR_REG_31__SCAN_IN), .A(n4537), .ZN(
        n4536) );
  INV_X1 U5020 ( .A(n4538), .ZN(n4537) );
  AOI21_X1 U5021 ( .B1(n4403), .B2(P2_IR_REG_31__SCAN_IN), .A(
        P2_IR_REG_18__SCAN_IN), .ZN(n4538) );
  NAND2_X1 U5022 ( .A1(n5150), .A2(n5024), .ZN(n5607) );
  AND2_X1 U5023 ( .A1(n5011), .A2(n5871), .ZN(n4889) );
  INV_X2 U5024 ( .A(n7077), .ZN(n4385) );
  OR2_X1 U5025 ( .A1(n5345), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5349) );
  NOR2_X1 U5026 ( .A1(n4401), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n5011) );
  NAND2_X1 U5027 ( .A1(n5187), .A2(n5188), .ZN(n6072) );
  NOR2_X1 U5028 ( .A1(n5873), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4572) );
  AND4_X1 U5029 ( .A1(n5386), .A2(n5146), .A3(n5366), .A4(n5145), .ZN(n5148)
         );
  INV_X1 U5030 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6436) );
  INV_X1 U5031 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4772) );
  INV_X1 U5032 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5025) );
  NOR2_X1 U5033 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4574) );
  INV_X1 U5034 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5366) );
  NOR2_X2 U5035 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5186) );
  OR2_X1 U5036 ( .A1(n6430), .A2(n4387), .ZN(n10112) );
  XNOR2_X1 U5037 ( .A(n6585), .B(n4383), .ZN(n10117) );
  NOR2_X4 U5038 ( .A1(n8473), .A2(n8654), .ZN(n8450) );
  INV_X1 U5039 ( .A(n4389), .ZN(n8473) );
  NAND3_X1 U5040 ( .A1(n4435), .A2(n4485), .A3(n5192), .ZN(n6296) );
  NAND4_X1 U5041 ( .A1(n4435), .A2(n4485), .A3(n4505), .A4(n5192), .ZN(n10073)
         );
  NAND2_X1 U5042 ( .A1(n4399), .A2(n8764), .ZN(n4390) );
  XNOR2_X2 U5043 ( .A(n4391), .B(n5169), .ZN(n5639) );
  XNOR2_X2 U5044 ( .A(n4392), .B(n5154), .ZN(n7533) );
  AND2_X2 U5045 ( .A1(n8634), .A2(n8640), .ZN(n8635) );
  NAND2_X1 U5046 ( .A1(n7346), .A2(n7474), .ZN(n7468) );
  AND2_X2 U5047 ( .A1(n8580), .A2(n8564), .ZN(n8559) );
  NOR2_X2 U5048 ( .A1(n4413), .A2(n8698), .ZN(n8580) );
  AND2_X2 U5049 ( .A1(n7153), .A2(n7207), .ZN(n4477) );
  NOR2_X2 U5050 ( .A1(n6845), .A2(n7008), .ZN(n7091) );
  NOR2_X4 U5051 ( .A1(n6944), .A2(n10003), .ZN(n6943) );
  INV_X1 U5053 ( .A(n5819), .ZN(n5816) );
  NOR2_X4 U5054 ( .A1(n4414), .A2(n9619), .ZN(n9178) );
  OR2_X2 U5055 ( .A1(n9193), .A2(n9201), .ZN(n4414) );
  NOR2_X4 U5056 ( .A1(n9148), .A2(n9603), .ZN(n9141) );
  NOR2_X2 U5057 ( .A1(n9163), .A2(n9609), .ZN(n4512) );
  NAND2_X1 U5058 ( .A1(n4398), .A2(n4498), .ZN(n4396) );
  NAND2_X1 U5059 ( .A1(n4399), .A2(n7743), .ZN(n4397) );
  NAND2_X1 U5060 ( .A1(n4398), .A2(n7743), .ZN(n5240) );
  NOR2_X2 U5061 ( .A1(n5917), .A2(n5853), .ZN(n5866) );
  CLKBUF_X2 U5062 ( .A(n6721), .Z(n8940) );
  NOR2_X1 U5063 ( .A1(n6750), .A2(n6721), .ZN(n6751) );
  NAND2_X1 U5064 ( .A1(n7533), .A2(n5639), .ZN(n6031) );
  NAND2_X2 U5065 ( .A1(n6408), .A2(n8604), .ZN(n6401) );
  NAND2_X1 U5066 ( .A1(n9171), .A2(n7826), .ZN(n4680) );
  NOR2_X1 U5067 ( .A1(n4758), .A2(n8566), .ZN(n4757) );
  INV_X1 U5068 ( .A(n4760), .ZN(n4758) );
  NAND2_X1 U5069 ( .A1(n8844), .A2(n4590), .ZN(n4588) );
  NAND2_X1 U5070 ( .A1(n5579), .A2(n5578), .ZN(n7562) );
  INV_X1 U5071 ( .A(n5343), .ZN(n5076) );
  INV_X1 U5072 ( .A(n8456), .ZN(n4739) );
  NAND2_X1 U5073 ( .A1(n4853), .A2(n4850), .ZN(n9491) );
  AOI21_X1 U5074 ( .B1(n4855), .B2(n4852), .A(n4851), .ZN(n4850) );
  INV_X1 U5075 ( .A(n4858), .ZN(n4852) );
  INV_X2 U5076 ( .A(n6813), .ZN(n7747) );
  NAND2_X1 U5077 ( .A1(n8076), .A2(n8065), .ZN(n4534) );
  NAND2_X1 U5078 ( .A1(n4421), .A2(n4673), .ZN(n4669) );
  NAND2_X1 U5079 ( .A1(n4468), .A2(n7779), .ZN(n4673) );
  AOI21_X1 U5080 ( .B1(n4539), .B2(n8150), .A(n8149), .ZN(n8156) );
  NAND2_X1 U5081 ( .A1(n4541), .A2(n4540), .ZN(n4539) );
  NOR2_X1 U5082 ( .A1(n8146), .A2(n4405), .ZN(n4540) );
  AND2_X1 U5083 ( .A1(n8430), .A2(n8164), .ZN(n4522) );
  NAND2_X1 U5084 ( .A1(n8827), .A2(n8828), .ZN(n8838) );
  OAI21_X1 U5085 ( .B1(n4691), .B2(n4695), .A(n4694), .ZN(n4690) );
  INV_X1 U5086 ( .A(n4680), .ZN(n4695) );
  NOR2_X1 U5087 ( .A1(n5761), .A2(n7218), .ZN(n4976) );
  OR2_X1 U5088 ( .A1(n7214), .A2(n7218), .ZN(n7355) );
  OR2_X1 U5089 ( .A1(n8418), .A2(n8020), .ZN(n8174) );
  AND2_X1 U5090 ( .A1(n8339), .A2(n8458), .ZN(n8152) );
  AND2_X1 U5091 ( .A1(n8661), .A2(n8254), .ZN(n5636) );
  AND2_X1 U5092 ( .A1(n8505), .A2(n5634), .ZN(n4801) );
  NOR2_X1 U5093 ( .A1(n8669), .A2(n4491), .ZN(n5635) );
  NOR2_X1 U5094 ( .A1(n8687), .A2(n8568), .ZN(n4750) );
  OR2_X1 U5095 ( .A1(n8709), .A2(n8623), .ZN(n8119) );
  AOI21_X1 U5096 ( .B1(n4794), .B2(n4793), .A(n4792), .ZN(n4791) );
  AND2_X1 U5097 ( .A1(n8109), .A2(n8108), .ZN(n4794) );
  NAND2_X1 U5098 ( .A1(n7563), .A2(n9696), .ZN(n6172) );
  AOI21_X1 U5099 ( .B1(n4883), .B2(n7850), .A(n4448), .ZN(n4882) );
  INV_X1 U5100 ( .A(n7808), .ZN(n4561) );
  NAND2_X1 U5101 ( .A1(n6926), .A2(n4843), .ZN(n7764) );
  NAND2_X1 U5102 ( .A1(n6726), .A2(n6725), .ZN(n9903) );
  OR2_X1 U5103 ( .A1(n7738), .A2(n9295), .ZN(n7742) );
  NAND2_X1 U5104 ( .A1(n5567), .A2(n5566), .ZN(n5579) );
  OAI21_X1 U5105 ( .B1(n5434), .B2(n5113), .A(n5112), .ZN(n5451) );
  NOR2_X1 U5106 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n4576) );
  NOR2_X1 U5107 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4575) );
  NAND2_X1 U5108 ( .A1(n4912), .A2(n4910), .ZN(n5344) );
  AOI21_X1 U5109 ( .B1(n4914), .B2(n4916), .A(n4911), .ZN(n4910) );
  INV_X1 U5110 ( .A(n5072), .ZN(n4911) );
  NAND2_X1 U5111 ( .A1(n5029), .A2(n6169), .ZN(n5031) );
  NAND2_X1 U5112 ( .A1(n6251), .A2(n4445), .ZN(n5029) );
  AND2_X1 U5113 ( .A1(n5638), .A2(n8228), .ZN(n8179) );
  NAND2_X1 U5114 ( .A1(n8219), .A2(n8218), .ZN(n4549) );
  OAI21_X1 U5115 ( .B1(n4957), .B2(n8406), .A(n4956), .ZN(n8388) );
  NAND2_X1 U5116 ( .A1(n4957), .A2(n8406), .ZN(n4956) );
  AND2_X1 U5117 ( .A1(n8444), .A2(n5637), .ZN(n8012) );
  OR2_X1 U5118 ( .A1(n8649), .A2(n8255), .ZN(n5637) );
  AOI21_X1 U5119 ( .B1(n4737), .B2(n4736), .A(n4743), .ZN(n4735) );
  INV_X1 U5120 ( .A(n4746), .ZN(n4736) );
  NAND2_X1 U5121 ( .A1(n8339), .A2(n8254), .ZN(n4744) );
  XNOR2_X1 U5122 ( .A(n8654), .B(n8341), .ZN(n8456) );
  OR2_X1 U5123 ( .A1(n8692), .A2(n8553), .ZN(n8139) );
  AOI21_X1 U5124 ( .B1(n4757), .B2(n4755), .A(n4457), .ZN(n4754) );
  INV_X1 U5125 ( .A(n4761), .ZN(n4755) );
  NAND2_X1 U5126 ( .A1(n8629), .A2(n4440), .ZN(n8601) );
  OAI21_X1 U5127 ( .B1(n7342), .B2(n8085), .A(n8089), .ZN(n7476) );
  INV_X1 U5128 ( .A(n5569), .ZN(n5469) );
  INV_X1 U5129 ( .A(n6031), .ZN(n5468) );
  INV_X1 U5130 ( .A(n4731), .ZN(n5604) );
  NAND2_X1 U5131 ( .A1(n8924), .A2(n8942), .ZN(n4579) );
  NAND2_X1 U5132 ( .A1(n4593), .A2(n4583), .ZN(n4582) );
  INV_X1 U5133 ( .A(n4586), .ZN(n4583) );
  NAND2_X1 U5134 ( .A1(n6101), .A2(n7563), .ZN(n6280) );
  NOR2_X1 U5135 ( .A1(n6322), .A2(n6323), .ZN(n6321) );
  XNOR2_X1 U5136 ( .A(n4635), .B(n4634), .ZN(n9123) );
  INV_X1 U5137 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n4634) );
  NOR2_X1 U5138 ( .A1(n9118), .A2(n4636), .ZN(n4635) );
  AND2_X1 U5139 ( .A1(n9119), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4636) );
  XNOR2_X1 U5140 ( .A(n9614), .B(n9056), .ZN(n9171) );
  AOI21_X1 U5141 ( .B1(n9537), .B2(n7592), .A(n7591), .ZN(n9524) );
  AND2_X1 U5142 ( .A1(n9651), .A2(n9569), .ZN(n7591) );
  INV_X1 U5143 ( .A(n4862), .ZN(n9575) );
  AOI21_X1 U5144 ( .B1(n4868), .B2(n7565), .A(n4874), .ZN(n4863) );
  NAND2_X1 U5145 ( .A1(n4865), .A2(n7565), .ZN(n4864) );
  OR2_X1 U5146 ( .A1(n9669), .A2(n8967), .ZN(n7709) );
  NAND2_X1 U5147 ( .A1(n7135), .A2(n7032), .ZN(n7189) );
  OR2_X1 U5148 ( .A1(n6904), .A2(n6854), .ZN(n6855) );
  NAND2_X1 U5149 ( .A1(n8010), .A2(n7747), .ZN(n7686) );
  AND2_X1 U5150 ( .A1(n4840), .A2(n4475), .ZN(n9606) );
  NAND2_X1 U5151 ( .A1(n4842), .A2(n4841), .ZN(n4840) );
  NAND2_X1 U5152 ( .A1(n8001), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6095) );
  XNOR2_X1 U5153 ( .A(n6097), .B(P1_IR_REG_29__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U5154 ( .A1(n6096), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U5155 ( .A1(n5568), .A2(n5579), .ZN(n7675) );
  OR2_X1 U5156 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  OAI21_X1 U5157 ( .B1(n8412), .B2(n8411), .A(n4963), .ZN(n4962) );
  AOI21_X1 U5158 ( .B1(n8413), .B2(n10050), .A(n10053), .ZN(n4963) );
  NAND2_X1 U5159 ( .A1(n4598), .A2(n9026), .ZN(n8915) );
  NAND2_X1 U5160 ( .A1(n4600), .A2(n4599), .ZN(n4598) );
  INV_X1 U5161 ( .A(n9028), .ZN(n4599) );
  NOR2_X1 U5162 ( .A1(n8064), .A2(n8173), .ZN(n4533) );
  NAND2_X1 U5163 ( .A1(n4535), .A2(n8062), .ZN(n8076) );
  NAND2_X1 U5164 ( .A1(n8057), .A2(n8056), .ZN(n4535) );
  NOR2_X1 U5165 ( .A1(n4678), .A2(n4677), .ZN(n4676) );
  AOI21_X1 U5166 ( .B1(n4527), .B2(n8135), .A(n8126), .ZN(n4526) );
  INV_X1 U5167 ( .A(n4529), .ZN(n4527) );
  AOI21_X1 U5168 ( .B1(n8124), .B2(n4530), .A(n8118), .ZN(n4529) );
  INV_X1 U5169 ( .A(n4667), .ZN(n4666) );
  OAI21_X1 U5170 ( .B1(n4668), .B2(n4421), .A(n4674), .ZN(n4667) );
  NAND2_X1 U5171 ( .A1(n7782), .A2(n4699), .ZN(n4674) );
  OAI211_X1 U5172 ( .C1(n8130), .C2(n8173), .A(n8145), .B(n4450), .ZN(n4541)
         );
  AOI21_X1 U5173 ( .B1(n4819), .B2(n4400), .A(n4818), .ZN(n4817) );
  INV_X1 U5174 ( .A(n4455), .ZN(n4818) );
  AOI21_X1 U5175 ( .B1(n8160), .B2(n8159), .A(n8158), .ZN(n4523) );
  NAND2_X1 U5176 ( .A1(n7251), .A2(n7232), .ZN(n8073) );
  NOR2_X1 U5177 ( .A1(n8974), .A2(n5002), .ZN(n5000) );
  NAND2_X1 U5178 ( .A1(n4688), .A2(n4437), .ZN(n4687) );
  NAND2_X1 U5179 ( .A1(n4689), .A2(n4691), .ZN(n4688) );
  OR2_X1 U5180 ( .A1(n7945), .A2(n7911), .ZN(n7954) );
  INV_X1 U5181 ( .A(n7854), .ZN(n7972) );
  INV_X1 U5182 ( .A(n7893), .ZN(n4831) );
  INV_X1 U5183 ( .A(n6892), .ZN(n4698) );
  NOR2_X1 U5184 ( .A1(n4479), .A2(n4909), .ZN(n4908) );
  INV_X1 U5185 ( .A(n5578), .ZN(n4909) );
  OR2_X1 U5186 ( .A1(n4479), .A2(n7561), .ZN(n4906) );
  INV_X1 U5187 ( .A(n7739), .ZN(n4905) );
  NOR2_X1 U5188 ( .A1(n4901), .A2(n4905), .ZN(n4898) );
  NAND2_X1 U5189 ( .A1(n4903), .A2(n4901), .ZN(n4900) );
  AOI21_X1 U5190 ( .B1(n4925), .B2(n4923), .A(n4922), .ZN(n4921) );
  INV_X1 U5191 ( .A(n5558), .ZN(n4922) );
  INV_X1 U5192 ( .A(n4927), .ZN(n4923) );
  INV_X1 U5193 ( .A(n4925), .ZN(n4924) );
  INV_X1 U5194 ( .A(n5065), .ZN(n4916) );
  NOR2_X1 U5195 ( .A1(n4969), .A2(n5815), .ZN(n4968) );
  INV_X1 U5196 ( .A(n4974), .ZN(n4969) );
  OR2_X1 U5197 ( .A1(n7229), .A2(n5743), .ZN(n4506) );
  OR2_X1 U5198 ( .A1(n8681), .A2(n8554), .ZN(n8131) );
  AND2_X1 U5199 ( .A1(n4756), .A2(n4428), .ZN(n4751) );
  NOR2_X1 U5200 ( .A1(n8551), .A2(n4781), .ZN(n4780) );
  INV_X1 U5201 ( .A(n8139), .ZN(n4781) );
  INV_X1 U5202 ( .A(n4729), .ZN(n4721) );
  NAND2_X1 U5203 ( .A1(n4730), .A2(n8103), .ZN(n4729) );
  INV_X1 U5204 ( .A(n5245), .ZN(n4703) );
  INV_X1 U5205 ( .A(n4800), .ZN(n4798) );
  OR2_X1 U5206 ( .A1(n4803), .A2(n4799), .ZN(n4492) );
  OAI21_X1 U5207 ( .B1(n4803), .B2(n8206), .A(n8150), .ZN(n4800) );
  AND2_X1 U5208 ( .A1(n8133), .A2(n8125), .ZN(n8576) );
  NOR2_X1 U5209 ( .A1(n8114), .A2(n4796), .ZN(n4795) );
  NAND2_X1 U5210 ( .A1(n7018), .A2(n8024), .ZN(n5690) );
  NAND2_X1 U5211 ( .A1(n5151), .A2(n5608), .ZN(n4715) );
  AND2_X1 U5212 ( .A1(n5153), .A2(n4990), .ZN(n4989) );
  INV_X1 U5213 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4990) );
  NOR2_X1 U5214 ( .A1(n5004), .A2(n5003), .ZN(n5002) );
  INV_X1 U5215 ( .A(n8965), .ZN(n5003) );
  INV_X1 U5216 ( .A(n8964), .ZN(n5004) );
  OR2_X1 U5217 ( .A1(n8840), .A2(n8839), .ZN(n8846) );
  INV_X1 U5218 ( .A(n4693), .ZN(n4692) );
  OAI21_X1 U5219 ( .B1(n7833), .B2(n7834), .A(n7955), .ZN(n4693) );
  AOI21_X1 U5220 ( .B1(n4661), .B2(n7814), .A(n4658), .ZN(n7817) );
  NOR2_X1 U5221 ( .A1(n4660), .A2(n4659), .ZN(n4658) );
  NOR2_X1 U5222 ( .A1(n5947), .A2(n6971), .ZN(n9069) );
  NOR2_X1 U5223 ( .A1(n9137), .A2(n9136), .ZN(n9135) );
  OR2_X1 U5224 ( .A1(n9598), .A2(n9134), .ZN(n7944) );
  OR2_X1 U5225 ( .A1(n9609), .A2(n9031), .ZN(n7948) );
  NAND2_X1 U5226 ( .A1(n7674), .A2(n4888), .ZN(n4886) );
  AND2_X1 U5227 ( .A1(n4887), .A2(n4879), .ZN(n4878) );
  AND2_X1 U5228 ( .A1(n4426), .A2(n9185), .ZN(n4887) );
  NAND2_X1 U5229 ( .A1(n4882), .A2(n4880), .ZN(n4879) );
  INV_X1 U5230 ( .A(n4883), .ZN(n4880) );
  INV_X1 U5231 ( .A(n4882), .ZN(n4881) );
  INV_X1 U5232 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4820) );
  OR2_X1 U5233 ( .A1(n9634), .A2(n9519), .ZN(n7813) );
  OR2_X1 U5234 ( .A1(n9634), .A2(n9479), .ZN(n7809) );
  AND2_X1 U5235 ( .A1(n9640), .A2(n9532), .ZN(n7618) );
  OR2_X1 U5236 ( .A1(n7270), .A2(n7046), .ZN(n7891) );
  INV_X1 U5237 ( .A(n6886), .ZN(n4846) );
  INV_X1 U5238 ( .A(n6934), .ZN(n4848) );
  NAND2_X1 U5239 ( .A1(n4890), .A2(n5011), .ZN(n5894) );
  NAND2_X1 U5240 ( .A1(n4889), .A2(n4890), .ZN(n6096) );
  NOR2_X1 U5241 ( .A1(n5544), .A2(n4928), .ZN(n4927) );
  INV_X1 U5242 ( .A(n5530), .ZN(n4928) );
  AOI21_X1 U5243 ( .B1(n4929), .B2(n4927), .A(n4926), .ZN(n4925) );
  INV_X1 U5244 ( .A(n5543), .ZN(n4926) );
  INV_X1 U5245 ( .A(n5528), .ZN(n4929) );
  NOR2_X1 U5246 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n6142) );
  INV_X1 U5247 ( .A(n5919), .ZN(n4614) );
  INV_X1 U5248 ( .A(n5384), .ZN(n5093) );
  XNOR2_X1 U5249 ( .A(n5073), .B(SI_11_), .ZN(n5343) );
  OAI21_X1 U5250 ( .B1(n5275), .B2(n4896), .A(n5289), .ZN(n4895) );
  INV_X1 U5251 ( .A(n5051), .ZN(n4896) );
  NAND2_X1 U5252 ( .A1(n9799), .A2(n4772), .ZN(n4770) );
  OR3_X1 U5253 ( .A1(n5552), .A2(n8287), .A3(n8333), .ZN(n5573) );
  OR2_X1 U5254 ( .A1(n4976), .A2(n4978), .ZN(n4975) );
  INV_X1 U5255 ( .A(n7362), .ZN(n4978) );
  INV_X1 U5256 ( .A(n4976), .ZN(n7357) );
  OR2_X1 U5257 ( .A1(n8304), .A2(n4986), .ZN(n4985) );
  INV_X1 U5258 ( .A(n5792), .ZN(n4986) );
  INV_X1 U5259 ( .A(n4985), .ZN(n4982) );
  OR2_X1 U5260 ( .A1(n5520), .A2(n5166), .ZN(n5522) );
  AOI21_X1 U5261 ( .B1(n7021), .B2(n7020), .A(n5732), .ZN(n7114) );
  AND2_X1 U5262 ( .A1(n5745), .A2(n5744), .ZN(n7218) );
  OR2_X1 U5263 ( .A1(n8283), .A2(n8282), .ZN(n4974) );
  OR2_X1 U5264 ( .A1(n8172), .A2(n8171), .ZN(n8177) );
  AND4_X1 U5265 ( .A1(n5429), .A2(n5428), .A3(n5427), .A4(n5426), .ZN(n8613)
         );
  AND4_X1 U5266 ( .A1(n5236), .A2(n5235), .A3(n5234), .A4(n5233), .ZN(n6550)
         );
  NAND2_X1 U5267 ( .A1(n5206), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U5268 ( .A1(n7510), .A2(n5980), .ZN(n8382) );
  OR2_X1 U5269 ( .A1(n8382), .A2(n8381), .ZN(n4946) );
  NAND2_X1 U5270 ( .A1(n8424), .A2(n8425), .ZN(n8423) );
  INV_X1 U5271 ( .A(n5636), .ZN(n8159) );
  NAND2_X1 U5272 ( .A1(n8466), .A2(n4806), .ZN(n8455) );
  AND2_X1 U5273 ( .A1(n4741), .A2(n5557), .ZN(n4740) );
  NAND2_X1 U5274 ( .A1(n8491), .A2(n4746), .ZN(n4741) );
  AND2_X1 U5275 ( .A1(n5551), .A2(n5550), .ZN(n8339) );
  OR2_X1 U5276 ( .A1(n8666), .A2(n8330), .ZN(n8468) );
  NAND2_X1 U5277 ( .A1(n4747), .A2(n8330), .ZN(n4746) );
  NOR2_X1 U5278 ( .A1(n8152), .A2(n5636), .ZN(n8467) );
  NAND2_X1 U5279 ( .A1(n4802), .A2(n4801), .ZN(n8504) );
  INV_X1 U5280 ( .A(n8514), .ZN(n4802) );
  NOR2_X2 U5281 ( .A1(n5635), .A2(n8146), .ZN(n8505) );
  NOR2_X1 U5282 ( .A1(n8681), .A2(n5512), .ZN(n5513) );
  NOR2_X1 U5283 ( .A1(n8515), .A2(n8524), .ZN(n8514) );
  NAND2_X1 U5284 ( .A1(n4782), .A2(n4779), .ZN(n8535) );
  AND2_X1 U5285 ( .A1(n8536), .A2(n8142), .ZN(n4779) );
  AND2_X1 U5286 ( .A1(n8131), .A2(n8143), .ZN(n8536) );
  INV_X1 U5287 ( .A(n4757), .ZN(n4756) );
  OR2_X1 U5288 ( .A1(n4763), .A2(n4422), .ZN(n4760) );
  AND2_X1 U5289 ( .A1(n5479), .A2(n4431), .ZN(n4763) );
  NOR2_X1 U5290 ( .A1(n4422), .A2(n4762), .ZN(n4761) );
  INV_X1 U5291 ( .A(n5461), .ZN(n4762) );
  AOI21_X1 U5292 ( .B1(n4787), .B2(n4790), .A(n4784), .ZN(n4783) );
  INV_X1 U5293 ( .A(n8119), .ZN(n4784) );
  NAND2_X1 U5294 ( .A1(n8635), .A2(n5649), .ZN(n8607) );
  NAND2_X1 U5295 ( .A1(n8601), .A2(n5449), .ZN(n8587) );
  AND2_X1 U5296 ( .A1(n8119), .A2(n8120), .ZN(n8609) );
  NAND2_X1 U5297 ( .A1(n5431), .A2(n5430), .ZN(n8629) );
  AND2_X1 U5298 ( .A1(n7237), .A2(n4476), .ZN(n4726) );
  NAND2_X1 U5299 ( .A1(n4723), .A2(n4729), .ZN(n4728) );
  AND2_X1 U5300 ( .A1(n5383), .A2(n4717), .ZN(n4716) );
  NOR2_X1 U5301 ( .A1(n4727), .A2(n5629), .ZN(n4717) );
  OR2_X1 U5302 ( .A1(n7464), .A2(n5378), .ZN(n7434) );
  NAND2_X1 U5303 ( .A1(n4766), .A2(n4765), .ZN(n7342) );
  AOI21_X1 U5304 ( .B1(n5627), .B2(n5626), .A(n4767), .ZN(n4766) );
  INV_X1 U5305 ( .A(n8087), .ZN(n4767) );
  OR2_X1 U5306 ( .A1(n5312), .A2(n9328), .ZN(n5336) );
  OAI21_X1 U5307 ( .B1(n6836), .B2(n4418), .A(n4705), .ZN(n7238) );
  INV_X1 U5308 ( .A(n4706), .ZN(n4705) );
  OAI21_X1 U5309 ( .B1(n4709), .B2(n4418), .A(n5322), .ZN(n4706) );
  AND2_X1 U5310 ( .A1(n8067), .A2(n8069), .ZN(n7151) );
  NOR2_X1 U5311 ( .A1(n5310), .A2(n4710), .ZN(n4709) );
  INV_X1 U5312 ( .A(n5293), .ZN(n4710) );
  OR2_X1 U5313 ( .A1(n5295), .A2(n5294), .ZN(n5312) );
  OR2_X2 U5314 ( .A1(n10064), .A2(n10105), .ZN(n8044) );
  AND4_X1 U5315 ( .A1(n5224), .A2(n5223), .A3(n5222), .A4(n5221), .ZN(n6604)
         );
  NAND2_X1 U5316 ( .A1(n5421), .A2(n5420), .ZN(n8712) );
  INV_X1 U5317 ( .A(n5690), .ZN(n10097) );
  NAND2_X1 U5318 ( .A1(n4712), .A2(n4711), .ZN(n5173) );
  NOR2_X1 U5319 ( .A1(n4713), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4711) );
  OR2_X1 U5320 ( .A1(n5437), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n4403) );
  NOR2_X1 U5321 ( .A1(n6482), .A2(n4993), .ZN(n4992) );
  INV_X1 U5322 ( .A(n6347), .ZN(n4993) );
  NOR2_X1 U5323 ( .A1(n6497), .A2(n6496), .ZN(n6498) );
  INV_X1 U5324 ( .A(n6537), .ZN(n6496) );
  NAND2_X1 U5325 ( .A1(n8851), .A2(n8854), .ZN(n8899) );
  AOI22_X1 U5326 ( .A1(n4589), .A2(n4587), .B1(n4415), .B2(n4586), .ZN(n4585)
         );
  OAI21_X1 U5327 ( .B1(n4589), .B2(n4415), .A(n8909), .ZN(n4581) );
  INV_X1 U5328 ( .A(n5002), .ZN(n4997) );
  NAND2_X1 U5329 ( .A1(n4579), .A2(n4577), .ZN(n6249) );
  OR2_X1 U5330 ( .A1(n8845), .A2(n8846), .ZN(n8999) );
  NOR2_X1 U5331 ( .A1(n8957), .A2(n5008), .ZN(n5007) );
  INV_X1 U5332 ( .A(n5010), .ZN(n5008) );
  AND2_X1 U5333 ( .A1(n8889), .A2(n8782), .ZN(n4991) );
  NAND2_X1 U5334 ( .A1(n4603), .A2(n8889), .ZN(n8786) );
  OR2_X1 U5335 ( .A1(n7985), .A2(n7984), .ZN(n7987) );
  OR2_X1 U5336 ( .A1(n7679), .A2(n6748), .ZN(n6266) );
  OR2_X1 U5337 ( .A1(n6280), .A2(n6100), .ZN(n6105) );
  NOR2_X1 U5338 ( .A1(n9888), .A2(n9887), .ZN(n9886) );
  OR2_X1 U5339 ( .A1(n9886), .A2(n4633), .ZN(n4632) );
  AND2_X1 U5340 ( .A1(n9899), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4633) );
  AND2_X1 U5341 ( .A1(n4632), .A2(n4631), .ZN(n6195) );
  INV_X1 U5342 ( .A(n6196), .ZN(n4631) );
  OR2_X1 U5343 ( .A1(n6321), .A2(n4480), .ZN(n4629) );
  AND2_X1 U5344 ( .A1(n4629), .A2(n4628), .ZN(n6445) );
  INV_X1 U5345 ( .A(n6446), .ZN(n4628) );
  NOR2_X1 U5346 ( .A1(n5951), .A2(n9344), .ZN(n9070) );
  NAND2_X1 U5347 ( .A1(n4622), .A2(n4621), .ZN(n4620) );
  INV_X1 U5348 ( .A(n9073), .ZN(n4621) );
  OR2_X1 U5349 ( .A1(n9102), .A2(n4639), .ZN(n4638) );
  AND2_X1 U5350 ( .A1(n9109), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4639) );
  AND2_X1 U5351 ( .A1(n4638), .A2(n4637), .ZN(n9118) );
  INV_X1 U5352 ( .A(n9104), .ZN(n4637) );
  INV_X1 U5353 ( .A(n7877), .ZN(n7715) );
  NAND2_X1 U5354 ( .A1(n7944), .A2(n7979), .ZN(n7877) );
  NAND2_X1 U5355 ( .A1(n4564), .A2(n4563), .ZN(n9154) );
  AOI21_X1 U5356 ( .B1(n4569), .B2(n4834), .A(n4832), .ZN(n4563) );
  NAND2_X1 U5357 ( .A1(n7946), .A2(n9171), .ZN(n4835) );
  NAND2_X1 U5358 ( .A1(n9182), .A2(n9032), .ZN(n4888) );
  NAND2_X1 U5359 ( .A1(n4565), .A2(n4568), .ZN(n9184) );
  NOR2_X1 U5360 ( .A1(n9184), .A2(n9185), .ZN(n9183) );
  NAND2_X1 U5361 ( .A1(n4877), .A2(n4882), .ZN(n9177) );
  NAND2_X1 U5362 ( .A1(n9476), .A2(n4883), .ZN(n4877) );
  NAND2_X1 U5363 ( .A1(n4820), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n9437) );
  NAND2_X1 U5364 ( .A1(n7642), .A2(n7747), .ZN(n4499) );
  NOR2_X2 U5365 ( .A1(n9508), .A2(n9634), .ZN(n9494) );
  NOR2_X1 U5366 ( .A1(n7618), .A2(n4859), .ZN(n4858) );
  INV_X1 U5367 ( .A(n7604), .ZN(n4859) );
  NAND2_X1 U5368 ( .A1(n4857), .A2(n4856), .ZN(n4855) );
  INV_X1 U5369 ( .A(n7618), .ZN(n4856) );
  INV_X1 U5370 ( .A(n4860), .ZN(n4857) );
  AOI21_X1 U5371 ( .B1(n4560), .B2(n4558), .A(n9506), .ZN(n4557) );
  INV_X1 U5372 ( .A(n4560), .ZN(n4559) );
  INV_X1 U5373 ( .A(n4416), .ZN(n4558) );
  OAI21_X1 U5374 ( .B1(n4562), .B2(n7913), .A(n4561), .ZN(n4560) );
  INV_X1 U5375 ( .A(n9531), .ZN(n4562) );
  AND2_X1 U5376 ( .A1(n9506), .A2(n4432), .ZN(n4860) );
  AND2_X1 U5377 ( .A1(n9651), .A2(n8994), .ZN(n7913) );
  AND2_X1 U5378 ( .A1(n9559), .A2(n9553), .ZN(n9547) );
  OR2_X1 U5379 ( .A1(n9563), .A2(n9543), .ZN(n5018) );
  NOR2_X2 U5380 ( .A1(n9576), .A2(n9655), .ZN(n9559) );
  NOR2_X1 U5381 ( .A1(n7315), .A2(n9415), .ZN(n7423) );
  NAND2_X1 U5382 ( .A1(n7867), .A2(n4871), .ZN(n4870) );
  NAND2_X1 U5383 ( .A1(n4873), .A2(n4871), .ZN(n4869) );
  NAND2_X1 U5384 ( .A1(n9768), .A2(n9042), .ZN(n4871) );
  OR2_X1 U5385 ( .A1(n7396), .A2(n7389), .ZN(n7328) );
  AND2_X1 U5386 ( .A1(n7324), .A2(n7865), .ZN(n7326) );
  NAND2_X1 U5387 ( .A1(n7028), .A2(n7027), .ZN(n7030) );
  AND2_X1 U5388 ( .A1(n7891), .A2(n7887), .ZN(n7862) );
  NAND2_X1 U5389 ( .A1(n7905), .A2(n7764), .ZN(n7856) );
  NAND2_X1 U5390 ( .A1(n6938), .A2(n6935), .ZN(n6878) );
  NAND2_X1 U5391 ( .A1(n4649), .A2(n4647), .ZN(n6904) );
  INV_X1 U5392 ( .A(n4648), .ZN(n4647) );
  OAI21_X1 U5393 ( .B1(n6852), .B2(n4651), .A(n6868), .ZN(n4648) );
  AND2_X1 U5394 ( .A1(n8942), .A2(n6750), .ZN(n6800) );
  OR2_X1 U5395 ( .A1(n8942), .A2(n9929), .ZN(n6801) );
  AND2_X1 U5396 ( .A1(n9800), .A2(n7845), .ZN(n9911) );
  NAND2_X1 U5397 ( .A1(n4552), .A2(n6512), .ZN(n10003) );
  INV_X1 U5398 ( .A(n6511), .ZN(n4552) );
  XNOR2_X1 U5399 ( .A(n7746), .B(n7745), .ZN(n8016) );
  NAND2_X1 U5400 ( .A1(n6144), .A2(n5849), .ZN(n4613) );
  XNOR2_X1 U5401 ( .A(n5402), .B(n5403), .ZN(n7412) );
  XNOR2_X1 U5402 ( .A(n5365), .B(n5364), .ZN(n7278) );
  OR2_X1 U5403 ( .A1(n5360), .A2(n5359), .ZN(n5362) );
  BUF_X1 U5404 ( .A(n5917), .Z(n5919) );
  NAND2_X1 U5405 ( .A1(n4913), .A2(n5065), .ZN(n5329) );
  NAND2_X1 U5406 ( .A1(n5319), .A2(n5020), .ZN(n4913) );
  XNOR2_X1 U5407 ( .A(n5049), .B(SI_6_), .ZN(n5275) );
  NAND2_X1 U5408 ( .A1(n5048), .A2(n5047), .ZN(n5276) );
  INV_X1 U5409 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5848) );
  XNOR2_X1 U5410 ( .A(n5039), .B(SI_3_), .ZN(n5226) );
  NAND2_X1 U5411 ( .A1(n5033), .A2(n5032), .ZN(n5212) );
  CLKBUF_X1 U5412 ( .A(n6251), .Z(n4498) );
  NAND2_X1 U5413 ( .A1(n7675), .A2(n8015), .ZN(n5571) );
  NAND2_X1 U5414 ( .A1(n8010), .A2(n8015), .ZN(n5582) );
  NAND2_X1 U5415 ( .A1(n5495), .A2(n5494), .ZN(n8687) );
  NAND2_X1 U5416 ( .A1(n5483), .A2(n5482), .ZN(n8692) );
  NAND2_X1 U5417 ( .A1(n8328), .A2(n8329), .ZN(n4509) );
  NAND2_X1 U5418 ( .A1(n4972), .A2(n4973), .ZN(n8328) );
  NOR2_X1 U5419 ( .A1(n8329), .A2(n4971), .ZN(n4970) );
  INV_X1 U5420 ( .A(n4973), .ZN(n4971) );
  INV_X1 U5421 ( .A(n8308), .ZN(n8568) );
  AND4_X1 U5422 ( .A1(n5491), .A2(n5490), .A3(n5489), .A4(n5488), .ZN(n8553)
         );
  INV_X1 U5423 ( .A(n7118), .ZN(n8352) );
  INV_X1 U5424 ( .A(n6604), .ZN(n8357) );
  NAND2_X1 U5425 ( .A1(n7511), .A2(n7453), .ZN(n7510) );
  OAI21_X1 U5426 ( .B1(n8417), .B2(n5025), .A(n8416), .ZN(n4961) );
  INV_X1 U5427 ( .A(n4956), .ZN(n8403) );
  AOI21_X1 U5428 ( .B1(n4502), .B2(n10077), .A(n8245), .ZN(n4501) );
  INV_X1 U5429 ( .A(n8247), .ZN(n4502) );
  INV_X1 U5430 ( .A(n5644), .ZN(n5645) );
  AND2_X1 U5431 ( .A1(n5453), .A2(n5452), .ZN(n8592) );
  OR2_X1 U5432 ( .A1(n5467), .A2(n5466), .ZN(n4550) );
  INV_X1 U5433 ( .A(n8429), .ZN(n8644) );
  NAND2_X1 U5434 ( .A1(n6478), .A2(n6477), .ZN(n6926) );
  NAND2_X1 U5435 ( .A1(n4584), .A2(n4589), .ZN(n8856) );
  OR2_X1 U5436 ( .A1(n8933), .A2(n4596), .ZN(n4595) );
  NAND2_X1 U5437 ( .A1(n4597), .A2(n8982), .ZN(n4596) );
  INV_X1 U5438 ( .A(n8932), .ZN(n4597) );
  AND2_X1 U5439 ( .A1(n8917), .A2(n8916), .ZN(n8914) );
  INV_X1 U5440 ( .A(n8935), .ZN(n4602) );
  INV_X1 U5441 ( .A(n9058), .ZN(n8967) );
  NAND2_X1 U5442 ( .A1(n4593), .A2(n4592), .ZN(n4591) );
  NAND2_X1 U5443 ( .A1(n7595), .A2(n7594), .ZN(n9644) );
  INV_X1 U5444 ( .A(n9196), .ZN(n9032) );
  NAND2_X1 U5445 ( .A1(n7663), .A2(n7747), .ZN(n7665) );
  NAND4_X1 U5446 ( .A1(n6507), .A2(n6506), .A3(n6505), .A4(n6504), .ZN(n9067)
         );
  NAND3_X1 U5447 ( .A1(n6355), .A2(n6354), .A3(n6353), .ZN(n9912) );
  AND2_X1 U5448 ( .A1(n6352), .A2(n6351), .ZN(n6353) );
  NOR2_X1 U5449 ( .A1(n5898), .A2(n5899), .ZN(n5938) );
  NAND2_X1 U5450 ( .A1(n9120), .A2(n4429), .ZN(n4641) );
  OR2_X1 U5451 ( .A1(n9121), .A2(n9896), .ZN(n4642) );
  OAI21_X1 U5452 ( .B1(n9880), .B2(n4772), .A(n9126), .ZN(n4644) );
  NAND2_X1 U5453 ( .A1(n4839), .A2(n10034), .ZN(n4838) );
  NOR2_X1 U5454 ( .A1(n10229), .A2(n10228), .ZN(n10227) );
  NOR2_X1 U5455 ( .A1(n10226), .A2(n10225), .ZN(n10224) );
  NAND2_X1 U5456 ( .A1(n8066), .A2(n8173), .ZN(n4531) );
  NAND2_X1 U5457 ( .A1(n4534), .A2(n4533), .ZN(n4532) );
  INV_X1 U5458 ( .A(n8116), .ZN(n4530) );
  NAND2_X1 U5459 ( .A1(n4468), .A2(n4672), .ZN(n4671) );
  NAND2_X1 U5460 ( .A1(n4468), .A2(n7896), .ZN(n4670) );
  NOR2_X1 U5461 ( .A1(n4676), .A2(n4675), .ZN(n4672) );
  NOR2_X1 U5462 ( .A1(n7770), .A2(n7835), .ZN(n4654) );
  NAND2_X1 U5463 ( .A1(n4528), .A2(n8124), .ZN(n8136) );
  NAND2_X1 U5464 ( .A1(n4543), .A2(n8173), .ZN(n4542) );
  INV_X1 U5465 ( .A(n8131), .ZN(n4543) );
  NAND2_X1 U5466 ( .A1(n4525), .A2(n4524), .ZN(n8129) );
  AOI21_X1 U5467 ( .B1(n4526), .B2(n4410), .A(n4459), .ZN(n4524) );
  OAI21_X1 U5468 ( .B1(n7784), .B2(n4668), .A(n4666), .ZN(n7787) );
  NOR2_X1 U5469 ( .A1(n7750), .A2(n4936), .ZN(n4935) );
  OAI21_X1 U5470 ( .B1(n4680), .B2(n4679), .A(n7829), .ZN(n4691) );
  INV_X1 U5471 ( .A(n7827), .ZN(n4679) );
  NOR2_X1 U5472 ( .A1(n7806), .A2(n4699), .ZN(n4664) );
  INV_X1 U5473 ( .A(n4908), .ZN(n4901) );
  AOI21_X1 U5474 ( .B1(n4817), .B2(n4816), .A(n4481), .ZN(n4815) );
  NOR2_X1 U5475 ( .A1(n4816), .A2(n9759), .ZN(n4814) );
  INV_X1 U5476 ( .A(n4801), .ZN(n4803) );
  NAND2_X1 U5477 ( .A1(n4510), .A2(n8838), .ZN(n8833) );
  NAND2_X1 U5478 ( .A1(n4937), .A2(n4934), .ZN(n7751) );
  NAND2_X1 U5479 ( .A1(n4942), .A2(n4938), .ZN(n4937) );
  NAND2_X1 U5480 ( .A1(n7982), .A2(n4935), .ZN(n4934) );
  NOR2_X1 U5481 ( .A1(n7750), .A2(n4944), .ZN(n4938) );
  INV_X1 U5482 ( .A(n7812), .ZN(n4660) );
  INV_X1 U5483 ( .A(n7813), .ZN(n4659) );
  NAND2_X1 U5484 ( .A1(n4665), .A2(n4662), .ZN(n4661) );
  NOR2_X1 U5485 ( .A1(n4664), .A2(n4663), .ZN(n4662) );
  OAI21_X1 U5486 ( .B1(n7801), .B2(n7935), .A(n4699), .ZN(n4665) );
  NAND2_X1 U5487 ( .A1(n9517), .A2(n9531), .ZN(n4663) );
  NOR2_X1 U5488 ( .A1(n7596), .A2(n8993), .ZN(n7608) );
  OR2_X1 U5489 ( .A1(n5012), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4401) );
  INV_X1 U5490 ( .A(n5492), .ZN(n4933) );
  INV_X1 U5491 ( .A(n5127), .ZN(n4932) );
  INV_X1 U5492 ( .A(n4915), .ZN(n4914) );
  OAI21_X1 U5493 ( .B1(n5020), .B2(n4916), .A(n5019), .ZN(n4915) );
  NAND2_X1 U5494 ( .A1(n5069), .A2(n5068), .ZN(n5072) );
  OR2_X1 U5495 ( .A1(n4811), .A2(n8214), .ZN(n4809) );
  AOI22_X1 U5496 ( .A1(n4815), .A2(n4812), .B1(n4814), .B2(n4819), .ZN(n4811)
         );
  INV_X1 U5497 ( .A(n4817), .ZN(n4812) );
  NOR2_X1 U5498 ( .A1(n4815), .A2(n4814), .ZN(n4813) );
  AOI21_X1 U5499 ( .B1(n4521), .B2(n4409), .A(n4520), .ZN(n8171) );
  NAND2_X1 U5500 ( .A1(n8169), .A2(n4441), .ZN(n4520) );
  OAI21_X1 U5501 ( .B1(n4523), .B2(n8165), .A(n4522), .ZN(n4521) );
  NAND2_X1 U5502 ( .A1(n4959), .A2(n4958), .ZN(n4957) );
  NAND2_X1 U5503 ( .A1(n8393), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4958) );
  INV_X1 U5504 ( .A(n8387), .ZN(n4959) );
  AND2_X1 U5505 ( .A1(n4788), .A2(n8609), .ZN(n4787) );
  NAND2_X1 U5506 ( .A1(n4791), .A2(n4789), .ZN(n4788) );
  INV_X1 U5507 ( .A(n4795), .ZN(n4789) );
  INV_X1 U5508 ( .A(n4791), .ZN(n4790) );
  AND2_X1 U5509 ( .A1(n8084), .A2(n7378), .ZN(n5627) );
  NAND2_X1 U5510 ( .A1(n4516), .A2(n4515), .ZN(n7345) );
  INV_X1 U5511 ( .A(n7372), .ZN(n4516) );
  INV_X1 U5512 ( .A(n5309), .ZN(n4707) );
  NAND2_X1 U5513 ( .A1(n8357), .A2(n4384), .ZN(n8051) );
  NAND2_X1 U5514 ( .A1(n6304), .A2(n10075), .ZN(n5615) );
  INV_X1 U5515 ( .A(n4733), .ZN(n4732) );
  OAI21_X1 U5516 ( .B1(n4735), .B2(n8430), .A(n4452), .ZN(n4733) );
  NAND2_X1 U5517 ( .A1(n4737), .A2(n8439), .ZN(n4734) );
  NAND2_X1 U5518 ( .A1(n5638), .A2(n7018), .ZN(n8025) );
  AND2_X1 U5519 ( .A1(n5679), .A2(n5678), .ZN(n5682) );
  OAI22_X1 U5520 ( .A1(n8768), .A2(n8767), .B1(n8766), .B2(n8765), .ZN(n8778)
         );
  NAND2_X1 U5521 ( .A1(n8831), .A2(n4592), .ZN(n4587) );
  NAND2_X1 U5522 ( .A1(n8844), .A2(n4592), .ZN(n4586) );
  INV_X1 U5523 ( .A(n4999), .ZN(n4998) );
  OAI21_X1 U5524 ( .B1(n8974), .B2(n4402), .A(n8799), .ZN(n4999) );
  NAND2_X1 U5525 ( .A1(n7982), .A2(n8004), .ZN(n4939) );
  OR2_X1 U5526 ( .A1(n7954), .A2(n7930), .ZN(n7978) );
  NAND2_X1 U5527 ( .A1(n7737), .A2(n4940), .ZN(n7982) );
  NOR2_X1 U5528 ( .A1(n7880), .A2(n4941), .ZN(n4940) );
  INV_X1 U5529 ( .A(n7736), .ZN(n4941) );
  OR2_X1 U5530 ( .A1(n9603), .A2(n9156), .ZN(n7943) );
  OAI21_X1 U5531 ( .B1(n4835), .B2(n4833), .A(n7906), .ZN(n4832) );
  INV_X1 U5532 ( .A(n9185), .ZN(n4833) );
  INV_X1 U5533 ( .A(n4835), .ZN(n4834) );
  NOR2_X1 U5534 ( .A1(n9194), .A2(n4567), .ZN(n4566) );
  INV_X1 U5535 ( .A(n7815), .ZN(n4567) );
  NOR2_X1 U5536 ( .A1(n7650), .A2(n7851), .ZN(n4883) );
  NOR2_X1 U5537 ( .A1(n9625), .A2(n9481), .ZN(n7650) );
  INV_X1 U5538 ( .A(n4855), .ZN(n4854) );
  INV_X1 U5539 ( .A(n9500), .ZN(n4851) );
  INV_X1 U5540 ( .A(n7584), .ZN(n7585) );
  NAND2_X1 U5541 ( .A1(n7585), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n7596) );
  INV_X1 U5542 ( .A(n4870), .ZN(n4865) );
  NOR2_X1 U5543 ( .A1(n4823), .A2(n7865), .ZN(n4822) );
  INV_X1 U5544 ( .A(n4828), .ZN(n4823) );
  AND2_X1 U5545 ( .A1(n4831), .A2(n7306), .ZN(n4828) );
  NAND2_X1 U5546 ( .A1(n4458), .A2(n4831), .ZN(n4826) );
  NAND2_X1 U5547 ( .A1(n7866), .A2(n7306), .ZN(n4830) );
  OR2_X1 U5548 ( .A1(n6640), .A2(n6639), .ZN(n6823) );
  OR2_X1 U5549 ( .A1(n6919), .A2(n10020), .ZN(n7765) );
  NOR2_X1 U5550 ( .A1(n6502), .A2(n6468), .ZN(n6527) );
  NAND2_X1 U5551 ( .A1(n10003), .A2(n4551), .ZN(n7762) );
  INV_X1 U5552 ( .A(n9067), .ZN(n4551) );
  NAND2_X1 U5553 ( .A1(n4696), .A2(n6938), .ZN(n4700) );
  NOR2_X1 U5554 ( .A1(n6936), .A2(n4698), .ZN(n4697) );
  OR2_X1 U5555 ( .A1(n9912), .A2(n9989), .ZN(n6894) );
  INV_X1 U5556 ( .A(n6866), .ZN(n6853) );
  NAND2_X1 U5557 ( .A1(n6851), .A2(n6729), .ZN(n4650) );
  OAI22_X1 U5558 ( .A1(n7966), .A2(n6801), .B1(n9970), .B2(n6723), .ZN(n6851)
         );
  INV_X1 U5559 ( .A(n6096), .ZN(n4573) );
  INV_X1 U5560 ( .A(n9135), .ZN(n4842) );
  INV_X1 U5561 ( .A(n4487), .ZN(n7403) );
  NOR2_X1 U5562 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n5871) );
  NAND2_X1 U5563 ( .A1(n4907), .A2(n4906), .ZN(n7740) );
  NAND2_X1 U5564 ( .A1(n5579), .A2(n4908), .ZN(n4907) );
  OAI211_X1 U5565 ( .C1(n5579), .C2(n4904), .A(n4899), .B(n4897), .ZN(n7738)
         );
  AND2_X1 U5566 ( .A1(n4900), .A2(n4902), .ZN(n4899) );
  OR2_X1 U5567 ( .A1(n4906), .A2(n4905), .ZN(n4902) );
  AOI21_X1 U5568 ( .B1(n4921), .B2(n4924), .A(n4919), .ZN(n4918) );
  INV_X1 U5569 ( .A(n5560), .ZN(n4919) );
  AND2_X1 U5570 ( .A1(n5089), .A2(n5088), .ZN(n5090) );
  OR2_X1 U5571 ( .A1(n5359), .A2(n5363), .ZN(n5091) );
  OR2_X1 U5572 ( .A1(n5363), .A2(n5361), .ZN(n5088) );
  NAND2_X1 U5573 ( .A1(n5062), .A2(n5061), .ZN(n5065) );
  INV_X1 U5574 ( .A(SI_4_), .ZN(n9244) );
  NAND2_X1 U5575 ( .A1(n5035), .A2(SI_2_), .ZN(n5036) );
  AND2_X2 U5576 ( .A1(n4769), .A2(n4768), .ZN(n6251) );
  NAND3_X1 U5577 ( .A1(n4820), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4768) );
  NAND2_X1 U5578 ( .A1(n5814), .A2(n4967), .ZN(n4966) );
  INV_X1 U5579 ( .A(n4970), .ZN(n4967) );
  AND2_X1 U5580 ( .A1(n5722), .A2(n5721), .ZN(n4988) );
  NAND2_X1 U5581 ( .A1(n4456), .A2(n4506), .ZN(n7257) );
  INV_X1 U5582 ( .A(n4506), .ZN(n5753) );
  INV_X1 U5583 ( .A(n5522), .ZN(n5167) );
  NAND2_X1 U5584 ( .A1(n4987), .A2(n5791), .ZN(n8266) );
  INV_X1 U5585 ( .A(n8269), .ZN(n4987) );
  NAND2_X1 U5586 ( .A1(n8283), .A2(n8282), .ZN(n4973) );
  AND2_X1 U5587 ( .A1(n5017), .A2(n5738), .ZN(n4977) );
  AND4_X1 U5588 ( .A1(n5477), .A2(n5476), .A3(n5475), .A4(n5474), .ZN(n8311)
         );
  AND4_X1 U5589 ( .A1(n5328), .A2(n5327), .A3(n5326), .A4(n5325), .ZN(n7232)
         );
  AND4_X1 U5590 ( .A1(n5198), .A2(n5197), .A3(n5196), .A4(n5195), .ZN(n5614)
         );
  NAND2_X1 U5591 ( .A1(n5970), .A2(n4948), .ZN(n9734) );
  NAND2_X1 U5592 ( .A1(n6072), .A2(n4949), .ZN(n4948) );
  NOR2_X1 U5593 ( .A1(n9734), .A2(n4947), .ZN(n9733) );
  NAND2_X1 U5594 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n4947) );
  OR2_X1 U5595 ( .A1(n6694), .A2(n6693), .ZN(n4954) );
  AND2_X1 U5596 ( .A1(n6782), .A2(n4964), .ZN(n7101) );
  NAND2_X1 U5597 ( .A1(n6018), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4964) );
  NAND2_X1 U5598 ( .A1(n7101), .A2(n7100), .ZN(n7099) );
  AND2_X1 U5599 ( .A1(n4946), .A2(n4945), .ZN(n5988) );
  NAND2_X1 U5600 ( .A1(n8376), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4945) );
  AND2_X1 U5601 ( .A1(n8026), .A2(n4400), .ZN(n8211) );
  AOI21_X1 U5602 ( .B1(n4805), .B2(n4806), .A(n4447), .ZN(n4804) );
  INV_X1 U5603 ( .A(n5022), .ZN(n4805) );
  AND2_X1 U5604 ( .A1(n5598), .A2(n5584), .ZN(n8435) );
  NAND2_X1 U5605 ( .A1(n4752), .A2(n4749), .ZN(n8528) );
  AOI21_X1 U5606 ( .B1(n4751), .B2(n4754), .A(n4750), .ZN(n4749) );
  AND2_X1 U5607 ( .A1(n4754), .A2(n4428), .ZN(n4753) );
  OR2_X1 U5608 ( .A1(n5496), .A2(n9451), .ZN(n5520) );
  OR2_X1 U5609 ( .A1(n5442), .A2(n7518), .ZN(n5455) );
  NAND2_X1 U5610 ( .A1(n4720), .A2(n5413), .ZN(n4719) );
  NOR2_X1 U5611 ( .A1(n4723), .A2(n4727), .ZN(n4722) );
  OAI21_X1 U5612 ( .B1(n7447), .B2(n8109), .A(n8108), .ZN(n8621) );
  INV_X1 U5613 ( .A(n8101), .ZN(n8197) );
  NAND2_X1 U5614 ( .A1(n8096), .A2(n8095), .ZN(n8101) );
  AND2_X1 U5615 ( .A1(n7462), .A2(n8101), .ZN(n7464) );
  AND2_X1 U5616 ( .A1(n5382), .A2(n8196), .ZN(n7462) );
  AND4_X1 U5617 ( .A1(n5377), .A2(n5376), .A3(n5375), .A4(n5374), .ZN(n7440)
         );
  AND2_X1 U5618 ( .A1(n8088), .A2(n8089), .ZN(n8196) );
  NAND2_X1 U5619 ( .A1(n4477), .A2(n10147), .ZN(n7372) );
  AND4_X1 U5620 ( .A1(n5342), .A2(n5341), .A3(n5340), .A4(n5339), .ZN(n7344)
         );
  AND4_X1 U5621 ( .A1(n5317), .A2(n5316), .A3(n5315), .A4(n5314), .ZN(n7243)
         );
  NAND2_X1 U5622 ( .A1(n6836), .A2(n5293), .ZN(n7080) );
  AND4_X1 U5623 ( .A1(n5268), .A2(n5267), .A3(n5266), .A4(n5265), .ZN(n6841)
         );
  AND4_X1 U5624 ( .A1(n5300), .A2(n5299), .A3(n5298), .A4(n5297), .ZN(n7118)
         );
  NOR2_X1 U5625 ( .A1(n5261), .A2(n4703), .ZN(n4702) );
  INV_X1 U5626 ( .A(n6423), .ZN(n8184) );
  NAND2_X1 U5627 ( .A1(n8051), .A2(n6599), .ZN(n6423) );
  OR2_X1 U5628 ( .A1(n10155), .A2(n8615), .ZN(n5831) );
  NAND2_X1 U5629 ( .A1(n5505), .A2(n5504), .ZN(n8681) );
  NAND2_X1 U5630 ( .A1(n4786), .A2(n4791), .ZN(n8610) );
  NAND2_X1 U5631 ( .A1(n7447), .A2(n4795), .ZN(n4786) );
  AND2_X1 U5632 ( .A1(n5352), .A2(n5351), .ZN(n10154) );
  NAND2_X1 U5633 ( .A1(n4408), .A2(n4714), .ZN(n4713) );
  INV_X1 U5634 ( .A(n4715), .ZN(n4714) );
  NOR2_X1 U5635 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4980) );
  AOI21_X1 U5636 ( .B1(n4608), .B2(n4611), .A(n4606), .ZN(n4605) );
  INV_X1 U5637 ( .A(n6979), .ZN(n4606) );
  AND2_X1 U5638 ( .A1(n8814), .A2(n8815), .ZN(n8907) );
  NAND2_X1 U5639 ( .A1(n8979), .A2(n8867), .ZN(n5010) );
  NOR2_X1 U5640 ( .A1(n7632), .A2(n9414), .ZN(n7645) );
  INV_X1 U5641 ( .A(n4609), .ZN(n4608) );
  OAI22_X1 U5642 ( .A1(n4417), .A2(n4610), .B1(n6624), .B2(n6632), .ZN(n4609)
         );
  INV_X1 U5643 ( .A(n6810), .ZN(n4610) );
  NOR2_X1 U5644 ( .A1(n6810), .A2(n6633), .ZN(n4611) );
  INV_X1 U5645 ( .A(n8907), .ZN(n4592) );
  NAND2_X1 U5646 ( .A1(n6249), .A2(n6248), .ZN(n6262) );
  NAND2_X1 U5647 ( .A1(n8936), .A2(n8938), .ZN(n8937) );
  AND2_X1 U5648 ( .A1(n7492), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7574) );
  NAND2_X1 U5649 ( .A1(n4681), .A2(n4683), .ZN(n4497) );
  OR2_X1 U5650 ( .A1(n6280), .A2(n6171), .ZN(n6176) );
  NAND2_X1 U5651 ( .A1(n6350), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6174) );
  AOI21_X1 U5652 ( .B1(n6336), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6039), .ZN(
        n9842) );
  OR2_X1 U5653 ( .A1(n9070), .A2(n9071), .ZN(n4622) );
  AND2_X1 U5654 ( .A1(n4620), .A2(n4619), .ZN(n9090) );
  NAND2_X1 U5655 ( .A1(n9092), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4619) );
  NAND2_X1 U5656 ( .A1(n7737), .A2(n7736), .ZN(n9128) );
  NAND2_X1 U5657 ( .A1(n4876), .A2(n4875), .ZN(n9147) );
  AOI21_X1 U5658 ( .B1(n4878), .B2(n4881), .A(n4454), .ZN(n4875) );
  AOI21_X1 U5659 ( .B1(n9515), .B2(n7917), .A(n7711), .ZN(n9477) );
  AND2_X1 U5660 ( .A1(n9538), .A2(n7852), .ZN(n9539) );
  NAND3_X1 U5661 ( .A1(n9587), .A2(n9585), .A3(n9586), .ZN(n9584) );
  AND2_X1 U5662 ( .A1(n9564), .A2(n7793), .ZN(n9585) );
  OR2_X1 U5663 ( .A1(n7296), .A2(n7295), .ZN(n7315) );
  NAND2_X1 U5664 ( .A1(n4821), .A2(n4824), .ZN(n7422) );
  INV_X1 U5665 ( .A(n4825), .ZN(n4824) );
  NAND2_X1 U5666 ( .A1(n4822), .A2(n7193), .ZN(n4821) );
  OAI21_X1 U5667 ( .B1(n4826), .B2(n7865), .A(n7778), .ZN(n4825) );
  NAND2_X1 U5668 ( .A1(n4827), .A2(n4826), .ZN(n7395) );
  NAND2_X1 U5669 ( .A1(n7193), .A2(n4828), .ZN(n4827) );
  NAND2_X1 U5670 ( .A1(n7395), .A2(n7396), .ZN(n7394) );
  NOR2_X1 U5671 ( .A1(n6997), .A2(n6996), .ZN(n7037) );
  AND2_X1 U5672 ( .A1(n7779), .A2(n7890), .ZN(n7863) );
  NAND2_X1 U5673 ( .A1(n4829), .A2(n7306), .ZN(n7309) );
  OR2_X1 U5674 ( .A1(n7193), .A2(n7866), .ZN(n4829) );
  NAND2_X1 U5675 ( .A1(n7036), .A2(n7035), .ZN(n7777) );
  NAND2_X1 U5676 ( .A1(n7133), .A2(n7887), .ZN(n7193) );
  AOI21_X1 U5677 ( .B1(n7044), .B2(n7860), .A(n7770), .ZN(n7134) );
  NAND2_X1 U5678 ( .A1(n7134), .A2(n7862), .ZN(n7133) );
  INV_X1 U5679 ( .A(n9065), .ZN(n6919) );
  AND2_X1 U5680 ( .A1(n6885), .A2(n7856), .ZN(n4847) );
  NAND2_X1 U5681 ( .A1(n4845), .A2(n4434), .ZN(n4844) );
  INV_X1 U5682 ( .A(n6959), .ZN(n4489) );
  NAND2_X1 U5683 ( .A1(n6918), .A2(n7764), .ZN(n6953) );
  NAND2_X1 U5684 ( .A1(n4555), .A2(n4554), .ZN(n7974) );
  NAND2_X1 U5685 ( .A1(n7858), .A2(n7755), .ZN(n4554) );
  NAND2_X1 U5686 ( .A1(n7854), .A2(n6891), .ZN(n4555) );
  NAND2_X1 U5687 ( .A1(n7974), .A2(n6898), .ZN(n6918) );
  AND3_X1 U5688 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6503) );
  AND2_X1 U5689 ( .A1(n7762), .A2(n7755), .ZN(n7753) );
  INV_X1 U5690 ( .A(n6476), .ZN(n6475) );
  NAND2_X1 U5691 ( .A1(n6894), .A2(n6892), .ZN(n6905) );
  NAND2_X1 U5692 ( .A1(n6868), .A2(n6893), .ZN(n9915) );
  CLKBUF_X1 U5693 ( .A(n6797), .Z(n6798) );
  AND2_X1 U5694 ( .A1(n10005), .A2(n9203), .ZN(n6235) );
  NAND2_X1 U5695 ( .A1(n4884), .A2(n7849), .ZN(n9192) );
  NAND2_X1 U5696 ( .A1(n7573), .A2(n7572), .ZN(n9655) );
  INV_X1 U5697 ( .A(n6926), .ZN(n10015) );
  XNOR2_X1 U5698 ( .A(n7738), .B(SI_30_), .ZN(n8014) );
  NAND2_X1 U5699 ( .A1(n5593), .A2(n7558), .ZN(n5595) );
  NAND2_X1 U5700 ( .A1(n4920), .A2(n4925), .ZN(n5559) );
  NAND2_X1 U5701 ( .A1(n5531), .A2(n4927), .ZN(n4920) );
  OAI21_X1 U5702 ( .B1(n5531), .B2(n4929), .A(n5530), .ZN(n5545) );
  NAND4_X1 U5703 ( .A1(n5852), .A2(n5851), .A3(n6142), .A4(n5944), .ZN(n5853)
         );
  NOR2_X1 U5704 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5851) );
  INV_X1 U5705 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5868) );
  INV_X1 U5706 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9407) );
  INV_X1 U5707 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9405) );
  NAND2_X1 U5708 ( .A1(n4614), .A2(n4419), .ZN(n6141) );
  OR2_X1 U5709 ( .A1(n5931), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5933) );
  AOI21_X1 U5710 ( .B1(n4894), .B2(n4896), .A(n4453), .ZN(n4891) );
  NAND2_X1 U5711 ( .A1(n5059), .A2(n5058), .ZN(n5304) );
  XNOR2_X1 U5712 ( .A(n5045), .B(SI_5_), .ZN(n5256) );
  XNOR2_X1 U5713 ( .A(n5042), .B(n9244), .ZN(n5241) );
  XNOR2_X1 U5714 ( .A(n5034), .B(SI_2_), .ZN(n5211) );
  XNOR2_X1 U5715 ( .A(n5031), .B(n5030), .ZN(n5190) );
  XNOR2_X1 U5716 ( .A(n5889), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U5717 ( .A1(n9437), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U5718 ( .A1(n5025), .A2(n4770), .ZN(n5026) );
  NAND2_X1 U5719 ( .A1(n6711), .A2(n5721), .ZN(n6773) );
  INV_X1 U5720 ( .A(n4975), .ZN(n7358) );
  NAND2_X1 U5721 ( .A1(n7112), .A2(n5738), .ZN(n7356) );
  OAI22_X1 U5722 ( .A1(n10072), .A2(n8232), .B1(n10096), .B2(n4504), .ZN(n6294) );
  INV_X1 U5723 ( .A(n4984), .ZN(n4983) );
  OAI21_X1 U5724 ( .B1(n4985), .B2(n5791), .A(n5795), .ZN(n4984) );
  INV_X1 U5725 ( .A(n10154), .ZN(n7350) );
  AND4_X1 U5726 ( .A1(n5412), .A2(n5411), .A3(n5410), .A4(n5409), .ZN(n8625)
         );
  NAND2_X1 U5727 ( .A1(n6412), .A2(n5709), .ZN(n6549) );
  NAND2_X1 U5728 ( .A1(n5156), .A2(n5155), .ZN(n8669) );
  NAND2_X1 U5729 ( .A1(n8266), .A2(n5792), .ZN(n8305) );
  NAND2_X1 U5730 ( .A1(n5369), .A2(n5368), .ZN(n8728) );
  INV_X1 U5731 ( .A(n8592), .ZN(n8702) );
  AND4_X1 U5732 ( .A1(n5286), .A2(n5285), .A3(n5284), .A4(n5283), .ZN(n7081)
         );
  NAND2_X1 U5733 ( .A1(n5408), .A2(n5407), .ZN(n8718) );
  NAND2_X1 U5734 ( .A1(n4549), .A2(n8220), .ZN(n4548) );
  INV_X1 U5735 ( .A(n8230), .ZN(n4545) );
  INV_X1 U5736 ( .A(n7232), .ZN(n8350) );
  INV_X1 U5737 ( .A(n6550), .ZN(n8356) );
  NAND2_X1 U5738 ( .A1(n5599), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5210) );
  INV_X1 U5739 ( .A(n5614), .ZN(n10067) );
  INV_X1 U5740 ( .A(n6072), .ZN(n9738) );
  NOR2_X1 U5741 ( .A1(n6060), .A2(n4955), .ZN(n6694) );
  AND2_X1 U5742 ( .A1(n5998), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4955) );
  INV_X1 U5743 ( .A(n4954), .ZN(n6692) );
  NOR2_X1 U5744 ( .A1(n6658), .A2(n6657), .ZN(n6656) );
  AND2_X1 U5745 ( .A1(n4954), .A2(n4953), .ZN(n6658) );
  NAND2_X1 U5746 ( .A1(n6697), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4953) );
  NOR2_X1 U5747 ( .A1(n6670), .A2(n6669), .ZN(n6668) );
  NOR2_X1 U5748 ( .A1(n6704), .A2(n4952), .ZN(n6670) );
  AND2_X1 U5749 ( .A1(n6709), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4952) );
  NOR2_X1 U5750 ( .A1(n6668), .A2(n4950), .ZN(n6558) );
  NOR2_X1 U5751 ( .A1(n4951), .A2(n7248), .ZN(n4950) );
  INV_X1 U5752 ( .A(n6673), .ZN(n4951) );
  NAND2_X1 U5753 ( .A1(n6558), .A2(n6559), .ZN(n6557) );
  OR2_X1 U5754 ( .A1(n6781), .A2(n6780), .ZN(n6782) );
  INV_X1 U5755 ( .A(n4946), .ZN(n8380) );
  INV_X1 U5756 ( .A(n8388), .ZN(n8390) );
  NAND2_X1 U5757 ( .A1(n8018), .A2(n8017), .ZN(n8418) );
  AOI21_X1 U5758 ( .B1(n8649), .B2(n8434), .A(n8433), .ZN(n8650) );
  OAI21_X1 U5759 ( .B1(n8481), .B2(n4738), .A(n4735), .ZN(n8431) );
  AND2_X1 U5760 ( .A1(n8461), .A2(n8460), .ZN(n8657) );
  AND2_X1 U5761 ( .A1(n8466), .A2(n8159), .ZN(n8457) );
  AND2_X1 U5762 ( .A1(n4745), .A2(n4744), .ZN(n8449) );
  NAND2_X1 U5763 ( .A1(n4742), .A2(n4740), .ZN(n4745) );
  OAI21_X1 U5764 ( .B1(n8481), .B2(n8491), .A(n4746), .ZN(n8465) );
  AND2_X1 U5765 ( .A1(n8510), .A2(n8509), .ZN(n8672) );
  INV_X1 U5766 ( .A(n8669), .ZN(n8503) );
  AND2_X1 U5767 ( .A1(n8539), .A2(n8538), .ZN(n8684) );
  AND2_X1 U5768 ( .A1(n4778), .A2(n8142), .ZN(n8537) );
  NAND2_X1 U5769 ( .A1(n8565), .A2(n8139), .ZN(n8550) );
  OAI21_X1 U5770 ( .B1(n8587), .B2(n4756), .A(n4754), .ZN(n8543) );
  NAND2_X1 U5771 ( .A1(n4759), .A2(n4760), .ZN(n8558) );
  NAND2_X1 U5772 ( .A1(n8587), .A2(n4761), .ZN(n4759) );
  AND2_X1 U5773 ( .A1(n4764), .A2(n4431), .ZN(n8575) );
  NAND2_X1 U5774 ( .A1(n8587), .A2(n5461), .ZN(n4764) );
  NAND2_X1 U5775 ( .A1(n5441), .A2(n5440), .ZN(n8709) );
  NAND2_X1 U5776 ( .A1(n8629), .A2(n5432), .ZN(n8603) );
  AND2_X1 U5777 ( .A1(n4725), .A2(n4724), .ZN(n7449) );
  OR2_X1 U5778 ( .A1(n4726), .A2(n4728), .ZN(n7450) );
  NAND2_X1 U5779 ( .A1(n4708), .A2(n5309), .ZN(n7150) );
  NAND2_X1 U5780 ( .A1(n6836), .A2(n4709), .ZN(n4708) );
  NAND2_X1 U5781 ( .A1(n4704), .A2(n5245), .ZN(n6583) );
  OR2_X1 U5782 ( .A1(n5191), .A2(n6339), .ZN(n5228) );
  AOI21_X1 U5783 ( .B1(n9759), .B2(n10137), .A(n9758), .ZN(n4517) );
  OR2_X1 U5784 ( .A1(n8247), .A2(n10132), .ZN(n4519) );
  OAI21_X1 U5785 ( .B1(n5438), .B2(n4403), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5464) );
  INV_X1 U5786 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6087) );
  INV_X1 U5787 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6081) );
  OAI21_X1 U5788 ( .B1(n6538), .B2(n4425), .A(n4616), .ZN(n6525) );
  INV_X1 U5789 ( .A(n4617), .ZN(n4616) );
  NAND2_X1 U5790 ( .A1(n7675), .A2(n7747), .ZN(n4493) );
  NAND2_X1 U5791 ( .A1(n6989), .A2(n6988), .ZN(n7270) );
  NAND2_X1 U5792 ( .A1(n7583), .A2(n7582), .ZN(n9651) );
  NAND2_X1 U5793 ( .A1(n6625), .A2(n4417), .ZN(n6811) );
  NAND2_X1 U5794 ( .A1(n4607), .A2(n6633), .ZN(n6812) );
  NAND2_X1 U5795 ( .A1(n6625), .A2(n6624), .ZN(n4607) );
  INV_X1 U5796 ( .A(n9062), .ZN(n7776) );
  NAND2_X1 U5797 ( .A1(n7174), .A2(n7173), .ZN(n7177) );
  NAND2_X1 U5798 ( .A1(n7485), .A2(n7484), .ZN(n9666) );
  OAI21_X1 U5799 ( .B1(n5001), .B2(n4996), .A(n4402), .ZN(n4995) );
  INV_X1 U5800 ( .A(n9038), .ZN(n5001) );
  NAND2_X1 U5801 ( .A1(n8787), .A2(n4997), .ZN(n4996) );
  NAND2_X1 U5802 ( .A1(n7569), .A2(n7568), .ZN(n9659) );
  AOI21_X1 U5803 ( .B1(n8981), .B2(n8980), .A(n8979), .ZN(n8984) );
  INV_X1 U5804 ( .A(n9929), .ZN(n6750) );
  NOR2_X1 U5805 ( .A1(n4580), .A2(n6225), .ZN(n6230) );
  INV_X1 U5806 ( .A(n4579), .ZN(n4580) );
  NAND2_X1 U5807 ( .A1(n8947), .A2(n8831), .ZN(n9000) );
  NAND2_X1 U5808 ( .A1(n7621), .A2(n7620), .ZN(n9634) );
  INV_X1 U5809 ( .A(n7777), .ZN(n9785) );
  NAND2_X1 U5810 ( .A1(n7059), .A2(n7058), .ZN(n7064) );
  AND2_X1 U5811 ( .A1(n6378), .A2(n6377), .ZN(n9045) );
  NAND2_X1 U5812 ( .A1(n5006), .A2(n4420), .ZN(n5005) );
  INV_X1 U5813 ( .A(n5007), .ZN(n5006) );
  NAND2_X1 U5814 ( .A1(n7415), .A2(n7414), .ZN(n9669) );
  OAI21_X1 U5815 ( .B1(n4495), .B2(n7961), .A(n4494), .ZN(n7962) );
  OR2_X1 U5816 ( .A1(n7960), .A2(n9203), .ZN(n4495) );
  NAND2_X1 U5817 ( .A1(n7961), .A2(n9203), .ZN(n4494) );
  NAND2_X1 U5818 ( .A1(n7988), .A2(n6177), .ZN(n4511) );
  NAND2_X1 U5819 ( .A1(n6177), .A2(n9124), .ZN(n7992) );
  NAND2_X1 U5820 ( .A1(n6350), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6268) );
  OR2_X1 U5821 ( .A1(n7679), .A2(n9801), .ZN(n6104) );
  NAND2_X1 U5822 ( .A1(n9861), .A2(n4469), .ZN(n5898) );
  NOR2_X1 U5823 ( .A1(n5938), .A2(n4627), .ZN(n9875) );
  NOR2_X1 U5824 ( .A1(n6509), .A2(n5877), .ZN(n4627) );
  NAND2_X1 U5825 ( .A1(n9875), .A2(n9874), .ZN(n9873) );
  INV_X1 U5826 ( .A(n4632), .ZN(n6197) );
  NOR2_X1 U5827 ( .A1(n6195), .A2(n4630), .ZN(n6208) );
  AND2_X1 U5828 ( .A1(n6987), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4630) );
  INV_X1 U5829 ( .A(n4629), .ZN(n6447) );
  INV_X1 U5830 ( .A(n4620), .ZN(n9087) );
  INV_X1 U5831 ( .A(n4622), .ZN(n9074) );
  INV_X1 U5832 ( .A(n4638), .ZN(n9105) );
  NAND2_X1 U5833 ( .A1(n7725), .A2(n7724), .ZN(n7726) );
  XNOR2_X1 U5834 ( .A(n4553), .B(n7715), .ZN(n7727) );
  XNOR2_X1 U5835 ( .A(n7708), .B(n7877), .ZN(n9602) );
  OR2_X1 U5836 ( .A1(n9183), .A2(n4835), .ZN(n9170) );
  INV_X1 U5837 ( .A(n9614), .ZN(n9169) );
  AOI21_X1 U5838 ( .B1(n9177), .B2(n9185), .A(n4885), .ZN(n9162) );
  INV_X1 U5839 ( .A(n4888), .ZN(n4885) );
  NAND2_X1 U5840 ( .A1(n4849), .A2(n4855), .ZN(n9492) );
  NAND2_X1 U5841 ( .A1(n9524), .A2(n4858), .ZN(n4849) );
  NAND2_X1 U5842 ( .A1(n4556), .A2(n4560), .ZN(n9516) );
  NAND2_X1 U5843 ( .A1(n9538), .A2(n4416), .ZN(n4556) );
  AND2_X1 U5844 ( .A1(n4861), .A2(n4432), .ZN(n9507) );
  NAND2_X1 U5845 ( .A1(n9524), .A2(n7604), .ZN(n4861) );
  INV_X1 U5846 ( .A(n9644), .ZN(n9530) );
  OAI21_X1 U5847 ( .B1(n7411), .B2(n4870), .A(n4867), .ZN(n7566) );
  NAND2_X1 U5848 ( .A1(n7411), .A2(n4872), .ZN(n4866) );
  NAND2_X1 U5849 ( .A1(n7164), .A2(n7163), .ZN(n7327) );
  NAND2_X1 U5850 ( .A1(n7030), .A2(n7029), .ZN(n7137) );
  NAND2_X1 U5851 ( .A1(n6816), .A2(n6815), .ZN(n7759) );
  NAND2_X1 U5852 ( .A1(n6932), .A2(n6886), .ZN(n6927) );
  INV_X1 U5853 ( .A(n10003), .ZN(n6946) );
  NAND2_X1 U5854 ( .A1(n6855), .A2(n6892), .ZN(n6937) );
  NAND2_X1 U5855 ( .A1(n6879), .A2(n6878), .ZN(n10001) );
  NOR2_X1 U5856 ( .A1(n5919), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U5857 ( .A1(n4893), .A2(n5051), .ZN(n5290) );
  NAND2_X1 U5858 ( .A1(n5276), .A2(n5275), .ZN(n4893) );
  NOR2_X1 U5859 ( .A1(n5885), .A2(n5884), .ZN(n9844) );
  AND2_X1 U5860 ( .A1(n5847), .A2(n5846), .ZN(n5881) );
  INV_X1 U5861 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9409) );
  NAND2_X1 U5862 ( .A1(n5883), .A2(n4626), .ZN(n4625) );
  OR2_X1 U5863 ( .A1(n5887), .A2(n4624), .ZN(n4623) );
  NAND2_X1 U5864 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4624) );
  NOR2_X1 U5865 ( .A1(n9717), .A2(n10209), .ZN(n10219) );
  NOR2_X1 U5866 ( .A1(n10219), .A2(n10218), .ZN(n10217) );
  NOR2_X1 U5867 ( .A1(n9723), .A2(n10224), .ZN(n10208) );
  AOI21_X1 U5868 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10206), .ZN(n10205) );
  NOR2_X1 U5869 ( .A1(n10205), .A2(n10204), .ZN(n10203) );
  NAND2_X1 U5870 ( .A1(n5702), .A2(n5701), .ZN(n6415) );
  OAI21_X1 U5871 ( .B1(n4449), .B2(n4508), .A(n4507), .ZN(P2_U3242) );
  AND2_X1 U5872 ( .A1(n8337), .A2(n4474), .ZN(n4507) );
  NAND2_X1 U5873 ( .A1(n4509), .A2(n8321), .ZN(n4508) );
  OAI21_X1 U5874 ( .B1(n8414), .B2(n5638), .A(n4960), .ZN(P2_U3264) );
  AOI21_X1 U5875 ( .B1(n4962), .B2(n5638), .A(n4961), .ZN(n4960) );
  NAND2_X1 U5876 ( .A1(n4404), .A2(n4436), .ZN(P2_U3267) );
  NAND2_X1 U5877 ( .A1(n8246), .A2(n8644), .ZN(n4500) );
  MUX2_X1 U5878 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n5688), .S(n10177), .Z(
        P2_U3549) );
  NOR2_X1 U5879 ( .A1(n4427), .A2(n4602), .ZN(n4601) );
  INV_X1 U5880 ( .A(n4644), .ZN(n4643) );
  NAND2_X1 U5881 ( .A1(n9125), .A2(n9124), .ZN(n4645) );
  NAND2_X1 U5882 ( .A1(n4641), .A2(n9203), .ZN(n4640) );
  NAND2_X1 U5883 ( .A1(n9676), .A2(n10049), .ZN(n4836) );
  NAND2_X1 U5884 ( .A1(n8240), .A2(n8442), .ZN(n4400) );
  INV_X2 U5885 ( .A(n6172), .ZN(n6350) );
  INV_X4 U5886 ( .A(n5194), .ZN(n5204) );
  NAND2_X2 U5887 ( .A1(n7653), .A2(n7652), .ZN(n9619) );
  MUX2_X1 U5888 ( .A(n9703), .B(n9806), .S(n6250), .Z(n9929) );
  NAND2_X1 U5889 ( .A1(n8077), .A2(n8073), .ZN(n5625) );
  OR2_X1 U5890 ( .A1(n8964), .A2(n8965), .ZN(n4402) );
  INV_X1 U5891 ( .A(n7251), .ZN(n10147) );
  OR2_X1 U5892 ( .A1(n8244), .A2(n8646), .ZN(n4404) );
  NAND2_X1 U5893 ( .A1(n6853), .A2(n6865), .ZN(n6868) );
  AND2_X1 U5894 ( .A1(n8147), .A2(n8173), .ZN(n4405) );
  AND2_X1 U5895 ( .A1(n4487), .A2(n4486), .ZN(n4406) );
  NAND2_X1 U5896 ( .A1(n7314), .A2(n7313), .ZN(n8774) );
  OR2_X1 U5897 ( .A1(n7962), .A2(n6177), .ZN(n4407) );
  NAND2_X1 U5898 ( .A1(n5009), .A2(n5010), .ZN(n8956) );
  AND3_X1 U5899 ( .A1(n4989), .A2(n5152), .A3(n5154), .ZN(n4408) );
  AND2_X1 U5900 ( .A1(n8712), .A2(n8613), .ZN(n8114) );
  INV_X1 U5901 ( .A(n8114), .ZN(n4793) );
  AND2_X1 U5902 ( .A1(n8211), .A2(n4444), .ZN(n4409) );
  INV_X1 U5903 ( .A(n8430), .ZN(n8439) );
  XNOR2_X1 U5904 ( .A(n8649), .B(n8459), .ZN(n8430) );
  OR2_X1 U5905 ( .A1(n8123), .A2(n8132), .ZN(n4410) );
  AND2_X1 U5906 ( .A1(n8113), .A2(n4793), .ZN(n8627) );
  INV_X1 U5907 ( .A(n8627), .ZN(n5430) );
  AND2_X1 U5908 ( .A1(n5542), .A2(n5541), .ZN(n8330) );
  OR2_X1 U5909 ( .A1(n8240), .A2(n8442), .ZN(n8026) );
  INV_X1 U5910 ( .A(n8026), .ZN(n4819) );
  INV_X1 U5911 ( .A(n4400), .ZN(n4816) );
  AND2_X1 U5912 ( .A1(n7031), .A2(n7029), .ZN(n4411) );
  AND2_X1 U5913 ( .A1(n5708), .A2(n5701), .ZN(n4412) );
  INV_X1 U5914 ( .A(n8103), .ZN(n8346) );
  AND4_X1 U5915 ( .A1(n5401), .A2(n5400), .A3(n5399), .A4(n5398), .ZN(n8103)
         );
  INV_X1 U5916 ( .A(n6883), .ZN(n9999) );
  INV_X1 U5917 ( .A(n10128), .ZN(n4513) );
  AND2_X1 U5918 ( .A1(n8847), .A2(n4588), .ZN(n4415) );
  NAND2_X1 U5919 ( .A1(n5178), .A2(n8763), .ZN(n5205) );
  INV_X1 U5920 ( .A(n8342), .ZN(n4491) );
  NAND2_X1 U5921 ( .A1(n4591), .A2(n8906), .ZN(n8947) );
  NAND2_X2 U5922 ( .A1(n6628), .A2(n4498), .ZN(n6476) );
  INV_X1 U5923 ( .A(n4943), .ZN(n7836) );
  AND2_X1 U5924 ( .A1(n7852), .A2(n4561), .ZN(n4416) );
  NAND2_X2 U5925 ( .A1(n7686), .A2(n7685), .ZN(n9603) );
  AND2_X1 U5926 ( .A1(n6624), .A2(n6632), .ZN(n4417) );
  INV_X1 U5927 ( .A(n8201), .ZN(n4727) );
  INV_X1 U5928 ( .A(n6251), .ZN(n5038) );
  NAND2_X1 U5929 ( .A1(n7780), .A2(n7778), .ZN(n7865) );
  NAND2_X1 U5930 ( .A1(n4740), .A2(n4739), .ZN(n4738) );
  OR2_X1 U5931 ( .A1(n7151), .A2(n4707), .ZN(n4418) );
  AND2_X1 U5932 ( .A1(n5944), .A2(n4615), .ZN(n4419) );
  NAND2_X1 U5933 ( .A1(n8873), .A2(n8872), .ZN(n4420) );
  NAND2_X1 U5934 ( .A1(n10147), .A2(n8350), .ZN(n8077) );
  AND3_X1 U5935 ( .A1(n4671), .A2(n4670), .A3(n7897), .ZN(n4421) );
  AND2_X1 U5936 ( .A1(n8468), .A2(n8157), .ZN(n8491) );
  INV_X1 U5937 ( .A(n8491), .ZN(n4748) );
  AND2_X1 U5938 ( .A1(n8698), .A2(n8596), .ZN(n4422) );
  OR2_X1 U5939 ( .A1(n8654), .A2(n8341), .ZN(n4423) );
  INV_X1 U5940 ( .A(n8109), .ZN(n4797) );
  NOR2_X1 U5941 ( .A1(n9539), .A2(n7913), .ZN(n4424) );
  NAND2_X1 U5942 ( .A1(n6517), .A2(n6573), .ZN(n4425) );
  NAND2_X1 U5943 ( .A1(n9614), .A2(n9056), .ZN(n4426) );
  AND3_X1 U5944 ( .A1(n8933), .A2(n8982), .A3(n8932), .ZN(n4427) );
  INV_X1 U5945 ( .A(n8108), .ZN(n4796) );
  NAND2_X1 U5946 ( .A1(n4399), .A2(n4498), .ZN(n5191) );
  OR2_X1 U5947 ( .A1(n8544), .A2(n8308), .ZN(n4428) );
  AND2_X1 U5948 ( .A1(n4642), .A2(n9818), .ZN(n4429) );
  NAND2_X1 U5949 ( .A1(n4582), .A2(n4415), .ZN(n8853) );
  AND4_X1 U5950 ( .A1(n4576), .A2(n4575), .A3(n4574), .A4(n5926), .ZN(n4430)
         );
  NAND2_X1 U5951 ( .A1(n8592), .A2(n8614), .ZN(n4431) );
  NAND2_X1 U5952 ( .A1(n9530), .A2(n9545), .ZN(n4432) );
  OAI211_X1 U5953 ( .C1(n6339), .C2(n6813), .A(n6338), .B(n6337), .ZN(n6865)
         );
  NAND2_X1 U5954 ( .A1(n8148), .A2(n5634), .ZN(n8524) );
  AND3_X1 U5955 ( .A1(n7842), .A2(n7841), .A3(n7843), .ZN(n4433) );
  NAND2_X1 U5956 ( .A1(n8174), .A2(n8170), .ZN(n8214) );
  INV_X1 U5957 ( .A(n4890), .ZN(n5864) );
  OR2_X1 U5958 ( .A1(n9066), .A2(n6926), .ZN(n4434) );
  OR2_X1 U5959 ( .A1(n5864), .A2(n5012), .ZN(n5858) );
  OR2_X1 U5960 ( .A1(n4399), .A2(n6072), .ZN(n4435) );
  AND2_X1 U5961 ( .A1(n4501), .A2(n4500), .ZN(n4436) );
  NAND2_X1 U5962 ( .A1(n7948), .A2(n7907), .ZN(n9155) );
  INV_X1 U5963 ( .A(n9155), .ZN(n4694) );
  AND2_X1 U5964 ( .A1(n7875), .A2(n7830), .ZN(n4437) );
  NAND2_X1 U5965 ( .A1(n4861), .A2(n4860), .ZN(n4438) );
  AND2_X1 U5966 ( .A1(n5009), .A2(n5007), .ZN(n4439) );
  NAND2_X1 U5967 ( .A1(n5537), .A2(n5536), .ZN(n8666) );
  INV_X1 U5968 ( .A(n8666), .ZN(n4747) );
  INV_X1 U5969 ( .A(n8649), .ZN(n8437) );
  NAND2_X1 U5970 ( .A1(n5582), .A2(n5581), .ZN(n8649) );
  AND2_X1 U5971 ( .A1(n5448), .A2(n5432), .ZN(n4440) );
  AND2_X1 U5972 ( .A1(n4455), .A2(n8170), .ZN(n4441) );
  AND2_X1 U5973 ( .A1(n7066), .A2(n7058), .ZN(n4442) );
  OR3_X1 U5974 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4443) );
  AND2_X1 U5975 ( .A1(n8168), .A2(n8167), .ZN(n4444) );
  NAND2_X1 U5976 ( .A1(n4650), .A2(n6852), .ZN(n6891) );
  AND2_X1 U5977 ( .A1(n5519), .A2(n5518), .ZN(n8522) );
  INV_X1 U5978 ( .A(n8522), .ZN(n8674) );
  AND2_X1 U5979 ( .A1(n8669), .A2(n4491), .ZN(n8146) );
  AND2_X1 U5980 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n4445) );
  NAND2_X1 U5981 ( .A1(n9498), .A2(n7617), .ZN(n9506) );
  AOI21_X1 U5982 ( .B1(n8014), .B2(n8015), .A(n8013), .ZN(n8425) );
  NAND2_X1 U5983 ( .A1(n8999), .A2(n9003), .ZN(n4446) );
  INV_X1 U5984 ( .A(n4868), .ZN(n4867) );
  OAI22_X1 U5985 ( .A1(n7786), .A2(n4869), .B1(n8967), .B2(n7481), .ZN(n4868)
         );
  INV_X1 U5986 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4626) );
  NOR2_X1 U5987 ( .A1(n8654), .A2(n8441), .ZN(n4447) );
  NOR2_X1 U5988 ( .A1(n9201), .A2(n9057), .ZN(n4448) );
  AND2_X1 U5989 ( .A1(n4972), .A2(n4970), .ZN(n4449) );
  AND2_X1 U5990 ( .A1(n8206), .A2(n4542), .ZN(n4450) );
  INV_X1 U5991 ( .A(n4807), .ZN(n4806) );
  NAND2_X1 U5992 ( .A1(n8159), .A2(n8456), .ZN(n4807) );
  INV_X1 U5993 ( .A(n4569), .ZN(n4568) );
  OAI21_X1 U5994 ( .B1(n9194), .B2(n4570), .A(n7821), .ZN(n4569) );
  OR2_X1 U5995 ( .A1(n5864), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n4451) );
  AND2_X1 U5996 ( .A1(n7709), .A2(n7923), .ZN(n7786) );
  OAI21_X1 U5997 ( .B1(n8456), .B2(n4744), .A(n4423), .ZN(n4743) );
  OR2_X1 U5998 ( .A1(n8649), .A2(n8459), .ZN(n4452) );
  AND2_X1 U5999 ( .A1(n5054), .A2(SI_7_), .ZN(n4453) );
  AND2_X1 U6000 ( .A1(n4426), .A2(n4886), .ZN(n4454) );
  NAND2_X1 U6001 ( .A1(n8425), .A2(n8340), .ZN(n4455) );
  NAND2_X1 U6002 ( .A1(n7227), .A2(n5752), .ZN(n4456) );
  INV_X1 U6003 ( .A(n4873), .ZN(n4872) );
  NOR2_X1 U6004 ( .A1(n9768), .A2(n9042), .ZN(n4873) );
  NOR2_X1 U6005 ( .A1(n8564), .A2(n8553), .ZN(n4457) );
  NAND2_X1 U6006 ( .A1(n7863), .A2(n4830), .ZN(n4458) );
  NAND2_X1 U6007 ( .A1(n8142), .A2(n8137), .ZN(n4459) );
  INV_X1 U6008 ( .A(n4738), .ZN(n4737) );
  OR2_X1 U6009 ( .A1(n5864), .A2(n4401), .ZN(n4460) );
  AND2_X1 U6010 ( .A1(n8990), .A2(n8833), .ZN(n8844) );
  INV_X1 U6011 ( .A(n8113), .ZN(n4792) );
  AND2_X1 U6012 ( .A1(n4989), .A2(n5152), .ZN(n4461) );
  NOR2_X1 U6013 ( .A1(n4813), .A2(n8214), .ZN(n4462) );
  NOR2_X1 U6014 ( .A1(n9183), .A2(n7712), .ZN(n4463) );
  INV_X1 U6015 ( .A(n6893), .ZN(n4651) );
  AND2_X1 U6016 ( .A1(n4419), .A2(n6142), .ZN(n4464) );
  INV_X1 U6017 ( .A(n7819), .ZN(n4570) );
  AND2_X1 U6018 ( .A1(n4834), .A2(n4566), .ZN(n4465) );
  AND2_X1 U6019 ( .A1(n7175), .A2(n7173), .ZN(n4466) );
  AND2_X1 U6020 ( .A1(n4420), .A2(n8867), .ZN(n4467) );
  NAND2_X1 U6021 ( .A1(n8418), .A2(n8020), .ZN(n8175) );
  AND2_X1 U6022 ( .A1(n7781), .A2(n7780), .ZN(n4468) );
  INV_X1 U6023 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5849) );
  OR2_X1 U6024 ( .A1(n9860), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4469) );
  INV_X1 U6025 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n4949) );
  NAND2_X1 U6026 ( .A1(n4785), .A2(n4783), .ZN(n8593) );
  NAND2_X1 U6027 ( .A1(n4866), .A2(n4871), .ZN(n7482) );
  NAND2_X1 U6028 ( .A1(n8787), .A2(n9038), .ZN(n8963) );
  INV_X1 U6029 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5013) );
  INV_X1 U6030 ( .A(n8906), .ZN(n4590) );
  NAND2_X1 U6031 ( .A1(n5615), .A2(n8043), .ZN(n8186) );
  OAI21_X1 U6032 ( .B1(n6288), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6312) );
  AND2_X1 U6033 ( .A1(n5658), .A2(n5152), .ZN(n5652) );
  NAND2_X1 U6034 ( .A1(n6839), .A2(n8065), .ZN(n7084) );
  OR2_X1 U6035 ( .A1(n5301), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n4470) );
  NAND2_X1 U6036 ( .A1(n4724), .A2(n4718), .ZN(n8626) );
  NAND2_X1 U6037 ( .A1(n4991), .A2(n4603), .ZN(n9037) );
  AND2_X1 U6038 ( .A1(n9172), .A2(n9913), .ZN(n4471) );
  OR2_X1 U6039 ( .A1(n5438), .A2(n5437), .ZN(n4472) );
  NAND2_X1 U6040 ( .A1(n5418), .A2(n5436), .ZN(n4473) );
  OR2_X1 U6041 ( .A1(n8339), .A2(n8338), .ZN(n4474) );
  NOR2_X1 U6042 ( .A1(n9138), .A2(n4471), .ZN(n4475) );
  AND2_X1 U6043 ( .A1(n5383), .A2(n8200), .ZN(n4476) );
  INV_X1 U6044 ( .A(n4995), .ZN(n8973) );
  INV_X1 U6045 ( .A(n8166), .ZN(n8173) );
  NAND2_X1 U6046 ( .A1(n7059), .A2(n4442), .ZN(n7174) );
  NAND2_X1 U6047 ( .A1(n5393), .A2(n5392), .ZN(n8723) );
  INV_X1 U6048 ( .A(n8723), .ZN(n4730) );
  NAND2_X1 U6049 ( .A1(n7282), .A2(n7281), .ZN(n7407) );
  INV_X1 U6050 ( .A(n7407), .ZN(n4486) );
  NAND2_X1 U6051 ( .A1(n5652), .A2(n5153), .ZN(n5655) );
  AOI21_X1 U6052 ( .B1(n6872), .B2(n6871), .A(n6870), .ZN(n6903) );
  AND2_X1 U6053 ( .A1(n7280), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4478) );
  NOR2_X1 U6054 ( .A1(n7560), .A2(n7559), .ZN(n4479) );
  OAI21_X1 U6055 ( .B1(n6625), .B2(n4611), .A(n4608), .ZN(n6980) );
  NAND2_X1 U6056 ( .A1(n4994), .A2(n6347), .ZN(n6483) );
  AND2_X1 U6057 ( .A1(n7162), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4480) );
  NAND2_X1 U6058 ( .A1(n6523), .A2(n6522), .ZN(n6625) );
  NAND2_X1 U6059 ( .A1(n4848), .A2(n6885), .ZN(n6932) );
  NOR2_X1 U6060 ( .A1(n8420), .A2(n8024), .ZN(n4481) );
  INV_X1 U6061 ( .A(n4904), .ZN(n4903) );
  NAND2_X1 U6062 ( .A1(n4906), .A2(n4905), .ZN(n4904) );
  NAND4_X1 U6063 ( .A1(n6473), .A2(n6472), .A3(n6471), .A4(n6470), .ZN(n9066)
         );
  INV_X1 U6064 ( .A(n9066), .ZN(n4843) );
  INV_X1 U6065 ( .A(n8004), .ZN(n4936) );
  INV_X1 U6066 ( .A(n10034), .ZN(n9995) );
  OR2_X1 U6067 ( .A1(n10049), .A2(n7687), .ZN(n4482) );
  INV_X1 U6068 ( .A(n5739), .ZN(n4515) );
  NAND2_X1 U6069 ( .A1(n6631), .A2(n6630), .ZN(n10020) );
  INV_X1 U6070 ( .A(n10020), .ZN(n4488) );
  XNOR2_X1 U6071 ( .A(n6262), .B(n6260), .ZN(n8936) );
  INV_X1 U6072 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4615) );
  NAND2_X1 U6073 ( .A1(n4613), .A2(n6147), .ZN(n9124) );
  INV_X1 U6074 ( .A(n9124), .ZN(n9203) );
  NOR2_X1 U6075 ( .A1(n5173), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8755) );
  OR2_X1 U6076 ( .A1(n8179), .A2(n10097), .ZN(n4483) );
  AOI21_X1 U6077 ( .B1(n5646), .B2(n10061), .A(n5645), .ZN(n8244) );
  MUX2_X1 U6078 ( .A(n7751), .B(n9055), .S(n7835), .Z(n7833) );
  NAND2_X1 U6079 ( .A1(n4669), .A2(n7835), .ZN(n4668) );
  INV_X1 U6080 ( .A(n7835), .ZN(n4699) );
  OR2_X1 U6081 ( .A1(n5910), .A2(P1_U3084), .ZN(n9833) );
  INV_X1 U6082 ( .A(n8950), .ZN(n4510) );
  OAI21_X1 U6083 ( .B1(n5463), .B2(n5462), .A(n5122), .ZN(n5481) );
  AOI21_X1 U6084 ( .B1(n8831), .B2(n4590), .A(n4446), .ZN(n4589) );
  NAND2_X1 U6085 ( .A1(n4484), .A2(n5005), .ZN(n9025) );
  NAND3_X1 U6086 ( .A1(n8980), .A2(n8981), .A3(n4467), .ZN(n4484) );
  INV_X1 U6087 ( .A(n6525), .ZN(n6523) );
  NAND2_X1 U6088 ( .A1(n4994), .A2(n4992), .ZN(n6538) );
  NAND2_X1 U6089 ( .A1(n4618), .A2(n4998), .ZN(n8805) );
  NOR2_X1 U6090 ( .A1(n6225), .A2(n4578), .ZN(n4577) );
  OR2_X1 U6091 ( .A1(n8909), .A2(n4587), .ZN(n4584) );
  NAND2_X1 U6092 ( .A1(n9606), .A2(n4837), .ZN(n9676) );
  OAI21_X1 U6093 ( .B1(n9575), .B2(n7570), .A(n7795), .ZN(n9558) );
  NAND2_X1 U6094 ( .A1(n9556), .A2(n5018), .ZN(n9537) );
  AOI21_X1 U6095 ( .B1(n4848), .B2(n4847), .A(n4844), .ZN(n6950) );
  NAND2_X2 U6096 ( .A1(n9491), .A2(n7813), .ZN(n9476) );
  OAI21_X1 U6097 ( .B1(n7411), .B2(n4864), .A(n4863), .ZN(n4862) );
  NOR2_X1 U6098 ( .A1(n7863), .A2(n7188), .ZN(n7325) );
  INV_X1 U6099 ( .A(n9607), .ZN(n4839) );
  NAND2_X2 U6100 ( .A1(n4571), .A2(n5872), .ZN(n6250) );
  NOR2_X2 U6101 ( .A1(n7199), .A2(n7327), .ZN(n4487) );
  INV_X1 U6102 ( .A(n4512), .ZN(n9148) );
  NAND2_X2 U6103 ( .A1(n4490), .A2(n9999), .ZN(n6944) );
  INV_X1 U6104 ( .A(n6912), .ZN(n4490) );
  NAND3_X1 U6105 ( .A1(n5025), .A2(n4772), .A3(n4771), .ZN(n4769) );
  OAI211_X1 U6106 ( .C1(n4483), .C2(n4549), .A(n4548), .B(n4547), .ZN(n4546)
         );
  AOI21_X1 U6107 ( .B1(n4810), .B2(n4462), .A(n4808), .ZN(n8021) );
  NAND2_X1 U6108 ( .A1(n4544), .A2(n8229), .ZN(P2_U3244) );
  OAI21_X1 U6109 ( .B1(n5385), .B2(n5093), .A(n5096), .ZN(n5402) );
  NAND2_X1 U6110 ( .A1(n4917), .A2(n4918), .ZN(n5567) );
  OAI21_X2 U6111 ( .B1(n5306), .B2(n5304), .A(n5059), .ZN(n5319) );
  NAND2_X1 U6112 ( .A1(n4496), .A2(n5043), .ZN(n5257) );
  NAND3_X1 U6113 ( .A1(n4775), .A2(n5241), .A3(n4773), .ZN(n4496) );
  NAND2_X2 U6114 ( .A1(n4499), .A2(n7643), .ZN(n9201) );
  OAI21_X1 U6115 ( .B1(n7963), .B2(n4407), .A(n4511), .ZN(n7999) );
  NOR2_X1 U6116 ( .A1(n4933), .A2(n4932), .ZN(n4931) );
  NAND2_X1 U6117 ( .A1(n4809), .A2(n8175), .ZN(n4808) );
  NAND2_X1 U6118 ( .A1(n4892), .A2(n4891), .ZN(n5306) );
  OAI21_X1 U6119 ( .B1(n8221), .B2(n4546), .A(n4545), .ZN(n4544) );
  NAND2_X1 U6120 ( .A1(n8223), .A2(n8222), .ZN(n4547) );
  OAI21_X1 U6121 ( .B1(n5402), .B2(n5403), .A(n5101), .ZN(n5415) );
  NAND2_X1 U6122 ( .A1(n5785), .A2(n5784), .ZN(n8269) );
  NAND2_X1 U6123 ( .A1(n5800), .A2(n5799), .ZN(n5801) );
  NOR2_X1 U6124 ( .A1(n5607), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U6125 ( .A1(n6712), .A2(n6713), .ZN(n6711) );
  NOR2_X1 U6126 ( .A1(n9135), .A2(n7714), .ZN(n4553) );
  NOR2_X1 U6127 ( .A1(n9153), .A2(n7713), .ZN(n9137) );
  NOR2_X1 U6128 ( .A1(n5811), .A2(n5810), .ZN(n8285) );
  OAI22_X1 U6129 ( .A1(n6303), .A2(n6302), .B1(n5697), .B2(n5696), .ZN(n6391)
         );
  NAND2_X2 U6130 ( .A1(n8450), .A2(n8437), .ZN(n8432) );
  XNOR2_X2 U6131 ( .A(n8423), .B(n8418), .ZN(n8648) );
  NAND2_X1 U6132 ( .A1(n5658), .A2(n4461), .ZN(n5664) );
  INV_X1 U6133 ( .A(n9025), .ZN(n4600) );
  NAND2_X1 U6134 ( .A1(n5128), .A2(n5127), .ZN(n5493) );
  MUX2_X1 U6135 ( .A(n7824), .B(n7911), .S(n7835), .Z(n7827) );
  INV_X1 U6136 ( .A(n4895), .ZN(n4894) );
  NAND2_X1 U6137 ( .A1(n5319), .A2(n4914), .ZN(n4912) );
  INV_X1 U6138 ( .A(n4690), .ZN(n4689) );
  NAND2_X1 U6139 ( .A1(n4930), .A2(n5131), .ZN(n5503) );
  NAND2_X1 U6140 ( .A1(n5415), .A2(n5414), .ZN(n5107) );
  NOR2_X1 U6141 ( .A1(n4573), .A2(n4572), .ZN(n4571) );
  NAND2_X1 U6142 ( .A1(n5854), .A2(n5013), .ZN(n5012) );
  NAND2_X1 U6143 ( .A1(n4979), .A2(n5255), .ZN(n5345) );
  NAND3_X1 U6144 ( .A1(n5651), .A2(n8244), .A3(n4519), .ZN(n5688) );
  NAND2_X1 U6145 ( .A1(n8117), .A2(n4526), .ZN(n4525) );
  NAND2_X1 U6146 ( .A1(n8117), .A2(n8116), .ZN(n4528) );
  NAND2_X1 U6147 ( .A1(n4532), .A2(n4531), .ZN(n8068) );
  INV_X1 U6148 ( .A(n4536), .ZN(n5465) );
  NOR2_X2 U6149 ( .A1(n5349), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5367) );
  AND2_X2 U6150 ( .A1(n5605), .A2(n4550), .ZN(n5638) );
  OAI21_X1 U6151 ( .B1(n9538), .B2(n4559), .A(n4557), .ZN(n9515) );
  NAND2_X1 U6152 ( .A1(n9477), .A2(n4465), .ZN(n4564) );
  NAND2_X1 U6153 ( .A1(n9477), .A2(n4566), .ZN(n4565) );
  AOI21_X1 U6154 ( .B1(n9477), .B2(n7815), .A(n7819), .ZN(n9195) );
  AND2_X2 U6155 ( .A1(n5866), .A2(n5868), .ZN(n4890) );
  INV_X1 U6156 ( .A(n6245), .ZN(n4578) );
  INV_X1 U6157 ( .A(n8909), .ZN(n4593) );
  NAND2_X1 U6158 ( .A1(n4581), .A2(n4585), .ZN(n8851) );
  NAND3_X1 U6159 ( .A1(n8934), .A2(n4601), .A3(n4594), .ZN(P1_U3218) );
  NAND2_X1 U6160 ( .A1(n6625), .A2(n4608), .ZN(n4604) );
  NAND2_X1 U6161 ( .A1(n4604), .A2(n4605), .ZN(n6985) );
  XNOR2_X2 U6162 ( .A(n4612), .B(n6145), .ZN(n6177) );
  NAND2_X1 U6163 ( .A1(n4614), .A2(n4464), .ZN(n6288) );
  NAND2_X1 U6164 ( .A1(n7174), .A2(n4466), .ZN(n7286) );
  OAI21_X1 U6165 ( .B1(n6498), .B2(n4425), .A(n6572), .ZN(n4617) );
  NAND3_X1 U6166 ( .A1(n8787), .A2(n5000), .A3(n9038), .ZN(n4618) );
  NAND3_X1 U6167 ( .A1(n5888), .A2(n4625), .A3(n4623), .ZN(n6077) );
  NAND3_X1 U6168 ( .A1(n4645), .A2(n4643), .A3(n4640), .ZN(P1_U3260) );
  AND2_X1 U6169 ( .A1(n6105), .A2(n6103), .ZN(n4646) );
  NAND2_X1 U6170 ( .A1(n6356), .A2(n8942), .ZN(n6229) );
  NAND3_X1 U6171 ( .A1(n6729), .A2(n6893), .A3(n6851), .ZN(n4649) );
  NAND2_X1 U6172 ( .A1(n4652), .A2(n7773), .ZN(n7775) );
  NAND2_X1 U6173 ( .A1(n4657), .A2(n4653), .ZN(n4652) );
  NAND2_X1 U6174 ( .A1(n4655), .A2(n4654), .ZN(n4653) );
  NAND2_X1 U6175 ( .A1(n4656), .A2(n7771), .ZN(n4655) );
  OAI21_X1 U6176 ( .B1(n7767), .B2(n7766), .A(n7765), .ZN(n4656) );
  AOI21_X1 U6177 ( .B1(n7772), .B2(n7835), .A(n7031), .ZN(n4657) );
  INV_X1 U6178 ( .A(n7779), .ZN(n4675) );
  INV_X1 U6179 ( .A(n7888), .ZN(n4677) );
  INV_X1 U6180 ( .A(n7890), .ZN(n4678) );
  INV_X1 U6181 ( .A(n4682), .ZN(n4681) );
  OAI21_X1 U6182 ( .B1(n4686), .B2(n4685), .A(n4692), .ZN(n4682) );
  NAND2_X1 U6183 ( .A1(n7828), .A2(n4684), .ZN(n4683) );
  INV_X1 U6184 ( .A(n4686), .ZN(n4684) );
  INV_X1 U6185 ( .A(n4687), .ZN(n4685) );
  NAND3_X1 U6186 ( .A1(n4890), .A2(n4889), .A3(n6094), .ZN(n8001) );
  NAND2_X1 U6187 ( .A1(n6855), .A2(n4697), .ZN(n4696) );
  XNOR2_X1 U6188 ( .A(n4700), .B(n4699), .ZN(n7754) );
  INV_X1 U6189 ( .A(n4700), .ZN(n7752) );
  NAND2_X1 U6190 ( .A1(n6595), .A2(n6601), .ZN(n4704) );
  NAND2_X1 U6191 ( .A1(n4704), .A2(n4702), .ZN(n4701) );
  NAND2_X1 U6192 ( .A1(n4701), .A2(n5260), .ZN(n6757) );
  AOI21_X1 U6193 ( .B1(n6757), .B2(n6759), .A(n5279), .ZN(n6835) );
  INV_X1 U6194 ( .A(n7238), .ZN(n5333) );
  NOR2_X1 U6195 ( .A1(n5607), .A2(n4713), .ZN(n5170) );
  INV_X1 U6196 ( .A(n5607), .ZN(n4712) );
  NAND2_X1 U6197 ( .A1(n5021), .A2(n8200), .ZN(n4723) );
  NAND2_X1 U6198 ( .A1(n7237), .A2(n4716), .ZN(n4724) );
  NAND2_X1 U6199 ( .A1(n4728), .A2(n8201), .ZN(n4725) );
  NOR2_X1 U6200 ( .A1(n4722), .A2(n4719), .ZN(n4718) );
  NAND2_X1 U6201 ( .A1(n8201), .A2(n4721), .ZN(n4720) );
  OAI21_X1 U6202 ( .B1(n8481), .B2(n4734), .A(n4732), .ZN(n4731) );
  NAND2_X1 U6203 ( .A1(n8481), .A2(n4746), .ZN(n4742) );
  NAND2_X1 U6204 ( .A1(n4753), .A2(n8587), .ZN(n4752) );
  INV_X1 U6205 ( .A(n5345), .ZN(n5150) );
  AND2_X2 U6206 ( .A1(n6751), .A2(n6725), .ZN(n9907) );
  OR2_X2 U6207 ( .A1(n9906), .A2(n6915), .ZN(n6912) );
  AOI21_X1 U6208 ( .B1(n9598), .B2(n7729), .A(n9127), .ZN(n9599) );
  NOR2_X2 U6209 ( .A1(n6961), .A2(n7759), .ZN(n7047) );
  NAND2_X1 U6210 ( .A1(n6835), .A2(n8060), .ZN(n6836) );
  AOI21_X1 U6211 ( .B1(n8528), .B2(n8208), .A(n5513), .ZN(n8525) );
  NAND3_X1 U6212 ( .A1(n7084), .A2(n5627), .A3(n8063), .ZN(n4765) );
  INV_X1 U6213 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4771) );
  NAND2_X1 U6214 ( .A1(n5037), .A2(n5036), .ZN(n5227) );
  NAND2_X1 U6215 ( .A1(n5041), .A2(n4774), .ZN(n4773) );
  INV_X1 U6216 ( .A(n5226), .ZN(n4774) );
  NAND3_X1 U6217 ( .A1(n5041), .A2(n5037), .A3(n5036), .ZN(n4775) );
  NAND2_X1 U6218 ( .A1(n4776), .A2(n5041), .ZN(n5242) );
  NAND2_X1 U6219 ( .A1(n5227), .A2(n5226), .ZN(n4776) );
  NAND2_X1 U6220 ( .A1(n4777), .A2(n8077), .ZN(n7378) );
  NAND3_X1 U6221 ( .A1(n8067), .A2(n8077), .A3(n8073), .ZN(n4777) );
  INV_X1 U6222 ( .A(n4777), .ZN(n8070) );
  NAND2_X1 U6223 ( .A1(n8565), .A2(n4780), .ZN(n4782) );
  CLKBUF_X1 U6224 ( .A(n4782), .Z(n4778) );
  INV_X1 U6225 ( .A(n4778), .ZN(n8549) );
  NAND2_X1 U6226 ( .A1(n7447), .A2(n4787), .ZN(n4785) );
  INV_X1 U6227 ( .A(n8515), .ZN(n4799) );
  NOR2_X1 U6228 ( .A1(n8514), .A2(n8147), .ZN(n8506) );
  OAI21_X2 U6229 ( .B1(n8489), .B2(n4807), .A(n4804), .ZN(n8438) );
  INV_X1 U6230 ( .A(n8012), .ZN(n4810) );
  NAND2_X1 U6231 ( .A1(n4836), .A2(n4482), .ZN(P1_U3551) );
  AOI21_X1 U6232 ( .B1(n9137), .B2(n9136), .A(n9588), .ZN(n4841) );
  MUX2_X1 U6233 ( .A(n6081), .B(n9409), .S(n5038), .Z(n5039) );
  MUX2_X1 U6234 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n7743), .Z(n5042) );
  MUX2_X1 U6235 ( .A(n6089), .B(n6510), .S(n7743), .Z(n5049) );
  MUX2_X1 U6236 ( .A(n6120), .B(n5060), .S(n7743), .Z(n5062) );
  MUX2_X1 U6237 ( .A(n9440), .B(n5077), .S(n7743), .Z(n5079) );
  NAND2_X1 U6238 ( .A1(n7856), .A2(n4846), .ZN(n4845) );
  AND2_X1 U6239 ( .A1(n9666), .A2(n9593), .ZN(n4874) );
  NAND2_X1 U6240 ( .A1(n9476), .A2(n4878), .ZN(n4876) );
  NAND2_X1 U6241 ( .A1(n7030), .A2(n4411), .ZN(n7135) );
  NAND2_X1 U6242 ( .A1(n5276), .A2(n4894), .ZN(n4892) );
  NAND2_X1 U6243 ( .A1(n5579), .A2(n4898), .ZN(n4897) );
  NAND2_X1 U6244 ( .A1(n5531), .A2(n4921), .ZN(n4917) );
  NAND2_X1 U6245 ( .A1(n5128), .A2(n4931), .ZN(n4930) );
  NAND2_X1 U6246 ( .A1(n8016), .A2(n7747), .ZN(n4942) );
  NAND2_X1 U6247 ( .A1(n4942), .A2(n7749), .ZN(n4943) );
  INV_X1 U6248 ( .A(n7749), .ZN(n4944) );
  NAND3_X1 U6249 ( .A1(n5026), .A2(n5027), .A3(n5028), .ZN(n6169) );
  NAND2_X1 U6250 ( .A1(n8285), .A2(n4968), .ZN(n4965) );
  NAND2_X1 U6251 ( .A1(n4965), .A2(n4966), .ZN(n8251) );
  NAND2_X1 U6252 ( .A1(n8285), .A2(n4974), .ZN(n4972) );
  AOI22_X2 U6253 ( .A1(n4975), .A2(n5767), .B1(n7112), .B2(n4977), .ZN(n7524)
         );
  OAI21_X2 U6254 ( .B1(n7524), .B2(n5773), .A(n5772), .ZN(n7539) );
  NAND2_X1 U6255 ( .A1(n5702), .A2(n4412), .ZN(n6412) );
  AND2_X1 U6256 ( .A1(n5144), .A2(n4980), .ZN(n4979) );
  NAND2_X1 U6257 ( .A1(n5255), .A2(n5144), .ZN(n5301) );
  NAND2_X1 U6258 ( .A1(n8269), .A2(n4982), .ZN(n4981) );
  NAND2_X1 U6259 ( .A1(n4981), .A2(n4983), .ZN(n8276) );
  NAND2_X1 U6260 ( .A1(n6711), .A2(n4988), .ZN(n5728) );
  NAND2_X1 U6261 ( .A1(n6383), .A2(n6384), .ZN(n4994) );
  NAND3_X1 U6262 ( .A1(n5846), .A2(n5847), .A3(n5848), .ZN(n5875) );
  NAND3_X1 U6263 ( .A1(n8981), .A2(n8980), .A3(n8867), .ZN(n5009) );
  NOR2_X1 U6264 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5143) );
  OR2_X1 U6266 ( .A1(n5203), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U6267 ( .A1(n8525), .A2(n8524), .ZN(n8676) );
  NAND2_X1 U6268 ( .A1(n8320), .A2(n8319), .ZN(n8318) );
  XNOR2_X1 U6269 ( .A(n5801), .B(n5802), .ZN(n8320) );
  AOI21_X2 U6270 ( .B1(n7476), .B2(n5632), .A(n5016), .ZN(n7447) );
  NOR2_X2 U6271 ( .A1(n8251), .A2(n8250), .ZN(n5825) );
  INV_X1 U6272 ( .A(n6727), .ZN(n6726) );
  XNOR2_X1 U6273 ( .A(n6722), .B(n9970), .ZN(n6797) );
  OAI222_X1 U6274 ( .A1(n4374), .A2(n8249), .B1(n4385), .B2(n8248), .C1(n9242), 
        .C2(n8761), .ZN(P2_U3328) );
  AND2_X2 U6275 ( .A1(n8249), .A2(n5175), .ZN(n5323) );
  NAND2_X1 U6276 ( .A1(n9903), .A2(n6728), .ZN(n6729) );
  OR2_X1 U6277 ( .A1(n6172), .A2(n6102), .ZN(n6103) );
  NAND2_X1 U6278 ( .A1(n7700), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6173) );
  AND2_X1 U6279 ( .A1(n8856), .A2(n8855), .ZN(n8857) );
  OR2_X1 U6280 ( .A1(n6349), .A2(n6098), .ZN(n6106) );
  AND2_X1 U6281 ( .A1(n5713), .A2(n5712), .ZN(n5015) );
  NOR2_X1 U6282 ( .A1(n5631), .A2(n5630), .ZN(n5016) );
  AND4_X1 U6283 ( .A1(n5511), .A2(n5510), .A3(n5509), .A4(n5508), .ZN(n8554)
         );
  INV_X1 U6284 ( .A(n8554), .ZN(n5512) );
  INV_X1 U6285 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6468) );
  NOR2_X1 U6286 ( .A1(n7355), .A2(n5768), .ZN(n5017) );
  INV_X1 U6287 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5684) );
  AND2_X1 U6288 ( .A1(n5072), .A2(n5071), .ZN(n5019) );
  AND2_X1 U6289 ( .A1(n5065), .A2(n5064), .ZN(n5020) );
  AND4_X1 U6290 ( .A1(n7694), .A2(n7693), .A3(n7692), .A4(n7691), .ZN(n9156)
         );
  NOR2_X1 U6291 ( .A1(n7434), .A2(n7433), .ZN(n5021) );
  OR3_X1 U6292 ( .A1(n5839), .A2(n5982), .A3(n10137), .ZN(n8316) );
  AND2_X1 U6293 ( .A1(n8467), .A2(n8468), .ZN(n5022) );
  NAND2_X1 U6294 ( .A1(n6800), .A2(n6797), .ZN(n6799) );
  INV_X1 U6295 ( .A(n8609), .ZN(n5448) );
  INV_X1 U6296 ( .A(n6587), .ZN(n5621) );
  AND2_X1 U6297 ( .A1(n5826), .A2(n8321), .ZN(n5023) );
  AND4_X1 U6298 ( .A1(n5149), .A2(n5148), .A3(n5147), .A4(n5416), .ZN(n5024)
         );
  AND2_X1 U6299 ( .A1(n6935), .A2(n6892), .ZN(n6896) );
  INV_X1 U6300 ( .A(n6526), .ZN(n6522) );
  INV_X1 U6301 ( .A(n8785), .ZN(n8782) );
  INV_X1 U6302 ( .A(n7862), .ZN(n7031) );
  INV_X1 U6303 ( .A(n8249), .ZN(n5178) );
  AOI22_X1 U6304 ( .A1(n8459), .A2(n10066), .B1(n8419), .B2(n8340), .ZN(n5644)
         );
  NAND2_X1 U6305 ( .A1(n5200), .A2(n6296), .ZN(n8043) );
  XNOR2_X1 U6306 ( .A(n6258), .B(n6247), .ZN(n6260) );
  AND2_X1 U6307 ( .A1(n8846), .A2(n8845), .ZN(n8847) );
  AND2_X1 U6308 ( .A1(n6127), .A2(n5960), .ZN(n9883) );
  INV_X1 U6309 ( .A(n7753), .ZN(n6885) );
  INV_X1 U6310 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5944) );
  INV_X1 U6311 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5926) );
  INV_X1 U6312 ( .A(n8268), .ZN(n5791) );
  OR2_X1 U6313 ( .A1(n5353), .A2(n9305), .ZN(n5371) );
  INV_X1 U6314 ( .A(n8536), .ZN(n8208) );
  OR2_X1 U6315 ( .A1(n5472), .A2(n8271), .ZN(n5485) );
  OR2_X1 U6316 ( .A1(n5395), .A2(n5394), .ZN(n5424) );
  AND2_X1 U6317 ( .A1(n7460), .A2(n8101), .ZN(n7433) );
  OR2_X1 U6318 ( .A1(n5280), .A2(n6774), .ZN(n5295) );
  NAND2_X1 U6319 ( .A1(n10064), .A2(n10105), .ZN(n8047) );
  INV_X1 U6320 ( .A(n6633), .ZN(n6632) );
  INV_X1 U6321 ( .A(n7065), .ZN(n7066) );
  NOR2_X1 U6322 ( .A1(n7655), .A2(n8958), .ZN(n7668) );
  OR2_X1 U6323 ( .A1(n7622), .A2(n9004), .ZN(n7632) );
  OR2_X1 U6324 ( .A1(n6823), .A2(n6822), .ZN(n6997) );
  INV_X1 U6325 ( .A(n9156), .ZN(n7695) );
  AND2_X1 U6326 ( .A1(n7423), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7492) );
  INV_X1 U6327 ( .A(n7865), .ZN(n7396) );
  NOR2_X1 U6328 ( .A1(n9154), .A2(n9155), .ZN(n9153) );
  NAND2_X1 U6329 ( .A1(n5056), .A2(n5055), .ZN(n5059) );
  XNOR2_X1 U6330 ( .A(n8503), .B(n5816), .ZN(n8296) );
  NAND2_X1 U6331 ( .A1(n5323), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5184) );
  OR2_X1 U6332 ( .A1(n5779), .A2(n5778), .ZN(n5780) );
  AND2_X1 U6333 ( .A1(n8217), .A2(n8024), .ZN(n8220) );
  AND4_X1 U6334 ( .A1(n5501), .A2(n5500), .A3(n5499), .A4(n5498), .ZN(n8308)
         );
  OR2_X1 U6335 ( .A1(n5194), .A2(n5232), .ZN(n5236) );
  AND2_X1 U6336 ( .A1(n8059), .A2(n8058), .ZN(n8185) );
  OR2_X1 U6337 ( .A1(n5831), .A2(n5829), .ZN(n8604) );
  INV_X1 U6338 ( .A(n6296), .ZN(n10075) );
  INV_X1 U6339 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5657) );
  INV_X1 U6340 ( .A(n9172), .ZN(n9031) );
  INV_X1 U6341 ( .A(n9057), .ZN(n9481) );
  INV_X1 U6342 ( .A(n9651), .ZN(n9553) );
  INV_X1 U6343 ( .A(n9669), .ZN(n7481) );
  AOI21_X1 U6344 ( .B1(n7407), .B2(n9060), .A(n7393), .ZN(n7411) );
  INV_X1 U6345 ( .A(n9063), .ZN(n7046) );
  AND2_X1 U6346 ( .A1(n5106), .A2(n5105), .ZN(n5414) );
  NAND2_X1 U6347 ( .A1(n5046), .A2(SI_5_), .ZN(n5047) );
  NAND2_X1 U6348 ( .A1(n5040), .A2(SI_3_), .ZN(n5041) );
  NAND2_X1 U6349 ( .A1(n5190), .A2(n5189), .ZN(n5033) );
  AND4_X1 U6350 ( .A1(n5447), .A2(n5446), .A3(n5445), .A4(n5444), .ZN(n8623)
         );
  INV_X1 U6351 ( .A(n10055), .ZN(n9744) );
  NOR2_X1 U6352 ( .A1(n8498), .A2(n8505), .ZN(n8499) );
  AND2_X1 U6353 ( .A1(n8139), .A2(n8137), .ZN(n8566) );
  AND2_X1 U6354 ( .A1(n5640), .A2(n5982), .ZN(n10066) );
  INV_X1 U6355 ( .A(n8185), .ZN(n6759) );
  INV_X1 U6356 ( .A(n8622), .ZN(n10065) );
  OR2_X1 U6357 ( .A1(n5650), .A2(n5690), .ZN(n10155) );
  AND2_X1 U6358 ( .A1(n8570), .A2(n8569), .ZN(n8695) );
  AND2_X1 U6359 ( .A1(n8630), .A2(n10142), .ZN(n10132) );
  AND2_X1 U6360 ( .A1(n5863), .A2(n10094), .ZN(n10081) );
  AND4_X1 U6361 ( .A1(n7707), .A2(n7706), .A3(n7705), .A4(n7704), .ZN(n9134)
         );
  OR2_X1 U6362 ( .A1(n6349), .A2(n6945), .ZN(n6505) );
  OR2_X1 U6363 ( .A1(n7703), .A2(n6348), .ZN(n6355) );
  NAND2_X1 U6364 ( .A1(n7943), .A2(n7910), .ZN(n9136) );
  NAND2_X1 U6365 ( .A1(n7946), .A2(n7825), .ZN(n9185) );
  NAND2_X1 U6366 ( .A1(n7802), .A2(n7932), .ZN(n9557) );
  AND2_X1 U6367 ( .A1(n9573), .A2(n10005), .ZN(n9909) );
  AND2_X1 U6368 ( .A1(n6177), .A2(n6232), .ZN(n10005) );
  XNOR2_X1 U6369 ( .A(n5053), .B(SI_7_), .ZN(n5289) );
  NOR2_X1 U6370 ( .A1(n9720), .A2(n10227), .ZN(n9721) );
  AND3_X1 U6371 ( .A1(n5602), .A2(n5601), .A3(n5600), .ZN(n8442) );
  AND2_X1 U6372 ( .A1(n6033), .A2(n6032), .ZN(n8417) );
  INV_X1 U6373 ( .A(n10177), .ZN(n10175) );
  INV_X1 U6374 ( .A(n10163), .ZN(n10161) );
  INV_X1 U6375 ( .A(n5650), .ZN(n8218) );
  INV_X1 U6376 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6089) );
  INV_X1 U6377 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6075) );
  INV_X1 U6378 ( .A(n8774), .ZN(n9768) );
  INV_X1 U6379 ( .A(n9201), .ZN(n9625) );
  OR2_X1 U6380 ( .A1(n6233), .A2(n6374), .ZN(n9052) );
  INV_X1 U6381 ( .A(n9128), .ZN(n9763) );
  NAND2_X1 U6382 ( .A1(n6235), .A2(n9691), .ZN(n9936) );
  INV_X1 U6383 ( .A(n10049), .ZN(n10047) );
  INV_X1 U6384 ( .A(n10037), .ZN(n10035) );
  INV_X1 U6385 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9302) );
  INV_X1 U6386 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6510) );
  INV_X1 U6387 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6078) );
  NOR2_X1 U6388 ( .A1(n10184), .A2(n10183), .ZN(n10182) );
  NOR2_X1 U6389 ( .A1(n10211), .A2(n10210), .ZN(n10209) );
  NOR2_X1 U6390 ( .A1(n10208), .A2(n10207), .ZN(n10206) );
  AND2_X1 U6391 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5028) );
  INV_X1 U6392 ( .A(SI_1_), .ZN(n5030) );
  MUX2_X1 U6393 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5038), .Z(n5189) );
  NAND2_X1 U6394 ( .A1(n5031), .A2(SI_1_), .ZN(n5032) );
  MUX2_X1 U6395 ( .A(n6075), .B(n6078), .S(n5038), .Z(n5034) );
  NAND2_X1 U6396 ( .A1(n5212), .A2(n5211), .ZN(n5037) );
  INV_X1 U6397 ( .A(n5034), .ZN(n5035) );
  INV_X1 U6398 ( .A(n5039), .ZN(n5040) );
  NAND2_X1 U6399 ( .A1(n5042), .A2(SI_4_), .ZN(n5043) );
  INV_X1 U6400 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5044) );
  INV_X8 U6401 ( .A(n6251), .ZN(n7743) );
  MUX2_X1 U6402 ( .A(n6087), .B(n5044), .S(n7743), .Z(n5045) );
  NAND2_X1 U6403 ( .A1(n5257), .A2(n5256), .ZN(n5048) );
  INV_X1 U6404 ( .A(n5045), .ZN(n5046) );
  INV_X1 U6405 ( .A(n5049), .ZN(n5050) );
  NAND2_X1 U6406 ( .A1(n5050), .A2(SI_6_), .ZN(n5051) );
  INV_X1 U6407 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6092) );
  INV_X1 U6408 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5052) );
  MUX2_X1 U6409 ( .A(n6092), .B(n5052), .S(n7743), .Z(n5053) );
  INV_X1 U6410 ( .A(n5053), .ZN(n5054) );
  INV_X1 U6411 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6093) );
  MUX2_X1 U6412 ( .A(n6093), .B(n9302), .S(n7743), .Z(n5056) );
  INV_X1 U6413 ( .A(SI_8_), .ZN(n5055) );
  INV_X1 U6414 ( .A(n5056), .ZN(n5057) );
  NAND2_X1 U6415 ( .A1(n5057), .A2(SI_8_), .ZN(n5058) );
  INV_X1 U6416 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6120) );
  INV_X1 U6417 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5060) );
  INV_X1 U6418 ( .A(SI_9_), .ZN(n5061) );
  INV_X1 U6419 ( .A(n5062), .ZN(n5063) );
  NAND2_X1 U6420 ( .A1(n5063), .A2(SI_9_), .ZN(n5064) );
  INV_X1 U6421 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5067) );
  INV_X1 U6422 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5066) );
  MUX2_X1 U6423 ( .A(n5067), .B(n5066), .S(n7743), .Z(n5069) );
  INV_X1 U6424 ( .A(SI_10_), .ZN(n5068) );
  INV_X1 U6425 ( .A(n5069), .ZN(n5070) );
  NAND2_X1 U6426 ( .A1(n5070), .A2(SI_10_), .ZN(n5071) );
  INV_X1 U6427 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6137) );
  INV_X1 U6428 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9329) );
  MUX2_X1 U6429 ( .A(n6137), .B(n9329), .S(n7743), .Z(n5073) );
  INV_X1 U6430 ( .A(n5073), .ZN(n5074) );
  NAND2_X1 U6431 ( .A1(n5074), .A2(SI_11_), .ZN(n5075) );
  INV_X1 U6432 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9440) );
  INV_X1 U6433 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5077) );
  INV_X1 U6434 ( .A(SI_12_), .ZN(n5078) );
  NAND2_X1 U6435 ( .A1(n5079), .A2(n5078), .ZN(n5361) );
  INV_X1 U6436 ( .A(n5079), .ZN(n5080) );
  NAND2_X1 U6437 ( .A1(n5080), .A2(SI_12_), .ZN(n5081) );
  NAND2_X1 U6438 ( .A1(n5361), .A2(n5081), .ZN(n5359) );
  INV_X1 U6439 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n5083) );
  INV_X1 U6440 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5082) );
  MUX2_X1 U6441 ( .A(n5083), .B(n5082), .S(n7743), .Z(n5085) );
  INV_X1 U6442 ( .A(SI_13_), .ZN(n5084) );
  NAND2_X1 U6443 ( .A1(n5085), .A2(n5084), .ZN(n5089) );
  INV_X1 U6444 ( .A(n5085), .ZN(n5086) );
  NAND2_X1 U6445 ( .A1(n5086), .A2(SI_13_), .ZN(n5087) );
  NAND2_X1 U6446 ( .A1(n5089), .A2(n5087), .ZN(n5363) );
  INV_X1 U6447 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n5092) );
  INV_X1 U6448 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6204) );
  MUX2_X1 U6449 ( .A(n5092), .B(n6204), .S(n7743), .Z(n5094) );
  XNOR2_X1 U6450 ( .A(n5094), .B(SI_14_), .ZN(n5384) );
  INV_X1 U6451 ( .A(n5094), .ZN(n5095) );
  NAND2_X1 U6452 ( .A1(n5095), .A2(SI_14_), .ZN(n5096) );
  INV_X1 U6453 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6311) );
  INV_X1 U6454 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6309) );
  MUX2_X1 U6455 ( .A(n6311), .B(n6309), .S(n7743), .Z(n5098) );
  INV_X1 U6456 ( .A(SI_15_), .ZN(n5097) );
  NAND2_X1 U6457 ( .A1(n5098), .A2(n5097), .ZN(n5101) );
  INV_X1 U6458 ( .A(n5098), .ZN(n5099) );
  NAND2_X1 U6459 ( .A1(n5099), .A2(SI_15_), .ZN(n5100) );
  NAND2_X1 U6460 ( .A1(n5101), .A2(n5100), .ZN(n5403) );
  INV_X1 U6461 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9288) );
  INV_X1 U6462 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6290) );
  MUX2_X1 U6463 ( .A(n9288), .B(n6290), .S(n7743), .Z(n5103) );
  INV_X1 U6464 ( .A(SI_16_), .ZN(n5102) );
  NAND2_X1 U6465 ( .A1(n5103), .A2(n5102), .ZN(n5106) );
  INV_X1 U6466 ( .A(n5103), .ZN(n5104) );
  NAND2_X1 U6467 ( .A1(n5104), .A2(SI_16_), .ZN(n5105) );
  NAND2_X1 U6468 ( .A1(n5107), .A2(n5106), .ZN(n5434) );
  INV_X1 U6469 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5109) );
  INV_X1 U6470 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5108) );
  MUX2_X1 U6471 ( .A(n5109), .B(n5108), .S(n7743), .Z(n5110) );
  XNOR2_X1 U6472 ( .A(n5110), .B(SI_17_), .ZN(n5433) );
  INV_X1 U6473 ( .A(n5433), .ZN(n5113) );
  INV_X1 U6474 ( .A(n5110), .ZN(n5111) );
  NAND2_X1 U6475 ( .A1(n5111), .A2(SI_17_), .ZN(n5112) );
  MUX2_X1 U6476 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7743), .Z(n5115) );
  XNOR2_X1 U6477 ( .A(n5115), .B(SI_18_), .ZN(n5450) );
  INV_X1 U6478 ( .A(n5450), .ZN(n5114) );
  NAND2_X1 U6479 ( .A1(n5451), .A2(n5114), .ZN(n5117) );
  NAND2_X1 U6480 ( .A1(n5115), .A2(SI_18_), .ZN(n5116) );
  NAND2_X1 U6481 ( .A1(n5117), .A2(n5116), .ZN(n5463) );
  INV_X1 U6482 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n9221) );
  INV_X1 U6483 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6555) );
  MUX2_X1 U6484 ( .A(n9221), .B(n6555), .S(n7743), .Z(n5119) );
  INV_X1 U6485 ( .A(SI_19_), .ZN(n5118) );
  NAND2_X1 U6486 ( .A1(n5119), .A2(n5118), .ZN(n5122) );
  INV_X1 U6487 ( .A(n5119), .ZN(n5120) );
  NAND2_X1 U6488 ( .A1(n5120), .A2(SI_19_), .ZN(n5121) );
  NAND2_X1 U6489 ( .A1(n5122), .A2(n5121), .ZN(n5462) );
  INV_X1 U6490 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6720) );
  INV_X1 U6491 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8007) );
  MUX2_X1 U6492 ( .A(n6720), .B(n8007), .S(n7743), .Z(n5124) );
  INV_X1 U6493 ( .A(SI_20_), .ZN(n5123) );
  NAND2_X1 U6494 ( .A1(n5124), .A2(n5123), .ZN(n5127) );
  INV_X1 U6495 ( .A(n5124), .ZN(n5125) );
  NAND2_X1 U6496 ( .A1(n5125), .A2(SI_20_), .ZN(n5126) );
  AND2_X1 U6497 ( .A1(n5127), .A2(n5126), .ZN(n5480) );
  NAND2_X1 U6498 ( .A1(n5481), .A2(n5480), .ZN(n5128) );
  MUX2_X1 U6499 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7743), .Z(n5130) );
  INV_X1 U6500 ( .A(SI_21_), .ZN(n5129) );
  XNOR2_X1 U6501 ( .A(n5130), .B(n5129), .ZN(n5492) );
  NAND2_X1 U6502 ( .A1(n5130), .A2(SI_21_), .ZN(n5131) );
  INV_X1 U6503 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n9358) );
  INV_X1 U6504 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7017) );
  MUX2_X1 U6505 ( .A(n9358), .B(n7017), .S(n7743), .Z(n5133) );
  INV_X1 U6506 ( .A(SI_22_), .ZN(n5132) );
  NAND2_X1 U6507 ( .A1(n5133), .A2(n5132), .ZN(n5136) );
  INV_X1 U6508 ( .A(n5133), .ZN(n5134) );
  NAND2_X1 U6509 ( .A1(n5134), .A2(SI_22_), .ZN(n5135) );
  NAND2_X1 U6510 ( .A1(n5136), .A2(n5135), .ZN(n5502) );
  INV_X1 U6511 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7079) );
  INV_X1 U6512 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5137) );
  MUX2_X1 U6513 ( .A(n7079), .B(n5137), .S(n7743), .Z(n5138) );
  INV_X1 U6514 ( .A(SI_23_), .ZN(n9448) );
  NAND2_X1 U6515 ( .A1(n5138), .A2(n9448), .ZN(n5141) );
  INV_X1 U6516 ( .A(n5138), .ZN(n5139) );
  NAND2_X1 U6517 ( .A1(n5139), .A2(SI_23_), .ZN(n5140) );
  AND2_X1 U6518 ( .A1(n5141), .A2(n5140), .ZN(n5514) );
  NAND2_X1 U6519 ( .A1(n5515), .A2(n5514), .ZN(n5517) );
  MUX2_X1 U6520 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7743), .Z(n5529) );
  INV_X1 U6521 ( .A(SI_24_), .ZN(n5142) );
  XNOR2_X1 U6522 ( .A(n5529), .B(n5142), .ZN(n5528) );
  NAND2_X1 U6523 ( .A1(n5186), .A2(n5143), .ZN(n5237) );
  NOR2_X2 U6524 ( .A1(n5237), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5255) );
  NOR3_X1 U6525 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .A3(
        P2_IR_REG_17__SCAN_IN), .ZN(n5149) );
  INV_X1 U6526 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5386) );
  INV_X1 U6527 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5146) );
  INV_X1 U6528 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5145) );
  NOR2_X1 U6529 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5147) );
  NOR2_X1 U6530 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5416) );
  INV_X1 U6531 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5151) );
  NOR2_X1 U6532 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5152) );
  INV_X1 U6533 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5153) );
  INV_X1 U6534 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5154) );
  INV_X1 U6535 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6536 ( .A1(n7642), .A2(n8015), .ZN(n5156) );
  INV_X1 U6537 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7125) );
  OR2_X1 U6538 ( .A1(n5569), .A2(n7125), .ZN(n5155) );
  NAND2_X1 U6539 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5248) );
  INV_X1 U6540 ( .A(n5248), .ZN(n5157) );
  NAND2_X1 U6541 ( .A1(n5157), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5263) );
  INV_X1 U6542 ( .A(n5263), .ZN(n5158) );
  NAND2_X1 U6543 ( .A1(n5158), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5280) );
  INV_X1 U6544 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6774) );
  INV_X1 U6545 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5294) );
  INV_X1 U6546 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9328) );
  INV_X1 U6547 ( .A(n5336), .ZN(n5160) );
  AND2_X1 U6548 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n5159) );
  NAND2_X1 U6549 ( .A1(n5160), .A2(n5159), .ZN(n5353) );
  INV_X1 U6550 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9305) );
  INV_X1 U6551 ( .A(n5371), .ZN(n5161) );
  NAND2_X1 U6552 ( .A1(n5161), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5395) );
  INV_X1 U6553 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5394) );
  INV_X1 U6554 ( .A(n5424), .ZN(n5163) );
  AND2_X1 U6555 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n5162) );
  NAND2_X1 U6556 ( .A1(n5163), .A2(n5162), .ZN(n5442) );
  INV_X1 U6557 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7518) );
  INV_X1 U6558 ( .A(n5455), .ZN(n5164) );
  NAND2_X1 U6559 ( .A1(n5164), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5472) );
  INV_X1 U6560 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8271) );
  INV_X1 U6561 ( .A(n5485), .ZN(n5165) );
  NAND2_X1 U6562 ( .A1(n5165), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5496) );
  INV_X1 U6563 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9451) );
  NAND2_X1 U6564 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n5166) );
  NAND2_X1 U6565 ( .A1(n5167), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5552) );
  INV_X1 U6566 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9460) );
  NAND2_X1 U6567 ( .A1(n5522), .A2(n9460), .ZN(n5168) );
  NAND2_X1 U6568 ( .A1(n5552), .A2(n5168), .ZN(n8500) );
  INV_X1 U6569 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5171) );
  XNOR2_X2 U6570 ( .A(n5172), .B(n5171), .ZN(n8249) );
  NAND2_X1 U6571 ( .A1(n5173), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5174) );
  XNOR2_X1 U6572 ( .A(n5174), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5175) );
  INV_X1 U6573 ( .A(n5175), .ZN(n8763) );
  OR2_X2 U6574 ( .A1(n8249), .A2(n8763), .ZN(n5203) );
  INV_X1 U6575 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9425) );
  OR2_X1 U6576 ( .A1(n6186), .A2(n9425), .ZN(n5177) );
  NAND2_X1 U6577 ( .A1(n8249), .A2(n8763), .ZN(n5194) );
  NAND2_X1 U6578 ( .A1(n5204), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5176) );
  AND2_X1 U6579 ( .A1(n5177), .A2(n5176), .ZN(n5180) );
  NAND2_X1 U6580 ( .A1(n5206), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5179) );
  OAI211_X1 U6581 ( .C1(n8500), .C2(n5203), .A(n5180), .B(n5179), .ZN(n8342)
         );
  INV_X1 U6582 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9453) );
  OR2_X1 U6583 ( .A1(n5203), .A2(n9453), .ZN(n5183) );
  OR2_X1 U6584 ( .A1(n4379), .A2(n4949), .ZN(n5182) );
  NAND2_X1 U6585 ( .A1(n5204), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5181) );
  NAND2_X1 U6586 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5185) );
  MUX2_X1 U6587 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5185), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5188) );
  INV_X1 U6588 ( .A(n5186), .ZN(n5187) );
  INV_X1 U6589 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6073) );
  XNOR2_X1 U6590 ( .A(n5190), .B(n5189), .ZN(n6255) );
  OR2_X1 U6591 ( .A1(n4396), .A2(n6255), .ZN(n5192) );
  INV_X1 U6592 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5193) );
  OR2_X1 U6593 ( .A1(n5194), .A2(n5193), .ZN(n5198) );
  NAND2_X1 U6594 ( .A1(n5323), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5197) );
  INV_X1 U6595 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6404) );
  OR2_X1 U6596 ( .A1(n5203), .A2(n6404), .ZN(n5196) );
  INV_X1 U6597 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10054) );
  OR2_X1 U6598 ( .A1(n4380), .A2(n10054), .ZN(n5195) );
  NAND2_X1 U6599 ( .A1(n4498), .A2(SI_0_), .ZN(n5199) );
  XNOR2_X1 U6600 ( .A(n5199), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U6601 ( .A1(n10067), .A2(n10096), .ZN(n10072) );
  NAND2_X1 U6602 ( .A1(n8186), .A2(n10072), .ZN(n5202) );
  NAND2_X1 U6603 ( .A1(n5200), .A2(n10075), .ZN(n5201) );
  NAND2_X1 U6604 ( .A1(n5202), .A2(n5201), .ZN(n6453) );
  NAND2_X1 U6605 ( .A1(n5323), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5209) );
  NAND2_X1 U6606 ( .A1(n5204), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5208) );
  OR2_X1 U6607 ( .A1(n5240), .A2(n6075), .ZN(n5217) );
  XNOR2_X1 U6608 ( .A(n5211), .B(n5212), .ZN(n6271) );
  OR2_X1 U6609 ( .A1(n5191), .A2(n6271), .ZN(n5216) );
  OR2_X1 U6610 ( .A1(n5186), .A2(n5657), .ZN(n5214) );
  INV_X1 U6611 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5213) );
  XNOR2_X1 U6612 ( .A(n5214), .B(n5213), .ZN(n6074) );
  OR2_X1 U6613 ( .A1(n4399), .A2(n6074), .ZN(n5215) );
  NAND2_X1 U6614 ( .A1(n8044), .A2(n8047), .ZN(n8187) );
  NAND2_X1 U6615 ( .A1(n6453), .A2(n8187), .ZN(n5219) );
  INV_X1 U6616 ( .A(n10105), .ZN(n6458) );
  OR2_X1 U6617 ( .A1(n10064), .A2(n6458), .ZN(n5218) );
  NAND2_X1 U6618 ( .A1(n5219), .A2(n5218), .ZN(n6420) );
  NAND2_X1 U6619 ( .A1(n5323), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5224) );
  INV_X1 U6620 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5220) );
  OR2_X1 U6621 ( .A1(n5194), .A2(n5220), .ZN(n5223) );
  INV_X1 U6622 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6429) );
  OR2_X1 U6623 ( .A1(n5205), .A2(n6429), .ZN(n5221) );
  NAND2_X1 U6624 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4443), .ZN(n5225) );
  XNOR2_X1 U6625 ( .A(n5225), .B(P2_IR_REG_3__SCAN_IN), .ZN(n5998) );
  INV_X1 U6626 ( .A(n5998), .ZN(n6080) );
  OR2_X1 U6627 ( .A1(n4397), .A2(n6081), .ZN(n5229) );
  XNOR2_X1 U6628 ( .A(n5227), .B(n5226), .ZN(n6339) );
  OAI211_X1 U6629 ( .C1(n4398), .C2(n6080), .A(n5229), .B(n5228), .ZN(n6433)
         );
  NAND2_X1 U6630 ( .A1(n6604), .A2(n6433), .ZN(n6599) );
  NAND2_X1 U6631 ( .A1(n6420), .A2(n6423), .ZN(n5231) );
  NAND2_X1 U6632 ( .A1(n6604), .A2(n4384), .ZN(n5230) );
  NAND2_X1 U6633 ( .A1(n5231), .A2(n5230), .ZN(n6595) );
  INV_X1 U6634 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5232) );
  INV_X1 U6635 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6002) );
  OR2_X1 U6636 ( .A1(n6186), .A2(n6002), .ZN(n5235) );
  OAI21_X1 U6637 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5248), .ZN(n6596) );
  OR2_X1 U6638 ( .A1(n5203), .A2(n6596), .ZN(n5234) );
  INV_X1 U6639 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5969) );
  OR2_X1 U6640 ( .A1(n5205), .A2(n5969), .ZN(n5233) );
  NAND2_X1 U6641 ( .A1(n5237), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5239) );
  INV_X1 U6642 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5238) );
  XNOR2_X1 U6643 ( .A(n5239), .B(n5238), .ZN(n6082) );
  INV_X1 U6644 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6083) );
  OR2_X1 U6645 ( .A1(n4397), .A2(n6083), .ZN(n5244) );
  XNOR2_X1 U6646 ( .A(n5241), .B(n5242), .ZN(n6359) );
  OR2_X1 U6647 ( .A1(n5191), .A2(n6359), .ZN(n5243) );
  OAI211_X1 U6648 ( .C1(n6031), .C2(n6082), .A(n5244), .B(n5243), .ZN(n10116)
         );
  NAND2_X1 U6649 ( .A1(n6550), .A2(n10116), .ZN(n8029) );
  NAND2_X1 U6650 ( .A1(n8356), .A2(n4383), .ZN(n8028) );
  NAND2_X1 U6651 ( .A1(n8029), .A2(n8028), .ZN(n6601) );
  NAND2_X1 U6652 ( .A1(n6550), .A2(n4383), .ZN(n5245) );
  NAND2_X1 U6653 ( .A1(n5206), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5254) );
  INV_X1 U6654 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5246) );
  OR2_X1 U6655 ( .A1(n5194), .A2(n5246), .ZN(n5253) );
  INV_X1 U6656 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U6657 ( .A1(n5248), .A2(n5247), .ZN(n5249) );
  NAND2_X1 U6658 ( .A1(n5263), .A2(n5249), .ZN(n6551) );
  OR2_X1 U6659 ( .A1(n5203), .A2(n6551), .ZN(n5252) );
  INV_X1 U6660 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5250) );
  OR2_X1 U6661 ( .A1(n6186), .A2(n5250), .ZN(n5251) );
  OR2_X1 U6662 ( .A1(n5255), .A2(n5657), .ZN(n5270) );
  XNOR2_X1 U6663 ( .A(n5270), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6661) );
  INV_X1 U6664 ( .A(n6661), .ZN(n6086) );
  XNOR2_X1 U6665 ( .A(n5257), .B(n5256), .ZN(n6486) );
  OR2_X1 U6666 ( .A1(n5191), .A2(n6486), .ZN(n5259) );
  OR2_X1 U6667 ( .A1(n5240), .A2(n6087), .ZN(n5258) );
  OAI211_X1 U6668 ( .C1(n6031), .C2(n6086), .A(n5259), .B(n5258), .ZN(n6584)
         );
  INV_X1 U6669 ( .A(n6584), .ZN(n10125) );
  AND2_X1 U6670 ( .A1(n6762), .A2(n10125), .ZN(n5261) );
  NAND2_X1 U6671 ( .A1(n6762), .A2(n6584), .ZN(n8033) );
  INV_X1 U6672 ( .A(n6762), .ZN(n8355) );
  NAND2_X1 U6673 ( .A1(n8355), .A2(n10125), .ZN(n8052) );
  NAND2_X1 U6674 ( .A1(n8033), .A2(n8052), .ZN(n6587) );
  OR2_X1 U6675 ( .A1(n6587), .A2(n10125), .ZN(n5260) );
  NAND2_X1 U6676 ( .A1(n5204), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5268) );
  INV_X1 U6677 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6005) );
  OR2_X1 U6678 ( .A1(n6186), .A2(n6005), .ZN(n5267) );
  INV_X1 U6679 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6680 ( .A1(n5263), .A2(n5262), .ZN(n5264) );
  NAND2_X1 U6681 ( .A1(n5280), .A2(n5264), .ZN(n6768) );
  OR2_X1 U6682 ( .A1(n5203), .A2(n6768), .ZN(n5266) );
  INV_X1 U6683 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6765) );
  OR2_X1 U6684 ( .A1(n4380), .A2(n6765), .ZN(n5265) );
  INV_X1 U6685 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U6686 ( .A1(n5270), .A2(n5269), .ZN(n5271) );
  NAND2_X1 U6687 ( .A1(n5271), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5273) );
  INV_X1 U6688 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6689 ( .A1(n5273), .A2(n5272), .ZN(n5287) );
  OR2_X1 U6690 ( .A1(n5273), .A2(n5272), .ZN(n5274) );
  NAND2_X1 U6691 ( .A1(n5287), .A2(n5274), .ZN(n6088) );
  XNOR2_X1 U6692 ( .A(n5276), .B(n5275), .ZN(n6508) );
  OR2_X1 U6693 ( .A1(n4503), .A2(n6508), .ZN(n5278) );
  OR2_X1 U6694 ( .A1(n5569), .A2(n6089), .ZN(n5277) );
  OAI211_X1 U6695 ( .C1(n6031), .C2(n6088), .A(n5278), .B(n5277), .ZN(n10128)
         );
  NAND2_X1 U6696 ( .A1(n6841), .A2(n10128), .ZN(n8059) );
  INV_X1 U6697 ( .A(n6841), .ZN(n8354) );
  NAND2_X1 U6698 ( .A1(n8354), .A2(n4513), .ZN(n8058) );
  NOR2_X1 U6699 ( .A1(n6841), .A2(n4513), .ZN(n5279) );
  NAND2_X1 U6700 ( .A1(n5204), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5286) );
  INV_X1 U6701 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9464) );
  OR2_X1 U6702 ( .A1(n4380), .A2(n9464), .ZN(n5285) );
  NAND2_X1 U6703 ( .A1(n5280), .A2(n6774), .ZN(n5281) );
  NAND2_X1 U6704 ( .A1(n5295), .A2(n5281), .ZN(n6846) );
  OR2_X1 U6705 ( .A1(n5203), .A2(n6846), .ZN(n5284) );
  INV_X1 U6706 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5282) );
  OR2_X1 U6707 ( .A1(n6186), .A2(n5282), .ZN(n5283) );
  NAND2_X1 U6708 ( .A1(n5287), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5288) );
  XNOR2_X1 U6709 ( .A(n5288), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6007) );
  INV_X1 U6710 ( .A(n6007), .ZN(n6091) );
  XNOR2_X1 U6711 ( .A(n5290), .B(n5289), .ZN(n6474) );
  OR2_X1 U6712 ( .A1(n4503), .A2(n6474), .ZN(n5292) );
  OR2_X1 U6713 ( .A1(n5569), .A2(n6092), .ZN(n5291) );
  OAI211_X1 U6714 ( .C1(n6031), .C2(n6091), .A(n5292), .B(n5291), .ZN(n7008)
         );
  NAND2_X1 U6715 ( .A1(n7081), .A2(n7008), .ZN(n8074) );
  INV_X1 U6716 ( .A(n7081), .ZN(n8353) );
  INV_X1 U6717 ( .A(n7008), .ZN(n6847) );
  NAND2_X1 U6718 ( .A1(n8353), .A2(n6847), .ZN(n5624) );
  NAND2_X1 U6719 ( .A1(n8074), .A2(n5624), .ZN(n8060) );
  NAND2_X1 U6720 ( .A1(n7081), .A2(n6847), .ZN(n5293) );
  NAND2_X1 U6721 ( .A1(n5204), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5300) );
  INV_X1 U6722 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7090) );
  OR2_X1 U6723 ( .A1(n4380), .A2(n7090), .ZN(n5299) );
  NAND2_X1 U6724 ( .A1(n5295), .A2(n5294), .ZN(n5296) );
  NAND2_X1 U6725 ( .A1(n5312), .A2(n5296), .ZN(n7093) );
  OR2_X1 U6726 ( .A1(n5203), .A2(n7093), .ZN(n5298) );
  INV_X1 U6727 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6008) );
  OR2_X1 U6728 ( .A1(n6186), .A2(n6008), .ZN(n5297) );
  NAND2_X1 U6729 ( .A1(n5301), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5303) );
  INV_X1 U6730 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5302) );
  XNOR2_X1 U6731 ( .A(n5303), .B(n5302), .ZN(n6621) );
  INV_X1 U6732 ( .A(n5304), .ZN(n5305) );
  XNOR2_X1 U6733 ( .A(n5306), .B(n5305), .ZN(n6626) );
  OR2_X1 U6734 ( .A1(n4503), .A2(n6626), .ZN(n5308) );
  OR2_X1 U6735 ( .A1(n5569), .A2(n6093), .ZN(n5307) );
  OAI211_X1 U6736 ( .C1(n6031), .C2(n6621), .A(n5308), .B(n5307), .ZN(n10136)
         );
  NAND2_X1 U6737 ( .A1(n7118), .A2(n10136), .ZN(n8063) );
  INV_X1 U6738 ( .A(n10136), .ZN(n7094) );
  NAND2_X1 U6739 ( .A1(n8352), .A2(n7094), .ZN(n8027) );
  NAND2_X1 U6740 ( .A1(n8063), .A2(n8027), .ZN(n8192) );
  INV_X1 U6741 ( .A(n8192), .ZN(n5310) );
  NAND2_X1 U6742 ( .A1(n8352), .A2(n10136), .ZN(n5309) );
  NAND2_X1 U6743 ( .A1(n5204), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5317) );
  INV_X1 U6744 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5311) );
  OR2_X1 U6745 ( .A1(n4380), .A2(n5311), .ZN(n5316) );
  NAND2_X1 U6746 ( .A1(n5312), .A2(n9328), .ZN(n5313) );
  NAND2_X1 U6747 ( .A1(n5336), .A2(n5313), .ZN(n7116) );
  OR2_X1 U6748 ( .A1(n5203), .A2(n7116), .ZN(n5315) );
  INV_X1 U6749 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6011) );
  OR2_X1 U6750 ( .A1(n6186), .A2(n6011), .ZN(n5314) );
  NAND2_X1 U6751 ( .A1(n4470), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5318) );
  XNOR2_X1 U6752 ( .A(n5318), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6709) );
  INV_X1 U6753 ( .A(n6709), .ZN(n6118) );
  XNOR2_X1 U6754 ( .A(n5319), .B(n5020), .ZN(n6814) );
  NAND2_X1 U6755 ( .A1(n6814), .A2(n8015), .ZN(n5321) );
  OR2_X1 U6756 ( .A1(n5569), .A2(n6120), .ZN(n5320) );
  OAI211_X1 U6757 ( .C1(n6031), .C2(n6118), .A(n5321), .B(n5320), .ZN(n7155)
         );
  NAND2_X1 U6758 ( .A1(n7243), .A2(n7155), .ZN(n8067) );
  INV_X1 U6759 ( .A(n7243), .ZN(n8351) );
  INV_X1 U6760 ( .A(n7155), .ZN(n7207) );
  NAND2_X1 U6761 ( .A1(n8351), .A2(n7207), .ZN(n8069) );
  NAND2_X1 U6762 ( .A1(n7243), .A2(n7207), .ZN(n5322) );
  NAND2_X1 U6763 ( .A1(n5323), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5328) );
  INV_X1 U6764 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5324) );
  OR2_X1 U6765 ( .A1(n5194), .A2(n5324), .ZN(n5327) );
  INV_X1 U6766 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5335) );
  XNOR2_X1 U6767 ( .A(n5336), .B(n5335), .ZN(n7247) );
  OR2_X1 U6768 ( .A1(n5203), .A2(n7247), .ZN(n5326) );
  INV_X1 U6769 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7248) );
  OR2_X1 U6770 ( .A1(n4380), .A2(n7248), .ZN(n5325) );
  XNOR2_X1 U6771 ( .A(n5329), .B(n5019), .ZN(n6986) );
  NAND2_X1 U6772 ( .A1(n6986), .A2(n8015), .ZN(n5332) );
  NAND2_X1 U6773 ( .A1(n5345), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5330) );
  XNOR2_X1 U6774 ( .A(n5330), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6673) );
  AOI22_X1 U6775 ( .A1(n5469), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5468), .B2(
        n6673), .ZN(n5331) );
  NAND2_X1 U6776 ( .A1(n5332), .A2(n5331), .ZN(n7251) );
  INV_X1 U6777 ( .A(n5625), .ZN(n7241) );
  NAND2_X1 U6778 ( .A1(n5333), .A2(n5625), .ZN(n7237) );
  NAND2_X1 U6779 ( .A1(n8350), .A2(n7251), .ZN(n7369) );
  NAND2_X1 U6780 ( .A1(n5323), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5342) );
  INV_X1 U6781 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9465) );
  OR2_X1 U6782 ( .A1(n5194), .A2(n9465), .ZN(n5341) );
  INV_X1 U6783 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5334) );
  OAI21_X1 U6784 ( .B1(n5336), .B2(n5335), .A(n5334), .ZN(n5337) );
  NAND2_X1 U6785 ( .A1(n5337), .A2(n5353), .ZN(n7373) );
  OR2_X1 U6786 ( .A1(n5203), .A2(n7373), .ZN(n5340) );
  INV_X1 U6787 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5338) );
  OR2_X1 U6788 ( .A1(n5205), .A2(n5338), .ZN(n5339) );
  INV_X1 U6789 ( .A(n7344), .ZN(n8349) );
  NAND2_X1 U6790 ( .A1(n7033), .A2(n8015), .ZN(n5348) );
  NAND2_X1 U6791 ( .A1(n5349), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5346) );
  XNOR2_X1 U6792 ( .A(n5346), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6016) );
  AOI22_X1 U6793 ( .A1(n5469), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5468), .B2(
        n6016), .ZN(n5347) );
  NAND2_X2 U6794 ( .A1(n5348), .A2(n5347), .ZN(n5739) );
  NAND2_X1 U6795 ( .A1(n8349), .A2(n5739), .ZN(n5380) );
  AND2_X1 U6796 ( .A1(n7369), .A2(n5380), .ZN(n7339) );
  XNOR2_X1 U6797 ( .A(n5360), .B(n5359), .ZN(n7161) );
  NAND2_X1 U6798 ( .A1(n7161), .A2(n8015), .ZN(n5352) );
  OR2_X1 U6799 ( .A1(n5367), .A2(n5657), .ZN(n5350) );
  XNOR2_X1 U6800 ( .A(n5350), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6018) );
  AOI22_X1 U6801 ( .A1(n5469), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5468), .B2(
        n6018), .ZN(n5351) );
  NAND2_X1 U6802 ( .A1(n5323), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U6803 ( .A1(n5353), .A2(n9305), .ZN(n5354) );
  NAND2_X1 U6804 ( .A1(n5371), .A2(n5354), .ZN(n7347) );
  OR2_X1 U6805 ( .A1(n5203), .A2(n7347), .ZN(n5357) );
  NAND2_X1 U6806 ( .A1(n5204), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6807 ( .A1(n5206), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5355) );
  NAND4_X1 U6808 ( .A1(n5358), .A2(n5357), .A3(n5356), .A4(n5355), .ZN(n8348)
         );
  INV_X1 U6809 ( .A(n8348), .ZN(n7231) );
  NAND2_X1 U6810 ( .A1(n10154), .A2(n7231), .ZN(n5382) );
  AND2_X1 U6811 ( .A1(n10154), .A2(n8348), .ZN(n8085) );
  INV_X1 U6812 ( .A(n8085), .ZN(n8088) );
  NAND2_X1 U6813 ( .A1(n7350), .A2(n7231), .ZN(n8089) );
  NAND2_X1 U6814 ( .A1(n5362), .A2(n5361), .ZN(n5365) );
  INV_X1 U6815 ( .A(n5363), .ZN(n5364) );
  NAND2_X1 U6816 ( .A1(n7278), .A2(n8015), .ZN(n5369) );
  NAND2_X1 U6817 ( .A1(n5367), .A2(n5366), .ZN(n5438) );
  NAND2_X1 U6818 ( .A1(n5438), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5387) );
  XNOR2_X1 U6819 ( .A(n5387), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7098) );
  AOI22_X1 U6820 ( .A1(n5469), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5468), .B2(
        n7098), .ZN(n5368) );
  NAND2_X1 U6821 ( .A1(n5204), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5377) );
  INV_X1 U6822 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6021) );
  OR2_X1 U6823 ( .A1(n6186), .A2(n6021), .ZN(n5376) );
  INV_X1 U6824 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6825 ( .A1(n5371), .A2(n5370), .ZN(n5372) );
  NAND2_X1 U6826 ( .A1(n5395), .A2(n5372), .ZN(n7471) );
  OR2_X1 U6827 ( .A1(n5203), .A2(n7471), .ZN(n5375) );
  INV_X1 U6828 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5373) );
  OR2_X1 U6829 ( .A1(n4380), .A2(n5373), .ZN(n5374) );
  OR2_X1 U6830 ( .A1(n8728), .A2(n7440), .ZN(n8096) );
  NAND2_X1 U6831 ( .A1(n8728), .A2(n7440), .ZN(n8095) );
  INV_X1 U6832 ( .A(n7440), .ZN(n8347) );
  AND2_X1 U6833 ( .A1(n8728), .A2(n8347), .ZN(n5378) );
  INV_X1 U6834 ( .A(n7434), .ZN(n5379) );
  AND2_X1 U6835 ( .A1(n7339), .A2(n5379), .ZN(n5383) );
  INV_X1 U6836 ( .A(n5380), .ZN(n5381) );
  OR2_X1 U6837 ( .A1(n7344), .A2(n5739), .ZN(n8087) );
  NAND2_X1 U6838 ( .A1(n5739), .A2(n7344), .ZN(n8084) );
  AND2_X1 U6839 ( .A1(n8087), .A2(n8084), .ZN(n8195) );
  INV_X1 U6840 ( .A(n8195), .ZN(n7380) );
  OR2_X1 U6841 ( .A1(n5381), .A2(n7380), .ZN(n7340) );
  AND2_X1 U6842 ( .A1(n7340), .A2(n5382), .ZN(n7460) );
  XNOR2_X1 U6843 ( .A(n5385), .B(n5384), .ZN(n7311) );
  NAND2_X1 U6844 ( .A1(n7311), .A2(n8015), .ZN(n5393) );
  NAND2_X1 U6845 ( .A1(n5387), .A2(n5386), .ZN(n5388) );
  NAND2_X1 U6846 ( .A1(n5388), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5390) );
  INV_X1 U6847 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U6848 ( .A1(n5390), .A2(n5389), .ZN(n5404) );
  OR2_X1 U6849 ( .A1(n5390), .A2(n5389), .ZN(n5391) );
  AND2_X1 U6850 ( .A1(n5404), .A2(n5391), .ZN(n8365) );
  AOI22_X1 U6851 ( .A1(n5469), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5468), .B2(
        n8365), .ZN(n5392) );
  NAND2_X1 U6852 ( .A1(n5204), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5401) );
  INV_X1 U6853 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5992) );
  OR2_X1 U6854 ( .A1(n6186), .A2(n5992), .ZN(n5400) );
  NAND2_X1 U6855 ( .A1(n5395), .A2(n5394), .ZN(n5396) );
  NAND2_X1 U6856 ( .A1(n5424), .A2(n5396), .ZN(n7364) );
  OR2_X1 U6857 ( .A1(n5203), .A2(n7364), .ZN(n5399) );
  INV_X1 U6858 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5397) );
  OR2_X1 U6859 ( .A1(n4379), .A2(n5397), .ZN(n5398) );
  XNOR2_X1 U6860 ( .A(n8723), .B(n8103), .ZN(n8200) );
  NAND2_X1 U6861 ( .A1(n7412), .A2(n8015), .ZN(n5408) );
  NAND2_X1 U6862 ( .A1(n5404), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5406) );
  INV_X1 U6863 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5405) );
  XNOR2_X1 U6864 ( .A(n5406), .B(n5405), .ZN(n7515) );
  INV_X1 U6865 ( .A(n7515), .ZN(n5979) );
  AOI22_X1 U6866 ( .A1(n5469), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5468), .B2(
        n5979), .ZN(n5407) );
  NAND2_X1 U6867 ( .A1(n5204), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5412) );
  INV_X1 U6868 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7506) );
  OR2_X1 U6869 ( .A1(n6186), .A2(n7506), .ZN(n5411) );
  INV_X1 U6870 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5423) );
  XNOR2_X1 U6871 ( .A(n5424), .B(n5423), .ZN(n7528) );
  OR2_X1 U6872 ( .A1(n5203), .A2(n7528), .ZN(n5410) );
  INV_X1 U6873 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7453) );
  OR2_X1 U6874 ( .A1(n4380), .A2(n7453), .ZN(n5409) );
  NOR2_X1 U6875 ( .A1(n8718), .A2(n8625), .ZN(n8109) );
  NAND2_X1 U6876 ( .A1(n8718), .A2(n8625), .ZN(n8108) );
  NAND2_X1 U6877 ( .A1(n4797), .A2(n8108), .ZN(n8201) );
  INV_X1 U6878 ( .A(n8625), .ZN(n8345) );
  OR2_X1 U6879 ( .A1(n8718), .A2(n8345), .ZN(n5413) );
  INV_X1 U6880 ( .A(n8626), .ZN(n5431) );
  XNOR2_X1 U6881 ( .A(n5415), .B(n5414), .ZN(n7483) );
  NAND2_X1 U6882 ( .A1(n7483), .A2(n8015), .ZN(n5421) );
  INV_X1 U6883 ( .A(n5438), .ZN(n5418) );
  INV_X1 U6884 ( .A(n5416), .ZN(n5417) );
  NOR2_X1 U6885 ( .A1(n5417), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U6886 ( .A1(n4473), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5419) );
  XNOR2_X1 U6887 ( .A(n5419), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8376) );
  AOI22_X1 U6888 ( .A1(n5469), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5468), .B2(
        n8376), .ZN(n5420) );
  NAND2_X1 U6889 ( .A1(n5204), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5429) );
  INV_X1 U6890 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n5991) );
  OR2_X1 U6891 ( .A1(n6186), .A2(n5991), .ZN(n5428) );
  INV_X1 U6892 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5422) );
  OAI21_X1 U6893 ( .B1(n5424), .B2(n5423), .A(n5422), .ZN(n5425) );
  NAND2_X1 U6894 ( .A1(n5425), .A2(n5442), .ZN(n7543) );
  OR2_X1 U6895 ( .A1(n5203), .A2(n7543), .ZN(n5427) );
  INV_X1 U6896 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5967) );
  OR2_X1 U6897 ( .A1(n4379), .A2(n5967), .ZN(n5426) );
  OR2_X1 U6898 ( .A1(n8712), .A2(n8613), .ZN(n8113) );
  INV_X1 U6899 ( .A(n8613), .ZN(n8344) );
  NAND2_X1 U6900 ( .A1(n8712), .A2(n8344), .ZN(n5432) );
  XNOR2_X1 U6901 ( .A(n5434), .B(n5433), .ZN(n7567) );
  NAND2_X1 U6902 ( .A1(n7567), .A2(n8015), .ZN(n5441) );
  INV_X1 U6903 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U6904 ( .A1(n5436), .A2(n5435), .ZN(n5437) );
  NAND2_X1 U6905 ( .A1(n4472), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5439) );
  XNOR2_X1 U6906 ( .A(n5439), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8393) );
  AOI22_X1 U6907 ( .A1(n5469), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5468), .B2(
        n8393), .ZN(n5440) );
  NAND2_X1 U6908 ( .A1(n5323), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5447) );
  INV_X1 U6909 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9461) );
  OR2_X1 U6910 ( .A1(n5194), .A2(n9461), .ZN(n5446) );
  NAND2_X1 U6911 ( .A1(n5442), .A2(n7518), .ZN(n5443) );
  NAND2_X1 U6912 ( .A1(n5455), .A2(n5443), .ZN(n8605) );
  OR2_X1 U6913 ( .A1(n5203), .A2(n8605), .ZN(n5445) );
  INV_X1 U6914 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8606) );
  OR2_X1 U6915 ( .A1(n4380), .A2(n8606), .ZN(n5444) );
  NAND2_X1 U6916 ( .A1(n8709), .A2(n8623), .ZN(n8120) );
  INV_X1 U6917 ( .A(n8623), .ZN(n8595) );
  OR2_X1 U6918 ( .A1(n8709), .A2(n8595), .ZN(n5449) );
  XNOR2_X1 U6919 ( .A(n5451), .B(n5450), .ZN(n7571) );
  NAND2_X1 U6920 ( .A1(n7571), .A2(n8015), .ZN(n5453) );
  XNOR2_X1 U6921 ( .A(n5464), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8406) );
  AOI22_X1 U6922 ( .A1(n5469), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5468), .B2(
        n8406), .ZN(n5452) );
  NAND2_X1 U6923 ( .A1(n5204), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5460) );
  INV_X1 U6924 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U6925 ( .A1(n5455), .A2(n5454), .ZN(n5456) );
  NAND2_X1 U6926 ( .A1(n5472), .A2(n5456), .ZN(n8589) );
  OR2_X1 U6927 ( .A1(n5203), .A2(n8589), .ZN(n5459) );
  NAND2_X1 U6928 ( .A1(n5206), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U6929 ( .A1(n5323), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5457) );
  NAND4_X1 U6930 ( .A1(n5460), .A2(n5459), .A3(n5458), .A4(n5457), .ZN(n8343)
         );
  INV_X1 U6931 ( .A(n8343), .ZN(n8614) );
  OR2_X1 U6932 ( .A1(n8592), .A2(n8614), .ZN(n5461) );
  XNOR2_X1 U6933 ( .A(n5463), .B(n5462), .ZN(n7581) );
  NAND2_X1 U6934 ( .A1(n7581), .A2(n8015), .ZN(n5471) );
  INV_X1 U6935 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U6936 ( .A1(n5467), .A2(n5466), .ZN(n5605) );
  AOI22_X1 U6937 ( .A1(n5469), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5468), .B2(
        n5638), .ZN(n5470) );
  INV_X1 U6938 ( .A(n8698), .ZN(n5478) );
  NAND2_X1 U6939 ( .A1(n5204), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5477) );
  INV_X1 U6940 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9421) );
  OR2_X1 U6941 ( .A1(n4380), .A2(n9421), .ZN(n5476) );
  NAND2_X1 U6942 ( .A1(n5472), .A2(n8271), .ZN(n5473) );
  NAND2_X1 U6943 ( .A1(n5485), .A2(n5473), .ZN(n8583) );
  OR2_X1 U6944 ( .A1(n5203), .A2(n8583), .ZN(n5475) );
  INV_X1 U6945 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9452) );
  OR2_X1 U6946 ( .A1(n6186), .A2(n9452), .ZN(n5474) );
  NAND2_X1 U6947 ( .A1(n5478), .A2(n8311), .ZN(n5479) );
  INV_X1 U6948 ( .A(n8311), .ZN(n8596) );
  XNOR2_X1 U6949 ( .A(n5481), .B(n5480), .ZN(n7593) );
  NAND2_X1 U6950 ( .A1(n7593), .A2(n8015), .ZN(n5483) );
  OR2_X1 U6951 ( .A1(n5569), .A2(n6720), .ZN(n5482) );
  NAND2_X1 U6952 ( .A1(n5204), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5491) );
  INV_X1 U6953 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5484) );
  OR2_X1 U6954 ( .A1(n4379), .A2(n5484), .ZN(n5490) );
  INV_X1 U6955 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8306) );
  NAND2_X1 U6956 ( .A1(n5485), .A2(n8306), .ZN(n5486) );
  NAND2_X1 U6957 ( .A1(n5496), .A2(n5486), .ZN(n8561) );
  OR2_X1 U6958 ( .A1(n5203), .A2(n8561), .ZN(n5489) );
  INV_X1 U6959 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n5487) );
  OR2_X1 U6960 ( .A1(n6186), .A2(n5487), .ZN(n5488) );
  NAND2_X1 U6961 ( .A1(n8692), .A2(n8553), .ZN(n8137) );
  INV_X1 U6962 ( .A(n8692), .ZN(n8564) );
  XNOR2_X1 U6963 ( .A(n5493), .B(n5492), .ZN(n7605) );
  NAND2_X1 U6964 ( .A1(n7605), .A2(n8015), .ZN(n5495) );
  INV_X1 U6965 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n9322) );
  OR2_X1 U6966 ( .A1(n5569), .A2(n9322), .ZN(n5494) );
  INV_X1 U6967 ( .A(n8687), .ZN(n8544) );
  NAND2_X1 U6968 ( .A1(n5204), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5501) );
  INV_X1 U6969 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9427) );
  OR2_X1 U6970 ( .A1(n6186), .A2(n9427), .ZN(n5500) );
  NAND2_X1 U6971 ( .A1(n5496), .A2(n9451), .ZN(n5497) );
  NAND2_X1 U6972 ( .A1(n5520), .A2(n5497), .ZN(n8545) );
  OR2_X1 U6973 ( .A1(n5203), .A2(n8545), .ZN(n5499) );
  INV_X1 U6974 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8546) );
  OR2_X1 U6975 ( .A1(n4380), .A2(n8546), .ZN(n5498) );
  XNOR2_X1 U6976 ( .A(n5503), .B(n5502), .ZN(n7619) );
  NAND2_X1 U6977 ( .A1(n7619), .A2(n8015), .ZN(n5505) );
  OR2_X1 U6978 ( .A1(n5569), .A2(n9358), .ZN(n5504) );
  NAND2_X1 U6979 ( .A1(n5204), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5511) );
  INV_X1 U6980 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n5506) );
  OR2_X1 U6981 ( .A1(n6186), .A2(n5506), .ZN(n5510) );
  INV_X1 U6982 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8324) );
  XNOR2_X1 U6983 ( .A(n5520), .B(n8324), .ZN(n8323) );
  OR2_X1 U6984 ( .A1(n5203), .A2(n8323), .ZN(n5509) );
  INV_X1 U6985 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5507) );
  OR2_X1 U6986 ( .A1(n4379), .A2(n5507), .ZN(n5508) );
  NAND2_X1 U6987 ( .A1(n8681), .A2(n8554), .ZN(n8143) );
  INV_X1 U6988 ( .A(n8681), .ZN(n8534) );
  OR2_X1 U6989 ( .A1(n5515), .A2(n5514), .ZN(n5516) );
  NAND2_X1 U6990 ( .A1(n5517), .A2(n5516), .ZN(n7629) );
  NAND2_X1 U6991 ( .A1(n7629), .A2(n8015), .ZN(n5519) );
  OR2_X1 U6992 ( .A1(n5569), .A2(n7079), .ZN(n5518) );
  NAND2_X1 U6993 ( .A1(n5204), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5526) );
  INV_X1 U6994 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9304) );
  OAI21_X1 U6995 ( .B1(n5520), .B2(n8324), .A(n9304), .ZN(n5521) );
  AND2_X1 U6996 ( .A1(n5522), .A2(n5521), .ZN(n8520) );
  NAND2_X1 U6997 ( .A1(n5599), .A2(n8520), .ZN(n5525) );
  NAND2_X1 U6998 ( .A1(n5206), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U6999 ( .A1(n5323), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5523) );
  NAND4_X1 U7000 ( .A1(n5526), .A2(n5525), .A3(n5524), .A4(n5523), .ZN(n8507)
         );
  NAND2_X1 U7001 ( .A1(n8522), .A2(n8507), .ZN(n8148) );
  INV_X1 U7002 ( .A(n8507), .ZN(n8299) );
  NAND2_X1 U7003 ( .A1(n8674), .A2(n8299), .ZN(n5634) );
  NAND2_X1 U7004 ( .A1(n8674), .A2(n8507), .ZN(n5527) );
  NAND2_X1 U7005 ( .A1(n8676), .A2(n5527), .ZN(n8498) );
  NAND2_X1 U7006 ( .A1(n5529), .A2(SI_24_), .ZN(n5530) );
  INV_X1 U7007 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7334) );
  INV_X1 U7008 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9376) );
  MUX2_X1 U7009 ( .A(n7334), .B(n9376), .S(n7743), .Z(n5533) );
  INV_X1 U7010 ( .A(SI_25_), .ZN(n5532) );
  NAND2_X1 U7011 ( .A1(n5533), .A2(n5532), .ZN(n5543) );
  INV_X1 U7012 ( .A(n5533), .ZN(n5534) );
  NAND2_X1 U7013 ( .A1(n5534), .A2(SI_25_), .ZN(n5535) );
  NAND2_X1 U7014 ( .A1(n5543), .A2(n5535), .ZN(n5544) );
  NAND2_X1 U7015 ( .A1(n7651), .A2(n8015), .ZN(n5537) );
  OR2_X1 U7016 ( .A1(n5569), .A2(n7334), .ZN(n5536) );
  XNOR2_X1 U7017 ( .A(n5552), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n8482) );
  NAND2_X1 U7018 ( .A1(n8482), .A2(n5599), .ZN(n5542) );
  INV_X1 U7019 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8484) );
  NAND2_X1 U7020 ( .A1(n5323), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U7021 ( .A1(n5204), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5538) );
  OAI211_X1 U7022 ( .C1(n8484), .C2(n4380), .A(n5539), .B(n5538), .ZN(n5540)
         );
  INV_X1 U7023 ( .A(n5540), .ZN(n5541) );
  NAND2_X1 U7024 ( .A1(n8666), .A2(n8330), .ZN(n8157) );
  INV_X1 U7025 ( .A(n8330), .ZN(n8508) );
  INV_X1 U7026 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7386) );
  INV_X1 U7027 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7337) );
  MUX2_X1 U7028 ( .A(n7386), .B(n7337), .S(n7743), .Z(n5547) );
  INV_X1 U7029 ( .A(SI_26_), .ZN(n5546) );
  NAND2_X1 U7030 ( .A1(n5547), .A2(n5546), .ZN(n5560) );
  INV_X1 U7031 ( .A(n5547), .ZN(n5548) );
  NAND2_X1 U7032 ( .A1(n5548), .A2(SI_26_), .ZN(n5549) );
  AND2_X1 U7033 ( .A1(n5560), .A2(n5549), .ZN(n5558) );
  NAND2_X1 U7034 ( .A1(n7663), .A2(n8015), .ZN(n5551) );
  OR2_X1 U7035 ( .A1(n5569), .A2(n7386), .ZN(n5550) );
  INV_X1 U7036 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n5556) );
  INV_X1 U7037 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8287) );
  INV_X1 U7038 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8333) );
  OAI21_X1 U7039 ( .B1(n5552), .B2(n8287), .A(n8333), .ZN(n5553) );
  AND2_X1 U7040 ( .A1(n5553), .A2(n5573), .ZN(n8475) );
  NAND2_X1 U7041 ( .A1(n8475), .A2(n5599), .ZN(n5555) );
  AOI22_X1 U7042 ( .A1(n5323), .A2(P2_REG1_REG_26__SCAN_IN), .B1(n5204), .B2(
        P2_REG0_REG_26__SCAN_IN), .ZN(n5554) );
  OAI211_X1 U7043 ( .C1(n4379), .C2(n5556), .A(n5555), .B(n5554), .ZN(n8458)
         );
  INV_X1 U7044 ( .A(n8458), .ZN(n8254) );
  INV_X1 U7045 ( .A(n8467), .ZN(n5557) );
  INV_X1 U7046 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9222) );
  INV_X1 U7047 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5561) );
  MUX2_X1 U7048 ( .A(n9222), .B(n5561), .S(n7743), .Z(n5563) );
  INV_X1 U7049 ( .A(SI_27_), .ZN(n5562) );
  NAND2_X1 U7050 ( .A1(n5563), .A2(n5562), .ZN(n5578) );
  INV_X1 U7051 ( .A(n5563), .ZN(n5564) );
  NAND2_X1 U7052 ( .A1(n5564), .A2(SI_27_), .ZN(n5565) );
  AND2_X1 U7053 ( .A1(n5578), .A2(n5565), .ZN(n5566) );
  OR2_X1 U7054 ( .A1(n5569), .A2(n9222), .ZN(n5570) );
  INV_X1 U7055 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5577) );
  INV_X1 U7056 ( .A(n5573), .ZN(n5572) );
  NAND2_X1 U7057 ( .A1(n5572), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5583) );
  INV_X1 U7058 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U7059 ( .A1(n5573), .A2(n9386), .ZN(n5574) );
  NAND2_X1 U7060 ( .A1(n5583), .A2(n5574), .ZN(n8451) );
  OR2_X1 U7061 ( .A1(n8451), .A2(n5203), .ZN(n5576) );
  AOI22_X1 U7062 ( .A1(n5323), .A2(P2_REG1_REG_27__SCAN_IN), .B1(n5204), .B2(
        P2_REG0_REG_27__SCAN_IN), .ZN(n5575) );
  OAI211_X1 U7063 ( .C1(n4379), .C2(n5577), .A(n5576), .B(n5575), .ZN(n8341)
         );
  INV_X1 U7064 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8011) );
  INV_X1 U7065 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5580) );
  MUX2_X1 U7066 ( .A(n8011), .B(n5580), .S(n7743), .Z(n5592) );
  XNOR2_X1 U7067 ( .A(n5592), .B(SI_28_), .ZN(n7554) );
  OR2_X1 U7068 ( .A1(n5569), .A2(n8011), .ZN(n5581) );
  INV_X1 U7069 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5837) );
  OR2_X1 U7070 ( .A1(n5583), .A2(n5837), .ZN(n5598) );
  NAND2_X1 U7071 ( .A1(n5583), .A2(n5837), .ZN(n5584) );
  NAND2_X1 U7072 ( .A1(n8435), .A2(n5599), .ZN(n5590) );
  INV_X1 U7073 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7074 ( .A1(n5206), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U7075 ( .A1(n5204), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5585) );
  OAI211_X1 U7076 ( .C1(n6186), .C2(n5587), .A(n5586), .B(n5585), .ZN(n5588)
         );
  INV_X1 U7077 ( .A(n5588), .ZN(n5589) );
  NAND2_X1 U7078 ( .A1(n5590), .A2(n5589), .ZN(n8459) );
  INV_X1 U7079 ( .A(n8459), .ZN(n8255) );
  NAND2_X1 U7080 ( .A1(n7562), .A2(n7554), .ZN(n5593) );
  INV_X1 U7081 ( .A(SI_28_), .ZN(n5591) );
  NAND2_X1 U7082 ( .A1(n5592), .A2(n5591), .ZN(n7558) );
  INV_X1 U7083 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8762) );
  INV_X1 U7084 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9697) );
  MUX2_X1 U7085 ( .A(n8762), .B(n9697), .S(n7743), .Z(n7553) );
  XNOR2_X1 U7086 ( .A(n7553), .B(SI_29_), .ZN(n5594) );
  NAND2_X1 U7087 ( .A1(n8760), .A2(n8015), .ZN(n5597) );
  OR2_X1 U7088 ( .A1(n5569), .A2(n8762), .ZN(n5596) );
  INV_X1 U7089 ( .A(n5598), .ZN(n8241) );
  NAND2_X1 U7090 ( .A1(n8241), .A2(n5599), .ZN(n5602) );
  AOI22_X1 U7091 ( .A1(n5323), .A2(P2_REG1_REG_29__SCAN_IN), .B1(n5204), .B2(
        P2_REG0_REG_29__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U7092 ( .A1(n5206), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5600) );
  INV_X1 U7093 ( .A(n8211), .ZN(n5603) );
  XNOR2_X1 U7094 ( .A(n5604), .B(n5603), .ZN(n8247) );
  XNOR2_X2 U7095 ( .A(n5606), .B(P2_IR_REG_20__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U7096 ( .A1(n5607), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5609) );
  INV_X1 U7097 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5608) );
  XNOR2_X1 U7098 ( .A(n5609), .B(n5608), .ZN(n8024) );
  OR2_X1 U7099 ( .A1(n5610), .A2(n5657), .ZN(n5611) );
  XNOR2_X1 U7100 ( .A(n5611), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8228) );
  INV_X1 U7101 ( .A(n8228), .ZN(n7018) );
  NAND2_X1 U7102 ( .A1(n6402), .A2(n7018), .ZN(n5613) );
  INV_X1 U7103 ( .A(n8024), .ZN(n8216) );
  AND2_X1 U7104 ( .A1(n8228), .A2(n8216), .ZN(n5982) );
  NOR2_X1 U7105 ( .A1(n5638), .A2(n5982), .ZN(n5612) );
  NAND2_X1 U7106 ( .A1(n5613), .A2(n5612), .ZN(n8630) );
  OR2_X1 U7107 ( .A1(n8025), .A2(n5650), .ZN(n10142) );
  NAND2_X1 U7108 ( .A1(n5614), .A2(n10096), .ZN(n10062) );
  NAND2_X1 U7109 ( .A1(n10062), .A2(n8043), .ZN(n8036) );
  NAND2_X1 U7110 ( .A1(n8036), .A2(n5615), .ZN(n6456) );
  INV_X1 U7111 ( .A(n6456), .ZN(n5617) );
  INV_X1 U7112 ( .A(n8187), .ZN(n5616) );
  NAND2_X1 U7113 ( .A1(n5617), .A2(n5616), .ZN(n6454) );
  NAND2_X1 U7114 ( .A1(n6454), .A2(n8044), .ZN(n5618) );
  NAND2_X1 U7115 ( .A1(n8184), .A2(n5618), .ZN(n6600) );
  INV_X1 U7116 ( .A(n6599), .ZN(n8031) );
  NOR2_X1 U7117 ( .A1(n6601), .A2(n8031), .ZN(n5619) );
  NAND2_X1 U7118 ( .A1(n6600), .A2(n5619), .ZN(n5620) );
  NAND2_X1 U7119 ( .A1(n6760), .A2(n8033), .ZN(n5622) );
  NAND2_X1 U7120 ( .A1(n5622), .A2(n8185), .ZN(n6758) );
  INV_X1 U7121 ( .A(n8059), .ZN(n8034) );
  NOR2_X1 U7122 ( .A1(n8060), .A2(n8034), .ZN(n5623) );
  NAND2_X1 U7123 ( .A1(n6758), .A2(n5623), .ZN(n6839) );
  INV_X1 U7124 ( .A(n5624), .ZN(n7082) );
  NOR2_X1 U7125 ( .A1(n8192), .A2(n7082), .ZN(n8065) );
  AND2_X1 U7126 ( .A1(n7151), .A2(n8077), .ZN(n7376) );
  INV_X1 U7127 ( .A(n7376), .ZN(n5626) );
  OR2_X1 U7128 ( .A1(n8723), .A2(n8103), .ZN(n5628) );
  AND2_X1 U7129 ( .A1(n8197), .A2(n5628), .ZN(n5632) );
  INV_X1 U7130 ( .A(n5628), .ZN(n5631) );
  INV_X1 U7131 ( .A(n8200), .ZN(n5629) );
  AND2_X1 U7132 ( .A1(n5629), .A2(n8095), .ZN(n5630) );
  NAND2_X1 U7133 ( .A1(n8702), .A2(n8614), .ZN(n8180) );
  AND2_X1 U7134 ( .A1(n8592), .A2(n8343), .ZN(n8118) );
  AOI21_X1 U7135 ( .B1(n8593), .B2(n8180), .A(n8118), .ZN(n8577) );
  OR2_X1 U7136 ( .A1(n8698), .A2(n8311), .ZN(n8133) );
  NAND2_X1 U7137 ( .A1(n8698), .A2(n8311), .ZN(n8125) );
  INV_X1 U7138 ( .A(n8125), .ZN(n5633) );
  AOI21_X2 U7139 ( .B1(n8577), .B2(n8576), .A(n5633), .ZN(n8567) );
  NAND2_X1 U7140 ( .A1(n8567), .A2(n8566), .ZN(n8565) );
  OR2_X1 U7141 ( .A1(n8687), .A2(n8308), .ZN(n8138) );
  NAND2_X1 U7142 ( .A1(n8687), .A2(n8308), .ZN(n8142) );
  NAND2_X1 U7143 ( .A1(n8138), .A2(n8142), .ZN(n8551) );
  NAND2_X1 U7144 ( .A1(n8535), .A2(n8131), .ZN(n8515) );
  INV_X1 U7145 ( .A(n5634), .ZN(n8147) );
  INV_X1 U7146 ( .A(n5635), .ZN(n8150) );
  INV_X1 U7147 ( .A(n8341), .ZN(n8441) );
  NAND2_X1 U7148 ( .A1(n8438), .A2(n8430), .ZN(n8444) );
  XNOR2_X1 U7149 ( .A(n8012), .B(n8211), .ZN(n5646) );
  NAND2_X1 U7150 ( .A1(n5650), .A2(n8216), .ZN(n8022) );
  INV_X1 U7151 ( .A(n8179), .ZN(n8178) );
  NAND2_X1 U7152 ( .A1(n8022), .A2(n8178), .ZN(n10061) );
  INV_X1 U7153 ( .A(n5639), .ZN(n5640) );
  INV_X1 U7154 ( .A(n7533), .ZN(n8225) );
  NAND2_X1 U7155 ( .A1(n5639), .A2(n5982), .ZN(n8622) );
  AOI21_X1 U7156 ( .B1(n8225), .B2(P2_B_REG_SCAN_IN), .A(n8622), .ZN(n8419) );
  INV_X1 U7157 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n5643) );
  NAND2_X1 U7158 ( .A1(n5206), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U7159 ( .A1(n5204), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5641) );
  OAI211_X1 U7160 ( .C1(n6186), .C2(n5643), .A(n5642), .B(n5641), .ZN(n8340)
         );
  NAND2_X1 U7161 ( .A1(n5647), .A2(n10105), .ZN(n6460) );
  NOR2_X1 U7162 ( .A1(n6584), .A2(n10116), .ZN(n5648) );
  NOR2_X2 U7163 ( .A1(n7345), .A2(n7350), .ZN(n7346) );
  INV_X1 U7164 ( .A(n8728), .ZN(n7474) );
  INV_X1 U7165 ( .A(n8712), .ZN(n8640) );
  INV_X1 U7166 ( .A(n8709), .ZN(n5649) );
  OR2_X2 U7167 ( .A1(n8531), .A2(n8681), .ZN(n8529) );
  OR2_X2 U7168 ( .A1(n8529), .A2(n8674), .ZN(n8518) );
  AOI21_X1 U7169 ( .B1(n8240), .B2(n8432), .A(n8424), .ZN(n8246) );
  INV_X1 U7170 ( .A(n10155), .ZN(n10138) );
  AND2_X2 U7171 ( .A1(n8224), .A2(n10097), .ZN(n10137) );
  AOI22_X1 U7172 ( .A1(n8246), .A2(n10138), .B1(n10137), .B2(n8240), .ZN(n5651) );
  NAND2_X1 U7173 ( .A1(n8224), .A2(n5982), .ZN(n5834) );
  NOR2_X1 U7174 ( .A1(n5652), .A2(n5657), .ZN(n5653) );
  MUX2_X1 U7175 ( .A(n5657), .B(n5653), .S(P2_IR_REG_25__SCAN_IN), .Z(n5654)
         );
  INV_X1 U7176 ( .A(n5654), .ZN(n5656) );
  NAND2_X1 U7177 ( .A1(n5656), .A2(n5655), .ZN(n7333) );
  OR2_X1 U7178 ( .A1(n5658), .A2(n5657), .ZN(n5667) );
  INV_X1 U7179 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5659) );
  NAND2_X1 U7180 ( .A1(n5667), .A2(n5659), .ZN(n5660) );
  NAND2_X1 U7181 ( .A1(n5660), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5662) );
  INV_X1 U7182 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5661) );
  XNOR2_X1 U7183 ( .A(n5662), .B(n5661), .ZN(n7127) );
  NOR2_X1 U7184 ( .A1(n7333), .A2(n7127), .ZN(n5666) );
  NAND2_X1 U7185 ( .A1(n5655), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5663) );
  MUX2_X1 U7186 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5663), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5665) );
  NAND2_X1 U7187 ( .A1(n5665), .A2(n5664), .ZN(n7388) );
  INV_X1 U7188 ( .A(n7388), .ZN(n5679) );
  NAND2_X1 U7189 ( .A1(n5666), .A2(n5679), .ZN(n5863) );
  XNOR2_X1 U7190 ( .A(n5667), .B(P2_IR_REG_23__SCAN_IN), .ZN(n5983) );
  NOR2_X1 U7191 ( .A1(n5983), .A2(P2_U3152), .ZN(n10094) );
  NOR4_X1 U7192 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5676) );
  INV_X1 U7193 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10083) );
  INV_X1 U7194 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n10084) );
  INV_X1 U7195 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10082) );
  INV_X1 U7196 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10085) );
  NAND4_X1 U7197 ( .A1(n10083), .A2(n10084), .A3(n10082), .A4(n10085), .ZN(
        n5673) );
  NOR4_X1 U7198 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5671) );
  NOR4_X1 U7199 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n5670) );
  NOR4_X1 U7200 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5669) );
  NOR4_X1 U7201 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5668) );
  NAND4_X1 U7202 ( .A1(n5671), .A2(n5670), .A3(n5669), .A4(n5668), .ZN(n5672)
         );
  NOR4_X1 U7203 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n5673), .A4(n5672), .ZN(n5675) );
  NOR4_X1 U7204 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n5674) );
  NAND3_X1 U7205 ( .A1(n5676), .A2(n5675), .A3(n5674), .ZN(n5680) );
  XNOR2_X1 U7206 ( .A(n7127), .B(P2_B_REG_SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7207 ( .A1(n7333), .A2(n5677), .ZN(n5678) );
  NAND2_X1 U7208 ( .A1(n5680), .A2(n5682), .ZN(n5822) );
  NAND3_X1 U7209 ( .A1(n5834), .A2(n10081), .A3(n5822), .ZN(n6396) );
  INV_X1 U7210 ( .A(n5682), .ZN(n10080) );
  NAND2_X1 U7211 ( .A1(n7388), .A2(n7333), .ZN(n10091) );
  OAI21_X1 U7212 ( .B1(P2_D_REG_1__SCAN_IN), .B2(n10080), .A(n10091), .ZN(
        n6398) );
  NAND2_X1 U7213 ( .A1(n6398), .A2(n5831), .ZN(n5681) );
  NOR2_X1 U7214 ( .A1(n6396), .A2(n5681), .ZN(n5687) );
  INV_X1 U7215 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10089) );
  AND2_X1 U7216 ( .A1(n7388), .A2(n7127), .ZN(n10090) );
  AOI21_X1 U7217 ( .B1(n5682), .B2(n10089), .A(n10090), .ZN(n6397) );
  INV_X1 U7218 ( .A(n6397), .ZN(n5683) );
  AND2_X2 U7219 ( .A1(n5687), .A2(n5683), .ZN(n10163) );
  NAND2_X1 U7220 ( .A1(n5688), .A2(n10163), .ZN(n5686) );
  OR2_X1 U7221 ( .A1(n10163), .A2(n5684), .ZN(n5685) );
  NAND2_X1 U7222 ( .A1(n5686), .A2(n5685), .ZN(P2_U3517) );
  AND2_X2 U7223 ( .A1(n5687), .A2(n6397), .ZN(n10177) );
  NAND2_X1 U7224 ( .A1(n5690), .A2(n8024), .ZN(n5689) );
  XNOR2_X1 U7225 ( .A(n4747), .B(n5816), .ZN(n8283) );
  OR2_X4 U7226 ( .A1(n8224), .A2(n5690), .ZN(n8023) );
  NAND2_X1 U7227 ( .A1(n8507), .A2(n8023), .ZN(n8294) );
  INV_X1 U7228 ( .A(n6294), .ZN(n5694) );
  XNOR2_X1 U7229 ( .A(n6296), .B(n4378), .ZN(n5692) );
  NAND2_X1 U7230 ( .A1(n5691), .A2(n5692), .ZN(n5695) );
  OAI21_X1 U7231 ( .B1(n5692), .B2(n5691), .A(n5695), .ZN(n6291) );
  INV_X1 U7232 ( .A(n6291), .ZN(n5693) );
  NAND2_X1 U7233 ( .A1(n5694), .A2(n5693), .ZN(n6292) );
  NAND2_X1 U7234 ( .A1(n6292), .A2(n5695), .ZN(n6303) );
  NAND2_X1 U7235 ( .A1(n10064), .A2(n8023), .ZN(n5696) );
  XNOR2_X1 U7236 ( .A(n5697), .B(n5696), .ZN(n6302) );
  NAND2_X1 U7237 ( .A1(n8357), .A2(n8023), .ZN(n5698) );
  XNOR2_X1 U7238 ( .A(n6433), .B(n4504), .ZN(n5699) );
  XNOR2_X1 U7239 ( .A(n5698), .B(n5699), .ZN(n6390) );
  NAND2_X1 U7240 ( .A1(n6391), .A2(n6390), .ZN(n5702) );
  INV_X1 U7241 ( .A(n5698), .ZN(n5700) );
  NAND2_X1 U7242 ( .A1(n5700), .A2(n5699), .ZN(n5701) );
  NAND2_X1 U7243 ( .A1(n8356), .A2(n8023), .ZN(n5703) );
  XNOR2_X1 U7244 ( .A(n10116), .B(n4378), .ZN(n5704) );
  NAND2_X1 U7245 ( .A1(n5703), .A2(n5704), .ZN(n5709) );
  INV_X1 U7246 ( .A(n5703), .ZN(n5706) );
  INV_X1 U7247 ( .A(n5704), .ZN(n5705) );
  NAND2_X1 U7248 ( .A1(n5706), .A2(n5705), .ZN(n5707) );
  NAND2_X1 U7249 ( .A1(n5709), .A2(n5707), .ZN(n6414) );
  INV_X1 U7250 ( .A(n6414), .ZN(n5708) );
  INV_X1 U7251 ( .A(n6549), .ZN(n5715) );
  NAND2_X1 U7252 ( .A1(n8355), .A2(n8023), .ZN(n5710) );
  XNOR2_X1 U7253 ( .A(n6584), .B(n5819), .ZN(n5711) );
  XNOR2_X1 U7254 ( .A(n5710), .B(n5711), .ZN(n6548) );
  INV_X1 U7255 ( .A(n6548), .ZN(n5714) );
  INV_X1 U7256 ( .A(n5710), .ZN(n5713) );
  INV_X1 U7257 ( .A(n5711), .ZN(n5712) );
  AOI21_X1 U7258 ( .B1(n5715), .B2(n5714), .A(n5015), .ZN(n6712) );
  NAND2_X1 U7259 ( .A1(n8354), .A2(n8023), .ZN(n5716) );
  XNOR2_X1 U7260 ( .A(n10128), .B(n5819), .ZN(n5717) );
  NAND2_X1 U7261 ( .A1(n5716), .A2(n5717), .ZN(n5721) );
  INV_X1 U7262 ( .A(n5716), .ZN(n5719) );
  INV_X1 U7263 ( .A(n5717), .ZN(n5718) );
  NAND2_X1 U7264 ( .A1(n5719), .A2(n5718), .ZN(n5720) );
  AND2_X1 U7265 ( .A1(n5721), .A2(n5720), .ZN(n6713) );
  NAND2_X1 U7266 ( .A1(n8353), .A2(n8023), .ZN(n5723) );
  XNOR2_X1 U7267 ( .A(n7008), .B(n5819), .ZN(n5724) );
  XNOR2_X1 U7268 ( .A(n5723), .B(n5724), .ZN(n6772) );
  INV_X1 U7269 ( .A(n6772), .ZN(n5722) );
  INV_X1 U7270 ( .A(n5723), .ZN(n5726) );
  INV_X1 U7271 ( .A(n5724), .ZN(n5725) );
  NAND2_X1 U7272 ( .A1(n5726), .A2(n5725), .ZN(n5727) );
  NAND2_X1 U7273 ( .A1(n8352), .A2(n8023), .ZN(n5729) );
  XNOR2_X1 U7274 ( .A(n10136), .B(n5816), .ZN(n5730) );
  XNOR2_X1 U7275 ( .A(n5729), .B(n5730), .ZN(n7020) );
  INV_X1 U7276 ( .A(n5729), .ZN(n5731) );
  AND2_X1 U7277 ( .A1(n5731), .A2(n5730), .ZN(n5732) );
  NAND2_X1 U7278 ( .A1(n8351), .A2(n8023), .ZN(n5733) );
  XNOR2_X1 U7279 ( .A(n7155), .B(n5819), .ZN(n5734) );
  NAND2_X1 U7280 ( .A1(n5733), .A2(n5734), .ZN(n5738) );
  INV_X1 U7281 ( .A(n5733), .ZN(n5736) );
  INV_X1 U7282 ( .A(n5734), .ZN(n5735) );
  NAND2_X1 U7283 ( .A1(n5736), .A2(n5735), .ZN(n5737) );
  AND2_X1 U7284 ( .A1(n5738), .A2(n5737), .ZN(n7113) );
  NAND2_X1 U7285 ( .A1(n8350), .A2(n8023), .ZN(n5748) );
  XNOR2_X1 U7286 ( .A(n7251), .B(n5819), .ZN(n5749) );
  XNOR2_X1 U7287 ( .A(n5748), .B(n5749), .ZN(n7226) );
  XNOR2_X1 U7288 ( .A(n5739), .B(n4504), .ZN(n5742) );
  NAND2_X1 U7289 ( .A1(n8349), .A2(n8023), .ZN(n5741) );
  INV_X1 U7290 ( .A(n5741), .ZN(n5740) );
  NAND2_X1 U7291 ( .A1(n5742), .A2(n5740), .ZN(n5752) );
  INV_X1 U7292 ( .A(n5752), .ZN(n5743) );
  XNOR2_X1 U7293 ( .A(n5742), .B(n5741), .ZN(n7229) );
  OR2_X1 U7294 ( .A1(n7226), .A2(n5753), .ZN(n7256) );
  XNOR2_X1 U7295 ( .A(n10154), .B(n5816), .ZN(n5755) );
  NAND2_X1 U7296 ( .A1(n8348), .A2(n8023), .ZN(n5756) );
  NAND2_X1 U7297 ( .A1(n5755), .A2(n5756), .ZN(n7254) );
  INV_X1 U7298 ( .A(n7254), .ZN(n5754) );
  OR2_X1 U7299 ( .A1(n7256), .A2(n5754), .ZN(n7214) );
  XNOR2_X1 U7300 ( .A(n8728), .B(n5816), .ZN(n5747) );
  INV_X1 U7301 ( .A(n5747), .ZN(n5745) );
  NOR2_X1 U7302 ( .A1(n7440), .A2(n8232), .ZN(n5746) );
  INV_X1 U7303 ( .A(n5746), .ZN(n5744) );
  XNOR2_X1 U7304 ( .A(n8723), .B(n5819), .ZN(n5762) );
  NAND2_X1 U7305 ( .A1(n8346), .A2(n8023), .ZN(n5763) );
  NAND2_X1 U7306 ( .A1(n5762), .A2(n5763), .ZN(n5767) );
  INV_X1 U7307 ( .A(n5767), .ZN(n5768) );
  AND2_X1 U7308 ( .A1(n5747), .A2(n5746), .ZN(n7217) );
  INV_X1 U7309 ( .A(n7217), .ZN(n5760) );
  INV_X1 U7310 ( .A(n5748), .ZN(n5751) );
  INV_X1 U7311 ( .A(n5749), .ZN(n5750) );
  NAND2_X1 U7312 ( .A1(n5751), .A2(n5750), .ZN(n7227) );
  OR2_X1 U7313 ( .A1(n5754), .A2(n7257), .ZN(n5759) );
  INV_X1 U7314 ( .A(n5755), .ZN(n5758) );
  INV_X1 U7315 ( .A(n5756), .ZN(n5757) );
  NAND2_X1 U7316 ( .A1(n5758), .A2(n5757), .ZN(n7255) );
  AND2_X1 U7317 ( .A1(n5759), .A2(n7255), .ZN(n7215) );
  AND2_X1 U7318 ( .A1(n5760), .A2(n7215), .ZN(n5761) );
  INV_X1 U7319 ( .A(n5762), .ZN(n5765) );
  INV_X1 U7320 ( .A(n5763), .ZN(n5764) );
  NAND2_X1 U7321 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  AND2_X1 U7322 ( .A1(n5767), .A2(n5766), .ZN(n7362) );
  XNOR2_X1 U7323 ( .A(n8718), .B(n5819), .ZN(n7523) );
  NAND2_X1 U7324 ( .A1(n8345), .A2(n8023), .ZN(n5769) );
  AND2_X1 U7325 ( .A1(n7523), .A2(n5769), .ZN(n5773) );
  XNOR2_X1 U7326 ( .A(n8712), .B(n5816), .ZN(n5774) );
  NAND2_X1 U7327 ( .A1(n8344), .A2(n8023), .ZN(n5775) );
  XNOR2_X1 U7328 ( .A(n5774), .B(n5775), .ZN(n7536) );
  INV_X1 U7329 ( .A(n7523), .ZN(n5770) );
  INV_X1 U7330 ( .A(n5769), .ZN(n7526) );
  NAND2_X1 U7331 ( .A1(n5770), .A2(n7526), .ZN(n5771) );
  AND2_X1 U7332 ( .A1(n7536), .A2(n5771), .ZN(n5772) );
  INV_X1 U7333 ( .A(n5774), .ZN(n5776) );
  NAND2_X1 U7334 ( .A1(n5776), .A2(n5775), .ZN(n5777) );
  NAND2_X1 U7335 ( .A1(n7539), .A2(n5777), .ZN(n7517) );
  XNOR2_X1 U7336 ( .A(n8709), .B(n5819), .ZN(n5779) );
  NAND2_X1 U7337 ( .A1(n8595), .A2(n8023), .ZN(n5778) );
  XNOR2_X1 U7338 ( .A(n5779), .B(n5778), .ZN(n7516) );
  XNOR2_X1 U7339 ( .A(n8592), .B(n5819), .ZN(n5783) );
  NAND2_X1 U7340 ( .A1(n8343), .A2(n8023), .ZN(n5781) );
  XNOR2_X1 U7341 ( .A(n5783), .B(n5781), .ZN(n7547) );
  NAND2_X1 U7342 ( .A1(n7548), .A2(n7547), .ZN(n5785) );
  INV_X1 U7343 ( .A(n5781), .ZN(n5782) );
  NAND2_X1 U7344 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  XNOR2_X1 U7345 ( .A(n8698), .B(n5819), .ZN(n5786) );
  NAND2_X1 U7346 ( .A1(n8596), .A2(n8023), .ZN(n5787) );
  NAND2_X1 U7347 ( .A1(n5786), .A2(n5787), .ZN(n5792) );
  INV_X1 U7348 ( .A(n5786), .ZN(n5789) );
  INV_X1 U7349 ( .A(n5787), .ZN(n5788) );
  NAND2_X1 U7350 ( .A1(n5789), .A2(n5788), .ZN(n5790) );
  NAND2_X1 U7351 ( .A1(n5792), .A2(n5790), .ZN(n8268) );
  XNOR2_X1 U7352 ( .A(n8692), .B(n5816), .ZN(n5794) );
  NOR2_X1 U7353 ( .A1(n8553), .A2(n8232), .ZN(n5793) );
  XNOR2_X1 U7354 ( .A(n5794), .B(n5793), .ZN(n8304) );
  NAND2_X1 U7355 ( .A1(n5794), .A2(n5793), .ZN(n5795) );
  XNOR2_X1 U7356 ( .A(n8687), .B(n5816), .ZN(n5798) );
  NAND2_X1 U7357 ( .A1(n8568), .A2(n8023), .ZN(n5796) );
  XNOR2_X1 U7358 ( .A(n5798), .B(n5796), .ZN(n8277) );
  NAND2_X1 U7359 ( .A1(n8276), .A2(n8277), .ZN(n5800) );
  INV_X1 U7360 ( .A(n5796), .ZN(n5797) );
  NAND2_X1 U7361 ( .A1(n5798), .A2(n5797), .ZN(n5799) );
  XNOR2_X1 U7362 ( .A(n8681), .B(n5819), .ZN(n5802) );
  NAND2_X1 U7363 ( .A1(n5512), .A2(n8023), .ZN(n8319) );
  INV_X1 U7364 ( .A(n5801), .ZN(n5803) );
  NAND2_X1 U7365 ( .A1(n5803), .A2(n5802), .ZN(n5804) );
  XNOR2_X1 U7366 ( .A(n8522), .B(n5816), .ZN(n5805) );
  NOR2_X1 U7367 ( .A1(n4491), .A2(n8232), .ZN(n8295) );
  INV_X1 U7368 ( .A(n8295), .ZN(n5809) );
  INV_X1 U7369 ( .A(n8296), .ZN(n5807) );
  NOR2_X1 U7370 ( .A1(n5806), .A2(n5805), .ZN(n8292) );
  OAI21_X1 U7371 ( .B1(n8295), .B2(n5807), .A(n8292), .ZN(n5808) );
  OAI21_X1 U7372 ( .B1(n8296), .B2(n5809), .A(n5808), .ZN(n5810) );
  NAND2_X1 U7373 ( .A1(n8508), .A2(n8023), .ZN(n8282) );
  XNOR2_X1 U7374 ( .A(n8339), .B(n5819), .ZN(n5813) );
  AND2_X1 U7375 ( .A1(n8458), .A2(n8023), .ZN(n5812) );
  NAND2_X1 U7376 ( .A1(n5813), .A2(n5812), .ZN(n5814) );
  OAI21_X1 U7377 ( .B1(n5813), .B2(n5812), .A(n5814), .ZN(n8329) );
  INV_X1 U7378 ( .A(n5814), .ZN(n5815) );
  XNOR2_X1 U7379 ( .A(n8654), .B(n5816), .ZN(n5818) );
  AND2_X1 U7380 ( .A1(n8341), .A2(n8023), .ZN(n5817) );
  NAND2_X1 U7381 ( .A1(n5818), .A2(n5817), .ZN(n5826) );
  OAI21_X1 U7382 ( .B1(n5818), .B2(n5817), .A(n5826), .ZN(n8250) );
  INV_X1 U7383 ( .A(n5825), .ZN(n8253) );
  NAND2_X1 U7384 ( .A1(n8459), .A2(n8023), .ZN(n5820) );
  XNOR2_X1 U7385 ( .A(n5820), .B(n5819), .ZN(n5821) );
  XNOR2_X1 U7386 ( .A(n8649), .B(n5821), .ZN(n5828) );
  INV_X1 U7387 ( .A(n5828), .ZN(n5824) );
  NAND2_X1 U7388 ( .A1(n5822), .A2(n6397), .ZN(n5823) );
  NOR2_X1 U7389 ( .A1(n6398), .A2(n5823), .ZN(n5830) );
  NAND2_X1 U7390 ( .A1(n5830), .A2(n10081), .ZN(n5839) );
  INV_X1 U7391 ( .A(n8316), .ZN(n8321) );
  NAND3_X1 U7392 ( .A1(n8253), .A2(n5824), .A3(n5023), .ZN(n5845) );
  NAND3_X1 U7393 ( .A1(n5825), .A2(n8321), .A3(n5828), .ZN(n5844) );
  INV_X1 U7394 ( .A(n5826), .ZN(n5827) );
  NAND3_X1 U7395 ( .A1(n5828), .A2(n5827), .A3(n8321), .ZN(n5843) );
  NAND2_X1 U7396 ( .A1(n5650), .A2(n10097), .ZN(n6406) );
  INV_X1 U7397 ( .A(n10081), .ZN(n5829) );
  OAI21_X1 U7398 ( .B1(n5839), .B2(n6406), .A(n8604), .ZN(n8237) );
  INV_X1 U7399 ( .A(n8435), .ZN(n5838) );
  INV_X1 U7400 ( .A(n5830), .ZN(n5832) );
  NAND2_X1 U7401 ( .A1(n5832), .A2(n5831), .ZN(n5836) );
  INV_X1 U7402 ( .A(n5983), .ZN(n5833) );
  AND3_X1 U7403 ( .A1(n5834), .A2(n5863), .A3(n5833), .ZN(n5835) );
  NAND2_X1 U7404 ( .A1(n5836), .A2(n5835), .ZN(n6295) );
  NAND2_X1 U7405 ( .A1(n6295), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8307) );
  OAI22_X1 U7406 ( .A1(n5838), .A2(n8307), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5837), .ZN(n5841) );
  NOR2_X1 U7407 ( .A1(n5839), .A2(n8224), .ZN(n8286) );
  NAND2_X1 U7408 ( .A1(n8286), .A2(n10065), .ZN(n8309) );
  NAND2_X1 U7409 ( .A1(n8286), .A2(n10066), .ZN(n8310) );
  OAI22_X1 U7410 ( .A1(n8442), .A2(n8309), .B1(n8441), .B2(n8310), .ZN(n5840)
         );
  AOI211_X1 U7411 ( .C1(n8649), .C2(n8314), .A(n5841), .B(n5840), .ZN(n5842)
         );
  NAND4_X1 U7412 ( .A1(n5845), .A2(n5844), .A3(n5843), .A4(n5842), .ZN(
        P2_U3222) );
  NOR2_X2 U7413 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5847) );
  NOR2_X2 U7414 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5846) );
  NAND2_X1 U7415 ( .A1(n5884), .A2(n4430), .ZN(n5917) );
  INV_X1 U7416 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5850) );
  AND4_X2 U7417 ( .A1(n5850), .A2(n4615), .A3(n6436), .A4(n5849), .ZN(n5852)
         );
  NOR2_X1 U7418 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5854) );
  NAND2_X1 U7419 ( .A1(n4460), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5855) );
  XNOR2_X1 U7420 ( .A(n5855), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7421 ( .A1(n4451), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5862) );
  INV_X1 U7422 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U7423 ( .A1(n5862), .A2(n5861), .ZN(n5856) );
  NAND2_X1 U7424 ( .A1(n5856), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5857) );
  XNOR2_X1 U7425 ( .A(n5857), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7426 ( .A1(n5858), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5859) );
  MUX2_X1 U7427 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5859), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5860) );
  AND2_X1 U7428 ( .A1(n5860), .A2(n4460), .ZN(n6152) );
  NAND3_X1 U7429 ( .A1(n6164), .A2(n6165), .A3(n6152), .ZN(n6223) );
  INV_X1 U7430 ( .A(n6223), .ZN(n6227) );
  XNOR2_X1 U7431 ( .A(n5862), .B(n5861), .ZN(n7074) );
  NAND2_X1 U7432 ( .A1(n6227), .A2(n7074), .ZN(n5910) );
  INV_X1 U7433 ( .A(n9833), .ZN(P1_U4006) );
  OR2_X1 U7434 ( .A1(n5863), .A2(n4374), .ZN(n5984) );
  NOR2_X2 U7435 ( .A1(n5984), .A2(n5983), .ZN(P2_U3966) );
  NAND2_X1 U7436 ( .A1(n5864), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5865) );
  XNOR2_X1 U7437 ( .A(n5865), .B(n5013), .ZN(n7844) );
  INV_X1 U7438 ( .A(n7844), .ZN(n7996) );
  INV_X1 U7439 ( .A(n5866), .ZN(n5867) );
  NAND2_X1 U7440 ( .A1(n5867), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5869) );
  XNOR2_X1 U7441 ( .A(n5869), .B(n5868), .ZN(n7967) );
  INV_X1 U7442 ( .A(n7967), .ZN(n7883) );
  AND2_X1 U7443 ( .A1(n7996), .A2(n7883), .ZN(n7845) );
  NAND2_X1 U7444 ( .A1(n7845), .A2(n7074), .ZN(n5870) );
  NAND2_X1 U7445 ( .A1(n5910), .A2(n5870), .ZN(n5913) );
  INV_X1 U7446 ( .A(n5871), .ZN(n5873) );
  NAND4_X1 U7447 ( .A1(n5894), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_IR_REG_28__SCAN_IN), .A4(P1_IR_REG_27__SCAN_IN), .ZN(n5872) );
  OR2_X1 U7448 ( .A1(n5913), .A2(n7279), .ZN(n9804) );
  NAND2_X1 U7449 ( .A1(n9804), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U7450 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5874) );
  NOR2_X1 U7451 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5874), .ZN(n6576) );
  INV_X1 U7452 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5877) );
  NOR2_X1 U7453 ( .A1(n5875), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5923) );
  OR2_X1 U7454 ( .A1(n5923), .A2(n5883), .ZN(n5876) );
  INV_X1 U7455 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5922) );
  XNOR2_X1 U7456 ( .A(n5876), .B(n5922), .ZN(n6509) );
  MUX2_X1 U7457 ( .A(n5877), .B(P1_REG2_REG_6__SCAN_IN), .S(n6509), .Z(n5878)
         );
  INV_X1 U7458 ( .A(n5878), .ZN(n5899) );
  NAND2_X1 U7459 ( .A1(n5875), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5879) );
  XNOR2_X1 U7460 ( .A(n5879), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9860) );
  NOR2_X1 U7461 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9860), .ZN(n5880) );
  AOI21_X1 U7462 ( .B1(n9860), .B2(P1_REG2_REG_5__SCAN_IN), .A(n5880), .ZN(
        n9863) );
  INV_X1 U7463 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5883) );
  NOR2_X1 U7464 ( .A1(n5881), .A2(n5883), .ZN(n5882) );
  MUX2_X1 U7465 ( .A(n5883), .B(n5882), .S(P1_IR_REG_4__SCAN_IN), .Z(n5885) );
  INV_X1 U7466 ( .A(n5875), .ZN(n5884) );
  INV_X1 U7467 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6910) );
  XNOR2_X1 U7468 ( .A(n9844), .B(n6910), .ZN(n9843) );
  NOR2_X1 U7469 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5887) );
  NAND2_X1 U7470 ( .A1(n4626), .A2(n5887), .ZN(n5888) );
  NAND2_X1 U7471 ( .A1(n5888), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5886) );
  XNOR2_X1 U7472 ( .A(n5886), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6336) );
  INV_X1 U7473 ( .A(n6077), .ZN(n9838) );
  NAND2_X1 U7474 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5889) );
  NAND2_X1 U7475 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9815) );
  NAND2_X1 U7476 ( .A1(n6252), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5890) );
  OAI21_X1 U7477 ( .B1(n6252), .B2(P1_REG2_REG_1__SCAN_IN), .A(n5890), .ZN(
        n9814) );
  NOR2_X1 U7478 ( .A1(n9815), .A2(n9814), .ZN(n9813) );
  AOI21_X1 U7479 ( .B1(n6252), .B2(P1_REG2_REG_1__SCAN_IN), .A(n9813), .ZN(
        n9830) );
  INV_X1 U7480 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6748) );
  MUX2_X1 U7481 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6748), .S(n6077), .Z(n9829)
         );
  NOR2_X1 U7482 ( .A1(n9830), .A2(n9829), .ZN(n9828) );
  AOI21_X1 U7483 ( .B1(n9838), .B2(P1_REG2_REG_2__SCAN_IN), .A(n9828), .ZN(
        n6041) );
  NAND2_X1 U7484 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n6336), .ZN(n5891) );
  OAI21_X1 U7485 ( .B1(n6336), .B2(P1_REG2_REG_3__SCAN_IN), .A(n5891), .ZN(
        n6040) );
  NOR2_X1 U7486 ( .A1(n6041), .A2(n6040), .ZN(n6039) );
  NAND2_X1 U7487 ( .A1(n9843), .A2(n9842), .ZN(n5893) );
  OR2_X1 U7488 ( .A1(n9844), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7489 ( .A1(n5893), .A2(n5892), .ZN(n9862) );
  NAND2_X1 U7490 ( .A1(n9863), .A2(n9862), .ZN(n9861) );
  NAND2_X1 U7491 ( .A1(n5894), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U7492 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n5895) );
  NAND2_X1 U7493 ( .A1(n5897), .A2(n5895), .ZN(n5896) );
  XNOR2_X1 U7494 ( .A(n5896), .B(P1_IR_REG_28__SCAN_IN), .ZN(n9800) );
  OR2_X1 U7495 ( .A1(n9800), .A2(P1_U3084), .ZN(n9700) );
  OR2_X1 U7496 ( .A1(n5913), .A2(n9700), .ZN(n5900) );
  XNOR2_X1 U7497 ( .A(n5897), .B(P1_IR_REG_27__SCAN_IN), .ZN(n9802) );
  INV_X1 U7498 ( .A(n9802), .ZN(n9831) );
  NOR2_X1 U7499 ( .A1(n5900), .A2(n9831), .ZN(n9891) );
  INV_X1 U7500 ( .A(n9891), .ZN(n9827) );
  AOI211_X1 U7501 ( .C1(n5899), .C2(n5898), .A(n5938), .B(n9827), .ZN(n5916)
         );
  INV_X1 U7502 ( .A(n5900), .ZN(n5901) );
  NAND2_X1 U7503 ( .A1(n5901), .A2(n9831), .ZN(n9896) );
  INV_X1 U7504 ( .A(n9896), .ZN(n9872) );
  INV_X1 U7505 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6348) );
  XNOR2_X1 U7506 ( .A(n9844), .B(n6348), .ZN(n9847) );
  INV_X1 U7507 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9806) );
  INV_X1 U7508 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7509 ( .A1(n6252), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5902) );
  OAI21_X1 U7510 ( .B1(n6252), .B2(P1_REG1_REG_1__SCAN_IN), .A(n5902), .ZN(
        n9811) );
  NOR3_X1 U7511 ( .A1(n9806), .A2(n6100), .A3(n9811), .ZN(n9810) );
  AOI21_X1 U7512 ( .B1(n6252), .B2(P1_REG1_REG_1__SCAN_IN), .A(n9810), .ZN(
        n9825) );
  INV_X1 U7513 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6264) );
  MUX2_X1 U7514 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6264), .S(n6077), .Z(n9824)
         );
  NOR2_X1 U7515 ( .A1(n9825), .A2(n9824), .ZN(n9823) );
  AOI21_X1 U7516 ( .B1(n9838), .B2(P1_REG1_REG_2__SCAN_IN), .A(n9823), .ZN(
        n6044) );
  NAND2_X1 U7517 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(n6336), .ZN(n5903) );
  OAI21_X1 U7518 ( .B1(n6336), .B2(P1_REG1_REG_3__SCAN_IN), .A(n5903), .ZN(
        n6043) );
  NOR2_X1 U7519 ( .A1(n6044), .A2(n6043), .ZN(n6042) );
  AOI21_X1 U7520 ( .B1(n6336), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6042), .ZN(
        n9846) );
  NOR2_X1 U7521 ( .A1(n9844), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5904) );
  AOI21_X1 U7522 ( .B1(n9847), .B2(n9846), .A(n5904), .ZN(n9855) );
  OR2_X1 U7523 ( .A1(n9860), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7524 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9860), .ZN(n5905) );
  AND2_X1 U7525 ( .A1(n5906), .A2(n5905), .ZN(n9854) );
  AND2_X1 U7526 ( .A1(n9855), .A2(n9854), .ZN(n9857) );
  AOI21_X1 U7527 ( .B1(n9860), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9857), .ZN(
        n5908) );
  INV_X1 U7528 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6501) );
  MUX2_X1 U7529 ( .A(n6501), .B(P1_REG1_REG_6__SCAN_IN), .S(n6509), .Z(n5907)
         );
  NAND2_X1 U7530 ( .A1(n5908), .A2(n5907), .ZN(n5957) );
  OAI21_X1 U7531 ( .B1(n5908), .B2(n5907), .A(n5957), .ZN(n5909) );
  AND2_X1 U7532 ( .A1(n9872), .A2(n5909), .ZN(n5915) );
  INV_X1 U7533 ( .A(P1_U3083), .ZN(n5911) );
  NAND2_X1 U7534 ( .A1(n5911), .A2(n5910), .ZN(n9880) );
  INV_X1 U7535 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9715) );
  AND2_X1 U7536 ( .A1(n9802), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7458) );
  NAND2_X1 U7537 ( .A1(n7458), .A2(n9800), .ZN(n5912) );
  OR2_X1 U7538 ( .A1(n5913), .A2(n5912), .ZN(n9818) );
  OAI22_X1 U7539 ( .A1(n9880), .A2(n9715), .B1(n6509), .B2(n9818), .ZN(n5914)
         );
  OR4_X1 U7540 ( .A1(n6576), .A2(n5916), .A3(n5915), .A4(n5914), .ZN(P1_U3247)
         );
  OR2_X1 U7541 ( .A1(n5945), .A2(n5883), .ZN(n5918) );
  XNOR2_X1 U7542 ( .A(n5918), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7280) );
  NAND2_X1 U7543 ( .A1(n5919), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5920) );
  XNOR2_X1 U7544 ( .A(n5920), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7162) );
  INV_X1 U7545 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7198) );
  NOR2_X1 U7546 ( .A1(n7162), .A2(n7198), .ZN(n5921) );
  AOI21_X1 U7547 ( .B1(n7162), .B2(n7198), .A(n5921), .ZN(n6323) );
  NAND2_X1 U7548 ( .A1(n5923), .A2(n5922), .ZN(n5935) );
  INV_X1 U7549 ( .A(n5935), .ZN(n5925) );
  INV_X1 U7550 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7551 ( .A1(n5925), .A2(n5924), .ZN(n5931) );
  OAI21_X1 U7552 ( .B1(n5933), .B2(P1_IR_REG_9__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U7553 ( .A1(n5929), .A2(n5926), .ZN(n5927) );
  NAND2_X1 U7554 ( .A1(n5927), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5928) );
  XNOR2_X1 U7555 ( .A(n5928), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7034) );
  INV_X1 U7556 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6999) );
  MUX2_X1 U7557 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n6999), .S(n7034), .Z(n6209)
         );
  XNOR2_X1 U7558 ( .A(n5929), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6987) );
  NAND2_X1 U7559 ( .A1(n5933), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5930) );
  XNOR2_X1 U7560 ( .A(n5930), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9899) );
  INV_X1 U7561 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6958) );
  NAND2_X1 U7562 ( .A1(n5931), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5932) );
  MUX2_X1 U7563 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5932), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5934) );
  NAND2_X1 U7564 ( .A1(n5934), .A2(n5933), .ZN(n6627) );
  MUX2_X1 U7565 ( .A(n6958), .B(P1_REG2_REG_8__SCAN_IN), .S(n6627), .Z(n6125)
         );
  NAND2_X1 U7566 ( .A1(n5935), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5936) );
  XNOR2_X1 U7567 ( .A(n5936), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9876) );
  NOR2_X1 U7568 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n9876), .ZN(n5937) );
  AOI21_X1 U7569 ( .B1(n9876), .B2(P1_REG2_REG_7__SCAN_IN), .A(n5937), .ZN(
        n9874) );
  INV_X1 U7570 ( .A(n6509), .ZN(n5958) );
  OAI21_X1 U7571 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n9876), .A(n9873), .ZN(
        n6126) );
  NAND2_X1 U7572 ( .A1(n6125), .A2(n6126), .ZN(n6124) );
  NAND2_X1 U7573 ( .A1(n6627), .A2(n6958), .ZN(n5939) );
  NAND2_X1 U7574 ( .A1(n6124), .A2(n5939), .ZN(n9888) );
  OR2_X1 U7575 ( .A1(n9899), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U7576 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n9899), .ZN(n5940) );
  NAND2_X1 U7577 ( .A1(n5941), .A2(n5940), .ZN(n9887) );
  NAND2_X1 U7578 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n6987), .ZN(n5942) );
  OAI21_X1 U7579 ( .B1(n6987), .B2(P1_REG2_REG_10__SCAN_IN), .A(n5942), .ZN(
        n6196) );
  NAND2_X1 U7580 ( .A1(n6209), .A2(n6208), .ZN(n6207) );
  OAI21_X1 U7581 ( .B1(n7034), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6207), .ZN(
        n6322) );
  NAND2_X1 U7582 ( .A1(n7280), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5943) );
  OAI21_X1 U7583 ( .B1(n7280), .B2(P1_REG2_REG_13__SCAN_IN), .A(n5943), .ZN(
        n6446) );
  NAND2_X1 U7584 ( .A1(n6141), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5948) );
  XNOR2_X1 U7585 ( .A(n5948), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7312) );
  INV_X1 U7586 ( .A(n7312), .ZN(n6970) );
  NOR2_X1 U7587 ( .A1(n5946), .A2(n6970), .ZN(n5947) );
  INV_X1 U7588 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6972) );
  XNOR2_X1 U7589 ( .A(n6970), .B(n5946), .ZN(n6973) );
  NOR2_X1 U7590 ( .A1(n6972), .A2(n6973), .ZN(n6971) );
  NAND2_X1 U7591 ( .A1(n5948), .A2(n9407), .ZN(n5949) );
  NAND2_X1 U7592 ( .A1(n5949), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5950) );
  XNOR2_X1 U7593 ( .A(n5950), .B(n9405), .ZN(n9076) );
  XNOR2_X1 U7594 ( .A(n9069), .B(n9076), .ZN(n5951) );
  INV_X1 U7595 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9344) );
  AOI211_X1 U7596 ( .C1(n5951), .C2(n9344), .A(n9070), .B(n9827), .ZN(n5966)
         );
  INV_X1 U7597 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n5952) );
  NOR2_X1 U7598 ( .A1(n9880), .A2(n5952), .ZN(n5965) );
  INV_X1 U7599 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9771) );
  NOR2_X1 U7600 ( .A1(n6970), .A2(n9771), .ZN(n5953) );
  AOI21_X1 U7601 ( .B1(n9771), .B2(n6970), .A(n5953), .ZN(n6968) );
  INV_X1 U7602 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9777) );
  INV_X1 U7603 ( .A(n7280), .ZN(n6444) );
  NOR2_X1 U7604 ( .A1(n6444), .A2(n9777), .ZN(n5954) );
  AOI21_X1 U7605 ( .B1(n9777), .B2(n6444), .A(n5954), .ZN(n6443) );
  INV_X1 U7606 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9784) );
  INV_X1 U7607 ( .A(n7162), .ZN(n6320) );
  NOR2_X1 U7608 ( .A1(n6320), .A2(n9784), .ZN(n5955) );
  AOI21_X1 U7609 ( .B1(n9784), .B2(n6320), .A(n5955), .ZN(n6318) );
  INV_X1 U7610 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6995) );
  MUX2_X1 U7611 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6995), .S(n7034), .Z(n6212)
         );
  INV_X1 U7612 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6821) );
  MUX2_X1 U7613 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6821), .S(n6987), .Z(n6193)
         );
  INV_X1 U7614 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10045) );
  MUX2_X1 U7615 ( .A(n10045), .B(P1_REG1_REG_8__SCAN_IN), .S(n6627), .Z(n6129)
         );
  OR2_X1 U7616 ( .A1(n9876), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5959) );
  NOR2_X1 U7617 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n9876), .ZN(n5956) );
  AOI21_X1 U7618 ( .B1(n9876), .B2(P1_REG1_REG_7__SCAN_IN), .A(n5956), .ZN(
        n9868) );
  OAI21_X1 U7619 ( .B1(n5958), .B2(P1_REG1_REG_6__SCAN_IN), .A(n5957), .ZN(
        n9869) );
  NAND2_X1 U7620 ( .A1(n9868), .A2(n9869), .ZN(n9867) );
  AND2_X1 U7621 ( .A1(n5959), .A2(n9867), .ZN(n6128) );
  NAND2_X1 U7622 ( .A1(n6129), .A2(n6128), .ZN(n6127) );
  INV_X1 U7623 ( .A(n6627), .ZN(n6130) );
  NAND2_X1 U7624 ( .A1(n6130), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5960) );
  NOR2_X1 U7625 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n9899), .ZN(n5961) );
  AOI21_X1 U7626 ( .B1(n9899), .B2(P1_REG1_REG_9__SCAN_IN), .A(n5961), .ZN(
        n9884) );
  NAND2_X1 U7627 ( .A1(n9883), .A2(n9884), .ZN(n9882) );
  OAI21_X1 U7628 ( .B1(n9899), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9882), .ZN(
        n6192) );
  NAND2_X1 U7629 ( .A1(n6193), .A2(n6192), .ZN(n6191) );
  OAI21_X1 U7630 ( .B1(n6987), .B2(P1_REG1_REG_10__SCAN_IN), .A(n6191), .ZN(
        n6211) );
  NAND2_X1 U7631 ( .A1(n6212), .A2(n6211), .ZN(n6210) );
  OAI21_X1 U7632 ( .B1(n7034), .B2(P1_REG1_REG_11__SCAN_IN), .A(n6210), .ZN(
        n6319) );
  NAND2_X1 U7633 ( .A1(n6318), .A2(n6319), .ZN(n6317) );
  OAI21_X1 U7634 ( .B1(n7162), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6317), .ZN(
        n6442) );
  NAND2_X1 U7635 ( .A1(n6443), .A2(n6442), .ZN(n6441) );
  OAI21_X1 U7636 ( .B1(n7280), .B2(P1_REG1_REG_13__SCAN_IN), .A(n6441), .ZN(
        n6967) );
  NAND2_X1 U7637 ( .A1(n6968), .A2(n6967), .ZN(n6966) );
  OAI21_X1 U7638 ( .B1(n7312), .B2(P1_REG1_REG_14__SCAN_IN), .A(n6966), .ZN(
        n9075) );
  XNOR2_X1 U7639 ( .A(n9076), .B(n9075), .ZN(n5962) );
  INV_X1 U7640 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9289) );
  NOR2_X1 U7641 ( .A1(n9289), .A2(n5962), .ZN(n9077) );
  AOI211_X1 U7642 ( .C1(n5962), .C2(n9289), .A(n9077), .B(n9896), .ZN(n5964)
         );
  NAND2_X1 U7643 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9041) );
  OAI21_X1 U7644 ( .B1(n9818), .B2(n9076), .A(n9041), .ZN(n5963) );
  OR4_X1 U7645 ( .A1(n5966), .A2(n5965), .A3(n5964), .A4(n5963), .ZN(P1_U3256)
         );
  MUX2_X1 U7646 ( .A(n5967), .B(P2_REG2_REG_16__SCAN_IN), .S(n8376), .Z(n8381)
         );
  MUX2_X1 U7647 ( .A(n5397), .B(P2_REG2_REG_14__SCAN_IN), .S(n8365), .Z(n5968)
         );
  INV_X1 U7648 ( .A(n5968), .ZN(n8360) );
  XNOR2_X1 U7649 ( .A(n6018), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n6780) );
  XNOR2_X1 U7650 ( .A(n6673), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n6669) );
  INV_X1 U7651 ( .A(n6621), .ZN(n5975) );
  INV_X1 U7652 ( .A(n6088), .ZN(n6685) );
  INV_X1 U7653 ( .A(n6082), .ZN(n6697) );
  XNOR2_X1 U7654 ( .A(n6082), .B(n5969), .ZN(n6693) );
  INV_X1 U7655 ( .A(n6074), .ZN(n9750) );
  INV_X1 U7656 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10059) );
  NAND2_X1 U7657 ( .A1(n9738), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5970) );
  AOI21_X1 U7658 ( .B1(n9738), .B2(P2_REG2_REG_1__SCAN_IN), .A(n9733), .ZN(
        n9747) );
  INV_X1 U7659 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5971) );
  MUX2_X1 U7660 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n5971), .S(n6074), .Z(n9746)
         );
  NOR2_X1 U7661 ( .A1(n9747), .A2(n9746), .ZN(n9745) );
  AOI21_X1 U7662 ( .B1(n9750), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9745), .ZN(
        n6062) );
  NAND2_X1 U7663 ( .A1(n5998), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5972) );
  OAI21_X1 U7664 ( .B1(n5998), .B2(P2_REG2_REG_3__SCAN_IN), .A(n5972), .ZN(
        n6061) );
  NOR2_X1 U7665 ( .A1(n6062), .A2(n6061), .ZN(n6060) );
  NAND2_X1 U7666 ( .A1(n6661), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5973) );
  OAI21_X1 U7667 ( .B1(n6661), .B2(P2_REG2_REG_5__SCAN_IN), .A(n5973), .ZN(
        n6657) );
  AOI21_X1 U7668 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n6661), .A(n6656), .ZN(
        n6682) );
  MUX2_X1 U7669 ( .A(n6765), .B(P2_REG2_REG_6__SCAN_IN), .S(n6088), .Z(n5974)
         );
  INV_X1 U7670 ( .A(n5974), .ZN(n6681) );
  NOR2_X1 U7671 ( .A1(n6682), .A2(n6681), .ZN(n6680) );
  AOI21_X1 U7672 ( .B1(n6685), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6680), .ZN(
        n6051) );
  MUX2_X1 U7673 ( .A(n9464), .B(P2_REG2_REG_7__SCAN_IN), .S(n6007), .Z(n6050)
         );
  NOR2_X1 U7674 ( .A1(n6051), .A2(n6050), .ZN(n6049) );
  AOI21_X1 U7675 ( .B1(n6007), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6049), .ZN(
        n6612) );
  MUX2_X1 U7676 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7090), .S(n6621), .Z(n6611)
         );
  NOR2_X1 U7677 ( .A1(n6612), .A2(n6611), .ZN(n6610) );
  AOI21_X1 U7678 ( .B1(n5975), .B2(P2_REG2_REG_8__SCAN_IN), .A(n6610), .ZN(
        n6706) );
  NAND2_X1 U7679 ( .A1(n6709), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5976) );
  OAI21_X1 U7680 ( .B1(n6709), .B2(P2_REG2_REG_9__SCAN_IN), .A(n5976), .ZN(
        n6705) );
  NOR2_X1 U7681 ( .A1(n6706), .A2(n6705), .ZN(n6704) );
  INV_X1 U7682 ( .A(n6016), .ZN(n6565) );
  AOI22_X1 U7683 ( .A1(n6016), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n5338), .B2(
        n6565), .ZN(n6559) );
  OAI21_X1 U7684 ( .B1(n6016), .B2(P2_REG2_REG_11__SCAN_IN), .A(n6557), .ZN(
        n6781) );
  NOR2_X1 U7685 ( .A1(n7098), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5977) );
  AOI21_X1 U7686 ( .B1(n7098), .B2(P2_REG2_REG_13__SCAN_IN), .A(n5977), .ZN(
        n7100) );
  OAI21_X1 U7687 ( .B1(n7098), .B2(P2_REG2_REG_13__SCAN_IN), .A(n7099), .ZN(
        n8361) );
  NAND2_X1 U7688 ( .A1(n8360), .A2(n8361), .ZN(n8359) );
  OAI21_X1 U7689 ( .B1(n8365), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8359), .ZN(
        n5978) );
  NAND2_X1 U7690 ( .A1(n7515), .A2(n5978), .ZN(n5980) );
  XNOR2_X1 U7691 ( .A(n5979), .B(n5978), .ZN(n7511) );
  NAND2_X1 U7692 ( .A1(n8393), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5981) );
  OAI21_X1 U7693 ( .B1(n8393), .B2(P2_REG2_REG_17__SCAN_IN), .A(n5981), .ZN(
        n5987) );
  NOR2_X1 U7694 ( .A1(n5988), .A2(n5987), .ZN(n8387) );
  INV_X2 U7695 ( .A(P2_U3966), .ZN(n8358) );
  INV_X1 U7696 ( .A(n5982), .ZN(n6029) );
  NAND2_X1 U7697 ( .A1(n10081), .A2(n6029), .ZN(n5985) );
  NAND2_X1 U7698 ( .A1(n5983), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8230) );
  NAND3_X1 U7699 ( .A1(n5985), .A2(n8230), .A3(n5984), .ZN(n5986) );
  NAND2_X1 U7700 ( .A1(n5986), .A2(n6031), .ZN(n6025) );
  NAND2_X1 U7701 ( .A1(n8358), .A2(n6025), .ZN(n5989) );
  NAND2_X1 U7702 ( .A1(n5989), .A2(n8225), .ZN(n8411) );
  NOR2_X1 U7703 ( .A1(n8411), .A2(n5639), .ZN(n10055) );
  AOI211_X1 U7704 ( .C1(n5988), .C2(n5987), .A(n8387), .B(n9744), .ZN(n6038)
         );
  AND2_X1 U7705 ( .A1(n5989), .A2(n5639), .ZN(n10053) );
  INV_X1 U7706 ( .A(n10053), .ZN(n8402) );
  INV_X1 U7707 ( .A(n8393), .ZN(n5990) );
  NOR2_X1 U7708 ( .A1(n8402), .A2(n5990), .ZN(n6037) );
  XNOR2_X1 U7709 ( .A(n8376), .B(n5991), .ZN(n8374) );
  XNOR2_X1 U7710 ( .A(n8365), .B(n5992), .ZN(n8367) );
  INV_X1 U7711 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10173) );
  MUX2_X1 U7712 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n10173), .S(n6673), .Z(n6665) );
  NAND2_X1 U7713 ( .A1(n6709), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6013) );
  OR2_X1 U7714 ( .A1(n6621), .A2(n6008), .ZN(n6010) );
  OR2_X1 U7715 ( .A1(n6661), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U7716 ( .A1(n6661), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6004) );
  AND2_X1 U7717 ( .A1(n5993), .A2(n6004), .ZN(n6653) );
  XNOR2_X1 U7718 ( .A(n6082), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n6689) );
  NAND2_X1 U7719 ( .A1(n5998), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6001) );
  INV_X1 U7720 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10164) );
  INV_X1 U7721 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5994) );
  NOR2_X1 U7722 ( .A1(n6072), .A2(n5994), .ZN(n5996) );
  INV_X1 U7723 ( .A(n5996), .ZN(n5995) );
  OAI21_X1 U7724 ( .B1(n9738), .B2(P2_REG1_REG_1__SCAN_IN), .A(n5995), .ZN(
        n9731) );
  NOR3_X1 U7725 ( .A1(n10059), .A2(n10164), .A3(n9731), .ZN(n9730) );
  NOR2_X1 U7726 ( .A1(n9730), .A2(n5996), .ZN(n9743) );
  INV_X1 U7727 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5997) );
  MUX2_X1 U7728 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n5997), .S(n6074), .Z(n9742)
         );
  NOR2_X1 U7729 ( .A1(n9743), .A2(n9742), .ZN(n9741) );
  AOI21_X1 U7730 ( .B1(n9750), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9741), .ZN(
        n6065) );
  INV_X1 U7731 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5999) );
  MUX2_X1 U7732 ( .A(n5999), .B(P2_REG1_REG_3__SCAN_IN), .S(n5998), .Z(n6064)
         );
  NOR2_X1 U7733 ( .A1(n6065), .A2(n6064), .ZN(n6063) );
  INV_X1 U7734 ( .A(n6063), .ZN(n6000) );
  NAND2_X1 U7735 ( .A1(n6001), .A2(n6000), .ZN(n6688) );
  NAND2_X1 U7736 ( .A1(n6689), .A2(n6688), .ZN(n6687) );
  OR2_X1 U7737 ( .A1(n6082), .A2(n6002), .ZN(n6003) );
  NAND2_X1 U7738 ( .A1(n6687), .A2(n6003), .ZN(n6652) );
  NAND2_X1 U7739 ( .A1(n6653), .A2(n6652), .ZN(n6651) );
  AND2_X1 U7740 ( .A1(n6651), .A2(n6004), .ZN(n6677) );
  MUX2_X1 U7741 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6005), .S(n6088), .Z(n6676)
         );
  NOR2_X1 U7742 ( .A1(n6677), .A2(n6676), .ZN(n6675) );
  AOI21_X1 U7743 ( .B1(n6685), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6675), .ZN(
        n6054) );
  NAND2_X1 U7744 ( .A1(n6007), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6006) );
  OAI21_X1 U7745 ( .B1(n6007), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6006), .ZN(
        n6053) );
  NOR2_X1 U7746 ( .A1(n6054), .A2(n6053), .ZN(n6052) );
  AOI21_X1 U7747 ( .B1(n6007), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6052), .ZN(
        n6616) );
  MUX2_X1 U7748 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6008), .S(n6621), .Z(n6615)
         );
  NOR2_X1 U7749 ( .A1(n6616), .A2(n6615), .ZN(n6614) );
  INV_X1 U7750 ( .A(n6614), .ZN(n6009) );
  AND2_X1 U7751 ( .A1(n6010), .A2(n6009), .ZN(n6700) );
  MUX2_X1 U7752 ( .A(n6011), .B(P2_REG1_REG_9__SCAN_IN), .S(n6709), .Z(n6701)
         );
  NOR2_X1 U7753 ( .A1(n6700), .A2(n6701), .ZN(n6699) );
  INV_X1 U7754 ( .A(n6699), .ZN(n6012) );
  NAND2_X1 U7755 ( .A1(n6013), .A2(n6012), .ZN(n6664) );
  NAND2_X1 U7756 ( .A1(n6665), .A2(n6664), .ZN(n6663) );
  NAND2_X1 U7757 ( .A1(n6673), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7758 ( .A1(n6663), .A2(n6014), .ZN(n6561) );
  INV_X1 U7759 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6015) );
  MUX2_X1 U7760 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n6015), .S(n6016), .Z(n6562)
         );
  NAND2_X1 U7761 ( .A1(n6561), .A2(n6562), .ZN(n6560) );
  NAND2_X1 U7762 ( .A1(n6016), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6017) );
  AND2_X1 U7763 ( .A1(n6560), .A2(n6017), .ZN(n6785) );
  INV_X1 U7764 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6019) );
  MUX2_X1 U7765 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6019), .S(n6018), .Z(n6786)
         );
  NAND2_X1 U7766 ( .A1(n6785), .A2(n6786), .ZN(n6790) );
  INV_X1 U7767 ( .A(n6018), .ZN(n6795) );
  NAND2_X1 U7768 ( .A1(n6795), .A2(n6019), .ZN(n6020) );
  NAND2_X1 U7769 ( .A1(n6790), .A2(n6020), .ZN(n7104) );
  MUX2_X1 U7770 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n6021), .S(n7098), .Z(n7105)
         );
  NAND2_X1 U7771 ( .A1(n7104), .A2(n7105), .ZN(n7103) );
  OR2_X1 U7772 ( .A1(n7098), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U7773 ( .A1(n7103), .A2(n6022), .ZN(n8368) );
  NAND2_X1 U7774 ( .A1(n8367), .A2(n8368), .ZN(n8366) );
  OAI21_X1 U7775 ( .B1(n8365), .B2(P2_REG1_REG_14__SCAN_IN), .A(n8366), .ZN(
        n6023) );
  NOR2_X1 U7776 ( .A1(n7515), .A2(n6023), .ZN(n6024) );
  XNOR2_X1 U7777 ( .A(n7515), .B(n6023), .ZN(n7507) );
  NOR2_X1 U7778 ( .A1(n7506), .A2(n7507), .ZN(n7505) );
  NOR2_X1 U7779 ( .A1(n6024), .A2(n7505), .ZN(n8375) );
  NAND2_X1 U7780 ( .A1(n8374), .A2(n8375), .ZN(n8373) );
  OAI21_X1 U7781 ( .B1(n8376), .B2(P2_REG1_REG_16__SCAN_IN), .A(n8373), .ZN(
        n6028) );
  XNOR2_X1 U7782 ( .A(n8393), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n6027) );
  NOR2_X1 U7783 ( .A1(n6027), .A2(n6028), .ZN(n8392) );
  INV_X1 U7784 ( .A(n6025), .ZN(n6026) );
  AND2_X1 U7785 ( .A1(n7533), .A2(n6026), .ZN(n10050) );
  INV_X1 U7786 ( .A(n10050), .ZN(n10051) );
  AOI211_X1 U7787 ( .C1(n6028), .C2(n6027), .A(n8392), .B(n10051), .ZN(n6036)
         );
  NAND2_X1 U7788 ( .A1(n6031), .A2(n6029), .ZN(n6030) );
  NAND2_X1 U7789 ( .A1(n6030), .A2(n10081), .ZN(n6033) );
  OR2_X1 U7790 ( .A1(n6031), .A2(n8230), .ZN(n6032) );
  INV_X1 U7791 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9367) );
  NAND2_X1 U7792 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(n4374), .ZN(n6034) );
  OAI21_X1 U7793 ( .B1(n8417), .B2(n9367), .A(n6034), .ZN(n6035) );
  OR4_X1 U7794 ( .A1(n6038), .A2(n6037), .A3(n6036), .A4(n6035), .ZN(P2_U3262)
         );
  AND2_X1 U7795 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6386) );
  AOI211_X1 U7796 ( .C1(n6041), .C2(n6040), .A(n6039), .B(n9827), .ZN(n6048)
         );
  AOI211_X1 U7797 ( .C1(n6044), .C2(n6043), .A(n6042), .B(n9896), .ZN(n6047)
         );
  INV_X1 U7798 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6045) );
  INV_X1 U7799 ( .A(n6336), .ZN(n6079) );
  OAI22_X1 U7800 ( .A1(n9880), .A2(n6045), .B1(n6079), .B2(n9818), .ZN(n6046)
         );
  OR4_X1 U7801 ( .A1(n6386), .A2(n6048), .A3(n6047), .A4(n6046), .ZN(P1_U3244)
         );
  AOI211_X1 U7802 ( .C1(n6051), .C2(n6050), .A(n6049), .B(n9744), .ZN(n6059)
         );
  NOR2_X1 U7803 ( .A1(n8402), .A2(n6091), .ZN(n6058) );
  AOI211_X1 U7804 ( .C1(n6054), .C2(n6053), .A(n6052), .B(n10051), .ZN(n6057)
         );
  INV_X1 U7805 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9718) );
  NAND2_X1 U7806 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3152), .ZN(n6055) );
  OAI21_X1 U7807 ( .B1(n8417), .B2(n9718), .A(n6055), .ZN(n6056) );
  OR4_X1 U7808 ( .A1(n6059), .A2(n6058), .A3(n6057), .A4(n6056), .ZN(P2_U3252)
         );
  AOI211_X1 U7809 ( .C1(n6062), .C2(n6061), .A(n6060), .B(n9744), .ZN(n6071)
         );
  NOR2_X1 U7810 ( .A1(n8402), .A2(n6080), .ZN(n6070) );
  AOI211_X1 U7811 ( .C1(n6065), .C2(n6064), .A(n6063), .B(n10051), .ZN(n6069)
         );
  INV_X1 U7812 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7813 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(n4374), .ZN(n6066) );
  OAI21_X1 U7814 ( .B1(n8417), .B2(n6067), .A(n6066), .ZN(n6068) );
  OR4_X1 U7815 ( .A1(n6071), .A2(n6070), .A3(n6069), .A4(n6068), .ZN(P2_U3248)
         );
  NOR2_X1 U7816 ( .A1(n4498), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8756) );
  INV_X1 U7817 ( .A(n8756), .ZN(n8761) );
  AND2_X1 U7818 ( .A1(n4498), .A2(n4374), .ZN(n7077) );
  OAI222_X1 U7819 ( .A1(n8761), .A2(n6073), .B1(n4385), .B2(n6255), .C1(
        P2_U3152), .C2(n6072), .ZN(P2_U3357) );
  OAI222_X1 U7820 ( .A1(n8761), .A2(n6075), .B1(n4385), .B2(n6271), .C1(n4374), 
        .C2(n6074), .ZN(P2_U3356) );
  NAND2_X1 U7821 ( .A1(n4498), .A2(P1_U3084), .ZN(n9698) );
  INV_X1 U7822 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7823 ( .A1(n7743), .A2(P1_U3084), .ZN(n8009) );
  INV_X1 U7824 ( .A(n6252), .ZN(n9819) );
  OAI222_X1 U7825 ( .A1(n9698), .A2(n6076), .B1(n9695), .B2(n6255), .C1(
        P1_U3084), .C2(n9819), .ZN(P1_U3352) );
  CLKBUF_X1 U7826 ( .A(n8009), .Z(n9695) );
  OAI222_X1 U7827 ( .A1(n9698), .A2(n6078), .B1(n9695), .B2(n6271), .C1(
        P1_U3084), .C2(n6077), .ZN(P1_U3351) );
  OAI222_X1 U7828 ( .A1(n9698), .A2(n9409), .B1(n9695), .B2(n6339), .C1(
        P1_U3084), .C2(n6079), .ZN(P1_U3350) );
  OAI222_X1 U7829 ( .A1(n8761), .A2(n6081), .B1(n4385), .B2(n6339), .C1(
        P2_U3152), .C2(n6080), .ZN(P2_U3355) );
  OAI222_X1 U7830 ( .A1(n8761), .A2(n6083), .B1(n4385), .B2(n6359), .C1(n4374), 
        .C2(n6082), .ZN(P2_U3354) );
  INV_X1 U7831 ( .A(n9698), .ZN(n9699) );
  AOI22_X1 U7832 ( .A1(n9844), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n9699), .ZN(n6084) );
  OAI21_X1 U7833 ( .B1(n6359), .B2(n9695), .A(n6084), .ZN(P1_U3349) );
  AOI22_X1 U7834 ( .A1(n9860), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9699), .ZN(n6085) );
  OAI21_X1 U7835 ( .B1(n6486), .B2(n8009), .A(n6085), .ZN(P1_U3348) );
  OAI222_X1 U7836 ( .A1(n8761), .A2(n6087), .B1(n4385), .B2(n6486), .C1(
        P2_U3152), .C2(n6086), .ZN(P2_U3353) );
  OAI222_X1 U7837 ( .A1(n9698), .A2(n6510), .B1(n9695), .B2(n6508), .C1(
        P1_U3084), .C2(n6509), .ZN(P1_U3347) );
  OAI222_X1 U7838 ( .A1(n8761), .A2(n6089), .B1(n4385), .B2(n6508), .C1(n4374), 
        .C2(n6088), .ZN(P2_U3352) );
  AOI22_X1 U7839 ( .A1(n9876), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9699), .ZN(n6090) );
  OAI21_X1 U7840 ( .B1(n6474), .B2(n8009), .A(n6090), .ZN(P1_U3346) );
  OAI222_X1 U7841 ( .A1(n8761), .A2(n6092), .B1(n4385), .B2(n6474), .C1(
        P2_U3152), .C2(n6091), .ZN(P2_U3351) );
  OAI222_X1 U7842 ( .A1(n8761), .A2(n6093), .B1(n4385), .B2(n6626), .C1(n4374), 
        .C2(n6621), .ZN(P2_U3350) );
  OAI222_X1 U7843 ( .A1(n9698), .A2(n9302), .B1(n9695), .B2(n6626), .C1(
        P1_U3084), .C2(n6627), .ZN(P1_U3345) );
  INV_X1 U7844 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6108) );
  INV_X1 U7845 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6094) );
  NAND2_X2 U7846 ( .A1(n6099), .A2(n6101), .ZN(n6349) );
  INV_X1 U7847 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6098) );
  INV_X1 U7848 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9801) );
  INV_X1 U7849 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7850 ( .A1(n8942), .A2(P1_U4006), .ZN(n6107) );
  OAI21_X1 U7851 ( .B1(P1_U4006), .B2(n6108), .A(n6107), .ZN(P1_U3555) );
  INV_X1 U7852 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6116) );
  INV_X1 U7853 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6109) );
  NOR2_X1 U7854 ( .A1(n7703), .A2(n6109), .ZN(n6114) );
  INV_X1 U7855 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6110) );
  NOR2_X1 U7856 ( .A1(n7679), .A2(n6110), .ZN(n6113) );
  INV_X1 U7857 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6111) );
  NOR2_X1 U7858 ( .A1(n7719), .A2(n6111), .ZN(n6112) );
  OR3_X1 U7859 ( .A1(n6114), .A2(n6113), .A3(n6112), .ZN(n8004) );
  NAND2_X1 U7860 ( .A1(n8004), .A2(P1_U4006), .ZN(n6115) );
  OAI21_X1 U7861 ( .B1(P1_U4006), .B2(n6116), .A(n6115), .ZN(P1_U3586) );
  INV_X1 U7862 ( .A(n6814), .ZN(n6119) );
  AOI22_X1 U7863 ( .A1(n9899), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9699), .ZN(n6117) );
  OAI21_X1 U7864 ( .B1(n6119), .B2(n8009), .A(n6117), .ZN(P1_U3344) );
  OAI222_X1 U7865 ( .A1(n8761), .A2(n6120), .B1(n4385), .B2(n6119), .C1(n6118), 
        .C2(n4374), .ZN(P2_U3349) );
  INV_X1 U7866 ( .A(n6986), .ZN(n6123) );
  AOI22_X1 U7867 ( .A1(n6987), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9699), .ZN(n6121) );
  OAI21_X1 U7868 ( .B1(n6123), .B2(n8009), .A(n6121), .ZN(P1_U3343) );
  AOI22_X1 U7869 ( .A1(n6673), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n8756), .ZN(n6122) );
  OAI21_X1 U7870 ( .B1(n6123), .B2(n4385), .A(n6122), .ZN(P2_U3348) );
  INV_X1 U7871 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6136) );
  OAI21_X1 U7872 ( .B1(n6126), .B2(n6125), .A(n6124), .ZN(n6134) );
  OAI21_X1 U7873 ( .B1(n6129), .B2(n6128), .A(n6127), .ZN(n6132) );
  INV_X1 U7874 ( .A(n9818), .ZN(n9898) );
  INV_X1 U7875 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9324) );
  NOR2_X1 U7876 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9324), .ZN(n6647) );
  AOI21_X1 U7877 ( .B1(n9898), .B2(n6130), .A(n6647), .ZN(n6131) );
  OAI21_X1 U7878 ( .B1(n9896), .B2(n6132), .A(n6131), .ZN(n6133) );
  AOI21_X1 U7879 ( .B1(n9891), .B2(n6134), .A(n6133), .ZN(n6135) );
  OAI21_X1 U7880 ( .B1(n9880), .B2(n6136), .A(n6135), .ZN(P1_U3249) );
  INV_X1 U7881 ( .A(n8417), .ZN(n10056) );
  NOR2_X1 U7882 ( .A1(n10056), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7883 ( .A(n7033), .ZN(n6138) );
  OAI222_X1 U7884 ( .A1(n8761), .A2(n6137), .B1(n4385), .B2(n6138), .C1(n6565), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U7885 ( .A(n7034), .ZN(n6215) );
  OAI222_X1 U7886 ( .A1(n9698), .A2(n9329), .B1(n6215), .B2(P1_U3084), .C1(
        n9695), .C2(n6138), .ZN(P1_U3342) );
  INV_X1 U7887 ( .A(n7161), .ZN(n6182) );
  AOI22_X1 U7888 ( .A1(n7162), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9699), .ZN(n6139) );
  OAI21_X1 U7889 ( .B1(n6182), .B2(n8009), .A(n6139), .ZN(P1_U3341) );
  NAND2_X1 U7890 ( .A1(n8358), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6140) );
  OAI21_X1 U7891 ( .B1(n8553), .B2(n8358), .A(n6140), .ZN(P2_U3572) );
  OAI21_X1 U7892 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U7893 ( .A1(n6312), .A2(n6143), .ZN(n6146) );
  INV_X1 U7894 ( .A(n6146), .ZN(n6144) );
  INV_X1 U7895 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7896 ( .A1(n6146), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7897 ( .A1(n7992), .A2(n7845), .ZN(n6149) );
  AND2_X1 U7898 ( .A1(n6223), .A2(n7074), .ZN(n6148) );
  AND2_X1 U7899 ( .A1(n6149), .A2(n6148), .ZN(n6373) );
  AND2_X1 U7900 ( .A1(n6373), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6735) );
  INV_X1 U7901 ( .A(n6152), .ZN(n7335) );
  NAND2_X1 U7902 ( .A1(n7335), .A2(P1_B_REG_SCAN_IN), .ZN(n6150) );
  MUX2_X1 U7903 ( .A(n6150), .B(P1_B_REG_SCAN_IN), .S(n6165), .Z(n6151) );
  NAND2_X1 U7904 ( .A1(n6151), .A2(n6164), .ZN(n9692) );
  OAI22_X1 U7905 ( .A1(n9692), .A2(P1_D_REG_1__SCAN_IN), .B1(n6164), .B2(n6152), .ZN(n6732) );
  AND2_X1 U7906 ( .A1(n7844), .A2(n7967), .ZN(n6232) );
  INV_X1 U7907 ( .A(n6235), .ZN(n6153) );
  AND3_X1 U7908 ( .A1(n6735), .A2(n6732), .A3(n6153), .ZN(n7268) );
  INV_X1 U7909 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9942) );
  INV_X1 U7910 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9939) );
  INV_X1 U7911 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9938) );
  INV_X1 U7912 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9946) );
  NAND4_X1 U7913 ( .A1(n9942), .A2(n9939), .A3(n9938), .A4(n9946), .ZN(n6156)
         );
  NOR4_X1 U7914 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6154) );
  INV_X1 U7915 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9965) );
  NAND2_X1 U7916 ( .A1(n6154), .A2(n9965), .ZN(n9420) );
  INV_X1 U7917 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9943) );
  INV_X1 U7918 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9945) );
  INV_X1 U7919 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n9950) );
  INV_X1 U7920 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9948) );
  NAND4_X1 U7921 ( .A1(n9943), .A2(n9945), .A3(n9950), .A4(n9948), .ZN(n6155)
         );
  NOR4_X1 U7922 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n6156), .A3(n9420), .A4(n6155), .ZN(n6162) );
  NOR4_X1 U7923 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6160) );
  NOR4_X1 U7924 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6159) );
  NOR4_X1 U7925 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6158) );
  NOR4_X1 U7926 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n6157) );
  AND4_X1 U7927 ( .A1(n6160), .A2(n6159), .A3(n6158), .A4(n6157), .ZN(n6161)
         );
  AND2_X1 U7928 ( .A1(n6162), .A2(n6161), .ZN(n6163) );
  NOR2_X1 U7929 ( .A1(n9692), .A2(n6163), .ZN(n6220) );
  INV_X1 U7930 ( .A(n6220), .ZN(n6734) );
  INV_X1 U7931 ( .A(n6164), .ZN(n7338) );
  INV_X1 U7932 ( .A(n6165), .ZN(n7124) );
  NAND2_X1 U7933 ( .A1(n7338), .A2(n7124), .ZN(n9693) );
  OAI21_X1 U7934 ( .B1(n9692), .B2(P1_D_REG_0__SCAN_IN), .A(n9693), .ZN(n6733)
         );
  AND2_X1 U7935 ( .A1(n6734), .A2(n6733), .ZN(n6166) );
  AND2_X2 U7936 ( .A1(n7268), .A2(n6166), .ZN(n10037) );
  INV_X1 U7937 ( .A(SI_0_), .ZN(n6168) );
  INV_X1 U7938 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6167) );
  OAI21_X1 U7939 ( .B1(n4498), .B2(n6168), .A(n6167), .ZN(n6170) );
  NAND2_X1 U7940 ( .A1(n6170), .A2(n6169), .ZN(n9703) );
  INV_X1 U7941 ( .A(n6232), .ZN(n6234) );
  INV_X1 U7942 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7943 ( .A1(n7635), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6175) );
  NAND4_X1 U7944 ( .A1(n6176), .A2(n6175), .A3(n6174), .A4(n6173), .ZN(n6722)
         );
  NAND2_X1 U7945 ( .A1(n8942), .A2(n9929), .ZN(n7968) );
  AND2_X1 U7946 ( .A1(n6801), .A2(n7968), .ZN(n7855) );
  INV_X1 U7947 ( .A(n6737), .ZN(n6179) );
  NAND2_X1 U7948 ( .A1(n9124), .A2(n7996), .ZN(n6246) );
  INV_X1 U7949 ( .A(n6246), .ZN(n6178) );
  AND2_X1 U7950 ( .A1(n6179), .A2(n6178), .ZN(n6876) );
  NOR3_X1 U7951 ( .A1(n7855), .A2(n6232), .A3(n6876), .ZN(n6180) );
  AOI21_X1 U7952 ( .B1(n9911), .B2(n6723), .A(n6180), .ZN(n9932) );
  OAI21_X1 U7953 ( .B1(n9929), .B2(n6234), .A(n9932), .ZN(n9674) );
  NAND2_X1 U7954 ( .A1(n9674), .A2(n10037), .ZN(n6181) );
  OAI21_X1 U7955 ( .B1(n10037), .B2(n6102), .A(n6181), .ZN(P1_U3454) );
  OAI222_X1 U7956 ( .A1(n8761), .A2(n9440), .B1(n4385), .B2(n6182), .C1(n4374), 
        .C2(n6795), .ZN(P2_U3346) );
  INV_X1 U7957 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9459) );
  INV_X1 U7958 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7959 ( .A1(n5206), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7960 ( .A1(n5204), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6183) );
  OAI211_X1 U7961 ( .C1(n6186), .C2(n6185), .A(n6184), .B(n6183), .ZN(n8420)
         );
  NAND2_X1 U7962 ( .A1(n8420), .A2(P2_U3966), .ZN(n6187) );
  OAI21_X1 U7963 ( .B1(P2_U3966), .B2(n9459), .A(n6187), .ZN(P2_U3583) );
  INV_X1 U7964 ( .A(n7278), .ZN(n6190) );
  AOI22_X1 U7965 ( .A1(n7280), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9699), .ZN(n6188) );
  OAI21_X1 U7966 ( .B1(n6190), .B2(n8009), .A(n6188), .ZN(P1_U3340) );
  AOI22_X1 U7967 ( .A1(n7098), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n8756), .ZN(n6189) );
  OAI21_X1 U7968 ( .B1(n6190), .B2(n4385), .A(n6189), .ZN(P2_U3345) );
  INV_X1 U7969 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6202) );
  OAI21_X1 U7970 ( .B1(n6193), .B2(n6192), .A(n6191), .ZN(n6200) );
  INV_X1 U7971 ( .A(n6987), .ZN(n6194) );
  NAND2_X1 U7972 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3084), .ZN(n6994) );
  OAI21_X1 U7973 ( .B1(n9818), .B2(n6194), .A(n6994), .ZN(n6199) );
  AOI211_X1 U7974 ( .C1(n6197), .C2(n6196), .A(n6195), .B(n9827), .ZN(n6198)
         );
  AOI211_X1 U7975 ( .C1(n9872), .C2(n6200), .A(n6199), .B(n6198), .ZN(n6201)
         );
  OAI21_X1 U7976 ( .B1(n9880), .B2(n6202), .A(n6201), .ZN(P1_U3251) );
  INV_X1 U7977 ( .A(n7311), .ZN(n6205) );
  AOI22_X1 U7978 ( .A1(n8365), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n8756), .ZN(n6203) );
  OAI21_X1 U7979 ( .B1(n6205), .B2(n4385), .A(n6203), .ZN(P2_U3344) );
  OAI222_X1 U7980 ( .A1(n9695), .A2(n6205), .B1(n6970), .B2(P1_U3084), .C1(
        n6204), .C2(n9698), .ZN(P1_U3339) );
  INV_X1 U7981 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6796) );
  NAND2_X1 U7982 ( .A1(n8568), .A2(P2_U3966), .ZN(n6206) );
  OAI21_X1 U7983 ( .B1(P2_U3966), .B2(n6796), .A(n6206), .ZN(P2_U3573) );
  INV_X1 U7984 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6219) );
  OAI21_X1 U7985 ( .B1(n6209), .B2(n6208), .A(n6207), .ZN(n6217) );
  OAI21_X1 U7986 ( .B1(n6212), .B2(n6211), .A(n6210), .ZN(n6213) );
  NAND2_X1 U7987 ( .A1(n9872), .A2(n6213), .ZN(n6214) );
  NAND2_X1 U7988 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3084), .ZN(n7068) );
  OAI211_X1 U7989 ( .C1(n9818), .C2(n6215), .A(n6214), .B(n7068), .ZN(n6216)
         );
  AOI21_X1 U7990 ( .B1(n9891), .B2(n6217), .A(n6216), .ZN(n6218) );
  OAI21_X1 U7991 ( .B1(n9880), .B2(n6219), .A(n6218), .ZN(P1_U3252) );
  INV_X1 U7992 ( .A(n6723), .ZN(n6244) );
  OR2_X1 U7993 ( .A1(n6733), .A2(n6220), .ZN(n7266) );
  NOR2_X1 U7994 ( .A1(n7266), .A2(n6732), .ZN(n6375) );
  AND2_X1 U7995 ( .A1(n7074), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6221) );
  AND2_X1 U7996 ( .A1(n6223), .A2(n6221), .ZN(n9691) );
  AND2_X1 U7997 ( .A1(n6375), .A2(n9691), .ZN(n6231) );
  AND2_X1 U7998 ( .A1(n6231), .A2(n6876), .ZN(n6277) );
  NAND2_X1 U7999 ( .A1(n6277), .A2(n9800), .ZN(n9046) );
  AND2_X1 U8000 ( .A1(n6737), .A2(n6223), .ZN(n6226) );
  OR2_X1 U8001 ( .A1(n7992), .A2(n7996), .ZN(n6222) );
  AND2_X4 U8002 ( .A1(n6226), .A2(n6222), .ZN(n8924) );
  NOR2_X2 U8003 ( .A1(n6737), .A2(n6227), .ZN(n6356) );
  INV_X1 U8004 ( .A(n6356), .ZN(n6224) );
  OAI22_X1 U8005 ( .A1(n9929), .A2(n6224), .B1(n6223), .B2(n9806), .ZN(n6225)
         );
  AOI22_X1 U8006 ( .A1(n6750), .A2(n6226), .B1(n6227), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n6228) );
  NAND2_X1 U8007 ( .A1(n6229), .A2(n6228), .ZN(n6245) );
  OAI21_X1 U8008 ( .B1(n6230), .B2(n6245), .A(n6249), .ZN(n9832) );
  INV_X1 U8009 ( .A(n6231), .ZN(n6233) );
  NAND2_X1 U8010 ( .A1(n7992), .A2(n6232), .ZN(n10027) );
  INV_X1 U8011 ( .A(n7845), .ZN(n6742) );
  NAND2_X1 U8012 ( .A1(n10027), .A2(n6742), .ZN(n6374) );
  INV_X1 U8013 ( .A(n9052), .ZN(n8982) );
  OR2_X1 U8014 ( .A1(n6177), .A2(n6234), .ZN(n6237) );
  INV_X1 U8015 ( .A(n6237), .ZN(n9200) );
  NAND3_X1 U8016 ( .A1(n6375), .A2(n9691), .A3(n9200), .ZN(n6236) );
  NAND2_X1 U8017 ( .A1(n6236), .A2(n9936), .ZN(n9050) );
  AOI22_X1 U8018 ( .A1(n9832), .A2(n8982), .B1(n6750), .B2(n9050), .ZN(n6243)
         );
  INV_X1 U8019 ( .A(n10027), .ZN(n10004) );
  INV_X1 U8020 ( .A(n6375), .ZN(n6241) );
  INV_X1 U8021 ( .A(n6876), .ZN(n6238) );
  NAND2_X1 U8022 ( .A1(n6238), .A2(n6237), .ZN(n6239) );
  AND2_X1 U8023 ( .A1(n6239), .A2(n9691), .ZN(n6240) );
  NAND2_X1 U8024 ( .A1(n6241), .A2(n6240), .ZN(n6377) );
  OAI211_X1 U8025 ( .C1(n6375), .C2(n10004), .A(n6735), .B(n6377), .ZN(n8941)
         );
  NAND2_X1 U8026 ( .A1(n8941), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6242) );
  OAI211_X1 U8027 ( .C1(n6244), .C2(n9046), .A(n6243), .B(n6242), .ZN(P1_U3230) );
  AND2_X2 U8028 ( .A1(n6737), .A2(n6246), .ZN(n8922) );
  NAND2_X1 U8029 ( .A1(n4578), .A2(n6247), .ZN(n6248) );
  NAND2_X1 U8030 ( .A1(n6723), .A2(n6356), .ZN(n6257) );
  NAND2_X1 U8031 ( .A1(n6475), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U8032 ( .A1(n7279), .A2(n6252), .ZN(n6253) );
  OAI211_X1 U8033 ( .C1(n6255), .C2(n6813), .A(n6254), .B(n6253), .ZN(n6721)
         );
  NAND2_X1 U8034 ( .A1(n8940), .A2(n6226), .ZN(n6256) );
  NAND2_X1 U8035 ( .A1(n6257), .A2(n6256), .ZN(n6258) );
  AND2_X1 U8036 ( .A1(n8940), .A2(n8919), .ZN(n6259) );
  AOI21_X1 U8037 ( .B1(n6723), .B2(n8924), .A(n6259), .ZN(n8938) );
  INV_X1 U8038 ( .A(n6260), .ZN(n6261) );
  NAND2_X1 U8039 ( .A1(n6262), .A2(n6261), .ZN(n6263) );
  NAND2_X1 U8040 ( .A1(n8937), .A2(n6263), .ZN(n6330) );
  INV_X1 U8041 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6753) );
  OR2_X1 U8042 ( .A1(n6349), .A2(n6753), .ZN(n6267) );
  OR2_X1 U8043 ( .A1(n6280), .A2(n6264), .ZN(n6265) );
  NAND4_X2 U8044 ( .A1(n6268), .A2(n6267), .A3(n6266), .A4(n6265), .ZN(n6727)
         );
  NAND2_X1 U8045 ( .A1(n6727), .A2(n8919), .ZN(n6273) );
  NAND2_X1 U8046 ( .A1(n6475), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U8047 ( .A1(n7279), .A2(n9838), .ZN(n6269) );
  OAI211_X2 U8048 ( .C1(n6271), .C2(n6813), .A(n6270), .B(n6269), .ZN(n9975)
         );
  NAND2_X1 U8049 ( .A1(n9975), .A2(n8918), .ZN(n6272) );
  NAND2_X1 U8050 ( .A1(n6273), .A2(n6272), .ZN(n6274) );
  XNOR2_X1 U8051 ( .A(n6274), .B(n6247), .ZN(n6331) );
  AND2_X1 U8052 ( .A1(n9975), .A2(n8919), .ZN(n6275) );
  AOI21_X1 U8053 ( .B1(n6727), .B2(n8924), .A(n6275), .ZN(n6332) );
  XNOR2_X1 U8054 ( .A(n6331), .B(n6332), .ZN(n6329) );
  XOR2_X1 U8055 ( .A(n6330), .B(n6329), .Z(n6287) );
  AOI22_X1 U8056 ( .A1(n8941), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n9050), .B2(
        n9975), .ZN(n6286) );
  INV_X1 U8057 ( .A(n9800), .ZN(n6276) );
  NAND2_X1 U8058 ( .A1(n6277), .A2(n6276), .ZN(n9043) );
  INV_X1 U8059 ( .A(n9043), .ZN(n8943) );
  INV_X1 U8060 ( .A(n9046), .ZN(n9021) );
  INV_X1 U8061 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6278) );
  OR2_X1 U8062 ( .A1(n7679), .A2(n6278), .ZN(n6284) );
  OR2_X1 U8063 ( .A1(n6349), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U8064 ( .A1(n6350), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6282) );
  INV_X1 U8065 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6279) );
  OR2_X1 U8066 ( .A1(n6280), .A2(n6279), .ZN(n6281) );
  AOI22_X1 U8067 ( .A1(n8943), .A2(n6723), .B1(n9021), .B2(n6866), .ZN(n6285)
         );
  OAI211_X1 U8068 ( .C1(n6287), .C2(n9052), .A(n6286), .B(n6285), .ZN(P1_U3235) );
  INV_X1 U8069 ( .A(n7483), .ZN(n6300) );
  NAND2_X1 U8070 ( .A1(n6288), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6289) );
  XNOR2_X1 U8071 ( .A(n6289), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9092) );
  INV_X1 U8072 ( .A(n9092), .ZN(n9083) );
  OAI222_X1 U8073 ( .A1(n9695), .A2(n6300), .B1(n9083), .B2(P1_U3084), .C1(
        n6290), .C2(n9698), .ZN(P1_U3337) );
  INV_X1 U8074 ( .A(n6292), .ZN(n6293) );
  AOI21_X1 U8075 ( .B1(n6291), .B2(n6294), .A(n6293), .ZN(n6299) );
  OR2_X1 U8076 ( .A1(n6295), .A2(P2_U3152), .ZN(n8236) );
  AOI22_X1 U8077 ( .A1(n8314), .A2(n6296), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8236), .ZN(n6298) );
  INV_X1 U8078 ( .A(n8310), .ZN(n6777) );
  INV_X1 U8079 ( .A(n8309), .ZN(n6305) );
  AOI22_X1 U8080 ( .A1(n6777), .A2(n10067), .B1(n6305), .B2(n10064), .ZN(n6297) );
  OAI211_X1 U8081 ( .C1(n6299), .C2(n8316), .A(n6298), .B(n6297), .ZN(P2_U3224) );
  INV_X1 U8082 ( .A(n8376), .ZN(n6301) );
  OAI222_X1 U8083 ( .A1(P2_U3152), .A2(n6301), .B1(n4385), .B2(n6300), .C1(
        n9288), .C2(n8761), .ZN(P2_U3342) );
  XNOR2_X1 U8084 ( .A(n6303), .B(n6302), .ZN(n6308) );
  AOI22_X1 U8085 ( .A1(n8314), .A2(n6458), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n8236), .ZN(n6307) );
  AOI22_X1 U8086 ( .A1(n6777), .A2(n6304), .B1(n6305), .B2(n8357), .ZN(n6306)
         );
  OAI211_X1 U8087 ( .C1(n6308), .C2(n8316), .A(n6307), .B(n6306), .ZN(P2_U3239) );
  INV_X1 U8088 ( .A(n7412), .ZN(n6310) );
  OAI222_X1 U8089 ( .A1(n9698), .A2(n6309), .B1(n9695), .B2(n6310), .C1(
        P1_U3084), .C2(n9076), .ZN(P1_U3338) );
  OAI222_X1 U8090 ( .A1(n8761), .A2(n6311), .B1(n4385), .B2(n6310), .C1(
        P2_U3152), .C2(n7515), .ZN(P2_U3343) );
  INV_X1 U8091 ( .A(n7567), .ZN(n6315) );
  XNOR2_X1 U8092 ( .A(n6312), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9109) );
  AOI22_X1 U8093 ( .A1(n9109), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9699), .ZN(n6313) );
  OAI21_X1 U8094 ( .B1(n6315), .B2(n8009), .A(n6313), .ZN(P1_U3336) );
  AOI22_X1 U8095 ( .A1(n8393), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n8756), .ZN(n6314) );
  OAI21_X1 U8096 ( .B1(n6315), .B2(n4385), .A(n6314), .ZN(P2_U3341) );
  NAND2_X1 U8097 ( .A1(n8358), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6316) );
  OAI21_X1 U8098 ( .B1(n8442), .B2(n8358), .A(n6316), .ZN(P2_U3581) );
  INV_X1 U8099 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6328) );
  OAI21_X1 U8100 ( .B1(n6319), .B2(n6318), .A(n6317), .ZN(n6326) );
  NAND2_X1 U8101 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n7179) );
  OAI21_X1 U8102 ( .B1(n9818), .B2(n6320), .A(n7179), .ZN(n6325) );
  AOI211_X1 U8103 ( .C1(n6323), .C2(n6322), .A(n6321), .B(n9827), .ZN(n6324)
         );
  AOI211_X1 U8104 ( .C1(n9872), .C2(n6326), .A(n6325), .B(n6324), .ZN(n6327)
         );
  OAI21_X1 U8105 ( .B1(n9880), .B2(n6328), .A(n6327), .ZN(P1_U3253) );
  NAND2_X1 U8106 ( .A1(n6330), .A2(n6329), .ZN(n6335) );
  INV_X1 U8107 ( .A(n6331), .ZN(n6333) );
  NAND2_X1 U8108 ( .A1(n6333), .A2(n6332), .ZN(n6334) );
  NAND2_X1 U8109 ( .A1(n6335), .A2(n6334), .ZN(n6383) );
  NAND2_X1 U8110 ( .A1(n6866), .A2(n8919), .ZN(n6341) );
  NAND2_X1 U8111 ( .A1(n6475), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U8112 ( .A1(n7279), .A2(n6336), .ZN(n6337) );
  NAND2_X1 U8113 ( .A1(n6865), .A2(n8918), .ZN(n6340) );
  NAND2_X1 U8114 ( .A1(n6341), .A2(n6340), .ZN(n6342) );
  XNOR2_X1 U8115 ( .A(n6342), .B(n6247), .ZN(n6344) );
  AND2_X1 U8116 ( .A1(n6865), .A2(n8919), .ZN(n6343) );
  AOI21_X1 U8117 ( .B1(n6866), .B2(n8924), .A(n6343), .ZN(n6345) );
  XNOR2_X1 U8118 ( .A(n6344), .B(n6345), .ZN(n6384) );
  INV_X1 U8119 ( .A(n6344), .ZN(n6346) );
  NAND2_X1 U8120 ( .A1(n6346), .A2(n6345), .ZN(n6347) );
  XNOR2_X1 U8121 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6909) );
  OR2_X1 U8122 ( .A1(n6349), .A2(n6909), .ZN(n6354) );
  NAND2_X1 U8123 ( .A1(n6350), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6352) );
  OR2_X1 U8124 ( .A1(n7679), .A2(n6910), .ZN(n6351) );
  NAND2_X1 U8125 ( .A1(n9912), .A2(n8925), .ZN(n6361) );
  NAND2_X1 U8126 ( .A1(n6475), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U8127 ( .A1(n7279), .A2(n9844), .ZN(n6357) );
  OAI211_X1 U8128 ( .C1(n6359), .C2(n6813), .A(n6358), .B(n6357), .ZN(n6915)
         );
  NAND2_X1 U8129 ( .A1(n6915), .A2(n8918), .ZN(n6360) );
  NAND2_X1 U8130 ( .A1(n6361), .A2(n6360), .ZN(n6362) );
  XNOR2_X1 U8131 ( .A(n6362), .B(n8922), .ZN(n6492) );
  AND2_X1 U8132 ( .A1(n6915), .A2(n8919), .ZN(n6363) );
  AOI21_X1 U8133 ( .B1(n9912), .B2(n8924), .A(n6363), .ZN(n6493) );
  XNOR2_X1 U8134 ( .A(n6492), .B(n6493), .ZN(n6364) );
  XNOR2_X1 U8135 ( .A(n6483), .B(n6364), .ZN(n6382) );
  AND2_X1 U8136 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9849) );
  INV_X1 U8137 ( .A(n9050), .ZN(n9024) );
  INV_X1 U8138 ( .A(n6915), .ZN(n9989) );
  NOR2_X1 U8139 ( .A1(n9024), .A2(n9989), .ZN(n6365) );
  AOI211_X1 U8140 ( .C1(n8943), .C2(n6866), .A(n9849), .B(n6365), .ZN(n6381)
         );
  AOI21_X1 U8141 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6366) );
  NOR2_X1 U8142 ( .A1(n6366), .A2(n6503), .ZN(n6858) );
  NAND2_X1 U8143 ( .A1(n7700), .A2(n6858), .ZN(n6372) );
  INV_X1 U8144 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6367) );
  OR2_X1 U8145 ( .A1(n7703), .A2(n6367), .ZN(n6371) );
  INV_X1 U8146 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6860) );
  OR2_X1 U8147 ( .A1(n7679), .A2(n6860), .ZN(n6370) );
  INV_X1 U8148 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6368) );
  OR2_X1 U8149 ( .A1(n7719), .A2(n6368), .ZN(n6369) );
  OAI21_X1 U8150 ( .B1(n6375), .B2(n6374), .A(n6373), .ZN(n6376) );
  NAND2_X1 U8151 ( .A1(n6376), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6378) );
  INV_X1 U8152 ( .A(n9045), .ZN(n6544) );
  INV_X1 U8153 ( .A(n6909), .ZN(n6379) );
  AOI22_X1 U8154 ( .A1(n9021), .A2(n9068), .B1(n6544), .B2(n6379), .ZN(n6380)
         );
  OAI211_X1 U8155 ( .C1(n6382), .C2(n9052), .A(n6381), .B(n6380), .ZN(P1_U3228) );
  XOR2_X1 U8156 ( .A(n6383), .B(n6384), .Z(n6389) );
  NOR2_X1 U8157 ( .A1(n9024), .A2(n9982), .ZN(n6385) );
  AOI211_X1 U8158 ( .C1(n8943), .C2(n6727), .A(n6386), .B(n6385), .ZN(n6388)
         );
  INV_X1 U8159 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9922) );
  AOI22_X1 U8160 ( .A1(n9021), .A2(n9912), .B1(n6544), .B2(n9922), .ZN(n6387)
         );
  OAI211_X1 U8161 ( .C1(n6389), .C2(n9052), .A(n6388), .B(n6387), .ZN(P1_U3216) );
  XNOR2_X1 U8162 ( .A(n6391), .B(n6390), .ZN(n6395) );
  AOI22_X1 U8163 ( .A1(n8356), .A2(n10065), .B1(n10066), .B2(n10064), .ZN(
        n6427) );
  INV_X1 U8164 ( .A(n6427), .ZN(n6392) );
  AOI22_X1 U8165 ( .A1(n6392), .A2(n8286), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3152), .ZN(n6394) );
  INV_X1 U8166 ( .A(n8307), .ZN(n8336) );
  INV_X1 U8167 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6428) );
  AOI22_X1 U8168 ( .A1(n6433), .A2(n8314), .B1(n8336), .B2(n6428), .ZN(n6393)
         );
  OAI211_X1 U8169 ( .C1(n6395), .C2(n8316), .A(n6394), .B(n6393), .ZN(P2_U3220) );
  NAND2_X1 U8170 ( .A1(n10067), .A2(n4505), .ZN(n8231) );
  NAND2_X1 U8171 ( .A1(n10062), .A2(n8231), .ZN(n10098) );
  AOI22_X1 U8172 ( .A1(n10098), .A2(n10061), .B1(n10065), .B2(n6304), .ZN(
        n10100) );
  INV_X1 U8173 ( .A(n6396), .ZN(n6400) );
  NOR2_X1 U8174 ( .A1(n6398), .A2(n6397), .ZN(n6399) );
  NAND2_X1 U8175 ( .A1(n6400), .A2(n6399), .ZN(n6408) );
  OR2_X1 U8176 ( .A1(n6402), .A2(n8615), .ZN(n6421) );
  NAND2_X1 U8177 ( .A1(n8630), .A2(n6421), .ZN(n6403) );
  NAND2_X1 U8178 ( .A1(n6401), .A2(n6403), .ZN(n8557) );
  INV_X1 U8179 ( .A(n8557), .ZN(n10077) );
  OAI22_X1 U8180 ( .A1(n6401), .A2(n10054), .B1(n6404), .B2(n8604), .ZN(n6405)
         );
  AOI21_X1 U8181 ( .B1(n10077), .B2(n10098), .A(n6405), .ZN(n6410) );
  INV_X1 U8182 ( .A(n6406), .ZN(n6407) );
  NAND2_X1 U8183 ( .A1(n6401), .A2(n6407), .ZN(n8639) );
  OR2_X1 U8184 ( .A1(n6408), .A2(n8023), .ZN(n8429) );
  NAND2_X1 U8185 ( .A1(n8639), .A2(n8429), .ZN(n10076) );
  NAND2_X1 U8186 ( .A1(n10076), .A2(n10096), .ZN(n6409) );
  OAI211_X1 U8187 ( .C1(n10100), .C2(n8646), .A(n6410), .B(n6409), .ZN(
        P2_U3296) );
  INV_X1 U8188 ( .A(n7571), .ZN(n6440) );
  AOI22_X1 U8189 ( .A1(n8406), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8756), .ZN(n6411) );
  OAI21_X1 U8190 ( .B1(n6440), .B2(n4385), .A(n6411), .ZN(P2_U3340) );
  INV_X1 U8191 ( .A(n6412), .ZN(n6413) );
  AOI21_X1 U8192 ( .B1(n6415), .B2(n6414), .A(n6413), .ZN(n6419) );
  NAND2_X1 U8193 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(n4374), .ZN(n6690) );
  OAI21_X1 U8194 ( .B1(n8307), .B2(n6596), .A(n6690), .ZN(n6417) );
  INV_X1 U8195 ( .A(n8237), .ZN(n8338) );
  OAI22_X1 U8196 ( .A1(n4383), .A2(n8338), .B1(n8309), .B2(n6762), .ZN(n6416)
         );
  AOI211_X1 U8197 ( .C1(n6777), .C2(n8357), .A(n6417), .B(n6416), .ZN(n6418)
         );
  OAI21_X1 U8198 ( .B1(n6419), .B2(n8316), .A(n6418), .ZN(P2_U3232) );
  XNOR2_X1 U8199 ( .A(n8184), .B(n6420), .ZN(n10111) );
  INV_X1 U8200 ( .A(n6421), .ZN(n6422) );
  NAND2_X1 U8201 ( .A1(n6401), .A2(n6422), .ZN(n8641) );
  INV_X1 U8202 ( .A(n6600), .ZN(n6425) );
  AND3_X1 U8203 ( .A1(n6454), .A2(n6423), .A3(n8044), .ZN(n6424) );
  OAI21_X1 U8204 ( .B1(n6425), .B2(n6424), .A(n10061), .ZN(n6426) );
  OAI211_X1 U8205 ( .C1(n10111), .C2(n8630), .A(n6427), .B(n6426), .ZN(n10113)
         );
  NAND2_X1 U8206 ( .A1(n10113), .A2(n6401), .ZN(n6435) );
  INV_X1 U8207 ( .A(n8639), .ZN(n8619) );
  OAI22_X1 U8208 ( .A1(n6401), .A2(n6429), .B1(n8604), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n6432) );
  AND2_X1 U8209 ( .A1(n6460), .A2(n6433), .ZN(n6430) );
  NOR2_X1 U8210 ( .A1(n10112), .A2(n8429), .ZN(n6431) );
  AOI211_X1 U8211 ( .C1(n8619), .C2(n6433), .A(n6432), .B(n6431), .ZN(n6434)
         );
  OAI211_X1 U8212 ( .C1(n10111), .C2(n8641), .A(n6435), .B(n6434), .ZN(
        P2_U3293) );
  INV_X1 U8213 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U8214 ( .A1(n6312), .A2(n6436), .ZN(n6437) );
  NAND2_X1 U8215 ( .A1(n6437), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6438) );
  XNOR2_X1 U8216 ( .A(n6438), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9119) );
  INV_X1 U8217 ( .A(n9119), .ZN(n6439) );
  OAI222_X1 U8218 ( .A1(n9698), .A2(n9229), .B1(n9695), .B2(n6440), .C1(
        P1_U3084), .C2(n6439), .ZN(P1_U3335) );
  INV_X1 U8219 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6452) );
  OAI21_X1 U8220 ( .B1(n6443), .B2(n6442), .A(n6441), .ZN(n6450) );
  NAND2_X1 U8221 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7293) );
  OAI21_X1 U8222 ( .B1(n9818), .B2(n6444), .A(n7293), .ZN(n6449) );
  AOI211_X1 U8223 ( .C1(n6447), .C2(n6446), .A(n6445), .B(n9827), .ZN(n6448)
         );
  AOI211_X1 U8224 ( .C1(n9872), .C2(n6450), .A(n6449), .B(n6448), .ZN(n6451)
         );
  OAI21_X1 U8225 ( .B1(n9880), .B2(n6452), .A(n6451), .ZN(P1_U3254) );
  XNOR2_X1 U8226 ( .A(n6453), .B(n8187), .ZN(n10109) );
  INV_X1 U8227 ( .A(n10109), .ZN(n6466) );
  INV_X1 U8228 ( .A(n10066), .ZN(n8624) );
  INV_X1 U8229 ( .A(n10061), .ZN(n8612) );
  INV_X1 U8230 ( .A(n6454), .ZN(n6455) );
  AOI21_X1 U8231 ( .B1(n8187), .B2(n6456), .A(n6455), .ZN(n6457) );
  OAI222_X1 U8232 ( .A1(n8622), .A2(n6604), .B1(n8624), .B2(n5200), .C1(n8612), 
        .C2(n6457), .ZN(n10107) );
  NOR2_X1 U8233 ( .A1(n8639), .A2(n10105), .ZN(n6464) );
  NAND2_X1 U8234 ( .A1(n6458), .A2(n10073), .ZN(n6459) );
  NAND2_X1 U8235 ( .A1(n6460), .A2(n6459), .ZN(n10106) );
  OR2_X1 U8236 ( .A1(n6401), .A2(n5971), .ZN(n6462) );
  INV_X1 U8237 ( .A(n8604), .ZN(n10071) );
  NAND2_X1 U8238 ( .A1(n10071), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6461) );
  OAI211_X1 U8239 ( .C1(n10106), .C2(n8429), .A(n6462), .B(n6461), .ZN(n6463)
         );
  AOI211_X1 U8240 ( .C1(n10107), .C2(n6401), .A(n6464), .B(n6463), .ZN(n6465)
         );
  OAI21_X1 U8241 ( .B1(n6466), .B2(n8557), .A(n6465), .ZN(P2_U3294) );
  NAND2_X1 U8242 ( .A1(n6350), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6473) );
  INV_X1 U8243 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6467) );
  OR2_X1 U8244 ( .A1(n7703), .A2(n6467), .ZN(n6472) );
  NAND2_X1 U8245 ( .A1(n6503), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6502) );
  AND2_X1 U8246 ( .A1(n6502), .A2(n6468), .ZN(n6469) );
  OR2_X1 U8247 ( .A1(n6469), .A2(n6527), .ZN(n6887) );
  OR2_X1 U8248 ( .A1(n6349), .A2(n6887), .ZN(n6471) );
  INV_X1 U8249 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6888) );
  OR2_X1 U8250 ( .A1(n7679), .A2(n6888), .ZN(n6470) );
  NAND2_X1 U8251 ( .A1(n9066), .A2(n8925), .ZN(n6480) );
  OR2_X1 U8252 ( .A1(n6474), .A2(n6813), .ZN(n6478) );
  AOI22_X1 U8253 ( .A1(n7748), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9876), .B2(
        n7279), .ZN(n6477) );
  NAND2_X1 U8254 ( .A1(n6926), .A2(n6226), .ZN(n6479) );
  NAND2_X1 U8255 ( .A1(n6480), .A2(n6479), .ZN(n6481) );
  XNOR2_X1 U8256 ( .A(n6481), .B(n8922), .ZN(n6623) );
  AOI22_X1 U8257 ( .A1(n9066), .A2(n8924), .B1(n6926), .B2(n8919), .ZN(n6622)
         );
  XNOR2_X1 U8258 ( .A(n6623), .B(n6622), .ZN(n6526) );
  AND2_X1 U8259 ( .A1(n6492), .A2(n6493), .ZN(n6482) );
  NAND2_X1 U8260 ( .A1(n9068), .A2(n8919), .ZN(n6488) );
  NAND2_X1 U8261 ( .A1(n7748), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6485) );
  NAND2_X1 U8262 ( .A1(n7279), .A2(n9860), .ZN(n6484) );
  OAI211_X1 U8263 ( .C1(n6486), .C2(n6813), .A(n6485), .B(n6484), .ZN(n6883)
         );
  NAND2_X1 U8264 ( .A1(n6883), .A2(n8918), .ZN(n6487) );
  NAND2_X1 U8265 ( .A1(n6488), .A2(n6487), .ZN(n6489) );
  XNOR2_X1 U8266 ( .A(n6489), .B(n6247), .ZN(n6499) );
  NAND2_X1 U8267 ( .A1(n9068), .A2(n8924), .ZN(n6491) );
  NAND2_X1 U8268 ( .A1(n6883), .A2(n8925), .ZN(n6490) );
  NAND2_X1 U8269 ( .A1(n6491), .A2(n6490), .ZN(n6542) );
  AND2_X1 U8270 ( .A1(n6499), .A2(n6542), .ZN(n6497) );
  INV_X1 U8271 ( .A(n6492), .ZN(n6495) );
  INV_X1 U8272 ( .A(n6493), .ZN(n6494) );
  NAND2_X1 U8273 ( .A1(n6495), .A2(n6494), .ZN(n6537) );
  INV_X1 U8274 ( .A(n6499), .ZN(n6539) );
  INV_X1 U8275 ( .A(n6542), .ZN(n6500) );
  NAND2_X1 U8276 ( .A1(n6539), .A2(n6500), .ZN(n6517) );
  NAND2_X1 U8277 ( .A1(n6350), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6507) );
  OR2_X1 U8278 ( .A1(n7703), .A2(n6501), .ZN(n6506) );
  OAI21_X1 U8279 ( .B1(n6503), .B2(P1_REG3_REG_6__SCAN_IN), .A(n6502), .ZN(
        n6945) );
  OR2_X1 U8280 ( .A1(n7679), .A2(n5877), .ZN(n6504) );
  NAND2_X1 U8281 ( .A1(n9067), .A2(n8919), .ZN(n6514) );
  OR2_X1 U8282 ( .A1(n6508), .A2(n6813), .ZN(n6512) );
  OAI22_X1 U8283 ( .A1(n6476), .A2(n6510), .B1(n6628), .B2(n6509), .ZN(n6511)
         );
  NAND2_X1 U8284 ( .A1(n10003), .A2(n8918), .ZN(n6513) );
  NAND2_X1 U8285 ( .A1(n6514), .A2(n6513), .ZN(n6515) );
  XNOR2_X1 U8286 ( .A(n6515), .B(n8922), .ZN(n6518) );
  AND2_X1 U8287 ( .A1(n10003), .A2(n8925), .ZN(n6516) );
  AOI21_X1 U8288 ( .B1(n9067), .B2(n8924), .A(n6516), .ZN(n6519) );
  NAND2_X1 U8289 ( .A1(n6518), .A2(n6519), .ZN(n6573) );
  INV_X1 U8290 ( .A(n6518), .ZN(n6521) );
  INV_X1 U8291 ( .A(n6519), .ZN(n6520) );
  NAND2_X1 U8292 ( .A1(n6521), .A2(n6520), .ZN(n6572) );
  INV_X1 U8293 ( .A(n6625), .ZN(n6524) );
  AOI21_X1 U8294 ( .B1(n6526), .B2(n6525), .A(n6524), .ZN(n6536) );
  NOR2_X1 U8295 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6468), .ZN(n9870) );
  NAND2_X1 U8296 ( .A1(n6350), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6532) );
  OR2_X1 U8297 ( .A1(n7703), .A2(n10045), .ZN(n6531) );
  NAND2_X1 U8298 ( .A1(n6527), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6640) );
  OR2_X1 U8299 ( .A1(n6527), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U8300 ( .A1(n6640), .A2(n6528), .ZN(n6957) );
  OR2_X1 U8301 ( .A1(n6349), .A2(n6957), .ZN(n6530) );
  OR2_X1 U8302 ( .A1(n7679), .A2(n6958), .ZN(n6529) );
  NAND4_X1 U8303 ( .A1(n6532), .A2(n6531), .A3(n6530), .A4(n6529), .ZN(n9065)
         );
  OAI22_X1 U8304 ( .A1(n6919), .A2(n9046), .B1(n9045), .B2(n6887), .ZN(n6533)
         );
  AOI211_X1 U8305 ( .C1(n8943), .C2(n9067), .A(n9870), .B(n6533), .ZN(n6535)
         );
  NAND2_X1 U8306 ( .A1(n9050), .A2(n6926), .ZN(n6534) );
  OAI211_X1 U8307 ( .C1(n6536), .C2(n9052), .A(n6535), .B(n6534), .ZN(P1_U3211) );
  AND2_X1 U8308 ( .A1(n6538), .A2(n6537), .ZN(n6540) );
  NAND2_X1 U8309 ( .A1(n6540), .A2(n6539), .ZN(n6569) );
  OAI21_X1 U8310 ( .B1(n6540), .B2(n6539), .A(n6569), .ZN(n6541) );
  NOR2_X1 U8311 ( .A1(n6541), .A2(n6542), .ZN(n6571) );
  AOI21_X1 U8312 ( .B1(n6542), .B2(n6541), .A(n6571), .ZN(n6547) );
  AND2_X1 U8313 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9859) );
  NOR2_X1 U8314 ( .A1(n9024), .A2(n9999), .ZN(n6543) );
  AOI211_X1 U8315 ( .C1(n8943), .C2(n9912), .A(n9859), .B(n6543), .ZN(n6546)
         );
  AOI22_X1 U8316 ( .A1(n9021), .A2(n9067), .B1(n6544), .B2(n6858), .ZN(n6545)
         );
  OAI211_X1 U8317 ( .C1(n6547), .C2(n9052), .A(n6546), .B(n6545), .ZN(P1_U3225) );
  XNOR2_X1 U8318 ( .A(n6549), .B(n6548), .ZN(n6554) );
  OAI22_X1 U8319 ( .A1(n6550), .A2(n8624), .B1(n6841), .B2(n8622), .ZN(n6588)
         );
  AOI22_X1 U8320 ( .A1(n6588), .A2(n8286), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        n4374), .ZN(n6553) );
  INV_X1 U8321 ( .A(n6551), .ZN(n6590) );
  AOI22_X1 U8322 ( .A1(n6584), .A2(n8314), .B1(n8336), .B2(n6590), .ZN(n6552)
         );
  OAI211_X1 U8323 ( .C1(n6554), .C2(n8316), .A(n6553), .B(n6552), .ZN(P2_U3229) );
  INV_X1 U8324 ( .A(n7581), .ZN(n6556) );
  OAI222_X1 U8325 ( .A1(n9698), .A2(n6555), .B1(n9695), .B2(n6556), .C1(
        P1_U3084), .C2(n9124), .ZN(P1_U3334) );
  OAI222_X1 U8326 ( .A1(n8761), .A2(n9221), .B1(n4385), .B2(n6556), .C1(n4374), 
        .C2(n8615), .ZN(P2_U3339) );
  OAI21_X1 U8327 ( .B1(n6559), .B2(n6558), .A(n6557), .ZN(n6567) );
  AOI22_X1 U8328 ( .A1(n10056), .A2(P2_ADDR_REG_11__SCAN_IN), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(P2_U3152), .ZN(n6564) );
  OAI211_X1 U8329 ( .C1(n6562), .C2(n6561), .A(n10050), .B(n6560), .ZN(n6563)
         );
  OAI211_X1 U8330 ( .C1(n8402), .C2(n6565), .A(n6564), .B(n6563), .ZN(n6566)
         );
  AOI21_X1 U8331 ( .B1(n10055), .B2(n6567), .A(n6566), .ZN(n6568) );
  INV_X1 U8332 ( .A(n6568), .ZN(P2_U3256) );
  INV_X1 U8333 ( .A(n6569), .ZN(n6570) );
  NOR2_X1 U8334 ( .A1(n6571), .A2(n6570), .ZN(n6575) );
  NAND2_X1 U8335 ( .A1(n6573), .A2(n6572), .ZN(n6574) );
  XNOR2_X1 U8336 ( .A(n6575), .B(n6574), .ZN(n6581) );
  AOI21_X1 U8337 ( .B1(n8943), .B2(n9068), .A(n6576), .ZN(n6579) );
  OAI22_X1 U8338 ( .A1(n9046), .A2(n4843), .B1(n6946), .B2(n9024), .ZN(n6577)
         );
  INV_X1 U8339 ( .A(n6577), .ZN(n6578) );
  OAI211_X1 U8340 ( .C1(n9045), .C2(n6945), .A(n6579), .B(n6578), .ZN(n6580)
         );
  AOI21_X1 U8341 ( .B1(n6581), .B2(n8982), .A(n6580), .ZN(n6582) );
  INV_X1 U8342 ( .A(n6582), .ZN(P1_U3237) );
  XOR2_X1 U8343 ( .A(n6587), .B(n6583), .Z(n10122) );
  OAI21_X1 U8344 ( .B1(n6585), .B2(n10116), .A(n6584), .ZN(n6586) );
  NAND3_X1 U8345 ( .A1(n6586), .A2(n10138), .A3(n6767), .ZN(n10123) );
  OAI21_X1 U8346 ( .B1(n5014), .B2(n5621), .A(n6760), .ZN(n6589) );
  AOI21_X1 U8347 ( .B1(n6589), .B2(n10061), .A(n6588), .ZN(n10124) );
  OAI21_X1 U8348 ( .B1(n5638), .B2(n10123), .A(n10124), .ZN(n6593) );
  AOI22_X1 U8349 ( .A1(n8646), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n6590), .B2(
        n10071), .ZN(n6591) );
  OAI21_X1 U8350 ( .B1(n10125), .B2(n8639), .A(n6591), .ZN(n6592) );
  AOI21_X1 U8351 ( .B1(n6593), .B2(n6401), .A(n6592), .ZN(n6594) );
  OAI21_X1 U8352 ( .B1(n10122), .B2(n8557), .A(n6594), .ZN(P2_U3291) );
  XOR2_X1 U8353 ( .A(n6601), .B(n6595), .Z(n10120) );
  INV_X1 U8354 ( .A(n6596), .ZN(n6597) );
  AOI22_X1 U8355 ( .A1(n8646), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n6597), .B2(
        n10071), .ZN(n6598) );
  OAI21_X1 U8356 ( .B1(n4383), .B2(n8639), .A(n6598), .ZN(n6608) );
  NAND2_X1 U8357 ( .A1(n6600), .A2(n6599), .ZN(n6603) );
  INV_X1 U8358 ( .A(n6601), .ZN(n6602) );
  XNOR2_X1 U8359 ( .A(n6603), .B(n6602), .ZN(n6606) );
  OAI22_X1 U8360 ( .A1(n6604), .A2(n8624), .B1(n6762), .B2(n8622), .ZN(n6605)
         );
  AOI21_X1 U8361 ( .B1(n6606), .B2(n10061), .A(n6605), .ZN(n10119) );
  NOR2_X1 U8362 ( .A1(n10119), .A2(n8646), .ZN(n6607) );
  AOI211_X1 U8363 ( .C1(n8644), .C2(n10117), .A(n6608), .B(n6607), .ZN(n6609)
         );
  OAI21_X1 U8364 ( .B1(n10120), .B2(n8557), .A(n6609), .ZN(P2_U3292) );
  AOI211_X1 U8365 ( .C1(n6612), .C2(n6611), .A(n6610), .B(n9744), .ZN(n6613)
         );
  INV_X1 U8366 ( .A(n6613), .ZN(n6620) );
  AOI21_X1 U8367 ( .B1(n6616), .B2(n6615), .A(n6614), .ZN(n6618) );
  INV_X1 U8368 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10229) );
  NAND2_X1 U8369 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(n4374), .ZN(n7022) );
  OAI21_X1 U8370 ( .B1(n8417), .B2(n10229), .A(n7022), .ZN(n6617) );
  AOI21_X1 U8371 ( .B1(n10050), .B2(n6618), .A(n6617), .ZN(n6619) );
  OAI211_X1 U8372 ( .C1(n8402), .C2(n6621), .A(n6620), .B(n6619), .ZN(P2_U3253) );
  NAND2_X1 U8373 ( .A1(n6623), .A2(n6622), .ZN(n6624) );
  OR2_X1 U8374 ( .A1(n6626), .A2(n6813), .ZN(n6631) );
  OAI22_X1 U8375 ( .A1(n6476), .A2(n9302), .B1(n6628), .B2(n6627), .ZN(n6629)
         );
  INV_X1 U8376 ( .A(n6629), .ZN(n6630) );
  AOI22_X1 U8377 ( .A1(n10020), .A2(n8925), .B1(n9065), .B2(n8924), .ZN(n6633)
         );
  NAND2_X1 U8378 ( .A1(n6811), .A2(n6812), .ZN(n6637) );
  NAND2_X1 U8379 ( .A1(n10020), .A2(n8918), .ZN(n6635) );
  NAND2_X1 U8380 ( .A1(n9065), .A2(n8919), .ZN(n6634) );
  NAND2_X1 U8381 ( .A1(n6635), .A2(n6634), .ZN(n6636) );
  XNOR2_X1 U8382 ( .A(n6636), .B(n8922), .ZN(n6810) );
  XNOR2_X1 U8383 ( .A(n6637), .B(n6810), .ZN(n6650) );
  NAND2_X1 U8384 ( .A1(n6350), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6645) );
  INV_X1 U8385 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6638) );
  OR2_X1 U8386 ( .A1(n7703), .A2(n6638), .ZN(n6644) );
  INV_X1 U8387 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6639) );
  NAND2_X1 U8388 ( .A1(n6640), .A2(n6639), .ZN(n6641) );
  NAND2_X1 U8389 ( .A1(n6823), .A2(n6641), .ZN(n6921) );
  OR2_X1 U8390 ( .A1(n6349), .A2(n6921), .ZN(n6643) );
  INV_X1 U8391 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6922) );
  OR2_X1 U8392 ( .A1(n7679), .A2(n6922), .ZN(n6642) );
  NAND4_X1 U8393 ( .A1(n6645), .A2(n6644), .A3(n6643), .A4(n6642), .ZN(n9064)
         );
  INV_X1 U8394 ( .A(n9064), .ZN(n7758) );
  OAI22_X1 U8395 ( .A1(n7758), .A2(n9046), .B1(n9045), .B2(n6957), .ZN(n6646)
         );
  AOI211_X1 U8396 ( .C1(n8943), .C2(n9066), .A(n6647), .B(n6646), .ZN(n6649)
         );
  NAND2_X1 U8397 ( .A1(n9050), .A2(n10020), .ZN(n6648) );
  OAI211_X1 U8398 ( .C1(n6650), .C2(n9052), .A(n6649), .B(n6648), .ZN(P1_U3219) );
  INV_X1 U8399 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9714) );
  OAI211_X1 U8400 ( .C1(n6653), .C2(n6652), .A(n10050), .B(n6651), .ZN(n6655)
         );
  NAND2_X1 U8401 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(n4374), .ZN(n6654) );
  OAI211_X1 U8402 ( .C1(n8417), .C2(n9714), .A(n6655), .B(n6654), .ZN(n6660)
         );
  AOI211_X1 U8403 ( .C1(n6658), .C2(n6657), .A(n6656), .B(n9744), .ZN(n6659)
         );
  AOI211_X1 U8404 ( .C1(n10053), .C2(n6661), .A(n6660), .B(n6659), .ZN(n6662)
         );
  INV_X1 U8405 ( .A(n6662), .ZN(P2_U3250) );
  INV_X1 U8406 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n6667) );
  OAI211_X1 U8407 ( .C1(n6665), .C2(n6664), .A(n10050), .B(n6663), .ZN(n6666)
         );
  NAND2_X1 U8408 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7128) );
  OAI211_X1 U8409 ( .C1(n8417), .C2(n6667), .A(n6666), .B(n7128), .ZN(n6672)
         );
  AOI211_X1 U8410 ( .C1(n6670), .C2(n6669), .A(n6668), .B(n9744), .ZN(n6671)
         );
  AOI211_X1 U8411 ( .C1(n10053), .C2(n6673), .A(n6672), .B(n6671), .ZN(n6674)
         );
  INV_X1 U8412 ( .A(n6674), .ZN(P2_U3255) );
  INV_X1 U8413 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10211) );
  AOI21_X1 U8414 ( .B1(n6677), .B2(n6676), .A(n6675), .ZN(n6678) );
  NAND2_X1 U8415 ( .A1(n10050), .A2(n6678), .ZN(n6679) );
  NAND2_X1 U8416 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n6714) );
  OAI211_X1 U8417 ( .C1(n8417), .C2(n10211), .A(n6679), .B(n6714), .ZN(n6684)
         );
  AOI211_X1 U8418 ( .C1(n6682), .C2(n6681), .A(n6680), .B(n9744), .ZN(n6683)
         );
  AOI211_X1 U8419 ( .C1(n10053), .C2(n6685), .A(n6684), .B(n6683), .ZN(n6686)
         );
  INV_X1 U8420 ( .A(n6686), .ZN(P2_U3251) );
  INV_X1 U8421 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9209) );
  OAI211_X1 U8422 ( .C1(n6689), .C2(n6688), .A(n10050), .B(n6687), .ZN(n6691)
         );
  OAI211_X1 U8423 ( .C1(n8417), .C2(n9209), .A(n6691), .B(n6690), .ZN(n6696)
         );
  AOI211_X1 U8424 ( .C1(n6694), .C2(n6693), .A(n6692), .B(n9744), .ZN(n6695)
         );
  AOI211_X1 U8425 ( .C1(n10053), .C2(n6697), .A(n6696), .B(n6695), .ZN(n6698)
         );
  INV_X1 U8426 ( .A(n6698), .ZN(P2_U3249) );
  INV_X1 U8427 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9722) );
  AOI21_X1 U8428 ( .B1(n6701), .B2(n6700), .A(n6699), .ZN(n6702) );
  NAND2_X1 U8429 ( .A1(n10050), .A2(n6702), .ZN(n6703) );
  NAND2_X1 U8430 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(n4374), .ZN(n7117) );
  OAI211_X1 U8431 ( .C1(n8417), .C2(n9722), .A(n6703), .B(n7117), .ZN(n6708)
         );
  AOI211_X1 U8432 ( .C1(n6706), .C2(n6705), .A(n6704), .B(n9744), .ZN(n6707)
         );
  AOI211_X1 U8433 ( .C1(n10053), .C2(n6709), .A(n6708), .B(n6707), .ZN(n6710)
         );
  INV_X1 U8434 ( .A(n6710), .ZN(P2_U3254) );
  OAI21_X1 U8435 ( .B1(n6713), .B2(n6712), .A(n6711), .ZN(n6718) );
  OAI22_X1 U8436 ( .A1(n4513), .A2(n8338), .B1(n8309), .B2(n7081), .ZN(n6717)
         );
  NAND2_X1 U8437 ( .A1(n6777), .A2(n8355), .ZN(n6715) );
  OAI211_X1 U8438 ( .C1(n8307), .C2(n6768), .A(n6715), .B(n6714), .ZN(n6716)
         );
  AOI211_X1 U8439 ( .C1(n6718), .C2(n8321), .A(n6717), .B(n6716), .ZN(n6719)
         );
  INV_X1 U8440 ( .A(n6719), .ZN(P2_U3241) );
  INV_X1 U8441 ( .A(n7593), .ZN(n8008) );
  OAI222_X1 U8442 ( .A1(n8761), .A2(n6720), .B1(n4385), .B2(n8008), .C1(n8218), 
        .C2(n4374), .ZN(P2_U3338) );
  INV_X1 U8443 ( .A(n8940), .ZN(n9970) );
  NAND2_X1 U8444 ( .A1(n6723), .A2(n8940), .ZN(n6724) );
  AND2_X1 U8445 ( .A1(n6799), .A2(n6724), .ZN(n6730) );
  INV_X2 U8446 ( .A(n9975), .ZN(n6725) );
  NAND2_X1 U8447 ( .A1(n6727), .A2(n9975), .ZN(n6728) );
  INV_X1 U8448 ( .A(n6729), .ZN(n6731) );
  NAND2_X1 U8449 ( .A1(n6731), .A2(n6730), .ZN(n6872) );
  OAI21_X1 U8450 ( .B1(n6730), .B2(n6731), .A(n6872), .ZN(n6746) );
  INV_X1 U8451 ( .A(n6746), .ZN(n9979) );
  INV_X1 U8452 ( .A(n6732), .ZN(n9690) );
  NAND4_X1 U8453 ( .A1(n6735), .A2(n9690), .A3(n6734), .A4(n6733), .ZN(n6749)
         );
  NAND2_X2 U8454 ( .A1(n6749), .A2(n9936), .ZN(n9926) );
  NOR2_X1 U8455 ( .A1(n6737), .A2(n9124), .ZN(n6736) );
  NAND2_X1 U8456 ( .A1(n9926), .A2(n6736), .ZN(n9905) );
  OR2_X1 U8457 ( .A1(n7992), .A2(n7967), .ZN(n6739) );
  NAND2_X1 U8458 ( .A1(n6737), .A2(n9124), .ZN(n6738) );
  MUX2_X1 U8459 ( .A(n6739), .B(n6738), .S(n7996), .Z(n9920) );
  INV_X1 U8460 ( .A(n9920), .ZN(n6747) );
  AND2_X1 U8461 ( .A1(n6723), .A2(n9970), .ZN(n7966) );
  XOR2_X1 U8462 ( .A(n6729), .B(n6851), .Z(n6744) );
  OR2_X1 U8463 ( .A1(n6177), .A2(n7967), .ZN(n6741) );
  NAND2_X1 U8464 ( .A1(n9203), .A2(n7996), .ZN(n6740) );
  NAND2_X1 U8465 ( .A1(n6741), .A2(n6740), .ZN(n9916) );
  INV_X1 U8466 ( .A(n9916), .ZN(n9588) );
  OR2_X1 U8467 ( .A1(n9800), .A2(n6742), .ZN(n9544) );
  INV_X1 U8468 ( .A(n9544), .ZN(n9913) );
  AOI22_X1 U8469 ( .A1(n9913), .A2(n6723), .B1(n6866), .B2(n9911), .ZN(n6743)
         );
  OAI21_X1 U8470 ( .B1(n6744), .B2(n9588), .A(n6743), .ZN(n6745) );
  AOI21_X1 U8471 ( .B1(n6747), .B2(n6746), .A(n6745), .ZN(n9978) );
  MUX2_X1 U8472 ( .A(n6748), .B(n9978), .S(n9926), .Z(n6756) );
  NOR2_X1 U8473 ( .A1(n6749), .A2(n9203), .ZN(n9573) );
  INV_X1 U8474 ( .A(n6751), .ZN(n6752) );
  AOI21_X1 U8475 ( .B1(n9975), .B2(n6752), .A(n9907), .ZN(n9976) );
  NAND2_X1 U8476 ( .A1(n9926), .A2(n9200), .ZN(n9930) );
  OAI22_X1 U8477 ( .A1(n9930), .A2(n6725), .B1(n6753), .B2(n9936), .ZN(n6754)
         );
  AOI21_X1 U8478 ( .B1(n9909), .B2(n9976), .A(n6754), .ZN(n6755) );
  OAI211_X1 U8479 ( .C1(n9979), .C2(n9905), .A(n6756), .B(n6755), .ZN(P1_U3289) );
  XNOR2_X1 U8480 ( .A(n6757), .B(n6759), .ZN(n10133) );
  NAND3_X1 U8481 ( .A1(n6760), .A2(n6759), .A3(n8033), .ZN(n6761) );
  NAND2_X1 U8482 ( .A1(n6758), .A2(n6761), .ZN(n6764) );
  OAI22_X1 U8483 ( .A1(n6762), .A2(n8624), .B1(n7081), .B2(n8622), .ZN(n6763)
         );
  AOI21_X1 U8484 ( .B1(n6764), .B2(n10061), .A(n6763), .ZN(n10131) );
  MUX2_X1 U8485 ( .A(n6765), .B(n10131), .S(n6401), .Z(n6771) );
  INV_X1 U8486 ( .A(n6845), .ZN(n6766) );
  AOI21_X1 U8487 ( .B1(n10128), .B2(n6767), .A(n6766), .ZN(n10129) );
  OAI22_X1 U8488 ( .A1(n8639), .A2(n4513), .B1(n8604), .B2(n6768), .ZN(n6769)
         );
  AOI21_X1 U8489 ( .B1(n10129), .B2(n8644), .A(n6769), .ZN(n6770) );
  OAI211_X1 U8490 ( .C1(n8557), .C2(n10133), .A(n6771), .B(n6770), .ZN(
        P2_U3290) );
  XNOR2_X1 U8491 ( .A(n6773), .B(n6772), .ZN(n6779) );
  OAI22_X1 U8492 ( .A1(n8307), .A2(n6846), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6774), .ZN(n6776) );
  OAI22_X1 U8493 ( .A1(n6847), .A2(n8338), .B1(n8309), .B2(n7118), .ZN(n6775)
         );
  AOI211_X1 U8494 ( .C1(n6777), .C2(n8354), .A(n6776), .B(n6775), .ZN(n6778)
         );
  OAI21_X1 U8495 ( .B1(n6779), .B2(n8316), .A(n6778), .ZN(P2_U3215) );
  INV_X1 U8496 ( .A(n6780), .ZN(n6784) );
  INV_X1 U8497 ( .A(n6781), .ZN(n6783) );
  OAI211_X1 U8498 ( .C1(n6784), .C2(n6783), .A(n10055), .B(n6782), .ZN(n6794)
         );
  INV_X1 U8499 ( .A(n6785), .ZN(n6788) );
  INV_X1 U8500 ( .A(n6786), .ZN(n6787) );
  NAND2_X1 U8501 ( .A1(n6788), .A2(n6787), .ZN(n6789) );
  NAND2_X1 U8502 ( .A1(n6790), .A2(n6789), .ZN(n6792) );
  INV_X1 U8503 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n9211) );
  NAND2_X1 U8504 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7261) );
  OAI21_X1 U8505 ( .B1(n8417), .B2(n9211), .A(n7261), .ZN(n6791) );
  AOI21_X1 U8506 ( .B1(n10050), .B2(n6792), .A(n6791), .ZN(n6793) );
  OAI211_X1 U8507 ( .C1(n8402), .C2(n6795), .A(n6794), .B(n6793), .ZN(P2_U3257) );
  INV_X1 U8508 ( .A(n7605), .ZN(n6834) );
  OAI222_X1 U8509 ( .A1(n9695), .A2(n6834), .B1(n9698), .B2(n6796), .C1(
        P1_U3084), .C2(n7967), .ZN(P1_U3332) );
  OAI21_X1 U8510 ( .B1(n6798), .B2(n6800), .A(n6799), .ZN(n9968) );
  AOI22_X1 U8511 ( .A1(n9913), .A2(n8942), .B1(n6727), .B2(n9911), .ZN(n6804)
         );
  XNOR2_X1 U8512 ( .A(n6798), .B(n6801), .ZN(n6802) );
  NAND2_X1 U8513 ( .A1(n6802), .A2(n9916), .ZN(n6803) );
  OAI211_X1 U8514 ( .C1(n9968), .C2(n9920), .A(n6804), .B(n6803), .ZN(n9971)
         );
  XNOR2_X1 U8515 ( .A(n8940), .B(n9929), .ZN(n6805) );
  NAND2_X1 U8516 ( .A1(n6805), .A2(n10005), .ZN(n9969) );
  INV_X1 U8517 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6806) );
  OAI22_X1 U8518 ( .A1(n9969), .A2(n9203), .B1(n9936), .B2(n6806), .ZN(n6807)
         );
  OAI21_X1 U8519 ( .B1(n9971), .B2(n6807), .A(n9926), .ZN(n6809) );
  INV_X1 U8520 ( .A(n9930), .ZN(n7408) );
  AOI22_X1 U8521 ( .A1(n7408), .A2(n8940), .B1(n4382), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6808) );
  OAI211_X1 U8522 ( .C1(n9968), .C2(n9905), .A(n6809), .B(n6808), .ZN(P1_U3290) );
  NAND2_X1 U8523 ( .A1(n6814), .A2(n7747), .ZN(n6816) );
  AOI22_X1 U8524 ( .A1(n7748), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9899), .B2(
        n7279), .ZN(n6815) );
  NAND2_X1 U8525 ( .A1(n7759), .A2(n8918), .ZN(n6818) );
  NAND2_X1 U8526 ( .A1(n9064), .A2(n8925), .ZN(n6817) );
  NAND2_X1 U8527 ( .A1(n6818), .A2(n6817), .ZN(n6819) );
  XNOR2_X1 U8528 ( .A(n6819), .B(n6247), .ZN(n6981) );
  AND2_X1 U8529 ( .A1(n9064), .A2(n8924), .ZN(n6820) );
  AOI21_X1 U8530 ( .B1(n7759), .B2(n8925), .A(n6820), .ZN(n6982) );
  XNOR2_X1 U8531 ( .A(n6981), .B(n6982), .ZN(n6979) );
  XOR2_X1 U8532 ( .A(n6980), .B(n6979), .Z(n6833) );
  NOR2_X1 U8533 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6639), .ZN(n9892) );
  NAND2_X1 U8534 ( .A1(n6350), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6829) );
  OR2_X1 U8535 ( .A1(n7703), .A2(n6821), .ZN(n6828) );
  INV_X1 U8536 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6822) );
  NAND2_X1 U8537 ( .A1(n6823), .A2(n6822), .ZN(n6824) );
  NAND2_X1 U8538 ( .A1(n6997), .A2(n6824), .ZN(n7143) );
  OR2_X1 U8539 ( .A1(n6349), .A2(n7143), .ZN(n6827) );
  INV_X1 U8540 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6825) );
  OR2_X1 U8541 ( .A1(n7679), .A2(n6825), .ZN(n6826) );
  NAND4_X1 U8542 ( .A1(n6829), .A2(n6828), .A3(n6827), .A4(n6826), .ZN(n9063)
         );
  OAI22_X1 U8543 ( .A1(n7046), .A2(n9046), .B1(n9045), .B2(n6921), .ZN(n6830)
         );
  AOI211_X1 U8544 ( .C1(n8943), .C2(n9065), .A(n9892), .B(n6830), .ZN(n6832)
         );
  NAND2_X1 U8545 ( .A1(n7759), .A2(n9050), .ZN(n6831) );
  OAI211_X1 U8546 ( .C1(n6833), .C2(n9052), .A(n6832), .B(n6831), .ZN(P1_U3229) );
  OAI222_X1 U8547 ( .A1(n8761), .A2(n9322), .B1(n4385), .B2(n6834), .C1(n8024), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  OAI21_X1 U8548 ( .B1(n6835), .B2(n8060), .A(n6836), .ZN(n6837) );
  INV_X1 U8549 ( .A(n6837), .ZN(n7012) );
  NAND2_X1 U8550 ( .A1(n6758), .A2(n8059), .ZN(n6838) );
  NAND2_X1 U8551 ( .A1(n6838), .A2(n8060), .ZN(n6840) );
  NAND3_X1 U8552 ( .A1(n6840), .A2(n10061), .A3(n6839), .ZN(n6844) );
  OAI22_X1 U8553 ( .A1(n6841), .A2(n8624), .B1(n7118), .B2(n8622), .ZN(n6842)
         );
  INV_X1 U8554 ( .A(n6842), .ZN(n6843) );
  AND2_X1 U8555 ( .A1(n6844), .A2(n6843), .ZN(n7011) );
  MUX2_X1 U8556 ( .A(n7011), .B(n9464), .S(n8646), .Z(n6850) );
  AOI21_X1 U8557 ( .B1(n7008), .B2(n6845), .A(n7091), .ZN(n7009) );
  OAI22_X1 U8558 ( .A1(n8639), .A2(n6847), .B1(n8604), .B2(n6846), .ZN(n6848)
         );
  AOI21_X1 U8559 ( .B1(n7009), .B2(n8644), .A(n6848), .ZN(n6849) );
  OAI211_X1 U8560 ( .C1(n7012), .C2(n8557), .A(n6850), .B(n6849), .ZN(P2_U3289) );
  OR2_X1 U8561 ( .A1(n9068), .A2(n9999), .ZN(n6938) );
  NAND2_X1 U8562 ( .A1(n9068), .A2(n9999), .ZN(n6935) );
  INV_X1 U8563 ( .A(n6878), .ZN(n6875) );
  OR2_X1 U8564 ( .A1(n6727), .A2(n6725), .ZN(n6852) );
  NAND2_X1 U8565 ( .A1(n6866), .A2(n9982), .ZN(n6893) );
  INV_X1 U8566 ( .A(n6894), .ZN(n6854) );
  NAND2_X1 U8567 ( .A1(n9912), .A2(n9989), .ZN(n6892) );
  XOR2_X1 U8568 ( .A(n6875), .B(n6937), .Z(n6856) );
  AOI222_X1 U8569 ( .A1(n9916), .A2(n6856), .B1(n9067), .B2(n9911), .C1(n9912), 
        .C2(n9913), .ZN(n9998) );
  NAND2_X1 U8570 ( .A1(n9907), .A2(n9982), .ZN(n9906) );
  INV_X1 U8571 ( .A(n10005), .ZN(n10029) );
  AOI21_X1 U8572 ( .B1(n6912), .B2(n6883), .A(n10029), .ZN(n6857) );
  NAND2_X1 U8573 ( .A1(n6857), .A2(n6944), .ZN(n9997) );
  INV_X1 U8574 ( .A(n9573), .ZN(n6863) );
  INV_X1 U8575 ( .A(n6858), .ZN(n6859) );
  OAI22_X1 U8576 ( .A1(n9926), .A2(n6860), .B1(n6859), .B2(n9936), .ZN(n6861)
         );
  AOI21_X1 U8577 ( .B1(n7408), .B2(n6883), .A(n6861), .ZN(n6862) );
  OAI21_X1 U8578 ( .B1(n9997), .B2(n6863), .A(n6862), .ZN(n6864) );
  INV_X1 U8579 ( .A(n6864), .ZN(n6882) );
  OR2_X1 U8580 ( .A1(n6866), .A2(n6865), .ZN(n6867) );
  AND2_X1 U8581 ( .A1(n9903), .A2(n6867), .ZN(n6871) );
  INV_X1 U8582 ( .A(n6867), .ZN(n6869) );
  NOR2_X1 U8583 ( .A1(n6869), .A2(n9915), .ZN(n6870) );
  NAND2_X1 U8584 ( .A1(n6903), .A2(n6905), .ZN(n6874) );
  OR2_X1 U8585 ( .A1(n9912), .A2(n6915), .ZN(n6873) );
  NAND2_X1 U8586 ( .A1(n6874), .A2(n6873), .ZN(n6877) );
  AND2_X1 U8587 ( .A1(n6877), .A2(n6875), .ZN(n9996) );
  INV_X1 U8588 ( .A(n9996), .ZN(n6880) );
  NOR2_X1 U8589 ( .A1(n6876), .A2(n8922), .ZN(n9205) );
  NAND2_X1 U8590 ( .A1(n9926), .A2(n9205), .ZN(n9597) );
  INV_X1 U8591 ( .A(n9597), .ZN(n7330) );
  INV_X1 U8592 ( .A(n6877), .ZN(n6879) );
  NAND3_X1 U8593 ( .A1(n6880), .A2(n7330), .A3(n10001), .ZN(n6881) );
  OAI211_X1 U8594 ( .C1(n9998), .C2(n4382), .A(n6882), .B(n6881), .ZN(P1_U3286) );
  NAND2_X1 U8595 ( .A1(n9068), .A2(n6883), .ZN(n6884) );
  NAND2_X1 U8596 ( .A1(n10001), .A2(n6884), .ZN(n6934) );
  NAND2_X1 U8597 ( .A1(n9067), .A2(n6946), .ZN(n7755) );
  OR2_X1 U8598 ( .A1(n9067), .A2(n10003), .ZN(n6886) );
  NAND2_X1 U8599 ( .A1(n10015), .A2(n9066), .ZN(n7905) );
  XNOR2_X1 U8600 ( .A(n6927), .B(n7856), .ZN(n10017) );
  NAND2_X1 U8601 ( .A1(n6943), .A2(n10015), .ZN(n6959) );
  OAI211_X1 U8602 ( .C1(n6943), .C2(n10015), .A(n10005), .B(n6959), .ZN(n10013) );
  OAI22_X1 U8603 ( .A1(n9926), .A2(n6888), .B1(n6887), .B2(n9936), .ZN(n6889)
         );
  AOI21_X1 U8604 ( .B1(n7408), .B2(n6926), .A(n6889), .ZN(n6890) );
  OAI21_X1 U8605 ( .B1(n10013), .B2(n6863), .A(n6890), .ZN(n6901) );
  INV_X1 U8606 ( .A(n6891), .ZN(n9914) );
  AND3_X1 U8607 ( .A1(n6896), .A2(n7755), .A3(n6893), .ZN(n7854) );
  NAND2_X1 U8608 ( .A1(n6894), .A2(n6868), .ZN(n6895) );
  NAND2_X1 U8609 ( .A1(n6896), .A2(n6895), .ZN(n6897) );
  NAND3_X1 U8610 ( .A1(n6897), .A2(n7762), .A3(n6938), .ZN(n7858) );
  INV_X1 U8611 ( .A(n7856), .ZN(n6898) );
  OAI21_X1 U8612 ( .B1(n7974), .B2(n6898), .A(n6918), .ZN(n6899) );
  AOI222_X1 U8613 ( .A1(n9916), .A2(n6899), .B1(n9065), .B2(n9911), .C1(n9067), 
        .C2(n9913), .ZN(n10014) );
  NOR2_X1 U8614 ( .A1(n10014), .A2(n4382), .ZN(n6900) );
  AOI211_X1 U8615 ( .C1(n7330), .C2(n10017), .A(n6901), .B(n6900), .ZN(n6902)
         );
  INV_X1 U8616 ( .A(n6902), .ZN(P1_U3284) );
  XOR2_X1 U8617 ( .A(n6905), .B(n6903), .Z(n9988) );
  AOI22_X1 U8618 ( .A1(n9913), .A2(n6866), .B1(n9068), .B2(n9911), .ZN(n6908)
         );
  XOR2_X1 U8619 ( .A(n6905), .B(n6904), .Z(n6906) );
  NAND2_X1 U8620 ( .A1(n6906), .A2(n9916), .ZN(n6907) );
  OAI211_X1 U8621 ( .C1(n9988), .C2(n9920), .A(n6908), .B(n6907), .ZN(n9991)
         );
  NAND2_X1 U8622 ( .A1(n9991), .A2(n9926), .ZN(n6917) );
  OAI22_X1 U8623 ( .A1(n9926), .A2(n6910), .B1(n6909), .B2(n9936), .ZN(n6914)
         );
  INV_X1 U8624 ( .A(n9909), .ZN(n9931) );
  NAND2_X1 U8625 ( .A1(n9906), .A2(n6915), .ZN(n6911) );
  NAND2_X1 U8626 ( .A1(n6912), .A2(n6911), .ZN(n9990) );
  NOR2_X1 U8627 ( .A1(n9931), .A2(n9990), .ZN(n6913) );
  AOI211_X1 U8628 ( .C1(n7408), .C2(n6915), .A(n6914), .B(n6913), .ZN(n6916)
         );
  OAI211_X1 U8629 ( .C1(n9988), .C2(n9905), .A(n6917), .B(n6916), .ZN(P1_U3287) );
  INV_X1 U8630 ( .A(n9911), .ZN(n9546) );
  NAND2_X1 U8631 ( .A1(n6919), .A2(n10020), .ZN(n7768) );
  NAND2_X1 U8632 ( .A1(n7765), .A2(n7768), .ZN(n7857) );
  OAI21_X1 U8633 ( .B1(n6953), .B2(n7857), .A(n7765), .ZN(n7044) );
  XNOR2_X1 U8634 ( .A(n7759), .B(n9064), .ZN(n7860) );
  XNOR2_X1 U8635 ( .A(n7044), .B(n7860), .ZN(n6920) );
  OAI222_X1 U8636 ( .A1(n9546), .A2(n7046), .B1(n6920), .B2(n9588), .C1(n9544), 
        .C2(n6919), .ZN(n10031) );
  INV_X1 U8637 ( .A(n10031), .ZN(n6931) );
  OAI22_X1 U8638 ( .A1(n9926), .A2(n6922), .B1(n6921), .B2(n9936), .ZN(n6925)
         );
  INV_X1 U8639 ( .A(n7759), .ZN(n10028) );
  INV_X1 U8640 ( .A(n6961), .ZN(n6923) );
  INV_X1 U8641 ( .A(n7047), .ZN(n7142) );
  OAI21_X1 U8642 ( .B1(n10028), .B2(n6923), .A(n7142), .ZN(n10030) );
  NOR2_X1 U8643 ( .A1(n10030), .A2(n9931), .ZN(n6924) );
  AOI211_X1 U8644 ( .C1(n7408), .C2(n7759), .A(n6925), .B(n6924), .ZN(n6930)
         );
  NAND2_X1 U8645 ( .A1(n6950), .A2(n7857), .ZN(n6952) );
  NAND2_X1 U8646 ( .A1(n10020), .A2(n9065), .ZN(n6928) );
  NAND2_X1 U8647 ( .A1(n6952), .A2(n6928), .ZN(n7028) );
  XNOR2_X1 U8648 ( .A(n7028), .B(n7860), .ZN(n10033) );
  NAND2_X1 U8649 ( .A1(n10033), .A2(n7330), .ZN(n6929) );
  OAI211_X1 U8650 ( .C1(n6931), .C2(n4382), .A(n6930), .B(n6929), .ZN(P1_U3282) );
  INV_X1 U8651 ( .A(n6932), .ZN(n6933) );
  AOI21_X1 U8652 ( .B1(n7753), .B2(n6934), .A(n6933), .ZN(n10010) );
  INV_X1 U8653 ( .A(n6935), .ZN(n6936) );
  XOR2_X1 U8654 ( .A(n7753), .B(n7752), .Z(n6942) );
  INV_X1 U8655 ( .A(n9068), .ZN(n6939) );
  OAI22_X1 U8656 ( .A1(n6939), .A2(n9544), .B1(n4843), .B2(n9546), .ZN(n6941)
         );
  NOR2_X1 U8657 ( .A1(n10010), .A2(n9920), .ZN(n6940) );
  AOI211_X1 U8658 ( .C1(n6942), .C2(n9916), .A(n6941), .B(n6940), .ZN(n10008)
         );
  MUX2_X1 U8659 ( .A(n5877), .B(n10008), .S(n9926), .Z(n6949) );
  AOI21_X1 U8660 ( .B1(n10003), .B2(n6944), .A(n6943), .ZN(n10006) );
  OAI22_X1 U8661 ( .A1(n9930), .A2(n6946), .B1(n9936), .B2(n6945), .ZN(n6947)
         );
  AOI21_X1 U8662 ( .B1(n10006), .B2(n9909), .A(n6947), .ZN(n6948) );
  OAI211_X1 U8663 ( .C1(n10010), .C2(n9905), .A(n6949), .B(n6948), .ZN(
        P1_U3285) );
  OR2_X1 U8664 ( .A1(n6950), .A2(n7857), .ZN(n6951) );
  NAND2_X1 U8665 ( .A1(n6952), .A2(n6951), .ZN(n10019) );
  AOI22_X1 U8666 ( .A1(n9913), .A2(n9066), .B1(n9064), .B2(n9911), .ZN(n6956)
         );
  XOR2_X1 U8667 ( .A(n7857), .B(n6953), .Z(n6954) );
  NAND2_X1 U8668 ( .A1(n6954), .A2(n9916), .ZN(n6955) );
  OAI211_X1 U8669 ( .C1(n10019), .C2(n9920), .A(n6956), .B(n6955), .ZN(n10022)
         );
  NAND2_X1 U8670 ( .A1(n10022), .A2(n9926), .ZN(n6965) );
  OAI22_X1 U8671 ( .A1(n9926), .A2(n6958), .B1(n6957), .B2(n9936), .ZN(n6963)
         );
  NAND2_X1 U8672 ( .A1(n6959), .A2(n10020), .ZN(n6960) );
  NAND2_X1 U8673 ( .A1(n6961), .A2(n6960), .ZN(n10021) );
  NOR2_X1 U8674 ( .A1(n10021), .A2(n9931), .ZN(n6962) );
  AOI211_X1 U8675 ( .C1(n7408), .C2(n10020), .A(n6963), .B(n6962), .ZN(n6964)
         );
  OAI211_X1 U8676 ( .C1(n10019), .C2(n9905), .A(n6965), .B(n6964), .ZN(
        P1_U3283) );
  INV_X1 U8677 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n6978) );
  OAI21_X1 U8678 ( .B1(n6968), .B2(n6967), .A(n6966), .ZN(n6976) );
  INV_X1 U8679 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9388) );
  NOR2_X1 U8680 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9388), .ZN(n8895) );
  INV_X1 U8681 ( .A(n8895), .ZN(n6969) );
  OAI21_X1 U8682 ( .B1(n9818), .B2(n6970), .A(n6969), .ZN(n6975) );
  AOI211_X1 U8683 ( .C1(n6973), .C2(n6972), .A(n6971), .B(n9827), .ZN(n6974)
         );
  AOI211_X1 U8684 ( .C1(n9872), .C2(n6976), .A(n6975), .B(n6974), .ZN(n6977)
         );
  OAI21_X1 U8685 ( .B1(n9880), .B2(n6978), .A(n6977), .ZN(P1_U3255) );
  INV_X1 U8686 ( .A(n6981), .ZN(n6983) );
  NAND2_X1 U8687 ( .A1(n6983), .A2(n6982), .ZN(n6984) );
  NAND2_X1 U8688 ( .A1(n6985), .A2(n6984), .ZN(n7054) );
  NAND2_X1 U8689 ( .A1(n6986), .A2(n7747), .ZN(n6989) );
  AOI22_X1 U8690 ( .A1(n7748), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6987), .B2(
        n7279), .ZN(n6988) );
  NAND2_X1 U8691 ( .A1(n7270), .A2(n8918), .ZN(n6991) );
  NAND2_X1 U8692 ( .A1(n9063), .A2(n8919), .ZN(n6990) );
  NAND2_X1 U8693 ( .A1(n6991), .A2(n6990), .ZN(n6992) );
  XNOR2_X1 U8694 ( .A(n6992), .B(n6247), .ZN(n7055) );
  AND2_X1 U8695 ( .A1(n9063), .A2(n8924), .ZN(n6993) );
  AOI21_X1 U8696 ( .B1(n7270), .B2(n8925), .A(n6993), .ZN(n7056) );
  XNOR2_X1 U8697 ( .A(n7055), .B(n7056), .ZN(n7053) );
  XOR2_X1 U8698 ( .A(n7054), .B(n7053), .Z(n7007) );
  OAI21_X1 U8699 ( .B1(n9043), .B2(n7758), .A(n6994), .ZN(n7005) );
  NAND2_X1 U8700 ( .A1(n6350), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7003) );
  OR2_X1 U8701 ( .A1(n7703), .A2(n6995), .ZN(n7002) );
  INV_X1 U8702 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6996) );
  AND2_X1 U8703 ( .A1(n6997), .A2(n6996), .ZN(n6998) );
  OR2_X1 U8704 ( .A1(n6998), .A2(n7037), .ZN(n7069) );
  OR2_X1 U8705 ( .A1(n6349), .A2(n7069), .ZN(n7001) );
  OR2_X1 U8706 ( .A1(n7679), .A2(n6999), .ZN(n7000) );
  NAND4_X1 U8707 ( .A1(n7003), .A2(n7002), .A3(n7001), .A4(n7000), .ZN(n9062)
         );
  OAI22_X1 U8708 ( .A1(n7776), .A2(n9046), .B1(n9045), .B2(n7143), .ZN(n7004)
         );
  AOI211_X1 U8709 ( .C1(n7270), .C2(n9050), .A(n7005), .B(n7004), .ZN(n7006)
         );
  OAI21_X1 U8710 ( .B1(n7007), .B2(n9052), .A(n7006), .ZN(P1_U3215) );
  INV_X1 U8711 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7014) );
  AOI22_X1 U8712 ( .A1(n7009), .A2(n10138), .B1(n10137), .B2(n7008), .ZN(n7010) );
  OAI211_X1 U8713 ( .C1(n7012), .C2(n10132), .A(n7011), .B(n7010), .ZN(n7015)
         );
  NAND2_X1 U8714 ( .A1(n7015), .A2(n10163), .ZN(n7013) );
  OAI21_X1 U8715 ( .B1(n10163), .B2(n7014), .A(n7013), .ZN(P2_U3472) );
  NAND2_X1 U8716 ( .A1(n7015), .A2(n10177), .ZN(n7016) );
  OAI21_X1 U8717 ( .B1(n10177), .B2(n5282), .A(n7016), .ZN(P2_U3527) );
  INV_X1 U8718 ( .A(n7619), .ZN(n7019) );
  OAI222_X1 U8719 ( .A1(n9698), .A2(n7017), .B1(n9695), .B2(n7019), .C1(
        P1_U3084), .C2(n7844), .ZN(P1_U3331) );
  OAI222_X1 U8720 ( .A1(n8761), .A2(n9358), .B1(n4385), .B2(n7019), .C1(
        P2_U3152), .C2(n7018), .ZN(P2_U3336) );
  XNOR2_X1 U8721 ( .A(n7021), .B(n7020), .ZN(n7026) );
  OAI21_X1 U8722 ( .B1(n8307), .B2(n7093), .A(n7022), .ZN(n7024) );
  OAI22_X1 U8723 ( .A1(n7081), .A2(n8310), .B1(n8309), .B2(n7243), .ZN(n7023)
         );
  AOI211_X1 U8724 ( .C1(n10136), .C2(n8314), .A(n7024), .B(n7023), .ZN(n7025)
         );
  OAI21_X1 U8725 ( .B1(n7026), .B2(n8316), .A(n7025), .ZN(P2_U3223) );
  OR2_X1 U8726 ( .A1(n7759), .A2(n9064), .ZN(n7027) );
  NAND2_X1 U8727 ( .A1(n7759), .A2(n9064), .ZN(n7029) );
  NAND2_X1 U8728 ( .A1(n7270), .A2(n7046), .ZN(n7887) );
  OR2_X1 U8729 ( .A1(n7270), .A2(n9063), .ZN(n7032) );
  NAND2_X1 U8730 ( .A1(n7033), .A2(n7747), .ZN(n7036) );
  AOI22_X1 U8731 ( .A1(n7748), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7034), .B2(
        n7279), .ZN(n7035) );
  XNOR2_X1 U8732 ( .A(n7777), .B(n7776), .ZN(n7866) );
  XNOR2_X1 U8733 ( .A(n7189), .B(n7866), .ZN(n9789) );
  INV_X1 U8734 ( .A(n9789), .ZN(n7052) );
  INV_X1 U8735 ( .A(n7679), .ZN(n7635) );
  NAND2_X1 U8736 ( .A1(n7635), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7043) );
  OR2_X1 U8737 ( .A1(n7703), .A2(n9784), .ZN(n7042) );
  NAND2_X1 U8738 ( .A1(n7037), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7296) );
  OR2_X1 U8739 ( .A1(n7037), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7038) );
  NAND2_X1 U8740 ( .A1(n7296), .A2(n7038), .ZN(n7197) );
  OR2_X1 U8741 ( .A1(n6349), .A2(n7197), .ZN(n7041) );
  INV_X1 U8742 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7039) );
  OR2_X1 U8743 ( .A1(n7719), .A2(n7039), .ZN(n7040) );
  NAND4_X1 U8744 ( .A1(n7043), .A2(n7042), .A3(n7041), .A4(n7040), .ZN(n9061)
         );
  INV_X1 U8745 ( .A(n9061), .ZN(n7397) );
  NOR2_X1 U8746 ( .A1(n7759), .A2(n7758), .ZN(n7770) );
  XNOR2_X1 U8747 ( .A(n7193), .B(n7866), .ZN(n7045) );
  OAI222_X1 U8748 ( .A1(n9546), .A2(n7397), .B1(n9544), .B2(n7046), .C1(n9588), 
        .C2(n7045), .ZN(n9787) );
  INV_X1 U8749 ( .A(n7270), .ZN(n7146) );
  AND2_X2 U8750 ( .A1(n7047), .A2(n7146), .ZN(n7141) );
  NAND2_X1 U8751 ( .A1(n7141), .A2(n9785), .ZN(n7199) );
  OAI21_X1 U8752 ( .B1(n7141), .B2(n9785), .A(n7199), .ZN(n9786) );
  OAI22_X1 U8753 ( .A1(n9926), .A2(n6999), .B1(n7069), .B2(n9936), .ZN(n7048)
         );
  AOI21_X1 U8754 ( .B1(n7777), .B2(n7408), .A(n7048), .ZN(n7049) );
  OAI21_X1 U8755 ( .B1(n9786), .B2(n9931), .A(n7049), .ZN(n7050) );
  AOI21_X1 U8756 ( .B1(n9787), .B2(n9926), .A(n7050), .ZN(n7051) );
  OAI21_X1 U8757 ( .B1(n9597), .B2(n7052), .A(n7051), .ZN(P1_U3280) );
  NAND2_X1 U8758 ( .A1(n7054), .A2(n7053), .ZN(n7059) );
  INV_X1 U8759 ( .A(n7055), .ZN(n7057) );
  NAND2_X1 U8760 ( .A1(n7057), .A2(n7056), .ZN(n7058) );
  NAND2_X1 U8761 ( .A1(n7777), .A2(n8918), .ZN(n7061) );
  NAND2_X1 U8762 ( .A1(n9062), .A2(n8925), .ZN(n7060) );
  NAND2_X1 U8763 ( .A1(n7061), .A2(n7060), .ZN(n7062) );
  XNOR2_X1 U8764 ( .A(n7062), .B(n8922), .ZN(n7169) );
  AND2_X1 U8765 ( .A1(n9062), .A2(n8924), .ZN(n7063) );
  AOI21_X1 U8766 ( .B1(n7777), .B2(n8919), .A(n7063), .ZN(n7170) );
  XNOR2_X1 U8767 ( .A(n7169), .B(n7170), .ZN(n7065) );
  AOI21_X1 U8768 ( .B1(n7064), .B2(n7065), .A(n9052), .ZN(n7067) );
  NAND2_X1 U8769 ( .A1(n7067), .A2(n7174), .ZN(n7073) );
  INV_X1 U8770 ( .A(n7068), .ZN(n7071) );
  OAI22_X1 U8771 ( .A1(n7397), .A2(n9046), .B1(n9045), .B2(n7069), .ZN(n7070)
         );
  AOI211_X1 U8772 ( .C1(n8943), .C2(n9063), .A(n7071), .B(n7070), .ZN(n7072)
         );
  OAI211_X1 U8773 ( .C1(n9785), .C2(n9024), .A(n7073), .B(n7072), .ZN(P1_U3234) );
  INV_X1 U8774 ( .A(n7629), .ZN(n7076) );
  NOR2_X1 U8775 ( .A1(n7074), .A2(P1_U3084), .ZN(n7991) );
  AOI21_X1 U8776 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9699), .A(n7991), .ZN(
        n7075) );
  OAI21_X1 U8777 ( .B1(n7076), .B2(n8009), .A(n7075), .ZN(P1_U3330) );
  NAND2_X1 U8778 ( .A1(n7629), .A2(n7077), .ZN(n7078) );
  OAI211_X1 U8779 ( .C1(n7079), .C2(n8761), .A(n7078), .B(n8230), .ZN(P2_U3335) );
  XNOR2_X1 U8780 ( .A(n7080), .B(n8192), .ZN(n7089) );
  INV_X1 U8781 ( .A(n7089), .ZN(n10143) );
  INV_X1 U8782 ( .A(n8630), .ZN(n7088) );
  OAI22_X1 U8783 ( .A1(n7081), .A2(n8624), .B1(n7243), .B2(n8622), .ZN(n7087)
         );
  INV_X1 U8784 ( .A(n6839), .ZN(n7083) );
  OAI21_X1 U8785 ( .B1(n7083), .B2(n7082), .A(n8192), .ZN(n7085) );
  AOI21_X1 U8786 ( .B1(n7085), .B2(n7084), .A(n8612), .ZN(n7086) );
  AOI211_X1 U8787 ( .C1(n7089), .C2(n7088), .A(n7087), .B(n7086), .ZN(n10141)
         );
  MUX2_X1 U8788 ( .A(n7090), .B(n10141), .S(n6401), .Z(n7097) );
  INV_X1 U8789 ( .A(n7091), .ZN(n7092) );
  AOI21_X1 U8790 ( .B1(n10136), .B2(n7092), .A(n7153), .ZN(n10139) );
  OAI22_X1 U8791 ( .A1(n8639), .A2(n7094), .B1(n8604), .B2(n7093), .ZN(n7095)
         );
  AOI21_X1 U8792 ( .B1(n10139), .B2(n8644), .A(n7095), .ZN(n7096) );
  OAI211_X1 U8793 ( .C1(n10143), .C2(n8641), .A(n7097), .B(n7096), .ZN(
        P2_U3288) );
  INV_X1 U8794 ( .A(n7098), .ZN(n7111) );
  OAI21_X1 U8795 ( .B1(n7101), .B2(n7100), .A(n7099), .ZN(n7102) );
  NAND2_X1 U8796 ( .A1(n10055), .A2(n7102), .ZN(n7110) );
  OAI21_X1 U8797 ( .B1(n7105), .B2(n7104), .A(n7103), .ZN(n7108) );
  INV_X1 U8798 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7106) );
  NAND2_X1 U8799 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(n4374), .ZN(n7221) );
  OAI21_X1 U8800 ( .B1(n8417), .B2(n7106), .A(n7221), .ZN(n7107) );
  AOI21_X1 U8801 ( .B1(n10050), .B2(n7108), .A(n7107), .ZN(n7109) );
  OAI211_X1 U8802 ( .C1(n8402), .C2(n7111), .A(n7110), .B(n7109), .ZN(P2_U3258) );
  OAI21_X1 U8803 ( .B1(n7114), .B2(n7113), .A(n7112), .ZN(n7115) );
  NAND2_X1 U8804 ( .A1(n7115), .A2(n8321), .ZN(n7122) );
  INV_X1 U8805 ( .A(n7116), .ZN(n7205) );
  INV_X1 U8806 ( .A(n7117), .ZN(n7120) );
  OAI22_X1 U8807 ( .A1(n7118), .A2(n8310), .B1(n8309), .B2(n7232), .ZN(n7119)
         );
  AOI211_X1 U8808 ( .C1(n7205), .C2(n8336), .A(n7120), .B(n7119), .ZN(n7121)
         );
  OAI211_X1 U8809 ( .C1(n7207), .C2(n8338), .A(n7122), .B(n7121), .ZN(P2_U3233) );
  INV_X1 U8810 ( .A(n7642), .ZN(n7126) );
  INV_X1 U8811 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7123) );
  OAI222_X1 U8812 ( .A1(n8009), .A2(n7126), .B1(P1_U3084), .B2(n7124), .C1(
        n7123), .C2(n9698), .ZN(P1_U3329) );
  OAI222_X1 U8813 ( .A1(n4374), .A2(n7127), .B1(n4385), .B2(n7126), .C1(n7125), 
        .C2(n8761), .ZN(P2_U3334) );
  XNOR2_X1 U8814 ( .A(n7356), .B(n7226), .ZN(n7132) );
  OAI21_X1 U8815 ( .B1(n8307), .B2(n7247), .A(n7128), .ZN(n7130) );
  OAI22_X1 U8816 ( .A1(n7243), .A2(n8310), .B1(n8309), .B2(n7344), .ZN(n7129)
         );
  AOI211_X1 U8817 ( .C1(n7251), .C2(n8314), .A(n7130), .B(n7129), .ZN(n7131)
         );
  OAI21_X1 U8818 ( .B1(n7132), .B2(n8316), .A(n7131), .ZN(P2_U3219) );
  OAI21_X1 U8819 ( .B1(n7862), .B2(n7134), .A(n7133), .ZN(n7140) );
  OAI22_X1 U8820 ( .A1(n7776), .A2(n9546), .B1(n7758), .B2(n9544), .ZN(n7139)
         );
  INV_X1 U8821 ( .A(n7135), .ZN(n7136) );
  AOI21_X1 U8822 ( .B1(n7862), .B2(n7137), .A(n7136), .ZN(n7273) );
  NOR2_X1 U8823 ( .A1(n7273), .A2(n9920), .ZN(n7138) );
  AOI211_X1 U8824 ( .C1(n9916), .C2(n7140), .A(n7139), .B(n7138), .ZN(n7272)
         );
  AOI211_X1 U8825 ( .C1(n7270), .C2(n7142), .A(n10029), .B(n7141), .ZN(n7269)
         );
  INV_X1 U8826 ( .A(n7143), .ZN(n7144) );
  INV_X1 U8827 ( .A(n9936), .ZN(n9923) );
  AOI22_X1 U8828 ( .A1(n4382), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7144), .B2(
        n9923), .ZN(n7145) );
  OAI21_X1 U8829 ( .B1(n7146), .B2(n9930), .A(n7145), .ZN(n7148) );
  NOR2_X1 U8830 ( .A1(n7273), .A2(n9905), .ZN(n7147) );
  AOI211_X1 U8831 ( .C1(n7269), .C2(n9573), .A(n7148), .B(n7147), .ZN(n7149)
         );
  OAI21_X1 U8832 ( .B1(n7272), .B2(n4382), .A(n7149), .ZN(P1_U3281) );
  INV_X1 U8833 ( .A(n7151), .ZN(n8193) );
  XNOR2_X1 U8834 ( .A(n7150), .B(n8193), .ZN(n7213) );
  NAND2_X1 U8835 ( .A1(n7084), .A2(n8063), .ZN(n7377) );
  NAND2_X1 U8836 ( .A1(n7377), .A2(n7151), .ZN(n7240) );
  OAI21_X1 U8837 ( .B1(n7151), .B2(n7377), .A(n7240), .ZN(n7152) );
  AOI222_X1 U8838 ( .A1(n10061), .A2(n7152), .B1(n8350), .B2(n10065), .C1(
        n8352), .C2(n10066), .ZN(n7208) );
  INV_X1 U8839 ( .A(n7153), .ZN(n7154) );
  AOI21_X1 U8840 ( .B1(n7155), .B2(n7154), .A(n4477), .ZN(n7211) );
  AOI22_X1 U8841 ( .A1(n7211), .A2(n10138), .B1(n10137), .B2(n7155), .ZN(n7156) );
  OAI211_X1 U8842 ( .C1(n10132), .C2(n7213), .A(n7208), .B(n7156), .ZN(n7158)
         );
  NAND2_X1 U8843 ( .A1(n7158), .A2(n10177), .ZN(n7157) );
  OAI21_X1 U8844 ( .B1(n10177), .B2(n6011), .A(n7157), .ZN(P2_U3529) );
  INV_X1 U8845 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7160) );
  NAND2_X1 U8846 ( .A1(n7158), .A2(n10163), .ZN(n7159) );
  OAI21_X1 U8847 ( .B1(n10163), .B2(n7160), .A(n7159), .ZN(P2_U3478) );
  NAND2_X1 U8848 ( .A1(n7161), .A2(n7747), .ZN(n7164) );
  AOI22_X1 U8849 ( .A1(n7748), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7162), .B2(
        n7279), .ZN(n7163) );
  NAND2_X1 U8850 ( .A1(n7327), .A2(n8918), .ZN(n7166) );
  NAND2_X1 U8851 ( .A1(n9061), .A2(n8925), .ZN(n7165) );
  NAND2_X1 U8852 ( .A1(n7166), .A2(n7165), .ZN(n7167) );
  XNOR2_X1 U8853 ( .A(n7167), .B(n8922), .ZN(n7284) );
  AND2_X1 U8854 ( .A1(n9061), .A2(n8924), .ZN(n7168) );
  AOI21_X1 U8855 ( .B1(n7327), .B2(n8919), .A(n7168), .ZN(n7283) );
  XNOR2_X1 U8856 ( .A(n7284), .B(n7283), .ZN(n7178) );
  INV_X1 U8857 ( .A(n7169), .ZN(n7172) );
  INV_X1 U8858 ( .A(n7170), .ZN(n7171) );
  NAND2_X1 U8859 ( .A1(n7172), .A2(n7171), .ZN(n7173) );
  INV_X1 U8860 ( .A(n7178), .ZN(n7175) );
  INV_X1 U8861 ( .A(n7286), .ZN(n7176) );
  AOI21_X1 U8862 ( .B1(n7178), .B2(n7177), .A(n7176), .ZN(n7187) );
  OAI21_X1 U8863 ( .B1(n9043), .B2(n7776), .A(n7179), .ZN(n7185) );
  NAND2_X1 U8864 ( .A1(n6350), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7183) );
  OR2_X1 U8865 ( .A1(n7703), .A2(n9777), .ZN(n7182) );
  INV_X1 U8866 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7294) );
  XNOR2_X1 U8867 ( .A(n7296), .B(n7294), .ZN(n7401) );
  OR2_X1 U8868 ( .A1(n6349), .A2(n7401), .ZN(n7181) );
  INV_X1 U8869 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7402) );
  OR2_X1 U8870 ( .A1(n7679), .A2(n7402), .ZN(n7180) );
  NAND4_X1 U8871 ( .A1(n7183), .A2(n7182), .A3(n7181), .A4(n7180), .ZN(n9060)
         );
  INV_X1 U8872 ( .A(n9060), .ZN(n7310) );
  OAI22_X1 U8873 ( .A1(n7310), .A2(n9046), .B1(n9045), .B2(n7197), .ZN(n7184)
         );
  AOI211_X1 U8874 ( .C1(n7327), .C2(n9050), .A(n7185), .B(n7184), .ZN(n7186)
         );
  OAI21_X1 U8875 ( .B1(n7187), .B2(n9052), .A(n7186), .ZN(P1_U3222) );
  OR2_X1 U8876 ( .A1(n7327), .A2(n7397), .ZN(n7779) );
  NAND2_X1 U8877 ( .A1(n7327), .A2(n7397), .ZN(n7890) );
  NAND2_X1 U8878 ( .A1(n7189), .A2(n9785), .ZN(n7190) );
  INV_X1 U8879 ( .A(n7190), .ZN(n7188) );
  NAND2_X1 U8880 ( .A1(n7325), .A2(n7324), .ZN(n7390) );
  NAND2_X1 U8881 ( .A1(n7324), .A2(n7190), .ZN(n7191) );
  NAND2_X1 U8882 ( .A1(n7191), .A2(n7863), .ZN(n7192) );
  NAND2_X1 U8883 ( .A1(n7390), .A2(n7192), .ZN(n9778) );
  OR2_X1 U8884 ( .A1(n7777), .A2(n7776), .ZN(n7306) );
  XOR2_X1 U8885 ( .A(n7863), .B(n7309), .Z(n7195) );
  OAI22_X1 U8886 ( .A1(n7310), .A2(n9546), .B1(n7776), .B2(n9544), .ZN(n7194)
         );
  AOI21_X1 U8887 ( .B1(n7195), .B2(n9916), .A(n7194), .ZN(n7196) );
  OAI21_X1 U8888 ( .B1(n9920), .B2(n9778), .A(n7196), .ZN(n9781) );
  NAND2_X1 U8889 ( .A1(n9781), .A2(n9926), .ZN(n7204) );
  OAI22_X1 U8890 ( .A1(n9926), .A2(n7198), .B1(n7197), .B2(n9936), .ZN(n7202)
         );
  INV_X1 U8891 ( .A(n7199), .ZN(n7200) );
  INV_X1 U8892 ( .A(n7327), .ZN(n9780) );
  OAI211_X1 U8893 ( .C1(n7200), .C2(n9780), .A(n10005), .B(n7403), .ZN(n9779)
         );
  NOR2_X1 U8894 ( .A1(n9779), .A2(n6863), .ZN(n7201) );
  AOI211_X1 U8895 ( .C1(n7408), .C2(n7327), .A(n7202), .B(n7201), .ZN(n7203)
         );
  OAI211_X1 U8896 ( .C1(n9778), .C2(n9905), .A(n7204), .B(n7203), .ZN(P1_U3279) );
  AOI22_X1 U8897 ( .A1(n8646), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7205), .B2(
        n10071), .ZN(n7206) );
  OAI21_X1 U8898 ( .B1(n7207), .B2(n8639), .A(n7206), .ZN(n7210) );
  NOR2_X1 U8899 ( .A1(n7208), .A2(n8646), .ZN(n7209) );
  AOI211_X1 U8900 ( .C1(n7211), .C2(n8644), .A(n7210), .B(n7209), .ZN(n7212)
         );
  OAI21_X1 U8901 ( .B1(n8557), .B2(n7213), .A(n7212), .ZN(P2_U3287) );
  OR2_X1 U8902 ( .A1(n7356), .A2(n7214), .ZN(n7216) );
  NAND2_X1 U8903 ( .A1(n7216), .A2(n7215), .ZN(n7220) );
  NOR2_X1 U8904 ( .A1(n7218), .A2(n7217), .ZN(n7219) );
  XNOR2_X1 U8905 ( .A(n7220), .B(n7219), .ZN(n7225) );
  OAI21_X1 U8906 ( .B1(n8307), .B2(n7471), .A(n7221), .ZN(n7223) );
  OAI22_X1 U8907 ( .A1(n7231), .A2(n8310), .B1(n8309), .B2(n8103), .ZN(n7222)
         );
  AOI211_X1 U8908 ( .C1(n8728), .C2(n8314), .A(n7223), .B(n7222), .ZN(n7224)
         );
  OAI21_X1 U8909 ( .B1(n7225), .B2(n8316), .A(n7224), .ZN(P2_U3236) );
  OR2_X1 U8910 ( .A1(n7356), .A2(n7226), .ZN(n7228) );
  NAND2_X1 U8911 ( .A1(n7228), .A2(n7227), .ZN(n7230) );
  XNOR2_X1 U8912 ( .A(n7230), .B(n7229), .ZN(n7236) );
  OAI22_X1 U8913 ( .A1(n8307), .A2(n7373), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5334), .ZN(n7234) );
  OAI22_X1 U8914 ( .A1(n7232), .A2(n8310), .B1(n8309), .B2(n7231), .ZN(n7233)
         );
  AOI211_X1 U8915 ( .C1(n5739), .C2(n8314), .A(n7234), .B(n7233), .ZN(n7235)
         );
  OAI21_X1 U8916 ( .B1(n7236), .B2(n8316), .A(n7235), .ZN(P2_U3238) );
  NAND2_X1 U8917 ( .A1(n7238), .A2(n7241), .ZN(n7239) );
  NAND2_X1 U8918 ( .A1(n7237), .A2(n7239), .ZN(n10146) );
  NAND2_X1 U8919 ( .A1(n7240), .A2(n8067), .ZN(n7242) );
  XNOR2_X1 U8920 ( .A(n7242), .B(n7241), .ZN(n7245) );
  OAI22_X1 U8921 ( .A1(n7243), .A2(n8624), .B1(n7344), .B2(n8622), .ZN(n7244)
         );
  AOI21_X1 U8922 ( .B1(n7245), .B2(n10061), .A(n7244), .ZN(n7246) );
  OAI21_X1 U8923 ( .B1(n10146), .B2(n8630), .A(n7246), .ZN(n10149) );
  NAND2_X1 U8924 ( .A1(n10149), .A2(n6401), .ZN(n7253) );
  OAI22_X1 U8925 ( .A1(n6401), .A2(n7248), .B1(n7247), .B2(n8604), .ZN(n7250)
         );
  OAI21_X1 U8926 ( .B1(n4477), .B2(n10147), .A(n7372), .ZN(n10148) );
  NOR2_X1 U8927 ( .A1(n10148), .A2(n8429), .ZN(n7249) );
  AOI211_X1 U8928 ( .C1(n8619), .C2(n7251), .A(n7250), .B(n7249), .ZN(n7252)
         );
  OAI211_X1 U8929 ( .C1(n10146), .C2(n8641), .A(n7253), .B(n7252), .ZN(
        P2_U3286) );
  NAND2_X1 U8930 ( .A1(n7255), .A2(n7254), .ZN(n7260) );
  OR2_X1 U8931 ( .A1(n7356), .A2(n7256), .ZN(n7258) );
  NAND2_X1 U8932 ( .A1(n7258), .A2(n7257), .ZN(n7259) );
  XOR2_X1 U8933 ( .A(n7260), .B(n7259), .Z(n7265) );
  OAI21_X1 U8934 ( .B1(n8307), .B2(n7347), .A(n7261), .ZN(n7263) );
  OAI22_X1 U8935 ( .A1(n7344), .A2(n8310), .B1(n8309), .B2(n7440), .ZN(n7262)
         );
  AOI211_X1 U8936 ( .C1(n7350), .C2(n8314), .A(n7263), .B(n7262), .ZN(n7264)
         );
  OAI21_X1 U8937 ( .B1(n7265), .B2(n8316), .A(n7264), .ZN(P2_U3226) );
  INV_X1 U8938 ( .A(n7266), .ZN(n7267) );
  AND2_X2 U8939 ( .A1(n7268), .A2(n7267), .ZN(n10049) );
  AND2_X1 U8940 ( .A1(n9203), .A2(n7844), .ZN(n7835) );
  NAND2_X1 U8941 ( .A1(n6177), .A2(n7835), .ZN(n10009) );
  AOI21_X1 U8942 ( .B1(n10004), .B2(n7270), .A(n7269), .ZN(n7271) );
  OAI211_X1 U8943 ( .C1(n7273), .C2(n10009), .A(n7272), .B(n7271), .ZN(n7275)
         );
  NAND2_X1 U8944 ( .A1(n7275), .A2(n10049), .ZN(n7274) );
  OAI21_X1 U8945 ( .B1(n10049), .B2(n6821), .A(n7274), .ZN(P1_U3533) );
  INV_X1 U8946 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7277) );
  NAND2_X1 U8947 ( .A1(n7275), .A2(n10037), .ZN(n7276) );
  OAI21_X1 U8948 ( .B1(n10037), .B2(n7277), .A(n7276), .ZN(P1_U3484) );
  NAND2_X1 U8949 ( .A1(n7278), .A2(n7747), .ZN(n7282) );
  AOI22_X1 U8950 ( .A1(n7748), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7280), .B2(
        n7279), .ZN(n7281) );
  NAND2_X1 U8951 ( .A1(n7284), .A2(n7283), .ZN(n7285) );
  NAND2_X1 U8952 ( .A1(n7286), .A2(n7285), .ZN(n8768) );
  AND2_X1 U8953 ( .A1(n9060), .A2(n8924), .ZN(n7287) );
  AOI21_X1 U8954 ( .B1(n7407), .B2(n8919), .A(n7287), .ZN(n8765) );
  NAND2_X1 U8955 ( .A1(n7407), .A2(n8918), .ZN(n7289) );
  NAND2_X1 U8956 ( .A1(n9060), .A2(n8925), .ZN(n7288) );
  NAND2_X1 U8957 ( .A1(n7289), .A2(n7288), .ZN(n7290) );
  XNOR2_X1 U8958 ( .A(n7290), .B(n8922), .ZN(n8766) );
  XOR2_X1 U8959 ( .A(n8765), .B(n8766), .Z(n7291) );
  XNOR2_X1 U8960 ( .A(n8768), .B(n7291), .ZN(n7292) );
  NAND2_X1 U8961 ( .A1(n7292), .A2(n8982), .ZN(n7305) );
  INV_X1 U8962 ( .A(n7293), .ZN(n7303) );
  NAND2_X1 U8963 ( .A1(n6350), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7301) );
  OR2_X1 U8964 ( .A1(n7703), .A2(n9771), .ZN(n7300) );
  OAI21_X1 U8965 ( .B1(n7296), .B2(n7294), .A(n9388), .ZN(n7297) );
  NAND2_X1 U8966 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG3_REG_14__SCAN_IN), 
        .ZN(n7295) );
  NAND2_X1 U8967 ( .A1(n7297), .A2(n7315), .ZN(n8893) );
  OR2_X1 U8968 ( .A1(n6349), .A2(n8893), .ZN(n7299) );
  OR2_X1 U8969 ( .A1(n7679), .A2(n6972), .ZN(n7298) );
  NAND4_X1 U8970 ( .A1(n7301), .A2(n7300), .A3(n7299), .A4(n7298), .ZN(n9059)
         );
  INV_X1 U8971 ( .A(n9059), .ZN(n9042) );
  OAI22_X1 U8972 ( .A1(n9042), .A2(n9046), .B1(n9045), .B2(n7401), .ZN(n7302)
         );
  AOI211_X1 U8973 ( .C1(n8943), .C2(n9061), .A(n7303), .B(n7302), .ZN(n7304)
         );
  OAI211_X1 U8974 ( .C1(n4486), .C2(n9024), .A(n7305), .B(n7304), .ZN(P1_U3232) );
  INV_X1 U8975 ( .A(n7306), .ZN(n7307) );
  NAND2_X1 U8976 ( .A1(n7890), .A2(n7307), .ZN(n7308) );
  NAND2_X1 U8977 ( .A1(n7308), .A2(n7779), .ZN(n7893) );
  OR2_X1 U8978 ( .A1(n7407), .A2(n7310), .ZN(n7780) );
  NAND2_X1 U8979 ( .A1(n7407), .A2(n7310), .ZN(n7778) );
  NAND2_X1 U8980 ( .A1(n7311), .A2(n7747), .ZN(n7314) );
  AOI22_X1 U8981 ( .A1(n7748), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7312), .B2(
        n7279), .ZN(n7313) );
  XNOR2_X1 U8982 ( .A(n8774), .B(n9042), .ZN(n7421) );
  INV_X1 U8983 ( .A(n7421), .ZN(n7868) );
  XNOR2_X1 U8984 ( .A(n7422), .B(n7868), .ZN(n7321) );
  NAND2_X1 U8985 ( .A1(n6350), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7320) );
  OR2_X1 U8986 ( .A1(n7703), .A2(n9289), .ZN(n7319) );
  OR2_X1 U8987 ( .A1(n7679), .A2(n9344), .ZN(n7318) );
  INV_X1 U8988 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9415) );
  AND2_X1 U8989 ( .A1(n7315), .A2(n9415), .ZN(n7316) );
  OR2_X1 U8990 ( .A1(n7316), .A2(n7423), .ZN(n9044) );
  OR2_X1 U8991 ( .A1(n6349), .A2(n9044), .ZN(n7317) );
  NAND4_X1 U8992 ( .A1(n7320), .A2(n7319), .A3(n7318), .A4(n7317), .ZN(n9058)
         );
  AOI222_X1 U8993 ( .A1(n9916), .A2(n7321), .B1(n9058), .B2(n9911), .C1(n9060), 
        .C2(n9913), .ZN(n9767) );
  OAI22_X1 U8994 ( .A1(n9926), .A2(n6972), .B1(n8893), .B2(n9936), .ZN(n7323)
         );
  AND2_X2 U8995 ( .A1(n4406), .A2(n9768), .ZN(n7416) );
  INV_X1 U8996 ( .A(n7416), .ZN(n7418) );
  OAI211_X1 U8997 ( .C1(n9768), .C2(n4406), .A(n7418), .B(n10005), .ZN(n9766)
         );
  NOR2_X1 U8998 ( .A1(n9766), .A2(n6863), .ZN(n7322) );
  AOI211_X1 U8999 ( .C1(n7408), .C2(n8774), .A(n7323), .B(n7322), .ZN(n7332)
         );
  NAND2_X1 U9000 ( .A1(n7326), .A2(n7325), .ZN(n7329) );
  NAND2_X1 U9001 ( .A1(n7327), .A2(n9061), .ZN(n7389) );
  NAND2_X1 U9002 ( .A1(n7329), .A2(n7328), .ZN(n7393) );
  XNOR2_X1 U9003 ( .A(n7411), .B(n7421), .ZN(n9770) );
  NAND2_X1 U9004 ( .A1(n9770), .A2(n7330), .ZN(n7331) );
  OAI211_X1 U9005 ( .C1(n9767), .C2(n4382), .A(n7332), .B(n7331), .ZN(P1_U3277) );
  INV_X1 U9006 ( .A(n7651), .ZN(n7336) );
  OAI222_X1 U9007 ( .A1(n8761), .A2(n7334), .B1(n4385), .B2(n7336), .C1(
        P2_U3152), .C2(n7333), .ZN(P2_U3333) );
  OAI222_X1 U9008 ( .A1(n9698), .A2(n9376), .B1(n9695), .B2(n7336), .C1(n7335), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9009 ( .A(n7663), .ZN(n7387) );
  OAI222_X1 U9010 ( .A1(n9695), .A2(n7387), .B1(P1_U3084), .B2(n7338), .C1(
        n7337), .C2(n9698), .ZN(P1_U3327) );
  NAND2_X1 U9011 ( .A1(n7237), .A2(n7339), .ZN(n7461) );
  AND2_X1 U9012 ( .A1(n7461), .A2(n7340), .ZN(n7341) );
  XNOR2_X1 U9013 ( .A(n7341), .B(n8196), .ZN(n10160) );
  INV_X1 U9014 ( .A(n10160), .ZN(n7354) );
  XNOR2_X1 U9015 ( .A(n7342), .B(n8196), .ZN(n7343) );
  OAI222_X1 U9016 ( .A1(n8622), .A2(n7440), .B1(n8624), .B2(n7344), .C1(n8612), 
        .C2(n7343), .ZN(n10157) );
  INV_X1 U9017 ( .A(n7345), .ZN(n7371) );
  INV_X1 U9018 ( .A(n7346), .ZN(n7470) );
  OAI21_X1 U9019 ( .B1(n10154), .B2(n7371), .A(n7470), .ZN(n10156) );
  INV_X1 U9020 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7348) );
  OAI22_X1 U9021 ( .A1(n6401), .A2(n7348), .B1(n7347), .B2(n8604), .ZN(n7349)
         );
  AOI21_X1 U9022 ( .B1(n7350), .B2(n8619), .A(n7349), .ZN(n7351) );
  OAI21_X1 U9023 ( .B1(n10156), .B2(n8429), .A(n7351), .ZN(n7352) );
  AOI21_X1 U9024 ( .B1(n10157), .B2(n6401), .A(n7352), .ZN(n7353) );
  OAI21_X1 U9025 ( .B1(n7354), .B2(n8557), .A(n7353), .ZN(P2_U3284) );
  OR2_X1 U9026 ( .A1(n7356), .A2(n7355), .ZN(n7359) );
  AND2_X1 U9027 ( .A1(n7359), .A2(n7357), .ZN(n7361) );
  NAND2_X1 U9028 ( .A1(n7359), .A2(n7358), .ZN(n7360) );
  OAI21_X1 U9029 ( .B1(n7362), .B2(n7361), .A(n7360), .ZN(n7363) );
  NAND2_X1 U9030 ( .A1(n7363), .A2(n8321), .ZN(n7368) );
  INV_X1 U9031 ( .A(n7364), .ZN(n7437) );
  NAND2_X1 U9032 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(n4374), .ZN(n8363) );
  INV_X1 U9033 ( .A(n8363), .ZN(n7366) );
  OAI22_X1 U9034 ( .A1(n7440), .A2(n8310), .B1(n8309), .B2(n8625), .ZN(n7365)
         );
  AOI211_X1 U9035 ( .C1(n7437), .C2(n8336), .A(n7366), .B(n7365), .ZN(n7367)
         );
  OAI211_X1 U9036 ( .C1(n4730), .C2(n8338), .A(n7368), .B(n7367), .ZN(P2_U3217) );
  NAND2_X1 U9037 ( .A1(n7237), .A2(n7369), .ZN(n7370) );
  XNOR2_X1 U9038 ( .A(n7370), .B(n7380), .ZN(n8736) );
  AOI21_X1 U9039 ( .B1(n5739), .B2(n7372), .A(n7371), .ZN(n8733) );
  INV_X1 U9040 ( .A(n7373), .ZN(n7374) );
  AOI22_X1 U9041 ( .A1(n8646), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7374), .B2(
        n10071), .ZN(n7375) );
  OAI21_X1 U9042 ( .B1(n4515), .B2(n8639), .A(n7375), .ZN(n7384) );
  NAND2_X1 U9043 ( .A1(n7377), .A2(n7376), .ZN(n7379) );
  AND2_X1 U9044 ( .A1(n7379), .A2(n7378), .ZN(n7381) );
  XNOR2_X1 U9045 ( .A(n7381), .B(n7380), .ZN(n7382) );
  AOI222_X1 U9046 ( .A1(n10061), .A2(n7382), .B1(n8348), .B2(n10065), .C1(
        n8350), .C2(n10066), .ZN(n8735) );
  NOR2_X1 U9047 ( .A1(n8735), .A2(n8646), .ZN(n7383) );
  AOI211_X1 U9048 ( .C1(n8733), .C2(n8644), .A(n7384), .B(n7383), .ZN(n7385)
         );
  OAI21_X1 U9049 ( .B1(n8557), .B2(n8736), .A(n7385), .ZN(P2_U3285) );
  OAI222_X1 U9050 ( .A1(P2_U3152), .A2(n7388), .B1(n4385), .B2(n7387), .C1(
        n7386), .C2(n8761), .ZN(P2_U3332) );
  NAND2_X1 U9051 ( .A1(n7390), .A2(n7389), .ZN(n7391) );
  NOR2_X1 U9052 ( .A1(n7391), .A2(n7865), .ZN(n7392) );
  OR2_X1 U9053 ( .A1(n7393), .A2(n7392), .ZN(n9772) );
  OAI21_X1 U9054 ( .B1(n7396), .B2(n7395), .A(n7394), .ZN(n7399) );
  OAI22_X1 U9055 ( .A1(n7397), .A2(n9544), .B1(n9042), .B2(n9546), .ZN(n7398)
         );
  AOI21_X1 U9056 ( .B1(n7399), .B2(n9916), .A(n7398), .ZN(n7400) );
  OAI21_X1 U9057 ( .B1(n9772), .B2(n9920), .A(n7400), .ZN(n9774) );
  NAND2_X1 U9058 ( .A1(n9774), .A2(n9926), .ZN(n7410) );
  OAI22_X1 U9059 ( .A1(n9926), .A2(n7402), .B1(n7401), .B2(n9936), .ZN(n7406)
         );
  AND2_X1 U9060 ( .A1(n7403), .A2(n7407), .ZN(n7404) );
  OR2_X1 U9061 ( .A1(n7404), .A2(n4406), .ZN(n9773) );
  NOR2_X1 U9062 ( .A1(n9773), .A2(n9931), .ZN(n7405) );
  AOI211_X1 U9063 ( .C1(n7408), .C2(n7407), .A(n7406), .B(n7405), .ZN(n7409)
         );
  OAI211_X1 U9064 ( .C1(n9772), .C2(n9905), .A(n7410), .B(n7409), .ZN(P1_U3278) );
  NAND2_X1 U9065 ( .A1(n7412), .A2(n7747), .ZN(n7415) );
  INV_X1 U9066 ( .A(n9076), .ZN(n7413) );
  AOI22_X1 U9067 ( .A1(n7748), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7413), .B2(
        n7279), .ZN(n7414) );
  NAND2_X1 U9068 ( .A1(n9669), .A2(n8967), .ZN(n7923) );
  XNOR2_X1 U9069 ( .A(n7482), .B(n7786), .ZN(n9673) );
  NAND2_X1 U9070 ( .A1(n7416), .A2(n7481), .ZN(n7487) );
  INV_X1 U9071 ( .A(n7487), .ZN(n7417) );
  AOI21_X1 U9072 ( .B1(n9669), .B2(n7418), .A(n7417), .ZN(n9670) );
  INV_X1 U9073 ( .A(n9044), .ZN(n7419) );
  AOI22_X1 U9074 ( .A1(n4382), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7419), .B2(
        n9923), .ZN(n7420) );
  OAI21_X1 U9075 ( .B1(n7481), .B2(n9930), .A(n7420), .ZN(n7431) );
  OR2_X1 U9076 ( .A1(n8774), .A2(n9042), .ZN(n7781) );
  OAI21_X1 U9077 ( .B1(n7422), .B2(n7421), .A(n7781), .ZN(n7500) );
  INV_X1 U9078 ( .A(n7786), .ZN(n7867) );
  XNOR2_X1 U9079 ( .A(n7500), .B(n7867), .ZN(n7429) );
  INV_X1 U9080 ( .A(n7703), .ZN(n7666) );
  NAND2_X1 U9081 ( .A1(n7666), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7428) );
  INV_X1 U9082 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9231) );
  OR2_X1 U9083 ( .A1(n7719), .A2(n9231), .ZN(n7427) );
  NOR2_X1 U9084 ( .A1(n7423), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7424) );
  OR2_X1 U9085 ( .A1(n7492), .A2(n7424), .ZN(n8968) );
  OR2_X1 U9086 ( .A1(n6349), .A2(n8968), .ZN(n7426) );
  INV_X1 U9087 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7489) );
  OR2_X1 U9088 ( .A1(n7679), .A2(n7489), .ZN(n7425) );
  NAND4_X1 U9089 ( .A1(n7428), .A2(n7427), .A3(n7426), .A4(n7425), .ZN(n9593)
         );
  AOI222_X1 U9090 ( .A1(n9916), .A2(n7429), .B1(n9593), .B2(n9911), .C1(n9059), 
        .C2(n9913), .ZN(n9672) );
  NOR2_X1 U9091 ( .A1(n9672), .A2(n4382), .ZN(n7430) );
  AOI211_X1 U9092 ( .C1(n9670), .C2(n9909), .A(n7431), .B(n7430), .ZN(n7432)
         );
  OAI21_X1 U9093 ( .B1(n9597), .B2(n9673), .A(n7432), .ZN(P1_U3276) );
  AND2_X1 U9094 ( .A1(n7461), .A2(n7433), .ZN(n7465) );
  OR2_X1 U9095 ( .A1(n7465), .A2(n7434), .ZN(n7435) );
  XNOR2_X1 U9096 ( .A(n7435), .B(n8200), .ZN(n8727) );
  INV_X1 U9097 ( .A(n7451), .ZN(n7436) );
  AOI21_X1 U9098 ( .B1(n8723), .B2(n7468), .A(n7436), .ZN(n8724) );
  AOI22_X1 U9099 ( .A1(n8646), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7437), .B2(
        n10071), .ZN(n7438) );
  OAI21_X1 U9100 ( .B1(n4730), .B2(n8639), .A(n7438), .ZN(n7445) );
  NAND2_X1 U9101 ( .A1(n7476), .A2(n8197), .ZN(n7475) );
  NAND2_X1 U9102 ( .A1(n7475), .A2(n8095), .ZN(n7439) );
  AOI21_X1 U9103 ( .B1(n7439), .B2(n8200), .A(n8612), .ZN(n7443) );
  OR2_X1 U9104 ( .A1(n7439), .A2(n8200), .ZN(n7442) );
  OAI22_X1 U9105 ( .A1(n7440), .A2(n8624), .B1(n8625), .B2(n8622), .ZN(n7441)
         );
  AOI21_X1 U9106 ( .B1(n7443), .B2(n7442), .A(n7441), .ZN(n8726) );
  NOR2_X1 U9107 ( .A1(n8726), .A2(n8646), .ZN(n7444) );
  AOI211_X1 U9108 ( .C1(n8724), .C2(n8644), .A(n7445), .B(n7444), .ZN(n7446)
         );
  OAI21_X1 U9109 ( .B1(n8727), .B2(n8557), .A(n7446), .ZN(P2_U3282) );
  XNOR2_X1 U9110 ( .A(n7447), .B(n8201), .ZN(n7448) );
  AOI222_X1 U9111 ( .A1(n10061), .A2(n7448), .B1(n8346), .B2(n10066), .C1(
        n8344), .C2(n10065), .ZN(n8721) );
  OAI21_X1 U9112 ( .B1(n7450), .B2(n8201), .A(n7449), .ZN(n8717) );
  NAND2_X1 U9113 ( .A1(n8717), .A2(n10077), .ZN(n7457) );
  AOI21_X1 U9114 ( .B1(n8718), .B2(n7451), .A(n8634), .ZN(n8719) );
  INV_X1 U9115 ( .A(n8718), .ZN(n7452) );
  NOR2_X1 U9116 ( .A1(n7452), .A2(n8639), .ZN(n7455) );
  OAI22_X1 U9117 ( .A1(n6401), .A2(n7453), .B1(n7528), .B2(n8604), .ZN(n7454)
         );
  AOI211_X1 U9118 ( .C1(n8719), .C2(n8644), .A(n7455), .B(n7454), .ZN(n7456)
         );
  OAI211_X1 U9119 ( .C1(n8646), .C2(n8721), .A(n7457), .B(n7456), .ZN(P2_U3281) );
  INV_X1 U9120 ( .A(n7675), .ZN(n7534) );
  AOI21_X1 U9121 ( .B1(n9699), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7458), .ZN(
        n7459) );
  OAI21_X1 U9122 ( .B1(n7534), .B2(n8009), .A(n7459), .ZN(P1_U3326) );
  AND2_X1 U9123 ( .A1(n7461), .A2(n7460), .ZN(n7463) );
  OR2_X1 U9124 ( .A1(n7463), .A2(n7462), .ZN(n7467) );
  NOR2_X1 U9125 ( .A1(n7465), .A2(n7464), .ZN(n7466) );
  OAI21_X1 U9126 ( .B1(n7467), .B2(n8101), .A(n7466), .ZN(n8732) );
  INV_X1 U9127 ( .A(n7468), .ZN(n7469) );
  AOI21_X1 U9128 ( .B1(n8728), .B2(n7470), .A(n7469), .ZN(n8729) );
  INV_X1 U9129 ( .A(n7471), .ZN(n7472) );
  AOI22_X1 U9130 ( .A1(n8646), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7472), .B2(
        n10071), .ZN(n7473) );
  OAI21_X1 U9131 ( .B1(n7474), .B2(n8639), .A(n7473), .ZN(n7479) );
  OAI21_X1 U9132 ( .B1(n8197), .B2(n7476), .A(n7475), .ZN(n7477) );
  AOI222_X1 U9133 ( .A1(n10061), .A2(n7477), .B1(n8346), .B2(n10065), .C1(
        n8348), .C2(n10066), .ZN(n8731) );
  NOR2_X1 U9134 ( .A1(n8731), .A2(n8646), .ZN(n7478) );
  AOI211_X1 U9135 ( .C1(n8729), .C2(n8644), .A(n7479), .B(n7478), .ZN(n7480)
         );
  OAI21_X1 U9136 ( .B1(n8557), .B2(n8732), .A(n7480), .ZN(P2_U3283) );
  NAND2_X1 U9137 ( .A1(n7483), .A2(n7747), .ZN(n7485) );
  AOI22_X1 U9138 ( .A1(n7748), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9092), .B2(
        n7279), .ZN(n7484) );
  INV_X1 U9139 ( .A(n9593), .ZN(n9047) );
  OR2_X1 U9140 ( .A1(n9666), .A2(n9047), .ZN(n7790) );
  NAND2_X1 U9141 ( .A1(n9666), .A2(n9047), .ZN(n9586) );
  NAND2_X1 U9142 ( .A1(n7790), .A2(n9586), .ZN(n7565) );
  XNOR2_X1 U9143 ( .A(n7566), .B(n7565), .ZN(n9668) );
  OR2_X2 U9144 ( .A1(n7487), .A2(n9666), .ZN(n9578) );
  INV_X1 U9145 ( .A(n9578), .ZN(n7486) );
  AOI211_X1 U9146 ( .C1(n9666), .C2(n7487), .A(n10029), .B(n7486), .ZN(n9665)
         );
  INV_X1 U9147 ( .A(n9666), .ZN(n7488) );
  NOR2_X1 U9148 ( .A1(n7488), .A2(n9930), .ZN(n7491) );
  OAI22_X1 U9149 ( .A1(n9926), .A2(n7489), .B1(n8968), .B2(n9936), .ZN(n7490)
         );
  AOI211_X1 U9150 ( .C1(n9665), .C2(n9573), .A(n7491), .B(n7490), .ZN(n7504)
         );
  NOR2_X1 U9151 ( .A1(n7492), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7493) );
  OR2_X1 U9152 ( .A1(n7574), .A2(n7493), .ZN(n9579) );
  OR2_X1 U9153 ( .A1(n6349), .A2(n9579), .ZN(n7499) );
  INV_X1 U9154 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9296) );
  OR2_X1 U9155 ( .A1(n7703), .A2(n9296), .ZN(n7498) );
  INV_X1 U9156 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n7494) );
  OR2_X1 U9157 ( .A1(n7719), .A2(n7494), .ZN(n7497) );
  INV_X1 U9158 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7495) );
  OR2_X1 U9159 ( .A1(n7679), .A2(n7495), .ZN(n7496) );
  NAND4_X1 U9160 ( .A1(n7499), .A2(n7498), .A3(n7497), .A4(n7496), .ZN(n9568)
         );
  INV_X1 U9161 ( .A(n9568), .ZN(n9019) );
  NAND2_X1 U9162 ( .A1(n7500), .A2(n7923), .ZN(n7710) );
  NAND2_X1 U9163 ( .A1(n7710), .A2(n7709), .ZN(n7501) );
  INV_X1 U9164 ( .A(n7565), .ZN(n7870) );
  XNOR2_X1 U9165 ( .A(n7501), .B(n7870), .ZN(n7502) );
  OAI222_X1 U9166 ( .A1(n9546), .A2(n9019), .B1(n9544), .B2(n8967), .C1(n9588), 
        .C2(n7502), .ZN(n9664) );
  NAND2_X1 U9167 ( .A1(n9664), .A2(n9926), .ZN(n7503) );
  OAI211_X1 U9168 ( .C1(n9668), .C2(n9597), .A(n7504), .B(n7503), .ZN(P1_U3275) );
  NAND2_X1 U9169 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n7527) );
  INV_X1 U9170 ( .A(n7527), .ZN(n7509) );
  AOI211_X1 U9171 ( .C1(n7507), .C2(n7506), .A(n7505), .B(n10051), .ZN(n7508)
         );
  AOI211_X1 U9172 ( .C1(n10056), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n7509), .B(
        n7508), .ZN(n7514) );
  OAI21_X1 U9173 ( .B1(n7511), .B2(n7453), .A(n7510), .ZN(n7512) );
  NAND2_X1 U9174 ( .A1(n10055), .A2(n7512), .ZN(n7513) );
  OAI211_X1 U9175 ( .C1(n8402), .C2(n7515), .A(n7514), .B(n7513), .ZN(P2_U3260) );
  XNOR2_X1 U9176 ( .A(n7517), .B(n7516), .ZN(n7522) );
  OAI22_X1 U9177 ( .A1(n8307), .A2(n8605), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7518), .ZN(n7520) );
  OAI22_X1 U9178 ( .A1(n8613), .A2(n8310), .B1(n8309), .B2(n8614), .ZN(n7519)
         );
  AOI211_X1 U9179 ( .C1(n8709), .C2(n8314), .A(n7520), .B(n7519), .ZN(n7521)
         );
  OAI21_X1 U9180 ( .B1(n7522), .B2(n8316), .A(n7521), .ZN(P2_U3230) );
  NAND2_X1 U9181 ( .A1(n7524), .A2(n7523), .ZN(n7535) );
  OAI21_X1 U9182 ( .B1(n7524), .B2(n7523), .A(n7535), .ZN(n7525) );
  NOR2_X1 U9183 ( .A1(n7525), .A2(n7526), .ZN(n7538) );
  AOI21_X1 U9184 ( .B1(n7526), .B2(n7525), .A(n7538), .ZN(n7532) );
  OAI21_X1 U9185 ( .B1(n8307), .B2(n7528), .A(n7527), .ZN(n7530) );
  OAI22_X1 U9186 ( .A1(n8613), .A2(n8309), .B1(n8310), .B2(n8103), .ZN(n7529)
         );
  AOI211_X1 U9187 ( .C1(n8718), .C2(n8314), .A(n7530), .B(n7529), .ZN(n7531)
         );
  OAI21_X1 U9188 ( .B1(n7532), .B2(n8316), .A(n7531), .ZN(P2_U3243) );
  OAI222_X1 U9189 ( .A1(n8761), .A2(n9222), .B1(n4385), .B2(n7534), .C1(n4374), 
        .C2(n7533), .ZN(P2_U3331) );
  INV_X1 U9190 ( .A(n7535), .ZN(n7537) );
  NOR3_X1 U9191 ( .A1(n7538), .A2(n7537), .A3(n7536), .ZN(n7542) );
  INV_X1 U9192 ( .A(n7539), .ZN(n7541) );
  OAI21_X1 U9193 ( .B1(n7542), .B2(n7541), .A(n8321), .ZN(n7546) );
  INV_X1 U9194 ( .A(n7543), .ZN(n8637) );
  AND2_X1 U9195 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8377) );
  OAI22_X1 U9196 ( .A1(n8625), .A2(n8310), .B1(n8309), .B2(n8623), .ZN(n7544)
         );
  AOI211_X1 U9197 ( .C1(n8336), .C2(n8637), .A(n8377), .B(n7544), .ZN(n7545)
         );
  OAI211_X1 U9198 ( .C1(n8640), .C2(n8338), .A(n7546), .B(n7545), .ZN(P2_U3228) );
  XNOR2_X1 U9199 ( .A(n7548), .B(n7547), .ZN(n7552) );
  NAND2_X1 U9200 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8396) );
  OAI21_X1 U9201 ( .B1(n8307), .B2(n8589), .A(n8396), .ZN(n7550) );
  OAI22_X1 U9202 ( .A1(n8623), .A2(n8310), .B1(n8309), .B2(n8311), .ZN(n7549)
         );
  AOI211_X1 U9203 ( .C1(n8702), .C2(n8314), .A(n7550), .B(n7549), .ZN(n7551)
         );
  OAI21_X1 U9204 ( .B1(n7552), .B2(n8316), .A(n7551), .ZN(P2_U3240) );
  INV_X1 U9205 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7564) );
  INV_X1 U9206 ( .A(n7553), .ZN(n7556) );
  NAND2_X1 U9207 ( .A1(n7556), .A2(SI_29_), .ZN(n7555) );
  AND2_X1 U9208 ( .A1(n7554), .A2(n7555), .ZN(n7561) );
  INV_X1 U9209 ( .A(n7555), .ZN(n7560) );
  OR2_X1 U9210 ( .A1(n7556), .A2(SI_29_), .ZN(n7557) );
  AND2_X1 U9211 ( .A1(n7558), .A2(n7557), .ZN(n7559) );
  MUX2_X1 U9212 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7743), .Z(n7739) );
  INV_X1 U9213 ( .A(n8014), .ZN(n8248) );
  OAI222_X1 U9214 ( .A1(n9698), .A2(n7564), .B1(n9695), .B2(n8248), .C1(
        P1_U3084), .C2(n7563), .ZN(P1_U3323) );
  NAND2_X1 U9215 ( .A1(n7567), .A2(n7747), .ZN(n7569) );
  AOI22_X1 U9216 ( .A1(n7748), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9109), .B2(
        n7279), .ZN(n7568) );
  NOR2_X1 U9217 ( .A1(n9659), .A2(n9568), .ZN(n7570) );
  NAND2_X1 U9218 ( .A1(n9659), .A2(n9568), .ZN(n7795) );
  NAND2_X1 U9219 ( .A1(n7571), .A2(n7747), .ZN(n7573) );
  AOI22_X1 U9220 ( .A1(n7748), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9119), .B2(
        n7279), .ZN(n7572) );
  OR2_X1 U9221 ( .A1(n7574), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7575) );
  NAND2_X1 U9222 ( .A1(n7574), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7584) );
  NAND2_X1 U9223 ( .A1(n7575), .A2(n7584), .ZN(n9560) );
  OR2_X1 U9224 ( .A1(n9560), .A2(n6349), .ZN(n7580) );
  INV_X1 U9225 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9253) );
  OR2_X1 U9226 ( .A1(n7719), .A2(n9253), .ZN(n7579) );
  INV_X1 U9227 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9286) );
  OR2_X1 U9228 ( .A1(n7703), .A2(n9286), .ZN(n7578) );
  INV_X1 U9229 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n7576) );
  OR2_X1 U9230 ( .A1(n7679), .A2(n7576), .ZN(n7577) );
  NAND4_X1 U9231 ( .A1(n7580), .A2(n7579), .A3(n7578), .A4(n7577), .ZN(n9583)
         );
  INV_X1 U9232 ( .A(n9583), .ZN(n9543) );
  OR2_X1 U9233 ( .A1(n9655), .A2(n9543), .ZN(n7802) );
  NAND2_X1 U9234 ( .A1(n9655), .A2(n9543), .ZN(n7932) );
  NAND2_X1 U9235 ( .A1(n9558), .A2(n9557), .ZN(n9556) );
  INV_X1 U9236 ( .A(n9655), .ZN(n9563) );
  NAND2_X1 U9237 ( .A1(n7581), .A2(n7747), .ZN(n7583) );
  AOI22_X1 U9238 ( .A1(n7748), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9203), .B2(
        n7279), .ZN(n7582) );
  OAI21_X1 U9239 ( .B1(n7585), .B2(P1_REG3_REG_19__SCAN_IN), .A(n7596), .ZN(
        n9549) );
  INV_X1 U9240 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n7586) );
  OR2_X1 U9241 ( .A1(n7719), .A2(n7586), .ZN(n7588) );
  INV_X1 U9242 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9403) );
  OR2_X1 U9243 ( .A1(n7703), .A2(n9403), .ZN(n7587) );
  AND2_X1 U9244 ( .A1(n7588), .A2(n7587), .ZN(n7590) );
  NAND2_X1 U9245 ( .A1(n7635), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7589) );
  OAI211_X1 U9246 ( .C1(n9549), .C2(n6349), .A(n7590), .B(n7589), .ZN(n9569)
         );
  INV_X1 U9247 ( .A(n9569), .ZN(n8994) );
  NAND2_X1 U9248 ( .A1(n9553), .A2(n8994), .ZN(n7592) );
  NAND2_X1 U9249 ( .A1(n7593), .A2(n7747), .ZN(n7595) );
  NAND2_X1 U9250 ( .A1(n7748), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7594) );
  INV_X1 U9251 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8993) );
  INV_X1 U9252 ( .A(n7608), .ZN(n7609) );
  NAND2_X1 U9253 ( .A1(n7596), .A2(n8993), .ZN(n7597) );
  NAND2_X1 U9254 ( .A1(n7609), .A2(n7597), .ZN(n9527) );
  OR2_X1 U9255 ( .A1(n9527), .A2(n6349), .ZN(n7603) );
  INV_X1 U9256 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n7600) );
  NAND2_X1 U9257 ( .A1(n7635), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n7599) );
  NAND2_X1 U9258 ( .A1(n6350), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7598) );
  OAI211_X1 U9259 ( .C1(n7703), .C2(n7600), .A(n7599), .B(n7598), .ZN(n7601)
         );
  INV_X1 U9260 ( .A(n7601), .ZN(n7602) );
  NAND2_X1 U9261 ( .A1(n7603), .A2(n7602), .ZN(n9518) );
  NAND2_X1 U9262 ( .A1(n9644), .A2(n9518), .ZN(n7604) );
  INV_X1 U9263 ( .A(n9518), .ZN(n9545) );
  NAND2_X1 U9264 ( .A1(n7605), .A2(n7747), .ZN(n7607) );
  NAND2_X1 U9265 ( .A1(n7748), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7606) );
  NAND2_X1 U9266 ( .A1(n7608), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7622) );
  INV_X1 U9267 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8951) );
  NAND2_X1 U9268 ( .A1(n7609), .A2(n8951), .ZN(n7610) );
  NAND2_X1 U9269 ( .A1(n7622), .A2(n7610), .ZN(n9511) );
  OR2_X1 U9270 ( .A1(n9511), .A2(n6349), .ZN(n7616) );
  INV_X1 U9271 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n7613) );
  NAND2_X1 U9272 ( .A1(n6350), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n7612) );
  NAND2_X1 U9273 ( .A1(n7635), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n7611) );
  OAI211_X1 U9274 ( .C1(n7703), .C2(n7613), .A(n7612), .B(n7611), .ZN(n7614)
         );
  INV_X1 U9275 ( .A(n7614), .ZN(n7615) );
  NAND2_X1 U9276 ( .A1(n7616), .A2(n7615), .ZN(n9532) );
  INV_X1 U9277 ( .A(n9532), .ZN(n9007) );
  NAND2_X1 U9278 ( .A1(n9640), .A2(n9007), .ZN(n9498) );
  OR2_X1 U9279 ( .A1(n9640), .A2(n9007), .ZN(n7617) );
  NAND2_X1 U9280 ( .A1(n7619), .A2(n7747), .ZN(n7621) );
  NAND2_X1 U9281 ( .A1(n7748), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7620) );
  INV_X1 U9282 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9004) );
  NAND2_X1 U9283 ( .A1(n7622), .A2(n9004), .ZN(n7623) );
  AND2_X1 U9284 ( .A1(n7632), .A2(n7623), .ZN(n9495) );
  NAND2_X1 U9285 ( .A1(n9495), .A2(n7700), .ZN(n7628) );
  INV_X1 U9286 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9390) );
  NAND2_X1 U9287 ( .A1(n6350), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n7625) );
  NAND2_X1 U9288 ( .A1(n7666), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n7624) );
  OAI211_X1 U9289 ( .C1(n9390), .C2(n7679), .A(n7625), .B(n7624), .ZN(n7626)
         );
  INV_X1 U9290 ( .A(n7626), .ZN(n7627) );
  NAND2_X1 U9291 ( .A1(n7628), .A2(n7627), .ZN(n9519) );
  INV_X1 U9292 ( .A(n9519), .ZN(n9479) );
  NAND2_X1 U9293 ( .A1(n9634), .A2(n9479), .ZN(n7936) );
  NAND2_X1 U9294 ( .A1(n7809), .A2(n7936), .ZN(n9500) );
  NAND2_X1 U9295 ( .A1(n7629), .A2(n7747), .ZN(n7631) );
  NAND2_X1 U9296 ( .A1(n7748), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7630) );
  INV_X1 U9297 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U9298 ( .A1(n7632), .A2(n9414), .ZN(n7634) );
  INV_X1 U9299 ( .A(n7645), .ZN(n7633) );
  NAND2_X1 U9300 ( .A1(n7634), .A2(n7633), .ZN(n9484) );
  OR2_X1 U9301 ( .A1(n9484), .A2(n6349), .ZN(n7641) );
  INV_X1 U9302 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n7638) );
  NAND2_X1 U9303 ( .A1(n6350), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n7637) );
  NAND2_X1 U9304 ( .A1(n7635), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7636) );
  OAI211_X1 U9305 ( .C1(n7703), .C2(n7638), .A(n7637), .B(n7636), .ZN(n7639)
         );
  INV_X1 U9306 ( .A(n7639), .ZN(n7640) );
  NAND2_X1 U9307 ( .A1(n7641), .A2(n7640), .ZN(n9502) );
  NOR2_X1 U9308 ( .A1(n9631), .A2(n9502), .ZN(n7850) );
  NAND2_X1 U9309 ( .A1(n9631), .A2(n9502), .ZN(n7849) );
  NAND2_X1 U9310 ( .A1(n7748), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7643) );
  NAND2_X1 U9311 ( .A1(n6350), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7649) );
  INV_X1 U9312 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n7644) );
  OR2_X1 U9313 ( .A1(n7703), .A2(n7644), .ZN(n7648) );
  NAND2_X1 U9314 ( .A1(n7645), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n7655) );
  OAI21_X1 U9315 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n7645), .A(n7655), .ZN(
        n9198) );
  OR2_X1 U9316 ( .A1(n6349), .A2(n9198), .ZN(n7647) );
  INV_X1 U9317 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9207) );
  OR2_X1 U9318 ( .A1(n7679), .A2(n9207), .ZN(n7646) );
  NAND4_X1 U9319 ( .A1(n7649), .A2(n7648), .A3(n7647), .A4(n7646), .ZN(n9057)
         );
  NAND2_X1 U9320 ( .A1(n7748), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7652) );
  NAND2_X1 U9321 ( .A1(n7666), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n7662) );
  INV_X1 U9322 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n7654) );
  OR2_X1 U9323 ( .A1(n7719), .A2(n7654), .ZN(n7661) );
  INV_X1 U9324 ( .A(n7655), .ZN(n7657) );
  INV_X1 U9325 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8958) );
  INV_X1 U9326 ( .A(n7668), .ZN(n7656) );
  OAI21_X1 U9327 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n7657), .A(n7656), .ZN(
        n9179) );
  OR2_X1 U9328 ( .A1(n6349), .A2(n9179), .ZN(n7660) );
  INV_X1 U9329 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n7658) );
  OR2_X1 U9330 ( .A1(n7679), .A2(n7658), .ZN(n7659) );
  NAND4_X1 U9331 ( .A1(n7662), .A2(n7661), .A3(n7660), .A4(n7659), .ZN(n9196)
         );
  OR2_X2 U9332 ( .A1(n9619), .A2(n9032), .ZN(n7946) );
  NAND2_X1 U9333 ( .A1(n9619), .A2(n9032), .ZN(n7825) );
  INV_X1 U9334 ( .A(n9619), .ZN(n9182) );
  NAND2_X1 U9335 ( .A1(n7748), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7664) );
  NAND2_X1 U9336 ( .A1(n7666), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n7673) );
  INV_X1 U9337 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n7667) );
  OR2_X1 U9338 ( .A1(n7719), .A2(n7667), .ZN(n7672) );
  NAND2_X1 U9339 ( .A1(n7668), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n7677) );
  OAI21_X1 U9340 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n7668), .A(n7677), .ZN(
        n9166) );
  OR2_X1 U9341 ( .A1(n6349), .A2(n9166), .ZN(n7671) );
  INV_X1 U9342 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n7669) );
  OR2_X1 U9343 ( .A1(n7679), .A2(n7669), .ZN(n7670) );
  NAND4_X1 U9344 ( .A1(n7673), .A2(n7672), .A3(n7671), .A4(n7670), .ZN(n9056)
         );
  INV_X1 U9345 ( .A(n9056), .ZN(n9186) );
  NAND2_X1 U9346 ( .A1(n9169), .A2(n9186), .ZN(n7674) );
  NAND2_X1 U9347 ( .A1(n7748), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7676) );
  INV_X1 U9348 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9454) );
  OR2_X1 U9349 ( .A1(n7719), .A2(n9454), .ZN(n7683) );
  INV_X1 U9350 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9326) );
  OR2_X1 U9351 ( .A1(n7703), .A2(n9326), .ZN(n7682) );
  INV_X1 U9352 ( .A(n7677), .ZN(n7678) );
  NAND2_X1 U9353 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n7678), .ZN(n7689) );
  OAI21_X1 U9354 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(n7678), .A(n7689), .ZN(
        n9149) );
  OR2_X1 U9355 ( .A1(n6349), .A2(n9149), .ZN(n7681) );
  INV_X1 U9356 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9422) );
  OR2_X1 U9357 ( .A1(n7679), .A2(n9422), .ZN(n7680) );
  NAND4_X1 U9358 ( .A1(n7683), .A2(n7682), .A3(n7681), .A4(n7680), .ZN(n9172)
         );
  NAND2_X1 U9359 ( .A1(n9609), .A2(n9031), .ZN(n7907) );
  NOR2_X1 U9360 ( .A1(n9609), .A2(n9172), .ZN(n7684) );
  AOI21_X1 U9361 ( .B1(n9147), .B2(n9155), .A(n7684), .ZN(n9133) );
  NAND2_X1 U9362 ( .A1(n7748), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n7685) );
  NAND2_X1 U9363 ( .A1(n6350), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7694) );
  INV_X1 U9364 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7687) );
  OR2_X1 U9365 ( .A1(n7703), .A2(n7687), .ZN(n7693) );
  INV_X1 U9366 ( .A(n7689), .ZN(n7688) );
  NAND2_X1 U9367 ( .A1(n7688), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n7730) );
  INV_X1 U9368 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8928) );
  NAND2_X1 U9369 ( .A1(n7689), .A2(n8928), .ZN(n7690) );
  NAND2_X1 U9370 ( .A1(n7730), .A2(n7690), .ZN(n9139) );
  OR2_X1 U9371 ( .A1(n6349), .A2(n9139), .ZN(n7692) );
  INV_X1 U9372 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9142) );
  OR2_X1 U9373 ( .A1(n7679), .A2(n9142), .ZN(n7691) );
  NAND2_X1 U9374 ( .A1(n9603), .A2(n9156), .ZN(n7910) );
  NAND2_X1 U9375 ( .A1(n9133), .A2(n9136), .ZN(n9132) );
  INV_X1 U9376 ( .A(n9603), .ZN(n9143) );
  NAND2_X1 U9377 ( .A1(n9603), .A2(n7695), .ZN(n7696) );
  NAND2_X1 U9378 ( .A1(n9132), .A2(n7696), .ZN(n7708) );
  NAND2_X1 U9379 ( .A1(n8760), .A2(n7747), .ZN(n7698) );
  NAND2_X1 U9380 ( .A1(n7748), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7697) );
  INV_X1 U9381 ( .A(n7730), .ZN(n7699) );
  NAND2_X1 U9382 ( .A1(n7700), .A2(n7699), .ZN(n7707) );
  INV_X1 U9383 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7701) );
  OR2_X1 U9384 ( .A1(n7719), .A2(n7701), .ZN(n7706) );
  INV_X1 U9385 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7702) );
  OR2_X1 U9386 ( .A1(n7703), .A2(n7702), .ZN(n7705) );
  INV_X1 U9387 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n7731) );
  OR2_X1 U9388 ( .A1(n7679), .A2(n7731), .ZN(n7704) );
  NAND2_X1 U9389 ( .A1(n9598), .A2(n9134), .ZN(n7979) );
  AND2_X1 U9390 ( .A1(n7790), .A2(n7709), .ZN(n7902) );
  NAND2_X1 U9391 ( .A1(n7710), .A2(n7902), .ZN(n9587) );
  OR2_X1 U9392 ( .A1(n9659), .A2(n9019), .ZN(n9564) );
  NAND2_X1 U9393 ( .A1(n9659), .A2(n9019), .ZN(n7793) );
  INV_X1 U9394 ( .A(n9557), .ZN(n9566) );
  NAND3_X1 U9395 ( .A1(n9584), .A2(n9566), .A3(n9564), .ZN(n9565) );
  NAND2_X1 U9396 ( .A1(n9565), .A2(n7932), .ZN(n9538) );
  NOR2_X1 U9397 ( .A1(n9651), .A2(n8994), .ZN(n7935) );
  NOR2_X1 U9398 ( .A1(n7935), .A2(n7913), .ZN(n7852) );
  XNOR2_X1 U9399 ( .A(n9644), .B(n9518), .ZN(n9531) );
  NOR2_X1 U9400 ( .A1(n9644), .A2(n9545), .ZN(n7808) );
  INV_X1 U9401 ( .A(n9506), .ZN(n9517) );
  AND2_X1 U9402 ( .A1(n7936), .A2(n9498), .ZN(n7917) );
  INV_X1 U9403 ( .A(n7809), .ZN(n7711) );
  INV_X1 U9404 ( .A(n9631), .ZN(n9488) );
  NAND2_X1 U9405 ( .A1(n9488), .A2(n9502), .ZN(n7815) );
  INV_X1 U9406 ( .A(n9502), .ZN(n9005) );
  AND2_X1 U9407 ( .A1(n9631), .A2(n9005), .ZN(n7819) );
  XNOR2_X1 U9408 ( .A(n9201), .B(n9481), .ZN(n9194) );
  NAND2_X1 U9409 ( .A1(n9201), .A2(n9481), .ZN(n7821) );
  INV_X1 U9410 ( .A(n7946), .ZN(n7712) );
  NAND2_X1 U9411 ( .A1(n9614), .A2(n9186), .ZN(n7906) );
  INV_X1 U9412 ( .A(n7948), .ZN(n7713) );
  INV_X1 U9413 ( .A(n7943), .ZN(n7714) );
  NAND2_X1 U9414 ( .A1(n7695), .A2(n9913), .ZN(n7725) );
  INV_X1 U9415 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n7716) );
  NOR2_X1 U9416 ( .A1(n7703), .A2(n7716), .ZN(n7722) );
  INV_X1 U9417 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n7717) );
  NOR2_X1 U9418 ( .A1(n7679), .A2(n7717), .ZN(n7721) );
  INV_X1 U9419 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n7718) );
  NOR2_X1 U9420 ( .A1(n7719), .A2(n7718), .ZN(n7720) );
  OR3_X1 U9421 ( .A1(n7722), .A2(n7721), .A3(n7720), .ZN(n9054) );
  NAND2_X1 U9422 ( .A1(n9802), .A2(P1_B_REG_SCAN_IN), .ZN(n7723) );
  AND2_X1 U9423 ( .A1(n9911), .A2(n7723), .ZN(n8003) );
  NAND2_X1 U9424 ( .A1(n9054), .A2(n8003), .ZN(n7724) );
  INV_X1 U9425 ( .A(n9601), .ZN(n7728) );
  NAND2_X1 U9426 ( .A1(n7728), .A2(n9926), .ZN(n7735) );
  OR2_X2 U9427 ( .A1(n9578), .A2(n9659), .ZN(n9576) );
  AND2_X2 U9428 ( .A1(n9547), .A2(n9530), .ZN(n9525) );
  INV_X1 U9429 ( .A(n9640), .ZN(n9514) );
  NAND2_X2 U9430 ( .A1(n9525), .A2(n9514), .ZN(n9508) );
  NAND2_X1 U9431 ( .A1(n9494), .A2(n9488), .ZN(n9193) );
  NAND2_X1 U9432 ( .A1(n9169), .A2(n9178), .ZN(n9163) );
  INV_X1 U9433 ( .A(n9141), .ZN(n7729) );
  INV_X1 U9434 ( .A(n9598), .ZN(n7750) );
  AND2_X2 U9435 ( .A1(n7750), .A2(n9141), .ZN(n9127) );
  NOR2_X1 U9436 ( .A1(n7750), .A2(n9930), .ZN(n7733) );
  OAI22_X1 U9437 ( .A1(n9926), .A2(n7731), .B1(n7730), .B2(n9936), .ZN(n7732)
         );
  OAI211_X1 U9438 ( .C1(n9597), .C2(n9602), .A(n7735), .B(n7734), .ZN(P1_U3355) );
  NAND2_X1 U9439 ( .A1(n8014), .A2(n7747), .ZN(n7737) );
  NAND2_X1 U9440 ( .A1(n7748), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7736) );
  INV_X1 U9441 ( .A(n9054), .ZN(n7880) );
  NAND2_X1 U9442 ( .A1(n7740), .A2(n7739), .ZN(n7741) );
  NAND2_X1 U9443 ( .A1(n7742), .A2(n7741), .ZN(n7746) );
  MUX2_X1 U9444 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7743), .Z(n7744) );
  XNOR2_X1 U9445 ( .A(n7744), .B(SI_31_), .ZN(n7745) );
  NAND2_X1 U9446 ( .A1(n7748), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7749) );
  INV_X1 U9447 ( .A(n9134), .ZN(n9055) );
  NOR3_X1 U9448 ( .A1(n7838), .A2(n9598), .A3(n9055), .ZN(n7834) );
  INV_X1 U9449 ( .A(n9659), .ZN(n9582) );
  NAND2_X1 U9450 ( .A1(n8774), .A2(n9042), .ZN(n7897) );
  NAND2_X1 U9451 ( .A1(n7897), .A2(n7778), .ZN(n7918) );
  NAND2_X1 U9452 ( .A1(n7918), .A2(n7781), .ZN(n7782) );
  NAND2_X1 U9453 ( .A1(n7754), .A2(n7753), .ZN(n7763) );
  NAND3_X1 U9454 ( .A1(n7763), .A2(n7755), .A3(n7905), .ZN(n7756) );
  AND2_X1 U9455 ( .A1(n7768), .A2(n7764), .ZN(n7920) );
  NAND2_X1 U9456 ( .A1(n7756), .A2(n7920), .ZN(n7760) );
  INV_X1 U9457 ( .A(n7765), .ZN(n7757) );
  NOR2_X1 U9458 ( .A1(n7770), .A2(n7757), .ZN(n7892) );
  NAND2_X1 U9459 ( .A1(n7759), .A2(n7758), .ZN(n7769) );
  INV_X1 U9460 ( .A(n7769), .ZN(n7885) );
  AOI21_X1 U9461 ( .B1(n7760), .B2(n7892), .A(n7885), .ZN(n7772) );
  INV_X1 U9462 ( .A(n7905), .ZN(n7761) );
  AOI21_X1 U9463 ( .B1(n7763), .B2(n7762), .A(n7761), .ZN(n7767) );
  INV_X1 U9464 ( .A(n7764), .ZN(n7766) );
  AND2_X1 U9465 ( .A1(n7769), .A2(n7768), .ZN(n7771) );
  MUX2_X1 U9466 ( .A(n7887), .B(n7891), .S(n4699), .Z(n7773) );
  INV_X1 U9467 ( .A(n7866), .ZN(n7774) );
  NAND2_X1 U9468 ( .A1(n7775), .A2(n7774), .ZN(n7784) );
  NAND2_X1 U9469 ( .A1(n7777), .A2(n7776), .ZN(n7888) );
  INV_X1 U9470 ( .A(n7778), .ZN(n7896) );
  NOR2_X1 U9471 ( .A1(n7893), .A2(n7835), .ZN(n7783) );
  OAI211_X1 U9472 ( .C1(n7784), .C2(n4678), .A(n4468), .B(n7783), .ZN(n7785)
         );
  NAND3_X1 U9473 ( .A1(n7787), .A2(n7786), .A3(n7785), .ZN(n7789) );
  AND2_X1 U9474 ( .A1(n9586), .A2(n7923), .ZN(n7899) );
  MUX2_X1 U9475 ( .A(n7902), .B(n7899), .S(n7835), .Z(n7788) );
  NAND2_X1 U9476 ( .A1(n7789), .A2(n7788), .ZN(n7792) );
  MUX2_X1 U9477 ( .A(n9586), .B(n7790), .S(n7835), .Z(n7791) );
  NAND2_X1 U9478 ( .A1(n7792), .A2(n7791), .ZN(n7797) );
  INV_X1 U9479 ( .A(n7797), .ZN(n7798) );
  NAND2_X1 U9480 ( .A1(n7802), .A2(n9564), .ZN(n7933) );
  NAND2_X1 U9481 ( .A1(n7932), .A2(n7793), .ZN(n7928) );
  INV_X1 U9482 ( .A(n7928), .ZN(n7796) );
  OAI21_X1 U9483 ( .B1(n7928), .B2(n9019), .A(n7835), .ZN(n7794) );
  AOI22_X1 U9484 ( .A1(n7797), .A2(n7796), .B1(n7795), .B2(n7794), .ZN(n7805)
         );
  AOI211_X1 U9485 ( .C1(n9582), .C2(n7798), .A(n7933), .B(n7805), .ZN(n7800)
         );
  INV_X1 U9486 ( .A(n7932), .ZN(n7799) );
  NOR3_X1 U9487 ( .A1(n7800), .A2(n7799), .A3(n7913), .ZN(n7801) );
  INV_X1 U9488 ( .A(n7802), .ZN(n7803) );
  NOR2_X1 U9489 ( .A1(n7935), .A2(n7803), .ZN(n7804) );
  AOI21_X1 U9490 ( .B1(n7805), .B2(n7804), .A(n7913), .ZN(n7806) );
  AND2_X1 U9491 ( .A1(n9644), .A2(n9545), .ZN(n7912) );
  INV_X1 U9492 ( .A(n7917), .ZN(n7807) );
  AOI21_X1 U9493 ( .B1(n7912), .B2(n9517), .A(n7807), .ZN(n7811) );
  OAI21_X1 U9494 ( .B1(n9506), .B2(n7808), .A(n9498), .ZN(n7810) );
  AND2_X1 U9495 ( .A1(n7810), .A2(n7809), .ZN(n7938) );
  MUX2_X1 U9496 ( .A(n7811), .B(n7938), .S(n7835), .Z(n7814) );
  INV_X1 U9497 ( .A(n9634), .ZN(n9497) );
  MUX2_X1 U9498 ( .A(n9497), .B(n9479), .S(n7835), .Z(n7812) );
  INV_X1 U9499 ( .A(n7821), .ZN(n7816) );
  OR2_X1 U9500 ( .A1(n9201), .A2(n9481), .ZN(n7820) );
  NAND2_X1 U9501 ( .A1(n7820), .A2(n7815), .ZN(n7942) );
  NOR4_X1 U9502 ( .A1(n7817), .A2(n7816), .A3(n7819), .A4(n7942), .ZN(n7828)
         );
  NAND2_X1 U9503 ( .A1(n7942), .A2(n7821), .ZN(n7818) );
  NAND2_X1 U9504 ( .A1(n7946), .A2(n7818), .ZN(n7824) );
  NAND2_X1 U9505 ( .A1(n7820), .A2(n7819), .ZN(n7822) );
  AND2_X1 U9506 ( .A1(n7822), .A2(n7821), .ZN(n7823) );
  NAND2_X1 U9507 ( .A1(n7823), .A2(n7825), .ZN(n7911) );
  MUX2_X1 U9508 ( .A(n7825), .B(n7946), .S(n7835), .Z(n7826) );
  OR2_X1 U9509 ( .A1(n9614), .A2(n9186), .ZN(n7947) );
  MUX2_X1 U9510 ( .A(n7947), .B(n7906), .S(n7835), .Z(n7829) );
  INV_X1 U9511 ( .A(n9136), .ZN(n7875) );
  MUX2_X1 U9512 ( .A(n7948), .B(n7907), .S(n7835), .Z(n7830) );
  MUX2_X1 U9513 ( .A(n7910), .B(n7943), .S(n7835), .Z(n7831) );
  NAND2_X1 U9514 ( .A1(n8004), .A2(n9054), .ZN(n7832) );
  NAND2_X1 U9515 ( .A1(n9128), .A2(n7832), .ZN(n7955) );
  NAND2_X1 U9516 ( .A1(n7838), .A2(n7835), .ZN(n7843) );
  NAND2_X1 U9517 ( .A1(n4943), .A2(n4936), .ZN(n7986) );
  INV_X1 U9518 ( .A(n7955), .ZN(n7837) );
  NAND3_X1 U9519 ( .A1(n7986), .A2(n7837), .A3(n4699), .ZN(n7842) );
  INV_X1 U9520 ( .A(n7838), .ZN(n7959) );
  NAND3_X1 U9521 ( .A1(n9598), .A2(n9134), .A3(n4699), .ZN(n7839) );
  OAI21_X1 U9522 ( .B1(n7944), .B2(n4699), .A(n7839), .ZN(n7840) );
  NAND3_X1 U9523 ( .A1(n7959), .A2(n7955), .A3(n7840), .ZN(n7841) );
  NAND2_X1 U9524 ( .A1(n7844), .A2(n7883), .ZN(n7847) );
  NOR2_X1 U9525 ( .A1(n4943), .A2(n4936), .ZN(n7957) );
  AOI21_X1 U9526 ( .B1(n9203), .B2(n7845), .A(n7848), .ZN(n7846) );
  AOI211_X1 U9527 ( .C1(n7848), .C2(n7847), .A(n7957), .B(n7846), .ZN(n7963)
         );
  INV_X1 U9528 ( .A(n7986), .ZN(n7879) );
  INV_X1 U9529 ( .A(n7982), .ZN(n7878) );
  INV_X1 U9530 ( .A(n7849), .ZN(n7851) );
  OR2_X1 U9531 ( .A1(n7851), .A2(n7850), .ZN(n9478) );
  INV_X1 U9532 ( .A(n7852), .ZN(n9540) );
  INV_X1 U9533 ( .A(n6798), .ZN(n7853) );
  NAND4_X1 U9534 ( .A1(n6729), .A2(n7855), .A3(n7854), .A4(n7853), .ZN(n7859)
         );
  NOR4_X1 U9535 ( .A1(n7859), .A2(n7858), .A3(n7857), .A4(n7856), .ZN(n7861)
         );
  NAND4_X1 U9536 ( .A1(n7863), .A2(n7862), .A3(n7861), .A4(n7860), .ZN(n7864)
         );
  NOR4_X1 U9537 ( .A1(n7867), .A2(n7866), .A3(n7865), .A4(n7864), .ZN(n7869)
         );
  NAND4_X1 U9538 ( .A1(n9585), .A2(n7870), .A3(n7869), .A4(n7868), .ZN(n7871)
         );
  NOR4_X1 U9539 ( .A1(n9506), .A2(n9540), .A3(n9557), .A4(n7871), .ZN(n7872)
         );
  NAND3_X1 U9540 ( .A1(n9478), .A2(n7872), .A3(n9531), .ZN(n7873) );
  NOR4_X1 U9541 ( .A1(n9185), .A2(n9194), .A3(n9500), .A4(n7873), .ZN(n7874)
         );
  NAND4_X1 U9542 ( .A1(n7875), .A2(n4694), .A3(n7874), .A4(n9171), .ZN(n7876)
         );
  NOR4_X1 U9543 ( .A1(n7879), .A2(n7878), .A3(n7877), .A4(n7876), .ZN(n7884)
         );
  INV_X1 U9544 ( .A(n7957), .ZN(n7882) );
  NAND2_X1 U9545 ( .A1(n9128), .A2(n7880), .ZN(n7881) );
  AND2_X1 U9546 ( .A1(n7882), .A2(n7881), .ZN(n7964) );
  AOI21_X1 U9547 ( .B1(n7884), .B2(n7964), .A(n7883), .ZN(n7961) );
  INV_X1 U9548 ( .A(n9586), .ZN(n7901) );
  NAND2_X1 U9549 ( .A1(n7891), .A2(n7885), .ZN(n7886) );
  AND3_X1 U9550 ( .A1(n7888), .A2(n7887), .A3(n7886), .ZN(n7889) );
  AND2_X1 U9551 ( .A1(n7890), .A2(n7889), .ZN(n7919) );
  NAND2_X1 U9552 ( .A1(n7892), .A2(n7891), .ZN(n7894) );
  AOI21_X1 U9553 ( .B1(n7919), .B2(n7894), .A(n7893), .ZN(n7895) );
  OAI21_X1 U9554 ( .B1(n7896), .B2(n7895), .A(n4468), .ZN(n7898) );
  NAND3_X1 U9555 ( .A1(n7899), .A2(n7898), .A3(n7897), .ZN(n7900) );
  OAI21_X1 U9556 ( .B1(n7902), .B2(n7901), .A(n7900), .ZN(n7903) );
  INV_X1 U9557 ( .A(n7903), .ZN(n7904) );
  OR2_X1 U9558 ( .A1(n7928), .A2(n7904), .ZN(n7926) );
  AND2_X1 U9559 ( .A1(n7926), .A2(n7905), .ZN(n7965) );
  NAND2_X1 U9560 ( .A1(n7907), .A2(n7906), .ZN(n7908) );
  NAND2_X1 U9561 ( .A1(n7908), .A2(n7948), .ZN(n7909) );
  NAND2_X1 U9562 ( .A1(n7910), .A2(n7909), .ZN(n7945) );
  INV_X1 U9563 ( .A(n7912), .ZN(n7915) );
  INV_X1 U9564 ( .A(n7913), .ZN(n7914) );
  AND2_X1 U9565 ( .A1(n7915), .A2(n7914), .ZN(n7916) );
  AND2_X1 U9566 ( .A1(n7917), .A2(n7916), .ZN(n7931) );
  INV_X1 U9567 ( .A(n7918), .ZN(n7925) );
  INV_X1 U9568 ( .A(n7919), .ZN(n7922) );
  INV_X1 U9569 ( .A(n7920), .ZN(n7921) );
  NOR2_X1 U9570 ( .A1(n7922), .A2(n7921), .ZN(n7924) );
  NAND4_X1 U9571 ( .A1(n9586), .A2(n7925), .A3(n7924), .A4(n7923), .ZN(n7927)
         );
  OAI21_X1 U9572 ( .B1(n7928), .B2(n7927), .A(n7926), .ZN(n7929) );
  NAND2_X1 U9573 ( .A1(n7931), .A2(n7929), .ZN(n7930) );
  AOI21_X1 U9574 ( .B1(n7965), .B2(n7974), .A(n7978), .ZN(n7956) );
  INV_X1 U9575 ( .A(n7931), .ZN(n7940) );
  AND2_X1 U9576 ( .A1(n7933), .A2(n7932), .ZN(n7934) );
  NOR2_X1 U9577 ( .A1(n7935), .A2(n7934), .ZN(n7939) );
  INV_X1 U9578 ( .A(n7936), .ZN(n7937) );
  OAI22_X1 U9579 ( .A1(n7940), .A2(n7939), .B1(n7938), .B2(n7937), .ZN(n7941)
         );
  NOR2_X1 U9580 ( .A1(n7942), .A2(n7941), .ZN(n7953) );
  AND2_X1 U9581 ( .A1(n7944), .A2(n7943), .ZN(n7952) );
  INV_X1 U9582 ( .A(n7945), .ZN(n7950) );
  NAND3_X1 U9583 ( .A1(n7948), .A2(n7947), .A3(n7946), .ZN(n7949) );
  NAND2_X1 U9584 ( .A1(n7950), .A2(n7949), .ZN(n7951) );
  OAI211_X1 U9585 ( .C1(n7954), .C2(n7953), .A(n7952), .B(n7951), .ZN(n7980)
         );
  OAI211_X1 U9586 ( .C1(n7956), .C2(n7980), .A(n7979), .B(n7955), .ZN(n7958)
         );
  AOI211_X1 U9587 ( .C1(n7959), .C2(n7958), .A(n7967), .B(n7957), .ZN(n7960)
         );
  INV_X1 U9588 ( .A(n7964), .ZN(n7985) );
  INV_X1 U9589 ( .A(n7965), .ZN(n7976) );
  INV_X1 U9590 ( .A(n7966), .ZN(n7970) );
  AOI21_X1 U9591 ( .B1(n6727), .B2(n6725), .A(n7967), .ZN(n7969) );
  NAND3_X1 U9592 ( .A1(n7970), .A2(n7969), .A3(n7968), .ZN(n7971) );
  NOR2_X1 U9593 ( .A1(n7972), .A2(n7971), .ZN(n7973) );
  NOR2_X1 U9594 ( .A1(n7974), .A2(n7973), .ZN(n7975) );
  NOR2_X1 U9595 ( .A1(n7976), .A2(n7975), .ZN(n7977) );
  NOR2_X1 U9596 ( .A1(n7978), .A2(n7977), .ZN(n7981) );
  OAI21_X1 U9597 ( .B1(n7981), .B2(n7980), .A(n7979), .ZN(n7983) );
  AND2_X1 U9598 ( .A1(n7983), .A2(n7982), .ZN(n7984) );
  NAND2_X1 U9599 ( .A1(n7987), .A2(n7986), .ZN(n7989) );
  NOR2_X1 U9600 ( .A1(n7989), .A2(n9124), .ZN(n7988) );
  INV_X1 U9601 ( .A(n7989), .ZN(n7990) );
  OAI21_X1 U9602 ( .B1(n7990), .B2(n7992), .A(n7991), .ZN(n7998) );
  INV_X1 U9603 ( .A(n7991), .ZN(n7995) );
  INV_X1 U9604 ( .A(n7992), .ZN(n7993) );
  NAND4_X1 U9605 ( .A1(n9913), .A2(n9691), .A3(n9802), .A4(n7993), .ZN(n7994)
         );
  OAI211_X1 U9606 ( .C1(n7996), .C2(n7995), .A(n7994), .B(P1_B_REG_SCAN_IN), 
        .ZN(n7997) );
  OAI21_X1 U9607 ( .B1(n7999), .B2(n7998), .A(n7997), .ZN(P1_U3240) );
  INV_X1 U9608 ( .A(n8016), .ZN(n8759) );
  INV_X1 U9609 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9240) );
  NAND3_X1 U9610 ( .A1(P1_STATE_REG_SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        n9240), .ZN(n8000) );
  OAI222_X1 U9611 ( .A1(n9698), .A2(n9459), .B1(n9695), .B2(n8759), .C1(n8001), 
        .C2(n8000), .ZN(P1_U3322) );
  NAND2_X1 U9612 ( .A1(n9763), .A2(n9127), .ZN(n8002) );
  XNOR2_X1 U9613 ( .A(n7836), .B(n8002), .ZN(n9754) );
  NAND2_X1 U9614 ( .A1(n9754), .A2(n9909), .ZN(n8006) );
  NAND2_X1 U9615 ( .A1(n8004), .A2(n8003), .ZN(n9762) );
  NOR2_X1 U9616 ( .A1(n4382), .A2(n9762), .ZN(n9129) );
  AOI21_X1 U9617 ( .B1(n4382), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9129), .ZN(
        n8005) );
  OAI211_X1 U9618 ( .C1(n7836), .C2(n9930), .A(n8006), .B(n8005), .ZN(P1_U3261) );
  OAI222_X1 U9619 ( .A1(n8009), .A2(n8008), .B1(n6177), .B2(P1_U3084), .C1(
        n8007), .C2(n9698), .ZN(P1_U3333) );
  INV_X1 U9620 ( .A(n8010), .ZN(n9702) );
  OAI222_X1 U9621 ( .A1(n5639), .A2(n4374), .B1(n4385), .B2(n9702), .C1(n8011), 
        .C2(n8761), .ZN(P2_U3330) );
  INV_X1 U9622 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9242) );
  NOR2_X1 U9623 ( .A1(n5569), .A2(n9242), .ZN(n8013) );
  INV_X1 U9624 ( .A(n8425), .ZN(n9759) );
  NAND2_X1 U9625 ( .A1(n8016), .A2(n8015), .ZN(n8018) );
  OR2_X1 U9626 ( .A1(n5569), .A2(n6116), .ZN(n8017) );
  INV_X1 U9627 ( .A(n8420), .ZN(n8020) );
  INV_X1 U9628 ( .A(n8340), .ZN(n8019) );
  NAND2_X1 U9629 ( .A1(n9759), .A2(n8019), .ZN(n8170) );
  XNOR2_X1 U9630 ( .A(n8021), .B(n8615), .ZN(n8223) );
  NAND2_X1 U9631 ( .A1(n8023), .A2(n8022), .ZN(n8222) );
  NAND2_X1 U9632 ( .A1(n8175), .A2(n4455), .ZN(n8213) );
  NOR2_X2 U9633 ( .A1(n8025), .A2(n8024), .ZN(n8166) );
  MUX2_X1 U9634 ( .A(n8213), .B(n8214), .S(n8166), .Z(n8172) );
  MUX2_X1 U9635 ( .A(n4400), .B(n8026), .S(n8166), .Z(n8169) );
  AND2_X1 U9636 ( .A1(n8069), .A2(n8027), .ZN(n8066) );
  AND2_X1 U9637 ( .A1(n8028), .A2(n8052), .ZN(n8183) );
  INV_X1 U9638 ( .A(n8183), .ZN(n8030) );
  NAND2_X1 U9639 ( .A1(n8033), .A2(n8029), .ZN(n8188) );
  MUX2_X1 U9640 ( .A(n8030), .B(n8188), .S(n8166), .Z(n8053) );
  NOR2_X1 U9641 ( .A1(n8188), .A2(n8031), .ZN(n8032) );
  AOI21_X1 U9642 ( .B1(n8053), .B2(n8033), .A(n8032), .ZN(n8035) );
  OAI21_X1 U9643 ( .B1(n8035), .B2(n8034), .A(n8173), .ZN(n8041) );
  INV_X1 U9644 ( .A(n8053), .ZN(n8039) );
  AND2_X1 U9645 ( .A1(n8231), .A2(n8216), .ZN(n8042) );
  OAI211_X1 U9646 ( .C1(n8036), .C2(n8042), .A(n8047), .B(n5615), .ZN(n8037)
         );
  NAND3_X1 U9647 ( .A1(n8037), .A2(n8044), .A3(n8173), .ZN(n8038) );
  NAND3_X1 U9648 ( .A1(n8039), .A2(n8184), .A3(n8038), .ZN(n8040) );
  NAND2_X1 U9649 ( .A1(n8041), .A2(n8040), .ZN(n8050) );
  INV_X1 U9650 ( .A(n8042), .ZN(n8046) );
  INV_X1 U9651 ( .A(n5615), .ZN(n8045) );
  OAI211_X1 U9652 ( .C1(n8046), .C2(n8045), .A(n8044), .B(n8043), .ZN(n8048)
         );
  NAND3_X1 U9653 ( .A1(n8048), .A2(n8166), .A3(n8047), .ZN(n8049) );
  NAND2_X1 U9654 ( .A1(n8050), .A2(n8049), .ZN(n8057) );
  AOI22_X1 U9655 ( .A1(n8053), .A2(n8052), .B1(n8183), .B2(n8051), .ZN(n8055)
         );
  INV_X1 U9656 ( .A(n8058), .ZN(n8054) );
  OAI21_X1 U9657 ( .B1(n8055), .B2(n8054), .A(n8166), .ZN(n8056) );
  MUX2_X1 U9658 ( .A(n8059), .B(n8058), .S(n8173), .Z(n8061) );
  INV_X1 U9659 ( .A(n8060), .ZN(n8190) );
  AND2_X1 U9660 ( .A1(n8061), .A2(n8190), .ZN(n8062) );
  INV_X1 U9661 ( .A(n8063), .ZN(n8064) );
  NAND2_X1 U9662 ( .A1(n8068), .A2(n8067), .ZN(n8072) );
  AND2_X1 U9663 ( .A1(n8077), .A2(n8069), .ZN(n8071) );
  MUX2_X1 U9664 ( .A(n8071), .B(n8070), .S(n8173), .Z(n8075) );
  NAND2_X1 U9665 ( .A1(n8072), .A2(n8075), .ZN(n8083) );
  NAND2_X1 U9666 ( .A1(n8084), .A2(n8073), .ZN(n8080) );
  NAND4_X1 U9667 ( .A1(n8076), .A2(n5310), .A3(n8075), .A4(n8074), .ZN(n8078)
         );
  NAND3_X1 U9668 ( .A1(n8078), .A2(n8087), .A3(n8077), .ZN(n8079) );
  MUX2_X1 U9669 ( .A(n8080), .B(n8079), .S(n8173), .Z(n8081) );
  INV_X1 U9670 ( .A(n8081), .ZN(n8082) );
  NAND2_X1 U9671 ( .A1(n8083), .A2(n8082), .ZN(n8092) );
  AND2_X1 U9672 ( .A1(n8089), .A2(n8084), .ZN(n8086) );
  AOI21_X1 U9673 ( .B1(n8092), .B2(n8086), .A(n8085), .ZN(n8094) );
  AND2_X1 U9674 ( .A1(n8088), .A2(n8087), .ZN(n8091) );
  INV_X1 U9675 ( .A(n8089), .ZN(n8090) );
  AOI21_X1 U9676 ( .B1(n8092), .B2(n8091), .A(n8090), .ZN(n8093) );
  MUX2_X1 U9677 ( .A(n8094), .B(n8093), .S(n8166), .Z(n8102) );
  INV_X1 U9678 ( .A(n8095), .ZN(n8098) );
  INV_X1 U9679 ( .A(n8096), .ZN(n8097) );
  MUX2_X1 U9680 ( .A(n8098), .B(n8097), .S(n8173), .Z(n8099) );
  NOR2_X1 U9681 ( .A1(n8200), .A2(n8099), .ZN(n8100) );
  OAI21_X1 U9682 ( .B1(n8102), .B2(n8101), .A(n8100), .ZN(n8107) );
  NAND2_X1 U9683 ( .A1(n8346), .A2(n8166), .ZN(n8105) );
  NAND2_X1 U9684 ( .A1(n8103), .A2(n8173), .ZN(n8104) );
  MUX2_X1 U9685 ( .A(n8105), .B(n8104), .S(n8723), .Z(n8106) );
  NAND3_X1 U9686 ( .A1(n8107), .A2(n4727), .A3(n8106), .ZN(n8112) );
  MUX2_X1 U9687 ( .A(n4796), .B(n8109), .S(n8173), .Z(n8110) );
  NOR2_X1 U9688 ( .A1(n5430), .A2(n8110), .ZN(n8111) );
  NAND2_X1 U9689 ( .A1(n8112), .A2(n8111), .ZN(n8117) );
  MUX2_X1 U9690 ( .A(n8114), .B(n4792), .S(n8166), .Z(n8115) );
  NOR2_X1 U9691 ( .A1(n5448), .A2(n8115), .ZN(n8116) );
  INV_X1 U9692 ( .A(n8118), .ZN(n8181) );
  NAND2_X1 U9693 ( .A1(n8181), .A2(n8119), .ZN(n8122) );
  INV_X1 U9694 ( .A(n8120), .ZN(n8121) );
  MUX2_X1 U9695 ( .A(n8122), .B(n8121), .S(n8166), .Z(n8123) );
  INV_X1 U9696 ( .A(n8123), .ZN(n8124) );
  NAND2_X1 U9697 ( .A1(n8125), .A2(n8180), .ZN(n8132) );
  NAND2_X1 U9698 ( .A1(n8139), .A2(n8133), .ZN(n8126) );
  AND2_X1 U9699 ( .A1(n8131), .A2(n8138), .ZN(n8128) );
  INV_X1 U9700 ( .A(n8143), .ZN(n8127) );
  AOI21_X1 U9701 ( .B1(n8129), .B2(n8128), .A(n8127), .ZN(n8130) );
  INV_X1 U9702 ( .A(n8524), .ZN(n8206) );
  INV_X1 U9703 ( .A(n8132), .ZN(n8135) );
  INV_X1 U9704 ( .A(n8133), .ZN(n8134) );
  AOI21_X1 U9705 ( .B1(n8136), .B2(n8135), .A(n8134), .ZN(n8141) );
  INV_X1 U9706 ( .A(n8137), .ZN(n8140) );
  OAI211_X1 U9707 ( .C1(n8141), .C2(n8140), .A(n8139), .B(n8138), .ZN(n8144)
         );
  NAND4_X1 U9708 ( .A1(n8144), .A2(n8143), .A3(n8142), .A4(n8173), .ZN(n8145)
         );
  AOI21_X1 U9709 ( .B1(n8150), .B2(n8148), .A(n8173), .ZN(n8149) );
  NAND3_X1 U9710 ( .A1(n8669), .A2(n4491), .A3(n8166), .ZN(n8151) );
  NAND2_X1 U9711 ( .A1(n8491), .A2(n8151), .ZN(n8155) );
  INV_X1 U9712 ( .A(n8152), .ZN(n8161) );
  INV_X1 U9713 ( .A(n8468), .ZN(n8153) );
  NAND2_X1 U9714 ( .A1(n8153), .A2(n8166), .ZN(n8154) );
  OAI211_X1 U9715 ( .C1(n8156), .C2(n8155), .A(n8161), .B(n8154), .ZN(n8160)
         );
  AOI21_X1 U9716 ( .B1(n8159), .B2(n8157), .A(n8166), .ZN(n8158) );
  OAI21_X1 U9717 ( .B1(n8166), .B2(n8161), .A(n8456), .ZN(n8165) );
  NAND2_X1 U9718 ( .A1(n8341), .A2(n8166), .ZN(n8163) );
  NAND2_X1 U9719 ( .A1(n8441), .A2(n8173), .ZN(n8162) );
  MUX2_X1 U9720 ( .A(n8163), .B(n8162), .S(n8654), .Z(n8164) );
  OR3_X1 U9721 ( .A1(n8649), .A2(n8255), .A3(n8166), .ZN(n8168) );
  NAND3_X1 U9722 ( .A1(n8649), .A2(n8255), .A3(n8166), .ZN(n8167) );
  MUX2_X1 U9723 ( .A(n8175), .B(n8174), .S(n8173), .Z(n8176) );
  NAND2_X1 U9724 ( .A1(n8177), .A2(n8176), .ZN(n8219) );
  NOR3_X1 U9725 ( .A1(n8219), .A2(n5650), .A3(n8178), .ZN(n8221) );
  INV_X1 U9726 ( .A(n8505), .ZN(n8209) );
  INV_X1 U9727 ( .A(n8551), .ZN(n8205) );
  INV_X1 U9728 ( .A(n8576), .ZN(n8574) );
  AND2_X1 U9729 ( .A1(n8181), .A2(n8180), .ZN(n8594) );
  AND2_X1 U9730 ( .A1(n8231), .A2(n5650), .ZN(n8182) );
  AND4_X1 U9731 ( .A1(n8185), .A2(n8184), .A3(n8183), .A4(n8182), .ZN(n8191)
         );
  INV_X1 U9732 ( .A(n10062), .ZN(n8234) );
  NOR2_X1 U9733 ( .A1(n8186), .A2(n8234), .ZN(n10069) );
  NOR2_X1 U9734 ( .A1(n8188), .A2(n8187), .ZN(n8189) );
  NAND4_X1 U9735 ( .A1(n8191), .A2(n8190), .A3(n10069), .A4(n8189), .ZN(n8194)
         );
  NOR4_X1 U9736 ( .A1(n8194), .A2(n5625), .A3(n8193), .A4(n8192), .ZN(n8198)
         );
  NAND4_X1 U9737 ( .A1(n8198), .A2(n8197), .A3(n8196), .A4(n8195), .ZN(n8199)
         );
  NOR3_X1 U9738 ( .A1(n8201), .A2(n8200), .A3(n8199), .ZN(n8202) );
  NAND4_X1 U9739 ( .A1(n8594), .A2(n8609), .A3(n8627), .A4(n8202), .ZN(n8203)
         );
  NOR2_X1 U9740 ( .A1(n8574), .A2(n8203), .ZN(n8204) );
  NAND4_X1 U9741 ( .A1(n8206), .A2(n8566), .A3(n8205), .A4(n8204), .ZN(n8207)
         );
  NOR4_X1 U9742 ( .A1(n4748), .A2(n8209), .A3(n8208), .A4(n8207), .ZN(n8210)
         );
  NAND4_X1 U9743 ( .A1(n8211), .A2(n8467), .A3(n8210), .A4(n8456), .ZN(n8212)
         );
  NOR4_X1 U9744 ( .A1(n8214), .A2(n8213), .A3(n8439), .A4(n8212), .ZN(n8215)
         );
  XNOR2_X1 U9745 ( .A(n8215), .B(n8615), .ZN(n8217) );
  INV_X1 U9746 ( .A(n8224), .ZN(n8226) );
  NAND4_X1 U9747 ( .A1(n8226), .A2(n8225), .A3(n10081), .A4(n10066), .ZN(n8227) );
  OAI211_X1 U9748 ( .C1(n8228), .C2(n8230), .A(n8227), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8229) );
  INV_X1 U9749 ( .A(n8231), .ZN(n8233) );
  MUX2_X1 U9750 ( .A(n8233), .B(n10096), .S(n8232), .Z(n8235) );
  OAI21_X1 U9751 ( .B1(n8235), .B2(n8234), .A(n8321), .ZN(n8239) );
  AOI22_X1 U9752 ( .A1(n8237), .A2(n10096), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8236), .ZN(n8238) );
  OAI211_X1 U9753 ( .C1(n5200), .C2(n8309), .A(n8239), .B(n8238), .ZN(P2_U3234) );
  INV_X1 U9754 ( .A(n8240), .ZN(n8243) );
  AOI22_X1 U9755 ( .A1(n8646), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8241), .B2(
        n10071), .ZN(n8242) );
  OAI21_X1 U9756 ( .B1(n8243), .B2(n8639), .A(n8242), .ZN(n8245) );
  AOI21_X1 U9757 ( .B1(n8251), .B2(n8250), .A(n8316), .ZN(n8252) );
  NAND2_X1 U9758 ( .A1(n8253), .A2(n8252), .ZN(n8259) );
  OAI22_X1 U9759 ( .A1(n8307), .A2(n8451), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9386), .ZN(n8257) );
  OAI22_X1 U9760 ( .A1(n8255), .A2(n8309), .B1(n8254), .B2(n8310), .ZN(n8256)
         );
  AOI211_X1 U9761 ( .C1(n8654), .C2(n8314), .A(n8257), .B(n8256), .ZN(n8258)
         );
  NAND2_X1 U9762 ( .A1(n8259), .A2(n8258), .ZN(P2_U3216) );
  XNOR2_X1 U9763 ( .A(n8260), .B(n8294), .ZN(n8265) );
  INV_X1 U9764 ( .A(n8520), .ZN(n8261) );
  OAI22_X1 U9765 ( .A1(n8307), .A2(n8261), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9304), .ZN(n8263) );
  OAI22_X1 U9766 ( .A1(n4491), .A2(n8309), .B1(n8310), .B2(n8554), .ZN(n8262)
         );
  AOI211_X1 U9767 ( .C1(n8674), .C2(n8314), .A(n8263), .B(n8262), .ZN(n8264)
         );
  OAI21_X1 U9768 ( .B1(n8265), .B2(n8316), .A(n8264), .ZN(P2_U3218) );
  INV_X1 U9769 ( .A(n8266), .ZN(n8267) );
  AOI21_X1 U9770 ( .B1(n8269), .B2(n8268), .A(n8267), .ZN(n8275) );
  NAND2_X1 U9771 ( .A1(n8343), .A2(n10066), .ZN(n8270) );
  OAI21_X1 U9772 ( .B1(n8553), .B2(n8622), .A(n8270), .ZN(n8578) );
  NOR2_X1 U9773 ( .A1(n8271), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8415) );
  AOI21_X1 U9774 ( .B1(n8286), .B2(n8578), .A(n8415), .ZN(n8272) );
  OAI21_X1 U9775 ( .B1(n8583), .B2(n8307), .A(n8272), .ZN(n8273) );
  AOI21_X1 U9776 ( .B1(n8698), .B2(n8314), .A(n8273), .ZN(n8274) );
  OAI21_X1 U9777 ( .B1(n8275), .B2(n8316), .A(n8274), .ZN(P2_U3221) );
  XNOR2_X1 U9778 ( .A(n8276), .B(n8277), .ZN(n8281) );
  OAI22_X1 U9779 ( .A1(n8307), .A2(n8545), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9451), .ZN(n8279) );
  OAI22_X1 U9780 ( .A1(n8553), .A2(n8310), .B1(n8309), .B2(n8554), .ZN(n8278)
         );
  AOI211_X1 U9781 ( .C1(n8687), .C2(n8314), .A(n8279), .B(n8278), .ZN(n8280)
         );
  OAI21_X1 U9782 ( .B1(n8281), .B2(n8316), .A(n8280), .ZN(P2_U3225) );
  XNOR2_X1 U9783 ( .A(n8283), .B(n8282), .ZN(n8284) );
  XNOR2_X1 U9784 ( .A(n8285), .B(n8284), .ZN(n8291) );
  AOI22_X1 U9785 ( .A1(n8458), .A2(n10065), .B1(n10066), .B2(n8342), .ZN(n8492) );
  INV_X1 U9786 ( .A(n8286), .ZN(n8334) );
  OAI22_X1 U9787 ( .A1(n8492), .A2(n8334), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8287), .ZN(n8289) );
  NOR2_X1 U9788 ( .A1(n4747), .A2(n8338), .ZN(n8288) );
  AOI211_X1 U9789 ( .C1(n8336), .C2(n8482), .A(n8289), .B(n8288), .ZN(n8290)
         );
  OAI21_X1 U9790 ( .B1(n8291), .B2(n8316), .A(n8290), .ZN(P2_U3227) );
  INV_X1 U9791 ( .A(n8292), .ZN(n8293) );
  OAI21_X1 U9792 ( .B1(n8260), .B2(n8294), .A(n8293), .ZN(n8298) );
  XNOR2_X1 U9793 ( .A(n8296), .B(n8295), .ZN(n8297) );
  XNOR2_X1 U9794 ( .A(n8298), .B(n8297), .ZN(n8303) );
  OAI22_X1 U9795 ( .A1(n8307), .A2(n8500), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9460), .ZN(n8301) );
  OAI22_X1 U9796 ( .A1(n8299), .A2(n8310), .B1(n8309), .B2(n8330), .ZN(n8300)
         );
  AOI211_X1 U9797 ( .C1(n8669), .C2(n8314), .A(n8301), .B(n8300), .ZN(n8302)
         );
  OAI21_X1 U9798 ( .B1(n8303), .B2(n8316), .A(n8302), .ZN(P2_U3231) );
  XNOR2_X1 U9799 ( .A(n8305), .B(n8304), .ZN(n8317) );
  OAI22_X1 U9800 ( .A1(n8307), .A2(n8561), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8306), .ZN(n8313) );
  OAI22_X1 U9801 ( .A1(n8311), .A2(n8310), .B1(n8309), .B2(n8308), .ZN(n8312)
         );
  AOI211_X1 U9802 ( .C1(n8692), .C2(n8314), .A(n8313), .B(n8312), .ZN(n8315)
         );
  OAI21_X1 U9803 ( .B1(n8317), .B2(n8316), .A(n8315), .ZN(P2_U3235) );
  OAI21_X1 U9804 ( .B1(n8320), .B2(n8319), .A(n8318), .ZN(n8322) );
  NAND2_X1 U9805 ( .A1(n8322), .A2(n8321), .ZN(n8327) );
  INV_X1 U9806 ( .A(n8323), .ZN(n8532) );
  AOI22_X1 U9807 ( .A1(n8568), .A2(n10066), .B1(n10065), .B2(n8507), .ZN(n8538) );
  OAI22_X1 U9808 ( .A1(n8538), .A2(n8334), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8324), .ZN(n8325) );
  AOI21_X1 U9809 ( .B1(n8532), .B2(n8336), .A(n8325), .ZN(n8326) );
  OAI211_X1 U9810 ( .C1(n8534), .C2(n8338), .A(n8327), .B(n8326), .ZN(P2_U3237) );
  NAND2_X1 U9811 ( .A1(n8341), .A2(n10065), .ZN(n8332) );
  OR2_X1 U9812 ( .A1(n8330), .A2(n8624), .ZN(n8331) );
  AND2_X1 U9813 ( .A1(n8332), .A2(n8331), .ZN(n8471) );
  OAI22_X1 U9814 ( .A1(n8471), .A2(n8334), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8333), .ZN(n8335) );
  AOI21_X1 U9815 ( .B1(n8475), .B2(n8336), .A(n8335), .ZN(n8337) );
  MUX2_X1 U9816 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8340), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9817 ( .A(n8459), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8358), .Z(
        P2_U3580) );
  MUX2_X1 U9818 ( .A(n8341), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8358), .Z(
        P2_U3579) );
  MUX2_X1 U9819 ( .A(n8458), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8358), .Z(
        P2_U3578) );
  MUX2_X1 U9820 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8508), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U9821 ( .A(n8342), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8358), .Z(
        P2_U3576) );
  MUX2_X1 U9822 ( .A(n8507), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8358), .Z(
        P2_U3575) );
  MUX2_X1 U9823 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n5512), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9824 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8596), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9825 ( .A(n8343), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8358), .Z(
        P2_U3570) );
  MUX2_X1 U9826 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8595), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9827 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8344), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9828 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8345), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9829 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8346), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9830 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8347), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9831 ( .A(n8348), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8358), .Z(
        P2_U3564) );
  MUX2_X1 U9832 ( .A(n8349), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8358), .Z(
        P2_U3563) );
  MUX2_X1 U9833 ( .A(n8350), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8358), .Z(
        P2_U3562) );
  MUX2_X1 U9834 ( .A(n8351), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8358), .Z(
        P2_U3561) );
  MUX2_X1 U9835 ( .A(n8352), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8358), .Z(
        P2_U3560) );
  MUX2_X1 U9836 ( .A(n8353), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8358), .Z(
        P2_U3559) );
  MUX2_X1 U9837 ( .A(n8354), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8358), .Z(
        P2_U3558) );
  MUX2_X1 U9838 ( .A(n8355), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8358), .Z(
        P2_U3557) );
  MUX2_X1 U9839 ( .A(n8356), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8358), .Z(
        P2_U3556) );
  MUX2_X1 U9840 ( .A(n8357), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8358), .Z(
        P2_U3555) );
  MUX2_X1 U9841 ( .A(n10064), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8358), .Z(
        P2_U3554) );
  MUX2_X1 U9842 ( .A(n6304), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8358), .Z(
        P2_U3553) );
  MUX2_X1 U9843 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n10067), .S(P2_U3966), .Z(
        P2_U3552) );
  OAI21_X1 U9844 ( .B1(n8361), .B2(n8360), .A(n8359), .ZN(n8362) );
  NAND2_X1 U9845 ( .A1(n10055), .A2(n8362), .ZN(n8372) );
  INV_X1 U9846 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9378) );
  OAI21_X1 U9847 ( .B1(n8417), .B2(n9378), .A(n8363), .ZN(n8364) );
  AOI21_X1 U9848 ( .B1(n10053), .B2(n8365), .A(n8364), .ZN(n8371) );
  OAI21_X1 U9849 ( .B1(n8368), .B2(n8367), .A(n8366), .ZN(n8369) );
  NAND2_X1 U9850 ( .A1(n10050), .A2(n8369), .ZN(n8370) );
  NAND3_X1 U9851 ( .A1(n8372), .A2(n8371), .A3(n8370), .ZN(P2_U3259) );
  OAI21_X1 U9852 ( .B1(n8375), .B2(n8374), .A(n8373), .ZN(n8385) );
  INV_X1 U9853 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9213) );
  NAND2_X1 U9854 ( .A1(n10053), .A2(n8376), .ZN(n8379) );
  INV_X1 U9855 ( .A(n8377), .ZN(n8378) );
  OAI211_X1 U9856 ( .C1(n8417), .C2(n9213), .A(n8379), .B(n8378), .ZN(n8384)
         );
  AOI211_X1 U9857 ( .C1(n8382), .C2(n8381), .A(n8380), .B(n9744), .ZN(n8383)
         );
  AOI211_X1 U9858 ( .C1(n8385), .C2(n10050), .A(n8384), .B(n8383), .ZN(n8386)
         );
  INV_X1 U9859 ( .A(n8386), .ZN(P2_U3261) );
  INV_X1 U9860 ( .A(n8406), .ZN(n8401) );
  INV_X1 U9861 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9426) );
  NOR2_X1 U9862 ( .A1(n8388), .A2(n9426), .ZN(n8404) );
  INV_X1 U9863 ( .A(n8404), .ZN(n8389) );
  OAI211_X1 U9864 ( .C1(n8390), .C2(P2_REG2_REG_18__SCAN_IN), .A(n8389), .B(
        n10055), .ZN(n8400) );
  INV_X1 U9865 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8391) );
  XNOR2_X1 U9866 ( .A(n8406), .B(n8391), .ZN(n8395) );
  AOI21_X1 U9867 ( .B1(n8393), .B2(P2_REG1_REG_17__SCAN_IN), .A(n8392), .ZN(
        n8394) );
  NAND2_X1 U9868 ( .A1(n8395), .A2(n8394), .ZN(n8408) );
  OAI21_X1 U9869 ( .B1(n8395), .B2(n8394), .A(n8408), .ZN(n8398) );
  INV_X1 U9870 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10222) );
  OAI21_X1 U9871 ( .B1(n8417), .B2(n10222), .A(n8396), .ZN(n8397) );
  AOI21_X1 U9872 ( .B1(n10050), .B2(n8398), .A(n8397), .ZN(n8399) );
  OAI211_X1 U9873 ( .C1(n8402), .C2(n8401), .A(n8400), .B(n8399), .ZN(P2_U3263) );
  NOR2_X1 U9874 ( .A1(n8404), .A2(n8403), .ZN(n8405) );
  XNOR2_X1 U9875 ( .A(n8405), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8412) );
  OR2_X1 U9876 ( .A1(n8406), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8407) );
  NAND2_X1 U9877 ( .A1(n8408), .A2(n8407), .ZN(n8409) );
  XNOR2_X1 U9878 ( .A(n8409), .B(n9452), .ZN(n8413) );
  INV_X1 U9879 ( .A(n8413), .ZN(n8410) );
  AOI22_X1 U9880 ( .A1(n8412), .A2(n10055), .B1(n8410), .B2(n10050), .ZN(n8414) );
  INV_X1 U9881 ( .A(n8415), .ZN(n8416) );
  NAND2_X1 U9882 ( .A1(n8420), .A2(n8419), .ZN(n9756) );
  NOR2_X1 U9883 ( .A1(n8646), .A2(n9756), .ZN(n8427) );
  AOI21_X1 U9884 ( .B1(n8646), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8427), .ZN(
        n8422) );
  NAND2_X1 U9885 ( .A1(n8418), .A2(n8619), .ZN(n8421) );
  OAI211_X1 U9886 ( .C1(n8648), .C2(n8429), .A(n8422), .B(n8421), .ZN(P2_U3265) );
  OAI21_X1 U9887 ( .B1(n8425), .B2(n8424), .A(n8423), .ZN(n9757) );
  NOR2_X1 U9888 ( .A1(n8425), .A2(n8639), .ZN(n8426) );
  AOI211_X1 U9889 ( .C1(n8646), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8427), .B(
        n8426), .ZN(n8428) );
  OAI21_X1 U9890 ( .B1(n8429), .B2(n9757), .A(n8428), .ZN(P2_U3266) );
  XNOR2_X1 U9891 ( .A(n8431), .B(n8430), .ZN(n8653) );
  INV_X1 U9892 ( .A(n8450), .ZN(n8434) );
  INV_X1 U9893 ( .A(n8432), .ZN(n8433) );
  AOI22_X1 U9894 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(n8646), .B1(n8435), .B2(
        n10071), .ZN(n8436) );
  OAI21_X1 U9895 ( .B1(n8437), .B2(n8639), .A(n8436), .ZN(n8447) );
  INV_X1 U9896 ( .A(n8438), .ZN(n8440) );
  AOI21_X1 U9897 ( .B1(n8440), .B2(n8439), .A(n8612), .ZN(n8445) );
  OAI22_X1 U9898 ( .A1(n8442), .A2(n8622), .B1(n8441), .B2(n8624), .ZN(n8443)
         );
  AOI21_X1 U9899 ( .B1(n8445), .B2(n8444), .A(n8443), .ZN(n8652) );
  NOR2_X1 U9900 ( .A1(n8652), .A2(n8646), .ZN(n8446) );
  AOI211_X1 U9901 ( .C1(n8644), .C2(n8650), .A(n8447), .B(n8446), .ZN(n8448)
         );
  OAI21_X1 U9902 ( .B1(n8653), .B2(n8557), .A(n8448), .ZN(P2_U3268) );
  XOR2_X1 U9903 ( .A(n8456), .B(n8449), .Z(n8658) );
  AOI21_X1 U9904 ( .B1(n8654), .B2(n8473), .A(n8450), .ZN(n8655) );
  INV_X1 U9905 ( .A(n8654), .ZN(n8454) );
  INV_X1 U9906 ( .A(n8451), .ZN(n8452) );
  AOI22_X1 U9907 ( .A1(n8646), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8452), .B2(
        n10071), .ZN(n8453) );
  OAI21_X1 U9908 ( .B1(n8454), .B2(n8639), .A(n8453), .ZN(n8463) );
  OAI211_X1 U9909 ( .C1(n8457), .C2(n8456), .A(n8455), .B(n10061), .ZN(n8461)
         );
  AOI22_X1 U9910 ( .A1(n8459), .A2(n10065), .B1(n10066), .B2(n8458), .ZN(n8460) );
  NOR2_X1 U9911 ( .A1(n8657), .A2(n8646), .ZN(n8462) );
  AOI211_X1 U9912 ( .C1(n8644), .C2(n8655), .A(n8463), .B(n8462), .ZN(n8464)
         );
  OAI21_X1 U9913 ( .B1(n8658), .B2(n8557), .A(n8464), .ZN(P2_U3269) );
  XNOR2_X1 U9914 ( .A(n8465), .B(n8467), .ZN(n8663) );
  AOI22_X1 U9915 ( .A1(n8661), .A2(n8619), .B1(n8646), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8480) );
  INV_X1 U9916 ( .A(n8466), .ZN(n8470) );
  AOI21_X1 U9917 ( .B1(n8489), .B2(n8468), .A(n8467), .ZN(n8469) );
  OAI21_X1 U9918 ( .B1(n8470), .B2(n8469), .A(n10061), .ZN(n8472) );
  NAND2_X1 U9919 ( .A1(n8472), .A2(n8471), .ZN(n8659) );
  INV_X1 U9920 ( .A(n8473), .ZN(n8474) );
  AOI211_X1 U9921 ( .C1(n8661), .C2(n8486), .A(n10155), .B(n8474), .ZN(n8660)
         );
  INV_X1 U9922 ( .A(n8660), .ZN(n8477) );
  INV_X1 U9923 ( .A(n8475), .ZN(n8476) );
  OAI22_X1 U9924 ( .A1(n8477), .A2(n5638), .B1(n8604), .B2(n8476), .ZN(n8478)
         );
  OAI21_X1 U9925 ( .B1(n8659), .B2(n8478), .A(n6401), .ZN(n8479) );
  OAI211_X1 U9926 ( .C1(n8663), .C2(n8557), .A(n8480), .B(n8479), .ZN(P2_U3270) );
  XNOR2_X1 U9927 ( .A(n8481), .B(n4748), .ZN(n8668) );
  INV_X1 U9928 ( .A(n8482), .ZN(n8483) );
  OAI22_X1 U9929 ( .A1(n6401), .A2(n8484), .B1(n8483), .B2(n8604), .ZN(n8496)
         );
  INV_X1 U9930 ( .A(n8485), .ZN(n8488) );
  INV_X1 U9931 ( .A(n8486), .ZN(n8487) );
  AOI211_X1 U9932 ( .C1(n8666), .C2(n8488), .A(n10155), .B(n8487), .ZN(n8665)
         );
  OAI211_X1 U9933 ( .C1(n8491), .C2(n8490), .A(n8489), .B(n10061), .ZN(n8493)
         );
  NAND2_X1 U9934 ( .A1(n8493), .A2(n8492), .ZN(n8664) );
  AOI21_X1 U9935 ( .B1(n8665), .B2(n8615), .A(n8664), .ZN(n8494) );
  NOR2_X1 U9936 ( .A1(n8494), .A2(n8646), .ZN(n8495) );
  AOI211_X1 U9937 ( .C1(n8619), .C2(n8666), .A(n8496), .B(n8495), .ZN(n8497)
         );
  OAI21_X1 U9938 ( .B1(n8668), .B2(n8557), .A(n8497), .ZN(P2_U3271) );
  AOI21_X1 U9939 ( .B1(n8505), .B2(n8498), .A(n8499), .ZN(n8673) );
  XNOR2_X1 U9940 ( .A(n8518), .B(n8503), .ZN(n8670) );
  INV_X1 U9941 ( .A(n8500), .ZN(n8501) );
  AOI22_X1 U9942 ( .A1(n8646), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8501), .B2(
        n10071), .ZN(n8502) );
  OAI21_X1 U9943 ( .B1(n8503), .B2(n8639), .A(n8502), .ZN(n8512) );
  OAI211_X1 U9944 ( .C1(n8506), .C2(n8505), .A(n8504), .B(n10061), .ZN(n8510)
         );
  AOI22_X1 U9945 ( .A1(n8508), .A2(n10065), .B1(n10066), .B2(n8507), .ZN(n8509) );
  NOR2_X1 U9946 ( .A1(n8672), .A2(n8646), .ZN(n8511) );
  AOI211_X1 U9947 ( .C1(n8670), .C2(n8644), .A(n8512), .B(n8511), .ZN(n8513)
         );
  OAI21_X1 U9948 ( .B1(n8673), .B2(n8557), .A(n8513), .ZN(P2_U3272) );
  AOI21_X1 U9949 ( .B1(n8524), .B2(n8515), .A(n8514), .ZN(n8516) );
  OAI222_X1 U9950 ( .A1(n8624), .A2(n8554), .B1(n8622), .B2(n4491), .C1(n8612), 
        .C2(n8516), .ZN(n8517) );
  INV_X1 U9951 ( .A(n8517), .ZN(n8680) );
  INV_X1 U9952 ( .A(n8518), .ZN(n8519) );
  AOI21_X1 U9953 ( .B1(n8674), .B2(n8529), .A(n8519), .ZN(n8675) );
  AOI22_X1 U9954 ( .A1(n8646), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8520), .B2(
        n10071), .ZN(n8521) );
  OAI21_X1 U9955 ( .B1(n8522), .B2(n8639), .A(n8521), .ZN(n8523) );
  AOI21_X1 U9956 ( .B1(n8675), .B2(n8644), .A(n8523), .ZN(n8527) );
  OR2_X1 U9957 ( .A1(n8525), .A2(n8524), .ZN(n8677) );
  NAND3_X1 U9958 ( .A1(n8677), .A2(n8676), .A3(n10077), .ZN(n8526) );
  OAI211_X1 U9959 ( .C1(n8680), .C2(n8646), .A(n8527), .B(n8526), .ZN(P2_U3273) );
  XNOR2_X1 U9960 ( .A(n8528), .B(n8536), .ZN(n8685) );
  INV_X1 U9961 ( .A(n8529), .ZN(n8530) );
  AOI21_X1 U9962 ( .B1(n8681), .B2(n8531), .A(n8530), .ZN(n8682) );
  AOI22_X1 U9963 ( .A1(n8646), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8532), .B2(
        n10071), .ZN(n8533) );
  OAI21_X1 U9964 ( .B1(n8534), .B2(n8639), .A(n8533), .ZN(n8541) );
  OAI211_X1 U9965 ( .C1(n8537), .C2(n8536), .A(n8535), .B(n10061), .ZN(n8539)
         );
  NOR2_X1 U9966 ( .A1(n8684), .A2(n8646), .ZN(n8540) );
  AOI211_X1 U9967 ( .C1(n8682), .C2(n8644), .A(n8541), .B(n8540), .ZN(n8542)
         );
  OAI21_X1 U9968 ( .B1(n8685), .B2(n8557), .A(n8542), .ZN(P2_U3274) );
  XNOR2_X1 U9969 ( .A(n8543), .B(n8551), .ZN(n8691) );
  XNOR2_X1 U9970 ( .A(n8559), .B(n8687), .ZN(n8688) );
  NOR2_X1 U9971 ( .A1(n8544), .A2(n8639), .ZN(n8548) );
  OAI22_X1 U9972 ( .A1(n6401), .A2(n8546), .B1(n8545), .B2(n8604), .ZN(n8547)
         );
  AOI211_X1 U9973 ( .C1(n8688), .C2(n8644), .A(n8548), .B(n8547), .ZN(n8556)
         );
  AOI21_X1 U9974 ( .B1(n8551), .B2(n8550), .A(n8549), .ZN(n8552) );
  OAI222_X1 U9975 ( .A1(n8622), .A2(n8554), .B1(n8624), .B2(n8553), .C1(n8612), 
        .C2(n8552), .ZN(n8686) );
  NAND2_X1 U9976 ( .A1(n8686), .A2(n6401), .ZN(n8555) );
  OAI211_X1 U9977 ( .C1(n8691), .C2(n8557), .A(n8556), .B(n8555), .ZN(P2_U3275) );
  XNOR2_X1 U9978 ( .A(n8558), .B(n8566), .ZN(n8696) );
  INV_X1 U9979 ( .A(n8580), .ZN(n8560) );
  AOI21_X1 U9980 ( .B1(n8692), .B2(n8560), .A(n8559), .ZN(n8693) );
  INV_X1 U9981 ( .A(n8561), .ZN(n8562) );
  AOI22_X1 U9982 ( .A1(n8646), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8562), .B2(
        n10071), .ZN(n8563) );
  OAI21_X1 U9983 ( .B1(n8564), .B2(n8639), .A(n8563), .ZN(n8572) );
  OAI211_X1 U9984 ( .C1(n8567), .C2(n8566), .A(n8565), .B(n10061), .ZN(n8570)
         );
  AOI22_X1 U9985 ( .A1(n10066), .A2(n8596), .B1(n8568), .B2(n10065), .ZN(n8569) );
  NOR2_X1 U9986 ( .A1(n8695), .A2(n8646), .ZN(n8571) );
  AOI211_X1 U9987 ( .C1(n8693), .C2(n8644), .A(n8572), .B(n8571), .ZN(n8573)
         );
  OAI21_X1 U9988 ( .B1(n8696), .B2(n8557), .A(n8573), .ZN(P2_U3276) );
  XNOR2_X1 U9989 ( .A(n8575), .B(n8574), .ZN(n8701) );
  XNOR2_X1 U9990 ( .A(n8577), .B(n8576), .ZN(n8579) );
  AOI21_X1 U9991 ( .B1(n8579), .B2(n10061), .A(n8578), .ZN(n8700) );
  AOI211_X1 U9992 ( .C1(n8698), .C2(n4413), .A(n10155), .B(n8580), .ZN(n8697)
         );
  NAND2_X1 U9993 ( .A1(n8697), .A2(n8615), .ZN(n8581) );
  OAI211_X1 U9994 ( .C1(n8701), .C2(n8630), .A(n8700), .B(n8581), .ZN(n8582)
         );
  NAND2_X1 U9995 ( .A1(n8582), .A2(n6401), .ZN(n8586) );
  OAI22_X1 U9996 ( .A1(n6401), .A2(n9421), .B1(n8583), .B2(n8604), .ZN(n8584)
         );
  AOI21_X1 U9997 ( .B1(n8698), .B2(n8619), .A(n8584), .ZN(n8585) );
  OAI211_X1 U9998 ( .C1(n8701), .C2(n8641), .A(n8586), .B(n8585), .ZN(P2_U3277) );
  XNOR2_X1 U9999 ( .A(n8587), .B(n8594), .ZN(n8706) );
  INV_X1 U10000 ( .A(n4413), .ZN(n8588) );
  AOI21_X1 U10001 ( .B1(n8702), .B2(n8607), .A(n8588), .ZN(n8703) );
  INV_X1 U10002 ( .A(n8589), .ZN(n8590) );
  AOI22_X1 U10003 ( .A1(n8646), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8590), .B2(
        n10071), .ZN(n8591) );
  OAI21_X1 U10004 ( .B1(n8592), .B2(n8639), .A(n8591), .ZN(n8599) );
  XOR2_X1 U10005 ( .A(n8594), .B(n8593), .Z(n8597) );
  AOI222_X1 U10006 ( .A1(n10061), .A2(n8597), .B1(n8596), .B2(n10065), .C1(
        n8595), .C2(n10066), .ZN(n8705) );
  NOR2_X1 U10007 ( .A1(n8705), .A2(n8646), .ZN(n8598) );
  AOI211_X1 U10008 ( .C1(n8703), .C2(n8644), .A(n8599), .B(n8598), .ZN(n8600)
         );
  OAI21_X1 U10009 ( .B1(n8706), .B2(n8557), .A(n8600), .ZN(P2_U3278) );
  INV_X1 U10010 ( .A(n8601), .ZN(n8602) );
  AOI21_X1 U10011 ( .B1(n8609), .B2(n8603), .A(n8602), .ZN(n8711) );
  OAI22_X1 U10012 ( .A1(n6401), .A2(n8606), .B1(n8605), .B2(n8604), .ZN(n8618)
         );
  INV_X1 U10013 ( .A(n8635), .ZN(n8608) );
  AOI211_X1 U10014 ( .C1(n8709), .C2(n8608), .A(n10155), .B(n4381), .ZN(n8708)
         );
  XNOR2_X1 U10015 ( .A(n8610), .B(n8609), .ZN(n8611) );
  OAI222_X1 U10016 ( .A1(n8622), .A2(n8614), .B1(n8624), .B2(n8613), .C1(n8612), .C2(n8611), .ZN(n8707) );
  AOI21_X1 U10017 ( .B1(n8708), .B2(n8615), .A(n8707), .ZN(n8616) );
  NOR2_X1 U10018 ( .A1(n8616), .A2(n8646), .ZN(n8617) );
  AOI211_X1 U10019 ( .C1(n8619), .C2(n8709), .A(n8618), .B(n8617), .ZN(n8620)
         );
  OAI21_X1 U10020 ( .B1(n8711), .B2(n8557), .A(n8620), .ZN(P2_U3279) );
  XNOR2_X1 U10021 ( .A(n8621), .B(n8627), .ZN(n8633) );
  OAI22_X1 U10022 ( .A1(n8625), .A2(n8624), .B1(n8623), .B2(n8622), .ZN(n8632)
         );
  NAND2_X1 U10023 ( .A1(n8626), .A2(n8627), .ZN(n8628) );
  NAND2_X1 U10024 ( .A1(n8629), .A2(n8628), .ZN(n8716) );
  NOR2_X1 U10025 ( .A1(n8716), .A2(n8630), .ZN(n8631) );
  AOI211_X1 U10026 ( .C1(n8633), .C2(n10061), .A(n8632), .B(n8631), .ZN(n8715)
         );
  INV_X1 U10027 ( .A(n8634), .ZN(n8636) );
  AOI21_X1 U10028 ( .B1(n8712), .B2(n8636), .A(n8635), .ZN(n8713) );
  AOI22_X1 U10029 ( .A1(n8646), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8637), .B2(
        n10071), .ZN(n8638) );
  OAI21_X1 U10030 ( .B1(n8640), .B2(n8639), .A(n8638), .ZN(n8643) );
  NOR2_X1 U10031 ( .A1(n8716), .A2(n8641), .ZN(n8642) );
  AOI211_X1 U10032 ( .C1(n8713), .C2(n8644), .A(n8643), .B(n8642), .ZN(n8645)
         );
  OAI21_X1 U10033 ( .B1(n8715), .B2(n8646), .A(n8645), .ZN(P2_U3280) );
  NAND2_X1 U10034 ( .A1(n8418), .A2(n10137), .ZN(n8647) );
  OAI211_X1 U10035 ( .C1(n8648), .C2(n10155), .A(n9756), .B(n8647), .ZN(n8737)
         );
  MUX2_X1 U10036 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8737), .S(n10177), .Z(
        P2_U3551) );
  AOI22_X1 U10037 ( .A1(n8650), .A2(n10138), .B1(n10137), .B2(n8649), .ZN(
        n8651) );
  OAI211_X1 U10038 ( .C1(n8653), .C2(n10132), .A(n8652), .B(n8651), .ZN(n8738)
         );
  MUX2_X1 U10039 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8738), .S(n10177), .Z(
        P2_U3548) );
  AOI22_X1 U10040 ( .A1(n8655), .A2(n10138), .B1(n10137), .B2(n8654), .ZN(
        n8656) );
  OAI211_X1 U10041 ( .C1(n8658), .C2(n10132), .A(n8657), .B(n8656), .ZN(n8739)
         );
  MUX2_X1 U10042 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8739), .S(n10177), .Z(
        P2_U3547) );
  AOI211_X1 U10043 ( .C1(n10137), .C2(n8661), .A(n8660), .B(n8659), .ZN(n8662)
         );
  OAI21_X1 U10044 ( .B1(n8663), .B2(n10132), .A(n8662), .ZN(n8740) );
  MUX2_X1 U10045 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8740), .S(n10177), .Z(
        P2_U3546) );
  AOI211_X1 U10046 ( .C1(n10137), .C2(n8666), .A(n8665), .B(n8664), .ZN(n8667)
         );
  OAI21_X1 U10047 ( .B1(n8668), .B2(n10132), .A(n8667), .ZN(n8741) );
  MUX2_X1 U10048 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8741), .S(n10177), .Z(
        P2_U3545) );
  AOI22_X1 U10049 ( .A1(n8670), .A2(n10138), .B1(n10137), .B2(n8669), .ZN(
        n8671) );
  OAI211_X1 U10050 ( .C1(n8673), .C2(n10132), .A(n8672), .B(n8671), .ZN(n8742)
         );
  MUX2_X1 U10051 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8742), .S(n10177), .Z(
        P2_U3544) );
  AOI22_X1 U10052 ( .A1(n8675), .A2(n10138), .B1(n10137), .B2(n8674), .ZN(
        n8679) );
  INV_X1 U10053 ( .A(n10132), .ZN(n10159) );
  NAND3_X1 U10054 ( .A1(n8677), .A2(n8676), .A3(n10159), .ZN(n8678) );
  NAND3_X1 U10055 ( .A1(n8680), .A2(n8679), .A3(n8678), .ZN(n8743) );
  MUX2_X1 U10056 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8743), .S(n10177), .Z(
        P2_U3543) );
  AOI22_X1 U10057 ( .A1(n8682), .A2(n10138), .B1(n10137), .B2(n8681), .ZN(
        n8683) );
  OAI211_X1 U10058 ( .C1(n8685), .C2(n10132), .A(n8684), .B(n8683), .ZN(n8744)
         );
  MUX2_X1 U10059 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8744), .S(n10177), .Z(
        P2_U3542) );
  INV_X1 U10060 ( .A(n8686), .ZN(n8690) );
  AOI22_X1 U10061 ( .A1(n8688), .A2(n10138), .B1(n10137), .B2(n8687), .ZN(
        n8689) );
  OAI211_X1 U10062 ( .C1(n8691), .C2(n10132), .A(n8690), .B(n8689), .ZN(n8745)
         );
  MUX2_X1 U10063 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8745), .S(n10177), .Z(
        P2_U3541) );
  AOI22_X1 U10064 ( .A1(n8693), .A2(n10138), .B1(n10137), .B2(n8692), .ZN(
        n8694) );
  OAI211_X1 U10065 ( .C1(n8696), .C2(n10132), .A(n8695), .B(n8694), .ZN(n8746)
         );
  MUX2_X1 U10066 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8746), .S(n10177), .Z(
        P2_U3540) );
  AOI21_X1 U10067 ( .B1(n10137), .B2(n8698), .A(n8697), .ZN(n8699) );
  OAI211_X1 U10068 ( .C1(n8701), .C2(n10132), .A(n8700), .B(n8699), .ZN(n8747)
         );
  MUX2_X1 U10069 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8747), .S(n10177), .Z(
        P2_U3539) );
  AOI22_X1 U10070 ( .A1(n8703), .A2(n10138), .B1(n10137), .B2(n8702), .ZN(
        n8704) );
  OAI211_X1 U10071 ( .C1(n8706), .C2(n10132), .A(n8705), .B(n8704), .ZN(n8748)
         );
  MUX2_X1 U10072 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8748), .S(n10177), .Z(
        P2_U3538) );
  AOI211_X1 U10073 ( .C1(n10137), .C2(n8709), .A(n8708), .B(n8707), .ZN(n8710)
         );
  OAI21_X1 U10074 ( .B1(n8711), .B2(n10132), .A(n8710), .ZN(n8749) );
  MUX2_X1 U10075 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8749), .S(n10177), .Z(
        P2_U3537) );
  AOI22_X1 U10076 ( .A1(n8713), .A2(n10138), .B1(n10137), .B2(n8712), .ZN(
        n8714) );
  OAI211_X1 U10077 ( .C1(n10142), .C2(n8716), .A(n8715), .B(n8714), .ZN(n8750)
         );
  MUX2_X1 U10078 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8750), .S(n10177), .Z(
        P2_U3536) );
  INV_X1 U10079 ( .A(n8717), .ZN(n8722) );
  AOI22_X1 U10080 ( .A1(n8719), .A2(n10138), .B1(n10137), .B2(n8718), .ZN(
        n8720) );
  OAI211_X1 U10081 ( .C1(n8722), .C2(n10132), .A(n8721), .B(n8720), .ZN(n8751)
         );
  MUX2_X1 U10082 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8751), .S(n10177), .Z(
        P2_U3535) );
  AOI22_X1 U10083 ( .A1(n8724), .A2(n10138), .B1(n10137), .B2(n8723), .ZN(
        n8725) );
  OAI211_X1 U10084 ( .C1(n8727), .C2(n10132), .A(n8726), .B(n8725), .ZN(n8752)
         );
  MUX2_X1 U10085 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8752), .S(n10177), .Z(
        P2_U3534) );
  AOI22_X1 U10086 ( .A1(n8729), .A2(n10138), .B1(n10137), .B2(n8728), .ZN(
        n8730) );
  OAI211_X1 U10087 ( .C1(n8732), .C2(n10132), .A(n8731), .B(n8730), .ZN(n8753)
         );
  MUX2_X1 U10088 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8753), .S(n10177), .Z(
        P2_U3533) );
  AOI22_X1 U10089 ( .A1(n8733), .A2(n10138), .B1(n10137), .B2(n5739), .ZN(
        n8734) );
  OAI211_X1 U10090 ( .C1(n8736), .C2(n10132), .A(n8735), .B(n8734), .ZN(n8754)
         );
  MUX2_X1 U10091 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8754), .S(n10177), .Z(
        P2_U3531) );
  MUX2_X1 U10092 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8737), .S(n10163), .Z(
        P2_U3519) );
  MUX2_X1 U10093 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8738), .S(n10163), .Z(
        P2_U3516) );
  MUX2_X1 U10094 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8739), .S(n10163), .Z(
        P2_U3515) );
  MUX2_X1 U10095 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8740), .S(n10163), .Z(
        P2_U3514) );
  MUX2_X1 U10096 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8741), .S(n10163), .Z(
        P2_U3513) );
  MUX2_X1 U10097 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8742), .S(n10163), .Z(
        P2_U3512) );
  MUX2_X1 U10098 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8743), .S(n10163), .Z(
        P2_U3511) );
  MUX2_X1 U10099 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8744), .S(n10163), .Z(
        P2_U3510) );
  MUX2_X1 U10100 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8745), .S(n10163), .Z(
        P2_U3509) );
  MUX2_X1 U10101 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8746), .S(n10163), .Z(
        P2_U3508) );
  MUX2_X1 U10102 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8747), .S(n10163), .Z(
        P2_U3507) );
  MUX2_X1 U10103 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8748), .S(n10163), .Z(
        P2_U3505) );
  MUX2_X1 U10104 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8749), .S(n10163), .Z(
        P2_U3502) );
  MUX2_X1 U10105 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8750), .S(n10163), .Z(
        P2_U3499) );
  MUX2_X1 U10106 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8751), .S(n10163), .Z(
        P2_U3496) );
  MUX2_X1 U10107 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8752), .S(n10163), .Z(
        P2_U3493) );
  MUX2_X1 U10108 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8753), .S(n10163), .Z(
        P2_U3490) );
  MUX2_X1 U10109 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n8754), .S(n10163), .Z(
        P2_U3484) );
  NAND4_X1 U10110 ( .A1(n8755), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .A4(n5171), .ZN(n8758) );
  NAND2_X1 U10111 ( .A1(n8756), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8757) );
  OAI211_X1 U10112 ( .C1(n8759), .C2(n4385), .A(n8758), .B(n8757), .ZN(
        P2_U3327) );
  INV_X1 U10113 ( .A(n8760), .ZN(n9694) );
  OAI222_X1 U10114 ( .A1(n8763), .A2(P2_U3152), .B1(n4385), .B2(n9694), .C1(
        n8762), .C2(n8761), .ZN(P2_U3329) );
  MUX2_X1 U10115 ( .A(n8764), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  AND2_X1 U10116 ( .A1(n8766), .A2(n8765), .ZN(n8767) );
  INV_X1 U10117 ( .A(n8778), .ZN(n8773) );
  NAND2_X1 U10118 ( .A1(n8774), .A2(n8918), .ZN(n8770) );
  NAND2_X1 U10119 ( .A1(n9059), .A2(n8925), .ZN(n8769) );
  NAND2_X1 U10120 ( .A1(n8770), .A2(n8769), .ZN(n8771) );
  XNOR2_X1 U10121 ( .A(n8771), .B(n6247), .ZN(n8777) );
  INV_X1 U10122 ( .A(n8777), .ZN(n8772) );
  NAND2_X1 U10123 ( .A1(n8773), .A2(n8772), .ZN(n8888) );
  NAND2_X1 U10124 ( .A1(n8774), .A2(n8925), .ZN(n8776) );
  NAND2_X1 U10125 ( .A1(n9059), .A2(n8924), .ZN(n8775) );
  NAND2_X1 U10126 ( .A1(n8776), .A2(n8775), .ZN(n8890) );
  NAND2_X1 U10127 ( .A1(n8778), .A2(n8777), .ZN(n8889) );
  NAND2_X1 U10128 ( .A1(n9669), .A2(n8918), .ZN(n8780) );
  NAND2_X1 U10129 ( .A1(n9058), .A2(n8925), .ZN(n8779) );
  NAND2_X1 U10130 ( .A1(n8780), .A2(n8779), .ZN(n8781) );
  XNOR2_X1 U10131 ( .A(n8781), .B(n6247), .ZN(n8785) );
  NAND2_X1 U10132 ( .A1(n9669), .A2(n8919), .ZN(n8784) );
  NAND2_X1 U10133 ( .A1(n9058), .A2(n8924), .ZN(n8783) );
  NAND2_X1 U10134 ( .A1(n8784), .A2(n8783), .ZN(n9039) );
  NAND2_X1 U10135 ( .A1(n9037), .A2(n9039), .ZN(n8787) );
  NAND2_X1 U10136 ( .A1(n8786), .A2(n8785), .ZN(n9038) );
  NAND2_X1 U10137 ( .A1(n9666), .A2(n8918), .ZN(n8789) );
  NAND2_X1 U10138 ( .A1(n9593), .A2(n8919), .ZN(n8788) );
  NAND2_X1 U10139 ( .A1(n8789), .A2(n8788), .ZN(n8790) );
  XNOR2_X1 U10140 ( .A(n8790), .B(n6247), .ZN(n8964) );
  NAND2_X1 U10141 ( .A1(n9666), .A2(n8919), .ZN(n8792) );
  NAND2_X1 U10142 ( .A1(n9593), .A2(n8924), .ZN(n8791) );
  NAND2_X1 U10143 ( .A1(n8792), .A2(n8791), .ZN(n8965) );
  NAND2_X1 U10144 ( .A1(n9659), .A2(n8918), .ZN(n8794) );
  NAND2_X1 U10145 ( .A1(n9568), .A2(n8925), .ZN(n8793) );
  NAND2_X1 U10146 ( .A1(n8794), .A2(n8793), .ZN(n8795) );
  XNOR2_X1 U10147 ( .A(n8795), .B(n8922), .ZN(n8798) );
  AND2_X1 U10148 ( .A1(n9568), .A2(n8924), .ZN(n8796) );
  AOI21_X1 U10149 ( .B1(n9659), .B2(n8925), .A(n8796), .ZN(n8797) );
  XNOR2_X1 U10150 ( .A(n8798), .B(n8797), .ZN(n8974) );
  NAND2_X1 U10151 ( .A1(n8798), .A2(n8797), .ZN(n8799) );
  NAND2_X1 U10152 ( .A1(n9655), .A2(n8918), .ZN(n8801) );
  NAND2_X1 U10153 ( .A1(n9583), .A2(n8925), .ZN(n8800) );
  NAND2_X1 U10154 ( .A1(n8801), .A2(n8800), .ZN(n8802) );
  XNOR2_X1 U10155 ( .A(n8802), .B(n8922), .ZN(n8806) );
  NAND2_X1 U10156 ( .A1(n8805), .A2(n8806), .ZN(n9013) );
  NAND2_X1 U10157 ( .A1(n9655), .A2(n8919), .ZN(n8804) );
  NAND2_X1 U10158 ( .A1(n9583), .A2(n8924), .ZN(n8803) );
  NAND2_X1 U10159 ( .A1(n8804), .A2(n8803), .ZN(n9012) );
  NAND2_X1 U10160 ( .A1(n9013), .A2(n9012), .ZN(n9017) );
  INV_X1 U10161 ( .A(n8805), .ZN(n8808) );
  INV_X1 U10162 ( .A(n8806), .ZN(n8807) );
  NAND2_X1 U10163 ( .A1(n9651), .A2(n8918), .ZN(n8810) );
  NAND2_X1 U10164 ( .A1(n9569), .A2(n8925), .ZN(n8809) );
  NAND2_X1 U10165 ( .A1(n8810), .A2(n8809), .ZN(n8811) );
  XNOR2_X1 U10166 ( .A(n8811), .B(n6247), .ZN(n8814) );
  NAND2_X1 U10167 ( .A1(n9651), .A2(n8919), .ZN(n8813) );
  NAND2_X1 U10168 ( .A1(n9569), .A2(n8924), .ZN(n8812) );
  NAND2_X1 U10169 ( .A1(n8813), .A2(n8812), .ZN(n8815) );
  INV_X1 U10170 ( .A(n8814), .ZN(n8817) );
  INV_X1 U10171 ( .A(n8815), .ZN(n8816) );
  NAND2_X1 U10172 ( .A1(n8817), .A2(n8816), .ZN(n8906) );
  NAND2_X1 U10173 ( .A1(n9644), .A2(n8918), .ZN(n8819) );
  NAND2_X1 U10174 ( .A1(n9518), .A2(n8925), .ZN(n8818) );
  NAND2_X1 U10175 ( .A1(n8819), .A2(n8818), .ZN(n8820) );
  XNOR2_X1 U10176 ( .A(n8820), .B(n6247), .ZN(n8834) );
  NAND2_X1 U10177 ( .A1(n9644), .A2(n8925), .ZN(n8822) );
  NAND2_X1 U10178 ( .A1(n9518), .A2(n8924), .ZN(n8821) );
  NAND2_X1 U10179 ( .A1(n8822), .A2(n8821), .ZN(n8835) );
  NAND2_X1 U10180 ( .A1(n8834), .A2(n8835), .ZN(n8990) );
  NAND2_X1 U10181 ( .A1(n9640), .A2(n8918), .ZN(n8824) );
  NAND2_X1 U10182 ( .A1(n9532), .A2(n8925), .ZN(n8823) );
  NAND2_X1 U10183 ( .A1(n8824), .A2(n8823), .ZN(n8825) );
  XNOR2_X1 U10184 ( .A(n8825), .B(n6247), .ZN(n8829) );
  INV_X1 U10185 ( .A(n8829), .ZN(n8827) );
  AND2_X1 U10186 ( .A1(n9532), .A2(n8924), .ZN(n8826) );
  AOI21_X1 U10187 ( .B1(n9640), .B2(n8925), .A(n8826), .ZN(n8828) );
  XNOR2_X1 U10188 ( .A(n8829), .B(n8828), .ZN(n8950) );
  AND2_X1 U10189 ( .A1(n9519), .A2(n8924), .ZN(n8830) );
  AOI21_X1 U10190 ( .B1(n9634), .B2(n8925), .A(n8830), .ZN(n8832) );
  AND2_X1 U10191 ( .A1(n8844), .A2(n8832), .ZN(n8831) );
  INV_X1 U10192 ( .A(n8832), .ZN(n8845) );
  INV_X1 U10193 ( .A(n8833), .ZN(n8840) );
  INV_X1 U10194 ( .A(n8834), .ZN(n8837) );
  INV_X1 U10195 ( .A(n8835), .ZN(n8836) );
  NAND2_X1 U10196 ( .A1(n8837), .A2(n8836), .ZN(n8991) );
  AND2_X1 U10197 ( .A1(n8991), .A2(n8838), .ZN(n8839) );
  NAND2_X1 U10198 ( .A1(n9634), .A2(n8918), .ZN(n8842) );
  NAND2_X1 U10199 ( .A1(n9519), .A2(n8925), .ZN(n8841) );
  NAND2_X1 U10200 ( .A1(n8842), .A2(n8841), .ZN(n8843) );
  XNOR2_X1 U10201 ( .A(n8843), .B(n6247), .ZN(n9003) );
  NAND2_X1 U10202 ( .A1(n9631), .A2(n8918), .ZN(n8849) );
  NAND2_X1 U10203 ( .A1(n9502), .A2(n8925), .ZN(n8848) );
  NAND2_X1 U10204 ( .A1(n8849), .A2(n8848), .ZN(n8850) );
  XNOR2_X1 U10205 ( .A(n8850), .B(n6247), .ZN(n8854) );
  AND2_X1 U10206 ( .A1(n9502), .A2(n8924), .ZN(n8852) );
  AOI21_X1 U10207 ( .B1(n9631), .B2(n8919), .A(n8852), .ZN(n8898) );
  INV_X1 U10208 ( .A(n8854), .ZN(n8855) );
  NAND2_X1 U10209 ( .A1(n9201), .A2(n8918), .ZN(n8859) );
  NAND2_X1 U10210 ( .A1(n9057), .A2(n8925), .ZN(n8858) );
  NAND2_X1 U10211 ( .A1(n8859), .A2(n8858), .ZN(n8860) );
  XNOR2_X1 U10212 ( .A(n8860), .B(n8922), .ZN(n8862) );
  AND2_X1 U10213 ( .A1(n9057), .A2(n8924), .ZN(n8861) );
  AOI21_X1 U10214 ( .B1(n9201), .B2(n8925), .A(n8861), .ZN(n8863) );
  NAND2_X1 U10215 ( .A1(n8862), .A2(n8863), .ZN(n8867) );
  INV_X1 U10216 ( .A(n8862), .ZN(n8865) );
  INV_X1 U10217 ( .A(n8863), .ZN(n8864) );
  NAND2_X1 U10218 ( .A1(n8865), .A2(n8864), .ZN(n8866) );
  NAND2_X1 U10219 ( .A1(n8867), .A2(n8866), .ZN(n8979) );
  AOI22_X1 U10220 ( .A1(n9619), .A2(n8925), .B1(n8924), .B2(n9196), .ZN(n8872)
         );
  NAND2_X1 U10221 ( .A1(n9619), .A2(n8918), .ZN(n8869) );
  NAND2_X1 U10222 ( .A1(n9196), .A2(n8925), .ZN(n8868) );
  NAND2_X1 U10223 ( .A1(n8869), .A2(n8868), .ZN(n8870) );
  XNOR2_X1 U10224 ( .A(n8870), .B(n6247), .ZN(n8871) );
  XOR2_X1 U10225 ( .A(n8872), .B(n8871), .Z(n8957) );
  INV_X1 U10226 ( .A(n8871), .ZN(n8873) );
  NAND2_X1 U10227 ( .A1(n9614), .A2(n8918), .ZN(n8875) );
  NAND2_X1 U10228 ( .A1(n9056), .A2(n8919), .ZN(n8874) );
  NAND2_X1 U10229 ( .A1(n8875), .A2(n8874), .ZN(n8876) );
  XNOR2_X1 U10230 ( .A(n8876), .B(n8922), .ZN(n8879) );
  AND2_X1 U10231 ( .A1(n9056), .A2(n8924), .ZN(n8877) );
  AOI21_X1 U10232 ( .B1(n9614), .B2(n8925), .A(n8877), .ZN(n8878) );
  NOR2_X1 U10233 ( .A1(n8879), .A2(n8878), .ZN(n9028) );
  NAND2_X1 U10234 ( .A1(n8879), .A2(n8878), .ZN(n9026) );
  AOI22_X1 U10235 ( .A1(n9609), .A2(n6226), .B1(n8925), .B2(n9172), .ZN(n8880)
         );
  XNOR2_X1 U10236 ( .A(n8880), .B(n6247), .ZN(n8917) );
  AND2_X1 U10237 ( .A1(n9172), .A2(n8924), .ZN(n8881) );
  AOI21_X1 U10238 ( .B1(n9609), .B2(n8925), .A(n8881), .ZN(n8916) );
  XNOR2_X1 U10239 ( .A(n8917), .B(n8916), .ZN(n8882) );
  XNOR2_X1 U10240 ( .A(n8915), .B(n8882), .ZN(n8887) );
  INV_X1 U10241 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8883) );
  OAI22_X1 U10242 ( .A1(n9043), .A2(n9186), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8883), .ZN(n8885) );
  OAI22_X1 U10243 ( .A1(n9156), .A2(n9046), .B1(n9045), .B2(n9149), .ZN(n8884)
         );
  AOI211_X1 U10244 ( .C1(n9609), .C2(n9050), .A(n8885), .B(n8884), .ZN(n8886)
         );
  OAI21_X1 U10245 ( .B1(n8887), .B2(n9052), .A(n8886), .ZN(P1_U3212) );
  NAND2_X1 U10246 ( .A1(n8888), .A2(n8889), .ZN(n8891) );
  XNOR2_X1 U10247 ( .A(n8891), .B(n8890), .ZN(n8892) );
  NAND2_X1 U10248 ( .A1(n8892), .A2(n8982), .ZN(n8897) );
  OAI22_X1 U10249 ( .A1(n8967), .A2(n9046), .B1(n9045), .B2(n8893), .ZN(n8894)
         );
  AOI211_X1 U10250 ( .C1(n8943), .C2(n9060), .A(n8895), .B(n8894), .ZN(n8896)
         );
  OAI211_X1 U10251 ( .C1(n9768), .C2(n9024), .A(n8897), .B(n8896), .ZN(
        P1_U3213) );
  INV_X1 U10252 ( .A(n8981), .ZN(n8901) );
  AOI21_X1 U10253 ( .B1(n8980), .B2(n8899), .A(n8898), .ZN(n8900) );
  AOI21_X1 U10254 ( .B1(n8901), .B2(n8980), .A(n8900), .ZN(n8905) );
  OAI22_X1 U10255 ( .A1(n9046), .A2(n9481), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9414), .ZN(n8903) );
  OAI22_X1 U10256 ( .A1(n9479), .A2(n9043), .B1(n9045), .B2(n9484), .ZN(n8902)
         );
  AOI211_X1 U10257 ( .C1(n9631), .C2(n9050), .A(n8903), .B(n8902), .ZN(n8904)
         );
  OAI21_X1 U10258 ( .B1(n8905), .B2(n9052), .A(n8904), .ZN(P1_U3214) );
  NOR2_X1 U10259 ( .A1(n4590), .A2(n8907), .ZN(n8908) );
  XNOR2_X1 U10260 ( .A(n8909), .B(n8908), .ZN(n8913) );
  NAND2_X1 U10261 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9126) );
  OAI21_X1 U10262 ( .B1(n9046), .B2(n9545), .A(n9126), .ZN(n8911) );
  OAI22_X1 U10263 ( .A1(n9543), .A2(n9043), .B1(n9045), .B2(n9549), .ZN(n8910)
         );
  AOI211_X1 U10264 ( .C1(n9651), .C2(n9050), .A(n8911), .B(n8910), .ZN(n8912)
         );
  OAI21_X1 U10265 ( .B1(n8913), .B2(n9052), .A(n8912), .ZN(P1_U3217) );
  NOR2_X1 U10266 ( .A1(n8917), .A2(n8916), .ZN(n8932) );
  NAND2_X1 U10267 ( .A1(n9603), .A2(n8918), .ZN(n8921) );
  OR2_X1 U10268 ( .A1(n9156), .A2(n6224), .ZN(n8920) );
  NAND2_X1 U10269 ( .A1(n8921), .A2(n8920), .ZN(n8923) );
  XNOR2_X1 U10270 ( .A(n8923), .B(n8922), .ZN(n8927) );
  AOI22_X1 U10271 ( .A1(n9603), .A2(n8925), .B1(n8924), .B2(n7695), .ZN(n8926)
         );
  XNOR2_X1 U10272 ( .A(n8927), .B(n8926), .ZN(n8933) );
  OAI22_X1 U10273 ( .A1(n9043), .A2(n9031), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8928), .ZN(n8930) );
  OAI22_X1 U10274 ( .A1(n9134), .A2(n9046), .B1(n9045), .B2(n9139), .ZN(n8929)
         );
  AOI211_X1 U10275 ( .C1(n9603), .C2(n9050), .A(n8930), .B(n8929), .ZN(n8935)
         );
  NAND3_X1 U10276 ( .A1(n8931), .A2(n8982), .A3(n8933), .ZN(n8934) );
  OAI21_X1 U10277 ( .B1(n8938), .B2(n8936), .A(n8937), .ZN(n8939) );
  NAND2_X1 U10278 ( .A1(n8939), .A2(n8982), .ZN(n8946) );
  AOI22_X1 U10279 ( .A1(n8941), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9050), .B2(
        n8940), .ZN(n8945) );
  AOI22_X1 U10280 ( .A1(n8943), .A2(n8942), .B1(n9021), .B2(n6727), .ZN(n8944)
         );
  NAND3_X1 U10281 ( .A1(n8946), .A2(n8945), .A3(n8944), .ZN(P1_U3220) );
  NAND2_X1 U10282 ( .A1(n8947), .A2(n8990), .ZN(n8948) );
  NAND2_X1 U10283 ( .A1(n8948), .A2(n8991), .ZN(n8949) );
  XOR2_X1 U10284 ( .A(n8950), .B(n8949), .Z(n8955) );
  OAI22_X1 U10285 ( .A1(n9043), .A2(n9545), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8951), .ZN(n8953) );
  OAI22_X1 U10286 ( .A1(n9479), .A2(n9046), .B1(n9045), .B2(n9511), .ZN(n8952)
         );
  AOI211_X1 U10287 ( .C1(n9640), .C2(n9050), .A(n8953), .B(n8952), .ZN(n8954)
         );
  OAI21_X1 U10288 ( .B1(n8955), .B2(n9052), .A(n8954), .ZN(P1_U3221) );
  AOI21_X1 U10289 ( .B1(n8956), .B2(n8957), .A(n4439), .ZN(n8962) );
  OAI22_X1 U10290 ( .A1(n9046), .A2(n9186), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8958), .ZN(n8960) );
  OAI22_X1 U10291 ( .A1(n9481), .A2(n9043), .B1(n9045), .B2(n9179), .ZN(n8959)
         );
  AOI211_X1 U10292 ( .C1(n9619), .C2(n9050), .A(n8960), .B(n8959), .ZN(n8961)
         );
  OAI21_X1 U10293 ( .B1(n8962), .B2(n9052), .A(n8961), .ZN(P1_U3223) );
  XOR2_X1 U10294 ( .A(n8965), .B(n8964), .Z(n8966) );
  XNOR2_X1 U10295 ( .A(n8963), .B(n8966), .ZN(n8972) );
  NAND2_X1 U10296 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9081) );
  OAI21_X1 U10297 ( .B1(n9043), .B2(n8967), .A(n9081), .ZN(n8970) );
  OAI22_X1 U10298 ( .A1(n9019), .A2(n9046), .B1(n9045), .B2(n8968), .ZN(n8969)
         );
  AOI211_X1 U10299 ( .C1(n9666), .C2(n9050), .A(n8970), .B(n8969), .ZN(n8971)
         );
  OAI21_X1 U10300 ( .B1(n8972), .B2(n9052), .A(n8971), .ZN(P1_U3224) );
  XOR2_X1 U10301 ( .A(n8973), .B(n8974), .Z(n8978) );
  NAND2_X1 U10302 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9095) );
  OAI21_X1 U10303 ( .B1(n9043), .B2(n9047), .A(n9095), .ZN(n8976) );
  OAI22_X1 U10304 ( .A1(n9543), .A2(n9046), .B1(n9045), .B2(n9579), .ZN(n8975)
         );
  AOI211_X1 U10305 ( .C1(n9659), .C2(n9050), .A(n8976), .B(n8975), .ZN(n8977)
         );
  OAI21_X1 U10306 ( .B1(n8978), .B2(n9052), .A(n8977), .ZN(P1_U3226) );
  AND3_X1 U10307 ( .A1(n8981), .A2(n8980), .A3(n8979), .ZN(n8983) );
  OAI21_X1 U10308 ( .B1(n8984), .B2(n8983), .A(n8982), .ZN(n8989) );
  NOR2_X1 U10309 ( .A1(n9046), .A2(n9032), .ZN(n8986) );
  OAI22_X1 U10310 ( .A1(n9005), .A2(n9043), .B1(n9045), .B2(n9198), .ZN(n8985)
         );
  AOI211_X1 U10311 ( .C1(P1_REG3_REG_24__SCAN_IN), .C2(P1_U3084), .A(n8986), 
        .B(n8985), .ZN(n8988) );
  OAI211_X1 U10312 ( .C1(n9625), .C2(n9024), .A(n8989), .B(n8988), .ZN(
        P1_U3227) );
  NAND2_X1 U10313 ( .A1(n8991), .A2(n8990), .ZN(n8992) );
  XNOR2_X1 U10314 ( .A(n8947), .B(n8992), .ZN(n8998) );
  OAI22_X1 U10315 ( .A1(n9046), .A2(n9007), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8993), .ZN(n8996) );
  OAI22_X1 U10316 ( .A1(n8994), .A2(n9043), .B1(n9045), .B2(n9527), .ZN(n8995)
         );
  AOI211_X1 U10317 ( .C1(n9644), .C2(n9050), .A(n8996), .B(n8995), .ZN(n8997)
         );
  OAI21_X1 U10318 ( .B1(n8998), .B2(n9052), .A(n8997), .ZN(P1_U3231) );
  AND2_X1 U10319 ( .A1(n9000), .A2(n8999), .ZN(n9001) );
  NAND2_X1 U10320 ( .A1(n8853), .A2(n9001), .ZN(n9002) );
  XOR2_X1 U10321 ( .A(n9003), .B(n9002), .Z(n9011) );
  OAI22_X1 U10322 ( .A1(n9005), .A2(n9046), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9004), .ZN(n9009) );
  INV_X1 U10323 ( .A(n9495), .ZN(n9006) );
  OAI22_X1 U10324 ( .A1(n9007), .A2(n9043), .B1(n9045), .B2(n9006), .ZN(n9008)
         );
  AOI211_X1 U10325 ( .C1(n9634), .C2(n9050), .A(n9009), .B(n9008), .ZN(n9010)
         );
  OAI21_X1 U10326 ( .B1(n9011), .B2(n9052), .A(n9010), .ZN(P1_U3233) );
  INV_X1 U10327 ( .A(n9014), .ZN(n9018) );
  AOI21_X1 U10328 ( .B1(n9014), .B2(n9013), .A(n9012), .ZN(n9015) );
  NOR2_X1 U10329 ( .A1(n9015), .A2(n9052), .ZN(n9016) );
  OAI21_X1 U10330 ( .B1(n9018), .B2(n9017), .A(n9016), .ZN(n9023) );
  AND2_X1 U10331 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9107) );
  OAI22_X1 U10332 ( .A1(n9019), .A2(n9043), .B1(n9045), .B2(n9560), .ZN(n9020)
         );
  AOI211_X1 U10333 ( .C1(n9021), .C2(n9569), .A(n9107), .B(n9020), .ZN(n9022)
         );
  OAI211_X1 U10334 ( .C1(n9563), .C2(n9024), .A(n9023), .B(n9022), .ZN(
        P1_U3236) );
  INV_X1 U10335 ( .A(n9026), .ZN(n9027) );
  NOR2_X1 U10336 ( .A1(n9028), .A2(n9027), .ZN(n9029) );
  XNOR2_X1 U10337 ( .A(n9025), .B(n9029), .ZN(n9036) );
  INV_X1 U10338 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9030) );
  OAI22_X1 U10339 ( .A1(n9046), .A2(n9031), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9030), .ZN(n9034) );
  OAI22_X1 U10340 ( .A1(n9032), .A2(n9043), .B1(n9045), .B2(n9166), .ZN(n9033)
         );
  AOI211_X1 U10341 ( .C1(n9614), .C2(n9050), .A(n9034), .B(n9033), .ZN(n9035)
         );
  OAI21_X1 U10342 ( .B1(n9036), .B2(n9052), .A(n9035), .ZN(P1_U3238) );
  NAND2_X1 U10343 ( .A1(n9037), .A2(n9038), .ZN(n9040) );
  XOR2_X1 U10344 ( .A(n9040), .B(n9039), .Z(n9053) );
  OAI21_X1 U10345 ( .B1(n9043), .B2(n9042), .A(n9041), .ZN(n9049) );
  OAI22_X1 U10346 ( .A1(n9047), .A2(n9046), .B1(n9045), .B2(n9044), .ZN(n9048)
         );
  AOI211_X1 U10347 ( .C1(n9669), .C2(n9050), .A(n9049), .B(n9048), .ZN(n9051)
         );
  OAI21_X1 U10348 ( .B1(n9053), .B2(n9052), .A(n9051), .ZN(P1_U3239) );
  MUX2_X1 U10349 ( .A(n9054), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9833), .Z(
        P1_U3585) );
  MUX2_X1 U10350 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9055), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10351 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n7695), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10352 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9172), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10353 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9056), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10354 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9196), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10355 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9057), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10356 ( .A(n9502), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9833), .Z(
        P1_U3578) );
  MUX2_X1 U10357 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9519), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10358 ( .A(n9532), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9833), .Z(
        P1_U3576) );
  MUX2_X1 U10359 ( .A(n9518), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9833), .Z(
        P1_U3575) );
  MUX2_X1 U10360 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9569), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10361 ( .A(n9583), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9833), .Z(
        P1_U3573) );
  MUX2_X1 U10362 ( .A(n9568), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9833), .Z(
        P1_U3572) );
  MUX2_X1 U10363 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9593), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10364 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9058), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10365 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9059), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10366 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9060), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10367 ( .A(n9061), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9833), .Z(
        P1_U3567) );
  MUX2_X1 U10368 ( .A(n9062), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9833), .Z(
        P1_U3566) );
  MUX2_X1 U10369 ( .A(n9063), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9833), .Z(
        P1_U3565) );
  MUX2_X1 U10370 ( .A(n9064), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9833), .Z(
        P1_U3564) );
  MUX2_X1 U10371 ( .A(n9065), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9833), .Z(
        P1_U3563) );
  MUX2_X1 U10372 ( .A(n9066), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9833), .Z(
        P1_U3562) );
  MUX2_X1 U10373 ( .A(n9067), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9833), .Z(
        P1_U3561) );
  MUX2_X1 U10374 ( .A(n9068), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9833), .Z(
        P1_U3560) );
  MUX2_X1 U10375 ( .A(n9912), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9833), .Z(
        P1_U3559) );
  MUX2_X1 U10376 ( .A(n6866), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9833), .Z(
        P1_U3558) );
  MUX2_X1 U10377 ( .A(n6727), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9833), .Z(
        P1_U3557) );
  MUX2_X1 U10378 ( .A(n6723), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9833), .Z(
        P1_U3556) );
  NOR2_X1 U10379 ( .A1(n9069), .A2(n9076), .ZN(n9071) );
  NAND2_X1 U10380 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9092), .ZN(n9072) );
  OAI21_X1 U10381 ( .B1(n9092), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9072), .ZN(
        n9073) );
  AOI211_X1 U10382 ( .C1(n9074), .C2(n9073), .A(n9087), .B(n9827), .ZN(n9086)
         );
  NOR2_X1 U10383 ( .A1(n9076), .A2(n9075), .ZN(n9078) );
  NOR2_X1 U10384 ( .A1(n9078), .A2(n9077), .ZN(n9080) );
  XNOR2_X1 U10385 ( .A(n9092), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9079) );
  NOR2_X1 U10386 ( .A1(n9080), .A2(n9079), .ZN(n9091) );
  AOI211_X1 U10387 ( .C1(n9080), .C2(n9079), .A(n9091), .B(n9896), .ZN(n9085)
         );
  INV_X1 U10388 ( .A(n9880), .ZN(n9900) );
  NAND2_X1 U10389 ( .A1(n9900), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9082) );
  OAI211_X1 U10390 ( .C1(n9818), .C2(n9083), .A(n9082), .B(n9081), .ZN(n9084)
         );
  OR3_X1 U10391 ( .A1(n9086), .A2(n9085), .A3(n9084), .ZN(P1_U3257) );
  INV_X1 U10392 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U10393 ( .A1(n9109), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9088) );
  OAI21_X1 U10394 ( .B1(n9109), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9088), .ZN(
        n9089) );
  NOR2_X1 U10395 ( .A1(n9090), .A2(n9089), .ZN(n9102) );
  AOI211_X1 U10396 ( .C1(n9090), .C2(n9089), .A(n9102), .B(n9827), .ZN(n9099)
         );
  AOI21_X1 U10397 ( .B1(n9092), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9091), .ZN(
        n9094) );
  XNOR2_X1 U10398 ( .A(n9109), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9093) );
  NOR2_X1 U10399 ( .A1(n9094), .A2(n9093), .ZN(n9108) );
  AOI211_X1 U10400 ( .C1(n9094), .C2(n9093), .A(n9108), .B(n9896), .ZN(n9098)
         );
  INV_X1 U10401 ( .A(n9109), .ZN(n9096) );
  OAI21_X1 U10402 ( .B1(n9818), .B2(n9096), .A(n9095), .ZN(n9097) );
  NOR3_X1 U10403 ( .A1(n9099), .A2(n9098), .A3(n9097), .ZN(n9100) );
  OAI21_X1 U10404 ( .B1(n9880), .B2(n9101), .A(n9100), .ZN(P1_U3258) );
  INV_X1 U10405 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9115) );
  NAND2_X1 U10406 ( .A1(n9119), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9103) );
  OAI21_X1 U10407 ( .B1(n9119), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9103), .ZN(
        n9104) );
  AOI211_X1 U10408 ( .C1(n9105), .C2(n9104), .A(n9118), .B(n9827), .ZN(n9106)
         );
  AOI211_X1 U10409 ( .C1(n9119), .C2(n9898), .A(n9107), .B(n9106), .ZN(n9114)
         );
  XNOR2_X1 U10410 ( .A(n9119), .B(n9286), .ZN(n9111) );
  AOI21_X1 U10411 ( .B1(n9109), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9108), .ZN(
        n9110) );
  NAND2_X1 U10412 ( .A1(n9111), .A2(n9110), .ZN(n9116) );
  OAI21_X1 U10413 ( .B1(n9111), .B2(n9110), .A(n9116), .ZN(n9112) );
  NAND2_X1 U10414 ( .A1(n9872), .A2(n9112), .ZN(n9113) );
  OAI211_X1 U10415 ( .C1(n9880), .C2(n9115), .A(n9114), .B(n9113), .ZN(
        P1_U3259) );
  OAI21_X1 U10416 ( .B1(n9119), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9116), .ZN(
        n9117) );
  XNOR2_X1 U10417 ( .A(n9117), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9121) );
  NAND2_X1 U10418 ( .A1(n9123), .A2(n9891), .ZN(n9120) );
  INV_X1 U10419 ( .A(n9121), .ZN(n9122) );
  OAI22_X1 U10420 ( .A1(n9123), .A2(n9827), .B1(n9896), .B2(n9122), .ZN(n9125)
         );
  XNOR2_X1 U10421 ( .A(n9128), .B(n9127), .ZN(n9765) );
  NAND2_X1 U10422 ( .A1(n9765), .A2(n9909), .ZN(n9131) );
  AOI21_X1 U10423 ( .B1(n4382), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9129), .ZN(
        n9130) );
  OAI211_X1 U10424 ( .C1(n9763), .C2(n9930), .A(n9131), .B(n9130), .ZN(
        P1_U3262) );
  OAI21_X1 U10425 ( .B1(n9133), .B2(n9136), .A(n9132), .ZN(n9607) );
  NOR2_X1 U10426 ( .A1(n9134), .A2(n9546), .ZN(n9138) );
  OAI21_X1 U10427 ( .B1(n9139), .B2(n9936), .A(n9606), .ZN(n9140) );
  NAND2_X1 U10428 ( .A1(n9140), .A2(n9926), .ZN(n9146) );
  AOI21_X1 U10429 ( .B1(n9603), .B2(n9148), .A(n9141), .ZN(n9604) );
  OAI22_X1 U10430 ( .A1(n9143), .A2(n9930), .B1(n9142), .B2(n9926), .ZN(n9144)
         );
  AOI21_X1 U10431 ( .B1(n9604), .B2(n9909), .A(n9144), .ZN(n9145) );
  OAI211_X1 U10432 ( .C1(n9607), .C2(n9597), .A(n9146), .B(n9145), .ZN(
        P1_U3263) );
  XOR2_X1 U10433 ( .A(n9147), .B(n9155), .Z(n9612) );
  AOI211_X1 U10434 ( .C1(n9609), .C2(n9163), .A(n10029), .B(n4512), .ZN(n9608)
         );
  INV_X1 U10435 ( .A(n9609), .ZN(n9152) );
  INV_X1 U10436 ( .A(n9149), .ZN(n9150) );
  AOI22_X1 U10437 ( .A1(n4382), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9150), .B2(
        n9923), .ZN(n9151) );
  OAI21_X1 U10438 ( .B1(n9152), .B2(n9930), .A(n9151), .ZN(n9160) );
  AOI211_X1 U10439 ( .C1(n9155), .C2(n9154), .A(n9588), .B(n9153), .ZN(n9158)
         );
  OAI22_X1 U10440 ( .A1(n9186), .A2(n9544), .B1(n9156), .B2(n9546), .ZN(n9157)
         );
  NOR2_X1 U10441 ( .A1(n9158), .A2(n9157), .ZN(n9611) );
  NOR2_X1 U10442 ( .A1(n9611), .A2(n4382), .ZN(n9159) );
  AOI211_X1 U10443 ( .C1(n9573), .C2(n9608), .A(n9160), .B(n9159), .ZN(n9161)
         );
  OAI21_X1 U10444 ( .B1(n9612), .B2(n9597), .A(n9161), .ZN(P1_U3264) );
  XOR2_X1 U10445 ( .A(n9171), .B(n9162), .Z(n9617) );
  INV_X1 U10446 ( .A(n9178), .ZN(n9165) );
  INV_X1 U10447 ( .A(n9163), .ZN(n9164) );
  AOI211_X1 U10448 ( .C1(n9614), .C2(n9165), .A(n10029), .B(n9164), .ZN(n9613)
         );
  INV_X1 U10449 ( .A(n9166), .ZN(n9167) );
  AOI22_X1 U10450 ( .A1(n4382), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9167), .B2(
        n9923), .ZN(n9168) );
  OAI21_X1 U10451 ( .B1(n9169), .B2(n9930), .A(n9168), .ZN(n9175) );
  OAI21_X1 U10452 ( .B1(n4463), .B2(n9171), .A(n9170), .ZN(n9173) );
  AOI222_X1 U10453 ( .A1(n9916), .A2(n9173), .B1(n9172), .B2(n9911), .C1(n9196), .C2(n9913), .ZN(n9616) );
  NOR2_X1 U10454 ( .A1(n9616), .A2(n4382), .ZN(n9174) );
  AOI211_X1 U10455 ( .C1(n9613), .C2(n9573), .A(n9175), .B(n9174), .ZN(n9176)
         );
  OAI21_X1 U10456 ( .B1(n9617), .B2(n9597), .A(n9176), .ZN(P1_U3265) );
  XOR2_X1 U10457 ( .A(n9177), .B(n9185), .Z(n9622) );
  AOI211_X1 U10458 ( .C1(n9619), .C2(n4414), .A(n10029), .B(n9178), .ZN(n9618)
         );
  INV_X1 U10459 ( .A(n9179), .ZN(n9180) );
  AOI22_X1 U10460 ( .A1(n4382), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9180), .B2(
        n9923), .ZN(n9181) );
  OAI21_X1 U10461 ( .B1(n9182), .B2(n9930), .A(n9181), .ZN(n9190) );
  AOI211_X1 U10462 ( .C1(n9185), .C2(n9184), .A(n9588), .B(n9183), .ZN(n9188)
         );
  OAI22_X1 U10463 ( .A1(n9481), .A2(n9544), .B1(n9186), .B2(n9546), .ZN(n9187)
         );
  NOR2_X1 U10464 ( .A1(n9188), .A2(n9187), .ZN(n9621) );
  NOR2_X1 U10465 ( .A1(n9621), .A2(n4382), .ZN(n9189) );
  AOI211_X1 U10466 ( .C1(n9618), .C2(n9573), .A(n9190), .B(n9189), .ZN(n9191)
         );
  OAI21_X1 U10467 ( .B1(n9622), .B2(n9597), .A(n9191), .ZN(P1_U3266) );
  XOR2_X1 U10468 ( .A(n9192), .B(n9194), .Z(n9627) );
  INV_X1 U10469 ( .A(n9193), .ZN(n9482) );
  OAI211_X1 U10470 ( .C1(n9625), .C2(n9482), .A(n10005), .B(n4414), .ZN(n9623)
         );
  XNOR2_X1 U10471 ( .A(n9195), .B(n9194), .ZN(n9197) );
  AOI222_X1 U10472 ( .A1(n9916), .A2(n9197), .B1(n9196), .B2(n9911), .C1(n9502), .C2(n9913), .ZN(n9624) );
  OAI21_X1 U10473 ( .B1(n9936), .B2(n9198), .A(n9926), .ZN(n9199) );
  AOI21_X1 U10474 ( .B1(n9201), .B2(n9200), .A(n9199), .ZN(n9202) );
  OAI211_X1 U10475 ( .C1(n9203), .C2(n9623), .A(n9624), .B(n9202), .ZN(n9204)
         );
  AOI21_X1 U10476 ( .B1(n9627), .B2(n9205), .A(n9204), .ZN(n9206) );
  AOI21_X1 U10477 ( .B1(n4382), .B2(n9207), .A(n9206), .ZN(n9475) );
  AOI22_X1 U10478 ( .A1(n9938), .A2(keyinput49), .B1(keyinput10), .B2(n9209), 
        .ZN(n9208) );
  OAI221_X1 U10479 ( .B1(n9938), .B2(keyinput49), .C1(n9209), .C2(keyinput10), 
        .A(n9208), .ZN(n9218) );
  AOI22_X1 U10480 ( .A1(n9427), .A2(keyinput7), .B1(keyinput34), .B2(n9211), 
        .ZN(n9210) );
  OAI221_X1 U10481 ( .B1(n9427), .B2(keyinput7), .C1(n9211), .C2(keyinput34), 
        .A(n9210), .ZN(n9217) );
  INV_X1 U10482 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n9958) );
  AOI22_X1 U10483 ( .A1(n9958), .A2(keyinput61), .B1(keyinput6), .B2(n9213), 
        .ZN(n9212) );
  OAI221_X1 U10484 ( .B1(n9958), .B2(keyinput61), .C1(n9213), .C2(keyinput6), 
        .A(n9212), .ZN(n9216) );
  AOI22_X1 U10485 ( .A1(n6995), .A2(keyinput57), .B1(keyinput126), .B2(n7090), 
        .ZN(n9214) );
  OAI221_X1 U10486 ( .B1(n6995), .B2(keyinput57), .C1(n7090), .C2(keyinput126), 
        .A(n9214), .ZN(n9215) );
  NOR4_X1 U10487 ( .A1(n9218), .A2(n9217), .A3(n9216), .A4(n9215), .ZN(n9236)
         );
  INV_X1 U10488 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9881) );
  AOI22_X1 U10489 ( .A1(n4615), .A2(keyinput82), .B1(keyinput114), .B2(n9881), 
        .ZN(n9219) );
  OAI221_X1 U10490 ( .B1(n4615), .B2(keyinput82), .C1(n9881), .C2(keyinput114), 
        .A(n9219), .ZN(n9227) );
  AOI22_X1 U10491 ( .A1(n9222), .A2(keyinput29), .B1(keyinput74), .B2(n9221), 
        .ZN(n9220) );
  OAI221_X1 U10492 ( .B1(n9222), .B2(keyinput29), .C1(n9221), .C2(keyinput74), 
        .A(n9220), .ZN(n9226) );
  INV_X1 U10493 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9224) );
  INV_X1 U10494 ( .A(SI_3_), .ZN(n9406) );
  AOI22_X1 U10495 ( .A1(n9224), .A2(keyinput68), .B1(n9406), .B2(keyinput8), 
        .ZN(n9223) );
  OAI221_X1 U10496 ( .B1(n9224), .B2(keyinput68), .C1(n9406), .C2(keyinput8), 
        .A(n9223), .ZN(n9225) );
  NOR3_X1 U10497 ( .A1(n9227), .A2(n9226), .A3(n9225), .ZN(n9235) );
  AOI22_X1 U10498 ( .A1(n9229), .A2(keyinput1), .B1(keyinput71), .B2(n10229), 
        .ZN(n9228) );
  OAI221_X1 U10499 ( .B1(n9229), .B2(keyinput1), .C1(n10229), .C2(keyinput71), 
        .A(n9228), .ZN(n9233) );
  INV_X1 U10500 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U10501 ( .A1(n9231), .A2(keyinput43), .B1(keyinput27), .B2(n10184), 
        .ZN(n9230) );
  OAI221_X1 U10502 ( .B1(n9231), .B2(keyinput43), .C1(n10184), .C2(keyinput27), 
        .A(n9230), .ZN(n9232) );
  NOR2_X1 U10503 ( .A1(n9233), .A2(n9232), .ZN(n9234) );
  NAND3_X1 U10504 ( .A1(n9236), .A2(n9235), .A3(n9234), .ZN(n9320) );
  INV_X1 U10505 ( .A(keyinput44), .ZN(n9238) );
  AOI22_X1 U10506 ( .A1(n9784), .A2(keyinput113), .B1(P2_WR_REG_SCAN_IN), .B2(
        n9238), .ZN(n9237) );
  OAI221_X1 U10507 ( .B1(n9784), .B2(keyinput113), .C1(n9238), .C2(
        P2_WR_REG_SCAN_IN), .A(n9237), .ZN(n9248) );
  AOI22_X1 U10508 ( .A1(n9403), .A2(keyinput108), .B1(n9240), .B2(keyinput64), 
        .ZN(n9239) );
  OAI221_X1 U10509 ( .B1(n9403), .B2(keyinput108), .C1(n9240), .C2(keyinput64), 
        .A(n9239), .ZN(n9247) );
  AOI22_X1 U10510 ( .A1(n9242), .A2(keyinput93), .B1(n5171), .B2(keyinput104), 
        .ZN(n9241) );
  OAI221_X1 U10511 ( .B1(n9242), .B2(keyinput93), .C1(n5171), .C2(keyinput104), 
        .A(n9241), .ZN(n9246) );
  AOI22_X1 U10512 ( .A1(n5999), .A2(keyinput86), .B1(n9244), .B2(keyinput55), 
        .ZN(n9243) );
  OAI221_X1 U10513 ( .B1(n5999), .B2(keyinput86), .C1(n9244), .C2(keyinput55), 
        .A(n9243), .ZN(n9245) );
  NOR4_X1 U10514 ( .A1(n9248), .A2(n9247), .A3(n9246), .A4(n9245), .ZN(n9251)
         );
  INV_X1 U10515 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9940) );
  XOR2_X1 U10516 ( .A(keyinput9), .B(n9940), .Z(n9250) );
  INV_X1 U10517 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9949) );
  XOR2_X1 U10518 ( .A(keyinput90), .B(n9949), .Z(n9249) );
  NAND3_X1 U10519 ( .A1(n9251), .A2(n9250), .A3(n9249), .ZN(n9319) );
  AOI22_X1 U10520 ( .A1(n6748), .A2(keyinput69), .B1(keyinput70), .B2(n9253), 
        .ZN(n9252) );
  OAI221_X1 U10521 ( .B1(n6748), .B2(keyinput69), .C1(n9253), .C2(keyinput70), 
        .A(n9252), .ZN(n9256) );
  AOI22_X1 U10522 ( .A1(n10084), .A2(keyinput50), .B1(n9440), .B2(keyinput99), 
        .ZN(n9254) );
  OAI221_X1 U10523 ( .B1(n10084), .B2(keyinput50), .C1(n9440), .C2(keyinput99), 
        .A(n9254), .ZN(n9255) );
  NOR2_X1 U10524 ( .A1(n9256), .A2(n9255), .ZN(n9284) );
  AOI22_X1 U10525 ( .A1(n6185), .A2(keyinput17), .B1(n9425), .B2(keyinput47), 
        .ZN(n9257) );
  OAI221_X1 U10526 ( .B1(n6185), .B2(keyinput17), .C1(n9425), .C2(keyinput47), 
        .A(n9257), .ZN(n9263) );
  XNOR2_X1 U10527 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput105), .ZN(n9261) );
  XNOR2_X1 U10528 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput77), .ZN(n9260) );
  XNOR2_X1 U10529 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput53), .ZN(n9259) );
  XNOR2_X1 U10530 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput78), .ZN(n9258) );
  NAND4_X1 U10531 ( .A1(n9261), .A2(n9260), .A3(n9259), .A4(n9258), .ZN(n9262)
         );
  NOR2_X1 U10532 ( .A1(n9263), .A2(n9262), .ZN(n9283) );
  XNOR2_X1 U10533 ( .A(SI_21_), .B(keyinput4), .ZN(n9267) );
  XNOR2_X1 U10534 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput81), .ZN(n9266) );
  XNOR2_X1 U10535 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput2), .ZN(n9265) );
  XNOR2_X1 U10536 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput38), .ZN(n9264) );
  NAND4_X1 U10537 ( .A1(n9267), .A2(n9266), .A3(n9265), .A4(n9264), .ZN(n9273)
         );
  XNOR2_X1 U10538 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput84), .ZN(n9271) );
  XNOR2_X1 U10539 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput124), .ZN(n9270)
         );
  XNOR2_X1 U10540 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput79), .ZN(n9269) );
  XNOR2_X1 U10541 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput94), .ZN(n9268) );
  NAND4_X1 U10542 ( .A1(n9271), .A2(n9270), .A3(n9269), .A4(n9268), .ZN(n9272)
         );
  NOR2_X1 U10543 ( .A1(n9273), .A2(n9272), .ZN(n9282) );
  AOI22_X1 U10544 ( .A1(n9965), .A2(keyinput36), .B1(keyinput122), .B2(n9461), 
        .ZN(n9274) );
  OAI221_X1 U10545 ( .B1(n9965), .B2(keyinput36), .C1(n9461), .C2(keyinput122), 
        .A(n9274), .ZN(n9280) );
  XNOR2_X1 U10546 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput41), .ZN(n9278) );
  XNOR2_X1 U10547 ( .A(P2_IR_REG_27__SCAN_IN), .B(keyinput80), .ZN(n9277) );
  XNOR2_X1 U10548 ( .A(keyinput60), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n9276) );
  XNOR2_X1 U10549 ( .A(keyinput120), .B(P1_REG3_REG_7__SCAN_IN), .ZN(n9275) );
  NAND4_X1 U10550 ( .A1(n9278), .A2(n9277), .A3(n9276), .A4(n9275), .ZN(n9279)
         );
  NOR2_X1 U10551 ( .A1(n9280), .A2(n9279), .ZN(n9281) );
  NAND4_X1 U10552 ( .A1(n9284), .A2(n9283), .A3(n9282), .A4(n9281), .ZN(n9318)
         );
  AOI22_X1 U10553 ( .A1(n9286), .A2(keyinput30), .B1(keyinput125), .B2(n6110), 
        .ZN(n9285) );
  OAI221_X1 U10554 ( .B1(n9286), .B2(keyinput30), .C1(n6110), .C2(keyinput125), 
        .A(n9285), .ZN(n9293) );
  AOI22_X1 U10555 ( .A1(n9289), .A2(keyinput83), .B1(n9288), .B2(keyinput72), 
        .ZN(n9287) );
  OAI221_X1 U10556 ( .B1(n9289), .B2(keyinput83), .C1(n9288), .C2(keyinput72), 
        .A(n9287), .ZN(n9292) );
  XNOR2_X1 U10557 ( .A(keyinput14), .B(n5324), .ZN(n9291) );
  XNOR2_X1 U10558 ( .A(keyinput42), .B(n5142), .ZN(n9290) );
  NOR4_X1 U10559 ( .A1(n9293), .A2(n9292), .A3(n9291), .A4(n9290), .ZN(n9316)
         );
  INV_X1 U10560 ( .A(SI_30_), .ZN(n9295) );
  AOI22_X1 U10561 ( .A1(n9296), .A2(keyinput67), .B1(keyinput96), .B2(n9295), 
        .ZN(n9294) );
  OAI221_X1 U10562 ( .B1(n9296), .B2(keyinput67), .C1(n9295), .C2(keyinput96), 
        .A(n9294), .ZN(n9299) );
  INV_X1 U10563 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10087) );
  AOI22_X1 U10564 ( .A1(n9718), .A2(keyinput121), .B1(n10087), .B2(keyinput0), 
        .ZN(n9297) );
  OAI221_X1 U10565 ( .B1(n9718), .B2(keyinput121), .C1(n10087), .C2(keyinput0), 
        .A(n9297), .ZN(n9298) );
  NOR2_X1 U10566 ( .A1(n9299), .A2(n9298), .ZN(n9315) );
  AOI22_X1 U10567 ( .A1(n9460), .A2(keyinput106), .B1(keyinput127), .B2(n6202), 
        .ZN(n9300) );
  OAI221_X1 U10568 ( .B1(n9460), .B2(keyinput106), .C1(n6202), .C2(keyinput127), .A(n9300), .ZN(n9308) );
  AOI22_X1 U10569 ( .A1(n9422), .A2(keyinput109), .B1(n9302), .B2(keyinput62), 
        .ZN(n9301) );
  OAI221_X1 U10570 ( .B1(n9422), .B2(keyinput109), .C1(n9302), .C2(keyinput62), 
        .A(n9301), .ZN(n9307) );
  AOI22_X1 U10571 ( .A1(n9305), .A2(keyinput115), .B1(n9304), .B2(keyinput35), 
        .ZN(n9303) );
  OAI221_X1 U10572 ( .B1(n9305), .B2(keyinput115), .C1(n9304), .C2(keyinput35), 
        .A(n9303), .ZN(n9306) );
  NOR3_X1 U10573 ( .A1(n9308), .A2(n9307), .A3(n9306), .ZN(n9314) );
  AOI22_X1 U10574 ( .A1(n9409), .A2(keyinput123), .B1(keyinput76), .B2(n5967), 
        .ZN(n9309) );
  OAI221_X1 U10575 ( .B1(n9409), .B2(keyinput123), .C1(n5967), .C2(keyinput76), 
        .A(n9309), .ZN(n9312) );
  AOI22_X1 U10576 ( .A1(n6098), .A2(keyinput22), .B1(keyinput97), .B2(n6102), 
        .ZN(n9310) );
  OAI221_X1 U10577 ( .B1(n6098), .B2(keyinput22), .C1(n6102), .C2(keyinput97), 
        .A(n9310), .ZN(n9311) );
  NOR2_X1 U10578 ( .A1(n9312), .A2(n9311), .ZN(n9313) );
  NAND4_X1 U10579 ( .A1(n9316), .A2(n9315), .A3(n9314), .A4(n9313), .ZN(n9317)
         );
  NOR4_X1 U10580 ( .A1(n9320), .A2(n9319), .A3(n9318), .A4(n9317), .ZN(n9355)
         );
  AOI22_X1 U10581 ( .A1(n8484), .A2(keyinput52), .B1(n9322), .B2(keyinput66), 
        .ZN(n9321) );
  OAI221_X1 U10582 ( .B1(n8484), .B2(keyinput52), .C1(n9322), .C2(keyinput66), 
        .A(n9321), .ZN(n9333) );
  INV_X1 U10583 ( .A(P1_RD_REG_SCAN_IN), .ZN(n9799) );
  AOI22_X1 U10584 ( .A1(n9799), .A2(keyinput54), .B1(keyinput39), .B2(n9324), 
        .ZN(n9323) );
  OAI221_X1 U10585 ( .B1(n9799), .B2(keyinput54), .C1(n9324), .C2(keyinput39), 
        .A(n9323), .ZN(n9332) );
  AOI22_X1 U10586 ( .A1(n9426), .A2(keyinput20), .B1(n9326), .B2(keyinput110), 
        .ZN(n9325) );
  OAI221_X1 U10587 ( .B1(n9426), .B2(keyinput20), .C1(n9326), .C2(keyinput110), 
        .A(n9325), .ZN(n9331) );
  AOI22_X1 U10588 ( .A1(n9329), .A2(keyinput107), .B1(keyinput100), .B2(n9328), 
        .ZN(n9327) );
  OAI221_X1 U10589 ( .B1(n9329), .B2(keyinput107), .C1(n9328), .C2(keyinput100), .A(n9327), .ZN(n9330) );
  NOR4_X1 U10590 ( .A1(n9333), .A2(n9332), .A3(n9331), .A4(n9330), .ZN(n9354)
         );
  AOI22_X1 U10591 ( .A1(n9464), .A2(keyinput45), .B1(n5269), .B2(keyinput46), 
        .ZN(n9334) );
  OAI221_X1 U10592 ( .B1(n9464), .B2(keyinput45), .C1(n5269), .C2(keyinput46), 
        .A(n9334), .ZN(n9341) );
  AOI22_X1 U10593 ( .A1(n9465), .A2(keyinput25), .B1(n9454), .B2(keyinput87), 
        .ZN(n9335) );
  OAI221_X1 U10594 ( .B1(n9465), .B2(keyinput25), .C1(n9454), .C2(keyinput87), 
        .A(n9335), .ZN(n9340) );
  AOI22_X1 U10595 ( .A1(n9453), .A2(keyinput13), .B1(keyinput51), .B2(n5193), 
        .ZN(n9336) );
  OAI221_X1 U10596 ( .B1(n9453), .B2(keyinput13), .C1(n5193), .C2(keyinput51), 
        .A(n9336), .ZN(n9339) );
  AOI22_X1 U10597 ( .A1(n5220), .A2(keyinput117), .B1(n9946), .B2(keyinput26), 
        .ZN(n9337) );
  OAI221_X1 U10598 ( .B1(n5220), .B2(keyinput117), .C1(n9946), .C2(keyinput26), 
        .A(n9337), .ZN(n9338) );
  NOR4_X1 U10599 ( .A1(n9341), .A2(n9340), .A3(n9339), .A4(n9338), .ZN(n9353)
         );
  AOI22_X1 U10600 ( .A1(n9771), .A2(keyinput92), .B1(n9448), .B2(keyinput118), 
        .ZN(n9342) );
  OAI221_X1 U10601 ( .B1(n9771), .B2(keyinput92), .C1(n9448), .C2(keyinput118), 
        .A(n9342), .ZN(n9351) );
  INV_X1 U10602 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10086) );
  AOI22_X1 U10603 ( .A1(n10086), .A2(keyinput23), .B1(n9344), .B2(keyinput65), 
        .ZN(n9343) );
  OAI221_X1 U10604 ( .B1(n10086), .B2(keyinput23), .C1(n9344), .C2(keyinput65), 
        .A(n9343), .ZN(n9350) );
  INV_X1 U10605 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9941) );
  AOI22_X1 U10606 ( .A1(n9414), .A2(keyinput95), .B1(n9941), .B2(keyinput18), 
        .ZN(n9345) );
  OAI221_X1 U10607 ( .B1(n9414), .B2(keyinput95), .C1(n9941), .C2(keyinput18), 
        .A(n9345), .ZN(n9349) );
  INV_X1 U10608 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n9347) );
  INV_X1 U10609 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n9937) );
  AOI22_X1 U10610 ( .A1(n9347), .A2(keyinput3), .B1(n9937), .B2(keyinput116), 
        .ZN(n9346) );
  OAI221_X1 U10611 ( .B1(n9347), .B2(keyinput3), .C1(n9937), .C2(keyinput116), 
        .A(n9346), .ZN(n9348) );
  NOR4_X1 U10612 ( .A1(n9351), .A2(n9350), .A3(n9349), .A4(n9348), .ZN(n9352)
         );
  NAND4_X1 U10613 ( .A1(n9355), .A2(n9354), .A3(n9353), .A4(n9352), .ZN(n9401)
         );
  AOI22_X1 U10614 ( .A1(n7198), .A2(keyinput85), .B1(keyinput16), .B2(n10054), 
        .ZN(n9356) );
  OAI221_X1 U10615 ( .B1(n7198), .B2(keyinput85), .C1(n10054), .C2(keyinput16), 
        .A(n9356), .ZN(n9364) );
  AOI22_X1 U10616 ( .A1(n10083), .A2(keyinput103), .B1(n9358), .B2(keyinput58), 
        .ZN(n9357) );
  OAI221_X1 U10617 ( .B1(n10083), .B2(keyinput103), .C1(n9358), .C2(keyinput58), .A(n9357), .ZN(n9363) );
  INV_X1 U10618 ( .A(P2_RD_REG_SCAN_IN), .ZN(n9798) );
  AOI22_X1 U10619 ( .A1(n9798), .A2(keyinput11), .B1(keyinput112), .B2(n10211), 
        .ZN(n9359) );
  OAI221_X1 U10620 ( .B1(n9798), .B2(keyinput11), .C1(n10211), .C2(keyinput112), .A(n9359), .ZN(n9362) );
  AOI22_X1 U10621 ( .A1(n9452), .A2(keyinput31), .B1(keyinput15), .B2(n9459), 
        .ZN(n9360) );
  OAI221_X1 U10622 ( .B1(n9452), .B2(keyinput31), .C1(n9459), .C2(keyinput15), 
        .A(n9360), .ZN(n9361) );
  NOR4_X1 U10623 ( .A1(n9364), .A2(n9363), .A3(n9362), .A4(n9361), .ZN(n9399)
         );
  INV_X1 U10624 ( .A(SI_14_), .ZN(n9441) );
  AOI22_X1 U10625 ( .A1(n5213), .A2(keyinput12), .B1(n9441), .B2(keyinput101), 
        .ZN(n9365) );
  OAI221_X1 U10626 ( .B1(n5213), .B2(keyinput12), .C1(n9441), .C2(keyinput101), 
        .A(n9365), .ZN(n9374) );
  INV_X1 U10627 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9368) );
  AOI22_X1 U10628 ( .A1(n9368), .A2(keyinput28), .B1(keyinput19), .B2(n9367), 
        .ZN(n9366) );
  OAI221_X1 U10629 ( .B1(n9368), .B2(keyinput28), .C1(n9367), .C2(keyinput19), 
        .A(n9366), .ZN(n9373) );
  AOI22_X1 U10630 ( .A1(n10082), .A2(keyinput73), .B1(keyinput33), .B2(n9421), 
        .ZN(n9369) );
  OAI221_X1 U10631 ( .B1(n10082), .B2(keyinput73), .C1(n9421), .C2(keyinput33), 
        .A(n9369), .ZN(n9372) );
  INV_X1 U10632 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9439) );
  AOI22_X1 U10633 ( .A1(n5684), .A2(keyinput37), .B1(keyinput24), .B2(n9439), 
        .ZN(n9370) );
  OAI221_X1 U10634 ( .B1(n5684), .B2(keyinput37), .C1(n9439), .C2(keyinput24), 
        .A(n9370), .ZN(n9371) );
  NOR4_X1 U10635 ( .A1(n9374), .A2(n9373), .A3(n9372), .A4(n9371), .ZN(n9398)
         );
  AOI22_X1 U10636 ( .A1(n10085), .A2(keyinput32), .B1(n9376), .B2(keyinput119), 
        .ZN(n9375) );
  OAI221_X1 U10637 ( .B1(n10085), .B2(keyinput32), .C1(n9376), .C2(keyinput119), .A(n9375), .ZN(n9384) );
  AOI22_X1 U10638 ( .A1(n9378), .A2(keyinput59), .B1(n10089), .B2(keyinput88), 
        .ZN(n9377) );
  OAI221_X1 U10639 ( .B1(n9378), .B2(keyinput59), .C1(n10089), .C2(keyinput88), 
        .A(n9377), .ZN(n9383) );
  INV_X1 U10640 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n9423) );
  AOI22_X1 U10641 ( .A1(P1_U3084), .A2(keyinput40), .B1(keyinput75), .B2(n9423), .ZN(n9379) );
  OAI221_X1 U10642 ( .B1(P1_U3084), .B2(keyinput40), .C1(n9423), .C2(
        keyinput75), .A(n9379), .ZN(n9382) );
  INV_X1 U10643 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9964) );
  AOI22_X1 U10644 ( .A1(n9964), .A2(keyinput21), .B1(keyinput5), .B2(n6958), 
        .ZN(n9380) );
  OAI221_X1 U10645 ( .B1(n9964), .B2(keyinput21), .C1(n6958), .C2(keyinput5), 
        .A(n9380), .ZN(n9381) );
  NOR4_X1 U10646 ( .A1(n9384), .A2(n9383), .A3(n9382), .A4(n9381), .ZN(n9397)
         );
  AOI22_X1 U10647 ( .A1(n9386), .A2(keyinput48), .B1(keyinput56), .B2(n5246), 
        .ZN(n9385) );
  OAI221_X1 U10648 ( .B1(n9386), .B2(keyinput48), .C1(n5246), .C2(keyinput56), 
        .A(n9385), .ZN(n9395) );
  AOI22_X1 U10649 ( .A1(n9388), .A2(keyinput98), .B1(keyinput63), .B2(n6821), 
        .ZN(n9387) );
  OAI221_X1 U10650 ( .B1(n9388), .B2(keyinput98), .C1(n6821), .C2(keyinput63), 
        .A(n9387), .ZN(n9394) );
  AOI22_X1 U10651 ( .A1(n9142), .A2(keyinput89), .B1(keyinput102), .B2(n9390), 
        .ZN(n9389) );
  OAI221_X1 U10652 ( .B1(n9142), .B2(keyinput89), .C1(n9390), .C2(keyinput102), 
        .A(n9389), .ZN(n9393) );
  AOI22_X1 U10653 ( .A1(n9415), .A2(keyinput111), .B1(n6639), .B2(keyinput91), 
        .ZN(n9391) );
  OAI221_X1 U10654 ( .B1(n9415), .B2(keyinput111), .C1(n6639), .C2(keyinput91), 
        .A(n9391), .ZN(n9392) );
  NOR4_X1 U10655 ( .A1(n9395), .A2(n9394), .A3(n9393), .A4(n9392), .ZN(n9396)
         );
  NAND4_X1 U10656 ( .A1(n9399), .A2(n9398), .A3(n9397), .A4(n9396), .ZN(n9400)
         );
  NOR2_X1 U10657 ( .A1(n9401), .A2(n9400), .ZN(n9473) );
  NOR4_X1 U10658 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(P1_REG1_REG_10__SCAN_IN), 
        .A3(P1_REG2_REG_8__SCAN_IN), .A4(n6748), .ZN(n9402) );
  NAND3_X1 U10659 ( .A1(P1_REG1_REG_14__SCAN_IN), .A2(P1_REG2_REG_12__SCAN_IN), 
        .A3(n9402), .ZN(n9419) );
  NAND4_X1 U10660 ( .A1(P1_REG2_REG_22__SCAN_IN), .A2(P1_REG1_REG_18__SCAN_IN), 
        .A3(P1_REG0_REG_18__SCAN_IN), .A4(n9403), .ZN(n9404) );
  NOR3_X1 U10661 ( .A1(P1_REG1_REG_17__SCAN_IN), .A2(P1_REG0_REG_16__SCAN_IN), 
        .A3(n9404), .ZN(n9417) );
  NOR4_X1 U10662 ( .A1(n9407), .A2(n9406), .A3(n9405), .A4(
        P1_IR_REG_22__SCAN_IN), .ZN(n9411) );
  NAND4_X1 U10663 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), 
        .A3(P1_IR_REG_29__SCAN_IN), .A4(P1_REG3_REG_7__SCAN_IN), .ZN(n9408) );
  NOR3_X1 U10664 ( .A1(n9409), .A2(P1_DATAO_REG_1__SCAN_IN), .A3(n9408), .ZN(
        n9410) );
  NAND4_X1 U10665 ( .A1(n9411), .A2(P1_IR_REG_12__SCAN_IN), .A3(
        P2_DATAO_REG_2__SCAN_IN), .A4(n9410), .ZN(n9413) );
  NAND4_X1 U10666 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .A3(P1_REG3_REG_14__SCAN_IN), .A4(n6639), .ZN(n9412) );
  NOR2_X1 U10667 ( .A1(n9413), .A2(n9412), .ZN(n9416) );
  NAND4_X1 U10668 ( .A1(n9417), .A2(n9416), .A3(n9415), .A4(n9414), .ZN(n9418)
         );
  NOR4_X1 U10669 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(P1_REG1_REG_15__SCAN_IN), 
        .A3(n9419), .A4(n9418), .ZN(n9436) );
  NOR4_X1 U10670 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(SI_30_), .A3(n10086), .A4(
        n9420), .ZN(n9435) );
  NOR4_X1 U10671 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9423), .A3(n9422), .A4(
        n9421), .ZN(n9424) );
  NAND3_X1 U10672 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_REG0_REG_29__SCAN_IN), 
        .A3(n9424), .ZN(n9433) );
  NOR4_X1 U10673 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .A3(P2_REG1_REG_31__SCAN_IN), .A4(n9425), .ZN(n9431) );
  NOR4_X1 U10674 ( .A1(P1_REG1_REG_27__SCAN_IN), .A2(P2_WR_REG_SCAN_IN), .A3(
        n8484), .A4(n9426), .ZN(n9430) );
  NOR4_X1 U10675 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(P2_REG0_REG_31__SCAN_IN), 
        .A3(n9427), .A4(n5213), .ZN(n9429) );
  NOR4_X1 U10676 ( .A1(P1_REG2_REG_28__SCAN_IN), .A2(P2_REG3_REG_27__SCAN_IN), 
        .A3(P2_REG2_REG_8__SCAN_IN), .A4(P2_REG0_REG_5__SCAN_IN), .ZN(n9428)
         );
  NAND4_X1 U10677 ( .A1(n9431), .A2(n9430), .A3(n9429), .A4(n9428), .ZN(n9432)
         );
  NOR4_X1 U10678 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(P2_D_REG_0__SCAN_IN), 
        .A3(n9433), .A4(n9432), .ZN(n9434) );
  NAND4_X1 U10679 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9436), .A3(n9435), .A4(
        n9434), .ZN(n9471) );
  NOR4_X1 U10680 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), 
        .A3(P2_ADDR_REG_8__SCAN_IN), .A4(n9437), .ZN(n9450) );
  NOR4_X1 U10681 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(P1_DATAO_REG_21__SCAN_IN), .A3(SI_21_), .A4(P1_DATAO_REG_19__SCAN_IN), .ZN(n9438) );
  NAND3_X1 U10682 ( .A1(P1_RD_REG_SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), .A3(
        n9438), .ZN(n9447) );
  NOR4_X1 U10683 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P2_ADDR_REG_14__SCAN_IN), 
        .A3(n6219), .A4(n9439), .ZN(n9445) );
  NOR4_X1 U10684 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .A3(P2_ADDR_REG_17__SCAN_IN), .A4(n9718), .ZN(n9444) );
  NOR4_X1 U10685 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(P2_DATAO_REG_8__SCAN_IN), 
        .A3(P2_DATAO_REG_7__SCAN_IN), .A4(SI_4_), .ZN(n9443) );
  NOR4_X1 U10686 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(P1_DATAO_REG_16__SCAN_IN), .A3(n9441), .A4(n9440), .ZN(n9442) );
  NAND4_X1 U10687 ( .A1(n9445), .A2(n9444), .A3(n9443), .A4(n9442), .ZN(n9446)
         );
  NOR4_X1 U10688 ( .A1(SI_24_), .A2(n9448), .A3(n9447), .A4(n9446), .ZN(n9449)
         );
  NAND4_X1 U10689 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .A3(n9450), .A4(n9449), .ZN(n9470) );
  NAND4_X1 U10690 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9458) );
  NAND4_X1 U10691 ( .A1(P1_STATE_REG_SCAN_IN), .A2(P1_REG1_REG_11__SCAN_IN), 
        .A3(P1_REG3_REG_0__SCAN_IN), .A4(P1_REG0_REG_0__SCAN_IN), .ZN(n9457)
         );
  NAND4_X1 U10692 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9452), .A4(n9451), .ZN(n9456) );
  NAND4_X1 U10693 ( .A1(P2_REG0_REG_3__SCAN_IN), .A2(P2_REG0_REG_0__SCAN_IN), 
        .A3(n9454), .A4(n9453), .ZN(n9455) );
  OR4_X1 U10694 ( .A1(n9458), .A2(n9457), .A3(n9456), .A4(n9455), .ZN(n9469)
         );
  NOR4_X1 U10695 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        n9460), .A4(n9459), .ZN(n9467) );
  NOR4_X1 U10696 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .A3(P2_REG0_REG_10__SCAN_IN), .A4(n9461), .ZN(n9463) );
  NOR4_X1 U10697 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P1_DATAO_REG_30__SCAN_IN), 
        .A3(P1_REG2_REG_31__SCAN_IN), .A4(n5999), .ZN(n9462) );
  AND4_X1 U10698 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(n9463), .A3(n9462), .A4(
        P2_IR_REG_5__SCAN_IN), .ZN(n9466) );
  NAND4_X1 U10699 ( .A1(n9467), .A2(n9466), .A3(n9465), .A4(n9464), .ZN(n9468)
         );
  NOR4_X1 U10700 ( .A1(n9471), .A2(n9470), .A3(n9469), .A4(n9468), .ZN(n9472)
         );
  XNOR2_X1 U10701 ( .A(n9473), .B(n9472), .ZN(n9474) );
  XNOR2_X1 U10702 ( .A(n9475), .B(n9474), .ZN(P1_U3267) );
  XNOR2_X1 U10703 ( .A(n9476), .B(n9478), .ZN(n9633) );
  XOR2_X1 U10704 ( .A(n9478), .B(n9477), .Z(n9480) );
  OAI222_X1 U10705 ( .A1(n9546), .A2(n9481), .B1(n9480), .B2(n9588), .C1(n9544), .C2(n9479), .ZN(n9629) );
  INV_X1 U10706 ( .A(n9494), .ZN(n9483) );
  AOI211_X1 U10707 ( .C1(n9631), .C2(n9483), .A(n10029), .B(n9482), .ZN(n9630)
         );
  NAND2_X1 U10708 ( .A1(n9630), .A2(n9573), .ZN(n9487) );
  INV_X1 U10709 ( .A(n9484), .ZN(n9485) );
  AOI22_X1 U10710 ( .A1(n9485), .A2(n9923), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n4382), .ZN(n9486) );
  OAI211_X1 U10711 ( .C1(n9488), .C2(n9930), .A(n9487), .B(n9486), .ZN(n9489)
         );
  AOI21_X1 U10712 ( .B1(n9629), .B2(n9926), .A(n9489), .ZN(n9490) );
  OAI21_X1 U10713 ( .B1(n9633), .B2(n9597), .A(n9490), .ZN(P1_U3268) );
  OAI21_X1 U10714 ( .B1(n9492), .B2(n9500), .A(n9491), .ZN(n9493) );
  INV_X1 U10715 ( .A(n9493), .ZN(n9638) );
  AOI21_X1 U10716 ( .B1(n9634), .B2(n9508), .A(n9494), .ZN(n9635) );
  AOI22_X1 U10717 ( .A1(n9495), .A2(n9923), .B1(n4382), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9496) );
  OAI21_X1 U10718 ( .B1(n9497), .B2(n9930), .A(n9496), .ZN(n9504) );
  NAND2_X1 U10719 ( .A1(n9515), .A2(n9498), .ZN(n9499) );
  XOR2_X1 U10720 ( .A(n9500), .B(n9499), .Z(n9501) );
  AOI222_X1 U10721 ( .A1(n9532), .A2(n9913), .B1(n9502), .B2(n9911), .C1(n9916), .C2(n9501), .ZN(n9637) );
  NOR2_X1 U10722 ( .A1(n9637), .A2(n4382), .ZN(n9503) );
  AOI211_X1 U10723 ( .C1(n9635), .C2(n9909), .A(n9504), .B(n9503), .ZN(n9505)
         );
  OAI21_X1 U10724 ( .B1(n9638), .B2(n9597), .A(n9505), .ZN(P1_U3269) );
  OAI21_X1 U10725 ( .B1(n9507), .B2(n9506), .A(n4438), .ZN(n9643) );
  INV_X1 U10726 ( .A(n9525), .ZN(n9510) );
  INV_X1 U10727 ( .A(n9508), .ZN(n9509) );
  AOI211_X1 U10728 ( .C1(n9640), .C2(n9510), .A(n10029), .B(n9509), .ZN(n9639)
         );
  INV_X1 U10729 ( .A(n9511), .ZN(n9512) );
  AOI22_X1 U10730 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(n4382), .B1(n9512), .B2(
        n9923), .ZN(n9513) );
  OAI21_X1 U10731 ( .B1(n9514), .B2(n9930), .A(n9513), .ZN(n9522) );
  OAI21_X1 U10732 ( .B1(n9517), .B2(n9516), .A(n9515), .ZN(n9520) );
  AOI222_X1 U10733 ( .A1(n9916), .A2(n9520), .B1(n9519), .B2(n9911), .C1(n9518), .C2(n9913), .ZN(n9642) );
  NOR2_X1 U10734 ( .A1(n9642), .A2(n4382), .ZN(n9521) );
  AOI211_X1 U10735 ( .C1(n9639), .C2(n9573), .A(n9522), .B(n9521), .ZN(n9523)
         );
  OAI21_X1 U10736 ( .B1(n9597), .B2(n9643), .A(n9523), .ZN(P1_U3270) );
  XNOR2_X1 U10737 ( .A(n9524), .B(n9531), .ZN(n9648) );
  INV_X1 U10738 ( .A(n9547), .ZN(n9526) );
  AOI21_X1 U10739 ( .B1(n9644), .B2(n9526), .A(n9525), .ZN(n9645) );
  INV_X1 U10740 ( .A(n9527), .ZN(n9528) );
  AOI22_X1 U10741 ( .A1(n4382), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9528), .B2(
        n9923), .ZN(n9529) );
  OAI21_X1 U10742 ( .B1(n9530), .B2(n9930), .A(n9529), .ZN(n9535) );
  XOR2_X1 U10743 ( .A(n9531), .B(n4424), .Z(n9533) );
  AOI222_X1 U10744 ( .A1(n9916), .A2(n9533), .B1(n9532), .B2(n9911), .C1(n9569), .C2(n9913), .ZN(n9647) );
  NOR2_X1 U10745 ( .A1(n9647), .A2(n4382), .ZN(n9534) );
  AOI211_X1 U10746 ( .C1(n9645), .C2(n9909), .A(n9535), .B(n9534), .ZN(n9536)
         );
  OAI21_X1 U10747 ( .B1(n9648), .B2(n9597), .A(n9536), .ZN(P1_U3271) );
  XNOR2_X1 U10748 ( .A(n9537), .B(n9540), .ZN(n9653) );
  INV_X1 U10749 ( .A(n9538), .ZN(n9541) );
  AOI21_X1 U10750 ( .B1(n9541), .B2(n9540), .A(n9539), .ZN(n9542) );
  OAI222_X1 U10751 ( .A1(n9546), .A2(n9545), .B1(n9544), .B2(n9543), .C1(n9588), .C2(n9542), .ZN(n9649) );
  INV_X1 U10752 ( .A(n9559), .ZN(n9548) );
  AOI211_X1 U10753 ( .C1(n9651), .C2(n9548), .A(n10029), .B(n9547), .ZN(n9650)
         );
  NAND2_X1 U10754 ( .A1(n9650), .A2(n9573), .ZN(n9552) );
  INV_X1 U10755 ( .A(n9549), .ZN(n9550) );
  AOI22_X1 U10756 ( .A1(n4382), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9923), .B2(
        n9550), .ZN(n9551) );
  OAI211_X1 U10757 ( .C1(n9553), .C2(n9930), .A(n9552), .B(n9551), .ZN(n9554)
         );
  AOI21_X1 U10758 ( .B1(n9649), .B2(n9926), .A(n9554), .ZN(n9555) );
  OAI21_X1 U10759 ( .B1(n9653), .B2(n9597), .A(n9555), .ZN(P1_U3272) );
  OAI21_X1 U10760 ( .B1(n9558), .B2(n9557), .A(n9556), .ZN(n9658) );
  AOI211_X1 U10761 ( .C1(n9655), .C2(n9576), .A(n10029), .B(n9559), .ZN(n9654)
         );
  INV_X1 U10762 ( .A(n9560), .ZN(n9561) );
  AOI22_X1 U10763 ( .A1(n4382), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9561), .B2(
        n9923), .ZN(n9562) );
  OAI21_X1 U10764 ( .B1(n9563), .B2(n9930), .A(n9562), .ZN(n9572) );
  AND2_X1 U10765 ( .A1(n9584), .A2(n9564), .ZN(n9567) );
  OAI21_X1 U10766 ( .B1(n9567), .B2(n9566), .A(n9565), .ZN(n9570) );
  AOI222_X1 U10767 ( .A1(n9916), .A2(n9570), .B1(n9569), .B2(n9911), .C1(n9568), .C2(n9913), .ZN(n9657) );
  NOR2_X1 U10768 ( .A1(n9657), .A2(n4382), .ZN(n9571) );
  AOI211_X1 U10769 ( .C1(n9654), .C2(n9573), .A(n9572), .B(n9571), .ZN(n9574)
         );
  OAI21_X1 U10770 ( .B1(n9597), .B2(n9658), .A(n9574), .ZN(P1_U3273) );
  XNOR2_X1 U10771 ( .A(n9575), .B(n9585), .ZN(n9663) );
  INV_X1 U10772 ( .A(n9576), .ZN(n9577) );
  AOI21_X1 U10773 ( .B1(n9659), .B2(n9578), .A(n9577), .ZN(n9660) );
  INV_X1 U10774 ( .A(n9579), .ZN(n9580) );
  AOI22_X1 U10775 ( .A1(n4382), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9580), .B2(
        n9923), .ZN(n9581) );
  OAI21_X1 U10776 ( .B1(n9582), .B2(n9930), .A(n9581), .ZN(n9595) );
  AND2_X1 U10777 ( .A1(n9583), .A2(n9911), .ZN(n9592) );
  INV_X1 U10778 ( .A(n9584), .ZN(n9590) );
  AOI21_X1 U10779 ( .B1(n9587), .B2(n9586), .A(n9585), .ZN(n9589) );
  NOR3_X1 U10780 ( .A1(n9590), .A2(n9589), .A3(n9588), .ZN(n9591) );
  AOI211_X1 U10781 ( .C1(n9913), .C2(n9593), .A(n9592), .B(n9591), .ZN(n9662)
         );
  NOR2_X1 U10782 ( .A1(n9662), .A2(n4382), .ZN(n9594) );
  AOI211_X1 U10783 ( .C1(n9660), .C2(n9909), .A(n9595), .B(n9594), .ZN(n9596)
         );
  OAI21_X1 U10784 ( .B1(n9597), .B2(n9663), .A(n9596), .ZN(P1_U3274) );
  NAND2_X1 U10785 ( .A1(n9920), .A2(n10009), .ZN(n10034) );
  OAI211_X1 U10786 ( .C1(n9602), .C2(n9995), .A(n9601), .B(n9600), .ZN(n9675)
         );
  MUX2_X1 U10787 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9675), .S(n10049), .Z(
        P1_U3552) );
  AOI22_X1 U10788 ( .A1(n9604), .A2(n10005), .B1(n10004), .B2(n9603), .ZN(
        n9605) );
  AOI21_X1 U10789 ( .B1(n10004), .B2(n9609), .A(n9608), .ZN(n9610) );
  OAI211_X1 U10790 ( .C1(n9612), .C2(n9995), .A(n9611), .B(n9610), .ZN(n9677)
         );
  MUX2_X1 U10791 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9677), .S(n10049), .Z(
        P1_U3550) );
  AOI21_X1 U10792 ( .B1(n10004), .B2(n9614), .A(n9613), .ZN(n9615) );
  OAI211_X1 U10793 ( .C1(n9617), .C2(n9995), .A(n9616), .B(n9615), .ZN(n9678)
         );
  MUX2_X1 U10794 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9678), .S(n10049), .Z(
        P1_U3549) );
  AOI21_X1 U10795 ( .B1(n10004), .B2(n9619), .A(n9618), .ZN(n9620) );
  OAI211_X1 U10796 ( .C1(n9622), .C2(n9995), .A(n9621), .B(n9620), .ZN(n9679)
         );
  MUX2_X1 U10797 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9679), .S(n10049), .Z(
        P1_U3548) );
  OAI211_X1 U10798 ( .C1(n9625), .C2(n10027), .A(n9624), .B(n9623), .ZN(n9626)
         );
  AOI21_X1 U10799 ( .B1(n9627), .B2(n10034), .A(n9626), .ZN(n9628) );
  INV_X1 U10800 ( .A(n9628), .ZN(n9680) );
  MUX2_X1 U10801 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9680), .S(n10049), .Z(
        P1_U3547) );
  AOI211_X1 U10802 ( .C1(n10004), .C2(n9631), .A(n9630), .B(n9629), .ZN(n9632)
         );
  OAI21_X1 U10803 ( .B1(n9633), .B2(n9995), .A(n9632), .ZN(n9681) );
  MUX2_X1 U10804 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9681), .S(n10049), .Z(
        P1_U3546) );
  AOI22_X1 U10805 ( .A1(n9635), .A2(n10005), .B1(n10004), .B2(n9634), .ZN(
        n9636) );
  OAI211_X1 U10806 ( .C1(n9638), .C2(n9995), .A(n9637), .B(n9636), .ZN(n9682)
         );
  MUX2_X1 U10807 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9682), .S(n10049), .Z(
        P1_U3545) );
  AOI21_X1 U10808 ( .B1(n10004), .B2(n9640), .A(n9639), .ZN(n9641) );
  OAI211_X1 U10809 ( .C1(n9643), .C2(n9995), .A(n9642), .B(n9641), .ZN(n9683)
         );
  MUX2_X1 U10810 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9683), .S(n10049), .Z(
        P1_U3544) );
  AOI22_X1 U10811 ( .A1(n9645), .A2(n10005), .B1(n10004), .B2(n9644), .ZN(
        n9646) );
  OAI211_X1 U10812 ( .C1(n9648), .C2(n9995), .A(n9647), .B(n9646), .ZN(n9684)
         );
  MUX2_X1 U10813 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9684), .S(n10049), .Z(
        P1_U3543) );
  AOI211_X1 U10814 ( .C1(n10004), .C2(n9651), .A(n9650), .B(n9649), .ZN(n9652)
         );
  OAI21_X1 U10815 ( .B1(n9995), .B2(n9653), .A(n9652), .ZN(n9685) );
  MUX2_X1 U10816 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9685), .S(n10049), .Z(
        P1_U3542) );
  AOI21_X1 U10817 ( .B1(n10004), .B2(n9655), .A(n9654), .ZN(n9656) );
  OAI211_X1 U10818 ( .C1(n9658), .C2(n9995), .A(n9657), .B(n9656), .ZN(n9686)
         );
  MUX2_X1 U10819 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9686), .S(n10049), .Z(
        P1_U3541) );
  AOI22_X1 U10820 ( .A1(n9660), .A2(n10005), .B1(n10004), .B2(n9659), .ZN(
        n9661) );
  OAI211_X1 U10821 ( .C1(n9663), .C2(n9995), .A(n9662), .B(n9661), .ZN(n9687)
         );
  MUX2_X1 U10822 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9687), .S(n10049), .Z(
        P1_U3540) );
  AOI211_X1 U10823 ( .C1(n10004), .C2(n9666), .A(n9665), .B(n9664), .ZN(n9667)
         );
  OAI21_X1 U10824 ( .B1(n9995), .B2(n9668), .A(n9667), .ZN(n9688) );
  MUX2_X1 U10825 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9688), .S(n10049), .Z(
        P1_U3539) );
  AOI22_X1 U10826 ( .A1(n9670), .A2(n10005), .B1(n10004), .B2(n9669), .ZN(
        n9671) );
  OAI211_X1 U10827 ( .C1(n9673), .C2(n9995), .A(n9672), .B(n9671), .ZN(n9689)
         );
  MUX2_X1 U10828 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9689), .S(n10049), .Z(
        P1_U3538) );
  MUX2_X1 U10829 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9674), .S(n10049), .Z(
        P1_U3523) );
  MUX2_X1 U10830 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9675), .S(n10037), .Z(
        P1_U3520) );
  MUX2_X1 U10831 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9676), .S(n10037), .Z(
        P1_U3519) );
  MUX2_X1 U10832 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9677), .S(n10037), .Z(
        P1_U3518) );
  MUX2_X1 U10833 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9678), .S(n10037), .Z(
        P1_U3517) );
  MUX2_X1 U10834 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9679), .S(n10037), .Z(
        P1_U3516) );
  MUX2_X1 U10835 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9680), .S(n10037), .Z(
        P1_U3515) );
  MUX2_X1 U10836 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9681), .S(n10037), .Z(
        P1_U3514) );
  MUX2_X1 U10837 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9682), .S(n10037), .Z(
        P1_U3513) );
  MUX2_X1 U10838 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9683), .S(n10037), .Z(
        P1_U3512) );
  MUX2_X1 U10839 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9684), .S(n10037), .Z(
        P1_U3511) );
  MUX2_X1 U10840 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9685), .S(n10037), .Z(
        P1_U3510) );
  MUX2_X1 U10841 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9686), .S(n10037), .Z(
        P1_U3508) );
  MUX2_X1 U10842 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9687), .S(n10037), .Z(
        P1_U3505) );
  MUX2_X1 U10843 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9688), .S(n10037), .Z(
        P1_U3502) );
  MUX2_X1 U10844 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9689), .S(n10037), .Z(
        P1_U3499) );
  MUX2_X1 U10845 ( .A(P1_D_REG_1__SCAN_IN), .B(n9690), .S(n9691), .Z(P1_U3441)
         );
  AND2_X2 U10846 ( .A1(n9692), .A2(n9691), .ZN(n9967) );
  MUX2_X1 U10847 ( .A(P1_D_REG_0__SCAN_IN), .B(n9693), .S(n9967), .Z(P1_U3440)
         );
  OAI222_X1 U10848 ( .A1(n9698), .A2(n9697), .B1(n9696), .B2(P1_U3084), .C1(
        n9695), .C2(n9694), .ZN(P1_U3324) );
  NAND2_X1 U10849 ( .A1(n9699), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9701) );
  OAI211_X1 U10850 ( .C1(n9702), .C2(n9695), .A(n9701), .B(n9700), .ZN(
        P1_U3325) );
  INV_X1 U10851 ( .A(n9703), .ZN(n9704) );
  MUX2_X1 U10852 ( .A(n9704), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  MUX2_X1 U10853 ( .A(n5025), .B(P2_ADDR_REG_19__SCAN_IN), .S(
        P1_ADDR_REG_19__SCAN_IN), .Z(n9729) );
  NOR2_X1 U10854 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9705) );
  AOI21_X1 U10855 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9705), .ZN(n10187) );
  NOR2_X1 U10856 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9706) );
  AOI21_X1 U10857 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9706), .ZN(n10190) );
  NOR2_X1 U10858 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9707) );
  AOI21_X1 U10859 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9707), .ZN(n10193) );
  NOR2_X1 U10860 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9708) );
  AOI21_X1 U10861 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9708), .ZN(n10196) );
  NOR2_X1 U10862 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9709) );
  AOI21_X1 U10863 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9709), .ZN(n10199) );
  NOR2_X1 U10864 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n9710) );
  AOI21_X1 U10865 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n9710), .ZN(n10238) );
  INV_X1 U10866 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10183) );
  INV_X1 U10867 ( .A(n10182), .ZN(n10180) );
  INV_X1 U10868 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10179) );
  NAND2_X1 U10869 ( .A1(n10180), .A2(n10179), .ZN(n10178) );
  AOI22_X1 U10870 ( .A1(n10182), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(n10178), .ZN(n10232) );
  NAND2_X1 U10871 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9711) );
  OAI21_X1 U10872 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n9711), .ZN(n10231) );
  NOR2_X1 U10873 ( .A1(n10232), .A2(n10231), .ZN(n10230) );
  AOI21_X1 U10874 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10230), .ZN(n10235) );
  NAND2_X1 U10875 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9712) );
  OAI21_X1 U10876 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n9712), .ZN(n10234) );
  NOR2_X1 U10877 ( .A1(n10235), .A2(n10234), .ZN(n10233) );
  AOI21_X1 U10878 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10233), .ZN(n10237) );
  NAND2_X1 U10879 ( .A1(n10238), .A2(n10237), .ZN(n10236) );
  OAI21_X1 U10880 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10236), .ZN(n9713) );
  NAND2_X1 U10881 ( .A1(n9714), .A2(n9713), .ZN(n10214) );
  INV_X1 U10882 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10216) );
  OR2_X1 U10883 ( .A1(n9714), .A2(n9713), .ZN(n10215) );
  NAND2_X1 U10884 ( .A1(n10216), .A2(n10215), .ZN(n10212) );
  NAND2_X1 U10885 ( .A1(n10214), .A2(n10212), .ZN(n9716) );
  NOR2_X1 U10886 ( .A1(n9716), .A2(n9715), .ZN(n9717) );
  XNOR2_X1 U10887 ( .A(n9716), .B(n9715), .ZN(n10210) );
  AOI22_X1 U10888 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9718), .B1(
        P2_ADDR_REG_7__SCAN_IN), .B2(n9881), .ZN(n10218) );
  AOI21_X1 U10889 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10217), .ZN(n9719) );
  NOR2_X1 U10890 ( .A1(n9719), .A2(n6136), .ZN(n9720) );
  XNOR2_X1 U10891 ( .A(n6136), .B(n9719), .ZN(n10228) );
  NOR2_X1 U10892 ( .A1(n9721), .A2(n9722), .ZN(n9723) );
  INV_X1 U10893 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10226) );
  XNOR2_X1 U10894 ( .A(n9722), .B(n9721), .ZN(n10225) );
  NAND2_X1 U10895 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9724) );
  OAI21_X1 U10896 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9724), .ZN(n10207) );
  NAND2_X1 U10897 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9725) );
  OAI21_X1 U10898 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9725), .ZN(n10204) );
  AOI21_X1 U10899 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10203), .ZN(n10202) );
  NOR2_X1 U10900 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9726) );
  AOI21_X1 U10901 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9726), .ZN(n10201) );
  NAND2_X1 U10902 ( .A1(n10202), .A2(n10201), .ZN(n10200) );
  OAI21_X1 U10903 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10200), .ZN(n10198) );
  NAND2_X1 U10904 ( .A1(n10199), .A2(n10198), .ZN(n10197) );
  OAI21_X1 U10905 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10197), .ZN(n10195) );
  NAND2_X1 U10906 ( .A1(n10196), .A2(n10195), .ZN(n10194) );
  OAI21_X1 U10907 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10194), .ZN(n10192) );
  NAND2_X1 U10908 ( .A1(n10193), .A2(n10192), .ZN(n10191) );
  OAI21_X1 U10909 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10191), .ZN(n10189) );
  NAND2_X1 U10910 ( .A1(n10190), .A2(n10189), .ZN(n10188) );
  OAI21_X1 U10911 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10188), .ZN(n10186) );
  NAND2_X1 U10912 ( .A1(n10187), .A2(n10186), .ZN(n10185) );
  OAI21_X1 U10913 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10185), .ZN(n10221) );
  NOR2_X1 U10914 ( .A1(n10222), .A2(n10221), .ZN(n9727) );
  NAND2_X1 U10915 ( .A1(n10222), .A2(n10221), .ZN(n10220) );
  OAI21_X1 U10916 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9727), .A(n10220), .ZN(
        n9728) );
  XOR2_X1 U10917 ( .A(n9729), .B(n9728), .Z(ADD_1071_U4) );
  AOI22_X1 U10918 ( .A1(n10056), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9740) );
  NAND2_X1 U10919 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9732) );
  AOI211_X1 U10920 ( .C1(n9732), .C2(n9731), .A(n9730), .B(n10051), .ZN(n9737)
         );
  NAND2_X1 U10921 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9735) );
  AOI211_X1 U10922 ( .C1(n9735), .C2(n9734), .A(n9733), .B(n9744), .ZN(n9736)
         );
  AOI211_X1 U10923 ( .C1(n10053), .C2(n9738), .A(n9737), .B(n9736), .ZN(n9739)
         );
  NAND2_X1 U10924 ( .A1(n9740), .A2(n9739), .ZN(P2_U3246) );
  AOI22_X1 U10925 ( .A1(n10056), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n4374), .ZN(n9752) );
  AOI211_X1 U10926 ( .C1(n9743), .C2(n9742), .A(n9741), .B(n10051), .ZN(n9749)
         );
  AOI211_X1 U10927 ( .C1(n9747), .C2(n9746), .A(n9745), .B(n9744), .ZN(n9748)
         );
  AOI211_X1 U10928 ( .C1(n10053), .C2(n9750), .A(n9749), .B(n9748), .ZN(n9751)
         );
  NAND2_X1 U10929 ( .A1(n9752), .A2(n9751), .ZN(P2_U3247) );
  OAI21_X1 U10930 ( .B1(n7836), .B2(n10027), .A(n9762), .ZN(n9753) );
  AOI21_X1 U10931 ( .B1(n9754), .B2(n10005), .A(n9753), .ZN(n9755) );
  AOI22_X1 U10932 ( .A1(n10049), .A2(n9755), .B1(n6109), .B2(n10047), .ZN(
        P1_U3554) );
  AOI22_X1 U10933 ( .A1(n10037), .A2(n9755), .B1(n6111), .B2(n10035), .ZN(
        P1_U3522) );
  INV_X1 U10934 ( .A(n9756), .ZN(n9758) );
  AOI22_X1 U10935 ( .A1(n10177), .A2(n9761), .B1(n5643), .B2(n10175), .ZN(
        P2_U3550) );
  INV_X1 U10936 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9760) );
  AOI22_X1 U10937 ( .A1(n10163), .A2(n9761), .B1(n9760), .B2(n10161), .ZN(
        P2_U3518) );
  OAI21_X1 U10938 ( .B1(n9763), .B2(n10027), .A(n9762), .ZN(n9764) );
  AOI21_X1 U10939 ( .B1(n10005), .B2(n9765), .A(n9764), .ZN(n9790) );
  AOI22_X1 U10940 ( .A1(n10049), .A2(n9790), .B1(n7716), .B2(n10047), .ZN(
        P1_U3553) );
  OAI211_X1 U10941 ( .C1(n9768), .C2(n10027), .A(n9767), .B(n9766), .ZN(n9769)
         );
  AOI21_X1 U10942 ( .B1(n10034), .B2(n9770), .A(n9769), .ZN(n9792) );
  AOI22_X1 U10943 ( .A1(n10049), .A2(n9792), .B1(n9771), .B2(n10047), .ZN(
        P1_U3537) );
  INV_X1 U10944 ( .A(n10009), .ZN(n10025) );
  INV_X1 U10945 ( .A(n9772), .ZN(n9776) );
  OAI22_X1 U10946 ( .A1(n9773), .A2(n10029), .B1(n4486), .B2(n10027), .ZN(
        n9775) );
  AOI211_X1 U10947 ( .C1(n10025), .C2(n9776), .A(n9775), .B(n9774), .ZN(n9794)
         );
  AOI22_X1 U10948 ( .A1(n10049), .A2(n9794), .B1(n9777), .B2(n10047), .ZN(
        P1_U3536) );
  INV_X1 U10949 ( .A(n9778), .ZN(n9783) );
  OAI21_X1 U10950 ( .B1(n9780), .B2(n10027), .A(n9779), .ZN(n9782) );
  AOI211_X1 U10951 ( .C1(n10025), .C2(n9783), .A(n9782), .B(n9781), .ZN(n9795)
         );
  AOI22_X1 U10952 ( .A1(n10049), .A2(n9795), .B1(n9784), .B2(n10047), .ZN(
        P1_U3535) );
  OAI22_X1 U10953 ( .A1(n9786), .A2(n10029), .B1(n9785), .B2(n10027), .ZN(
        n9788) );
  AOI211_X1 U10954 ( .C1(n9789), .C2(n10034), .A(n9788), .B(n9787), .ZN(n9797)
         );
  AOI22_X1 U10955 ( .A1(n10049), .A2(n9797), .B1(n6995), .B2(n10047), .ZN(
        P1_U3534) );
  AOI22_X1 U10956 ( .A1(n10037), .A2(n9790), .B1(n7718), .B2(n10035), .ZN(
        P1_U3521) );
  INV_X1 U10957 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9791) );
  AOI22_X1 U10958 ( .A1(n10037), .A2(n9792), .B1(n9791), .B2(n10035), .ZN(
        P1_U3496) );
  INV_X1 U10959 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9793) );
  AOI22_X1 U10960 ( .A1(n10037), .A2(n9794), .B1(n9793), .B2(n10035), .ZN(
        P1_U3493) );
  AOI22_X1 U10961 ( .A1(n10037), .A2(n9795), .B1(n7039), .B2(n10035), .ZN(
        P1_U3490) );
  INV_X1 U10962 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9796) );
  AOI22_X1 U10963 ( .A1(n10037), .A2(n9797), .B1(n9796), .B2(n10035), .ZN(
        P1_U3487) );
  XNOR2_X1 U10964 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  AOI22_X1 U10965 ( .A1(P2_RD_REG_SCAN_IN), .A2(n9799), .B1(P1_RD_REG_SCAN_IN), 
        .B2(n9798), .ZN(U126) );
  AOI21_X1 U10966 ( .B1(n9802), .B2(n9815), .A(n9800), .ZN(n9835) );
  NAND2_X1 U10967 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(n9806), .ZN(n9805) );
  AOI21_X1 U10968 ( .B1(n9802), .B2(n9801), .A(n9800), .ZN(n9803) );
  NOR2_X1 U10969 ( .A1(n9803), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n9834) );
  AOI211_X1 U10970 ( .C1(n9835), .C2(n9805), .A(n9804), .B(n9834), .ZN(n9808)
         );
  NOR3_X1 U10971 ( .A1(n9896), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n9806), .ZN(
        n9807) );
  AOI221_X1 U10972 ( .B1(n9808), .B2(P1_STATE_REG_SCAN_IN), .C1(
        P1_REG3_REG_0__SCAN_IN), .C2(P1_U3084), .A(n9807), .ZN(n9809) );
  OAI21_X1 U10973 ( .B1(n10184), .B2(n9880), .A(n9809), .ZN(P1_U3241) );
  NAND2_X1 U10974 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9812) );
  AOI211_X1 U10975 ( .C1(n9812), .C2(n9811), .A(n9810), .B(n9896), .ZN(n9817)
         );
  AOI211_X1 U10976 ( .C1(n9815), .C2(n9814), .A(n9813), .B(n9827), .ZN(n9816)
         );
  AOI211_X1 U10977 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(P1_U3084), .A(n9817), 
        .B(n9816), .ZN(n9822) );
  OAI22_X1 U10978 ( .A1(n9880), .A2(n10179), .B1(n9819), .B2(n9818), .ZN(n9820) );
  INV_X1 U10979 ( .A(n9820), .ZN(n9821) );
  NAND2_X1 U10980 ( .A1(n9822), .A2(n9821), .ZN(P1_U3242) );
  INV_X1 U10981 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9841) );
  AOI211_X1 U10982 ( .C1(n9825), .C2(n9824), .A(n9823), .B(n9896), .ZN(n9826)
         );
  AOI21_X1 U10983 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(P1_U3084), .A(n9826), 
        .ZN(n9840) );
  AOI211_X1 U10984 ( .C1(n9830), .C2(n9829), .A(n9828), .B(n9827), .ZN(n9837)
         );
  NAND2_X1 U10985 ( .A1(n9832), .A2(n9831), .ZN(n9836) );
  AOI211_X1 U10986 ( .C1(n9836), .C2(n9835), .A(n9834), .B(n9833), .ZN(n9848)
         );
  AOI211_X1 U10987 ( .C1(n9898), .C2(n9838), .A(n9837), .B(n9848), .ZN(n9839)
         );
  OAI211_X1 U10988 ( .C1(n9880), .C2(n9841), .A(n9840), .B(n9839), .ZN(
        P1_U3243) );
  INV_X1 U10989 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9853) );
  XNOR2_X1 U10990 ( .A(n9843), .B(n9842), .ZN(n9845) );
  AOI22_X1 U10991 ( .A1(n9891), .A2(n9845), .B1(n9844), .B2(n9898), .ZN(n9852)
         );
  XNOR2_X1 U10992 ( .A(n9847), .B(n9846), .ZN(n9850) );
  AOI211_X1 U10993 ( .C1(n9872), .C2(n9850), .A(n9849), .B(n9848), .ZN(n9851)
         );
  OAI211_X1 U10994 ( .C1(n9880), .C2(n9853), .A(n9852), .B(n9851), .ZN(
        P1_U3245) );
  NOR2_X1 U10995 ( .A1(n9855), .A2(n9854), .ZN(n9856) );
  NOR3_X1 U10996 ( .A1(n9896), .A2(n9857), .A3(n9856), .ZN(n9858) );
  AOI211_X1 U10997 ( .C1(n9898), .C2(n9860), .A(n9859), .B(n9858), .ZN(n9866)
         );
  OAI21_X1 U10998 ( .B1(n9863), .B2(n9862), .A(n9861), .ZN(n9864) );
  NAND2_X1 U10999 ( .A1(n9891), .A2(n9864), .ZN(n9865) );
  OAI211_X1 U11000 ( .C1(n10216), .C2(n9880), .A(n9866), .B(n9865), .ZN(
        P1_U3246) );
  OAI21_X1 U11001 ( .B1(n9869), .B2(n9868), .A(n9867), .ZN(n9871) );
  AOI21_X1 U11002 ( .B1(n9872), .B2(n9871), .A(n9870), .ZN(n9879) );
  OAI21_X1 U11003 ( .B1(n9875), .B2(n9874), .A(n9873), .ZN(n9877) );
  AOI22_X1 U11004 ( .A1(n9891), .A2(n9877), .B1(n9876), .B2(n9898), .ZN(n9878)
         );
  OAI211_X1 U11005 ( .C1(n9881), .C2(n9880), .A(n9879), .B(n9878), .ZN(
        P1_U3248) );
  OAI21_X1 U11006 ( .B1(n9884), .B2(n9883), .A(n9882), .ZN(n9885) );
  INV_X1 U11007 ( .A(n9885), .ZN(n9895) );
  INV_X1 U11008 ( .A(n9886), .ZN(n9890) );
  NAND2_X1 U11009 ( .A1(n9888), .A2(n9887), .ZN(n9889) );
  NAND3_X1 U11010 ( .A1(n9891), .A2(n9890), .A3(n9889), .ZN(n9894) );
  INV_X1 U11011 ( .A(n9892), .ZN(n9893) );
  OAI211_X1 U11012 ( .C1(n9896), .C2(n9895), .A(n9894), .B(n9893), .ZN(n9897)
         );
  INV_X1 U11013 ( .A(n9897), .ZN(n9902) );
  AOI22_X1 U11014 ( .A1(n9900), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n9899), .B2(
        n9898), .ZN(n9901) );
  NAND2_X1 U11015 ( .A1(n9902), .A2(n9901), .ZN(P1_U3250) );
  NAND2_X1 U11016 ( .A1(n6872), .A2(n9903), .ZN(n9904) );
  XOR2_X1 U11017 ( .A(n9915), .B(n9904), .Z(n9921) );
  INV_X1 U11018 ( .A(n9921), .ZN(n9986) );
  INV_X1 U11019 ( .A(n9905), .ZN(n9910) );
  OAI21_X1 U11020 ( .B1(n9907), .B2(n9982), .A(n9906), .ZN(n9983) );
  INV_X1 U11021 ( .A(n9983), .ZN(n9908) );
  AOI22_X1 U11022 ( .A1(n9986), .A2(n9910), .B1(n9909), .B2(n9908), .ZN(n9928)
         );
  AOI22_X1 U11023 ( .A1(n9913), .A2(n6727), .B1(n9912), .B2(n9911), .ZN(n9919)
         );
  XNOR2_X1 U11024 ( .A(n9915), .B(n9914), .ZN(n9917) );
  NAND2_X1 U11025 ( .A1(n9917), .A2(n9916), .ZN(n9918) );
  OAI211_X1 U11026 ( .C1(n9921), .C2(n9920), .A(n9919), .B(n9918), .ZN(n9984)
         );
  AOI22_X1 U11027 ( .A1(n4382), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9923), .B2(
        n9922), .ZN(n9924) );
  OAI21_X1 U11028 ( .B1(n9982), .B2(n9930), .A(n9924), .ZN(n9925) );
  AOI21_X1 U11029 ( .B1(n9984), .B2(n9926), .A(n9925), .ZN(n9927) );
  NAND2_X1 U11030 ( .A1(n9928), .A2(n9927), .ZN(P1_U3288) );
  AOI21_X1 U11031 ( .B1(n9931), .B2(n9930), .A(n9929), .ZN(n9934) );
  NOR2_X1 U11032 ( .A1(n9932), .A2(n4382), .ZN(n9933) );
  AOI211_X1 U11033 ( .C1(n4382), .C2(P1_REG2_REG_0__SCAN_IN), .A(n9934), .B(
        n9933), .ZN(n9935) );
  OAI21_X1 U11034 ( .B1(n9936), .B2(n6098), .A(n9935), .ZN(P1_U3291) );
  NOR2_X1 U11035 ( .A1(n9967), .A2(n9937), .ZN(P1_U3292) );
  NOR2_X1 U11036 ( .A1(n9967), .A2(n9938), .ZN(P1_U3293) );
  NOR2_X1 U11037 ( .A1(n9967), .A2(n9939), .ZN(P1_U3294) );
  NOR2_X1 U11038 ( .A1(n9967), .A2(n9940), .ZN(P1_U3295) );
  NOR2_X1 U11039 ( .A1(n9967), .A2(n9941), .ZN(P1_U3296) );
  NOR2_X1 U11040 ( .A1(n9967), .A2(n9942), .ZN(P1_U3297) );
  NOR2_X1 U11041 ( .A1(n9967), .A2(n9943), .ZN(P1_U3298) );
  INV_X1 U11042 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9944) );
  NOR2_X1 U11043 ( .A1(n9967), .A2(n9944), .ZN(P1_U3299) );
  NOR2_X1 U11044 ( .A1(n9967), .A2(n9945), .ZN(P1_U3300) );
  NOR2_X1 U11045 ( .A1(n9967), .A2(n9946), .ZN(P1_U3301) );
  INV_X1 U11046 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9947) );
  NOR2_X1 U11047 ( .A1(n9967), .A2(n9947), .ZN(P1_U3302) );
  NOR2_X1 U11048 ( .A1(n9967), .A2(n9948), .ZN(P1_U3303) );
  NOR2_X1 U11049 ( .A1(n9967), .A2(n9949), .ZN(P1_U3304) );
  NOR2_X1 U11050 ( .A1(n9967), .A2(n9950), .ZN(P1_U3305) );
  INV_X1 U11051 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9951) );
  NOR2_X1 U11052 ( .A1(n9967), .A2(n9951), .ZN(P1_U3306) );
  INV_X1 U11053 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9952) );
  NOR2_X1 U11054 ( .A1(n9967), .A2(n9952), .ZN(P1_U3307) );
  INV_X1 U11055 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n9953) );
  NOR2_X1 U11056 ( .A1(n9967), .A2(n9953), .ZN(P1_U3308) );
  INV_X1 U11057 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9954) );
  NOR2_X1 U11058 ( .A1(n9967), .A2(n9954), .ZN(P1_U3309) );
  INV_X1 U11059 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9955) );
  NOR2_X1 U11060 ( .A1(n9967), .A2(n9955), .ZN(P1_U3310) );
  INV_X1 U11061 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9956) );
  NOR2_X1 U11062 ( .A1(n9967), .A2(n9956), .ZN(P1_U3311) );
  INV_X1 U11063 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9957) );
  NOR2_X1 U11064 ( .A1(n9967), .A2(n9957), .ZN(P1_U3312) );
  NOR2_X1 U11065 ( .A1(n9967), .A2(n9958), .ZN(P1_U3313) );
  INV_X1 U11066 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9959) );
  NOR2_X1 U11067 ( .A1(n9967), .A2(n9959), .ZN(P1_U3314) );
  INV_X1 U11068 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9960) );
  NOR2_X1 U11069 ( .A1(n9967), .A2(n9960), .ZN(P1_U3315) );
  INV_X1 U11070 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9961) );
  NOR2_X1 U11071 ( .A1(n9967), .A2(n9961), .ZN(P1_U3316) );
  INV_X1 U11072 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9962) );
  NOR2_X1 U11073 ( .A1(n9967), .A2(n9962), .ZN(P1_U3317) );
  INV_X1 U11074 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9963) );
  NOR2_X1 U11075 ( .A1(n9967), .A2(n9963), .ZN(P1_U3318) );
  NOR2_X1 U11076 ( .A1(n9967), .A2(n9964), .ZN(P1_U3319) );
  NOR2_X1 U11077 ( .A1(n9967), .A2(n9965), .ZN(P1_U3320) );
  INV_X1 U11078 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n9966) );
  NOR2_X1 U11079 ( .A1(n9967), .A2(n9966), .ZN(P1_U3321) );
  INV_X1 U11080 ( .A(n9968), .ZN(n9973) );
  OAI21_X1 U11081 ( .B1(n9970), .B2(n10027), .A(n9969), .ZN(n9972) );
  AOI211_X1 U11082 ( .C1(n10025), .C2(n9973), .A(n9972), .B(n9971), .ZN(n10038) );
  INV_X1 U11083 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U11084 ( .A1(n10037), .A2(n10038), .B1(n9974), .B2(n10035), .ZN(
        P1_U3457) );
  AOI22_X1 U11085 ( .A1(n9976), .A2(n10005), .B1(n10004), .B2(n9975), .ZN(
        n9977) );
  OAI211_X1 U11086 ( .C1(n9979), .C2(n10009), .A(n9978), .B(n9977), .ZN(n9980)
         );
  INV_X1 U11087 ( .A(n9980), .ZN(n10039) );
  INV_X1 U11088 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9981) );
  AOI22_X1 U11089 ( .A1(n10037), .A2(n10039), .B1(n9981), .B2(n10035), .ZN(
        P1_U3460) );
  OAI22_X1 U11090 ( .A1(n9983), .A2(n10029), .B1(n9982), .B2(n10027), .ZN(
        n9985) );
  AOI211_X1 U11091 ( .C1(n10025), .C2(n9986), .A(n9985), .B(n9984), .ZN(n10040) );
  INV_X1 U11092 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9987) );
  AOI22_X1 U11093 ( .A1(n10037), .A2(n10040), .B1(n9987), .B2(n10035), .ZN(
        P1_U3463) );
  INV_X1 U11094 ( .A(n9988), .ZN(n9993) );
  OAI22_X1 U11095 ( .A1(n9990), .A2(n10029), .B1(n9989), .B2(n10027), .ZN(
        n9992) );
  AOI211_X1 U11096 ( .C1(n10025), .C2(n9993), .A(n9992), .B(n9991), .ZN(n10041) );
  INV_X1 U11097 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9994) );
  AOI22_X1 U11098 ( .A1(n10037), .A2(n10041), .B1(n9994), .B2(n10035), .ZN(
        P1_U3466) );
  NOR2_X1 U11099 ( .A1(n9996), .A2(n9995), .ZN(n10002) );
  OAI211_X1 U11100 ( .C1(n9999), .C2(n10027), .A(n9998), .B(n9997), .ZN(n10000) );
  AOI21_X1 U11101 ( .B1(n10002), .B2(n10001), .A(n10000), .ZN(n10042) );
  AOI22_X1 U11102 ( .A1(n10037), .A2(n10042), .B1(n6368), .B2(n10035), .ZN(
        P1_U3469) );
  AOI22_X1 U11103 ( .A1(n10006), .A2(n10005), .B1(n10004), .B2(n10003), .ZN(
        n10007) );
  OAI211_X1 U11104 ( .C1(n10010), .C2(n10009), .A(n10008), .B(n10007), .ZN(
        n10011) );
  INV_X1 U11105 ( .A(n10011), .ZN(n10043) );
  INV_X1 U11106 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10012) );
  AOI22_X1 U11107 ( .A1(n10037), .A2(n10043), .B1(n10012), .B2(n10035), .ZN(
        P1_U3472) );
  OAI211_X1 U11108 ( .C1(n10015), .C2(n10027), .A(n10014), .B(n10013), .ZN(
        n10016) );
  AOI21_X1 U11109 ( .B1(n10034), .B2(n10017), .A(n10016), .ZN(n10044) );
  INV_X1 U11110 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10018) );
  AOI22_X1 U11111 ( .A1(n10037), .A2(n10044), .B1(n10018), .B2(n10035), .ZN(
        P1_U3475) );
  INV_X1 U11112 ( .A(n10019), .ZN(n10024) );
  OAI22_X1 U11113 ( .A1(n10021), .A2(n10029), .B1(n4488), .B2(n10027), .ZN(
        n10023) );
  AOI211_X1 U11114 ( .C1(n10025), .C2(n10024), .A(n10023), .B(n10022), .ZN(
        n10046) );
  INV_X1 U11115 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10026) );
  AOI22_X1 U11116 ( .A1(n10037), .A2(n10046), .B1(n10026), .B2(n10035), .ZN(
        P1_U3478) );
  OAI22_X1 U11117 ( .A1(n10030), .A2(n10029), .B1(n10028), .B2(n10027), .ZN(
        n10032) );
  AOI211_X1 U11118 ( .C1(n10034), .C2(n10033), .A(n10032), .B(n10031), .ZN(
        n10048) );
  INV_X1 U11119 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10036) );
  AOI22_X1 U11120 ( .A1(n10037), .A2(n10048), .B1(n10036), .B2(n10035), .ZN(
        P1_U3481) );
  AOI22_X1 U11121 ( .A1(n10049), .A2(n10038), .B1(n6171), .B2(n10047), .ZN(
        P1_U3524) );
  AOI22_X1 U11122 ( .A1(n10049), .A2(n10039), .B1(n6264), .B2(n10047), .ZN(
        P1_U3525) );
  AOI22_X1 U11123 ( .A1(n10049), .A2(n10040), .B1(n6279), .B2(n10047), .ZN(
        P1_U3526) );
  AOI22_X1 U11124 ( .A1(n10049), .A2(n10041), .B1(n6348), .B2(n10047), .ZN(
        P1_U3527) );
  AOI22_X1 U11125 ( .A1(n10049), .A2(n10042), .B1(n6367), .B2(n10047), .ZN(
        P1_U3528) );
  AOI22_X1 U11126 ( .A1(n10049), .A2(n10043), .B1(n6501), .B2(n10047), .ZN(
        P1_U3529) );
  AOI22_X1 U11127 ( .A1(n10049), .A2(n10044), .B1(n6467), .B2(n10047), .ZN(
        P1_U3530) );
  AOI22_X1 U11128 ( .A1(n10049), .A2(n10046), .B1(n10045), .B2(n10047), .ZN(
        P1_U3531) );
  AOI22_X1 U11129 ( .A1(n10049), .A2(n10048), .B1(n6638), .B2(n10047), .ZN(
        P1_U3532) );
  AOI22_X1 U11130 ( .A1(n10055), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10050), .ZN(n10060) );
  NOR2_X1 U11131 ( .A1(n10051), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10052) );
  AOI211_X1 U11132 ( .C1(n10055), .C2(n10054), .A(n10053), .B(n10052), .ZN(
        n10058) );
  AOI22_X1 U11133 ( .A1(n10056), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(n4374), .ZN(n10057) );
  OAI221_X1 U11134 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10060), .C1(n10059), .C2(
        n10058), .A(n10057), .ZN(P2_U3245) );
  INV_X1 U11135 ( .A(n8186), .ZN(n10063) );
  OAI21_X1 U11136 ( .B1(n10063), .B2(n10062), .A(n10061), .ZN(n10070) );
  AOI22_X1 U11137 ( .A1(n10067), .A2(n10066), .B1(n10065), .B2(n10064), .ZN(
        n10068) );
  OAI21_X1 U11138 ( .B1(n10070), .B2(n10069), .A(n10068), .ZN(n10101) );
  AOI21_X1 U11139 ( .B1(n10071), .B2(P2_REG3_REG_1__SCAN_IN), .A(n10101), .ZN(
        n10079) );
  XNOR2_X1 U11140 ( .A(n8186), .B(n10072), .ZN(n10103) );
  INV_X1 U11141 ( .A(n10137), .ZN(n10153) );
  OAI211_X1 U11142 ( .C1(n10075), .C2(n4505), .A(n10138), .B(n10073), .ZN(
        n10074) );
  OAI21_X1 U11143 ( .B1(n10075), .B2(n10153), .A(n10074), .ZN(n10102) );
  AOI22_X1 U11144 ( .A1(n10103), .A2(n10077), .B1(n10102), .B2(n10076), .ZN(
        n10078) );
  OAI221_X1 U11145 ( .B1(n8646), .B2(n10079), .C1(n6401), .C2(n4949), .A(
        n10078), .ZN(P2_U3295) );
  NAND2_X1 U11146 ( .A1(n10081), .A2(n10080), .ZN(n10092) );
  AND2_X1 U11147 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10092), .ZN(P2_U3297) );
  AND2_X1 U11148 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10092), .ZN(P2_U3298) );
  INV_X1 U11149 ( .A(n10092), .ZN(n10088) );
  NOR2_X1 U11150 ( .A1(n10088), .A2(n10082), .ZN(P2_U3299) );
  AND2_X1 U11151 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10092), .ZN(P2_U3300) );
  AND2_X1 U11152 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10092), .ZN(P2_U3301) );
  NOR2_X1 U11153 ( .A1(n10088), .A2(n10083), .ZN(P2_U3302) );
  AND2_X1 U11154 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10092), .ZN(P2_U3303) );
  AND2_X1 U11155 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10092), .ZN(P2_U3304) );
  AND2_X1 U11156 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10092), .ZN(P2_U3305) );
  AND2_X1 U11157 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10092), .ZN(P2_U3306) );
  AND2_X1 U11158 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10092), .ZN(P2_U3307) );
  AND2_X1 U11159 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10092), .ZN(P2_U3308) );
  AND2_X1 U11160 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10092), .ZN(P2_U3309) );
  NOR2_X1 U11161 ( .A1(n10088), .A2(n10084), .ZN(P2_U3310) );
  AND2_X1 U11162 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10092), .ZN(P2_U3311) );
  AND2_X1 U11163 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10092), .ZN(P2_U3312) );
  AND2_X1 U11164 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10092), .ZN(P2_U3313) );
  AND2_X1 U11165 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10092), .ZN(P2_U3314) );
  AND2_X1 U11166 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10092), .ZN(P2_U3315) );
  NOR2_X1 U11167 ( .A1(n10088), .A2(n10085), .ZN(P2_U3316) );
  AND2_X1 U11168 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10092), .ZN(P2_U3317) );
  AND2_X1 U11169 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10092), .ZN(P2_U3318) );
  AND2_X1 U11170 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10092), .ZN(P2_U3319) );
  AND2_X1 U11171 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10092), .ZN(P2_U3320) );
  NOR2_X1 U11172 ( .A1(n10088), .A2(n10086), .ZN(P2_U3321) );
  AND2_X1 U11173 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10092), .ZN(P2_U3322) );
  AND2_X1 U11174 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10092), .ZN(P2_U3323) );
  AND2_X1 U11175 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10092), .ZN(P2_U3324) );
  AND2_X1 U11176 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10092), .ZN(P2_U3325) );
  NOR2_X1 U11177 ( .A1(n10088), .A2(n10087), .ZN(P2_U3326) );
  AOI22_X1 U11178 ( .A1(n10090), .A2(n10094), .B1(n10089), .B2(n10092), .ZN(
        P2_U3437) );
  INV_X1 U11179 ( .A(n10091), .ZN(n10095) );
  INV_X1 U11180 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10093) );
  AOI22_X1 U11181 ( .A1(n10095), .A2(n10094), .B1(n10093), .B2(n10092), .ZN(
        P2_U3438) );
  AOI22_X1 U11182 ( .A1(n10098), .A2(n10159), .B1(n10097), .B2(n10096), .ZN(
        n10099) );
  AND2_X1 U11183 ( .A1(n10100), .A2(n10099), .ZN(n10165) );
  AOI22_X1 U11184 ( .A1(n10163), .A2(n10165), .B1(n5193), .B2(n10161), .ZN(
        P2_U3451) );
  AOI211_X1 U11185 ( .C1(n10159), .C2(n10103), .A(n10102), .B(n10101), .ZN(
        n10166) );
  INV_X1 U11186 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10104) );
  AOI22_X1 U11187 ( .A1(n10163), .A2(n10166), .B1(n10104), .B2(n10161), .ZN(
        P2_U3454) );
  OAI22_X1 U11188 ( .A1(n10106), .A2(n10155), .B1(n10105), .B2(n10153), .ZN(
        n10108) );
  AOI211_X1 U11189 ( .C1(n10159), .C2(n10109), .A(n10108), .B(n10107), .ZN(
        n10167) );
  INV_X1 U11190 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10110) );
  AOI22_X1 U11191 ( .A1(n10163), .A2(n10167), .B1(n10110), .B2(n10161), .ZN(
        P2_U3457) );
  INV_X1 U11192 ( .A(n10142), .ZN(n10152) );
  INV_X1 U11193 ( .A(n10111), .ZN(n10115) );
  OAI22_X1 U11194 ( .A1(n10112), .A2(n10155), .B1(n4384), .B2(n10153), .ZN(
        n10114) );
  AOI211_X1 U11195 ( .C1(n10152), .C2(n10115), .A(n10114), .B(n10113), .ZN(
        n10168) );
  AOI22_X1 U11196 ( .A1(n10163), .A2(n10168), .B1(n5220), .B2(n10161), .ZN(
        P2_U3460) );
  AOI22_X1 U11197 ( .A1(n10117), .A2(n10138), .B1(n10137), .B2(n10116), .ZN(
        n10118) );
  OAI211_X1 U11198 ( .C1(n10120), .C2(n10132), .A(n10119), .B(n10118), .ZN(
        n10121) );
  INV_X1 U11199 ( .A(n10121), .ZN(n10169) );
  AOI22_X1 U11200 ( .A1(n10163), .A2(n10169), .B1(n5232), .B2(n10161), .ZN(
        P2_U3463) );
  INV_X1 U11201 ( .A(n10122), .ZN(n10127) );
  OAI211_X1 U11202 ( .C1(n10125), .C2(n10153), .A(n10124), .B(n10123), .ZN(
        n10126) );
  AOI21_X1 U11203 ( .B1(n10159), .B2(n10127), .A(n10126), .ZN(n10170) );
  AOI22_X1 U11204 ( .A1(n10163), .A2(n10170), .B1(n5246), .B2(n10161), .ZN(
        P2_U3466) );
  AOI22_X1 U11205 ( .A1(n10129), .A2(n10138), .B1(n10137), .B2(n10128), .ZN(
        n10130) );
  OAI211_X1 U11206 ( .C1(n10133), .C2(n10132), .A(n10131), .B(n10130), .ZN(
        n10134) );
  INV_X1 U11207 ( .A(n10134), .ZN(n10171) );
  INV_X1 U11208 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10135) );
  AOI22_X1 U11209 ( .A1(n10163), .A2(n10171), .B1(n10135), .B2(n10161), .ZN(
        P2_U3469) );
  AOI22_X1 U11210 ( .A1(n10139), .A2(n10138), .B1(n10137), .B2(n10136), .ZN(
        n10140) );
  OAI211_X1 U11211 ( .C1(n10143), .C2(n10142), .A(n10141), .B(n10140), .ZN(
        n10144) );
  INV_X1 U11212 ( .A(n10144), .ZN(n10172) );
  INV_X1 U11213 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10145) );
  AOI22_X1 U11214 ( .A1(n10163), .A2(n10172), .B1(n10145), .B2(n10161), .ZN(
        P2_U3475) );
  INV_X1 U11215 ( .A(n10146), .ZN(n10151) );
  OAI22_X1 U11216 ( .A1(n10148), .A2(n10155), .B1(n10147), .B2(n10153), .ZN(
        n10150) );
  AOI211_X1 U11217 ( .C1(n10152), .C2(n10151), .A(n10150), .B(n10149), .ZN(
        n10174) );
  AOI22_X1 U11218 ( .A1(n10163), .A2(n10174), .B1(n5324), .B2(n10161), .ZN(
        P2_U3481) );
  OAI22_X1 U11219 ( .A1(n10156), .A2(n10155), .B1(n10154), .B2(n10153), .ZN(
        n10158) );
  AOI211_X1 U11220 ( .C1(n10160), .C2(n10159), .A(n10158), .B(n10157), .ZN(
        n10176) );
  INV_X1 U11221 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U11222 ( .A1(n10163), .A2(n10176), .B1(n10162), .B2(n10161), .ZN(
        P2_U3487) );
  AOI22_X1 U11223 ( .A1(n10177), .A2(n10165), .B1(n10164), .B2(n10175), .ZN(
        P2_U3520) );
  AOI22_X1 U11224 ( .A1(n10177), .A2(n10166), .B1(n5994), .B2(n10175), .ZN(
        P2_U3521) );
  AOI22_X1 U11225 ( .A1(n10177), .A2(n10167), .B1(n5997), .B2(n10175), .ZN(
        P2_U3522) );
  AOI22_X1 U11226 ( .A1(n10177), .A2(n10168), .B1(n5999), .B2(n10175), .ZN(
        P2_U3523) );
  AOI22_X1 U11227 ( .A1(n10177), .A2(n10169), .B1(n6002), .B2(n10175), .ZN(
        P2_U3524) );
  AOI22_X1 U11228 ( .A1(n10177), .A2(n10170), .B1(n5250), .B2(n10175), .ZN(
        P2_U3525) );
  AOI22_X1 U11229 ( .A1(n10177), .A2(n10171), .B1(n6005), .B2(n10175), .ZN(
        P2_U3526) );
  AOI22_X1 U11230 ( .A1(n10177), .A2(n10172), .B1(n6008), .B2(n10175), .ZN(
        P2_U3528) );
  AOI22_X1 U11231 ( .A1(n10177), .A2(n10174), .B1(n10173), .B2(n10175), .ZN(
        P2_U3530) );
  AOI22_X1 U11232 ( .A1(n10177), .A2(n10176), .B1(n6019), .B2(n10175), .ZN(
        P2_U3532) );
  OAI21_X1 U11233 ( .B1(n10180), .B2(n10179), .A(n10178), .ZN(n10181) );
  XNOR2_X1 U11234 ( .A(n10181), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(ADD_1071_U5)
         );
  AOI21_X1 U11235 ( .B1(n10184), .B2(n10183), .A(n10182), .ZN(ADD_1071_U46) );
  OAI21_X1 U11236 ( .B1(n10187), .B2(n10186), .A(n10185), .ZN(ADD_1071_U56) );
  OAI21_X1 U11237 ( .B1(n10190), .B2(n10189), .A(n10188), .ZN(ADD_1071_U57) );
  OAI21_X1 U11238 ( .B1(n10193), .B2(n10192), .A(n10191), .ZN(ADD_1071_U58) );
  OAI21_X1 U11239 ( .B1(n10196), .B2(n10195), .A(n10194), .ZN(ADD_1071_U59) );
  OAI21_X1 U11240 ( .B1(n10199), .B2(n10198), .A(n10197), .ZN(ADD_1071_U60) );
  OAI21_X1 U11241 ( .B1(n10202), .B2(n10201), .A(n10200), .ZN(ADD_1071_U61) );
  AOI21_X1 U11242 ( .B1(n10205), .B2(n10204), .A(n10203), .ZN(ADD_1071_U62) );
  AOI21_X1 U11243 ( .B1(n10208), .B2(n10207), .A(n10206), .ZN(ADD_1071_U63) );
  AOI21_X1 U11244 ( .B1(n10211), .B2(n10210), .A(n10209), .ZN(ADD_1071_U50) );
  INV_X1 U11245 ( .A(n10214), .ZN(n10213) );
  OAI222_X1 U11246 ( .A1(n10216), .A2(n10215), .B1(n10216), .B2(n10214), .C1(
        n10213), .C2(n10212), .ZN(ADD_1071_U51) );
  AOI21_X1 U11247 ( .B1(n10219), .B2(n10218), .A(n10217), .ZN(ADD_1071_U49) );
  OAI21_X1 U11248 ( .B1(n10222), .B2(n10221), .A(n10220), .ZN(n10223) );
  XNOR2_X1 U11249 ( .A(n10223), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11250 ( .B1(n10226), .B2(n10225), .A(n10224), .ZN(ADD_1071_U47) );
  AOI21_X1 U11251 ( .B1(n10229), .B2(n10228), .A(n10227), .ZN(ADD_1071_U48) );
  AOI21_X1 U11252 ( .B1(n10232), .B2(n10231), .A(n10230), .ZN(ADD_1071_U54) );
  AOI21_X1 U11253 ( .B1(n10235), .B2(n10234), .A(n10233), .ZN(ADD_1071_U53) );
  OAI21_X1 U11254 ( .B1(n10238), .B2(n10237), .A(n10236), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4895 ( .A(n5191), .Z(n4503) );
  XNOR2_X1 U4919 ( .A(n5806), .B(n5805), .ZN(n8260) );
endmodule

