

module b22_C_SARLock_k_128_10 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6575, n6576, n6577, n6578, n6579, n6580, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410;

  XNOR2_X1 U7323 ( .A(n8196), .B(n8195), .ZN(n11883) );
  INV_X4 U7324 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  XNOR2_X1 U7325 ( .A(n12091), .B(n12090), .ZN(n9967) );
  OAI21_X1 U7326 ( .B1(n14463), .B2(n8174), .A(n8175), .ZN(n11749) );
  INV_X1 U7327 ( .A(n11597), .ZN(n12064) );
  AND2_X1 U7328 ( .A1(n10979), .A2(n8163), .ZN(n7534) );
  OR3_X1 U7329 ( .A1(n14305), .A2(n11695), .A3(n14301), .ZN(n10260) );
  NAND2_X2 U7330 ( .A1(n7676), .A2(n7675), .ZN(n10869) );
  NAND2_X1 U7332 ( .A1(n7162), .A2(n9235), .ZN(n9262) );
  INV_X1 U7333 ( .A(n11082), .ZN(n15080) );
  INV_X1 U7334 ( .A(n13085), .ZN(n10460) );
  INV_X1 U7335 ( .A(n9119), .ZN(n7947) );
  INV_X1 U7336 ( .A(n10167), .ZN(n7946) );
  NAND4_X2 U7337 ( .A1(n7612), .A2(n7611), .A3(n7610), .A4(n7609), .ZN(n13084)
         );
  NAND4_X2 U7338 ( .A1(n7589), .A2(n7588), .A3(n7587), .A4(n7586), .ZN(n13085)
         );
  CLKBUF_X2 U7339 ( .A(n7605), .Z(n7640) );
  AND2_X1 U7340 ( .A1(n9179), .A2(n11262), .ZN(n9856) );
  INV_X1 U7341 ( .A(n9859), .ZN(n8156) );
  INV_X1 U7342 ( .A(n9179), .ZN(n11373) );
  NAND2_X1 U7343 ( .A1(n8203), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8135) );
  MUX2_X1 U7344 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8140), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n8142) );
  AND2_X1 U7345 ( .A1(n7672), .A2(n7671), .ZN(n7801) );
  CLKBUF_X1 U7346 ( .A(n14747), .Z(n6575) );
  NOR2_X1 U7347 ( .A1(n14157), .A2(n10937), .ZN(n14747) );
  OAI21_X2 U7348 ( .B1(n11473), .B2(n7180), .A(n7177), .ZN(n9759) );
  OAI21_X2 U7349 ( .B1(n13255), .B2(n8189), .A(n8188), .ZN(n13245) );
  XNOR2_X1 U7350 ( .A(n10745), .B(n7235), .ZN(n10739) );
  CLKBUF_X1 U7351 ( .A(n11074), .Z(n6576) );
  NOR2_X1 U7352 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n9204) );
  INV_X1 U7353 ( .A(n12200), .ZN(n10834) );
  INV_X1 U7354 ( .A(n12448), .ZN(n12473) );
  AND2_X2 U7355 ( .A1(n9857), .A2(n9989), .ZN(n6580) );
  INV_X1 U7356 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8132) );
  NAND3_X1 U7358 ( .A1(n11936), .A2(n6596), .A3(n14564), .ZN(n14147) );
  INV_X1 U7359 ( .A(n8767), .ZN(n8613) );
  NAND2_X1 U7360 ( .A1(n7771), .A2(n7770), .ZN(n7774) );
  OR2_X1 U7361 ( .A1(n15139), .A2(n15140), .ZN(n15141) );
  INV_X1 U7362 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9231) );
  NAND2_X1 U7363 ( .A1(n12992), .A2(n9965), .ZN(n12091) );
  INV_X1 U7364 ( .A(n14465), .ZN(n9942) );
  OAI21_X1 U7365 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n8864), .A(n8863), .ZN(
        n8873) );
  AND2_X1 U7366 ( .A1(n9701), .A2(n9700), .ZN(n12654) );
  XNOR2_X1 U7367 ( .A(n8288), .B(n8287), .ZN(n8290) );
  XNOR2_X1 U7368 ( .A(n8827), .B(n8826), .ZN(n11695) );
  AND2_X2 U7369 ( .A1(n9857), .A2(n9989), .ZN(n6579) );
  AND2_X2 U7370 ( .A1(n9988), .A2(n15052), .ZN(n13358) );
  OAI222_X1 U7371 ( .A1(P3_U3151), .A2(n10631), .B1(n12961), .B2(n10028), .C1(
        n10027), .C2(n12962), .ZN(P3_U3293) );
  NAND4_X4 U7372 ( .A1(n8334), .A2(n8333), .A3(n8332), .A4(n8331), .ZN(n13898)
         );
  AOI21_X2 U7373 ( .B1(n15270), .B2(n9753), .A(n6637), .ZN(n15263) );
  NOR2_X2 U7374 ( .A1(n13182), .A2(n7533), .ZN(n8130) );
  NOR2_X2 U7375 ( .A1(n9503), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9523) );
  OAI21_X2 U7376 ( .B1(n7774), .B2(n6893), .A(n6891), .ZN(n7816) );
  NAND2_X2 U7377 ( .A1(n7555), .A2(n7557), .ZN(n7605) );
  AOI21_X2 U7378 ( .B1(n15257), .B2(n15256), .A(n9357), .ZN(n15245) );
  OAI21_X2 U7379 ( .B1(n11230), .B2(n7150), .A(n7148), .ZN(n15257) );
  NOR2_X2 U7380 ( .A1(n14260), .A2(n14147), .ZN(n14135) );
  NAND2_X2 U7381 ( .A1(n14057), .A2(n11931), .ZN(n14042) );
  OAI21_X2 U7382 ( .B1(n14089), .B2(n14091), .A(n11927), .ZN(n14078) );
  NAND2_X2 U7383 ( .A1(n11926), .A2(n11925), .ZN(n14089) );
  INV_X1 U7384 ( .A(n11597), .ZN(n6577) );
  INV_X1 U7385 ( .A(n11597), .ZN(n6578) );
  AND2_X1 U7386 ( .A1(n10260), .A2(n10779), .ZN(n10391) );
  INV_X1 U7387 ( .A(n10391), .ZN(n12035) );
  NAND2_X2 U7388 ( .A1(n7270), .A2(n7268), .ZN(n14697) );
  NAND2_X2 U7389 ( .A1(n13475), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7551) );
  NOR2_X2 U7390 ( .A1(n8856), .A2(n8855), .ZN(n8878) );
  BUF_X1 U7391 ( .A(n8345), .Z(n6582) );
  CLKBUF_X3 U7392 ( .A(n8345), .Z(n6583) );
  BUF_X2 U7393 ( .A(n8345), .Z(n6584) );
  NAND2_X1 U7394 ( .A1(n11966), .A2(n8290), .ZN(n8345) );
  NAND2_X1 U7395 ( .A1(n12079), .A2(n14745), .ZN(n6585) );
  NAND2_X1 U7396 ( .A1(n12079), .A2(n14745), .ZN(n6586) );
  BUF_X4 U7397 ( .A(n8484), .Z(n6588) );
  NAND2_X2 U7398 ( .A1(n7660), .A2(n7659), .ZN(n11242) );
  OAI21_X2 U7399 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n13670), .A(n8858), .ZN(
        n8874) );
  XNOR2_X2 U7400 ( .A(n13084), .B(n9871), .ZN(n10583) );
  NAND2_X2 U7401 ( .A1(n7781), .A2(n7780), .ZN(n11551) );
  NOR2_X2 U7402 ( .A1(n6746), .A2(n9254), .ZN(n10435) );
  XOR2_X2 U7403 ( .A(n8873), .B(n8872), .Z(n14621) );
  CLKBUF_X1 U7404 ( .A(n8182), .Z(n6751) );
  AOI21_X1 U7405 ( .B1(n9943), .B2(n7375), .A(n7374), .ZN(n11823) );
  NAND2_X1 U7406 ( .A1(n7792), .A2(n7791), .ZN(n11484) );
  NAND2_X1 U7407 ( .A1(n12079), .A2(n14745), .ZN(n12034) );
  INV_X2 U7408 ( .A(n10299), .ZN(n10781) );
  INV_X8 U7409 ( .A(n12036), .ZN(n12079) );
  CLKBUF_X2 U7410 ( .A(n8477), .Z(n8766) );
  NAND2_X2 U7411 ( .A1(n10260), .A2(n10388), .ZN(n12036) );
  CLKBUF_X3 U7412 ( .A(n7535), .Z(n6589) );
  CLKBUF_X2 U7413 ( .A(n7757), .Z(n9100) );
  NAND2_X1 U7415 ( .A1(n8133), .A2(n8132), .ZN(n8203) );
  NAND4_X1 U7416 ( .A1(n9207), .A2(n9206), .A3(n9205), .A4(n9204), .ZN(n9208)
         );
  OR2_X1 U7417 ( .A1(n14212), .A2(n14211), .ZN(n14273) );
  AND2_X1 U7418 ( .A1(n13051), .A2(n6897), .ZN(n13060) );
  NAND2_X1 U7419 ( .A1(n7369), .A2(n7367), .ZN(n12965) );
  NAND2_X1 U7420 ( .A1(n8020), .A2(n8019), .ZN(n13240) );
  OR2_X1 U7421 ( .A1(n14017), .A2(n14203), .ZN(n11960) );
  NAND2_X1 U7422 ( .A1(n8746), .A2(n8745), .ZN(n14203) );
  XNOR2_X1 U7423 ( .A(n12324), .B(n12637), .ZN(n12455) );
  NAND2_X1 U7424 ( .A1(n12983), .A2(n9959), .ZN(n13035) );
  NAND2_X1 U7425 ( .A1(n8721), .A2(n8720), .ZN(n14214) );
  NAND2_X1 U7426 ( .A1(n8065), .A2(n8064), .ZN(n13387) );
  NAND2_X1 U7427 ( .A1(n8708), .A2(n8707), .ZN(n14221) );
  XNOR2_X1 U7428 ( .A(n11993), .B(n11991), .ZN(n14542) );
  XNOR2_X1 U7429 ( .A(n12555), .B(n12554), .ZN(n14351) );
  AND3_X1 U7430 ( .A1(n7228), .A2(n7229), .A3(n12585), .ZN(n12555) );
  AND2_X1 U7431 ( .A1(n7215), .A2(n7214), .ZN(n14624) );
  NAND2_X1 U7432 ( .A1(n8647), .A2(n8646), .ZN(n14246) );
  OR2_X1 U7433 ( .A1(n15193), .A2(n7230), .ZN(n7228) );
  NAND2_X1 U7434 ( .A1(n7949), .A2(n7948), .ZN(n13426) );
  NAND2_X1 U7435 ( .A1(n11063), .A2(n6634), .ZN(n7365) );
  AOI21_X1 U7436 ( .B1(n11174), .B2(n6724), .A(n6906), .ZN(n6905) );
  NAND2_X1 U7437 ( .A1(n7926), .A2(n7925), .ZN(n13429) );
  NAND2_X1 U7438 ( .A1(n7804), .A2(n7803), .ZN(n14482) );
  NOR2_X1 U7439 ( .A1(n9693), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9710) );
  NAND2_X1 U7440 ( .A1(n8515), .A2(n8514), .ZN(n11799) );
  NAND2_X1 U7441 ( .A1(n10526), .A2(n10527), .ZN(n10525) );
  NAND2_X1 U7442 ( .A1(n7742), .A2(n7741), .ZN(n11339) );
  NAND2_X1 U7443 ( .A1(n7719), .A2(n7718), .ZN(n11052) );
  AOI21_X1 U7444 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n13653), .A(n8857), .ZN(
        n8910) );
  NAND2_X1 U7445 ( .A1(n10657), .A2(n15312), .ZN(n15330) );
  NAND2_X1 U7446 ( .A1(n9157), .A2(n9995), .ZN(n9993) );
  INV_X1 U7447 ( .A(n7405), .ZN(n9157) );
  CLKBUF_X2 U7448 ( .A(n10834), .Z(n12157) );
  INV_X1 U7449 ( .A(n15293), .ZN(n9277) );
  INV_X1 U7450 ( .A(n15260), .ZN(n12523) );
  AND4_X2 U7451 ( .A1(n9252), .A2(n9251), .A3(n9250), .A4(n9249), .ZN(n12819)
         );
  NAND4_X1 U7452 ( .A1(n9246), .A2(n9245), .A3(n9244), .A4(n9243), .ZN(n12817)
         );
  AND2_X1 U7453 ( .A1(n8311), .A2(n8310), .ZN(n8315) );
  BUF_X4 U7454 ( .A(n9942), .Z(n9935) );
  INV_X1 U7455 ( .A(n6812), .ZN(n14776) );
  OAI211_X1 U7456 ( .C1(n10167), .C2(n13090), .A(n7623), .B(n7622), .ZN(n9871)
         );
  NAND2_X1 U7457 ( .A1(n8337), .A2(n6611), .ZN(n6812) );
  NAND2_X1 U7458 ( .A1(n8197), .A2(n11192), .ZN(n9857) );
  BUF_X1 U7459 ( .A(n9226), .Z(n9738) );
  MUX2_X1 U7460 ( .A(n10790), .B(n11261), .S(n8777), .Z(n8544) );
  AND2_X2 U7461 ( .A1(n8290), .A2(n8298), .ZN(n8484) );
  BUF_X2 U7462 ( .A(n7583), .Z(n10167) );
  INV_X1 U7463 ( .A(n8291), .ZN(n11966) );
  MUX2_X1 U7464 ( .A(n13777), .B(n13778), .S(n7583), .Z(n10407) );
  XNOR2_X1 U7465 ( .A(n7521), .B(P1_IR_REG_30__SCAN_IN), .ZN(n8291) );
  NAND2_X1 U7466 ( .A1(n8271), .A2(n8282), .ZN(n11360) );
  INV_X1 U7467 ( .A(n8199), .ZN(n11192) );
  NAND2_X1 U7468 ( .A1(n7309), .A2(n7307), .ZN(n14650) );
  NAND2_X1 U7469 ( .A1(n14287), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7521) );
  XNOR2_X1 U7470 ( .A(n7531), .B(n9232), .ZN(n11871) );
  NAND2_X1 U7471 ( .A1(n8276), .A2(n8275), .ZN(n11261) );
  NAND2_X2 U7472 ( .A1(n8142), .A2(n8209), .ZN(n11262) );
  AND2_X2 U7473 ( .A1(n8137), .A2(n8203), .ZN(n9179) );
  OR2_X1 U7474 ( .A1(n8286), .A2(n8592), .ZN(n8288) );
  MUX2_X1 U7475 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8136), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n8137) );
  NAND2_X2 U7476 ( .A1(n8655), .A2(P1_U3086), .ZN(n14298) );
  OAI21_X1 U7477 ( .B1(n6945), .B2(n6944), .A(n8280), .ZN(n13984) );
  XNOR2_X1 U7478 ( .A(n7554), .B(n7553), .ZN(n11865) );
  NAND2_X1 U7479 ( .A1(n9784), .A2(n6594), .ZN(n6734) );
  AOI21_X1 U7480 ( .B1(n6843), .B2(n8887), .A(n6841), .ZN(n8884) );
  NOR2_X1 U7481 ( .A1(n9208), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n7161) );
  AND2_X1 U7482 ( .A1(n8263), .A2(n8261), .ZN(n7519) );
  AND2_X1 U7483 ( .A1(n7159), .A2(n9254), .ZN(n7461) );
  AND2_X1 U7484 ( .A1(n9209), .A2(n7163), .ZN(n7159) );
  AND2_X1 U7485 ( .A1(n8335), .A2(n8255), .ZN(n8352) );
  NAND4_X1 U7486 ( .A1(n7548), .A2(n8230), .A3(n8134), .A4(n8132), .ZN(n8208)
         );
  AND4_X1 U7487 ( .A1(n8254), .A2(n8253), .A3(n8252), .A4(n8251), .ZN(n8258)
         );
  AND2_X1 U7488 ( .A1(n8492), .A2(n8256), .ZN(n8257) );
  INV_X1 U7489 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7445) );
  NOR2_X1 U7490 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8492) );
  NOR2_X1 U7491 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n8251) );
  NOR2_X1 U7492 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n8253) );
  NOR2_X1 U7493 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n8252) );
  INV_X1 U7494 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8277) );
  INV_X1 U7495 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8823) );
  NOR2_X1 U7496 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n9206) );
  NOR2_X1 U7497 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n9205) );
  NOR2_X1 U7498 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n7542) );
  NOR2_X1 U7499 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7541) );
  INV_X1 U7500 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n9535) );
  INV_X1 U7501 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9496) );
  INV_X4 U7502 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7503 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n9209) );
  NOR2_X2 U7504 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n9254) );
  NOR2_X2 U7505 ( .A1(n12817), .A2(n10575), .ZN(n12822) );
  NAND3_X1 U7506 ( .A1(n11590), .A2(n8199), .A3(n11262), .ZN(n10308) );
  AND2_X2 U7507 ( .A1(n7550), .A2(n7423), .ZN(n7110) );
  NOR2_X2 U7508 ( .A1(n8208), .A2(n7549), .ZN(n7550) );
  INV_X4 U7509 ( .A(n7682), .ZN(n8109) );
  INV_X2 U7510 ( .A(n12304), .ZN(n9279) );
  NAND2_X1 U7511 ( .A1(n7978), .A2(n7439), .ZN(n7436) );
  AND2_X1 U7512 ( .A1(n11812), .A2(n11811), .ZN(n7471) );
  INV_X1 U7513 ( .A(n11871), .ZN(n7162) );
  NAND2_X1 U7514 ( .A1(n12651), .A2(n9683), .ZN(n9685) );
  NAND2_X1 U7515 ( .A1(n9215), .A2(n7476), .ZN(n7475) );
  INV_X1 U7516 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7476) );
  NOR2_X1 U7517 ( .A1(n7475), .A2(P3_IR_REG_26__SCAN_IN), .ZN(n7474) );
  NAND2_X1 U7518 ( .A1(n8190), .A2(n13246), .ZN(n7049) );
  INV_X1 U7519 ( .A(n12063), .ZN(n7503) );
  NOR2_X1 U7520 ( .A1(n11575), .A2(n6820), .ZN(n6819) );
  INV_X1 U7521 ( .A(n11535), .ZN(n6820) );
  NAND2_X1 U7522 ( .A1(n7030), .A2(n8044), .ZN(n8062) );
  NAND2_X2 U7523 ( .A1(n11871), .A2(n12959), .ZN(n12304) );
  OAI21_X1 U7524 ( .B1(n10739), .B2(n9305), .A(n6666), .ZN(n7234) );
  OR2_X1 U7525 ( .A1(n12628), .A2(n12637), .ZN(n7527) );
  OAI21_X1 U7526 ( .B1(n12762), .B2(n7157), .A(n7155), .ZN(n12739) );
  AOI21_X1 U7527 ( .B1(n7156), .B2(n12492), .A(n6645), .ZN(n7155) );
  OR2_X1 U7528 ( .A1(n9568), .A2(n9581), .ZN(n7315) );
  AND2_X1 U7529 ( .A1(n13879), .A2(n7502), .ZN(n7501) );
  OR2_X1 U7530 ( .A1(n13815), .A2(n7503), .ZN(n7502) );
  INV_X1 U7531 ( .A(n8482), .ZN(n7242) );
  AND2_X1 U7532 ( .A1(n8518), .A2(n6987), .ZN(n6986) );
  INV_X1 U7533 ( .A(n8516), .ZN(n6987) );
  INV_X1 U7534 ( .A(n8625), .ZN(n6953) );
  OAI21_X1 U7535 ( .B1(n12460), .B2(n12455), .A(n7010), .ZN(n7009) );
  AND2_X1 U7536 ( .A1(n12454), .A2(n12453), .ZN(n7010) );
  NOR2_X1 U7537 ( .A1(n7202), .A2(n7200), .ZN(n7199) );
  AND2_X1 U7538 ( .A1(n12465), .A2(n7201), .ZN(n7200) );
  NAND2_X1 U7539 ( .A1(n12901), .A2(n12612), .ZN(n6807) );
  OR2_X1 U7540 ( .A1(n7605), .A2(n10458), .ZN(n7562) );
  AND2_X1 U7541 ( .A1(n6704), .A2(n7251), .ZN(n7250) );
  NAND2_X1 U7542 ( .A1(n8722), .A2(n8725), .ZN(n7251) );
  AOI21_X1 U7543 ( .B1(n7439), .B2(n7977), .A(n7438), .ZN(n7437) );
  INV_X1 U7544 ( .A(n7994), .ZN(n7438) );
  OR2_X1 U7545 ( .A1(n7487), .A2(n12162), .ZN(n7481) );
  NAND2_X1 U7546 ( .A1(n7488), .A2(n7490), .ZN(n7487) );
  AND2_X1 U7547 ( .A1(n7468), .A2(n6685), .ZN(n7466) );
  OR2_X1 U7548 ( .A1(n12253), .A2(n12730), .ZN(n12434) );
  INV_X1 U7549 ( .A(n7141), .ZN(n7140) );
  OAI21_X1 U7550 ( .B1(n12489), .B2(n7142), .A(n9509), .ZN(n7141) );
  INV_X1 U7551 ( .A(n7183), .ZN(n7179) );
  INV_X1 U7552 ( .A(n7146), .ZN(n7145) );
  NAND2_X1 U7553 ( .A1(n12507), .A2(n12589), .ZN(n9226) );
  INV_X1 U7554 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9215) );
  INV_X1 U7555 ( .A(n9479), .ZN(n7022) );
  NAND2_X1 U7556 ( .A1(n9312), .A2(n9311), .ZN(n6797) );
  NAND2_X1 U7557 ( .A1(n9942), .A2(n13085), .ZN(n9866) );
  OR2_X1 U7558 ( .A1(n13451), .A2(n13168), .ZN(n9148) );
  NAND2_X1 U7559 ( .A1(n7583), .A2(n10005), .ZN(n8032) );
  XNOR2_X1 U7560 ( .A(n7564), .B(n7563), .ZN(n8144) );
  BUF_X1 U7561 ( .A(n8291), .Z(n8298) );
  AND2_X1 U7562 ( .A1(n7300), .A2(n11956), .ZN(n7299) );
  OR2_X1 U7563 ( .A1(n11948), .A2(n14007), .ZN(n7300) );
  NAND2_X1 U7564 ( .A1(n14118), .A2(n7386), .ZN(n7384) );
  INV_X1 U7565 ( .A(n11915), .ZN(n7266) );
  AOI21_X1 U7566 ( .B1(n7283), .B2(n7281), .A(n6669), .ZN(n7280) );
  INV_X1 U7567 ( .A(n7286), .ZN(n7281) );
  OR2_X1 U7568 ( .A1(n14537), .A2(n14834), .ZN(n6995) );
  NAND2_X1 U7569 ( .A1(n7261), .A2(n6812), .ZN(n10798) );
  NAND2_X1 U7570 ( .A1(n14776), .A2(n13898), .ZN(n8340) );
  AND2_X1 U7571 ( .A1(n10053), .A2(n10052), .ZN(n10273) );
  INV_X1 U7572 ( .A(n7974), .ZN(n7975) );
  NAND2_X1 U7573 ( .A1(n7963), .A2(n7962), .ZN(n7978) );
  AND2_X1 U7574 ( .A1(n7918), .A2(n7896), .ZN(n7916) );
  NAND2_X1 U7575 ( .A1(n7876), .A2(n7875), .ZN(n7892) );
  AOI21_X1 U7576 ( .B1(n7038), .B2(n6592), .A(n7036), .ZN(n7035) );
  INV_X1 U7577 ( .A(n7039), .ZN(n7038) );
  OAI21_X1 U7578 ( .B1(n7042), .B2(n6592), .A(n7852), .ZN(n7039) );
  INV_X1 U7579 ( .A(n6892), .ZN(n6891) );
  OAI21_X1 U7580 ( .B1(n6894), .B2(n6893), .A(n7532), .ZN(n6892) );
  INV_X1 U7581 ( .A(n7796), .ZN(n6893) );
  NAND2_X1 U7582 ( .A1(n6879), .A2(n6612), .ZN(n7771) );
  AOI21_X1 U7583 ( .B1(n7046), .B2(n7048), .A(n6668), .ZN(n7044) );
  NAND2_X1 U7584 ( .A1(n6880), .A2(n7715), .ZN(n7731) );
  NAND2_X1 U7585 ( .A1(n7713), .A2(n7712), .ZN(n6880) );
  OAI22_X1 U7586 ( .A1(n8901), .A2(n8853), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n8852), .ZN(n8854) );
  INV_X1 U7587 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n8852) );
  XNOR2_X1 U7588 ( .A(n10788), .B(n13984), .ZN(n8777) );
  NAND2_X1 U7589 ( .A1(n7490), .A2(n7492), .ZN(n7486) );
  NAND2_X1 U7590 ( .A1(n10821), .A2(n10820), .ZN(n10822) );
  NAND2_X1 U7591 ( .A1(n10850), .A2(n7463), .ZN(n10995) );
  NOR2_X1 U7592 ( .A1(n10853), .A2(n7464), .ZN(n7463) );
  INV_X1 U7593 ( .A(n10849), .ZN(n7464) );
  NAND2_X1 U7594 ( .A1(n9226), .A2(n10005), .ZN(n9430) );
  INV_X1 U7595 ( .A(n9262), .ZN(n9723) );
  AND2_X1 U7596 ( .A1(n10671), .A2(n10670), .ZN(n10672) );
  NAND2_X1 U7597 ( .A1(n12635), .A2(n9715), .ZN(n9837) );
  AOI21_X1 U7598 ( .B1(n12665), .B2(n9668), .A(n6616), .ZN(n12667) );
  AOI21_X1 U7599 ( .B1(n12715), .B2(n9627), .A(n6658), .ZN(n12700) );
  AOI21_X2 U7600 ( .B1(n12778), .B2(n12779), .A(n6707), .ZN(n12762) );
  AOI21_X1 U7601 ( .B1(n7149), .B2(n12358), .A(n6624), .ZN(n7148) );
  AND4_X1 U7602 ( .A1(n9331), .A2(n9330), .A3(n9329), .A4(n9328), .ZN(n15260)
         );
  AND4_X1 U7603 ( .A1(n9266), .A2(n9265), .A3(n9264), .A4(n9263), .ZN(n15293)
         );
  OR2_X1 U7604 ( .A1(n9281), .A2(n10437), .ZN(n9251) );
  NAND2_X1 U7605 ( .A1(n12473), .A2(n10839), .ZN(n15294) );
  OR2_X1 U7606 ( .A1(n10839), .A2(n12448), .ZN(n15292) );
  INV_X1 U7607 ( .A(n10819), .ZN(n12340) );
  NAND2_X2 U7608 ( .A1(n12509), .A2(n12340), .ZN(n12448) );
  INV_X4 U7609 ( .A(n9430), .ZN(n12319) );
  NOR2_X1 U7610 ( .A1(n9792), .A2(n11610), .ZN(n10203) );
  AND2_X1 U7611 ( .A1(n9791), .A2(n11504), .ZN(n9792) );
  OAI21_X1 U7612 ( .B1(n9718), .B2(n6774), .A(n6772), .ZN(n12315) );
  AOI21_X1 U7613 ( .B1(n6775), .B2(n6773), .A(n6607), .ZN(n6772) );
  INV_X1 U7614 ( .A(n6775), .ZN(n6774) );
  OAI21_X1 U7615 ( .B1(n7323), .B2(n6804), .A(n6802), .ZN(n9716) );
  INV_X1 U7616 ( .A(n6803), .ZN(n6802) );
  OAI21_X1 U7617 ( .B1(n6805), .B2(n6804), .A(n9705), .ZN(n6803) );
  AND2_X1 U7618 ( .A1(n9214), .A2(n7474), .ZN(n7160) );
  OAI21_X1 U7619 ( .B1(n9656), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n9655), .ZN(
        n9671) );
  XNOR2_X1 U7620 ( .A(n9732), .B(n9731), .ZN(n9809) );
  INV_X1 U7621 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n9731) );
  NAND2_X1 U7622 ( .A1(n9776), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9732) );
  NOR2_X1 U7623 ( .A1(n7027), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6786) );
  AND2_X1 U7624 ( .A1(n9615), .A2(n9599), .ZN(n9600) );
  INV_X1 U7625 ( .A(n6784), .ZN(n6783) );
  OAI21_X1 U7626 ( .B1(n6606), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n6785), .ZN(
        n6784) );
  NAND2_X1 U7627 ( .A1(n6787), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6785) );
  NAND2_X1 U7628 ( .A1(n9566), .A2(n9565), .ZN(n9568) );
  INV_X1 U7629 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n13665) );
  INV_X1 U7630 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9412) );
  NAND2_X1 U7631 ( .A1(n6795), .A2(n7340), .ZN(n9388) );
  AOI21_X1 U7632 ( .B1(n7342), .B2(n7345), .A(n7341), .ZN(n7340) );
  NAND2_X1 U7633 ( .A1(n6797), .A2(n6794), .ZN(n6795) );
  INV_X1 U7634 ( .A(n9366), .ZN(n7341) );
  INV_X1 U7635 ( .A(n9332), .ZN(n7347) );
  NAND2_X1 U7636 ( .A1(n11064), .A2(n11065), .ZN(n11063) );
  XNOR2_X1 U7637 ( .A(n6580), .B(n10869), .ZN(n9891) );
  AND2_X1 U7638 ( .A1(n9195), .A2(n9179), .ZN(n10166) );
  INV_X1 U7639 ( .A(n11865), .ZN(n7557) );
  INV_X1 U7640 ( .A(n7638), .ZN(n7757) );
  AOI21_X1 U7641 ( .B1(n7413), .B2(n7412), .A(n6630), .ZN(n7411) );
  INV_X1 U7642 ( .A(n8190), .ZN(n7412) );
  AND2_X1 U7643 ( .A1(n7523), .A2(n8008), .ZN(n7083) );
  NOR2_X1 U7644 ( .A1(n8184), .A2(n7422), .ZN(n7421) );
  INV_X1 U7645 ( .A(n8181), .ZN(n7422) );
  NAND2_X1 U7646 ( .A1(n9124), .A2(n8143), .ZN(n14456) );
  NAND2_X2 U7647 ( .A1(n7583), .A2(n7076), .ZN(n9119) );
  NAND2_X2 U7648 ( .A1(n8144), .A2(n13484), .ZN(n7583) );
  AND2_X1 U7649 ( .A1(n8212), .A2(n13768), .ZN(n15067) );
  XNOR2_X1 U7650 ( .A(n7945), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8199) );
  OAI21_X1 U7651 ( .B1(n7944), .B2(n7943), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7945) );
  AOI21_X1 U7652 ( .B1(n7501), .B2(n7503), .A(n6652), .ZN(n7499) );
  AOI21_X1 U7653 ( .B1(n7499), .B2(n6918), .A(n6917), .ZN(n6916) );
  INV_X1 U7654 ( .A(n13780), .ZN(n6917) );
  INV_X1 U7655 ( .A(n7501), .ZN(n6918) );
  OR2_X1 U7656 ( .A1(n6583), .A2(n8301), .ZN(n8303) );
  INV_X1 U7657 ( .A(n6932), .ZN(n6931) );
  AND2_X1 U7658 ( .A1(n11792), .A2(n6929), .ZN(n6928) );
  NAND2_X1 U7659 ( .A1(n6932), .A2(n6930), .ZN(n6929) );
  INV_X1 U7660 ( .A(n11638), .ZN(n6930) );
  NOR2_X1 U7661 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n8335) );
  NAND2_X1 U7662 ( .A1(n6830), .A2(n6829), .ZN(n14004) );
  AOI21_X1 U7663 ( .B1(n7391), .B2(n6646), .A(n6597), .ZN(n6829) );
  OR2_X1 U7664 ( .A1(n14075), .A2(n6831), .ZN(n6830) );
  AND2_X1 U7665 ( .A1(n14008), .A2(n14007), .ZN(n14010) );
  NAND2_X1 U7666 ( .A1(n14075), .A2(n6593), .ZN(n14052) );
  INV_X1 U7667 ( .A(n7387), .ZN(n7386) );
  OAI22_X1 U7668 ( .A1(n14132), .A2(n7388), .B1(n14260), .B2(n14146), .ZN(
        n7387) );
  NAND2_X1 U7669 ( .A1(n11896), .A2(n11895), .ZN(n7388) );
  INV_X1 U7670 ( .A(n6819), .ZN(n6818) );
  AOI21_X1 U7671 ( .B1(n6817), .B2(n6819), .A(n6656), .ZN(n6816) );
  INV_X1 U7672 ( .A(n6822), .ZN(n6817) );
  NAND2_X1 U7673 ( .A1(n6808), .A2(n11330), .ZN(n11413) );
  INV_X1 U7675 ( .A(n8683), .ZN(n8477) );
  INV_X1 U7676 ( .A(n13984), .ZN(n10937) );
  NAND2_X2 U7677 ( .A1(n8835), .A2(n14650), .ZN(n10064) );
  INV_X1 U7678 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8284) );
  AND2_X1 U7679 ( .A1(n7519), .A2(n6697), .ZN(n7396) );
  INV_X1 U7680 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7399) );
  OAI22_X1 U7681 ( .A1(n8080), .A2(n8079), .B1(n8078), .B2(n11609), .ZN(n8093)
         );
  AOI21_X1 U7682 ( .B1(n8025), .B2(n8024), .A(n8023), .ZN(n8027) );
  AND2_X1 U7683 ( .A1(n8273), .A2(n8261), .ZN(n8270) );
  AOI21_X1 U7684 ( .B1(n14954), .B2(n8911), .A(n14330), .ZN(n8913) );
  OR2_X1 U7685 ( .A1(n14620), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6858) );
  NAND2_X1 U7686 ( .A1(n10064), .A2(n10005), .ZN(n8767) );
  INV_X1 U7687 ( .A(n6583), .ZN(n8770) );
  NAND2_X1 U7688 ( .A1(n13868), .A2(n11400), .ZN(n11401) );
  MUX2_X1 U7689 ( .A(n8359), .B(n10799), .S(n8544), .Z(n8360) );
  NAND2_X1 U7690 ( .A1(n6967), .A2(n6965), .ZN(n6964) );
  NAND2_X1 U7691 ( .A1(n8469), .A2(n6966), .ZN(n6965) );
  NAND2_X1 U7692 ( .A1(n6970), .A2(n8468), .ZN(n6967) );
  INV_X1 U7693 ( .A(n8455), .ZN(n6966) );
  INV_X1 U7694 ( .A(n6972), .ZN(n6963) );
  AND2_X1 U7695 ( .A1(n8483), .A2(n7242), .ZN(n7241) );
  INV_X1 U7696 ( .A(n8432), .ZN(n7258) );
  OR2_X1 U7697 ( .A1(n6972), .A2(n6969), .ZN(n6968) );
  NOR2_X1 U7698 ( .A1(n8468), .A2(n8469), .ZN(n6969) );
  NAND2_X1 U7699 ( .A1(n9026), .A2(n9028), .ZN(n7112) );
  NAND2_X1 U7700 ( .A1(n8516), .A2(n6985), .ZN(n6984) );
  NAND2_X1 U7701 ( .A1(n6980), .A2(n6978), .ZN(n8558) );
  AND2_X1 U7702 ( .A1(n6979), .A2(n6988), .ZN(n6978) );
  NAND2_X1 U7703 ( .A1(n12447), .A2(n6635), .ZN(n12460) );
  NAND2_X1 U7704 ( .A1(n7012), .A2(n12473), .ZN(n7011) );
  NAND2_X1 U7705 ( .A1(n8697), .A2(n6948), .ZN(n6947) );
  INV_X1 U7706 ( .A(n8696), .ZN(n6948) );
  INV_X1 U7707 ( .A(n7432), .ZN(n7431) );
  OAI21_X1 U7708 ( .B1(n7891), .B2(n7433), .A(n7916), .ZN(n7432) );
  AOI21_X1 U7709 ( .B1(n7199), .B2(n7203), .A(n6664), .ZN(n7198) );
  NAND2_X1 U7710 ( .A1(n7320), .A2(n6650), .ZN(n12472) );
  OAI21_X1 U7711 ( .B1(n7321), .B2(n12463), .A(n12499), .ZN(n7320) );
  NAND2_X1 U7712 ( .A1(n9277), .A2(n10928), .ZN(n12352) );
  INV_X1 U7713 ( .A(n7335), .ZN(n7334) );
  OAI21_X1 U7714 ( .B1(n7337), .B2(n7336), .A(n9641), .ZN(n7335) );
  INV_X1 U7715 ( .A(n9628), .ZN(n7336) );
  NOR2_X1 U7716 ( .A1(n10308), .A2(n11373), .ZN(n7535) );
  NOR2_X1 U7717 ( .A1(n11573), .A2(n7284), .ZN(n7283) );
  INV_X1 U7718 ( .A(n11524), .ZN(n7284) );
  AND2_X1 U7719 ( .A1(n7046), .A2(n6882), .ZN(n6881) );
  NAND2_X1 U7720 ( .A1(n7711), .A2(n7715), .ZN(n6882) );
  NAND2_X1 U7721 ( .A1(n7443), .A2(n7442), .ZN(n7596) );
  INV_X1 U7722 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7029) );
  AOI21_X1 U7723 ( .B1(n7198), .B2(n7196), .A(n7195), .ZN(n7194) );
  INV_X1 U7724 ( .A(n7199), .ZN(n7196) );
  INV_X1 U7725 ( .A(n7198), .ZN(n7197) );
  INV_X1 U7726 ( .A(n12465), .ZN(n7203) );
  OAI21_X1 U7727 ( .B1(n7194), .B2(n6591), .A(n9836), .ZN(n6800) );
  OAI21_X1 U7728 ( .B1(n10674), .B2(n10554), .A(n10673), .ZN(n10675) );
  INV_X1 U7729 ( .A(n12404), .ZN(n7175) );
  NOR2_X1 U7730 ( .A1(n9451), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9469) );
  INV_X1 U7731 ( .A(n14422), .ZN(n7178) );
  OR2_X1 U7732 ( .A1(n9402), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9432) );
  AND2_X1 U7733 ( .A1(n12366), .A2(n12367), .ZN(n15272) );
  OR3_X1 U7734 ( .A1(n9809), .A2(n12608), .A3(n10820), .ZN(n9813) );
  NAND2_X1 U7735 ( .A1(n12352), .A2(n15286), .ZN(n9750) );
  AND3_X1 U7736 ( .A1(n9258), .A2(n9257), .A3(n9256), .ZN(n10831) );
  NAND2_X1 U7737 ( .A1(n7171), .A2(n12333), .ZN(n12707) );
  NAND2_X1 U7738 ( .A1(n12719), .A2(n12332), .ZN(n7171) );
  NOR2_X1 U7739 ( .A1(n11610), .A2(n9789), .ZN(n9985) );
  OAI21_X1 U7740 ( .B1(n9807), .B2(n9806), .A(n10203), .ZN(n9825) );
  INV_X1 U7741 ( .A(n7316), .ZN(n6787) );
  INV_X1 U7742 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n9571) );
  INV_X1 U7743 ( .A(n9570), .ZN(n9572) );
  INV_X1 U7744 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7163) );
  NAND2_X1 U7745 ( .A1(n9459), .A2(n9458), .ZN(n9460) );
  INV_X1 U7746 ( .A(n9419), .ZN(n7326) );
  INV_X1 U7747 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6748) );
  OR2_X1 U7748 ( .A1(n12108), .A2(n12107), .ZN(n12109) );
  XNOR2_X1 U7749 ( .A(n9864), .B(n11082), .ZN(n9867) );
  OR2_X1 U7750 ( .A1(n7608), .A2(n7558), .ZN(n7559) );
  NAND2_X1 U7751 ( .A1(n13202), .A2(n7103), .ZN(n7102) );
  INV_X1 U7752 ( .A(n13387), .ZN(n7103) );
  AND2_X1 U7753 ( .A1(n13230), .A2(n7066), .ZN(n7065) );
  OR2_X1 U7754 ( .A1(n13246), .A2(n7067), .ZN(n7066) );
  INV_X1 U7755 ( .A(n8043), .ZN(n7067) );
  AND2_X1 U7756 ( .A1(n13310), .A2(n7059), .ZN(n7058) );
  NAND2_X1 U7757 ( .A1(n7060), .A2(n7957), .ZN(n7059) );
  INV_X1 U7758 ( .A(n7956), .ZN(n7060) );
  NOR2_X1 U7759 ( .A1(n13437), .A2(n11829), .ZN(n7092) );
  NAND2_X1 U7760 ( .A1(n6667), .A2(n7813), .ZN(n7071) );
  NOR2_X1 U7761 ( .A1(n7073), .A2(n11459), .ZN(n7072) );
  INV_X1 U7762 ( .A(n7793), .ZN(n7073) );
  AOI21_X1 U7763 ( .B1(n11459), .B2(n7403), .A(n8170), .ZN(n7402) );
  INV_X1 U7764 ( .A(n8169), .ZN(n7403) );
  NOR2_X1 U7766 ( .A1(n13234), .A2(n7102), .ZN(n13199) );
  NOR2_X1 U7767 ( .A1(n13234), .A2(n13387), .ZN(n13221) );
  INV_X1 U7768 ( .A(n11752), .ZN(n11769) );
  INV_X1 U7769 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7423) );
  AND2_X1 U7770 ( .A1(n7373), .A2(n8131), .ZN(n6739) );
  NAND2_X1 U7771 ( .A1(n11169), .A2(n7526), .ZN(n11173) );
  AND2_X1 U7772 ( .A1(n7448), .A2(n8711), .ZN(n7447) );
  INV_X1 U7773 ( .A(n8709), .ZN(n7448) );
  NAND2_X1 U7774 ( .A1(n8748), .A2(n6977), .ZN(n6976) );
  AOI21_X1 U7775 ( .B1(n7250), .B2(n7252), .A(n6590), .ZN(n7248) );
  NAND2_X1 U7776 ( .A1(n8761), .A2(n7245), .ZN(n7244) );
  INV_X1 U7777 ( .A(n8760), .ZN(n7245) );
  OR2_X1 U7778 ( .A1(n14203), .A2(n8786), .ZN(n8787) );
  AND2_X1 U7779 ( .A1(n14041), .A2(n11902), .ZN(n7394) );
  INV_X1 U7780 ( .A(n7389), .ZN(n7382) );
  AND2_X1 U7781 ( .A1(n14132), .A2(n11920), .ZN(n7306) );
  INV_X1 U7782 ( .A(n14575), .ZN(n6990) );
  INV_X1 U7783 ( .A(n11888), .ZN(n6827) );
  INV_X1 U7784 ( .A(n7283), .ZN(n7282) );
  NOR2_X1 U7785 ( .A1(n7287), .A2(n11525), .ZN(n7286) );
  INV_X1 U7786 ( .A(n11409), .ZN(n7287) );
  AND2_X1 U7787 ( .A1(n11313), .A2(n7273), .ZN(n7272) );
  NAND2_X1 U7788 ( .A1(n7277), .A2(n7275), .ZN(n7273) );
  INV_X1 U7789 ( .A(n11315), .ZN(n7269) );
  NAND2_X1 U7790 ( .A1(n14811), .A2(n13893), .ZN(n7275) );
  NAND2_X1 U7791 ( .A1(n10781), .A2(n10392), .ZN(n10796) );
  NAND2_X1 U7792 ( .A1(n6828), .A2(n11686), .ZN(n11889) );
  INV_X1 U7793 ( .A(n11688), .ZN(n6828) );
  AND2_X1 U7794 ( .A1(n14770), .A2(n10953), .ZN(n10955) );
  NAND2_X1 U7795 ( .A1(n8269), .A2(n6943), .ZN(n6942) );
  INV_X1 U7796 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6943) );
  INV_X1 U7797 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8261) );
  NOR2_X1 U7798 ( .A1(n8578), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n8593) );
  INV_X1 U7799 ( .A(n7729), .ZN(n7730) );
  NAND2_X1 U7800 ( .A1(n7695), .A2(n7694), .ZN(n7713) );
  XNOR2_X1 U7801 ( .A(n6844), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n8885) );
  NOR2_X1 U7802 ( .A1(n8842), .A2(n8841), .ZN(n8844) );
  AND2_X1 U7803 ( .A1(n8840), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n8841) );
  NOR2_X1 U7804 ( .A1(n8847), .A2(n8846), .ZN(n8849) );
  INV_X1 U7805 ( .A(n7211), .ZN(n8845) );
  XNOR2_X1 U7806 ( .A(n8849), .B(n8848), .ZN(n8897) );
  AND3_X1 U7807 ( .A1(n9356), .A2(n9355), .A3(n9354), .ZN(n11203) );
  NOR2_X1 U7808 ( .A1(n7481), .A2(n12701), .ZN(n7479) );
  INV_X1 U7809 ( .A(n7481), .ZN(n7480) );
  AND3_X1 U7810 ( .A1(n9276), .A2(n9275), .A3(n9274), .ZN(n10843) );
  INV_X1 U7811 ( .A(n12455), .ZN(n12497) );
  AND2_X1 U7812 ( .A1(n6870), .A2(n12149), .ZN(n6869) );
  NAND2_X1 U7813 ( .A1(n12255), .A2(n6871), .ZN(n6870) );
  INV_X1 U7814 ( .A(n12255), .ZN(n6872) );
  INV_X1 U7815 ( .A(n11305), .ZN(n7459) );
  INV_X1 U7816 ( .A(n7458), .ZN(n7457) );
  OAI21_X1 U7817 ( .B1(n11302), .B2(n7459), .A(n11423), .ZN(n7458) );
  NAND2_X1 U7818 ( .A1(n6863), .A2(n7465), .ZN(n11710) );
  AOI21_X1 U7819 ( .B1(n11445), .B2(n11430), .A(n6661), .ZN(n7465) );
  NAND2_X1 U7820 ( .A1(n11429), .A2(n11445), .ZN(n6863) );
  INV_X1 U7821 ( .A(n7493), .ZN(n7491) );
  NAND2_X1 U7822 ( .A1(n7493), .A2(n12161), .ZN(n7492) );
  NAND2_X1 U7823 ( .A1(n6859), .A2(n12132), .ZN(n12287) );
  NAND2_X1 U7824 ( .A1(n7467), .A2(n7466), .ZN(n6859) );
  OR2_X1 U7825 ( .A1(n12304), .A2(n9236), .ZN(n9237) );
  OR2_X1 U7826 ( .A1(n9304), .A2(n10656), .ZN(n9244) );
  AND2_X1 U7827 ( .A1(n10428), .A2(n10546), .ZN(n10541) );
  OAI21_X1 U7828 ( .B1(n12572), .B2(n12571), .A(n12570), .ZN(n15168) );
  NAND2_X1 U7829 ( .A1(n15168), .A2(n15167), .ZN(n15166) );
  NAND2_X1 U7830 ( .A1(n15141), .A2(n12549), .ZN(n6741) );
  NOR2_X1 U7831 ( .A1(n12529), .A2(n11626), .ZN(n6749) );
  XOR2_X1 U7832 ( .A(n12537), .B(n15199), .Z(n15196) );
  AND2_X1 U7833 ( .A1(n15187), .A2(n12578), .ZN(n15204) );
  NAND2_X1 U7834 ( .A1(n14367), .A2(n6722), .ZN(n7219) );
  NAND2_X1 U7835 ( .A1(n7221), .A2(n6722), .ZN(n7220) );
  OR2_X1 U7836 ( .A1(n12618), .A2(n9711), .ZN(n12626) );
  NOR2_X1 U7837 ( .A1(n6622), .A2(n7168), .ZN(n7167) );
  NAND2_X1 U7838 ( .A1(n12707), .A2(n12706), .ZN(n12709) );
  OR2_X1 U7839 ( .A1(n9632), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9647) );
  AND2_X1 U7840 ( .A1(n12335), .A2(n12334), .ZN(n12732) );
  NOR2_X1 U7841 ( .A1(n12744), .A2(n7191), .ZN(n7190) );
  INV_X1 U7842 ( .A(n12430), .ZN(n7191) );
  NAND2_X1 U7843 ( .A1(n12762), .A2(n9562), .ZN(n12761) );
  AND4_X1 U7844 ( .A1(n9561), .A2(n9560), .A3(n9559), .A4(n9558), .ZN(n12781)
         );
  OR2_X1 U7845 ( .A1(n12944), .A2(n12791), .ZN(n12794) );
  AOI21_X1 U7846 ( .B1(n7140), .B2(n7142), .A(n6714), .ZN(n7138) );
  AND2_X1 U7847 ( .A1(n12794), .A2(n12409), .ZN(n12808) );
  NAND2_X1 U7848 ( .A1(n11740), .A2(n12489), .ZN(n11739) );
  OR2_X1 U7849 ( .A1(n11667), .A2(n9761), .ZN(n7174) );
  NAND2_X1 U7850 ( .A1(n7134), .A2(n7135), .ZN(n11664) );
  AOI21_X1 U7851 ( .B1(n9457), .B2(n7136), .A(n6711), .ZN(n7135) );
  NAND2_X1 U7852 ( .A1(n7137), .A2(n6608), .ZN(n11619) );
  INV_X1 U7853 ( .A(n14423), .ZN(n7137) );
  NOR2_X1 U7854 ( .A1(n7184), .A2(n9758), .ZN(n7183) );
  INV_X1 U7855 ( .A(n12381), .ZN(n7184) );
  AOI21_X1 U7856 ( .B1(n7183), .B2(n9757), .A(n7182), .ZN(n7181) );
  INV_X1 U7857 ( .A(n12384), .ZN(n7182) );
  AND2_X1 U7858 ( .A1(n12390), .A2(n12389), .ZN(n14422) );
  NAND2_X1 U7859 ( .A1(n9756), .A2(n12377), .ZN(n11473) );
  AND3_X1 U7860 ( .A1(n9374), .A2(n9373), .A3(n9372), .ZN(n15251) );
  AOI21_X2 U7861 ( .B1(n15291), .B2(n15290), .A(n7524), .ZN(n11230) );
  NAND2_X1 U7862 ( .A1(n11230), .A2(n9323), .ZN(n11229) );
  INV_X1 U7863 ( .A(n7152), .ZN(n7151) );
  OAI21_X1 U7864 ( .B1(n9430), .B2(n10032), .A(n7154), .ZN(n7152) );
  INV_X1 U7865 ( .A(n15299), .ZN(n15319) );
  NAND2_X1 U7866 ( .A1(n9605), .A2(n9604), .ZN(n12209) );
  OR2_X1 U7867 ( .A1(n10934), .A2(n9603), .ZN(n9605) );
  NAND2_X1 U7868 ( .A1(n9589), .A2(n9588), .ZN(n12253) );
  OR2_X1 U7869 ( .A1(n10752), .A2(n9603), .ZN(n9589) );
  INV_X1 U7870 ( .A(SI_15_), .ZN(n9500) );
  OR2_X1 U7871 ( .A1(n12951), .A2(n9985), .ZN(n10654) );
  INV_X1 U7872 ( .A(n15294), .ZN(n15322) );
  NOR2_X1 U7873 ( .A1(n9686), .A2(n6806), .ZN(n6805) );
  INV_X1 U7874 ( .A(n9672), .ZN(n6806) );
  INV_X1 U7875 ( .A(n7475), .ZN(n7473) );
  NAND2_X1 U7876 ( .A1(n9671), .A2(n9670), .ZN(n7323) );
  AOI21_X1 U7877 ( .B1(n7315), .B2(n6783), .A(n6780), .ZN(n6779) );
  NAND2_X1 U7878 ( .A1(n6781), .A2(n9600), .ZN(n6780) );
  NAND2_X1 U7879 ( .A1(n6783), .A2(n6786), .ZN(n6781) );
  INV_X1 U7880 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9734) );
  NAND2_X1 U7881 ( .A1(n7315), .A2(n6606), .ZN(n9585) );
  OAI21_X1 U7882 ( .B1(n6782), .B2(n6787), .A(P1_DATAO_REG_20__SCAN_IN), .ZN(
        n9597) );
  INV_X1 U7883 ( .A(n7315), .ZN(n6782) );
  NAND2_X1 U7884 ( .A1(n6790), .A2(n6788), .ZN(n9566) );
  AOI21_X1 U7885 ( .B1(n6791), .B2(n6793), .A(n6789), .ZN(n6788) );
  INV_X1 U7886 ( .A(n9551), .ZN(n6789) );
  AND2_X1 U7887 ( .A1(n9532), .A2(n9514), .ZN(n9515) );
  NAND2_X1 U7888 ( .A1(n9516), .A2(n9515), .ZN(n9533) );
  NAND2_X1 U7889 ( .A1(n7020), .A2(n7019), .ZN(n9511) );
  AND2_X1 U7890 ( .A1(n7018), .A2(n9493), .ZN(n7019) );
  NAND2_X1 U7891 ( .A1(n7311), .A2(n7021), .ZN(n7020) );
  OR2_X1 U7892 ( .A1(n9476), .A2(n7022), .ZN(n7018) );
  AND2_X1 U7893 ( .A1(n9512), .A2(n9495), .ZN(n9510) );
  NAND2_X1 U7894 ( .A1(n9460), .A2(n10321), .ZN(n9476) );
  NAND2_X1 U7895 ( .A1(n9477), .A2(n9476), .ZN(n9480) );
  AND2_X1 U7896 ( .A1(n9493), .A2(n9478), .ZN(n9479) );
  INV_X1 U7897 ( .A(n9461), .ZN(n7311) );
  INV_X1 U7898 ( .A(n9208), .ZN(n7462) );
  NAND2_X1 U7899 ( .A1(n7311), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9477) );
  NAND2_X1 U7900 ( .A1(n7006), .A2(n9476), .ZN(n9461) );
  NAND2_X1 U7901 ( .A1(n7007), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7006) );
  INV_X1 U7902 ( .A(n9460), .ZN(n7007) );
  AOI21_X1 U7903 ( .B1(n9392), .B2(n7329), .A(n7328), .ZN(n7327) );
  INV_X1 U7904 ( .A(n9409), .ZN(n7328) );
  INV_X1 U7905 ( .A(n9389), .ZN(n7329) );
  INV_X1 U7906 ( .A(n9392), .ZN(n7330) );
  NAND2_X1 U7907 ( .A1(n9388), .A2(n9387), .ZN(n9390) );
  AOI21_X1 U7908 ( .B1(n9333), .B2(n7346), .A(n6602), .ZN(n7345) );
  INV_X1 U7909 ( .A(n9334), .ZN(n7349) );
  NAND2_X1 U7910 ( .A1(n6797), .A2(n9313), .ZN(n9334) );
  NAND2_X1 U7911 ( .A1(n9292), .A2(n9291), .ZN(n9312) );
  INV_X1 U7912 ( .A(n9929), .ZN(n7363) );
  AND2_X1 U7913 ( .A1(n9870), .A2(n9863), .ZN(n7353) );
  AOI21_X1 U7914 ( .B1(n9877), .B2(n9876), .A(n7525), .ZN(n13020) );
  AND2_X1 U7915 ( .A1(n9922), .A2(n9916), .ZN(n7364) );
  INV_X1 U7916 ( .A(n11590), .ZN(n9195) );
  AOI21_X1 U7917 ( .B1(n14988), .B2(P2_REG1_REG_14__SCAN_IN), .A(n14980), .ZN(
        n13133) );
  AND2_X1 U7918 ( .A1(n7101), .A2(n7097), .ZN(n13172) );
  INV_X1 U7919 ( .A(n13234), .ZN(n7101) );
  AND2_X1 U7920 ( .A1(n7100), .A2(n7098), .ZN(n7097) );
  INV_X1 U7921 ( .A(n7102), .ZN(n7100) );
  NOR3_X1 U7922 ( .A1(n7104), .A2(n7102), .A3(n13234), .ZN(n13188) );
  OR2_X1 U7923 ( .A1(n13387), .A2(n13065), .ZN(n7034) );
  AND2_X1 U7924 ( .A1(n7411), .A2(n6684), .ZN(n6737) );
  NAND2_X1 U7925 ( .A1(n8034), .A2(n8033), .ZN(n13249) );
  NAND2_X1 U7926 ( .A1(n6752), .A2(n7414), .ZN(n13243) );
  INV_X1 U7927 ( .A(n13246), .ZN(n7414) );
  XNOR2_X1 U7928 ( .A(n13249), .B(n13067), .ZN(n13246) );
  OR2_X1 U7929 ( .A1(n7093), .A2(n13426), .ZN(n13321) );
  NAND2_X1 U7930 ( .A1(n7934), .A2(n7933), .ZN(n13318) );
  OR2_X1 U7931 ( .A1(n14464), .A2(n11841), .ZN(n11752) );
  NAND2_X1 U7932 ( .A1(n6743), .A2(n7072), .ZN(n11462) );
  AOI21_X1 U7933 ( .B1(n7408), .B2(n7410), .A(n6625), .ZN(n7407) );
  NAND2_X1 U7934 ( .A1(n11210), .A2(n7749), .ZN(n11344) );
  NAND2_X1 U7935 ( .A1(n7534), .A2(n11045), .ZN(n11044) );
  NAND2_X1 U7936 ( .A1(n9121), .A2(n9120), .ZN(n13165) );
  NAND2_X1 U7937 ( .A1(n7998), .A2(n7997), .ZN(n13409) );
  NAND3_X1 U7938 ( .A1(n8138), .A2(n7110), .A3(n7563), .ZN(n7109) );
  INV_X1 U7939 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7553) );
  NAND4_X1 U7940 ( .A1(n7599), .A2(n7108), .A3(n7107), .A4(n7106), .ZN(n7631)
         );
  INV_X1 U7941 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7108) );
  INV_X1 U7942 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7107) );
  INV_X1 U7943 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7106) );
  INV_X2 U7944 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7599) );
  NAND2_X1 U7945 ( .A1(n11639), .A2(n11638), .ZN(n6933) );
  AOI21_X1 U7946 ( .B1(n6916), .B2(n6919), .A(n6654), .ZN(n6914) );
  INV_X1 U7947 ( .A(n7499), .ZN(n6919) );
  AND2_X1 U7948 ( .A1(n10394), .A2(n10393), .ZN(n10395) );
  OR2_X1 U7949 ( .A1(n10781), .A2(n6585), .ZN(n10394) );
  XNOR2_X1 U7950 ( .A(n6903), .B(n10389), .ZN(n10396) );
  OAI22_X1 U7951 ( .A1(n12035), .A2(n10781), .B1(n14770), .B2(n12036), .ZN(
        n6903) );
  NAND2_X1 U7952 ( .A1(n6935), .A2(n6600), .ZN(n13805) );
  NAND2_X1 U7953 ( .A1(n7511), .A2(n6936), .ZN(n6935) );
  INV_X1 U7954 ( .A(n14506), .ZN(n7497) );
  NOR2_X1 U7955 ( .A1(n7497), .A2(n7498), .ZN(n7496) );
  INV_X1 U7956 ( .A(n14543), .ZN(n7498) );
  AND2_X1 U7957 ( .A1(n13787), .A2(n7507), .ZN(n7506) );
  OR2_X1 U7958 ( .A1(n13852), .A2(n7508), .ZN(n7507) );
  INV_X1 U7959 ( .A(n12042), .ZN(n7508) );
  XNOR2_X1 U7960 ( .A(n11173), .B(n11171), .ZN(n11254) );
  NAND2_X1 U7961 ( .A1(n10269), .A2(n10268), .ZN(n10270) );
  INV_X1 U7962 ( .A(n10267), .ZN(n10268) );
  NAND2_X1 U7963 ( .A1(n10266), .A2(n10265), .ZN(n10269) );
  OAI22_X1 U7964 ( .A1(n12035), .A2(n10953), .B1(n10260), .B2(n13900), .ZN(
        n10267) );
  NAND2_X1 U7965 ( .A1(n13860), .A2(n13861), .ZN(n7511) );
  NAND2_X1 U7966 ( .A1(n10395), .A2(n10396), .ZN(n10496) );
  NAND2_X1 U7967 ( .A1(n6921), .A2(n6925), .ZN(n6924) );
  INV_X1 U7968 ( .A(n10502), .ZN(n6925) );
  NAND2_X1 U7969 ( .A1(n14498), .A2(n11987), .ZN(n11993) );
  OR2_X1 U7970 ( .A1(n8701), .A2(n11250), .ZN(n8370) );
  NAND2_X1 U7971 ( .A1(n8769), .A2(n8768), .ZN(n13998) );
  NAND2_X1 U7972 ( .A1(n8759), .A2(n8758), .ZN(n11937) );
  AND2_X1 U7973 ( .A1(n7299), .A2(n11935), .ZN(n7289) );
  NAND2_X1 U7974 ( .A1(n7293), .A2(n7295), .ZN(n7292) );
  INV_X1 U7975 ( .A(n7299), .ZN(n7293) );
  INV_X1 U7976 ( .A(n11935), .ZN(n7295) );
  AOI21_X1 U7977 ( .B1(n7299), .B2(n11948), .A(n7298), .ZN(n7297) );
  INV_X1 U7978 ( .A(n11934), .ZN(n7298) );
  INV_X1 U7979 ( .A(n14007), .ZN(n11904) );
  NAND2_X1 U7980 ( .A1(n14052), .A2(n7394), .ZN(n14040) );
  INV_X1 U7981 ( .A(n14077), .ZN(n11899) );
  OAI21_X1 U7982 ( .B1(n14114), .B2(n11923), .A(n11897), .ZN(n14092) );
  NAND2_X1 U7983 ( .A1(n14092), .A2(n14091), .ZN(n14090) );
  NOR2_X1 U7984 ( .A1(n14132), .A2(n7390), .ZN(n7389) );
  INV_X1 U7985 ( .A(n7384), .ZN(n7383) );
  AND2_X1 U7986 ( .A1(n8635), .A2(n8634), .ZN(n13799) );
  NAND2_X1 U7987 ( .A1(n11921), .A2(n7306), .ZN(n14131) );
  NAND2_X1 U7988 ( .A1(n11893), .A2(n11892), .ZN(n14153) );
  NAND2_X1 U7989 ( .A1(n14162), .A2(n11918), .ZN(n14144) );
  AOI21_X1 U7990 ( .B1(n7265), .B2(n14567), .A(n6653), .ZN(n7264) );
  OR2_X1 U7991 ( .A1(n14592), .A2(n14493), .ZN(n11915) );
  NAND2_X1 U7992 ( .A1(n11913), .A2(n11912), .ZN(n14563) );
  NAND2_X1 U7993 ( .A1(n6816), .A2(n6818), .ZN(n6815) );
  NOR2_X1 U7994 ( .A1(n11533), .A2(n6823), .ZN(n6822) );
  INV_X1 U7995 ( .A(n11414), .ZN(n6823) );
  NAND2_X1 U7996 ( .A1(n11410), .A2(n7286), .ZN(n7285) );
  NAND2_X1 U7997 ( .A1(n6810), .A2(n11110), .ZN(n11264) );
  NAND2_X1 U7998 ( .A1(n10796), .A2(n10794), .ZN(n10958) );
  NOR2_X1 U7999 ( .A1(n8285), .A2(n7308), .ZN(n7307) );
  OR2_X1 U8000 ( .A1(n7397), .A2(n7310), .ZN(n7309) );
  NOR2_X1 U8001 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n7308) );
  OR2_X1 U8002 ( .A1(n6997), .A2(n13999), .ZN(n6996) );
  INV_X1 U8003 ( .A(n6998), .ZN(n6997) );
  AOI21_X1 U8004 ( .B1(n11960), .B2(n11937), .A(n14745), .ZN(n6998) );
  AND2_X1 U8005 ( .A1(n11961), .A2(n11960), .ZN(n14202) );
  NAND2_X1 U8006 ( .A1(n8615), .A2(n8614), .ZN(n14260) );
  NAND2_X1 U8007 ( .A1(n8481), .A2(n8480), .ZN(n14834) );
  AND2_X1 U8008 ( .A1(n8467), .A2(n8466), .ZN(n14825) );
  AND2_X1 U8009 ( .A1(n10275), .A2(n10274), .ZN(n11583) );
  AND2_X1 U8010 ( .A1(n10260), .A2(n10054), .ZN(n10302) );
  OR2_X1 U8011 ( .A1(n8763), .A2(n8762), .ZN(n8765) );
  INV_X1 U8012 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8287) );
  OR2_X1 U8013 ( .A1(n8285), .A2(n8592), .ZN(n8264) );
  XNOR2_X1 U8014 ( .A(n8099), .B(n8115), .ZN(n11876) );
  NAND2_X1 U8015 ( .A1(n8119), .A2(n8117), .ZN(n8099) );
  NOR2_X1 U8016 ( .A1(n8828), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n7397) );
  OAI21_X1 U8017 ( .B1(n8062), .B2(n8061), .A(n8060), .ZN(n8080) );
  NAND2_X1 U8018 ( .A1(n8030), .A2(n8029), .ZN(n7030) );
  NOR2_X1 U8019 ( .A1(n6942), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n6941) );
  NAND2_X1 U8020 ( .A1(n8283), .A2(n6662), .ZN(n10788) );
  INV_X1 U8021 ( .A(n7976), .ZN(n7440) );
  OR2_X1 U8022 ( .A1(n7978), .A2(n7977), .ZN(n7441) );
  CLKBUF_X1 U8023 ( .A(n8272), .Z(n8273) );
  NAND2_X1 U8024 ( .A1(n7430), .A2(n7893), .ZN(n7917) );
  NAND2_X1 U8025 ( .A1(n7892), .A2(n7891), .ZN(n7430) );
  OAI21_X1 U8026 ( .B1(n7816), .B2(n6592), .A(n7038), .ZN(n7874) );
  XNOR2_X1 U8027 ( .A(n8522), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11281) );
  NAND2_X1 U8028 ( .A1(n7041), .A2(n7832), .ZN(n7854) );
  NAND2_X1 U8029 ( .A1(n7816), .A2(n7042), .ZN(n7041) );
  INV_X1 U8030 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8255) );
  INV_X2 U8031 ( .A(n7076), .ZN(n8655) );
  XNOR2_X1 U8032 ( .A(n7592), .B(SI_1_), .ZN(n7590) );
  AND2_X1 U8033 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n6842), .ZN(n8887) );
  NAND2_X1 U8034 ( .A1(n15397), .A2(n15396), .ZN(n8895) );
  NAND2_X1 U8035 ( .A1(n6839), .A2(n6838), .ZN(n8918) );
  NAND2_X1 U8036 ( .A1(n14618), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n6838) );
  NAND2_X1 U8037 ( .A1(n6837), .A2(n6647), .ZN(n6839) );
  AOI22_X1 U8038 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n8866), .B1(n8873), .B2(
        n8865), .ZN(n8922) );
  AOI21_X1 U8039 ( .B1(n15031), .B2(n8930), .A(n14346), .ZN(n8935) );
  NAND2_X1 U8040 ( .A1(n11201), .A2(n11200), .ZN(n11303) );
  NAND2_X1 U8041 ( .A1(n9692), .A2(n9691), .ZN(n12836) );
  AND2_X1 U8042 ( .A1(n9654), .A2(n9653), .ZN(n12244) );
  NAND2_X1 U8043 ( .A1(n7026), .A2(n9631), .ZN(n12705) );
  NAND2_X1 U8044 ( .A1(n11195), .A2(n12318), .ZN(n7026) );
  NAND2_X1 U8045 ( .A1(n11427), .A2(n11426), .ZN(n11448) );
  INV_X1 U8046 ( .A(n11429), .ZN(n11427) );
  AND2_X1 U8047 ( .A1(n9416), .A2(n9415), .ZN(n11454) );
  AND3_X1 U8048 ( .A1(n9594), .A2(n9593), .A3(n9592), .ZN(n12730) );
  NAND2_X1 U8049 ( .A1(n12192), .A2(n12191), .ZN(n12190) );
  NAND2_X1 U8050 ( .A1(n9708), .A2(n9707), .ZN(n12324) );
  NAND2_X1 U8051 ( .A1(n9659), .A2(n9658), .ZN(n12845) );
  NAND2_X1 U8052 ( .A1(n12288), .A2(n12135), .ZN(n12226) );
  NAND2_X1 U8053 ( .A1(n10996), .A2(n10997), .ZN(n11139) );
  AND2_X1 U8054 ( .A1(n9667), .A2(n9666), .ZN(n12653) );
  NAND2_X1 U8055 ( .A1(n10836), .A2(n10884), .ZN(n10850) );
  AND3_X1 U8056 ( .A1(n9580), .A2(n9579), .A3(n9578), .ZN(n12741) );
  INV_X1 U8057 ( .A(n12687), .ZN(n12717) );
  NAND2_X1 U8058 ( .A1(n9618), .A2(n9617), .ZN(n12720) );
  NAND2_X1 U8059 ( .A1(n10885), .A2(n10886), .ZN(n10884) );
  AND4_X1 U8060 ( .A1(n9347), .A2(n9346), .A3(n9345), .A4(n9344), .ZN(n11309)
         );
  NAND2_X1 U8061 ( .A1(n6865), .A2(n7490), .ZN(n6864) );
  NAND2_X1 U8062 ( .A1(n7494), .A2(n7484), .ZN(n6865) );
  INV_X1 U8063 ( .A(n7492), .ZN(n7484) );
  INV_X1 U8064 ( .A(n12298), .ZN(n12282) );
  NAND2_X1 U8065 ( .A1(n10475), .A2(n10474), .ZN(n12285) );
  AND4_X1 U8066 ( .A1(n9529), .A2(n9528), .A3(n9527), .A4(n9526), .ZN(n12807)
         );
  OR2_X1 U8067 ( .A1(n12322), .A2(n12323), .ZN(n7025) );
  NAND2_X1 U8068 ( .A1(n9682), .A2(n9681), .ZN(n12670) );
  INV_X1 U8069 ( .A(n12653), .ZN(n12688) );
  INV_X1 U8070 ( .A(n12244), .ZN(n12702) );
  INV_X1 U8071 ( .A(n12730), .ZN(n12752) );
  INV_X1 U8072 ( .A(n12781), .ZN(n12751) );
  INV_X1 U8073 ( .A(n15233), .ZN(n15247) );
  INV_X1 U8074 ( .A(n11309), .ZN(n15277) );
  OAI22_X1 U8075 ( .A1(n10536), .A2(n10535), .B1(n10534), .B2(n10546), .ZN(
        n10720) );
  INV_X1 U8076 ( .A(n10543), .ZN(n7233) );
  XNOR2_X1 U8077 ( .A(n6741), .B(n15163), .ZN(n15158) );
  INV_X1 U8078 ( .A(n12601), .ZN(n7222) );
  NAND2_X1 U8079 ( .A1(n12597), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7224) );
  AND2_X1 U8080 ( .A1(n10432), .A2(n10424), .ZN(n15151) );
  NAND2_X1 U8081 ( .A1(n14405), .A2(n6764), .ZN(n6763) );
  OR2_X1 U8082 ( .A1(n14404), .A2(n12563), .ZN(n6764) );
  OR2_X1 U8083 ( .A1(n12604), .A2(n15184), .ZN(n6732) );
  NOR2_X1 U8084 ( .A1(n12607), .A2(n6731), .ZN(n6730) );
  AND2_X1 U8085 ( .A1(n15149), .A2(n12608), .ZN(n6731) );
  OR2_X1 U8086 ( .A1(n9842), .A2(n9841), .ZN(n12625) );
  NAND2_X1 U8087 ( .A1(n9675), .A2(n9674), .ZN(n12840) );
  AND3_X1 U8088 ( .A1(n9399), .A2(n9398), .A3(n9397), .ZN(n11480) );
  NAND2_X1 U8089 ( .A1(n12301), .A2(n12300), .ZN(n12901) );
  INV_X1 U8090 ( .A(n12324), .ZN(n12628) );
  NAND2_X1 U8091 ( .A1(n9542), .A2(n9541), .ZN(n12939) );
  NAND2_X1 U8092 ( .A1(n9485), .A2(n9484), .ZN(n12948) );
  AND2_X1 U8093 ( .A1(n9795), .A2(n9794), .ZN(n12950) );
  AOI21_X1 U8094 ( .B1(n10203), .B2(n9796), .A(n6655), .ZN(n12952) );
  INV_X1 U8095 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7204) );
  MUX2_X1 U8096 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9216), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n9218) );
  OR2_X1 U8097 ( .A1(n9221), .A2(n9231), .ZN(n9216) );
  MUX2_X1 U8098 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9220), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n9222) );
  INV_X1 U8099 ( .A(n9809), .ZN(n12509) );
  OR2_X1 U8100 ( .A1(n7638), .A2(n10173), .ZN(n7580) );
  OR2_X1 U8101 ( .A1(n7608), .A2(n10174), .ZN(n7577) );
  OR2_X1 U8102 ( .A1(n9944), .A2(n11699), .ZN(n7375) );
  AND2_X1 U8103 ( .A1(n9944), .A2(n11699), .ZN(n7374) );
  NAND2_X1 U8104 ( .A1(n7966), .A2(n7965), .ZN(n13420) );
  NAND2_X1 U8105 ( .A1(n10406), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14453) );
  NAND2_X1 U8106 ( .A1(n9972), .A2(n15052), .ZN(n14451) );
  INV_X1 U8107 ( .A(n13053), .ZN(n13064) );
  OR2_X1 U8108 ( .A1(n7605), .A2(n10450), .ZN(n7588) );
  OAI21_X1 U8109 ( .B1(n15050), .B2(n13638), .A(n13164), .ZN(n6758) );
  CLKBUF_X1 U8110 ( .A(n8199), .Z(n13161) );
  INV_X1 U8111 ( .A(n8152), .ZN(n8153) );
  AOI21_X1 U8112 ( .B1(n13063), .B2(n13335), .A(n8151), .ZN(n8152) );
  NAND2_X1 U8113 ( .A1(n8046), .A2(n8045), .ZN(n13392) );
  OR3_X1 U8114 ( .A1(n13358), .A2(n6579), .A3(n11014), .ZN(n13365) );
  OR2_X1 U8115 ( .A1(n13358), .A2(n9999), .ZN(n13360) );
  INV_X1 U8116 ( .A(n15061), .ZN(n14467) );
  NAND2_X1 U8117 ( .A1(n9099), .A2(n9098), .ZN(n13451) );
  NAND2_X1 U8118 ( .A1(n7077), .A2(n7076), .ZN(n7075) );
  AND2_X1 U8119 ( .A1(n8235), .A2(n8234), .ZN(n15074) );
  NAND2_X1 U8120 ( .A1(n8675), .A2(n8674), .ZN(n14235) );
  NAND2_X1 U8121 ( .A1(n6927), .A2(n6639), .ZN(n11972) );
  NOR2_X1 U8122 ( .A1(n11804), .A2(n7513), .ZN(n7512) );
  NAND4_X1 U8123 ( .A1(n8305), .A2(n8304), .A3(n8303), .A4(n8302), .ZN(n10299)
         );
  OR2_X1 U8124 ( .A1(n8740), .A2(n8300), .ZN(n8304) );
  OR2_X1 U8125 ( .A1(n8577), .A2(n8576), .ZN(n14546) );
  AND4_X1 U8126 ( .A1(n8538), .A2(n8537), .A3(n8536), .A4(n8535), .ZN(n14494)
         );
  OR2_X1 U8127 ( .A1(n8740), .A2(n8329), .ZN(n8332) );
  OR2_X1 U8128 ( .A1(n8364), .A2(n10915), .ZN(n8313) );
  OR2_X1 U8129 ( .A1(n8740), .A2(n8312), .ZN(n8314) );
  NAND2_X1 U8130 ( .A1(n8267), .A2(n8266), .ZN(n13996) );
  XNOR2_X1 U8131 ( .A(n6834), .B(n11935), .ZN(n14201) );
  NOR2_X1 U8132 ( .A1(n11954), .A2(n6835), .ZN(n6834) );
  AND2_X1 U8133 ( .A1(n14203), .A2(n14011), .ZN(n6835) );
  NAND2_X1 U8134 ( .A1(n8734), .A2(n8733), .ZN(n14020) );
  INV_X1 U8135 ( .A(n14252), .ZN(n14125) );
  NAND2_X1 U8136 ( .A1(n8907), .A2(n6854), .ZN(n6853) );
  NOR2_X1 U8137 ( .A1(n8908), .A2(n6856), .ZN(n6854) );
  XNOR2_X1 U8138 ( .A(n8913), .B(n8912), .ZN(n14334) );
  OR2_X1 U8139 ( .A1(n14334), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n6837) );
  INV_X1 U8140 ( .A(n6858), .ZN(n8920) );
  NAND2_X1 U8141 ( .A1(n6857), .A2(n7212), .ZN(n14625) );
  NAND2_X1 U8142 ( .A1(n14621), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7212) );
  NAND2_X1 U8143 ( .A1(n6672), .A2(n6858), .ZN(n6857) );
  NAND2_X1 U8144 ( .A1(n14629), .A2(n14630), .ZN(n14628) );
  NAND2_X1 U8145 ( .A1(n7209), .A2(n14628), .ZN(n14633) );
  OAI21_X1 U8146 ( .B1(n14629), .B2(n14630), .A(P2_ADDR_REG_15__SCAN_IN), .ZN(
        n7209) );
  NAND2_X1 U8147 ( .A1(n6847), .A2(n6846), .ZN(n7206) );
  INV_X1 U8148 ( .A(n14634), .ZN(n6846) );
  INV_X1 U8149 ( .A(n14633), .ZN(n6847) );
  MUX2_X1 U8150 ( .A(n10408), .B(n9156), .S(n9122), .Z(n8943) );
  MUX2_X1 U8151 ( .A(n13085), .B(n11082), .S(n9122), .Z(n8952) );
  NAND2_X1 U8152 ( .A1(n7125), .A2(n8984), .ZN(n7124) );
  NAND2_X1 U8153 ( .A1(n8994), .A2(n8996), .ZN(n7114) );
  NAND2_X1 U8154 ( .A1(n9005), .A2(n7117), .ZN(n7116) );
  OAI22_X1 U8155 ( .A1(n8394), .A2(n6954), .B1(n7254), .B2(n8395), .ZN(n8413)
         );
  NOR2_X1 U8156 ( .A1(n8393), .A2(n8396), .ZN(n6954) );
  NAND2_X1 U8157 ( .A1(n8413), .A2(n8414), .ZN(n8412) );
  NAND2_X1 U8158 ( .A1(n9017), .A2(n9015), .ZN(n7127) );
  NAND2_X1 U8159 ( .A1(n6971), .A2(n8455), .ZN(n6970) );
  INV_X1 U8160 ( .A(n8469), .ZN(n6971) );
  NOR2_X1 U8161 ( .A1(n8432), .A2(n8435), .ZN(n7259) );
  INV_X1 U8162 ( .A(n6962), .ZN(n6960) );
  NOR2_X1 U8163 ( .A1(n8456), .A2(n6968), .ZN(n6961) );
  OAI21_X1 U8164 ( .B1(n7241), .B2(n6964), .A(n6963), .ZN(n6962) );
  NAND2_X1 U8165 ( .A1(n6983), .A2(n6984), .ZN(n8561) );
  NOR2_X1 U8166 ( .A1(n8557), .A2(n6982), .ZN(n6981) );
  INV_X1 U8167 ( .A(n6984), .ZN(n6982) );
  NAND2_X1 U8168 ( .A1(n6981), .A2(n6986), .ZN(n6979) );
  NAND2_X1 U8169 ( .A1(n6673), .A2(n8544), .ZN(n6988) );
  NAND2_X1 U8170 ( .A1(n9052), .A2(n9054), .ZN(n7119) );
  AOI21_X1 U8171 ( .B1(n8583), .B2(n6959), .A(n6713), .ZN(n6958) );
  AND2_X1 U8172 ( .A1(n7522), .A2(n6957), .ZN(n6956) );
  NAND2_X1 U8173 ( .A1(n8582), .A2(n8584), .ZN(n6957) );
  NAND2_X1 U8174 ( .A1(n6951), .A2(n6641), .ZN(n8653) );
  NAND2_X1 U8175 ( .A1(n8626), .A2(n6952), .ZN(n6951) );
  AOI21_X1 U8176 ( .B1(n8638), .B2(n8639), .A(n6953), .ZN(n6952) );
  INV_X1 U8177 ( .A(n12449), .ZN(n7012) );
  NAND2_X1 U8178 ( .A1(n9071), .A2(n7122), .ZN(n7121) );
  INV_X1 U8179 ( .A(n7424), .ZN(n7257) );
  NAND2_X1 U8180 ( .A1(n7426), .A2(n7425), .ZN(n7424) );
  NAND2_X1 U8181 ( .A1(n13788), .A2(n8780), .ZN(n7425) );
  NAND2_X1 U8182 ( .A1(n14101), .A2(n8775), .ZN(n7426) );
  INV_X1 U8183 ( .A(n12453), .ZN(n7201) );
  NAND2_X1 U8184 ( .A1(n7008), .A2(n7322), .ZN(n7321) );
  NAND2_X1 U8185 ( .A1(n12456), .A2(n12448), .ZN(n7322) );
  NAND2_X1 U8186 ( .A1(n7009), .A2(n12473), .ZN(n7008) );
  INV_X1 U8187 ( .A(n7893), .ZN(n7433) );
  INV_X1 U8188 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7446) );
  INV_X1 U8189 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7028) );
  NAND2_X1 U8190 ( .A1(n12901), .A2(n12466), .ZN(n12469) );
  OAI21_X1 U8191 ( .B1(n9400), .B2(n7147), .A(n15232), .ZN(n7146) );
  NAND2_X1 U8192 ( .A1(n12525), .A2(n15310), .ZN(n12345) );
  AOI21_X1 U8193 ( .B1(n9582), .B2(n7318), .A(n7317), .ZN(n7316) );
  INV_X1 U8194 ( .A(n9584), .ZN(n7317) );
  INV_X1 U8195 ( .A(n9567), .ZN(n7318) );
  NAND2_X1 U8196 ( .A1(n6950), .A2(n8696), .ZN(n6949) );
  AND2_X1 U8197 ( .A1(n7253), .A2(n8724), .ZN(n7252) );
  OR2_X1 U8198 ( .A1(n11695), .A2(P1_B_REG_SCAN_IN), .ZN(n10051) );
  NAND2_X1 U8199 ( .A1(n7429), .A2(n7427), .ZN(n7938) );
  AOI21_X1 U8200 ( .B1(n7431), .B2(n7433), .A(n7428), .ZN(n7427) );
  NAND2_X1 U8201 ( .A1(n7892), .A2(n7431), .ZN(n7429) );
  INV_X1 U8202 ( .A(n7918), .ZN(n7428) );
  INV_X1 U8203 ( .A(n7873), .ZN(n7036) );
  INV_X1 U8204 ( .A(n7733), .ZN(n7048) );
  INV_X1 U8205 ( .A(n7715), .ZN(n6883) );
  OAI21_X1 U8206 ( .B1(n8893), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6663), .ZN(
        n7211) );
  INV_X1 U8207 ( .A(n12146), .ZN(n6871) );
  NAND2_X1 U8208 ( .A1(n12163), .A2(n12653), .ZN(n7493) );
  AOI21_X1 U8209 ( .B1(n12472), .B2(n12471), .A(n12448), .ZN(n7016) );
  NAND2_X1 U8210 ( .A1(n12474), .A2(n12448), .ZN(n7017) );
  AND2_X1 U8211 ( .A1(n12472), .A2(n12469), .ZN(n12474) );
  NAND2_X1 U8212 ( .A1(n10724), .A2(n6632), .ZN(n10551) );
  NAND2_X1 U8213 ( .A1(n12536), .A2(n15176), .ZN(n12537) );
  INV_X1 U8214 ( .A(n12556), .ZN(n7221) );
  OR2_X1 U8215 ( .A1(n12840), .A2(n12636), .ZN(n12449) );
  INV_X1 U8216 ( .A(n12333), .ZN(n7169) );
  NOR2_X1 U8217 ( .A1(n7170), .A2(n7166), .ZN(n7165) );
  INV_X1 U8218 ( .A(n12332), .ZN(n7166) );
  INV_X1 U8219 ( .A(n12327), .ZN(n7168) );
  OR2_X1 U8220 ( .A1(n12720), .A2(n12731), .ZN(n12333) );
  INV_X1 U8221 ( .A(n12434), .ZN(n7187) );
  INV_X1 U8222 ( .A(n9492), .ZN(n7142) );
  INV_X1 U8223 ( .A(n6608), .ZN(n7136) );
  OR2_X1 U8224 ( .A1(n9432), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9451) );
  NAND2_X1 U8225 ( .A1(n12819), .A2(n10831), .ZN(n12344) );
  NAND2_X1 U8226 ( .A1(n9226), .A2(n7153), .ZN(n7154) );
  AND2_X1 U8227 ( .A1(n7076), .A2(n10031), .ZN(n7153) );
  NAND2_X1 U8228 ( .A1(n10876), .A2(n10491), .ZN(n7133) );
  NAND2_X1 U8229 ( .A1(n9248), .A2(n12827), .ZN(n12341) );
  INV_X1 U8230 ( .A(n15256), .ZN(n15262) );
  NOR2_X1 U8231 ( .A1(n11868), .A2(n6776), .ZN(n6775) );
  INV_X1 U8232 ( .A(n9720), .ZN(n6776) );
  INV_X1 U8233 ( .A(n9717), .ZN(n6773) );
  NAND2_X1 U8234 ( .A1(n6725), .A2(n9689), .ZN(n6804) );
  AOI21_X1 U8235 ( .B1(n7334), .B2(n7336), .A(n6720), .ZN(n7332) );
  OR2_X1 U8236 ( .A1(n9643), .A2(n13595), .ZN(n9655) );
  NAND2_X1 U8237 ( .A1(n9733), .A2(n9734), .ZN(n9776) );
  INV_X1 U8238 ( .A(n6792), .ZN(n6791) );
  OAI21_X1 U8239 ( .B1(n9515), .B2(n6793), .A(n9549), .ZN(n6792) );
  INV_X1 U8240 ( .A(n9532), .ZN(n6793) );
  NOR2_X1 U8241 ( .A1(n7343), .A2(n6796), .ZN(n6794) );
  INV_X1 U8242 ( .A(n9313), .ZN(n6796) );
  NAND2_X1 U8243 ( .A1(n7345), .A2(n7344), .ZN(n7343) );
  INV_X1 U8244 ( .A(n9367), .ZN(n7344) );
  NOR2_X1 U8245 ( .A1(n7346), .A2(n9367), .ZN(n7342) );
  OR2_X1 U8246 ( .A1(n9370), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9395) );
  NAND2_X1 U8247 ( .A1(n13083), .A2(n9935), .ZN(n9879) );
  NAND2_X1 U8248 ( .A1(n9091), .A2(n9089), .ZN(n7129) );
  AOI21_X1 U8249 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n15027), .A(n15021), .ZN(
        n13135) );
  NOR2_X1 U8250 ( .A1(n7104), .A2(n7099), .ZN(n7098) );
  OR2_X1 U8251 ( .A1(n7421), .A2(n7420), .ZN(n7418) );
  INV_X1 U8252 ( .A(n8183), .ZN(n7420) );
  NOR2_X1 U8253 ( .A1(n13295), .A2(n13409), .ZN(n7089) );
  NOR2_X1 U8254 ( .A1(n7865), .A2(n7864), .ZN(n7907) );
  NOR2_X1 U8255 ( .A1(n14482), .A2(n11551), .ZN(n7095) );
  AND2_X1 U8256 ( .A1(n11353), .A2(n15093), .ZN(n11352) );
  AND2_X1 U8257 ( .A1(n7409), .A2(n11213), .ZN(n7408) );
  OR2_X1 U8258 ( .A1(n11045), .A2(n7410), .ZN(n7409) );
  INV_X1 U8259 ( .A(n8164), .ZN(n7410) );
  NAND2_X1 U8260 ( .A1(n7584), .A2(n7574), .ZN(n7405) );
  INV_X1 U8261 ( .A(n11076), .ZN(n11072) );
  XNOR2_X1 U8262 ( .A(n8231), .B(n8230), .ZN(n10165) );
  INV_X1 U8263 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8210) );
  INV_X1 U8264 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7540) );
  OR2_X1 U8265 ( .A1(n7716), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n7734) );
  NAND2_X1 U8266 ( .A1(n6936), .A2(n6938), .ZN(n6934) );
  INV_X1 U8267 ( .A(n12034), .ZN(n10265) );
  AND2_X1 U8268 ( .A1(n7392), .A2(n14023), .ZN(n7391) );
  OR2_X1 U8269 ( .A1(n7394), .A2(n7393), .ZN(n7392) );
  NOR2_X1 U8270 ( .A1(n14068), .A2(n7002), .ZN(n7001) );
  INV_X1 U8271 ( .A(n7003), .ZN(n7002) );
  NOR2_X1 U8272 ( .A1(n14235), .A2(n7004), .ZN(n7003) );
  NOR2_X1 U8273 ( .A1(n14592), .A2(n14184), .ZN(n6991) );
  NAND2_X1 U8274 ( .A1(n6809), .A2(n11329), .ZN(n14699) );
  NOR2_X1 U8275 ( .A1(n14811), .A2(n13893), .ZN(n7277) );
  NAND2_X1 U8276 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n7310) );
  NOR2_X1 U8277 ( .A1(n14214), .A2(n14043), .ZN(n14035) );
  INV_X1 U8278 ( .A(n11261), .ZN(n10789) );
  AOI21_X1 U8279 ( .B1(n10273), .B2(n10272), .A(n10271), .ZN(n11567) );
  INV_X1 U8280 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7398) );
  NAND2_X1 U8281 ( .A1(n8121), .A2(n8120), .ZN(n8242) );
  NAND2_X1 U8282 ( .A1(n8093), .A2(n8092), .ZN(n8119) );
  NAND2_X1 U8283 ( .A1(n7436), .A2(n6710), .ZN(n7051) );
  INV_X1 U8284 ( .A(SI_22_), .ZN(n7435) );
  INV_X1 U8285 ( .A(n6942), .ZN(n6940) );
  INV_X1 U8286 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8269) );
  XNOR2_X1 U8287 ( .A(n7938), .B(SI_18_), .ZN(n7937) );
  NAND4_X1 U8288 ( .A1(n8258), .A2(n6989), .A3(n8352), .A4(n8257), .ZN(n8578)
         );
  AND2_X1 U8289 ( .A1(n7893), .A2(n7879), .ZN(n7891) );
  INV_X1 U8290 ( .A(n7832), .ZN(n7040) );
  NOR2_X1 U8291 ( .A1(n7833), .A2(n7043), .ZN(n7042) );
  NOR2_X1 U8292 ( .A1(n7794), .A2(n6895), .ZN(n6894) );
  INV_X1 U8293 ( .A(n7773), .ZN(n6895) );
  OR2_X1 U8294 ( .A1(n8389), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n8405) );
  NAND2_X1 U8295 ( .A1(n7620), .A2(n7619), .ZN(n7627) );
  INV_X1 U8296 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8840) );
  INV_X1 U8297 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n8843) );
  XNOR2_X1 U8298 ( .A(n7211), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n8881) );
  INV_X1 U8299 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n13653) );
  INV_X1 U8300 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n8875) );
  OR2_X1 U8301 ( .A1(n14618), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n6840) );
  AOI21_X1 U8302 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n8862), .A(n8861), .ZN(
        n8917) );
  INV_X1 U8303 ( .A(n11360), .ZN(n10790) );
  AOI21_X1 U8304 ( .B1(n7470), .B2(n7469), .A(n6629), .ZN(n7468) );
  INV_X1 U8305 ( .A(n11811), .ZN(n7469) );
  NAND2_X1 U8306 ( .A1(n6860), .A2(n7470), .ZN(n7467) );
  CLKBUF_X1 U8307 ( .A(n9248), .Z(n10827) );
  NAND2_X1 U8308 ( .A1(n9607), .A2(n9606), .ZN(n9619) );
  INV_X1 U8309 ( .A(n12318), .ZN(n9603) );
  AND3_X1 U8310 ( .A1(n9322), .A2(n9321), .A3(n9320), .ZN(n11000) );
  AND2_X1 U8311 ( .A1(n9590), .A2(n12258), .ZN(n9607) );
  NAND2_X1 U8312 ( .A1(n6862), .A2(n6861), .ZN(n11725) );
  INV_X1 U8313 ( .A(n11709), .ZN(n6861) );
  XNOR2_X1 U8314 ( .A(n10831), .B(n10834), .ZN(n10832) );
  OR2_X1 U8315 ( .A1(n9556), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9576) );
  NAND2_X1 U8316 ( .A1(n9543), .A2(n12235), .ZN(n9556) );
  NAND2_X1 U8317 ( .A1(n7483), .A2(n7482), .ZN(n7494) );
  INV_X1 U8318 ( .A(n12162), .ZN(n7482) );
  XNOR2_X1 U8319 ( .A(n6798), .B(n10513), .ZN(n12322) );
  NAND2_X1 U8320 ( .A1(n6591), .A2(n7203), .ZN(n7193) );
  NAND2_X1 U8321 ( .A1(n7194), .A2(n7197), .ZN(n6799) );
  NAND2_X1 U8322 ( .A1(n7014), .A2(n7013), .ZN(n12478) );
  NAND2_X1 U8323 ( .A1(n7195), .A2(n12513), .ZN(n7013) );
  NAND2_X1 U8324 ( .A1(n7017), .A2(n7015), .ZN(n7014) );
  NOR2_X1 U8325 ( .A1(n7016), .A2(n12475), .ZN(n7015) );
  NAND2_X1 U8326 ( .A1(n12478), .A2(n12477), .ZN(n12506) );
  OR2_X1 U8327 ( .A1(n12504), .A2(n10817), .ZN(n12505) );
  INV_X1 U8328 ( .A(n9304), .ZN(n9741) );
  AND4_X1 U8329 ( .A1(n9508), .A2(n9507), .A3(n9506), .A4(n9505), .ZN(n12175)
         );
  AND4_X1 U8330 ( .A1(n9385), .A2(n9384), .A3(n9383), .A4(n9382), .ZN(n15233)
         );
  OAI21_X1 U8331 ( .B1(n12589), .B2(n10635), .A(n6733), .ZN(n10417) );
  NAND2_X1 U8332 ( .A1(n12589), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n6733) );
  XNOR2_X1 U8333 ( .A(n10547), .B(n6765), .ZN(n10439) );
  NAND2_X1 U8334 ( .A1(n10439), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10548) );
  NAND2_X1 U8335 ( .A1(n14321), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7236) );
  XNOR2_X1 U8336 ( .A(n10551), .B(n10552), .ZN(n10741) );
  NOR2_X1 U8337 ( .A1(n12531), .A2(n9361), .ZN(n7238) );
  INV_X1 U8338 ( .A(n12544), .ZN(n7239) );
  XNOR2_X1 U8339 ( .A(n12532), .B(n12568), .ZN(n15129) );
  NAND2_X1 U8340 ( .A1(n15129), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n15128) );
  XNOR2_X1 U8341 ( .A(n12534), .B(n12574), .ZN(n15160) );
  NAND2_X1 U8342 ( .A1(n15160), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n15159) );
  NAND2_X1 U8343 ( .A1(n15166), .A2(n12576), .ZN(n15185) );
  NAND2_X1 U8344 ( .A1(n7231), .A2(n12583), .ZN(n7229) );
  INV_X1 U8345 ( .A(n6609), .ZN(n7231) );
  OR2_X1 U8346 ( .A1(n15210), .A2(n15194), .ZN(n7230) );
  OR2_X1 U8347 ( .A1(n15193), .A2(n15194), .ZN(n7232) );
  OR2_X1 U8348 ( .A1(n14387), .A2(n12559), .ZN(n7227) );
  NAND2_X1 U8349 ( .A1(n7227), .A2(n7226), .ZN(n7225) );
  INV_X1 U8350 ( .A(n14413), .ZN(n7226) );
  NAND2_X1 U8351 ( .A1(n9770), .A2(n12497), .ZN(n9836) );
  OR2_X1 U8352 ( .A1(n9676), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9693) );
  NAND2_X1 U8353 ( .A1(n9685), .A2(n9684), .ZN(n12633) );
  AND2_X1 U8354 ( .A1(n9703), .A2(n9684), .ZN(n7143) );
  NOR2_X1 U8355 ( .A1(n9647), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9660) );
  OR2_X1 U8356 ( .A1(n9619), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9632) );
  NAND2_X1 U8357 ( .A1(n12726), .A2(n9614), .ZN(n12715) );
  NAND2_X1 U8358 ( .A1(n9767), .A2(n12335), .ZN(n12719) );
  OAI21_X1 U8359 ( .B1(n9766), .B2(n7189), .A(n7186), .ZN(n12733) );
  INV_X1 U8360 ( .A(n7190), .ZN(n7189) );
  AOI21_X1 U8361 ( .B1(n7190), .B2(n7188), .A(n7187), .ZN(n7186) );
  INV_X1 U8362 ( .A(n12429), .ZN(n7188) );
  NOR2_X1 U8363 ( .A1(n7175), .A2(n7173), .ZN(n7172) );
  INV_X1 U8364 ( .A(n12400), .ZN(n7173) );
  NAND2_X1 U8365 ( .A1(n11664), .A2(n12490), .ZN(n11663) );
  INV_X1 U8366 ( .A(n7181), .ZN(n7180) );
  AOI21_X1 U8367 ( .B1(n7181), .B2(n7179), .A(n7178), .ZN(n7177) );
  AND4_X1 U8368 ( .A1(n9408), .A2(n9407), .A3(n9406), .A4(n9405), .ZN(n14425)
         );
  AND2_X1 U8369 ( .A1(n12380), .A2(n12381), .ZN(n12482) );
  NAND2_X1 U8370 ( .A1(n11475), .A2(n9400), .ZN(n11474) );
  INV_X1 U8371 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10681) );
  INV_X1 U8372 ( .A(n15246), .ZN(n15242) );
  NOR2_X1 U8373 ( .A1(n9341), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9358) );
  OR2_X1 U8374 ( .A1(n9325), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9341) );
  AND2_X1 U8375 ( .A1(n12356), .A2(n15290), .ZN(n9751) );
  AND3_X1 U8376 ( .A1(n9298), .A2(n9297), .A3(n9296), .ZN(n15302) );
  NAND2_X1 U8377 ( .A1(n15315), .A2(n6613), .ZN(n10923) );
  NAND2_X1 U8378 ( .A1(n15315), .A2(n9260), .ZN(n10921) );
  NAND2_X1 U8379 ( .A1(n9775), .A2(n9813), .ZN(n15297) );
  INV_X1 U8380 ( .A(n9750), .ZN(n12480) );
  INV_X1 U8381 ( .A(n10831), .ZN(n15310) );
  OR2_X1 U8382 ( .A1(n10654), .A2(n10514), .ZN(n12508) );
  NOR2_X1 U8383 ( .A1(n9827), .A2(n9826), .ZN(n10488) );
  INV_X1 U8384 ( .A(n15368), .ZN(n15301) );
  INV_X1 U8385 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7472) );
  INV_X1 U8386 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9217) );
  INV_X1 U8387 ( .A(n6734), .ZN(n9221) );
  NAND2_X1 U8388 ( .A1(n9221), .A2(n9217), .ZN(n9230) );
  AND2_X1 U8389 ( .A1(n9783), .A2(n6626), .ZN(n9790) );
  NOR2_X1 U8390 ( .A1(n9629), .A2(n7338), .ZN(n7337) );
  INV_X1 U8391 ( .A(n9615), .ZN(n7338) );
  XNOR2_X1 U8392 ( .A(n9778), .B(n9777), .ZN(n10422) );
  INV_X1 U8393 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9777) );
  OAI21_X1 U8394 ( .B1(n9776), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9778) );
  XNOR2_X1 U8395 ( .A(n9737), .B(P3_IR_REG_20__SCAN_IN), .ZN(n9820) );
  AND2_X1 U8396 ( .A1(n9518), .A2(n9535), .ZN(n6873) );
  AND2_X1 U8397 ( .A1(n9482), .A2(n9518), .ZN(n9536) );
  AND2_X1 U8398 ( .A1(n9458), .A2(n9442), .ZN(n9443) );
  NAND2_X1 U8399 ( .A1(n9444), .A2(n9443), .ZN(n9459) );
  AOI21_X1 U8400 ( .B1(n7327), .B2(n7330), .A(n7326), .ZN(n7325) );
  AND2_X1 U8401 ( .A1(n9440), .A2(n9423), .ZN(n9424) );
  OR2_X1 U8402 ( .A1(n9351), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n9370) );
  NAND2_X1 U8403 ( .A1(n9254), .A2(n9209), .ZN(n9315) );
  NAND2_X1 U8404 ( .A1(n6770), .A2(n9270), .ZN(n9290) );
  XNOR2_X1 U8405 ( .A(n10006), .B(P1_DATAO_REG_2__SCAN_IN), .ZN(n9267) );
  NAND2_X1 U8406 ( .A1(n9253), .A2(n6771), .ZN(n9269) );
  NAND2_X1 U8407 ( .A1(n10233), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6771) );
  NOR2_X1 U8408 ( .A1(n7005), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9224) );
  XNOR2_X1 U8409 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9225) );
  NAND2_X1 U8410 ( .A1(n6748), .A2(n9231), .ZN(n6747) );
  INV_X1 U8411 ( .A(n7368), .ZN(n7367) );
  OAI21_X1 U8412 ( .B1(n7370), .B2(n13000), .A(n12109), .ZN(n7368) );
  NAND2_X1 U8413 ( .A1(n6615), .A2(n7359), .ZN(n7358) );
  INV_X1 U8414 ( .A(n11845), .ZN(n7359) );
  NAND2_X1 U8415 ( .A1(n7360), .A2(n6615), .ZN(n7357) );
  NAND2_X1 U8416 ( .A1(n13041), .A2(n9951), .ZN(n7360) );
  INV_X1 U8417 ( .A(n6580), .ZN(n12116) );
  XNOR2_X1 U8418 ( .A(n6579), .B(n10595), .ZN(n9860) );
  NOR2_X1 U8419 ( .A1(n11822), .A2(n9948), .ZN(n11843) );
  NAND2_X1 U8420 ( .A1(n6896), .A2(n7355), .ZN(n12983) );
  AND2_X1 U8421 ( .A1(n7356), .A2(n12984), .ZN(n7355) );
  NAND2_X1 U8422 ( .A1(n11843), .A2(n7357), .ZN(n6896) );
  NAND2_X1 U8423 ( .A1(n7357), .A2(n7358), .ZN(n7356) );
  NAND2_X1 U8424 ( .A1(n11380), .A2(n11381), .ZN(n11379) );
  NOR2_X1 U8425 ( .A1(n8000), .A2(n9978), .ZN(n8013) );
  INV_X1 U8426 ( .A(n9911), .ZN(n7366) );
  NAND2_X1 U8427 ( .A1(n13052), .A2(n7371), .ZN(n7370) );
  INV_X1 U8428 ( .A(n12105), .ZN(n7371) );
  INV_X1 U8429 ( .A(n9140), .ZN(n9110) );
  NAND2_X1 U8430 ( .A1(n11192), .A2(n11262), .ZN(n9193) );
  AND2_X1 U8431 ( .A1(n9149), .A2(n9148), .ZN(n9191) );
  AND4_X1 U8432 ( .A1(n8113), .A2(n8112), .A3(n8111), .A4(n8110), .ZN(n12969)
         );
  AND4_X1 U8433 ( .A1(n8090), .A2(n8089), .A3(n8088), .A4(n8087), .ZN(n13053)
         );
  CLKBUF_X1 U8434 ( .A(n7682), .Z(n9101) );
  AOI21_X1 U8436 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n14964), .A(n14957), .ZN(
        n10357) );
  AOI21_X1 U8437 ( .B1(n7065), .B2(n7067), .A(n6633), .ZN(n7063) );
  NAND2_X1 U8438 ( .A1(n13256), .A2(n13397), .ZN(n13247) );
  AND2_X1 U8439 ( .A1(n13305), .A2(n7087), .ZN(n13256) );
  AND2_X1 U8440 ( .A1(n7088), .A2(n7089), .ZN(n7087) );
  OAI21_X1 U8441 ( .B1(n8182), .B2(n7419), .A(n7416), .ZN(n13281) );
  INV_X1 U8442 ( .A(n7417), .ZN(n7416) );
  OR2_X1 U8443 ( .A1(n13290), .A2(n7420), .ZN(n7419) );
  OAI21_X1 U8444 ( .B1(n13290), .B2(n7418), .A(n8185), .ZN(n7417) );
  NAND2_X1 U8445 ( .A1(n13305), .A2(n13469), .ZN(n13292) );
  NAND2_X1 U8446 ( .A1(n13305), .A2(n7089), .ZN(n13274) );
  AOI21_X1 U8447 ( .B1(n7058), .B2(n7061), .A(n6628), .ZN(n7055) );
  INV_X1 U8448 ( .A(n7957), .ZN(n7061) );
  NOR2_X1 U8449 ( .A1(n13429), .A2(n7091), .ZN(n7090) );
  INV_X1 U8450 ( .A(n7092), .ZN(n7091) );
  OAI21_X1 U8451 ( .B1(n13362), .B2(n9038), .A(n9155), .ZN(n13328) );
  NAND2_X1 U8452 ( .A1(n11769), .A2(n7092), .ZN(n13353) );
  NAND2_X1 U8453 ( .A1(n11769), .A2(n13445), .ZN(n13355) );
  NAND2_X1 U8454 ( .A1(n7094), .A2(n14472), .ZN(n14464) );
  OR2_X1 U8455 ( .A1(n7843), .A2(n7842), .ZN(n7865) );
  NOR2_X1 U8456 ( .A1(n7070), .A2(n7069), .ZN(n7068) );
  NOR2_X1 U8457 ( .A1(n14477), .A2(n13074), .ZN(n7069) );
  NOR2_X1 U8458 ( .A1(n7072), .A2(n7071), .ZN(n7070) );
  INV_X1 U8459 ( .A(n7402), .ZN(n7400) );
  NAND2_X1 U8460 ( .A1(n11352), .A2(n7095), .ZN(n11559) );
  NAND2_X1 U8461 ( .A1(n6743), .A2(n7793), .ZN(n11460) );
  NAND2_X1 U8462 ( .A1(n11352), .A2(n11548), .ZN(n11491) );
  OR2_X1 U8463 ( .A1(n7743), .A2(n13748), .ZN(n7760) );
  NAND2_X1 U8464 ( .A1(n6754), .A2(n6753), .ZN(n11210) );
  INV_X1 U8465 ( .A(n11213), .ZN(n6753) );
  NOR2_X1 U8466 ( .A1(n11216), .A2(n11339), .ZN(n11353) );
  OR2_X1 U8467 ( .A1(n11053), .A2(n11052), .ZN(n11216) );
  NAND2_X1 U8468 ( .A1(n10986), .A2(n10990), .ZN(n11053) );
  NOR2_X1 U8469 ( .A1(n10899), .A2(n10869), .ZN(n10986) );
  NAND2_X1 U8470 ( .A1(n7086), .A2(n7085), .ZN(n10899) );
  AND2_X1 U8471 ( .A1(n10166), .A2(n8146), .ZN(n13335) );
  NAND2_X1 U8472 ( .A1(n11075), .A2(n11076), .ZN(n11074) );
  NOR2_X1 U8473 ( .A1(n8155), .A2(n11012), .ZN(n9992) );
  OR2_X1 U8474 ( .A1(n10308), .A2(n9179), .ZN(n9973) );
  CLKBUF_X1 U8475 ( .A(n9857), .Z(n8198) );
  INV_X1 U8476 ( .A(n9856), .ZN(n9989) );
  AOI21_X1 U8477 ( .B1(n13184), .B2(n7539), .A(n13183), .ZN(n13379) );
  OR2_X1 U8478 ( .A1(n13188), .A2(n13187), .ZN(n13378) );
  OR2_X1 U8479 ( .A1(n13199), .A2(n13198), .ZN(n13383) );
  NAND2_X1 U8480 ( .A1(n7084), .A2(n8008), .ZN(n13260) );
  AND2_X1 U8481 ( .A1(n8232), .A2(n10165), .ZN(n9975) );
  OR2_X1 U8482 ( .A1(n9853), .A2(n9851), .ZN(n8232) );
  CLKBUF_X1 U8483 ( .A(n8144), .Z(n8145) );
  NAND2_X1 U8484 ( .A1(n7568), .A2(n7565), .ZN(n13484) );
  MUX2_X1 U8485 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7567), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n7568) );
  INV_X1 U8486 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7444) );
  XNOR2_X1 U8487 ( .A(n8211), .B(n8210), .ZN(n9851) );
  OAI21_X1 U8488 ( .B1(n8208), .B2(n8209), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8211) );
  BUF_X1 U8489 ( .A(n8141), .Z(n8209) );
  OR2_X1 U8490 ( .A1(n7818), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n7858) );
  OR2_X1 U8491 ( .A1(n7734), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n7736) );
  AND2_X1 U8492 ( .A1(n6619), .A2(n11644), .ZN(n6932) );
  NOR2_X1 U8493 ( .A1(n13795), .A2(n7510), .ZN(n7509) );
  INV_X1 U8494 ( .A(n12016), .ZN(n7510) );
  NOR2_X1 U8495 ( .A1(n8627), .A2(n13834), .ZN(n8641) );
  INV_X1 U8496 ( .A(n11797), .ZN(n7513) );
  NAND2_X1 U8497 ( .A1(n6928), .A2(n6931), .ZN(n6926) );
  OR2_X1 U8498 ( .A1(n8573), .A2(n8572), .ZN(n8597) );
  AOI21_X1 U8499 ( .B1(n8319), .B2(n12079), .A(n10262), .ZN(n10263) );
  AND2_X1 U8500 ( .A1(n10261), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10262) );
  INV_X1 U8501 ( .A(n12024), .ZN(n6938) );
  INV_X1 U8502 ( .A(n6937), .ZN(n6936) );
  OAI21_X1 U8503 ( .B1(n7509), .B2(n6938), .A(n13830), .ZN(n6937) );
  OR2_X1 U8504 ( .A1(n8506), .A2(n10368), .ZN(n8532) );
  NAND2_X1 U8505 ( .A1(n8659), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U8506 ( .A1(n13851), .A2(n13852), .ZN(n13850) );
  AND2_X1 U8507 ( .A1(n8471), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8485) );
  NAND2_X1 U8508 ( .A1(n10064), .A2(n6599), .ZN(n6811) );
  NOR2_X1 U8509 ( .A1(n8597), .A2(n13944), .ZN(n8598) );
  NAND2_X1 U8510 ( .A1(n6905), .A2(n6904), .ZN(n13870) );
  INV_X1 U8511 ( .A(n11392), .ZN(n6906) );
  AND2_X1 U8512 ( .A1(n7244), .A2(n6975), .ZN(n6974) );
  NAND2_X1 U8513 ( .A1(n8747), .A2(n8749), .ZN(n6975) );
  NAND2_X1 U8514 ( .A1(n7247), .A2(n8760), .ZN(n7246) );
  AND4_X1 U8515 ( .A1(n8531), .A2(n8530), .A3(n8529), .A4(n8528), .ZN(n14556)
         );
  OR2_X1 U8516 ( .A1(n8512), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8513) );
  NAND2_X1 U8517 ( .A1(n14108), .A2(n6999), .ZN(n14043) );
  AND2_X1 U8518 ( .A1(n7001), .A2(n7000), .ZN(n6999) );
  NAND2_X1 U8519 ( .A1(n14108), .A2(n7001), .ZN(n14065) );
  NAND2_X1 U8520 ( .A1(n14108), .A2(n14101), .ZN(n14093) );
  OAI21_X1 U8521 ( .B1(n14153), .B2(n7384), .A(n7381), .ZN(n14114) );
  AOI21_X1 U8522 ( .B1(n14118), .B2(n7380), .A(n6659), .ZN(n7381) );
  AND2_X1 U8523 ( .A1(n7386), .A2(n7382), .ZN(n7380) );
  INV_X1 U8524 ( .A(n14095), .ZN(n14108) );
  INV_X1 U8525 ( .A(n7303), .ZN(n7302) );
  OAI22_X1 U8526 ( .A1(n7306), .A2(n7304), .B1(n14125), .B2(n13799), .ZN(n7303) );
  NAND2_X1 U8527 ( .A1(n7305), .A2(n11922), .ZN(n7304) );
  NAND2_X1 U8528 ( .A1(n14564), .A2(n6991), .ZN(n14176) );
  NAND2_X1 U8529 ( .A1(n6824), .A2(n6825), .ZN(n14175) );
  AOI21_X1 U8530 ( .B1(n11687), .B2(n6826), .A(n6601), .ZN(n6825) );
  NAND2_X1 U8531 ( .A1(n14175), .A2(n14174), .ZN(n14173) );
  AND2_X1 U8532 ( .A1(n14564), .A2(n14561), .ZN(n14565) );
  NOR2_X1 U8533 ( .A1(n8534), .A2(n8525), .ZN(n8549) );
  OR2_X1 U8534 ( .A1(n8532), .A2(n13746), .ZN(n8534) );
  NOR2_X1 U8535 ( .A1(n6995), .A2(n11799), .ZN(n6994) );
  INV_X1 U8536 ( .A(n14708), .ZN(n6993) );
  NAND2_X1 U8537 ( .A1(n6992), .A2(n11973), .ZN(n11679) );
  NAND2_X1 U8538 ( .A1(n7278), .A2(n7279), .ZN(n11676) );
  AOI21_X1 U8539 ( .B1(n7280), .B2(n7282), .A(n11536), .ZN(n7278) );
  OAI21_X1 U8540 ( .B1(n11410), .B2(n7282), .A(n7280), .ZN(n11528) );
  OR2_X1 U8541 ( .A1(n14707), .A2(n14705), .ZN(n14708) );
  NOR2_X1 U8542 ( .A1(n14708), .A2(n14834), .ZN(n11417) );
  NOR2_X1 U8543 ( .A1(n8457), .A2(n13580), .ZN(n8471) );
  INV_X1 U8544 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n13580) );
  AOI21_X1 U8545 ( .B1(n7272), .B2(n7274), .A(n7269), .ZN(n7268) );
  INV_X1 U8546 ( .A(n7275), .ZN(n7274) );
  NAND2_X1 U8547 ( .A1(n7271), .A2(n7275), .ZN(n11314) );
  NAND2_X1 U8548 ( .A1(n11271), .A2(n7276), .ZN(n7271) );
  INV_X1 U8549 ( .A(n7277), .ZN(n7276) );
  NAND2_X1 U8550 ( .A1(n8431), .A2(n8430), .ZN(n11390) );
  NOR2_X1 U8551 ( .A1(n11266), .A2(n11390), .ZN(n11265) );
  OR2_X1 U8552 ( .A1(n14724), .A2(n13872), .ZN(n11266) );
  NAND2_X1 U8553 ( .A1(n11109), .A2(n11108), .ZN(n7376) );
  NAND2_X1 U8554 ( .A1(n7301), .A2(n11095), .ZN(n11118) );
  NAND2_X1 U8555 ( .A1(n6723), .A2(n14796), .ZN(n14724) );
  INV_X1 U8556 ( .A(n14745), .ZN(n14725) );
  NAND2_X1 U8557 ( .A1(n10787), .A2(n10786), .ZN(n11104) );
  INV_X1 U8558 ( .A(n14555), .ZN(n14178) );
  NOR2_X1 U8559 ( .A1(n14746), .A2(n14782), .ZN(n14744) );
  OR2_X1 U8560 ( .A1(n10938), .A2(n10937), .ZN(n14734) );
  INV_X1 U8561 ( .A(n10936), .ZN(n10941) );
  INV_X1 U8562 ( .A(n8320), .ZN(n10266) );
  INV_X1 U8563 ( .A(n13996), .ZN(n14191) );
  INV_X1 U8564 ( .A(n14020), .ZN(n11907) );
  NAND2_X1 U8565 ( .A1(n11889), .A2(n11888), .ZN(n14568) );
  INV_X1 U8566 ( .A(n14833), .ZN(n14824) );
  AND2_X1 U8567 ( .A1(n14734), .A2(n14786), .ZN(n14793) );
  AND2_X1 U8568 ( .A1(n8765), .A2(n8764), .ZN(n11874) );
  NAND2_X1 U8569 ( .A1(n7052), .A2(n7051), .ZN(n8656) );
  NAND2_X1 U8570 ( .A1(n8270), .A2(n8269), .ZN(n8282) );
  AND2_X1 U8571 ( .A1(n8541), .A2(n8540), .ZN(n10688) );
  AOI21_X1 U8572 ( .B1(n6891), .B2(n6893), .A(n7043), .ZN(n6889) );
  NAND2_X1 U8573 ( .A1(n7045), .A2(n7733), .ZN(n7752) );
  NAND2_X1 U8574 ( .A1(n7731), .A2(n7730), .ZN(n7045) );
  OR2_X1 U8575 ( .A1(n8436), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8438) );
  XNOR2_X1 U8576 ( .A(n7713), .B(n7711), .ZN(n10057) );
  NAND2_X1 U8577 ( .A1(n6886), .A2(n7656), .ZN(n7667) );
  OR2_X1 U8578 ( .A1(n10005), .A2(n6688), .ZN(n8317) );
  INV_X1 U8579 ( .A(n8887), .ZN(n8886) );
  AND2_X1 U8580 ( .A1(n6844), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6841) );
  INV_X1 U8581 ( .A(n8885), .ZN(n6843) );
  XNOR2_X1 U8582 ( .A(n8844), .B(n8843), .ZN(n8893) );
  XNOR2_X1 U8583 ( .A(n8881), .B(n7210), .ZN(n8882) );
  INV_X1 U8584 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7210) );
  INV_X1 U8585 ( .A(n6845), .ZN(n8900) );
  INV_X1 U8586 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n13648) );
  NOR2_X1 U8587 ( .A1(n8851), .A2(n8850), .ZN(n8901) );
  OR2_X1 U8588 ( .A1(n14621), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7213) );
  OAI21_X1 U8589 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n8868), .A(n8867), .ZN(
        n8925) );
  AOI21_X1 U8590 ( .B1(n12156), .B2(n7480), .A(n7485), .ZN(n7478) );
  NAND2_X1 U8591 ( .A1(n12263), .A2(n7479), .ZN(n7477) );
  OAI22_X1 U8592 ( .A1(n7486), .A2(n12278), .B1(n12670), .B2(n12165), .ZN(
        n7485) );
  NAND2_X1 U8593 ( .A1(n7467), .A2(n7468), .ZN(n12173) );
  NAND2_X1 U8594 ( .A1(n11448), .A2(n11445), .ZN(n11708) );
  NAND2_X1 U8595 ( .A1(n7456), .A2(n11305), .ZN(n11424) );
  NAND2_X1 U8596 ( .A1(n11303), .A2(n11302), .ZN(n7456) );
  AND2_X1 U8597 ( .A1(n10828), .A2(n10830), .ZN(n7449) );
  NAND2_X1 U8598 ( .A1(n10834), .A2(n6755), .ZN(n10828) );
  NOR2_X1 U8599 ( .A1(n10827), .A2(n10876), .ZN(n6755) );
  AOI21_X1 U8600 ( .B1(n6869), .B2(n6872), .A(n6868), .ZN(n6867) );
  INV_X1 U8601 ( .A(n12211), .ZN(n6868) );
  OAI21_X1 U8602 ( .B1(n12190), .B2(n6872), .A(n6869), .ZN(n12212) );
  NAND2_X1 U8603 ( .A1(n7450), .A2(n7451), .ZN(n12224) );
  AND2_X1 U8604 ( .A1(n12225), .A2(n7452), .ZN(n7451) );
  NAND2_X1 U8605 ( .A1(n12287), .A2(n12135), .ZN(n7450) );
  NAND2_X1 U8606 ( .A1(n12286), .A2(n12135), .ZN(n7452) );
  INV_X1 U8607 ( .A(n12522), .ZN(n15259) );
  NAND2_X1 U8608 ( .A1(n7455), .A2(n7454), .ZN(n11429) );
  AOI21_X1 U8609 ( .B1(n7457), .B2(n7459), .A(n6627), .ZN(n7454) );
  NAND2_X1 U8610 ( .A1(n12256), .A2(n12255), .ZN(n12254) );
  NAND2_X1 U8611 ( .A1(n12190), .A2(n12146), .ZN(n12256) );
  AND4_X1 U8612 ( .A1(n9456), .A2(n9455), .A3(n9454), .A4(n9453), .ZN(n14426)
         );
  INV_X1 U8613 ( .A(n12285), .ZN(n12269) );
  NAND2_X1 U8614 ( .A1(n11139), .A2(n6643), .ZN(n11201) );
  NAND2_X1 U8615 ( .A1(n11139), .A2(n11138), .ZN(n11140) );
  OR3_X1 U8616 ( .A1(n10493), .A2(n15368), .A3(n10654), .ZN(n12298) );
  NAND2_X1 U8617 ( .A1(n7453), .A2(n12133), .ZN(n12288) );
  INV_X1 U8618 ( .A(n12287), .ZN(n7453) );
  INV_X1 U8619 ( .A(n12512), .ZN(n7314) );
  AND2_X1 U8620 ( .A1(n12310), .A2(n9728), .ZN(n12205) );
  INV_X1 U8621 ( .A(n12654), .ZN(n12514) );
  NAND2_X1 U8622 ( .A1(n9639), .A2(n9638), .ZN(n12687) );
  INV_X1 U8623 ( .A(n12742), .ZN(n12515) );
  INV_X1 U8624 ( .A(n12741), .ZN(n12763) );
  INV_X1 U8625 ( .A(n12807), .ZN(n12516) );
  INV_X1 U8626 ( .A(n14426), .ZN(n12519) );
  INV_X1 U8627 ( .A(n14425), .ZN(n12521) );
  INV_X1 U8628 ( .A(n10841), .ZN(n12524) );
  INV_X1 U8629 ( .A(n12819), .ZN(n12525) );
  OR2_X2 U8630 ( .A1(n12951), .A2(n10481), .ZN(n12526) );
  INV_X1 U8631 ( .A(n7234), .ZN(n10544) );
  INV_X1 U8632 ( .A(n7240), .ZN(n12545) );
  NOR2_X1 U8633 ( .A1(n9381), .A2(n15118), .ZN(n15117) );
  INV_X1 U8634 ( .A(n6741), .ZN(n12550) );
  OR2_X1 U8635 ( .A1(n15185), .A2(n15186), .ZN(n15187) );
  NAND2_X1 U8636 ( .A1(n7228), .A2(n7229), .ZN(n15209) );
  AND2_X1 U8637 ( .A1(n15202), .A2(n12582), .ZN(n15225) );
  NOR2_X1 U8638 ( .A1(n14350), .A2(n12556), .ZN(n14368) );
  XNOR2_X1 U8639 ( .A(n12558), .B(n12594), .ZN(n14388) );
  INV_X1 U8640 ( .A(n7227), .ZN(n14414) );
  INV_X1 U8641 ( .A(n15108), .ZN(n15220) );
  OAI21_X1 U8642 ( .B1(n9748), .B2(n15299), .A(n9747), .ZN(n12617) );
  AND2_X1 U8643 ( .A1(n12672), .A2(n12671), .ZN(n12848) );
  NOR2_X1 U8644 ( .A1(n12684), .A2(n12683), .ZN(n12850) );
  NAND2_X1 U8645 ( .A1(n9646), .A2(n9645), .ZN(n12849) );
  NAND2_X1 U8646 ( .A1(n9596), .A2(n9595), .ZN(n12728) );
  NAND2_X1 U8647 ( .A1(n7192), .A2(n12430), .ZN(n12743) );
  NAND2_X1 U8648 ( .A1(n9766), .A2(n12429), .ZN(n7192) );
  NAND2_X1 U8649 ( .A1(n12761), .A2(n7156), .ZN(n12750) );
  NAND2_X1 U8650 ( .A1(n11739), .A2(n9492), .ZN(n12804) );
  NAND2_X1 U8651 ( .A1(n7174), .A2(n12400), .ZN(n11743) );
  NAND2_X1 U8652 ( .A1(n11619), .A2(n9457), .ZN(n11620) );
  NAND2_X1 U8653 ( .A1(n7176), .A2(n7181), .ZN(n14420) );
  NAND2_X1 U8654 ( .A1(n11473), .A2(n7183), .ZN(n7176) );
  NAND2_X1 U8655 ( .A1(n7185), .A2(n12381), .ZN(n15230) );
  OR2_X1 U8656 ( .A1(n11473), .A2(n9757), .ZN(n7185) );
  NAND2_X1 U8657 ( .A1(n11229), .A2(n7149), .ZN(n15274) );
  INV_X1 U8658 ( .A(n11236), .ZN(n15305) );
  AND2_X1 U8659 ( .A1(n10820), .A2(n12608), .ZN(n15313) );
  OR3_X1 U8660 ( .A1(n10654), .A2(n12476), .A3(n15368), .ZN(n15312) );
  INV_X1 U8661 ( .A(n15312), .ZN(n15253) );
  INV_X1 U8662 ( .A(n12253), .ZN(n12930) );
  NAND2_X1 U8663 ( .A1(n9502), .A2(n9501), .ZN(n12944) );
  NAND2_X1 U8664 ( .A1(n10422), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12951) );
  XNOR2_X1 U8665 ( .A(n12315), .B(n11870), .ZN(n12299) );
  NAND2_X1 U8666 ( .A1(n7205), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7531) );
  NAND2_X1 U8667 ( .A1(n6777), .A2(n9720), .ZN(n11869) );
  NAND2_X1 U8668 ( .A1(n6801), .A2(n9689), .ZN(n9704) );
  INV_X1 U8669 ( .A(SI_26_), .ZN(n11609) );
  NAND2_X1 U8670 ( .A1(n9219), .A2(n9780), .ZN(n11610) );
  NAND2_X1 U8671 ( .A1(n7323), .A2(n9672), .ZN(n9687) );
  XNOR2_X1 U8672 ( .A(n9642), .B(n9641), .ZN(n11195) );
  NAND2_X1 U8673 ( .A1(n7333), .A2(n9628), .ZN(n9642) );
  NAND2_X1 U8674 ( .A1(n9616), .A2(n7337), .ZN(n7333) );
  NAND2_X1 U8675 ( .A1(n9616), .A2(n9615), .ZN(n9630) );
  OAI21_X1 U8676 ( .B1(n7315), .B2(n6786), .A(n6783), .ZN(n9601) );
  NAND2_X1 U8677 ( .A1(n6876), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9735) );
  INV_X1 U8678 ( .A(SI_20_), .ZN(n10751) );
  NAND2_X1 U8679 ( .A1(n6671), .A2(n9597), .ZN(n9598) );
  NAND2_X1 U8680 ( .A1(n9597), .A2(n9585), .ZN(n9586) );
  INV_X1 U8681 ( .A(n9820), .ZN(n10820) );
  NAND2_X1 U8682 ( .A1(n9568), .A2(n9567), .ZN(n9583) );
  NAND2_X1 U8683 ( .A1(n9533), .A2(n9532), .ZN(n9550) );
  INV_X1 U8684 ( .A(SI_16_), .ZN(n13582) );
  OAI21_X1 U8685 ( .B1(n7311), .B2(n7023), .A(n7021), .ZN(n9494) );
  INV_X1 U8686 ( .A(n9476), .ZN(n7023) );
  INV_X1 U8687 ( .A(SI_13_), .ZN(n13723) );
  AND2_X1 U8688 ( .A1(n7461), .A2(n7462), .ZN(n9463) );
  INV_X1 U8689 ( .A(SI_12_), .ZN(n10056) );
  INV_X1 U8690 ( .A(SI_11_), .ZN(n10044) );
  XNOR2_X1 U8691 ( .A(n9414), .B(n13665), .ZN(n12571) );
  OAI21_X1 U8692 ( .B1(n9390), .B2(n7330), .A(n7327), .ZN(n9420) );
  NAND2_X1 U8693 ( .A1(n9393), .A2(n9392), .ZN(n9410) );
  NAND2_X1 U8694 ( .A1(n9390), .A2(n9389), .ZN(n9393) );
  NAND2_X1 U8695 ( .A1(n7339), .A2(n7345), .ZN(n9368) );
  NAND2_X1 U8696 ( .A1(n9334), .A2(n7346), .ZN(n7339) );
  NAND2_X1 U8697 ( .A1(n7348), .A2(n9332), .ZN(n9349) );
  NAND2_X1 U8698 ( .A1(n7349), .A2(n7350), .ZN(n7348) );
  XNOR2_X1 U8699 ( .A(n9336), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10674) );
  OR3_X1 U8700 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n9271) );
  OR2_X1 U8701 ( .A1(n9254), .A2(n9231), .ZN(n9255) );
  OR3_X1 U8702 ( .A1(n9853), .A2(n9852), .A3(n9851), .ZN(n10170) );
  NAND2_X1 U8703 ( .A1(n6760), .A2(n7361), .ZN(n14446) );
  NAND2_X1 U8704 ( .A1(n7362), .A2(n9934), .ZN(n7361) );
  OR2_X1 U8705 ( .A1(n11436), .A2(n7363), .ZN(n7362) );
  NAND2_X1 U8706 ( .A1(n14446), .A2(n14447), .ZN(n14445) );
  AND2_X1 U8707 ( .A1(n9980), .A2(n9979), .ZN(n14450) );
  INV_X1 U8708 ( .A(n9869), .ZN(n7354) );
  XNOR2_X1 U8709 ( .A(n9860), .B(n9862), .ZN(n10457) );
  NOR2_X1 U8710 ( .A1(n11846), .A2(n11845), .ZN(n11844) );
  NAND2_X1 U8711 ( .A1(n7902), .A2(n7901), .ZN(n13437) );
  INV_X1 U8712 ( .A(n13249), .ZN(n13397) );
  NAND2_X1 U8713 ( .A1(n13088), .A2(n11012), .ZN(n10408) );
  NAND2_X1 U8714 ( .A1(n11379), .A2(n9929), .ZN(n11437) );
  NAND2_X1 U8715 ( .A1(n7365), .A2(n9916), .ZN(n11364) );
  CLKBUF_X1 U8716 ( .A(n8156), .Z(n6745) );
  NAND2_X1 U8717 ( .A1(n10448), .A2(n10449), .ZN(n10447) );
  INV_X1 U8718 ( .A(n13059), .ZN(n14448) );
  NAND2_X1 U8719 ( .A1(n6899), .A2(n6898), .ZN(n6897) );
  INV_X1 U8720 ( .A(n13052), .ZN(n6898) );
  OR2_X1 U8721 ( .A1(n13005), .A2(n12105), .ZN(n6899) );
  OR2_X1 U8722 ( .A1(n13005), .A2(n7370), .ZN(n13051) );
  XNOR2_X1 U8723 ( .A(n9943), .B(n9944), .ZN(n11700) );
  NAND2_X1 U8724 ( .A1(n9183), .A2(n9182), .ZN(n9184) );
  INV_X1 U8725 ( .A(n12969), .ZN(n13063) );
  NOR2_X1 U8726 ( .A1(n14947), .A2(n14946), .ZN(n14949) );
  AOI21_X1 U8727 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n14976), .A(n14971), .ZN(
        n14982) );
  NOR2_X1 U8728 ( .A1(n13134), .A2(n14994), .ZN(n15005) );
  AND2_X1 U8729 ( .A1(n15017), .A2(n15016), .ZN(n15020) );
  AND2_X1 U8730 ( .A1(n10172), .A2(n6740), .ZN(n15041) );
  NAND2_X1 U8731 ( .A1(n13179), .A2(n13178), .ZN(n13380) );
  NAND2_X1 U8732 ( .A1(n7033), .A2(n8192), .ZN(n13205) );
  NAND2_X1 U8733 ( .A1(n7032), .A2(n7411), .ZN(n13214) );
  NAND2_X1 U8734 ( .A1(n13243), .A2(n8190), .ZN(n13229) );
  NAND2_X1 U8735 ( .A1(n7064), .A2(n8043), .ZN(n13226) );
  NAND2_X1 U8736 ( .A1(n13240), .A2(n13246), .ZN(n7064) );
  NAND2_X1 U8737 ( .A1(n7415), .A2(n8183), .ZN(n13291) );
  NAND2_X1 U8738 ( .A1(n6751), .A2(n7421), .ZN(n7415) );
  NAND2_X1 U8739 ( .A1(n6751), .A2(n8181), .ZN(n13311) );
  NAND2_X1 U8740 ( .A1(n7057), .A2(n7957), .ZN(n13302) );
  NAND2_X1 U8741 ( .A1(n13318), .A2(n7956), .ZN(n7057) );
  CLKBUF_X1 U8742 ( .A(n13315), .Z(n13316) );
  CLKBUF_X1 U8743 ( .A(n13362), .Z(n13364) );
  NAND2_X1 U8744 ( .A1(n11462), .A2(n7813), .ZN(n11554) );
  OAI21_X1 U8745 ( .B1(n11483), .B2(n8167), .A(n8169), .ZN(n11458) );
  CLKBUF_X1 U8746 ( .A(n11342), .Z(n11343) );
  NAND2_X1 U8747 ( .A1(n7756), .A2(n7755), .ZN(n11356) );
  NAND2_X1 U8748 ( .A1(n11044), .A2(n8164), .ZN(n11209) );
  INV_X1 U8749 ( .A(n13365), .ZN(n15063) );
  AND2_X2 U8750 ( .A1(n11590), .A2(n11373), .ZN(n11005) );
  INV_X1 U8751 ( .A(n10407), .ZN(n11012) );
  NAND2_X1 U8752 ( .A1(n15103), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7081) );
  INV_X1 U8753 ( .A(n13165), .ZN(n13457) );
  OAI211_X1 U8754 ( .C1(n13380), .C2(n13440), .A(n13378), .B(n13379), .ZN(
        n13458) );
  NAND2_X1 U8755 ( .A1(n7863), .A2(n7862), .ZN(n11841) );
  NOR2_X1 U8756 ( .A1(n15076), .A2(n15067), .ZN(n15073) );
  INV_X1 U8757 ( .A(n15078), .ZN(n15076) );
  AND2_X1 U8758 ( .A1(n9975), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15078) );
  NAND2_X1 U8759 ( .A1(n7109), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7554) );
  CLKBUF_X1 U8760 ( .A(n13484), .Z(n6740) );
  INV_X1 U8761 ( .A(n9851), .ZN(n13768) );
  XNOR2_X1 U8762 ( .A(n8206), .B(P2_IR_REG_25__SCAN_IN), .ZN(n13773) );
  XNOR2_X1 U8763 ( .A(n8204), .B(P2_IR_REG_24__SCAN_IN), .ZN(n11696) );
  INV_X1 U8764 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13595) );
  INV_X1 U8765 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11591) );
  INV_X1 U8766 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11135) );
  INV_X1 U8767 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n13735) );
  INV_X1 U8768 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10774) );
  INV_X1 U8769 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10416) );
  INV_X1 U8770 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10315) );
  INV_X1 U8771 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10202) );
  INV_X1 U8772 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10047) );
  INV_X1 U8773 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10014) );
  CLKBUF_X1 U8774 ( .A(n7631), .Z(n7632) );
  INV_X1 U8775 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10003) );
  XNOR2_X1 U8776 ( .A(n7571), .B(n7570), .ZN(n14868) );
  AND2_X1 U8777 ( .A1(n7582), .A2(n7581), .ZN(n13778) );
  CLKBUF_X1 U8778 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n13777) );
  NAND2_X1 U8779 ( .A1(n6915), .A2(n7499), .ZN(n13779) );
  NAND2_X1 U8780 ( .A1(n8524), .A2(n8523), .ZN(n14598) );
  NAND2_X1 U8781 ( .A1(n13850), .A2(n12042), .ZN(n13786) );
  NOR2_X1 U8782 ( .A1(n6923), .A2(n7529), .ZN(n6922) );
  INV_X1 U8783 ( .A(n10766), .ZN(n6923) );
  NAND2_X1 U8784 ( .A1(n7511), .A2(n7509), .ZN(n13797) );
  NAND2_X1 U8785 ( .A1(n7511), .A2(n12016), .ZN(n13796) );
  NAND2_X1 U8786 ( .A1(n6912), .A2(n6911), .ZN(n6910) );
  NAND2_X1 U8787 ( .A1(n6914), .A2(n12083), .ZN(n6913) );
  NAND2_X1 U8788 ( .A1(n7516), .A2(n7517), .ZN(n11596) );
  NOR2_X1 U8789 ( .A1(n11514), .A2(n11513), .ZN(n11515) );
  NAND2_X1 U8790 ( .A1(n13829), .A2(n12028), .ZN(n13807) );
  NAND2_X1 U8791 ( .A1(n14531), .A2(n11797), .ZN(n11803) );
  INV_X1 U8792 ( .A(n11174), .ZN(n6908) );
  NAND2_X1 U8793 ( .A1(n11254), .A2(n11255), .ZN(n6907) );
  INV_X1 U8794 ( .A(n6902), .ZN(n6901) );
  OAI21_X1 U8795 ( .B1(n11994), .B2(n7497), .A(n12001), .ZN(n6902) );
  AOI21_X1 U8796 ( .B1(n7506), .B2(n7508), .A(n6651), .ZN(n7504) );
  AOI21_X1 U8797 ( .B1(n7517), .B2(n7515), .A(n6660), .ZN(n7514) );
  INV_X1 U8798 ( .A(n11402), .ZN(n7515) );
  OAI21_X1 U8799 ( .B1(n7511), .B2(n6938), .A(n6936), .ZN(n13829) );
  NAND2_X1 U8800 ( .A1(n13797), .A2(n12024), .ZN(n13831) );
  NOR2_X1 U8801 ( .A1(n10498), .A2(n10497), .ZN(n10503) );
  INV_X1 U8802 ( .A(n6924), .ZN(n10761) );
  AND2_X1 U8803 ( .A1(n10778), .A2(n11583), .ZN(n14517) );
  NAND2_X1 U8804 ( .A1(n10303), .A2(n14739), .ZN(n14536) );
  NAND2_X1 U8805 ( .A1(n7500), .A2(n12063), .ZN(n13878) );
  NAND2_X1 U8806 ( .A1(n13814), .A2(n13815), .ZN(n7500) );
  NAND2_X1 U8807 ( .A1(n14542), .A2(n14543), .ZN(n14541) );
  OR3_X1 U8808 ( .A1(n8294), .A2(n8293), .A3(n8292), .ZN(n13994) );
  OAI211_X1 U8809 ( .C1(n14137), .C2(n8701), .A(n8619), .B(n8618), .ZN(n14146)
         );
  INV_X1 U8810 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10237) );
  AND4_X1 U8811 ( .A1(n8462), .A2(n8461), .A3(n8460), .A4(n8459), .ZN(n11598)
         );
  INV_X1 U8812 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10235) );
  AND4_X1 U8813 ( .A1(n8452), .A2(n8451), .A3(n8450), .A4(n8449), .ZN(n11600)
         );
  NAND4_X1 U8814 ( .A1(n8372), .A2(n8371), .A3(n8370), .A4(n8369), .ZN(n13896)
         );
  NAND2_X1 U8815 ( .A1(n8258), .A2(n6836), .ZN(n8545) );
  AND2_X1 U8816 ( .A1(n8257), .A2(n8352), .ZN(n6836) );
  INV_X1 U8817 ( .A(n13998), .ZN(n14194) );
  INV_X1 U8818 ( .A(n6996), .ZN(n14199) );
  NAND2_X1 U8819 ( .A1(n7297), .A2(n7295), .ZN(n7294) );
  NAND2_X1 U8820 ( .A1(n11952), .A2(n11951), .ZN(n11953) );
  AND2_X1 U8821 ( .A1(n14006), .A2(n14005), .ZN(n14207) );
  NAND2_X1 U8822 ( .A1(n14040), .A2(n11903), .ZN(n14024) );
  AND2_X1 U8823 ( .A1(n14075), .A2(n11900), .ZN(n14053) );
  NAND2_X1 U8824 ( .A1(n14090), .A2(n11898), .ZN(n14073) );
  NAND2_X1 U8825 ( .A1(n7385), .A2(n7386), .ZN(n14120) );
  NAND2_X1 U8826 ( .A1(n14153), .A2(n7389), .ZN(n7385) );
  NAND2_X1 U8827 ( .A1(n14131), .A2(n11922), .ZN(n14119) );
  OAI21_X1 U8828 ( .B1(n14153), .B2(n11896), .A(n11895), .ZN(n14130) );
  NAND2_X1 U8829 ( .A1(n8596), .A2(n8595), .ZN(n14575) );
  NAND2_X1 U8830 ( .A1(n7262), .A2(n7264), .ZN(n14158) );
  NAND2_X1 U8831 ( .A1(n7267), .A2(n11915), .ZN(n14172) );
  NAND2_X1 U8832 ( .A1(n14563), .A2(n11914), .ZN(n7267) );
  OAI21_X1 U8833 ( .B1(n11415), .B2(n6818), .A(n6816), .ZN(n11537) );
  NAND2_X1 U8834 ( .A1(n6821), .A2(n11535), .ZN(n11574) );
  NAND2_X1 U8835 ( .A1(n11415), .A2(n6822), .ZN(n6821) );
  NAND2_X1 U8836 ( .A1(n7285), .A2(n11524), .ZN(n11576) );
  NAND2_X1 U8837 ( .A1(n11410), .A2(n11409), .ZN(n11526) );
  INV_X1 U8838 ( .A(n14825), .ZN(n14705) );
  NAND2_X1 U8839 ( .A1(n10302), .A2(n11582), .ZN(n14739) );
  NAND2_X1 U8840 ( .A1(n7379), .A2(n10782), .ZN(n10935) );
  NAND2_X1 U8841 ( .A1(n10958), .A2(n10952), .ZN(n7379) );
  OR2_X1 U8842 ( .A1(n14157), .A2(n14560), .ZN(n14337) );
  NAND2_X1 U8843 ( .A1(n10064), .A2(n6598), .ZN(n7395) );
  INV_X1 U8844 ( .A(n14339), .ZN(n14570) );
  NOR2_X1 U8845 ( .A1(n14157), .A2(n14837), .ZN(n14571) );
  INV_X1 U8846 ( .A(n14337), .ZN(n14743) );
  AND2_X2 U8847 ( .A1(n11585), .A2(n11571), .ZN(n14858) );
  OAI21_X1 U8848 ( .B1(n14201), .B2(n14793), .A(n6750), .ZN(n14271) );
  AOI21_X1 U8849 ( .B1(n14200), .B2(n14738), .A(n6735), .ZN(n6750) );
  NAND2_X1 U8850 ( .A1(n6996), .A2(n6736), .ZN(n6735) );
  INV_X1 U8851 ( .A(n14198), .ZN(n6736) );
  AND2_X2 U8852 ( .A1(n11585), .A2(n11584), .ZN(n14844) );
  INV_X1 U8853 ( .A(n10054), .ZN(n10072) );
  XNOR2_X1 U8854 ( .A(n8250), .B(n8249), .ZN(n14285) );
  AND2_X1 U8855 ( .A1(n8284), .A2(n8287), .ZN(n7520) );
  NOR2_X1 U8856 ( .A1(n8265), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n8286) );
  CLKBUF_X1 U8857 ( .A(n8835), .Z(n11878) );
  XNOR2_X1 U8858 ( .A(n8093), .B(n8081), .ZN(n14293) );
  NAND2_X1 U8859 ( .A1(n8831), .A2(n8830), .ZN(n14301) );
  INV_X1 U8860 ( .A(n7397), .ZN(n8831) );
  XNOR2_X1 U8861 ( .A(n8080), .B(n8063), .ZN(n14297) );
  XNOR2_X1 U8862 ( .A(n8824), .B(n8823), .ZN(n14305) );
  NAND2_X1 U8863 ( .A1(n6939), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8824) );
  NAND2_X1 U8864 ( .A1(n7030), .A2(n8031), .ZN(n11697) );
  AND2_X1 U8865 ( .A1(n7076), .A2(P1_U3086), .ZN(n14292) );
  XNOR2_X1 U8866 ( .A(n8657), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14308) );
  OR2_X1 U8867 ( .A1(n8656), .A2(n8655), .ZN(n8657) );
  INV_X1 U8868 ( .A(n10788), .ZN(n14307) );
  NAND2_X1 U8869 ( .A1(n7441), .A2(n7439), .ZN(n7995) );
  NAND2_X1 U8870 ( .A1(n7441), .A2(n7976), .ZN(n7981) );
  INV_X1 U8871 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n13560) );
  NAND2_X1 U8872 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n6944) );
  NOR2_X1 U8873 ( .A1(n8588), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n6945) );
  INV_X1 U8874 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11132) );
  INV_X1 U8875 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10773) );
  INV_X1 U8876 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10717) );
  INV_X1 U8877 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10414) );
  INV_X1 U8878 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10312) );
  INV_X1 U8879 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10199) );
  INV_X1 U8880 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10161) );
  INV_X1 U8881 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n13553) );
  INV_X1 U8882 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10075) );
  INV_X1 U8883 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10059) );
  INV_X1 U8884 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10048) );
  INV_X1 U8885 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10041) );
  XNOR2_X1 U8886 ( .A(n7590), .B(n7591), .ZN(n10009) );
  XNOR2_X1 U8887 ( .A(n8900), .B(n14914), .ZN(n14323) );
  AND2_X1 U8888 ( .A1(n6851), .A2(n6853), .ZN(n14332) );
  OAI21_X1 U8889 ( .B1(n8907), .B2(n6850), .A(n6849), .ZN(n6851) );
  INV_X1 U8890 ( .A(n14626), .ZN(n7214) );
  INV_X1 U8891 ( .A(n14625), .ZN(n7215) );
  AND2_X1 U8892 ( .A1(n7207), .A2(n7206), .ZN(n14348) );
  NAND2_X1 U8893 ( .A1(n7208), .A2(n15015), .ZN(n7207) );
  NAND2_X1 U8894 ( .A1(n14633), .A2(n14634), .ZN(n7208) );
  NOR2_X1 U8895 ( .A1(n14348), .A2(n14347), .ZN(n14346) );
  NAND2_X1 U8896 ( .A1(n10850), .A2(n10849), .ZN(n10854) );
  XNOR2_X1 U8897 ( .A(n6864), .B(n7488), .ZN(n12284) );
  NAND2_X1 U8898 ( .A1(n7313), .A2(n7312), .ZN(P3_U3296) );
  OR2_X1 U8899 ( .A1(n12511), .A2(n12510), .ZN(n7312) );
  NAND2_X1 U8900 ( .A1(n7024), .A2(n7314), .ZN(n7313) );
  XNOR2_X1 U8901 ( .A(n6763), .B(n6728), .ZN(n12610) );
  OAI21_X1 U8902 ( .B1(n12628), .B2(n12949), .A(n7528), .ZN(n9848) );
  OR4_X1 U8903 ( .A1(n9984), .A2(n9983), .A3(n9982), .A4(n9981), .ZN(P2_U3207)
         );
  NAND2_X1 U8904 ( .A1(n10525), .A2(n9889), .ZN(n10567) );
  INV_X1 U8905 ( .A(n6758), .ZN(n6757) );
  NAND2_X1 U8906 ( .A1(n13162), .A2(n13161), .ZN(n6759) );
  NAND2_X1 U8907 ( .A1(n13163), .A2(n11192), .ZN(n6756) );
  AOI21_X1 U8908 ( .B1(n11885), .B2(n14467), .A(n11884), .ZN(n6762) );
  NAND2_X1 U8909 ( .A1(n7082), .A2(n7079), .ZN(P2_U3527) );
  INV_X1 U8910 ( .A(n7080), .ZN(n7079) );
  NAND2_X1 U8911 ( .A1(n13458), .A2(n15105), .ZN(n7082) );
  OAI21_X1 U8912 ( .B1(n13459), .B2(n13418), .A(n7081), .ZN(n7080) );
  INV_X1 U8913 ( .A(n6767), .ZN(P2_U3495) );
  AOI21_X1 U8914 ( .B1(n13458), .B2(n15099), .A(n6768), .ZN(n6767) );
  OAI21_X1 U8915 ( .B1(n13459), .B2(n13468), .A(n6769), .ZN(n6768) );
  NAND2_X1 U8916 ( .A1(n15098), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6769) );
  NAND2_X1 U8917 ( .A1(n6833), .A2(n6832), .ZN(P1_U3525) );
  OR2_X1 U8918 ( .A1(n14844), .A2(n8750), .ZN(n6832) );
  NAND2_X1 U8919 ( .A1(n14271), .A2(n14844), .ZN(n6833) );
  NAND2_X1 U8920 ( .A1(n6855), .A2(n6853), .ZN(n14329) );
  NOR2_X1 U8921 ( .A1(n6708), .A2(n14618), .ZN(n14617) );
  NOR2_X1 U8922 ( .A1(n8920), .A2(n8921), .ZN(n14622) );
  INV_X1 U8923 ( .A(n7206), .ZN(n14632) );
  XNOR2_X1 U8924 ( .A(n7218), .B(n7217), .ZN(SUB_1596_U4) );
  XNOR2_X1 U8925 ( .A(n8941), .B(n6729), .ZN(n7217) );
  OAI21_X1 U8926 ( .B1(n14311), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6642), .ZN(
        n7218) );
  AND2_X1 U8927 ( .A1(n8735), .A2(n8737), .ZN(n6590) );
  INV_X2 U8928 ( .A(n7535), .ZN(n9122) );
  AND2_X1 U8929 ( .A1(n7199), .A2(n12612), .ZN(n6591) );
  OR2_X1 U8930 ( .A1(n7853), .A2(n7040), .ZN(n6592) );
  INV_X1 U8931 ( .A(n14118), .ZN(n7305) );
  NAND2_X1 U8932 ( .A1(n9784), .A2(n6649), .ZN(n7205) );
  AOI21_X1 U8933 ( .B1(n9476), .B2(n10319), .A(n7022), .ZN(n7021) );
  INV_X1 U8934 ( .A(n9333), .ZN(n7350) );
  AND4_X1 U8935 ( .A1(n9287), .A2(n9286), .A3(n9285), .A4(n9284), .ZN(n10841)
         );
  AND2_X1 U8936 ( .A1(n14054), .A2(n11900), .ZN(n6593) );
  AND2_X1 U8937 ( .A1(n7474), .A2(n7472), .ZN(n6594) );
  AND2_X1 U8938 ( .A1(n11459), .A2(n8168), .ZN(n6595) );
  AND2_X1 U8939 ( .A1(n8101), .A2(n8100), .ZN(n13459) );
  INV_X1 U8940 ( .A(n13459), .ZN(n7104) );
  AND2_X1 U8941 ( .A1(n12418), .A2(n12422), .ZN(n12492) );
  AND2_X1 U8942 ( .A1(n6991), .A2(n6990), .ZN(n6596) );
  AND2_X1 U8943 ( .A1(n14214), .A2(n14012), .ZN(n6597) );
  AND2_X1 U8944 ( .A1(n10005), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6598) );
  AND2_X1 U8945 ( .A1(n8655), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U8946 ( .A1(n8548), .A2(n8547), .ZN(n14592) );
  INV_X1 U8947 ( .A(n11973), .ZN(n13847) );
  AND2_X1 U8948 ( .A1(n8543), .A2(n8542), .ZN(n11973) );
  AND2_X1 U8949 ( .A1(n6670), .A2(n6934), .ZN(n6600) );
  NOR2_X1 U8950 ( .A1(n14592), .A2(n14507), .ZN(n6601) );
  AND2_X1 U8951 ( .A1(n10047), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6602) );
  NAND2_X1 U8952 ( .A1(n7821), .A2(n7820), .ZN(n11563) );
  AND2_X1 U8953 ( .A1(n6724), .A2(n11255), .ZN(n6603) );
  AND2_X1 U8954 ( .A1(n6873), .A2(n9539), .ZN(n6604) );
  AND2_X1 U8955 ( .A1(n12506), .A2(n12505), .ZN(n6605) );
  NAND2_X1 U8956 ( .A1(n6933), .A2(n6932), .ZN(n11793) );
  AND2_X1 U8957 ( .A1(n12310), .A2(n12309), .ZN(n12612) );
  AND2_X1 U8958 ( .A1(n7316), .A2(n7319), .ZN(n6606) );
  INV_X1 U8959 ( .A(n7096), .ZN(n7094) );
  INV_X1 U8960 ( .A(n11242), .ZN(n7085) );
  AND2_X1 U8961 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n6778), .ZN(n6607) );
  INV_X1 U8962 ( .A(n10391), .ZN(n11597) );
  NAND2_X1 U8963 ( .A1(n11719), .A2(n12520), .ZN(n6608) );
  OR2_X1 U8964 ( .A1(n12580), .A2(n12553), .ZN(n6609) );
  XNOR2_X1 U8965 ( .A(n9735), .B(n9734), .ZN(n10819) );
  INV_X1 U8966 ( .A(n11895), .ZN(n7390) );
  XNOR2_X1 U8967 ( .A(n12705), .B(n12687), .ZN(n12706) );
  INV_X1 U8968 ( .A(n12706), .ZN(n7170) );
  INV_X1 U8969 ( .A(n13898), .ZN(n7261) );
  NOR2_X1 U8970 ( .A1(n7347), .A2(n9348), .ZN(n7346) );
  AND2_X1 U8971 ( .A1(n14108), .A2(n7003), .ZN(n6610) );
  AND2_X1 U8972 ( .A1(n6813), .A2(n6811), .ZN(n6611) );
  AND2_X1 U8973 ( .A1(n6878), .A2(n7044), .ZN(n6612) );
  AND2_X1 U8974 ( .A1(n9750), .A2(n9260), .ZN(n6613) );
  OR2_X1 U8975 ( .A1(n8913), .A2(n8912), .ZN(n6614) );
  NAND2_X1 U8976 ( .A1(n9955), .A2(n9954), .ZN(n6615) );
  NOR2_X1 U8977 ( .A1(n12673), .A2(n12666), .ZN(n6616) );
  NOR2_X1 U8978 ( .A1(n12491), .A2(n12794), .ZN(n6617) );
  AND2_X1 U8979 ( .A1(n10264), .A2(n10263), .ZN(n6618) );
  NAND2_X1 U8980 ( .A1(n7505), .A2(n7504), .ZN(n13822) );
  NAND2_X1 U8981 ( .A1(n11637), .A2(n11636), .ZN(n6619) );
  OR2_X1 U8982 ( .A1(n10428), .A2(n10546), .ZN(n6620) );
  NAND2_X1 U8983 ( .A1(n14541), .A2(n11994), .ZN(n14505) );
  NAND2_X1 U8984 ( .A1(n9482), .A2(n7160), .ZN(n9219) );
  AND2_X1 U8985 ( .A1(n9571), .A2(n6875), .ZN(n6621) );
  INV_X1 U8986 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U8987 ( .A1(n7984), .A2(n7983), .ZN(n13295) );
  INV_X1 U8988 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n10731) );
  AND2_X1 U8989 ( .A1(n7884), .A2(n7883), .ZN(n13445) );
  INV_X1 U8990 ( .A(n13445), .ZN(n11829) );
  AND2_X1 U8991 ( .A1(n12706), .A2(n7169), .ZN(n6622) );
  AND2_X1 U8992 ( .A1(n12129), .A2(n12127), .ZN(n6623) );
  AND2_X1 U8993 ( .A1(n12523), .A2(n15281), .ZN(n6624) );
  INV_X1 U8994 ( .A(n9006), .ZN(n7117) );
  INV_X1 U8995 ( .A(n9072), .ZN(n7122) );
  AND2_X1 U8996 ( .A1(n11339), .A2(n13078), .ZN(n6625) );
  NAND2_X1 U8997 ( .A1(n9784), .A2(n7473), .ZN(n6626) );
  INV_X1 U8998 ( .A(n12083), .ZN(n6920) );
  NAND2_X1 U8999 ( .A1(n7597), .A2(n7599), .ZN(n7613) );
  NAND2_X1 U9000 ( .A1(n8685), .A2(n8684), .ZN(n14068) );
  NAND2_X1 U9001 ( .A1(n9229), .A2(n7151), .ZN(n12827) );
  INV_X1 U9002 ( .A(n12827), .ZN(n10876) );
  AND2_X1 U9003 ( .A1(n11425), .A2(n12522), .ZN(n6627) );
  AND2_X1 U9004 ( .A1(n13420), .A2(n7973), .ZN(n6628) );
  INV_X1 U9005 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6844) );
  AND2_X1 U9006 ( .A1(n12130), .A2(n12518), .ZN(n6629) );
  NAND2_X1 U9007 ( .A1(n8272), .A2(n7396), .ZN(n8265) );
  INV_X1 U9008 ( .A(n8265), .ZN(n8285) );
  AND2_X1 U9009 ( .A1(n13392), .A2(n13066), .ZN(n6630) );
  NAND2_X1 U9010 ( .A1(n8581), .A2(n8580), .ZN(n14184) );
  NOR2_X1 U9011 ( .A1(n9043), .A2(n9045), .ZN(n6631) );
  OR2_X1 U9012 ( .A1(n10550), .A2(n9280), .ZN(n6632) );
  AND2_X1 U9013 ( .A1(n13392), .A2(n8057), .ZN(n6633) );
  NOR2_X1 U9014 ( .A1(n11150), .A2(n7366), .ZN(n6634) );
  INV_X1 U9015 ( .A(n7815), .ZN(n7043) );
  INV_X1 U9016 ( .A(n11903), .ZN(n7393) );
  AND2_X1 U9017 ( .A1(n12640), .A2(n7011), .ZN(n6635) );
  AND2_X1 U9018 ( .A1(n8649), .A2(n8648), .ZN(n6636) );
  NOR2_X1 U9019 ( .A1(n12363), .A2(n15272), .ZN(n6637) );
  NOR2_X1 U9020 ( .A1(n14368), .A2(n14367), .ZN(n6638) );
  NAND2_X1 U9021 ( .A1(n7840), .A2(n7839), .ZN(n14461) );
  AND2_X1 U9022 ( .A1(n7512), .A2(n6926), .ZN(n6639) );
  INV_X1 U9023 ( .A(n8985), .ZN(n7125) );
  AND2_X1 U9024 ( .A1(n7192), .A2(n7190), .ZN(n6640) );
  OR2_X1 U9025 ( .A1(n8638), .A2(n8639), .ZN(n6641) );
  OR2_X1 U9026 ( .A1(n8935), .A2(n8936), .ZN(n6642) );
  AND2_X1 U9027 ( .A1(n11142), .A2(n11138), .ZN(n6643) );
  AND2_X1 U9028 ( .A1(n7656), .A2(n7629), .ZN(n6644) );
  AND2_X1 U9029 ( .A1(n12189), .A2(n12763), .ZN(n6645) );
  NAND2_X1 U9030 ( .A1(n6593), .A2(n11903), .ZN(n6646) );
  AND2_X1 U9031 ( .A1(n6614), .A2(n6840), .ZN(n6647) );
  AND2_X1 U9032 ( .A1(n9217), .A2(n7204), .ZN(n6648) );
  AND2_X1 U9033 ( .A1(n6594), .A2(n6648), .ZN(n6649) );
  AND2_X1 U9034 ( .A1(n12467), .A2(n12468), .ZN(n6650) );
  AND2_X1 U9035 ( .A1(n12048), .A2(n12047), .ZN(n6651) );
  AND2_X1 U9036 ( .A1(n12070), .A2(n12069), .ZN(n6652) );
  INV_X1 U9037 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8826) );
  INV_X1 U9038 ( .A(n11512), .ZN(n11513) );
  AND2_X1 U9039 ( .A1(n14184), .A2(n14558), .ZN(n6653) );
  AND2_X1 U9040 ( .A1(n12076), .A2(n12075), .ZN(n6654) );
  AND2_X1 U9041 ( .A1(n8123), .A2(n8122), .ZN(n11882) );
  INV_X1 U9042 ( .A(n11882), .ZN(n7099) );
  AND2_X1 U9043 ( .A1(n11610), .A2(n11378), .ZN(n6655) );
  NOR2_X1 U9044 ( .A1(n11799), .A2(n13890), .ZN(n6656) );
  OR2_X1 U9045 ( .A1(n9185), .A2(n9184), .ZN(n6657) );
  NOR2_X1 U9046 ( .A1(n12720), .A2(n12701), .ZN(n6658) );
  NOR2_X1 U9047 ( .A1(n14252), .A2(n13799), .ZN(n6659) );
  NOR2_X1 U9048 ( .A1(n11595), .A2(n11594), .ZN(n6660) );
  INV_X1 U9049 ( .A(n8393), .ZN(n7254) );
  AND2_X1 U9050 ( .A1(n12521), .A2(n11707), .ZN(n6661) );
  NAND2_X1 U9051 ( .A1(n8270), .A2(n6940), .ZN(n6662) );
  OR2_X1 U9052 ( .A1(n8844), .A2(n8843), .ZN(n6663) );
  OR2_X1 U9053 ( .A1(n12470), .A2(n12612), .ZN(n6664) );
  AND4_X1 U9054 ( .A1(n8260), .A2(n6989), .A3(n8259), .A4(n8277), .ZN(n6665)
         );
  OR2_X1 U9055 ( .A1(n10552), .A2(n10542), .ZN(n6666) );
  NOR2_X1 U9056 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7597) );
  OR2_X1 U9057 ( .A1(n11563), .A2(n14442), .ZN(n6667) );
  AND2_X1 U9058 ( .A1(n7753), .A2(SI_9_), .ZN(n6668) );
  NOR2_X1 U9059 ( .A1(n11799), .A2(n14527), .ZN(n6669) );
  INV_X1 U9060 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8822) );
  INV_X1 U9061 ( .A(n7150), .ZN(n7149) );
  NAND2_X1 U9062 ( .A1(n15275), .A2(n9324), .ZN(n7150) );
  INV_X1 U9063 ( .A(n7157), .ZN(n7156) );
  NAND2_X1 U9064 ( .A1(n7537), .A2(n9563), .ZN(n7157) );
  INV_X1 U9065 ( .A(n7518), .ZN(n7517) );
  NAND2_X1 U9066 ( .A1(n11516), .A2(n11512), .ZN(n7518) );
  AND2_X1 U9067 ( .A1(n8083), .A2(n8082), .ZN(n13202) );
  INV_X1 U9068 ( .A(n13202), .ZN(n7105) );
  AND2_X1 U9069 ( .A1(n12030), .A2(n12028), .ZN(n6670) );
  AND2_X1 U9070 ( .A1(n9585), .A2(n7027), .ZN(n6671) );
  AND2_X1 U9071 ( .A1(n7216), .A2(n7213), .ZN(n6672) );
  INV_X1 U9072 ( .A(n8747), .ZN(n6977) );
  INV_X1 U9073 ( .A(n8735), .ZN(n7434) );
  NAND2_X1 U9074 ( .A1(n11915), .A2(n11912), .ZN(n6673) );
  INV_X1 U9075 ( .A(n8697), .ZN(n6950) );
  INV_X1 U9076 ( .A(n8761), .ZN(n7247) );
  AND2_X1 U9077 ( .A1(n6916), .A2(n6920), .ZN(n6674) );
  OR2_X1 U9078 ( .A1(n8899), .A2(n8898), .ZN(n6675) );
  NAND2_X1 U9079 ( .A1(n8497), .A2(n8496), .ZN(n14537) );
  OR2_X1 U9080 ( .A1(n10676), .A2(n10672), .ZN(n6676) );
  AND2_X1 U9081 ( .A1(n6815), .A2(n11536), .ZN(n6677) );
  AND2_X1 U9082 ( .A1(n11095), .A2(n11096), .ZN(n6678) );
  OR2_X1 U9083 ( .A1(n6916), .A2(n6920), .ZN(n6679) );
  AND2_X1 U9084 ( .A1(n7248), .A2(n6976), .ZN(n6680) );
  AND2_X1 U9085 ( .A1(n9934), .A2(n11381), .ZN(n6681) );
  AND2_X1 U9086 ( .A1(n6941), .A2(n8826), .ZN(n6682) );
  AND2_X1 U9087 ( .A1(n11916), .A2(n7264), .ZN(n6683) );
  NAND2_X1 U9088 ( .A1(n13387), .A2(n13065), .ZN(n6684) );
  NAND2_X1 U9089 ( .A1(n12171), .A2(n12517), .ZN(n6685) );
  INV_X1 U9090 ( .A(n9401), .ZN(n7147) );
  NOR2_X1 U9091 ( .A1(n11914), .A2(n6827), .ZN(n6826) );
  AND2_X1 U9092 ( .A1(n14477), .A2(n7095), .ZN(n6686) );
  NOR2_X1 U9093 ( .A1(n14174), .A2(n7266), .ZN(n7265) );
  AND2_X1 U9094 ( .A1(n9890), .A2(n9889), .ZN(n6687) );
  NAND2_X1 U9095 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n6688) );
  AND2_X1 U9096 ( .A1(n14052), .A2(n11902), .ZN(n6689) );
  AND2_X1 U9097 ( .A1(n11899), .A2(n11898), .ZN(n6690) );
  AND2_X1 U9098 ( .A1(n9613), .A2(n9595), .ZN(n6691) );
  INV_X1 U9099 ( .A(n8518), .ZN(n6985) );
  OR2_X1 U9100 ( .A1(n9054), .A2(n9052), .ZN(n6692) );
  OR2_X1 U9101 ( .A1(n8984), .A2(n7125), .ZN(n6693) );
  OR2_X1 U9102 ( .A1(n9091), .A2(n9089), .ZN(n6694) );
  OR2_X1 U9103 ( .A1(n8996), .A2(n8994), .ZN(n6695) );
  OR2_X1 U9104 ( .A1(n7117), .A2(n9005), .ZN(n6696) );
  AND2_X1 U9105 ( .A1(n7399), .A2(n7398), .ZN(n6697) );
  AND2_X1 U9106 ( .A1(n6732), .A2(n6730), .ZN(n6698) );
  OR2_X1 U9107 ( .A1(n9015), .A2(n9017), .ZN(n6699) );
  OR2_X1 U9108 ( .A1(n9026), .A2(n9028), .ZN(n6700) );
  OR2_X1 U9109 ( .A1(n9071), .A2(n7122), .ZN(n6701) );
  AND2_X1 U9110 ( .A1(n6621), .A2(n6874), .ZN(n6702) );
  INV_X1 U9111 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8131) );
  INV_X1 U9112 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7621) );
  INV_X1 U9113 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9464) );
  AND2_X1 U9114 ( .A1(n8191), .A2(n7049), .ZN(n7413) );
  OR2_X1 U9115 ( .A1(n8668), .A2(n7257), .ZN(n6703) );
  NAND2_X1 U9116 ( .A1(n8591), .A2(n8590), .ZN(n14265) );
  NAND2_X1 U9117 ( .A1(n8736), .A2(n7434), .ZN(n6704) );
  INV_X1 U9118 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n6875) );
  OR2_X1 U9119 ( .A1(n12478), .A2(n12476), .ZN(n6705) );
  INV_X1 U9120 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n6874) );
  INV_X1 U9121 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6989) );
  INV_X1 U9122 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7054) );
  INV_X1 U9123 ( .A(n12278), .ZN(n7488) );
  INV_X1 U9124 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n7005) );
  NAND2_X1 U9125 ( .A1(n14308), .A2(n10064), .ZN(n14101) );
  INV_X1 U9126 ( .A(n14101), .ZN(n7004) );
  NAND2_X1 U9127 ( .A1(n8012), .A2(n8011), .ZN(n13404) );
  INV_X1 U9128 ( .A(n13404), .ZN(n7088) );
  NAND2_X1 U9129 ( .A1(n14564), .A2(n6596), .ZN(n6706) );
  NOR2_X1 U9130 ( .A1(n12939), .A2(n12228), .ZN(n6707) );
  INV_X1 U9131 ( .A(n12531), .ZN(n12564) );
  AND2_X1 U9132 ( .A1(n6837), .A2(n6614), .ZN(n6708) );
  NAND2_X1 U9133 ( .A1(n11474), .A2(n9401), .ZN(n15231) );
  INV_X1 U9134 ( .A(n14221), .ZN(n7000) );
  OAI21_X1 U9135 ( .B1(n11639), .B2(n6931), .A(n6928), .ZN(n14531) );
  INV_X1 U9136 ( .A(n12701), .ZN(n12731) );
  NAND2_X1 U9137 ( .A1(n9482), .A2(n6873), .ZN(n9538) );
  AND2_X1 U9138 ( .A1(n11921), .A2(n11920), .ZN(n6709) );
  AND2_X1 U9139 ( .A1(n7437), .A2(n7435), .ZN(n6710) );
  NOR2_X1 U9140 ( .A1(n7980), .A2(n7440), .ZN(n7439) );
  AND2_X1 U9141 ( .A1(n11736), .A2(n12519), .ZN(n6711) );
  INV_X1 U9142 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10319) );
  NOR2_X1 U9143 ( .A1(n6623), .A2(n7471), .ZN(n7470) );
  INV_X1 U9144 ( .A(n8921), .ZN(n7216) );
  NAND2_X1 U9145 ( .A1(n12321), .A2(n12320), .ZN(n12897) );
  INV_X1 U9146 ( .A(n12897), .ZN(n7195) );
  OR2_X1 U9147 ( .A1(n7491), .A2(n12218), .ZN(n7490) );
  AND2_X1 U9148 ( .A1(n7385), .A2(n7383), .ZN(n6712) );
  NOR2_X1 U9149 ( .A1(n11915), .A2(n8780), .ZN(n6713) );
  NOR2_X1 U9150 ( .A1(n12944), .A2(n12175), .ZN(n6714) );
  INV_X1 U9151 ( .A(n7516), .ZN(n11514) );
  NAND2_X1 U9152 ( .A1(n11401), .A2(n11402), .ZN(n7516) );
  INV_X1 U9153 ( .A(n8582), .ZN(n6959) );
  NOR2_X1 U9154 ( .A1(n14622), .A2(n14621), .ZN(n6715) );
  AND2_X1 U9155 ( .A1(n12761), .A2(n9563), .ZN(n6716) );
  AND2_X1 U9156 ( .A1(n7232), .A2(n6609), .ZN(n6717) );
  AND2_X1 U9157 ( .A1(n6933), .A2(n6619), .ZN(n6718) );
  OR2_X1 U9158 ( .A1(n14708), .A2(n6995), .ZN(n6719) );
  AND2_X1 U9159 ( .A1(n6908), .A2(n6907), .ZN(n11393) );
  INV_X1 U9160 ( .A(n12529), .ZN(n15181) );
  NAND2_X1 U9161 ( .A1(n6993), .A2(n6994), .ZN(n11579) );
  INV_X1 U9162 ( .A(n11579), .ZN(n6992) );
  NAND2_X1 U9163 ( .A1(n10995), .A2(n10994), .ZN(n10996) );
  AND2_X1 U9164 ( .A1(n11613), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6720) );
  AND2_X1 U9165 ( .A1(n11229), .A2(n9324), .ZN(n6721) );
  INV_X1 U9166 ( .A(n8906), .ZN(n6856) );
  INV_X1 U9167 ( .A(n15395), .ZN(n15392) );
  NAND2_X1 U9168 ( .A1(n10756), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14554) );
  INV_X1 U9169 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n6778) );
  OR2_X1 U9170 ( .A1(n14372), .A2(n12557), .ZN(n6722) );
  AND2_X1 U9171 ( .A1(n14744), .A2(n11091), .ZN(n6723) );
  INV_X1 U9172 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7027) );
  OR2_X1 U9173 ( .A1(n11181), .A2(n11180), .ZN(n6724) );
  INV_X1 U9174 ( .A(n11038), .ZN(n7086) );
  NAND2_X1 U9175 ( .A1(n13486), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6725) );
  INV_X1 U9176 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n6852) );
  INV_X1 U9177 ( .A(n10546), .ZN(n6765) );
  AND2_X1 U9178 ( .A1(n8655), .A2(P2_U3088), .ZN(n6726) );
  AND2_X1 U9179 ( .A1(n8655), .A2(P3_U3151), .ZN(n6727) );
  XOR2_X1 U9180 ( .A(n12608), .B(P3_REG1_REG_19__SCAN_IN), .Z(n6728) );
  INV_X1 U9181 ( .A(n7555), .ZN(n11875) );
  XOR2_X1 U9182 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n6729) );
  INV_X1 U9183 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6842) );
  INV_X1 U9184 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9223) );
  NAND2_X1 U9185 ( .A1(n15204), .A2(n15203), .ZN(n15202) );
  NAND2_X1 U9186 ( .A1(n15223), .A2(n12586), .ZN(n12587) );
  AOI21_X1 U9187 ( .B1(n15120), .B2(n15123), .A(n15119), .ZN(n15146) );
  NOR2_X1 U9188 ( .A1(n14394), .A2(n14395), .ZN(n14393) );
  AOI21_X1 U9189 ( .B1(n12588), .B2(n12554), .A(n14360), .ZN(n14383) );
  XNOR2_X1 U9190 ( .A(n12597), .B(n12598), .ZN(n14410) );
  NAND2_X4 U9191 ( .A1(n9222), .A2(n6734), .ZN(n12589) );
  NAND2_X1 U9192 ( .A1(n8166), .A2(n8165), .ZN(n11483) );
  NAND2_X1 U9193 ( .A1(n11027), .A2(n11026), .ZN(n11029) );
  NAND2_X1 U9194 ( .A1(n10862), .A2(n10866), .ZN(n10861) );
  OAI211_X2 U9195 ( .C1(n8032), .C2(n10007), .A(n7602), .B(n7601), .ZN(n11082)
         );
  NAND2_X1 U9196 ( .A1(n10457), .A2(n10456), .ZN(n10455) );
  OR2_X1 U9198 ( .A1(n10167), .A2(n14879), .ZN(n7602) );
  NAND2_X1 U9199 ( .A1(n7110), .A2(n8138), .ZN(n7565) );
  NAND2_X1 U9200 ( .A1(n7051), .A2(n8009), .ZN(n7050) );
  INV_X1 U9201 ( .A(n11909), .ZN(n11956) );
  NAND2_X1 U9202 ( .A1(n7297), .A2(n7292), .ZN(n7291) );
  NAND2_X1 U9203 ( .A1(n7032), .A2(n6737), .ZN(n7031) );
  NAND2_X1 U9204 ( .A1(n6752), .A2(n7413), .ZN(n7032) );
  NAND2_X1 U9205 ( .A1(n10968), .A2(n9905), .ZN(n11064) );
  NAND2_X1 U9206 ( .A1(n13007), .A2(n13009), .ZN(n13008) );
  NAND2_X1 U9207 ( .A1(n12113), .A2(n12112), .ZN(n12966) );
  NAND2_X1 U9208 ( .A1(n12994), .A2(n12993), .ZN(n12992) );
  NAND2_X1 U9209 ( .A1(n6744), .A2(n9895), .ZN(n10809) );
  INV_X1 U9210 ( .A(n7943), .ZN(n6738) );
  NAND2_X1 U9211 ( .A1(n10525), .A2(n6687), .ZN(n6744) );
  NAND2_X1 U9212 ( .A1(n13018), .A2(n9883), .ZN(n10526) );
  NAND3_X1 U9213 ( .A1(n7672), .A2(n6739), .A3(n6738), .ZN(n8141) );
  NOR2_X1 U9214 ( .A1(n11823), .A2(n11824), .ZN(n11822) );
  NAND2_X1 U9215 ( .A1(n7139), .A2(n7138), .ZN(n12790) );
  AOI21_X1 U9216 ( .B1(n15366), .B2(n12622), .A(n12617), .ZN(n9830) );
  NOR2_X1 U9217 ( .A1(n14351), .A2(n14352), .ZN(n14350) );
  NAND2_X1 U9218 ( .A1(n7225), .A2(n7224), .ZN(n7223) );
  NAND2_X1 U9219 ( .A1(n7234), .A2(n7233), .ZN(n10671) );
  NOR2_X1 U9220 ( .A1(n14388), .A2(n14389), .ZN(n14387) );
  NAND2_X1 U9221 ( .A1(n6766), .A2(n6620), .ZN(n10540) );
  AOI21_X1 U9222 ( .B1(n7237), .B2(P3_REG2_REG_3__SCAN_IN), .A(n10541), .ZN(
        n10723) );
  AOI21_X1 U9223 ( .B1(n7240), .B2(n7239), .A(n7238), .ZN(n12546) );
  NOR2_X1 U9224 ( .A1(n15173), .A2(n6749), .ZN(n12553) );
  NOR2_X1 U9225 ( .A1(n12551), .A2(n15157), .ZN(n15175) );
  NAND2_X1 U9226 ( .A1(n7296), .A2(n7299), .ZN(n11950) );
  NAND2_X1 U9227 ( .A1(n7262), .A2(n6683), .ZN(n14162) );
  OAI21_X2 U9228 ( .B1(n11921), .B2(n7304), .A(n7302), .ZN(n14104) );
  OAI21_X1 U9229 ( .B1(n14042), .B2(n14041), .A(n11932), .ZN(n14026) );
  NAND2_X1 U9230 ( .A1(n14729), .A2(n10800), .ZN(n10801) );
  OAI21_X1 U9231 ( .B1(n14697), .B2(n14698), .A(n11316), .ZN(n11317) );
  AOI21_X2 U9232 ( .B1(n6742), .B2(n14738), .A(n11953), .ZN(n14205) );
  NAND2_X1 U9233 ( .A1(n11949), .A2(n11950), .ZN(n6742) );
  NAND2_X2 U9234 ( .A1(n14025), .A2(n11933), .ZN(n14008) );
  NAND2_X1 U9235 ( .A1(n14715), .A2(n11094), .ZN(n7301) );
  AND2_X2 U9236 ( .A1(n7604), .A2(n7603), .ZN(n11076) );
  AND2_X2 U9237 ( .A1(n13181), .A2(n13180), .ZN(n13182) );
  OAI211_X1 U9238 ( .C1(n13440), .C2(n11883), .A(n11887), .B(n8202), .ZN(
        n13377) );
  AOI21_X1 U9239 ( .B1(n7401), .B2(n6595), .A(n7400), .ZN(n11558) );
  NAND3_X1 U9240 ( .A1(n6884), .A2(n6885), .A3(n7666), .ZN(n7670) );
  INV_X1 U9241 ( .A(n8141), .ZN(n8133) );
  NAND2_X1 U9242 ( .A1(n10638), .A2(n7530), .ZN(n10616) );
  INV_X1 U9243 ( .A(n7225), .ZN(n14415) );
  OAI21_X1 U9244 ( .B1(n9227), .B2(n6748), .A(n6747), .ZN(n6746) );
  INV_X1 U9245 ( .A(n10541), .ZN(n6766) );
  INV_X1 U9246 ( .A(n10540), .ZN(n7237) );
  NAND4_X1 U9247 ( .A1(n14416), .A2(n14418), .A3(n14417), .A4(n14419), .ZN(
        P3_U3200) );
  OAI21_X1 U9248 ( .B1(n10723), .B2(n10722), .A(n7236), .ZN(n7235) );
  OAI21_X1 U9249 ( .B1(n10705), .B2(n9343), .A(n6676), .ZN(n7240) );
  NAND2_X1 U9250 ( .A1(n6890), .A2(n7796), .ZN(n7814) );
  INV_X1 U9251 ( .A(n7047), .ZN(n7046) );
  NAND2_X1 U9252 ( .A1(n7263), .A2(n7265), .ZN(n7262) );
  NAND2_X1 U9253 ( .A1(n6881), .A2(n6883), .ZN(n6878) );
  NAND2_X1 U9254 ( .A1(n6644), .A2(n7630), .ZN(n6885) );
  OAI21_X1 U9255 ( .B1(n7730), .B2(n7048), .A(n7751), .ZN(n7047) );
  NAND2_X1 U9256 ( .A1(n7941), .A2(n7940), .ZN(n7960) );
  NAND2_X1 U9257 ( .A1(n7050), .A2(n7052), .ZN(n8025) );
  INV_X2 U9258 ( .A(n7596), .ZN(n10005) );
  NAND2_X1 U9259 ( .A1(n7816), .A2(n7038), .ZN(n7037) );
  NAND2_X1 U9260 ( .A1(n7037), .A2(n7035), .ZN(n7876) );
  OAI21_X1 U9261 ( .B1(n11935), .B2(n7297), .A(n7291), .ZN(n7290) );
  OR2_X2 U9262 ( .A1(n7555), .A2(n11865), .ZN(n7608) );
  NAND2_X1 U9263 ( .A1(n8173), .A2(n8172), .ZN(n14463) );
  NAND2_X1 U9264 ( .A1(n13315), .A2(n8180), .ZN(n8182) );
  NAND2_X1 U9265 ( .A1(n13328), .A2(n13332), .ZN(n13330) );
  NAND2_X1 U9266 ( .A1(n13442), .A2(n8177), .ZN(n13362) );
  AOI21_X1 U9267 ( .B1(n11749), .B2(n11750), .A(n8176), .ZN(n11773) );
  INV_X1 U9268 ( .A(n13245), .ZN(n6752) );
  NOR2_X2 U9269 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7546) );
  INV_X1 U9270 ( .A(n9992), .ZN(n7404) );
  NAND2_X1 U9271 ( .A1(n6877), .A2(n9223), .ZN(n7581) );
  NAND2_X2 U9272 ( .A1(n11361), .A2(n9923), .ZN(n11380) );
  NAND2_X1 U9273 ( .A1(n7352), .A2(n7351), .ZN(n9877) );
  NOR2_X2 U9274 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7544) );
  NOR2_X2 U9275 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7545) );
  NAND2_X1 U9276 ( .A1(n9993), .A2(n7584), .ZN(n11075) );
  INV_X1 U9277 ( .A(n11212), .ZN(n6754) );
  OAI21_X2 U9278 ( .B1(n11765), .B2(n7889), .A(n7890), .ZN(n13350) );
  OAI21_X2 U9279 ( .B1(n13287), .B2(n7993), .A(n7992), .ZN(n13270) );
  OAI21_X2 U9280 ( .B1(n11484), .B2(n7071), .A(n7068), .ZN(n14454) );
  INV_X2 U9281 ( .A(n7573), .ZN(n10595) );
  NAND2_X1 U9282 ( .A1(n7078), .A2(n7572), .ZN(n7573) );
  AOI21_X2 U9283 ( .B1(n8154), .B2(n14456), .A(n8153), .ZN(n11887) );
  XNOR2_X1 U9284 ( .A(n15086), .B(n13083), .ZN(n11026) );
  NAND2_X2 U9285 ( .A1(n7637), .A2(n7636), .ZN(n13022) );
  NAND2_X1 U9286 ( .A1(n11030), .A2(n7646), .ZN(n10902) );
  INV_X1 U9287 ( .A(n11486), .ZN(n7792) );
  NAND2_X1 U9288 ( .A1(n11032), .A2(n11031), .ZN(n11030) );
  NAND2_X1 U9289 ( .A1(n8155), .A2(n10407), .ZN(n9156) );
  NAND2_X1 U9290 ( .A1(n7494), .A2(n12161), .ZN(n12217) );
  NAND2_X1 U9291 ( .A1(n12210), .A2(n12152), .ZN(n12155) );
  INV_X1 U9292 ( .A(n9790), .ZN(n11504) );
  INV_X1 U9293 ( .A(n11710), .ZN(n6862) );
  INV_X1 U9294 ( .A(n11813), .ZN(n6860) );
  INV_X1 U9295 ( .A(n12242), .ZN(n7483) );
  NAND3_X1 U9296 ( .A1(n6759), .A2(n6757), .A3(n6756), .ZN(P2_U3233) );
  NAND2_X1 U9297 ( .A1(n11380), .A2(n6681), .ZN(n6760) );
  INV_X4 U9298 ( .A(n10005), .ZN(n7076) );
  NAND2_X1 U9299 ( .A1(n13283), .A2(n8187), .ZN(n13255) );
  NAND2_X1 U9300 ( .A1(n13179), .A2(n8194), .ZN(n8196) );
  NAND2_X1 U9301 ( .A1(n7405), .A2(n7404), .ZN(n9990) );
  NAND2_X1 U9302 ( .A1(n9859), .A2(n10595), .ZN(n7574) );
  INV_X1 U9303 ( .A(n6761), .ZN(n11886) );
  OAI21_X1 U9304 ( .B1(n11883), .B2(n13365), .A(n6762), .ZN(n6761) );
  NAND2_X1 U9305 ( .A1(n9990), .A2(n8157), .ZN(n11073) );
  INV_X1 U9306 ( .A(n7109), .ZN(n7552) );
  NAND2_X1 U9307 ( .A1(n9762), .A2(n12405), .ZN(n12809) );
  XNOR2_X1 U9308 ( .A(n7223), .B(n7222), .ZN(n12562) );
  INV_X1 U9309 ( .A(n7235), .ZN(n10542) );
  OAI21_X1 U9310 ( .B1(n14350), .B2(n7220), .A(n7219), .ZN(n12558) );
  AND2_X4 U9311 ( .A1(n9226), .A2(n7076), .ZN(n12318) );
  NAND2_X1 U9312 ( .A1(n13270), .A2(n13280), .ZN(n7084) );
  NAND2_X1 U9313 ( .A1(n7872), .A2(n7871), .ZN(n11765) );
  NAND2_X1 U9314 ( .A1(n7056), .A2(n7055), .ZN(n13287) );
  INV_X1 U9315 ( .A(n13350), .ZN(n7913) );
  NAND2_X1 U9316 ( .A1(n9269), .A2(n9268), .ZN(n6770) );
  NAND2_X1 U9317 ( .A1(n9225), .A2(n9224), .ZN(n9253) );
  NAND2_X1 U9318 ( .A1(n9718), .A2(n9717), .ZN(n6777) );
  INV_X1 U9319 ( .A(n6779), .ZN(n9616) );
  NAND2_X1 U9320 ( .A1(n9516), .A2(n6791), .ZN(n6790) );
  NAND3_X1 U9321 ( .A1(n6800), .A2(n7193), .A3(n6799), .ZN(n6798) );
  NAND2_X1 U9322 ( .A1(n7323), .A2(n6805), .ZN(n6801) );
  NAND3_X1 U9323 ( .A1(n12469), .A2(n12464), .A3(n6807), .ZN(n7202) );
  NAND2_X1 U9324 ( .A1(n14699), .A2(n14698), .ZN(n6808) );
  NAND2_X1 U9325 ( .A1(n11327), .A2(n11326), .ZN(n6809) );
  NAND2_X1 U9326 ( .A1(n11264), .A2(n11272), .ZN(n11112) );
  NAND2_X1 U9327 ( .A1(n7376), .A2(n11117), .ZN(n6810) );
  NAND3_X1 U9328 ( .A1(n8835), .A2(n14650), .A3(n14649), .ZN(n6813) );
  NAND2_X1 U9329 ( .A1(n11415), .A2(n6816), .ZN(n6814) );
  NAND2_X1 U9330 ( .A1(n6677), .A2(n6814), .ZN(n11685) );
  NAND2_X1 U9331 ( .A1(n11415), .A2(n11414), .ZN(n11534) );
  NAND2_X1 U9332 ( .A1(n11688), .A2(n6826), .ZN(n6824) );
  INV_X1 U9333 ( .A(n7391), .ZN(n6831) );
  AND4_X2 U9334 ( .A1(n8258), .A2(n8257), .A3(n8352), .A4(n6665), .ZN(n8272)
         );
  OAI21_X1 U9335 ( .B1(n15398), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6675), .ZN(
        n6845) );
  XNOR2_X1 U9336 ( .A(n8898), .B(n8899), .ZN(n15398) );
  NAND2_X1 U9337 ( .A1(n6848), .A2(n8908), .ZN(n6855) );
  NAND2_X1 U9338 ( .A1(n8907), .A2(n8906), .ZN(n6848) );
  AOI21_X1 U9339 ( .B1(n6856), .B2(n8908), .A(P2_ADDR_REG_8__SCAN_IN), .ZN(
        n6849) );
  INV_X1 U9340 ( .A(n8908), .ZN(n6850) );
  NAND2_X1 U9341 ( .A1(n12190), .A2(n6869), .ZN(n6866) );
  NAND2_X1 U9342 ( .A1(n6866), .A2(n6867), .ZN(n12210) );
  NAND2_X1 U9343 ( .A1(n9482), .A2(n6604), .ZN(n9570) );
  NAND2_X1 U9344 ( .A1(n9572), .A2(n6621), .ZN(n9736) );
  NAND2_X1 U9345 ( .A1(n9572), .A2(n6702), .ZN(n6876) );
  NAND2_X1 U9346 ( .A1(n9572), .A2(n9571), .ZN(n9730) );
  INV_X1 U9347 ( .A(n6876), .ZN(n9733) );
  NAND2_X1 U9348 ( .A1(n7076), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7077) );
  NAND2_X1 U9349 ( .A1(n7076), .A2(SI_0_), .ZN(n8316) );
  NOR2_X1 U9350 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8655), .ZN(n14325) );
  NAND2_X1 U9351 ( .A1(n8655), .A2(SI_0_), .ZN(n6877) );
  MUX2_X1 U9352 ( .A(n10893), .B(n13735), .S(n8655), .Z(n7894) );
  MUX2_X1 U9353 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n8655), .Z(n7974) );
  MUX2_X1 U9354 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n8655), .Z(n7961) );
  MUX2_X1 U9355 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n8655), .Z(n7979) );
  MUX2_X1 U9356 ( .A(n11132), .B(n11135), .S(n8655), .Z(n7935) );
  MUX2_X1 U9357 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n8655), .Z(n8010) );
  MUX2_X1 U9358 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n8655), .Z(n8009) );
  MUX2_X1 U9359 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n8655), .Z(n8058) );
  MUX2_X1 U9360 ( .A(n14299), .B(n9688), .S(n8655), .Z(n8078) );
  MUX2_X1 U9361 ( .A(n14296), .B(n13486), .S(n8655), .Z(n8094) );
  MUX2_X1 U9362 ( .A(n11877), .B(n9719), .S(n8655), .Z(n8096) );
  MUX2_X1 U9363 ( .A(n6778), .B(n11867), .S(n8655), .Z(n8243) );
  MUX2_X1 U9364 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8655), .Z(n8246) );
  MUX2_X1 U9365 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8655), .Z(n8248) );
  AND2_X1 U9366 ( .A1(P2_U3088), .A2(n7076), .ZN(n13769) );
  NAND2_X1 U9367 ( .A1(n10064), .A2(n7076), .ZN(n8683) );
  NAND2_X1 U9368 ( .A1(n7713), .A2(n6881), .ZN(n6879) );
  NAND2_X1 U9369 ( .A1(n7653), .A2(n7656), .ZN(n6884) );
  INV_X1 U9370 ( .A(n7653), .ZN(n6887) );
  NAND2_X1 U9371 ( .A1(n7630), .A2(n7629), .ZN(n7654) );
  NAND2_X1 U9372 ( .A1(n6887), .A2(n7654), .ZN(n6886) );
  NAND2_X1 U9373 ( .A1(n14445), .A2(n9941), .ZN(n9943) );
  NAND2_X1 U9374 ( .A1(n7774), .A2(n6891), .ZN(n6888) );
  NAND2_X1 U9375 ( .A1(n6888), .A2(n6889), .ZN(n7834) );
  NAND2_X1 U9376 ( .A1(n7774), .A2(n6894), .ZN(n6890) );
  NAND2_X1 U9377 ( .A1(n7774), .A2(n7773), .ZN(n7795) );
  NAND2_X1 U9378 ( .A1(n14515), .A2(n14516), .ZN(n12009) );
  NAND2_X1 U9379 ( .A1(n6901), .A2(n6900), .ZN(n14515) );
  NAND2_X1 U9380 ( .A1(n14542), .A2(n7496), .ZN(n6900) );
  NAND2_X1 U9381 ( .A1(n11254), .A2(n6603), .ZN(n6904) );
  NAND2_X1 U9382 ( .A1(n13870), .A2(n13869), .ZN(n13868) );
  NAND2_X1 U9383 ( .A1(n13814), .A2(n7501), .ZN(n6915) );
  OAI211_X1 U9384 ( .C1(n13814), .C2(n6913), .A(n6910), .B(n6909), .ZN(n12089)
         );
  NAND2_X1 U9385 ( .A1(n13814), .A2(n6674), .ZN(n6909) );
  NAND2_X1 U9386 ( .A1(n6914), .A2(n6679), .ZN(n6911) );
  OR2_X1 U9387 ( .A1(n6914), .A2(n6920), .ZN(n6912) );
  INV_X1 U9388 ( .A(n10503), .ZN(n6921) );
  NAND2_X1 U9389 ( .A1(n6924), .A2(n6922), .ZN(n11169) );
  NOR2_X1 U9390 ( .A1(n10761), .A2(n7529), .ZN(n10767) );
  NAND2_X1 U9391 ( .A1(n11639), .A2(n6928), .ZN(n6927) );
  NAND2_X1 U9392 ( .A1(n8270), .A2(n6941), .ZN(n8825) );
  NAND2_X1 U9393 ( .A1(n8270), .A2(n6682), .ZN(n6939) );
  NAND2_X1 U9394 ( .A1(n6946), .A2(n6949), .ZN(n8710) );
  NAND3_X1 U9395 ( .A1(n8682), .A2(n6947), .A3(n8681), .ZN(n6946) );
  INV_X1 U9396 ( .A(n8653), .ZN(n8650) );
  NAND2_X1 U9397 ( .A1(n6955), .A2(n6956), .ZN(n8622) );
  NAND2_X1 U9398 ( .A1(n8569), .A2(n6958), .ZN(n6955) );
  NOR2_X1 U9399 ( .A1(n6961), .A2(n6960), .ZN(n8500) );
  NOR2_X1 U9400 ( .A1(n7242), .A2(n8483), .ZN(n6972) );
  NAND2_X1 U9401 ( .A1(n6973), .A2(n6974), .ZN(n7243) );
  NAND2_X1 U9402 ( .A1(n7249), .A2(n6680), .ZN(n6973) );
  OR2_X1 U9403 ( .A1(n8517), .A2(n6986), .ZN(n6983) );
  NAND2_X1 U9404 ( .A1(n8517), .A2(n6981), .ZN(n6980) );
  NAND3_X1 U9405 ( .A1(n8835), .A2(n14650), .A3(n13904), .ZN(n8307) );
  NAND3_X1 U9406 ( .A1(n6605), .A2(n7025), .A3(n6705), .ZN(n7024) );
  NAND4_X1 U9407 ( .A1(n7029), .A2(n7028), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7442) );
  NAND2_X1 U9408 ( .A1(n7031), .A2(n7034), .ZN(n13207) );
  INV_X1 U9409 ( .A(n13207), .ZN(n7033) );
  NAND2_X1 U9410 ( .A1(n7996), .A2(SI_22_), .ZN(n7052) );
  XNOR2_X1 U9411 ( .A(n7628), .B(SI_3_), .ZN(n7625) );
  OAI21_X1 U9412 ( .B1(n10005), .B2(n7054), .A(n7053), .ZN(n7628) );
  NAND2_X1 U9413 ( .A1(n10005), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7053) );
  NAND2_X1 U9414 ( .A1(n10902), .A2(n7661), .ZN(n7664) );
  NAND2_X1 U9415 ( .A1(n10582), .A2(n7624), .ZN(n11032) );
  NAND2_X1 U9416 ( .A1(n13318), .A2(n7058), .ZN(n7056) );
  NAND2_X1 U9417 ( .A1(n13240), .A2(n7065), .ZN(n7062) );
  NAND2_X1 U9418 ( .A1(n7062), .A2(n7063), .ZN(n13210) );
  NAND3_X1 U9419 ( .A1(n7074), .A2(n10167), .A3(n7075), .ZN(n7078) );
  NAND2_X1 U9420 ( .A1(n10009), .A2(n7077), .ZN(n7074) );
  NAND2_X1 U9421 ( .A1(n7084), .A2(n7083), .ZN(n8020) );
  OAI21_X2 U9422 ( .B1(n11344), .B2(n7767), .A(n7768), .ZN(n11486) );
  NAND2_X1 U9423 ( .A1(n11769), .A2(n7090), .ZN(n7093) );
  NAND2_X1 U9424 ( .A1(n11352), .A2(n6686), .ZN(n7096) );
  AND3_X2 U9425 ( .A1(n7373), .A2(n7372), .A3(n7634), .ZN(n8138) );
  NAND2_X1 U9426 ( .A1(n7111), .A2(n7112), .ZN(n9030) );
  NAND3_X1 U9427 ( .A1(n9025), .A2(n6700), .A3(n9024), .ZN(n7111) );
  NAND2_X1 U9428 ( .A1(n7113), .A2(n7114), .ZN(n8999) );
  NAND3_X1 U9429 ( .A1(n8993), .A2(n6695), .A3(n8992), .ZN(n7113) );
  NAND2_X1 U9430 ( .A1(n7115), .A2(n7116), .ZN(n9009) );
  NAND3_X1 U9431 ( .A1(n9004), .A2(n6696), .A3(n9003), .ZN(n7115) );
  NAND3_X1 U9432 ( .A1(n9051), .A2(n9050), .A3(n6692), .ZN(n7118) );
  NAND2_X1 U9433 ( .A1(n7118), .A2(n7119), .ZN(n9057) );
  NAND2_X1 U9434 ( .A1(n7120), .A2(n7121), .ZN(n9075) );
  NAND3_X1 U9435 ( .A1(n9070), .A2(n6701), .A3(n9069), .ZN(n7120) );
  NAND3_X1 U9436 ( .A1(n8983), .A2(n8982), .A3(n6693), .ZN(n7123) );
  NAND2_X1 U9437 ( .A1(n7123), .A2(n7124), .ZN(n8988) );
  NAND2_X1 U9438 ( .A1(n7126), .A2(n7127), .ZN(n9020) );
  NAND3_X1 U9439 ( .A1(n9014), .A2(n6699), .A3(n9013), .ZN(n7126) );
  NAND2_X1 U9440 ( .A1(n7128), .A2(n7129), .ZN(n9094) );
  NAND3_X1 U9441 ( .A1(n9088), .A2(n6694), .A3(n9087), .ZN(n7128) );
  NAND2_X1 U9442 ( .A1(n7130), .A2(n7132), .ZN(n8962) );
  NAND3_X1 U9443 ( .A1(n8956), .A2(n7131), .A3(n8955), .ZN(n7130) );
  OR2_X1 U9444 ( .A1(n8957), .A2(n8959), .ZN(n7131) );
  NAND2_X1 U9445 ( .A1(n8957), .A2(n8959), .ZN(n7132) );
  INV_X1 U9446 ( .A(n7133), .ZN(n12337) );
  NAND2_X2 U9447 ( .A1(n12341), .A2(n7133), .ZN(n12823) );
  NAND2_X1 U9448 ( .A1(n12822), .A2(n7133), .ZN(n10825) );
  NAND2_X1 U9449 ( .A1(n14421), .A2(n9457), .ZN(n7134) );
  NAND2_X1 U9450 ( .A1(n9596), .A2(n6691), .ZN(n12726) );
  NAND2_X1 U9451 ( .A1(n11740), .A2(n7140), .ZN(n7139) );
  NAND2_X1 U9452 ( .A1(n9685), .A2(n7143), .ZN(n12635) );
  INV_X1 U9453 ( .A(n9376), .ZN(n11475) );
  NAND2_X1 U9454 ( .A1(n7144), .A2(n7145), .ZN(n9418) );
  NAND2_X1 U9455 ( .A1(n9376), .A2(n9401), .ZN(n7144) );
  NAND2_X1 U9456 ( .A1(n9259), .A2(n15309), .ZN(n15315) );
  NOR2_X2 U9457 ( .A1(n7158), .A2(n9208), .ZN(n9482) );
  NAND3_X1 U9458 ( .A1(n7159), .A2(n9254), .A3(n9464), .ZN(n7158) );
  AND3_X2 U9459 ( .A1(n7161), .A2(n7461), .A3(n9214), .ZN(n9784) );
  NAND2_X1 U9460 ( .A1(n12700), .A2(n7170), .ZN(n12699) );
  AOI21_X2 U9461 ( .B1(n13194), .B2(n13206), .A(n8091), .ZN(n13181) );
  NAND2_X1 U9462 ( .A1(n12823), .A2(n12816), .ZN(n15318) );
  NAND2_X1 U9463 ( .A1(n11074), .A2(n7604), .ZN(n10584) );
  OAI21_X2 U9464 ( .B1(n10983), .B2(n10980), .A(n7710), .ZN(n11048) );
  NOR2_X2 U9465 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n7548) );
  NAND2_X4 U9466 ( .A1(n7162), .A2(n12959), .ZN(n9304) );
  INV_X1 U9467 ( .A(n15309), .ZN(n15317) );
  NAND2_X1 U9468 ( .A1(n12345), .A2(n12344), .ZN(n15309) );
  NAND2_X1 U9469 ( .A1(n15317), .A2(n15308), .ZN(n9749) );
  NAND2_X1 U9470 ( .A1(n12719), .A2(n7165), .ZN(n7164) );
  NAND2_X1 U9471 ( .A1(n7164), .A2(n7167), .ZN(n12680) );
  NAND2_X1 U9472 ( .A1(n7174), .A2(n7172), .ZN(n9762) );
  NAND2_X1 U9473 ( .A1(n9836), .A2(n12453), .ZN(n12311) );
  INV_X1 U9474 ( .A(n7232), .ZN(n15192) );
  NAND2_X1 U9475 ( .A1(n8500), .A2(n8501), .ZN(n8499) );
  NAND2_X1 U9476 ( .A1(n7243), .A2(n7246), .ZN(n8785) );
  NAND2_X1 U9477 ( .A1(n8723), .A2(n7250), .ZN(n7249) );
  INV_X1 U9478 ( .A(n8722), .ZN(n7253) );
  NAND2_X1 U9479 ( .A1(n8654), .A2(n6703), .ZN(n7255) );
  OAI21_X1 U9480 ( .B1(n6636), .B2(n7255), .A(n7256), .ZN(n8680) );
  OR2_X1 U9481 ( .A1(n8669), .A2(n7424), .ZN(n7256) );
  OAI22_X1 U9482 ( .A1(n8433), .A2(n7259), .B1(n7258), .B2(n8434), .ZN(n7260)
         );
  NAND2_X1 U9483 ( .A1(n7260), .A2(n8453), .ZN(n8456) );
  INV_X2 U9484 ( .A(n8544), .ZN(n8775) );
  MUX2_X1 U9485 ( .A(n8341), .B(n8342), .S(n8544), .Z(n8343) );
  NAND2_X2 U9486 ( .A1(n10798), .A2(n8340), .ZN(n10936) );
  INV_X1 U9487 ( .A(n14563), .ZN(n7263) );
  NAND2_X1 U9488 ( .A1(n11271), .A2(n7272), .ZN(n7270) );
  NAND2_X1 U9489 ( .A1(n11410), .A2(n7280), .ZN(n7279) );
  OR2_X1 U9490 ( .A1(n14008), .A2(n11948), .ZN(n7296) );
  OAI211_X1 U9491 ( .C1(n14008), .C2(n7294), .A(n7290), .B(n7288), .ZN(n14200)
         );
  NAND2_X1 U9492 ( .A1(n14008), .A2(n7289), .ZN(n7288) );
  NAND2_X1 U9493 ( .A1(n7301), .A2(n6678), .ZN(n11121) );
  INV_X1 U9494 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7319) );
  NAND2_X1 U9495 ( .A1(n9390), .A2(n7327), .ZN(n7324) );
  NAND2_X1 U9496 ( .A1(n7324), .A2(n7325), .ZN(n9422) );
  NAND2_X1 U9497 ( .A1(n9616), .A2(n7334), .ZN(n7331) );
  NAND2_X1 U9498 ( .A1(n7331), .A2(n7332), .ZN(n9643) );
  INV_X1 U9499 ( .A(n9877), .ZN(n10519) );
  NAND2_X1 U9500 ( .A1(n7354), .A2(n9870), .ZN(n7351) );
  NAND2_X1 U9501 ( .A1(n7353), .A2(n10455), .ZN(n7352) );
  AND2_X1 U9502 ( .A1(n9870), .A2(n9869), .ZN(n10449) );
  NAND2_X1 U9503 ( .A1(n10455), .A2(n9863), .ZN(n10448) );
  OAI21_X1 U9504 ( .B1(n11846), .B2(n7358), .A(n7357), .ZN(n12985) );
  NOR2_X1 U9505 ( .A1(n11844), .A2(n9952), .ZN(n13042) );
  NAND2_X1 U9506 ( .A1(n7365), .A2(n7364), .ZN(n11361) );
  NAND2_X1 U9507 ( .A1(n11063), .A2(n9911), .ZN(n11151) );
  AND2_X1 U9508 ( .A1(n12999), .A2(n13000), .ZN(n13005) );
  OR2_X2 U9509 ( .A1(n12999), .A2(n7370), .ZN(n7369) );
  INV_X1 U9510 ( .A(n7942), .ZN(n7372) );
  AND3_X1 U9511 ( .A1(n7544), .A2(n7545), .A3(n7546), .ZN(n7800) );
  XNOR2_X1 U9512 ( .A(n7376), .B(n11117), .ZN(n14806) );
  OAI211_X1 U9513 ( .C1(n10952), .C2(n7378), .A(n10936), .B(n7377), .ZN(n10784) );
  NAND3_X1 U9514 ( .A1(n10796), .A2(n10782), .A3(n10794), .ZN(n7377) );
  INV_X1 U9515 ( .A(n10782), .ZN(n7378) );
  NAND2_X1 U9516 ( .A1(n14090), .A2(n6690), .ZN(n14075) );
  AND3_X2 U9517 ( .A1(n8307), .A2(n7395), .A3(n8308), .ZN(n14770) );
  NAND2_X1 U9518 ( .A1(n8272), .A2(n7519), .ZN(n8828) );
  INV_X1 U9519 ( .A(n11483), .ZN(n7401) );
  NAND2_X1 U9520 ( .A1(n7534), .A2(n7408), .ZN(n7406) );
  NAND2_X1 U9521 ( .A1(n7406), .A2(n7407), .ZN(n11342) );
  NAND2_X1 U9522 ( .A1(n8138), .A2(n7550), .ZN(n7566) );
  NAND2_X1 U9523 ( .A1(n7436), .A2(n7437), .ZN(n7996) );
  NAND4_X1 U9524 ( .A1(n7446), .A2(n7445), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n13724), .ZN(n7443) );
  OAI22_X1 U9525 ( .A1(n8710), .A2(n7447), .B1(n8711), .B2(n7448), .ZN(n8723)
         );
  OAI211_X1 U9526 ( .C1(n7449), .C2(n12816), .A(n10880), .B(n10879), .ZN(
        n10881) );
  NAND2_X1 U9527 ( .A1(n10829), .A2(n7449), .ZN(n10880) );
  NAND2_X1 U9528 ( .A1(n11303), .A2(n7457), .ZN(n7455) );
  NAND2_X1 U9529 ( .A1(n7462), .A2(n7460), .ZN(n9446) );
  INV_X1 U9530 ( .A(n9315), .ZN(n7460) );
  OAI21_X1 U9531 ( .B1(n11813), .B2(n11812), .A(n11811), .ZN(n12128) );
  NAND2_X1 U9532 ( .A1(n9784), .A2(n9215), .ZN(n9781) );
  NAND2_X1 U9533 ( .A1(n12263), .A2(n12731), .ZN(n7489) );
  NAND2_X1 U9534 ( .A1(n7478), .A2(n7477), .ZN(n12199) );
  AND2_X1 U9535 ( .A1(n7489), .A2(n7495), .ZN(n12242) );
  INV_X1 U9536 ( .A(n12156), .ZN(n7495) );
  NAND2_X1 U9537 ( .A1(n13851), .A2(n7506), .ZN(n7505) );
  OAI21_X2 U9538 ( .B1(n11401), .B2(n7518), .A(n7514), .ZN(n11639) );
  NAND2_X1 U9539 ( .A1(n8285), .A2(n7520), .ZN(n14287) );
  NAND2_X1 U9540 ( .A1(n9768), .A2(n12328), .ZN(n12650) );
  NAND2_X1 U9541 ( .A1(n8978), .A2(n8977), .ZN(n8974) );
  MUX2_X1 U9542 ( .A(n14273), .B(P1_REG1_REG_27__SCAN_IN), .S(n14856), .Z(
        P1_U3555) );
  MUX2_X1 U9543 ( .A(n14273), .B(P1_REG0_REG_27__SCAN_IN), .S(n14842), .Z(
        P1_U3523) );
  INV_X1 U9544 ( .A(n8970), .ZN(n8973) );
  CLKBUF_X1 U9545 ( .A(n11227), .Z(n11228) );
  NAND2_X1 U9546 ( .A1(n11725), .A2(n11711), .ZN(n11714) );
  INV_X1 U9547 ( .A(n9248), .ZN(n10491) );
  AND4_X2 U9548 ( .A1(n9240), .A2(n9239), .A3(n9238), .A4(n9237), .ZN(n9248)
         );
  CLKBUF_X1 U9549 ( .A(n9157), .Z(n9994) );
  OR2_X1 U9550 ( .A1(n7606), .A2(n7585), .ZN(n7587) );
  OR2_X1 U9551 ( .A1(n7606), .A2(n7575), .ZN(n7579) );
  OR2_X1 U9552 ( .A1(n7606), .A2(n7556), .ZN(n7560) );
  NAND2_X1 U9553 ( .A1(n7565), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7564) );
  CLKBUF_X1 U9554 ( .A(n11843), .Z(n11846) );
  NAND2_X1 U9555 ( .A1(n12978), .A2(n12977), .ZN(n12976) );
  NAND2_X1 U9556 ( .A1(n7555), .A2(n11865), .ZN(n7638) );
  XNOR2_X2 U9557 ( .A(n8264), .B(n8284), .ZN(n8835) );
  CLKBUF_X1 U9558 ( .A(n14421), .Z(n14423) );
  NAND2_X1 U9559 ( .A1(n10266), .A2(n10391), .ZN(n10264) );
  NAND2_X1 U9560 ( .A1(n8309), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8310) );
  NAND2_X1 U9561 ( .A1(n10819), .A2(n9820), .ZN(n10817) );
  INV_X1 U9562 ( .A(n12095), .ZN(n12097) );
  XNOR2_X1 U9563 ( .A(n12095), .B(n12096), .ZN(n12978) );
  NAND2_X1 U9564 ( .A1(n9218), .A2(n9230), .ZN(n12507) );
  NOR2_X1 U9565 ( .A1(n10270), .A2(n6618), .ZN(n10390) );
  AOI21_X2 U9566 ( .B1(n10809), .B2(n10808), .A(n9899), .ZN(n10970) );
  NOR2_X2 U9567 ( .A1(n9967), .A2(n9968), .ZN(n12093) );
  INV_X1 U9568 ( .A(n14265), .ZN(n11936) );
  AND2_X1 U9569 ( .A1(n8602), .A2(n11916), .ZN(n7522) );
  INV_X1 U9570 ( .A(n11096), .ZN(n11117) );
  INV_X1 U9571 ( .A(n8273), .ZN(n8278) );
  OR2_X1 U9572 ( .A1(n13404), .A2(n12094), .ZN(n7523) );
  AND2_X2 U9573 ( .A1(n11941), .A2(n14739), .ZN(n14157) );
  OR2_X1 U9575 ( .A1(n15378), .A2(n15368), .ZN(n12949) );
  INV_X1 U9576 ( .A(n12949), .ZN(n9832) );
  INV_X2 U9577 ( .A(n15330), .ZN(n15333) );
  BUF_X1 U9578 ( .A(n7634), .Z(n7672) );
  AND2_X1 U9579 ( .A1(n12524), .A2(n15302), .ZN(n7524) );
  AND2_X1 U9580 ( .A1(n9875), .A2(n9874), .ZN(n7525) );
  OR2_X1 U9581 ( .A1(n11168), .A2(n11167), .ZN(n7526) );
  OR2_X1 U9582 ( .A1(n15379), .A2(n13549), .ZN(n7528) );
  AND2_X1 U9583 ( .A1(n10760), .A2(n10759), .ZN(n7529) );
  INV_X1 U9584 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n8880) );
  CLKBUF_X2 U9585 ( .A(P1_U4016), .Z(n14655) );
  OR3_X1 U9586 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n10656), .ZN(n7530) );
  CLKBUF_X3 U9587 ( .A(n8364), .Z(n8701) );
  INV_X1 U9588 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13476) );
  AND2_X1 U9589 ( .A1(n7815), .A2(n7799), .ZN(n7532) );
  AND2_X1 U9590 ( .A1(n13459), .A2(n13063), .ZN(n7533) );
  INV_X1 U9591 ( .A(n13358), .ZN(n15055) );
  INV_X1 U9592 ( .A(n9817), .ZN(n12620) );
  INV_X1 U9593 ( .A(n12302), .ZN(n9281) );
  OR2_X1 U9594 ( .A1(n6580), .A2(n10407), .ZN(n7536) );
  NAND2_X1 U9595 ( .A1(n12429), .A2(n12430), .ZN(n7537) );
  OR2_X1 U9596 ( .A1(n13437), .A2(n13046), .ZN(n7538) );
  OR2_X1 U9597 ( .A1(n13181), .A2(n13180), .ZN(n7539) );
  MUX2_X1 U9598 ( .A(n11082), .B(n13085), .S(n9122), .Z(n8949) );
  NAND2_X1 U9599 ( .A1(n8954), .A2(n8953), .ZN(n8955) );
  INV_X1 U9600 ( .A(n8971), .ZN(n8972) );
  NAND2_X1 U9601 ( .A1(n8973), .A2(n8972), .ZN(n8977) );
  AND2_X1 U9602 ( .A1(n8620), .A2(n14132), .ZN(n8621) );
  INV_X1 U9603 ( .A(n9027), .ZN(n9028) );
  AOI21_X1 U9604 ( .B1(n9049), .B2(n9044), .A(n6631), .ZN(n9051) );
  INV_X1 U9605 ( .A(n8676), .ZN(n8677) );
  OR2_X1 U9606 ( .A1(n8680), .A2(n8679), .ZN(n8681) );
  INV_X1 U9607 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8259) );
  INV_X1 U9608 ( .A(n12732), .ZN(n9613) );
  INV_X1 U9609 ( .A(n12358), .ZN(n9323) );
  INV_X1 U9610 ( .A(n9963), .ZN(n9964) );
  INV_X1 U9611 ( .A(n11487), .ZN(n7791) );
  INV_X1 U9612 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7563) );
  INV_X1 U9613 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n13624) );
  NOR2_X1 U9614 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7547) );
  INV_X1 U9615 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7671) );
  INV_X1 U9616 ( .A(n13887), .ZN(n11906) );
  INV_X1 U9617 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9468) );
  NAND2_X1 U9618 ( .A1(n15217), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12585) );
  INV_X1 U9619 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12557) );
  INV_X1 U9620 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9378) );
  INV_X1 U9621 ( .A(n12482), .ZN(n9400) );
  INV_X1 U9622 ( .A(n12952), .ZN(n9797) );
  NOR2_X1 U9623 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n9518) );
  INV_X1 U9624 ( .A(n9866), .ZN(n9868) );
  NAND2_X1 U9625 ( .A1(n9114), .A2(n9115), .ZN(n9109) );
  INV_X1 U9626 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n13748) );
  INV_X1 U9627 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7864) );
  AND2_X1 U9628 ( .A1(n7782), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7805) );
  NOR2_X1 U9629 ( .A1(n8203), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8228) );
  INV_X1 U9630 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8446) );
  AND2_X1 U9631 ( .A1(n14528), .A2(n14529), .ZN(n11792) );
  BUF_X1 U9632 ( .A(n8544), .Z(n8780) );
  NOR2_X1 U9633 ( .A1(n8689), .A2(n8688), .ZN(n8699) );
  AND2_X1 U9634 ( .A1(P1_REG3_REG_21__SCAN_IN), .A2(n8641), .ZN(n8659) );
  NAND2_X1 U9635 ( .A1(n11907), .A2(n11906), .ZN(n11908) );
  INV_X1 U9636 ( .A(n11687), .ZN(n11686) );
  AND4_X1 U9637 ( .A1(n8262), .A2(n8823), .A3(n8826), .A4(n8822), .ZN(n8263)
         );
  INV_X1 U9638 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n9522) );
  OR2_X1 U9639 ( .A1(n9304), .A2(n10635), .ZN(n9240) );
  OAI22_X1 U9640 ( .A1(n12637), .A2(n15292), .B1(n12611), .B2(n12466), .ZN(
        n9746) );
  INV_X1 U9641 ( .A(n12492), .ZN(n9562) );
  OR2_X1 U9642 ( .A1(n9486), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9503) );
  OR2_X1 U9643 ( .A1(n12448), .A2(n12477), .ZN(n10480) );
  INV_X1 U9644 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n9539) );
  AND2_X1 U9645 ( .A1(n7805), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7822) );
  NAND2_X1 U9646 ( .A1(n12097), .A2(n12096), .ZN(n12098) );
  INV_X1 U9647 ( .A(n11363), .ZN(n9922) );
  INV_X1 U9648 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9688) );
  NAND2_X1 U9649 ( .A1(n9186), .A2(n9180), .ZN(n9183) );
  NOR2_X1 U9650 ( .A1(n7950), .A2(n12988), .ZN(n7967) );
  INV_X1 U9651 ( .A(n7606), .ZN(n7682) );
  INV_X1 U9652 ( .A(n9174), .ZN(n8195) );
  INV_X1 U9653 ( .A(n13206), .ZN(n8192) );
  OR2_X1 U9654 ( .A1(n15077), .A2(n9966), .ZN(n9974) );
  INV_X1 U9655 ( .A(n13426), .ZN(n8200) );
  OR2_X1 U9656 ( .A1(n7721), .A2(n7720), .ZN(n7743) );
  OR2_X1 U9657 ( .A1(n11039), .A2(n13022), .ZN(n11038) );
  AND2_X1 U9658 ( .A1(n15067), .A2(n8223), .ZN(n9966) );
  INV_X1 U9659 ( .A(n12035), .ZN(n12078) );
  OR2_X1 U9660 ( .A1(n8447), .A2(n8446), .ZN(n8457) );
  OR2_X1 U9661 ( .A1(n11796), .A2(n11795), .ZN(n11797) );
  AND2_X1 U9662 ( .A1(n11173), .A2(n11172), .ZN(n11174) );
  AND2_X1 U9663 ( .A1(n8699), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8714) );
  INV_X1 U9664 ( .A(n8290), .ZN(n8297) );
  INV_X1 U9665 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n13746) );
  AND2_X1 U9666 ( .A1(n10291), .A2(n10788), .ZN(n10300) );
  AND2_X1 U9667 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8383) );
  OR2_X1 U9668 ( .A1(n14246), .A2(n14121), .ZN(n14095) );
  INV_X1 U9669 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n13671) );
  INV_X1 U9670 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n13670) );
  INV_X1 U9671 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n8868) );
  INV_X1 U9672 ( .A(n11430), .ZN(n11426) );
  NOR2_X1 U9673 ( .A1(n9576), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9590) );
  AND2_X1 U9674 ( .A1(n9523), .A2(n9522), .ZN(n9543) );
  INV_X1 U9675 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n12258) );
  OR2_X1 U9676 ( .A1(n10840), .A2(n10839), .ZN(n12257) );
  AND2_X1 U9677 ( .A1(n9710), .A2(n9709), .ZN(n12618) );
  INV_X1 U9678 ( .A(n15163), .ZN(n12574) );
  INV_X1 U9679 ( .A(n14328), .ZN(n12554) );
  INV_X1 U9680 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14375) );
  INV_X1 U9681 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n12235) );
  INV_X1 U9682 ( .A(n9746), .ZN(n9747) );
  INV_X1 U9683 ( .A(n12670), .ZN(n12636) );
  AND2_X1 U9684 ( .A1(n12333), .A2(n12332), .ZN(n12718) );
  AND2_X1 U9685 ( .A1(n9358), .A2(n10681), .ZN(n9379) );
  AOI21_X1 U9686 ( .B1(n15287), .B2(n9752), .A(n9751), .ZN(n11227) );
  INV_X1 U9687 ( .A(n12950), .ZN(n10647) );
  AND2_X1 U9688 ( .A1(n12950), .A2(n12952), .ZN(n9823) );
  AND2_X1 U9689 ( .A1(n9821), .A2(n12323), .ZN(n15299) );
  INV_X1 U9690 ( .A(n15297), .ZN(n15327) );
  INV_X1 U9691 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n9317) );
  NAND2_X1 U9692 ( .A1(n12976), .A2(n12098), .ZN(n13007) );
  INV_X1 U9693 ( .A(n14450), .ZN(n13012) );
  AND2_X1 U9694 ( .A1(n7967), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7985) );
  OR2_X1 U9695 ( .A1(n7928), .A2(n7927), .ZN(n7950) );
  AND2_X1 U9696 ( .A1(n10179), .A2(n13481), .ZN(n10172) );
  INV_X1 U9697 ( .A(n15041), .ZN(n15022) );
  INV_X1 U9698 ( .A(n15028), .ZN(n15046) );
  NOR2_X1 U9699 ( .A1(n9974), .A2(n15076), .ZN(n9987) );
  INV_X1 U9700 ( .A(n13335), .ZN(n14441) );
  NAND2_X1 U9701 ( .A1(n10166), .A2(n9193), .ZN(n10381) );
  INV_X1 U9702 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9719) );
  INV_X1 U9703 ( .A(n9166), .ZN(n14462) );
  INV_X1 U9704 ( .A(n14456), .ZN(n13340) );
  INV_X1 U9705 ( .A(n9871), .ZN(n11855) );
  OAI21_X1 U9706 ( .B1(n8205), .B2(P2_IR_REG_24__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8206) );
  OR2_X1 U9707 ( .A1(n7944), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n7818) );
  INV_X1 U9708 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8525) );
  INV_X1 U9709 ( .A(n14547), .ZN(n14526) );
  INV_X1 U9710 ( .A(n10302), .ZN(n10288) );
  AND2_X1 U9711 ( .A1(n8598), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8616) );
  INV_X1 U9712 ( .A(n8740), .ZN(n8363) );
  INV_X1 U9713 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10368) );
  OR2_X1 U9714 ( .A1(n10611), .A2(n10612), .ZN(n10690) );
  INV_X1 U9715 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n13944) );
  NAND2_X1 U9716 ( .A1(n13887), .A2(n14178), .ZN(n11951) );
  INV_X1 U9717 ( .A(n11901), .ZN(n14054) );
  INV_X1 U9718 ( .A(n10389), .ZN(n11786) );
  NAND2_X1 U9719 ( .A1(n10292), .A2(n14560), .ZN(n14833) );
  INV_X1 U9720 ( .A(n14184), .ZN(n14584) );
  NAND2_X1 U9721 ( .A1(n14653), .A2(n10296), .ZN(n14555) );
  INV_X1 U9722 ( .A(n11107), .ZN(n14714) );
  OR2_X1 U9723 ( .A1(n11572), .A2(n13984), .ZN(n14786) );
  NOR2_X1 U9724 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n8279) );
  AND2_X1 U9725 ( .A1(n7875), .A2(n7857), .ZN(n7873) );
  INV_X1 U9726 ( .A(n12257), .ZN(n12291) );
  NAND2_X1 U9727 ( .A1(n10816), .A2(n12512), .ZN(n12295) );
  AOI21_X1 U9728 ( .B1(n12734), .B2(n9723), .A(n9612), .ZN(n12742) );
  OR2_X1 U9729 ( .A1(n9262), .A2(n9241), .ZN(n9245) );
  INV_X1 U9730 ( .A(n15184), .ZN(n15222) );
  INV_X1 U9731 ( .A(n15292), .ZN(n15323) );
  AND2_X1 U9732 ( .A1(n15330), .A2(n15250), .ZN(n15265) );
  AND2_X1 U9733 ( .A1(n12340), .A2(n15313), .ZN(n15329) );
  OAI22_X1 U9734 ( .A1(n12628), .A2(n12896), .B1(n15395), .B2(n9843), .ZN(
        n9844) );
  NOR3_X1 U9735 ( .A1(n10654), .A2(n9823), .A3(n9808), .ZN(n10652) );
  NAND2_X1 U9736 ( .A1(n9809), .A2(n10819), .ZN(n15368) );
  OR2_X1 U9737 ( .A1(n15297), .A2(n15377), .ZN(n15366) );
  AND2_X1 U9738 ( .A1(n9809), .A2(n15313), .ZN(n15377) );
  NOR2_X1 U9739 ( .A1(n12951), .A2(n10203), .ZN(n10205) );
  INV_X1 U9740 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n9232) );
  AND2_X1 U9741 ( .A1(n9551), .A2(n9534), .ZN(n9549) );
  AND2_X1 U9742 ( .A1(n9421), .A2(n9411), .ZN(n9419) );
  OAI21_X1 U9743 ( .B1(n13035), .B2(n13031), .A(n13032), .ZN(n12994) );
  INV_X1 U9744 ( .A(n14453), .ZN(n13014) );
  AND4_X1 U9745 ( .A1(n7888), .A2(n7887), .A3(n7886), .A4(n7885), .ZN(n11847)
         );
  INV_X1 U9746 ( .A(n15018), .ZN(n15035) );
  AND2_X1 U9747 ( .A1(n10179), .A2(n10175), .ZN(n15028) );
  INV_X1 U9748 ( .A(n14443), .ZN(n13336) );
  NAND2_X1 U9749 ( .A1(n15078), .A2(n9971), .ZN(n15052) );
  INV_X1 U9750 ( .A(n13360), .ZN(n15058) );
  INV_X1 U9751 ( .A(n15074), .ZN(n10383) );
  AND2_X1 U9752 ( .A1(n11005), .A2(n9193), .ZN(n14481) );
  AND2_X1 U9753 ( .A1(n8198), .A2(n10308), .ZN(n13440) );
  INV_X1 U9754 ( .A(n13440), .ZN(n14479) );
  NOR2_X1 U9755 ( .A1(n15074), .A2(n8236), .ZN(n9986) );
  INV_X1 U9756 ( .A(n14532), .ZN(n14551) );
  AND4_X1 U9757 ( .A1(n8667), .A2(n8666), .A3(n8665), .A4(n8664), .ZN(n13788)
         );
  AND4_X1 U9758 ( .A1(n8556), .A2(n8555), .A3(n8554), .A4(n8553), .ZN(n14493)
         );
  OR2_X1 U9759 ( .A1(n10086), .A2(n14653), .ZN(n14673) );
  AND2_X1 U9760 ( .A1(n10104), .A2(n14650), .ZN(n14684) );
  INV_X1 U9761 ( .A(n14132), .ZN(n14129) );
  AND2_X1 U9762 ( .A1(n11878), .A2(n10296), .ZN(n14177) );
  NOR2_X1 U9763 ( .A1(n14745), .A2(n13984), .ZN(n11582) );
  INV_X1 U9764 ( .A(n14734), .ZN(n14719) );
  INV_X1 U9765 ( .A(n14157), .ZN(n14741) );
  AND2_X1 U9766 ( .A1(n11583), .A2(n11570), .ZN(n11571) );
  INV_X1 U9767 ( .A(n14738), .ZN(n14837) );
  NAND2_X1 U9768 ( .A1(n10792), .A2(n10791), .ZN(n14738) );
  INV_X1 U9769 ( .A(n14793), .ZN(n14840) );
  INV_X1 U9770 ( .A(n14786), .ZN(n14830) );
  XNOR2_X1 U9771 ( .A(n8820), .B(n8822), .ZN(n10062) );
  AND2_X1 U9772 ( .A1(n8478), .A2(n8465), .ZN(n10189) );
  AND2_X1 U9773 ( .A1(n10431), .A2(n10430), .ZN(n15215) );
  INV_X1 U9774 ( .A(n12295), .ZN(n12178) );
  AND2_X1 U9775 ( .A1(n12310), .A2(n9745), .ZN(n12466) );
  NAND2_X1 U9776 ( .A1(n9626), .A2(n9625), .ZN(n12701) );
  INV_X1 U9777 ( .A(n12175), .ZN(n12791) );
  OR2_X1 U9778 ( .A1(n12526), .A2(n10420), .ZN(n15184) );
  INV_X1 U9779 ( .A(n15151), .ZN(n15228) );
  NAND2_X1 U9780 ( .A1(n15305), .A2(n15301), .ZN(n12812) );
  INV_X1 U9781 ( .A(n12901), .ZN(n12835) );
  NAND2_X1 U9782 ( .A1(n15395), .A2(n15301), .ZN(n12896) );
  AND3_X2 U9783 ( .A1(n10652), .A2(n9815), .A3(n9814), .ZN(n15395) );
  NAND2_X1 U9784 ( .A1(n9817), .A2(n9832), .ZN(n9833) );
  INV_X1 U9785 ( .A(n12209), .ZN(n12926) );
  INV_X2 U9786 ( .A(n15378), .ZN(n15379) );
  AND2_X1 U9787 ( .A1(n9829), .A2(n9828), .ZN(n15378) );
  OR2_X1 U9788 ( .A1(n10422), .A2(P3_U3151), .ZN(n12512) );
  INV_X1 U9789 ( .A(SI_17_), .ZN(n10316) );
  INV_X1 U9790 ( .A(SI_14_), .ZN(n10163) );
  NOR2_X1 U9791 ( .A1(n10179), .A2(P2_U3088), .ZN(n14872) );
  INV_X1 U9792 ( .A(n14451), .ZN(n13017) );
  OR3_X1 U9793 ( .A1(n9970), .A2(n10166), .A3(n14481), .ZN(n13059) );
  INV_X1 U9794 ( .A(n12120), .ZN(n13062) );
  OAI21_X1 U9795 ( .B1(n13306), .B2(n7640), .A(n7972), .ZN(n13069) );
  OR3_X1 U9796 ( .A1(n7912), .A2(n7911), .A3(n7910), .ZN(n13334) );
  INV_X1 U9797 ( .A(n14872), .ZN(n15050) );
  OR2_X1 U9798 ( .A1(n13358), .A2(n13161), .ZN(n15061) );
  NAND2_X1 U9799 ( .A1(n15105), .A2(n14481), .ZN(n13418) );
  OR3_X1 U9800 ( .A1(n10384), .A2(n10383), .A3(n10382), .ZN(n15103) );
  INV_X2 U9801 ( .A(n15103), .ZN(n15105) );
  INV_X1 U9802 ( .A(n13295), .ZN(n13469) );
  OR3_X1 U9803 ( .A1(n13448), .A2(n13447), .A3(n13446), .ZN(n13474) );
  INV_X1 U9804 ( .A(n15099), .ZN(n15098) );
  AND2_X2 U9805 ( .A1(n8237), .A2(n9986), .ZN(n15099) );
  INV_X1 U9806 ( .A(n15073), .ZN(n15071) );
  INV_X1 U9807 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10719) );
  INV_X1 U9808 ( .A(n14536), .ZN(n14549) );
  NAND2_X1 U9809 ( .A1(n10301), .A2(n10293), .ZN(n14532) );
  NAND4_X1 U9810 ( .A1(n8732), .A2(n8731), .A3(n8730), .A4(n8729), .ZN(n13887)
         );
  INV_X1 U9811 ( .A(n13799), .ZN(n14107) );
  INV_X1 U9812 ( .A(n14556), .ZN(n14544) );
  OR2_X1 U9813 ( .A1(n10086), .A2(n10085), .ZN(n14690) );
  INV_X1 U9814 ( .A(n14675), .ZN(n14695) );
  INV_X1 U9815 ( .A(n6575), .ZN(n14186) );
  INV_X1 U9816 ( .A(n14571), .ZN(n14189) );
  OR2_X1 U9817 ( .A1(n14157), .A2(n10938), .ZN(n14339) );
  INV_X1 U9818 ( .A(n14858), .ZN(n14856) );
  AND3_X1 U9819 ( .A1(n14581), .A2(n14580), .A3(n14579), .ZN(n14611) );
  AND2_X1 U9820 ( .A1(n14808), .A2(n14807), .ZN(n14852) );
  INV_X1 U9821 ( .A(n14844), .ZN(n14842) );
  INV_X1 U9822 ( .A(n14760), .ZN(n14759) );
  AND2_X1 U9823 ( .A1(n10062), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10054) );
  INV_X1 U9824 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10893) );
  INV_X1 U9825 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10321) );
  XNOR2_X1 U9826 ( .A(n8882), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15397) );
  XNOR2_X1 U9827 ( .A(n8940), .B(n12606), .ZN(n8941) );
  INV_X1 U9828 ( .A(n12526), .ZN(P3_U3897) );
  AND2_X1 U9829 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9854), .ZN(P2_U3947) );
  NAND2_X1 U9830 ( .A1(n8240), .A2(n8239), .ZN(P2_U3496) );
  NOR2_X1 U9831 ( .A1(n10260), .A2(n10072), .ZN(P1_U4016) );
  NOR2_X2 U9832 ( .A1(n7631), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n7634) );
  NOR2_X1 U9833 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n7543) );
  NAND4_X1 U9834 ( .A1(n7543), .A2(n7542), .A3(n7541), .A4(n7540), .ZN(n7942)
         );
  INV_X2 U9835 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8230) );
  INV_X2 U9836 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8134) );
  NAND2_X1 U9837 ( .A1(n8131), .A2(n8210), .ZN(n7549) );
  NAND2_X1 U9838 ( .A1(n7552), .A2(n7553), .ZN(n13475) );
  XNOR2_X2 U9839 ( .A(n7551), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7555) );
  INV_X1 U9840 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10458) );
  NAND2_X1 U9841 ( .A1(n7757), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7561) );
  NAND2_X2 U9842 ( .A1(n11875), .A2(n11865), .ZN(n7606) );
  INV_X1 U9843 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7556) );
  INV_X1 U9844 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7558) );
  NAND4_X1 U9845 ( .A1(n7560), .A2(n7561), .A3(n7562), .A4(n7559), .ZN(n9859)
         );
  NAND2_X1 U9846 ( .A1(n7566), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7567) );
  INV_X1 U9847 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10233) );
  INV_X1 U9848 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10008) );
  MUX2_X1 U9849 ( .A(n10233), .B(n10008), .S(n7596), .Z(n7592) );
  AND2_X1 U9850 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7569) );
  NAND2_X1 U9851 ( .A1(n10005), .A2(n7569), .ZN(n7582) );
  NAND2_X1 U9852 ( .A1(n7582), .A2(n8317), .ZN(n7591) );
  INV_X1 U9853 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7571) );
  NAND2_X1 U9854 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n13777), .ZN(n7570) );
  OR2_X1 U9855 ( .A1(n7583), .A2(n14868), .ZN(n7572) );
  NAND2_X1 U9856 ( .A1(n8156), .A2(n7573), .ZN(n7584) );
  INV_X1 U9857 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10173) );
  INV_X1 U9858 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7575) );
  INV_X1 U9859 ( .A(n7605), .ZN(n7576) );
  NAND2_X1 U9860 ( .A1(n7576), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7578) );
  INV_X1 U9861 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10174) );
  AND4_X2 U9862 ( .A1(n7580), .A2(n7579), .A3(n7578), .A4(n7577), .ZN(n8155)
         );
  INV_X1 U9863 ( .A(n9156), .ZN(n9995) );
  NAND2_X1 U9864 ( .A1(n7757), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7589) );
  INV_X1 U9865 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10450) );
  INV_X1 U9866 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7585) );
  INV_X1 U9867 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10341) );
  OR2_X1 U9868 ( .A1(n7608), .A2(n10341), .ZN(n7586) );
  NAND2_X1 U9869 ( .A1(n7591), .A2(n7590), .ZN(n7595) );
  INV_X1 U9870 ( .A(n7592), .ZN(n7593) );
  NAND2_X1 U9871 ( .A1(n7593), .A2(SI_1_), .ZN(n7594) );
  NAND2_X1 U9872 ( .A1(n7595), .A2(n7594), .ZN(n7617) );
  MUX2_X1 U9873 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n7596), .Z(n7618) );
  INV_X1 U9874 ( .A(SI_2_), .ZN(n10027) );
  XNOR2_X1 U9875 ( .A(n7618), .B(n10027), .ZN(n7616) );
  XNOR2_X1 U9876 ( .A(n7617), .B(n7616), .ZN(n10007) );
  INV_X1 U9877 ( .A(n7597), .ZN(n7598) );
  NAND2_X1 U9878 ( .A1(n7598), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7600) );
  XNOR2_X1 U9879 ( .A(n7600), .B(n7599), .ZN(n14879) );
  OR2_X1 U9880 ( .A1(n9119), .A2(n10003), .ZN(n7601) );
  NAND2_X1 U9881 ( .A1(n10460), .A2(n11082), .ZN(n7604) );
  NAND2_X1 U9882 ( .A1(n13085), .A2(n15080), .ZN(n7603) );
  NAND2_X1 U9883 ( .A1(n9100), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7612) );
  OR2_X1 U9884 ( .A1(n7640), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7611) );
  INV_X1 U9885 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7607) );
  OR2_X1 U9886 ( .A1(n8109), .A2(n7607), .ZN(n7610) );
  INV_X1 U9887 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10343) );
  OR2_X1 U9888 ( .A1(n9105), .A2(n10343), .ZN(n7609) );
  NAND2_X1 U9889 ( .A1(n7613), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7615) );
  INV_X1 U9890 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7614) );
  XNOR2_X1 U9891 ( .A(n7615), .B(n7614), .ZN(n13090) );
  NAND2_X1 U9892 ( .A1(n7617), .A2(n7616), .ZN(n7620) );
  NAND2_X1 U9893 ( .A1(n7618), .A2(SI_2_), .ZN(n7619) );
  XNOR2_X1 U9894 ( .A(n7627), .B(n7625), .ZN(n10004) );
  INV_X4 U9895 ( .A(n8032), .ZN(n9118) );
  NAND2_X1 U9896 ( .A1(n10004), .A2(n9118), .ZN(n7623) );
  OR2_X1 U9897 ( .A1(n9119), .A2(n7621), .ZN(n7622) );
  NAND2_X1 U9898 ( .A1(n10584), .A2(n10583), .ZN(n10582) );
  INV_X1 U9899 ( .A(n13084), .ZN(n11077) );
  NAND2_X1 U9900 ( .A1(n11077), .A2(n9871), .ZN(n7624) );
  INV_X1 U9901 ( .A(n7625), .ZN(n7626) );
  NAND2_X1 U9902 ( .A1(n7627), .A2(n7626), .ZN(n7630) );
  NAND2_X1 U9903 ( .A1(n7628), .A2(SI_3_), .ZN(n7629) );
  MUX2_X1 U9904 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n7076), .Z(n7655) );
  XNOR2_X1 U9905 ( .A(n7655), .B(SI_4_), .ZN(n7653) );
  XNOR2_X1 U9906 ( .A(n7654), .B(n7653), .ZN(n10013) );
  NAND2_X1 U9907 ( .A1(n10013), .A2(n9118), .ZN(n7637) );
  NAND2_X1 U9908 ( .A1(n7632), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7633) );
  MUX2_X1 U9909 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7633), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n7635) );
  INV_X1 U9910 ( .A(n7672), .ZN(n7657) );
  NAND2_X1 U9911 ( .A1(n7635), .A2(n7657), .ZN(n10345) );
  INV_X1 U9912 ( .A(n10345), .ZN(n14893) );
  AOI22_X1 U9913 ( .A1(n7947), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7946), .B2(
        n14893), .ZN(n7636) );
  INV_X1 U9914 ( .A(n13022), .ZN(n15086) );
  INV_X2 U9915 ( .A(n9105), .ZN(n8084) );
  NAND2_X1 U9916 ( .A1(n8084), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7645) );
  INV_X1 U9917 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7639) );
  OR2_X1 U9918 ( .A1(n8125), .A2(n7639), .ZN(n7644) );
  NAND2_X1 U9919 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7680) );
  OAI21_X1 U9920 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n7680), .ZN(n13024) );
  OR2_X1 U9921 ( .A1(n7640), .A2(n13024), .ZN(n7643) );
  INV_X1 U9922 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7641) );
  OR2_X1 U9923 ( .A1(n8109), .A2(n7641), .ZN(n7642) );
  NAND4_X2 U9924 ( .A1(n7645), .A2(n7644), .A3(n7643), .A4(n7642), .ZN(n13083)
         );
  INV_X1 U9925 ( .A(n11026), .ZN(n11031) );
  INV_X1 U9926 ( .A(n13083), .ZN(n10528) );
  NAND2_X1 U9927 ( .A1(n10528), .A2(n13022), .ZN(n7646) );
  NAND2_X1 U9928 ( .A1(n8084), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7652) );
  INV_X1 U9929 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7647) );
  OR2_X1 U9930 ( .A1(n8125), .A2(n7647), .ZN(n7651) );
  INV_X1 U9931 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7678) );
  XNOR2_X1 U9932 ( .A(n7680), .B(n7678), .ZN(n11240) );
  OR2_X1 U9933 ( .A1(n7640), .A2(n11240), .ZN(n7650) );
  INV_X1 U9934 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7648) );
  OR2_X1 U9935 ( .A1(n8109), .A2(n7648), .ZN(n7649) );
  NAND4_X1 U9936 ( .A1(n7652), .A2(n7651), .A3(n7650), .A4(n7649), .ZN(n13082)
         );
  INV_X1 U9937 ( .A(n13082), .ZN(n7662) );
  NAND2_X1 U9938 ( .A1(n7655), .A2(SI_4_), .ZN(n7656) );
  MUX2_X1 U9939 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7076), .Z(n7668) );
  XNOR2_X1 U9940 ( .A(n7668), .B(SI_5_), .ZN(n7665) );
  XNOR2_X1 U9941 ( .A(n7667), .B(n7665), .ZN(n10038) );
  NAND2_X1 U9942 ( .A1(n10038), .A2(n9118), .ZN(n7660) );
  NAND2_X1 U9943 ( .A1(n7657), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7658) );
  XNOR2_X1 U9944 ( .A(n7658), .B(P2_IR_REG_5__SCAN_IN), .ZN(n13104) );
  AOI22_X1 U9945 ( .A1(n7947), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7946), .B2(
        n13104), .ZN(n7659) );
  OR2_X1 U9946 ( .A1(n7662), .A2(n11242), .ZN(n7661) );
  NAND2_X1 U9947 ( .A1(n11242), .A2(n7662), .ZN(n7663) );
  NAND2_X1 U9948 ( .A1(n7664), .A2(n7663), .ZN(n10865) );
  INV_X1 U9949 ( .A(n7665), .ZN(n7666) );
  NAND2_X1 U9950 ( .A1(n7668), .A2(SI_5_), .ZN(n7669) );
  NAND2_X1 U9951 ( .A1(n7670), .A2(n7669), .ZN(n7692) );
  MUX2_X1 U9952 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7076), .Z(n7693) );
  XNOR2_X1 U9953 ( .A(n7693), .B(SI_6_), .ZN(n7690) );
  XNOR2_X1 U9954 ( .A(n7692), .B(n7690), .ZN(n10045) );
  NAND2_X1 U9955 ( .A1(n10045), .A2(n9118), .ZN(n7676) );
  INV_X1 U9956 ( .A(n7801), .ZN(n7673) );
  NAND2_X1 U9957 ( .A1(n7673), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7674) );
  XNOR2_X1 U9958 ( .A(n7674), .B(P2_IR_REG_6__SCAN_IN), .ZN(n14907) );
  AOI22_X1 U9959 ( .A1(n7947), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7946), .B2(
        n14907), .ZN(n7675) );
  NAND2_X1 U9960 ( .A1(n8084), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7687) );
  INV_X1 U9961 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11018) );
  OR2_X1 U9962 ( .A1(n8125), .A2(n11018), .ZN(n7686) );
  INV_X1 U9963 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7677) );
  OAI21_X1 U9964 ( .B1(n7680), .B2(n7678), .A(n7677), .ZN(n7681) );
  NAND2_X1 U9965 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_5__SCAN_IN), 
        .ZN(n7679) );
  NOR2_X1 U9966 ( .A1(n7680), .A2(n7679), .ZN(n7700) );
  INV_X1 U9967 ( .A(n7700), .ZN(n7702) );
  NAND2_X1 U9968 ( .A1(n7681), .A2(n7702), .ZN(n11019) );
  OR2_X1 U9969 ( .A1(n7640), .A2(n11019), .ZN(n7685) );
  INV_X1 U9970 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7683) );
  OR2_X1 U9971 ( .A1(n8109), .A2(n7683), .ZN(n7684) );
  NAND4_X1 U9972 ( .A1(n7687), .A2(n7686), .A3(n7685), .A4(n7684), .ZN(n13081)
         );
  XNOR2_X1 U9973 ( .A(n10869), .B(n13081), .ZN(n9161) );
  NAND2_X1 U9974 ( .A1(n10865), .A2(n9161), .ZN(n7689) );
  INV_X1 U9975 ( .A(n13081), .ZN(n10811) );
  NAND2_X1 U9976 ( .A1(n10869), .A2(n10811), .ZN(n7688) );
  NAND2_X1 U9977 ( .A1(n7689), .A2(n7688), .ZN(n10983) );
  INV_X1 U9978 ( .A(n7690), .ZN(n7691) );
  NAND2_X1 U9979 ( .A1(n7692), .A2(n7691), .ZN(n7695) );
  NAND2_X1 U9980 ( .A1(n7693), .A2(SI_6_), .ZN(n7694) );
  MUX2_X1 U9981 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7076), .Z(n7714) );
  XNOR2_X1 U9982 ( .A(n7714), .B(SI_7_), .ZN(n7711) );
  NAND2_X1 U9983 ( .A1(n10057), .A2(n9118), .ZN(n7699) );
  INV_X1 U9984 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7696) );
  NAND2_X1 U9985 ( .A1(n7801), .A2(n7696), .ZN(n7716) );
  NAND2_X1 U9986 ( .A1(n7716), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7697) );
  XNOR2_X1 U9987 ( .A(n7697), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U9988 ( .A1(n7947), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7946), .B2(
        n10349), .ZN(n7698) );
  NAND2_X1 U9989 ( .A1(n7699), .A2(n7698), .ZN(n15057) );
  NAND2_X1 U9990 ( .A1(n9101), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7708) );
  INV_X1 U9991 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n15054) );
  OR2_X1 U9992 ( .A1(n8125), .A2(n15054), .ZN(n7707) );
  NAND2_X1 U9993 ( .A1(n7700), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7721) );
  INV_X1 U9994 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7701) );
  NAND2_X1 U9995 ( .A1(n7702), .A2(n7701), .ZN(n7703) );
  NAND2_X1 U9996 ( .A1(n7721), .A2(n7703), .ZN(n15053) );
  OR2_X1 U9997 ( .A1(n7640), .A2(n15053), .ZN(n7706) );
  INV_X1 U9998 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7704) );
  OR2_X1 U9999 ( .A1(n9105), .A2(n7704), .ZN(n7705) );
  NAND4_X1 U10000 ( .A1(n7708), .A2(n7707), .A3(n7706), .A4(n7705), .ZN(n13080) );
  XNOR2_X1 U10001 ( .A(n15057), .B(n13080), .ZN(n10982) );
  INV_X1 U10002 ( .A(n10982), .ZN(n10980) );
  INV_X1 U10003 ( .A(n13080), .ZN(n7709) );
  OR2_X1 U10004 ( .A1(n15057), .A2(n7709), .ZN(n7710) );
  INV_X1 U10005 ( .A(n7711), .ZN(n7712) );
  NAND2_X1 U10006 ( .A1(n7714), .A2(SI_7_), .ZN(n7715) );
  MUX2_X1 U10007 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n7076), .Z(n7732) );
  XNOR2_X1 U10008 ( .A(n7732), .B(SI_8_), .ZN(n7729) );
  XNOR2_X1 U10009 ( .A(n7731), .B(n7729), .ZN(n10074) );
  NAND2_X1 U10010 ( .A1(n10074), .A2(n9118), .ZN(n7719) );
  NAND2_X1 U10011 ( .A1(n7734), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7717) );
  XNOR2_X1 U10012 ( .A(n7717), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10351) );
  AOI22_X1 U10013 ( .A1(n7947), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7946), .B2(
        n10351), .ZN(n7718) );
  NAND2_X1 U10014 ( .A1(n8084), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7727) );
  INV_X1 U10015 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11051) );
  OR2_X1 U10016 ( .A1(n8125), .A2(n11051), .ZN(n7726) );
  INV_X1 U10017 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7720) );
  NAND2_X1 U10018 ( .A1(n7721), .A2(n7720), .ZN(n7722) );
  NAND2_X1 U10019 ( .A1(n7743), .A2(n7722), .ZN(n11055) );
  OR2_X1 U10020 ( .A1(n7640), .A2(n11055), .ZN(n7725) );
  INV_X1 U10021 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7723) );
  OR2_X1 U10022 ( .A1(n8109), .A2(n7723), .ZN(n7724) );
  NAND4_X1 U10023 ( .A1(n7727), .A2(n7726), .A3(n7725), .A4(n7724), .ZN(n13079) );
  INV_X1 U10024 ( .A(n13079), .ZN(n10810) );
  XNOR2_X1 U10025 ( .A(n11052), .B(n10810), .ZN(n11045) );
  INV_X1 U10026 ( .A(n11045), .ZN(n11047) );
  NAND2_X1 U10027 ( .A1(n11048), .A2(n11047), .ZN(n11046) );
  OR2_X1 U10028 ( .A1(n11052), .A2(n10810), .ZN(n7728) );
  NAND2_X1 U10029 ( .A1(n11046), .A2(n7728), .ZN(n11212) );
  NAND2_X1 U10030 ( .A1(n7732), .A2(SI_8_), .ZN(n7733) );
  MUX2_X1 U10031 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n7076), .Z(n7753) );
  XNOR2_X1 U10032 ( .A(n7753), .B(SI_9_), .ZN(n7750) );
  XNOR2_X1 U10033 ( .A(n7752), .B(n7750), .ZN(n10078) );
  NAND2_X1 U10034 ( .A1(n10078), .A2(n9118), .ZN(n7742) );
  NAND2_X1 U10035 ( .A1(n7736), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7735) );
  MUX2_X1 U10036 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7735), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n7739) );
  INV_X1 U10037 ( .A(n7736), .ZN(n7738) );
  INV_X1 U10038 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7737) );
  NAND2_X1 U10039 ( .A1(n7738), .A2(n7737), .ZN(n7778) );
  NAND2_X1 U10040 ( .A1(n7739), .A2(n7778), .ZN(n10354) );
  OAI22_X1 U10041 ( .A1(n9119), .A2(n10237), .B1(n10354), .B2(n10167), .ZN(
        n7740) );
  INV_X1 U10042 ( .A(n7740), .ZN(n7741) );
  NAND2_X1 U10043 ( .A1(n9101), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7748) );
  INV_X1 U10044 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10333) );
  OR2_X1 U10045 ( .A1(n8125), .A2(n10333), .ZN(n7747) );
  NAND2_X1 U10046 ( .A1(n7743), .A2(n13748), .ZN(n7744) );
  NAND2_X1 U10047 ( .A1(n7760), .A2(n7744), .ZN(n11219) );
  OR2_X1 U10048 ( .A1(n7640), .A2(n11219), .ZN(n7746) );
  INV_X1 U10049 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10353) );
  OR2_X1 U10050 ( .A1(n9105), .A2(n10353), .ZN(n7745) );
  NAND4_X1 U10051 ( .A1(n7748), .A2(n7747), .A3(n7746), .A4(n7745), .ZN(n13078) );
  INV_X1 U10052 ( .A(n13078), .ZN(n11346) );
  XNOR2_X1 U10053 ( .A(n11339), .B(n11346), .ZN(n11213) );
  NAND2_X1 U10054 ( .A1(n11339), .A2(n11346), .ZN(n7749) );
  INV_X1 U10055 ( .A(n7750), .ZN(n7751) );
  MUX2_X1 U10056 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n7076), .Z(n7772) );
  XNOR2_X1 U10057 ( .A(n7772), .B(SI_10_), .ZN(n7769) );
  XNOR2_X1 U10058 ( .A(n7771), .B(n7769), .ZN(n10157) );
  NAND2_X1 U10059 ( .A1(n10157), .A2(n9118), .ZN(n7756) );
  NAND2_X1 U10060 ( .A1(n7778), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7754) );
  XNOR2_X1 U10061 ( .A(n7754), .B(P2_IR_REG_10__SCAN_IN), .ZN(n14964) );
  AOI22_X1 U10062 ( .A1(n14964), .A2(n7946), .B1(n7947), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n7755) );
  NAND2_X1 U10063 ( .A1(n9100), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7766) );
  INV_X1 U10064 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7758) );
  OR2_X1 U10065 ( .A1(n9105), .A2(n7758), .ZN(n7765) );
  INV_X1 U10066 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7759) );
  NOR2_X1 U10067 ( .A1(n7760), .A2(n7759), .ZN(n7782) );
  INV_X1 U10068 ( .A(n7782), .ZN(n7784) );
  NAND2_X1 U10069 ( .A1(n7760), .A2(n7759), .ZN(n7761) );
  NAND2_X1 U10070 ( .A1(n7784), .A2(n7761), .ZN(n11350) );
  OR2_X1 U10071 ( .A1(n7640), .A2(n11350), .ZN(n7764) );
  INV_X1 U10072 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7762) );
  OR2_X1 U10073 ( .A1(n8109), .A2(n7762), .ZN(n7763) );
  NAND4_X1 U10074 ( .A1(n7766), .A2(n7765), .A3(n7764), .A4(n7763), .ZN(n13077) );
  INV_X1 U10075 ( .A(n13077), .ZN(n11367) );
  AND2_X1 U10076 ( .A1(n11356), .A2(n11367), .ZN(n7767) );
  OR2_X1 U10077 ( .A1(n11356), .A2(n11367), .ZN(n7768) );
  INV_X1 U10078 ( .A(n7769), .ZN(n7770) );
  NAND2_X1 U10079 ( .A1(n7772), .A2(SI_10_), .ZN(n7773) );
  MUX2_X1 U10080 ( .A(n10202), .B(n10199), .S(n7076), .Z(n7775) );
  NAND2_X1 U10081 ( .A1(n7775), .A2(n10044), .ZN(n7796) );
  INV_X1 U10082 ( .A(n7775), .ZN(n7776) );
  NAND2_X1 U10083 ( .A1(n7776), .A2(SI_11_), .ZN(n7777) );
  NAND2_X1 U10084 ( .A1(n7796), .A2(n7777), .ZN(n7794) );
  XNOR2_X1 U10085 ( .A(n7795), .B(n7794), .ZN(n10198) );
  NAND2_X1 U10086 ( .A1(n10198), .A2(n9118), .ZN(n7781) );
  OAI21_X1 U10087 ( .B1(n7778), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7779) );
  XNOR2_X1 U10088 ( .A(n7779), .B(P2_IR_REG_11__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U10089 ( .A1(n13122), .A2(n7946), .B1(n7947), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n7780) );
  NAND2_X1 U10090 ( .A1(n8084), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7790) );
  INV_X1 U10091 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11495) );
  OR2_X1 U10092 ( .A1(n8125), .A2(n11495), .ZN(n7789) );
  INV_X1 U10093 ( .A(n7805), .ZN(n7807) );
  INV_X1 U10094 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7783) );
  NAND2_X1 U10095 ( .A1(n7784), .A2(n7783), .ZN(n7785) );
  NAND2_X1 U10096 ( .A1(n7807), .A2(n7785), .ZN(n11494) );
  OR2_X1 U10097 ( .A1(n7640), .A2(n11494), .ZN(n7788) );
  INV_X1 U10098 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7786) );
  OR2_X1 U10099 ( .A1(n8109), .A2(n7786), .ZN(n7787) );
  NAND4_X1 U10100 ( .A1(n7790), .A2(n7789), .A3(n7788), .A4(n7787), .ZN(n13076) );
  INV_X1 U10101 ( .A(n13076), .ZN(n11383) );
  XNOR2_X1 U10102 ( .A(n11551), .B(n11383), .ZN(n11487) );
  NAND2_X1 U10103 ( .A1(n11551), .A2(n11383), .ZN(n7793) );
  MUX2_X1 U10104 ( .A(n10315), .B(n10312), .S(n7076), .Z(n7797) );
  NAND2_X1 U10105 ( .A1(n7797), .A2(n10056), .ZN(n7815) );
  INV_X1 U10106 ( .A(n7797), .ZN(n7798) );
  NAND2_X1 U10107 ( .A1(n7798), .A2(SI_12_), .ZN(n7799) );
  XNOR2_X1 U10108 ( .A(n7814), .B(n7532), .ZN(n10311) );
  NAND2_X1 U10109 ( .A1(n10311), .A2(n9118), .ZN(n7804) );
  NAND2_X1 U10110 ( .A1(n7801), .A2(n7800), .ZN(n7944) );
  NAND2_X1 U10111 ( .A1(n7944), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7802) );
  XNOR2_X1 U10112 ( .A(n7802), .B(P2_IR_REG_12__SCAN_IN), .ZN(n13139) );
  AOI22_X1 U10113 ( .A1(n7947), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7946), 
        .B2(n13139), .ZN(n7803) );
  NAND2_X1 U10114 ( .A1(n9101), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7812) );
  INV_X1 U10115 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n13115) );
  OR2_X1 U10116 ( .A1(n9105), .A2(n13115), .ZN(n7811) );
  INV_X1 U10117 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n13120) );
  OR2_X1 U10118 ( .A1(n8125), .A2(n13120), .ZN(n7810) );
  INV_X1 U10119 ( .A(n7822), .ZN(n7823) );
  INV_X1 U10120 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7806) );
  NAND2_X1 U10121 ( .A1(n7807), .A2(n7806), .ZN(n7808) );
  NAND2_X1 U10122 ( .A1(n7823), .A2(n7808), .ZN(n11468) );
  OR2_X1 U10123 ( .A1(n7640), .A2(n11468), .ZN(n7809) );
  NAND4_X1 U10124 ( .A1(n7812), .A2(n7811), .A3(n7810), .A4(n7809), .ZN(n13075) );
  INV_X1 U10125 ( .A(n13075), .ZN(n11366) );
  XNOR2_X1 U10126 ( .A(n14482), .B(n11366), .ZN(n11459) );
  OR2_X1 U10127 ( .A1(n14482), .A2(n11366), .ZN(n7813) );
  MUX2_X1 U10128 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7076), .Z(n7831) );
  XNOR2_X1 U10129 ( .A(n7831), .B(n13723), .ZN(n7830) );
  XNOR2_X1 U10130 ( .A(n7834), .B(n7830), .ZN(n10318) );
  NAND2_X1 U10131 ( .A1(n10318), .A2(n9118), .ZN(n7821) );
  NAND2_X1 U10132 ( .A1(n7818), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7817) );
  MUX2_X1 U10133 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7817), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n7819) );
  NAND2_X1 U10134 ( .A1(n7819), .A2(n7858), .ZN(n13141) );
  INV_X1 U10135 ( .A(n13141), .ZN(n14976) );
  AOI22_X1 U10136 ( .A1(n7947), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7946), 
        .B2(n14976), .ZN(n7820) );
  NAND2_X1 U10137 ( .A1(n9100), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7829) );
  NAND2_X1 U10138 ( .A1(n7822), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7843) );
  INV_X1 U10139 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n13632) );
  NAND2_X1 U10140 ( .A1(n7823), .A2(n13632), .ZN(n7824) );
  NAND2_X1 U10141 ( .A1(n7843), .A2(n7824), .ZN(n11561) );
  OR2_X1 U10142 ( .A1(n7640), .A2(n11561), .ZN(n7828) );
  INV_X1 U10143 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7825) );
  OR2_X1 U10144 ( .A1(n8109), .A2(n7825), .ZN(n7827) );
  INV_X1 U10145 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n13131) );
  OR2_X1 U10146 ( .A1(n9105), .A2(n13131), .ZN(n7826) );
  NAND4_X1 U10147 ( .A1(n7829), .A2(n7828), .A3(n7827), .A4(n7826), .ZN(n13074) );
  INV_X1 U10148 ( .A(n13074), .ZN(n14442) );
  INV_X1 U10149 ( .A(n11563), .ZN(n14477) );
  INV_X1 U10150 ( .A(n7830), .ZN(n7833) );
  NAND2_X1 U10151 ( .A1(n7831), .A2(SI_13_), .ZN(n7832) );
  MUX2_X1 U10152 ( .A(n10416), .B(n10414), .S(n7076), .Z(n7835) );
  NAND2_X1 U10153 ( .A1(n7835), .A2(n10163), .ZN(n7852) );
  INV_X1 U10154 ( .A(n7835), .ZN(n7836) );
  NAND2_X1 U10155 ( .A1(n7836), .A2(SI_14_), .ZN(n7837) );
  NAND2_X1 U10156 ( .A1(n7852), .A2(n7837), .ZN(n7853) );
  XNOR2_X1 U10157 ( .A(n7854), .B(n7853), .ZN(n10413) );
  NAND2_X1 U10158 ( .A1(n10413), .A2(n9118), .ZN(n7840) );
  NAND2_X1 U10159 ( .A1(n7858), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7838) );
  XNOR2_X1 U10160 ( .A(n7838), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14988) );
  AOI22_X1 U10161 ( .A1(n7947), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7946), 
        .B2(n14988), .ZN(n7839) );
  NAND2_X1 U10162 ( .A1(n9100), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7848) );
  INV_X1 U10163 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7841) );
  OR2_X1 U10164 ( .A1(n8109), .A2(n7841), .ZN(n7847) );
  INV_X1 U10165 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n13132) );
  OR2_X1 U10166 ( .A1(n9105), .A2(n13132), .ZN(n7846) );
  INV_X1 U10167 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7842) );
  NAND2_X1 U10168 ( .A1(n7843), .A2(n7842), .ZN(n7844) );
  NAND2_X1 U10169 ( .A1(n7865), .A2(n7844), .ZN(n14458) );
  OR2_X1 U10170 ( .A1(n7640), .A2(n14458), .ZN(n7845) );
  NAND4_X1 U10171 ( .A1(n7848), .A2(n7847), .A3(n7846), .A4(n7845), .ZN(n13073) );
  INV_X1 U10172 ( .A(n13073), .ZN(n7849) );
  XNOR2_X1 U10173 ( .A(n14461), .B(n7849), .ZN(n9166) );
  NAND2_X1 U10174 ( .A1(n14454), .A2(n14462), .ZN(n7851) );
  NAND2_X1 U10175 ( .A1(n14461), .A2(n7849), .ZN(n7850) );
  NAND2_X1 U10176 ( .A1(n7851), .A2(n7850), .ZN(n11757) );
  MUX2_X1 U10177 ( .A(n10719), .B(n10717), .S(n7076), .Z(n7855) );
  NAND2_X1 U10178 ( .A1(n7855), .A2(n9500), .ZN(n7875) );
  INV_X1 U10179 ( .A(n7855), .ZN(n7856) );
  NAND2_X1 U10180 ( .A1(n7856), .A2(SI_15_), .ZN(n7857) );
  XNOR2_X1 U10181 ( .A(n7874), .B(n7873), .ZN(n10716) );
  NAND2_X1 U10182 ( .A1(n10716), .A2(n9118), .ZN(n7863) );
  INV_X1 U10183 ( .A(n7858), .ZN(n7860) );
  INV_X1 U10184 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7859) );
  NAND2_X1 U10185 ( .A1(n7860), .A2(n7859), .ZN(n7880) );
  NAND2_X1 U10186 ( .A1(n7880), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7861) );
  XNOR2_X1 U10187 ( .A(n7861), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14999) );
  AOI22_X1 U10188 ( .A1(n14999), .A2(n7946), .B1(n7947), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n7862) );
  NAND2_X1 U10189 ( .A1(n9101), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7870) );
  INV_X1 U10190 ( .A(n7907), .ZN(n7905) );
  NAND2_X1 U10191 ( .A1(n7865), .A2(n7864), .ZN(n7866) );
  NAND2_X1 U10192 ( .A1(n7905), .A2(n7866), .ZN(n11753) );
  OR2_X1 U10193 ( .A1(n11753), .A2(n7640), .ZN(n7869) );
  INV_X1 U10194 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14995) );
  OR2_X1 U10195 ( .A1(n9105), .A2(n14995), .ZN(n7868) );
  INV_X1 U10196 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n11754) );
  OR2_X1 U10197 ( .A1(n8125), .A2(n11754), .ZN(n7867) );
  NAND4_X1 U10198 ( .A1(n7870), .A2(n7869), .A3(n7868), .A4(n7867), .ZN(n13072) );
  XNOR2_X1 U10199 ( .A(n11841), .B(n13072), .ZN(n11758) );
  NAND2_X1 U10200 ( .A1(n11757), .A2(n11758), .ZN(n7872) );
  INV_X1 U10201 ( .A(n13072), .ZN(n14444) );
  NAND2_X1 U10202 ( .A1(n11841), .A2(n14444), .ZN(n7871) );
  MUX2_X1 U10203 ( .A(n10774), .B(n10773), .S(n7076), .Z(n7877) );
  NAND2_X1 U10204 ( .A1(n7877), .A2(n13582), .ZN(n7893) );
  INV_X1 U10205 ( .A(n7877), .ZN(n7878) );
  NAND2_X1 U10206 ( .A1(n7878), .A2(SI_16_), .ZN(n7879) );
  XNOR2_X1 U10207 ( .A(n7892), .B(n7891), .ZN(n10772) );
  NAND2_X1 U10208 ( .A1(n10772), .A2(n9118), .ZN(n7884) );
  NOR2_X1 U10209 ( .A1(n7880), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n7898) );
  INV_X1 U10210 ( .A(n7898), .ZN(n7881) );
  NAND2_X1 U10211 ( .A1(n7881), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7882) );
  XNOR2_X1 U10212 ( .A(n7882), .B(P2_IR_REG_16__SCAN_IN), .ZN(n15012) );
  AOI22_X1 U10213 ( .A1(n15012), .A2(n7946), .B1(n7947), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n7883) );
  XNOR2_X1 U10214 ( .A(n7905), .B(P2_REG3_REG_16__SCAN_IN), .ZN(n11825) );
  NAND2_X1 U10215 ( .A1(n11825), .A2(n7576), .ZN(n7888) );
  NAND2_X1 U10216 ( .A1(n8084), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7887) );
  NAND2_X1 U10217 ( .A1(n9100), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7886) );
  NAND2_X1 U10218 ( .A1(n9101), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7885) );
  INV_X1 U10219 ( .A(n11847), .ZN(n13071) );
  NOR2_X1 U10220 ( .A1(n13445), .A2(n13071), .ZN(n7889) );
  NAND2_X1 U10221 ( .A1(n13445), .A2(n13071), .ZN(n7890) );
  NAND2_X1 U10222 ( .A1(n7894), .A2(n10316), .ZN(n7918) );
  INV_X1 U10223 ( .A(n7894), .ZN(n7895) );
  NAND2_X1 U10224 ( .A1(n7895), .A2(SI_17_), .ZN(n7896) );
  XNOR2_X1 U10225 ( .A(n7917), .B(n7916), .ZN(n10892) );
  NAND2_X1 U10226 ( .A1(n10892), .A2(n9118), .ZN(n7902) );
  INV_X1 U10227 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7897) );
  NAND2_X1 U10228 ( .A1(n7898), .A2(n7897), .ZN(n7899) );
  NAND2_X1 U10229 ( .A1(n7899), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7920) );
  XNOR2_X1 U10230 ( .A(n7920), .B(P2_IR_REG_17__SCAN_IN), .ZN(n15027) );
  NOR2_X1 U10231 ( .A1(n9119), .A2(n13735), .ZN(n7900) );
  AOI21_X1 U10232 ( .B1(n15027), .B2(n7946), .A(n7900), .ZN(n7901) );
  INV_X1 U10233 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7904) );
  INV_X1 U10234 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7903) );
  OAI21_X1 U10235 ( .B1(n7905), .B2(n7904), .A(n7903), .ZN(n7908) );
  AND2_X1 U10236 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n7906) );
  NAND2_X1 U10237 ( .A1(n7907), .A2(n7906), .ZN(n7928) );
  NAND2_X1 U10238 ( .A1(n7908), .A2(n7928), .ZN(n13356) );
  NOR2_X1 U10239 ( .A1(n13356), .A2(n7640), .ZN(n7912) );
  INV_X1 U10240 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n7909) );
  NOR2_X1 U10241 ( .A1(n8109), .A2(n7909), .ZN(n7911) );
  INV_X1 U10242 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13611) );
  INV_X1 U10243 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13150) );
  OAI22_X1 U10244 ( .A1(n9105), .A2(n13611), .B1(n8125), .B2(n13150), .ZN(
        n7910) );
  INV_X1 U10245 ( .A(n13334), .ZN(n13046) );
  NAND2_X1 U10246 ( .A1(n7913), .A2(n7538), .ZN(n7915) );
  NAND2_X1 U10247 ( .A1(n13437), .A2(n13046), .ZN(n7914) );
  NAND2_X1 U10248 ( .A1(n7915), .A2(n7914), .ZN(n13331) );
  XNOR2_X1 U10249 ( .A(n7937), .B(n7935), .ZN(n11131) );
  NAND2_X1 U10250 ( .A1(n11131), .A2(n9118), .ZN(n7926) );
  INV_X1 U10251 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7919) );
  NAND2_X1 U10252 ( .A1(n7920), .A2(n7919), .ZN(n7921) );
  NAND2_X1 U10253 ( .A1(n7921), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7923) );
  INV_X1 U10254 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7922) );
  XNOR2_X1 U10255 ( .A(n7923), .B(n7922), .ZN(n15045) );
  OAI22_X1 U10256 ( .A1(n15045), .A2(n10167), .B1(n9119), .B2(n11135), .ZN(
        n7924) );
  INV_X1 U10257 ( .A(n7924), .ZN(n7925) );
  INV_X1 U10258 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7927) );
  NAND2_X1 U10259 ( .A1(n7928), .A2(n7927), .ZN(n7929) );
  NAND2_X1 U10260 ( .A1(n7950), .A2(n7929), .ZN(n13342) );
  AOI22_X1 U10261 ( .A1(n8084), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n9100), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n7931) );
  NAND2_X1 U10262 ( .A1(n9101), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7930) );
  OAI211_X1 U10263 ( .C1(n13342), .C2(n7640), .A(n7931), .B(n7930), .ZN(n13070) );
  INV_X1 U10264 ( .A(n13070), .ZN(n8178) );
  OR2_X1 U10265 ( .A1(n13429), .A2(n8178), .ZN(n7932) );
  NAND2_X1 U10266 ( .A1(n13331), .A2(n7932), .ZN(n7934) );
  NAND2_X1 U10267 ( .A1(n13429), .A2(n8178), .ZN(n7933) );
  INV_X1 U10268 ( .A(n7935), .ZN(n7936) );
  NAND2_X1 U10269 ( .A1(n7937), .A2(n7936), .ZN(n7941) );
  INV_X1 U10270 ( .A(n7938), .ZN(n7939) );
  NAND2_X1 U10271 ( .A1(n7939), .A2(SI_18_), .ZN(n7940) );
  XNOR2_X1 U10272 ( .A(n7961), .B(SI_19_), .ZN(n7958) );
  XNOR2_X1 U10273 ( .A(n7960), .B(n7958), .ZN(n11191) );
  NAND2_X1 U10274 ( .A1(n11191), .A2(n9118), .ZN(n7949) );
  AOI22_X1 U10276 ( .A1(n7947), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7946), 
        .B2(n13161), .ZN(n7948) );
  INV_X1 U10277 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n7955) );
  INV_X1 U10278 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n12988) );
  INV_X1 U10279 ( .A(n7967), .ZN(n7952) );
  NAND2_X1 U10280 ( .A1(n7950), .A2(n12988), .ZN(n7951) );
  NAND2_X1 U10281 ( .A1(n7952), .A2(n7951), .ZN(n12987) );
  OR2_X1 U10282 ( .A1(n12987), .A2(n7640), .ZN(n7954) );
  AOI22_X1 U10283 ( .A1(n8084), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n9100), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n7953) );
  OAI211_X1 U10284 ( .C1(n8109), .C2(n7955), .A(n7954), .B(n7953), .ZN(n13337)
         );
  INV_X1 U10285 ( .A(n13337), .ZN(n13043) );
  OR2_X1 U10286 ( .A1(n13426), .A2(n13043), .ZN(n7956) );
  NAND2_X1 U10287 ( .A1(n13426), .A2(n13043), .ZN(n7957) );
  INV_X1 U10288 ( .A(n7958), .ZN(n7959) );
  NAND2_X1 U10289 ( .A1(n7960), .A2(n7959), .ZN(n7963) );
  NAND2_X1 U10290 ( .A1(n7961), .A2(SI_19_), .ZN(n7962) );
  XNOR2_X1 U10291 ( .A(n7974), .B(SI_20_), .ZN(n7964) );
  XNOR2_X1 U10292 ( .A(n7978), .B(n7964), .ZN(n11260) );
  NAND2_X1 U10293 ( .A1(n11260), .A2(n9118), .ZN(n7966) );
  OR2_X1 U10294 ( .A1(n9119), .A2(n7319), .ZN(n7965) );
  NOR2_X1 U10295 ( .A1(n7967), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7968) );
  OR2_X1 U10296 ( .A1(n7985), .A2(n7968), .ZN(n13306) );
  INV_X1 U10297 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n13637) );
  NAND2_X1 U10298 ( .A1(n8084), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n7970) );
  NAND2_X1 U10299 ( .A1(n9100), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n7969) );
  OAI211_X1 U10300 ( .C1(n13637), .C2(n8109), .A(n7970), .B(n7969), .ZN(n7971)
         );
  INV_X1 U10301 ( .A(n7971), .ZN(n7972) );
  XNOR2_X1 U10302 ( .A(n13420), .B(n13069), .ZN(n13310) );
  INV_X1 U10303 ( .A(n13069), .ZN(n7973) );
  NOR2_X1 U10304 ( .A1(n7975), .A2(n10751), .ZN(n7977) );
  NAND2_X1 U10305 ( .A1(n7975), .A2(n10751), .ZN(n7976) );
  NAND2_X1 U10306 ( .A1(n7979), .A2(SI_21_), .ZN(n7994) );
  OAI21_X1 U10307 ( .B1(n7979), .B2(SI_21_), .A(n7994), .ZN(n7980) );
  NAND2_X1 U10308 ( .A1(n7981), .A2(n7980), .ZN(n7982) );
  NAND2_X1 U10309 ( .A1(n7995), .A2(n7982), .ZN(n11372) );
  OR2_X1 U10310 ( .A1(n11372), .A2(n8032), .ZN(n7984) );
  INV_X1 U10311 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11374) );
  OR2_X1 U10312 ( .A1(n9119), .A2(n11374), .ZN(n7983) );
  OR2_X1 U10313 ( .A1(n7985), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U10314 ( .A1(n7985), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8000) );
  AND2_X1 U10315 ( .A1(n7986), .A2(n8000), .ZN(n13296) );
  NAND2_X1 U10316 ( .A1(n13296), .A2(n7576), .ZN(n7991) );
  INV_X1 U10317 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13709) );
  NAND2_X1 U10318 ( .A1(n8084), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n7988) );
  NAND2_X1 U10319 ( .A1(n9100), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7987) );
  OAI211_X1 U10320 ( .C1(n13709), .C2(n8109), .A(n7988), .B(n7987), .ZN(n7989)
         );
  INV_X1 U10321 ( .A(n7989), .ZN(n7990) );
  NAND2_X1 U10322 ( .A1(n7991), .A2(n7990), .ZN(n13272) );
  INV_X1 U10323 ( .A(n13272), .ZN(n13036) );
  AND2_X1 U10324 ( .A1(n13295), .A2(n13036), .ZN(n7993) );
  OR2_X1 U10325 ( .A1(n13295), .A2(n13036), .ZN(n7992) );
  XNOR2_X1 U10326 ( .A(n8656), .B(n8009), .ZN(n11588) );
  NAND2_X1 U10327 ( .A1(n11588), .A2(n9118), .ZN(n7998) );
  OR2_X1 U10328 ( .A1(n9119), .A2(n11591), .ZN(n7997) );
  NAND2_X1 U10329 ( .A1(n8084), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8007) );
  INV_X1 U10330 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n7999) );
  OR2_X1 U10331 ( .A1(n8125), .A2(n7999), .ZN(n8006) );
  INV_X1 U10332 ( .A(n8000), .ZN(n8002) );
  INV_X1 U10333 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9978) );
  INV_X1 U10334 ( .A(n8013), .ZN(n8001) );
  OAI21_X1 U10335 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(n8002), .A(n8001), .ZN(
        n13276) );
  OR2_X1 U10336 ( .A1(n7640), .A2(n13276), .ZN(n8005) );
  INV_X1 U10337 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8003) );
  OR2_X1 U10338 ( .A1(n8109), .A2(n8003), .ZN(n8004) );
  NAND4_X1 U10339 ( .A1(n8007), .A2(n8006), .A3(n8005), .A4(n8004), .ZN(n13068) );
  INV_X1 U10340 ( .A(n13068), .ZN(n13263) );
  XNOR2_X1 U10341 ( .A(n13409), .B(n13263), .ZN(n13269) );
  INV_X1 U10342 ( .A(n13269), .ZN(n13280) );
  OR2_X1 U10343 ( .A1(n13409), .A2(n13263), .ZN(n8008) );
  NAND2_X1 U10344 ( .A1(n8010), .A2(SI_23_), .ZN(n8022) );
  OAI21_X1 U10345 ( .B1(n8010), .B2(SI_23_), .A(n8022), .ZN(n8021) );
  XNOR2_X1 U10346 ( .A(n8025), .B(n8021), .ZN(n11614) );
  NAND2_X1 U10347 ( .A1(n11614), .A2(n9118), .ZN(n8012) );
  INV_X1 U10348 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11613) );
  OR2_X1 U10349 ( .A1(n9119), .A2(n11613), .ZN(n8011) );
  NAND2_X1 U10350 ( .A1(n8084), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8018) );
  INV_X1 U10351 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13257) );
  OR2_X1 U10352 ( .A1(n8125), .A2(n13257), .ZN(n8017) );
  NAND2_X1 U10353 ( .A1(n8013), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8036) );
  OAI21_X1 U10354 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n8013), .A(n8036), .ZN(
        n13265) );
  OR2_X1 U10355 ( .A1(n7640), .A2(n13265), .ZN(n8016) );
  INV_X1 U10356 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8014) );
  OR2_X1 U10357 ( .A1(n8109), .A2(n8014), .ZN(n8015) );
  NAND4_X1 U10358 ( .A1(n8018), .A2(n8017), .A3(n8016), .A4(n8015), .ZN(n13271) );
  INV_X1 U10359 ( .A(n13271), .ZN(n12094) );
  NAND2_X1 U10360 ( .A1(n13404), .A2(n12094), .ZN(n8019) );
  INV_X1 U10361 ( .A(n8021), .ZN(n8024) );
  INV_X1 U10362 ( .A(n8022), .ZN(n8023) );
  MUX2_X1 U10363 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7076), .Z(n8026) );
  NAND2_X1 U10364 ( .A1(n8026), .A2(SI_24_), .ZN(n8044) );
  OAI21_X1 U10365 ( .B1(n8026), .B2(SI_24_), .A(n8044), .ZN(n8028) );
  NAND2_X1 U10366 ( .A1(n8027), .A2(n8028), .ZN(n8031) );
  INV_X1 U10367 ( .A(n8027), .ZN(n8030) );
  INV_X1 U10368 ( .A(n8028), .ZN(n8029) );
  OR2_X1 U10369 ( .A1(n11697), .A2(n8032), .ZN(n8034) );
  OR2_X1 U10370 ( .A1(n9119), .A2(n13595), .ZN(n8033) );
  NAND2_X1 U10371 ( .A1(n9100), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8042) );
  INV_X1 U10372 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8035) );
  OR2_X1 U10373 ( .A1(n9105), .A2(n8035), .ZN(n8041) );
  INV_X1 U10374 ( .A(n8036), .ZN(n8037) );
  NAND2_X1 U10375 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n8037), .ZN(n8050) );
  OAI21_X1 U10376 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n8037), .A(n8050), .ZN(
        n13010) );
  OR2_X1 U10377 ( .A1(n7640), .A2(n13010), .ZN(n8040) );
  INV_X1 U10378 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8038) );
  OR2_X1 U10379 ( .A1(n8109), .A2(n8038), .ZN(n8039) );
  NAND4_X1 U10380 ( .A1(n8042), .A2(n8041), .A3(n8040), .A4(n8039), .ZN(n13067) );
  INV_X1 U10381 ( .A(n13067), .ZN(n13262) );
  NAND2_X1 U10382 ( .A1(n13249), .A2(n13262), .ZN(n8043) );
  XNOR2_X1 U10383 ( .A(n8058), .B(SI_25_), .ZN(n8061) );
  XNOR2_X1 U10384 ( .A(n8062), .B(n8061), .ZN(n13772) );
  NAND2_X1 U10385 ( .A1(n13772), .A2(n9118), .ZN(n8046) );
  INV_X1 U10386 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13775) );
  OR2_X1 U10387 ( .A1(n9119), .A2(n13775), .ZN(n8045) );
  NAND2_X1 U10388 ( .A1(n8084), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8056) );
  INV_X1 U10389 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8047) );
  OR2_X1 U10390 ( .A1(n8125), .A2(n8047), .ZN(n8055) );
  INV_X1 U10391 ( .A(n8050), .ZN(n8048) );
  NAND2_X1 U10392 ( .A1(n8048), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8068) );
  INV_X1 U10393 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U10394 ( .A1(n8050), .A2(n8049), .ZN(n8051) );
  NAND2_X1 U10395 ( .A1(n8068), .A2(n8051), .ZN(n13232) );
  OR2_X1 U10396 ( .A1(n7640), .A2(n13232), .ZN(n8054) );
  INV_X1 U10397 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8052) );
  OR2_X1 U10398 ( .A1(n8109), .A2(n8052), .ZN(n8053) );
  NAND4_X1 U10399 ( .A1(n8056), .A2(n8055), .A3(n8054), .A4(n8053), .ZN(n13066) );
  XNOR2_X1 U10400 ( .A(n13392), .B(n13066), .ZN(n13230) );
  INV_X1 U10401 ( .A(n13066), .ZN(n8057) );
  INV_X1 U10402 ( .A(n8058), .ZN(n8059) );
  INV_X1 U10403 ( .A(SI_25_), .ZN(n11502) );
  NAND2_X1 U10404 ( .A1(n8059), .A2(n11502), .ZN(n8060) );
  INV_X1 U10405 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14299) );
  XNOR2_X1 U10406 ( .A(n8078), .B(SI_26_), .ZN(n8063) );
  NAND2_X1 U10407 ( .A1(n14297), .A2(n9118), .ZN(n8065) );
  OR2_X1 U10408 ( .A1(n9119), .A2(n9688), .ZN(n8064) );
  NAND2_X1 U10409 ( .A1(n8084), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8074) );
  INV_X1 U10410 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8066) );
  OR2_X1 U10411 ( .A1(n8125), .A2(n8066), .ZN(n8073) );
  INV_X1 U10412 ( .A(n8068), .ZN(n8067) );
  NAND2_X1 U10413 ( .A1(n8067), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8104) );
  INV_X1 U10414 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13707) );
  NAND2_X1 U10415 ( .A1(n8068), .A2(n13707), .ZN(n8069) );
  NAND2_X1 U10416 ( .A1(n8104), .A2(n8069), .ZN(n13217) );
  OR2_X1 U10417 ( .A1(n7640), .A2(n13217), .ZN(n8072) );
  INV_X1 U10418 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8070) );
  OR2_X1 U10419 ( .A1(n8109), .A2(n8070), .ZN(n8071) );
  NAND4_X1 U10420 ( .A1(n8074), .A2(n8073), .A3(n8072), .A4(n8071), .ZN(n13065) );
  INV_X1 U10421 ( .A(n13065), .ZN(n13001) );
  XNOR2_X1 U10422 ( .A(n13387), .B(n13001), .ZN(n13215) );
  INV_X1 U10423 ( .A(n13215), .ZN(n13211) );
  NAND2_X1 U10424 ( .A1(n13210), .A2(n13211), .ZN(n8076) );
  NAND2_X1 U10425 ( .A1(n13387), .A2(n13001), .ZN(n8075) );
  NAND2_X1 U10426 ( .A1(n8076), .A2(n8075), .ZN(n13194) );
  INV_X1 U10427 ( .A(n8078), .ZN(n8077) );
  NOR2_X1 U10428 ( .A1(n8077), .A2(SI_26_), .ZN(n8079) );
  INV_X1 U10429 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13486) );
  INV_X1 U10430 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14296) );
  XNOR2_X1 U10431 ( .A(n8094), .B(SI_27_), .ZN(n8092) );
  INV_X1 U10432 ( .A(n8092), .ZN(n8081) );
  NAND2_X1 U10433 ( .A1(n14293), .A2(n9118), .ZN(n8083) );
  OR2_X1 U10434 ( .A1(n9119), .A2(n13486), .ZN(n8082) );
  NAND2_X1 U10435 ( .A1(n8084), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8090) );
  INV_X1 U10436 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8085) );
  OR2_X1 U10437 ( .A1(n8125), .A2(n8085), .ZN(n8089) );
  INV_X1 U10438 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12972) );
  XNOR2_X1 U10439 ( .A(n8104), .B(n12972), .ZN(n12968) );
  OR2_X1 U10440 ( .A1(n7640), .A2(n12968), .ZN(n8088) );
  INV_X1 U10441 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8086) );
  OR2_X1 U10442 ( .A1(n8109), .A2(n8086), .ZN(n8087) );
  XNOR2_X1 U10443 ( .A(n7105), .B(n13064), .ZN(n13206) );
  NOR2_X1 U10444 ( .A1(n13202), .A2(n13064), .ZN(n8091) );
  INV_X1 U10445 ( .A(n8094), .ZN(n8095) );
  NAND2_X1 U10446 ( .A1(n8095), .A2(SI_27_), .ZN(n8117) );
  INV_X1 U10447 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11877) );
  INV_X1 U10448 ( .A(SI_28_), .ZN(n11723) );
  NAND2_X1 U10449 ( .A1(n8096), .A2(n11723), .ZN(n8120) );
  INV_X1 U10450 ( .A(n8096), .ZN(n8097) );
  NAND2_X1 U10451 ( .A1(n8097), .A2(SI_28_), .ZN(n8098) );
  NAND2_X1 U10452 ( .A1(n8120), .A2(n8098), .ZN(n8115) );
  NAND2_X1 U10453 ( .A1(n11876), .A2(n9118), .ZN(n8101) );
  OR2_X1 U10454 ( .A1(n9119), .A2(n9719), .ZN(n8100) );
  NAND2_X1 U10455 ( .A1(n9100), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8113) );
  INV_X1 U10456 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8102) );
  OR2_X1 U10457 ( .A1(n9105), .A2(n8102), .ZN(n8112) );
  INV_X1 U10458 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8103) );
  OAI21_X1 U10459 ( .B1(n8104), .B2(n12972), .A(n8103), .ZN(n8107) );
  INV_X1 U10460 ( .A(n8104), .ZN(n8106) );
  AND2_X1 U10461 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n8105) );
  NAND2_X1 U10462 ( .A1(n8106), .A2(n8105), .ZN(n11879) );
  NAND2_X1 U10463 ( .A1(n8107), .A2(n11879), .ZN(n13185) );
  OR2_X1 U10464 ( .A1(n7640), .A2(n13185), .ZN(n8111) );
  INV_X1 U10465 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8108) );
  OR2_X1 U10466 ( .A1(n8109), .A2(n8108), .ZN(n8110) );
  NAND2_X1 U10467 ( .A1(n7104), .A2(n13063), .ZN(n8194) );
  OR2_X1 U10468 ( .A1(n7104), .A2(n13063), .ZN(n8114) );
  NAND2_X1 U10469 ( .A1(n8194), .A2(n8114), .ZN(n13180) );
  INV_X1 U10470 ( .A(n8115), .ZN(n8116) );
  AND2_X1 U10471 ( .A1(n8117), .A2(n8116), .ZN(n8118) );
  NAND2_X1 U10472 ( .A1(n8119), .A2(n8118), .ZN(n8121) );
  INV_X1 U10473 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n11867) );
  XNOR2_X1 U10474 ( .A(n8243), .B(SI_29_), .ZN(n8241) );
  XNOR2_X1 U10475 ( .A(n8242), .B(n8241), .ZN(n11864) );
  NAND2_X1 U10476 ( .A1(n11864), .A2(n9118), .ZN(n8123) );
  OR2_X1 U10477 ( .A1(n9119), .A2(n11867), .ZN(n8122) );
  NAND2_X1 U10478 ( .A1(n9101), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8129) );
  INV_X1 U10479 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n13663) );
  OR2_X1 U10480 ( .A1(n9105), .A2(n13663), .ZN(n8128) );
  INV_X1 U10481 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8124) );
  OR2_X1 U10482 ( .A1(n8125), .A2(n8124), .ZN(n8127) );
  OR2_X1 U10483 ( .A1(n7640), .A2(n11879), .ZN(n8126) );
  AND4_X1 U10484 ( .A1(n8129), .A2(n8128), .A3(n8127), .A4(n8126), .ZN(n12120)
         );
  XNOR2_X1 U10485 ( .A(n7099), .B(n13062), .ZN(n9174) );
  XNOR2_X1 U10486 ( .A(n8130), .B(n9174), .ZN(n8154) );
  XNOR2_X2 U10487 ( .A(n8135), .B(n8134), .ZN(n11590) );
  NAND2_X1 U10488 ( .A1(n9195), .A2(n13161), .ZN(n9124) );
  NAND2_X1 U10489 ( .A1(n8141), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8136) );
  INV_X1 U10490 ( .A(n8138), .ZN(n8139) );
  NAND2_X1 U10491 ( .A1(n8139), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8140) );
  INV_X1 U10492 ( .A(n11262), .ZN(n9123) );
  NAND2_X1 U10493 ( .A1(n9179), .A2(n9123), .ZN(n8143) );
  INV_X1 U10494 ( .A(n8145), .ZN(n8146) );
  INV_X1 U10495 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13375) );
  NAND2_X1 U10496 ( .A1(n9100), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8148) );
  NAND2_X1 U10497 ( .A1(n9101), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8147) );
  OAI211_X1 U10498 ( .C1(n9105), .C2(n13375), .A(n8148), .B(n8147), .ZN(n13061) );
  NAND2_X1 U10499 ( .A1(n10166), .A2(n8145), .ZN(n14443) );
  INV_X1 U10500 ( .A(P2_B_REG_SCAN_IN), .ZN(n8149) );
  NOR2_X1 U10501 ( .A1(n6740), .A2(n8149), .ZN(n8150) );
  NOR2_X1 U10502 ( .A1(n14443), .A2(n8150), .ZN(n13167) );
  AND2_X1 U10503 ( .A1(n13061), .A2(n13167), .ZN(n8151) );
  NAND2_X1 U10504 ( .A1(n8156), .A2(n10595), .ZN(n8157) );
  NAND2_X1 U10505 ( .A1(n11073), .A2(n11072), .ZN(n11071) );
  NAND2_X1 U10506 ( .A1(n10460), .A2(n15080), .ZN(n8158) );
  NAND2_X1 U10507 ( .A1(n11071), .A2(n8158), .ZN(n10579) );
  INV_X1 U10508 ( .A(n10583), .ZN(n10578) );
  NAND2_X1 U10509 ( .A1(n10579), .A2(n10578), .ZN(n10581) );
  NAND2_X1 U10510 ( .A1(n11077), .A2(n11855), .ZN(n8159) );
  NAND2_X1 U10511 ( .A1(n10581), .A2(n8159), .ZN(n11027) );
  NAND2_X1 U10512 ( .A1(n10528), .A2(n15086), .ZN(n8160) );
  NAND2_X1 U10513 ( .A1(n11029), .A2(n8160), .ZN(n10896) );
  XNOR2_X1 U10514 ( .A(n11242), .B(n13082), .ZN(n9160) );
  INV_X1 U10515 ( .A(n9160), .ZN(n10901) );
  NAND2_X1 U10516 ( .A1(n10896), .A2(n10901), .ZN(n10898) );
  OR2_X1 U10517 ( .A1(n11242), .A2(n13082), .ZN(n8161) );
  NAND2_X1 U10518 ( .A1(n10898), .A2(n8161), .ZN(n10862) );
  INV_X1 U10519 ( .A(n9161), .ZN(n10866) );
  OR2_X1 U10520 ( .A1(n10869), .A2(n13081), .ZN(n8162) );
  NAND2_X1 U10521 ( .A1(n10861), .A2(n8162), .ZN(n10981) );
  NAND2_X1 U10522 ( .A1(n10981), .A2(n10980), .ZN(n10979) );
  OR2_X1 U10523 ( .A1(n15057), .A2(n13080), .ZN(n8163) );
  NAND2_X1 U10524 ( .A1(n11052), .A2(n13079), .ZN(n8164) );
  XNOR2_X1 U10525 ( .A(n11356), .B(n11367), .ZN(n11345) );
  NAND2_X1 U10526 ( .A1(n11342), .A2(n11345), .ZN(n8166) );
  NAND2_X1 U10527 ( .A1(n11356), .A2(n13077), .ZN(n8165) );
  AND2_X1 U10528 ( .A1(n11551), .A2(n13076), .ZN(n8167) );
  INV_X1 U10529 ( .A(n8167), .ZN(n8168) );
  OR2_X1 U10530 ( .A1(n11551), .A2(n13076), .ZN(n8169) );
  NOR2_X1 U10531 ( .A1(n14482), .A2(n13075), .ZN(n8170) );
  OR2_X1 U10532 ( .A1(n11563), .A2(n13074), .ZN(n8171) );
  NAND2_X1 U10533 ( .A1(n11558), .A2(n8171), .ZN(n8173) );
  NAND2_X1 U10534 ( .A1(n11563), .A2(n13074), .ZN(n8172) );
  AND2_X1 U10535 ( .A1(n14461), .A2(n13073), .ZN(n8174) );
  OR2_X1 U10536 ( .A1(n14461), .A2(n13073), .ZN(n8175) );
  INV_X1 U10537 ( .A(n11758), .ZN(n11750) );
  NOR2_X1 U10538 ( .A1(n11841), .A2(n13072), .ZN(n8176) );
  XNOR2_X1 U10539 ( .A(n11829), .B(n13071), .ZN(n11764) );
  INV_X1 U10540 ( .A(n11764), .ZN(n11772) );
  NAND2_X1 U10541 ( .A1(n11773), .A2(n11772), .ZN(n13442) );
  OR2_X1 U10542 ( .A1(n13445), .A2(n11847), .ZN(n8177) );
  NAND2_X1 U10543 ( .A1(n13437), .A2(n13334), .ZN(n9154) );
  INV_X1 U10544 ( .A(n9154), .ZN(n9038) );
  NOR2_X1 U10545 ( .A1(n13437), .A2(n13334), .ZN(n9035) );
  INV_X1 U10546 ( .A(n9035), .ZN(n9155) );
  XNOR2_X1 U10547 ( .A(n13429), .B(n8178), .ZN(n13332) );
  OR2_X1 U10548 ( .A1(n13429), .A2(n13070), .ZN(n8179) );
  NAND2_X1 U10549 ( .A1(n13330), .A2(n8179), .ZN(n13315) );
  NAND2_X1 U10550 ( .A1(n13426), .A2(n13337), .ZN(n8180) );
  OR2_X1 U10551 ( .A1(n13426), .A2(n13337), .ZN(n8181) );
  NOR2_X1 U10552 ( .A1(n13420), .A2(n13069), .ZN(n8184) );
  NAND2_X1 U10553 ( .A1(n13420), .A2(n13069), .ZN(n8183) );
  XNOR2_X1 U10554 ( .A(n13295), .B(n13272), .ZN(n13290) );
  OR2_X1 U10555 ( .A1(n13295), .A2(n13272), .ZN(n8185) );
  INV_X1 U10556 ( .A(n13281), .ZN(n8186) );
  NAND2_X1 U10557 ( .A1(n8186), .A2(n13269), .ZN(n13283) );
  NAND2_X1 U10558 ( .A1(n13409), .A2(n13068), .ZN(n8187) );
  AND2_X1 U10559 ( .A1(n13404), .A2(n13271), .ZN(n8189) );
  OR2_X1 U10560 ( .A1(n13404), .A2(n13271), .ZN(n8188) );
  NAND2_X1 U10561 ( .A1(n13249), .A2(n13067), .ZN(n8190) );
  OR2_X1 U10562 ( .A1(n13392), .A2(n13066), .ZN(n8191) );
  OR2_X1 U10563 ( .A1(n13202), .A2(n13053), .ZN(n8193) );
  NAND2_X1 U10564 ( .A1(n13205), .A2(n8193), .ZN(n13177) );
  INV_X1 U10565 ( .A(n13180), .ZN(n13176) );
  NAND2_X1 U10566 ( .A1(n13177), .A2(n13176), .ZN(n13179) );
  XNOR2_X1 U10567 ( .A(n11590), .B(n9856), .ZN(n8197) );
  INV_X1 U10568 ( .A(n14461), .ZN(n14472) );
  NAND2_X1 U10569 ( .A1(n11012), .A2(n10595), .ZN(n11083) );
  NOR2_X1 U10570 ( .A1(n11083), .A2(n11082), .ZN(n11086) );
  NAND2_X1 U10571 ( .A1(n11086), .A2(n11855), .ZN(n11039) );
  INV_X1 U10572 ( .A(n15057), .ZN(n10990) );
  INV_X1 U10573 ( .A(n11356), .ZN(n15093) );
  INV_X1 U10574 ( .A(n11551), .ZN(n11548) );
  NOR2_X1 U10575 ( .A1(n13420), .A2(n13321), .ZN(n13305) );
  OR2_X2 U10576 ( .A1(n13392), .A2(n13247), .ZN(n13234) );
  INV_X1 U10577 ( .A(n13188), .ZN(n8201) );
  AND2_X4 U10578 ( .A1(n11005), .A2(n11262), .ZN(n14465) );
  AOI211_X1 U10579 ( .C1(n7099), .C2(n8201), .A(n9935), .B(n13172), .ZN(n11885) );
  AOI21_X1 U10580 ( .B1(n14481), .B2(n7099), .A(n11885), .ZN(n8202) );
  NAND2_X1 U10581 ( .A1(n8228), .A2(n8230), .ZN(n8205) );
  NAND2_X1 U10582 ( .A1(n8205), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8204) );
  XNOR2_X1 U10583 ( .A(n11696), .B(P2_B_REG_SCAN_IN), .ZN(n8207) );
  OR2_X1 U10584 ( .A1(n8207), .A2(n13773), .ZN(n8212) );
  NOR4_X1 U10585 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n8216) );
  NOR4_X1 U10586 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n8215) );
  NOR4_X1 U10587 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8214) );
  NOR4_X1 U10588 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8213) );
  AND4_X1 U10589 ( .A1(n8216), .A2(n8215), .A3(n8214), .A4(n8213), .ZN(n8222)
         );
  NOR2_X1 U10590 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .ZN(
        n8220) );
  NOR4_X1 U10591 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n8219) );
  NOR4_X1 U10592 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n8218) );
  NOR4_X1 U10593 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n8217) );
  AND4_X1 U10594 ( .A1(n8220), .A2(n8219), .A3(n8218), .A4(n8217), .ZN(n8221)
         );
  NAND2_X1 U10595 ( .A1(n8222), .A2(n8221), .ZN(n8223) );
  INV_X1 U10596 ( .A(n9966), .ZN(n8227) );
  INV_X1 U10597 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n8224) );
  NAND2_X1 U10598 ( .A1(n15067), .A2(n8224), .ZN(n8226) );
  OR2_X1 U10599 ( .A1(n13773), .A2(n13768), .ZN(n8225) );
  NAND2_X1 U10600 ( .A1(n8226), .A2(n8225), .ZN(n15077) );
  NAND3_X1 U10601 ( .A1(n8227), .A2(n15077), .A3(n9973), .ZN(n10384) );
  NAND2_X1 U10602 ( .A1(n13773), .A2(n11696), .ZN(n9853) );
  INV_X1 U10603 ( .A(n8228), .ZN(n8229) );
  NAND2_X1 U10604 ( .A1(n8229), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8231) );
  NOR2_X1 U10605 ( .A1(n10384), .A2(n15076), .ZN(n8237) );
  INV_X1 U10606 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n8233) );
  NAND2_X1 U10607 ( .A1(n15067), .A2(n8233), .ZN(n8235) );
  OR2_X1 U10608 ( .A1(n11696), .A2(n13768), .ZN(n8234) );
  INV_X1 U10609 ( .A(n10381), .ZN(n8236) );
  NAND2_X1 U10610 ( .A1(n13377), .A2(n15099), .ZN(n8240) );
  INV_X1 U10611 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8238) );
  OR2_X1 U10612 ( .A1(n15099), .A2(n8238), .ZN(n8239) );
  NAND2_X1 U10613 ( .A1(n8242), .A2(n8241), .ZN(n8245) );
  NAND2_X1 U10614 ( .A1(n8243), .A2(n13652), .ZN(n8244) );
  NAND2_X1 U10615 ( .A1(n8245), .A2(n8244), .ZN(n8763) );
  NAND2_X1 U10616 ( .A1(n8246), .A2(SI_30_), .ZN(n8247) );
  OAI21_X1 U10617 ( .B1(SI_30_), .B2(n8246), .A(n8247), .ZN(n8762) );
  NAND2_X1 U10618 ( .A1(n8765), .A2(n8247), .ZN(n8250) );
  XNOR2_X1 U10619 ( .A(n8248), .B(SI_31_), .ZN(n8249) );
  NOR2_X1 U10620 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), 
        .ZN(n8254) );
  NOR2_X1 U10621 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8256) );
  NOR2_X1 U10622 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), 
        .ZN(n8260) );
  NOR2_X1 U10623 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n8262) );
  NAND2_X1 U10624 ( .A1(n14285), .A2(n8766), .ZN(n8267) );
  INV_X1 U10625 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14290) );
  OR2_X1 U10626 ( .A1(n8767), .A2(n14290), .ZN(n8266) );
  INV_X1 U10627 ( .A(n8270), .ZN(n8275) );
  NAND2_X1 U10628 ( .A1(n8275), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8268) );
  MUX2_X1 U10629 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8268), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n8271) );
  NAND2_X1 U10630 ( .A1(n8278), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8274) );
  MUX2_X1 U10631 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8274), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n8276) );
  NAND2_X1 U10632 ( .A1(n8593), .A2(n8277), .ZN(n8588) );
  NOR2_X1 U10633 ( .A1(n8273), .A2(n8279), .ZN(n8280) );
  NAND2_X1 U10634 ( .A1(n8282), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8281) );
  MUX2_X1 U10635 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8281), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n8283) );
  NOR2_X1 U10636 ( .A1(n13996), .A2(n8775), .ZN(n8809) );
  NAND2_X4 U10637 ( .A1(n11966), .A2(n8297), .ZN(n8740) );
  INV_X1 U10638 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8289) );
  NOR2_X1 U10639 ( .A1(n8740), .A2(n8289), .ZN(n8294) );
  INV_X2 U10640 ( .A(n6587), .ZN(n8713) );
  INV_X1 U10641 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n13992) );
  NOR2_X1 U10642 ( .A1(n8713), .A2(n13992), .ZN(n8293) );
  INV_X1 U10643 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n13630) );
  NOR2_X1 U10644 ( .A1(n6584), .A2(n13630), .ZN(n8292) );
  NAND2_X1 U10645 ( .A1(n14307), .A2(n10790), .ZN(n8832) );
  NAND2_X1 U10646 ( .A1(n10788), .A2(n11261), .ZN(n11572) );
  NAND2_X1 U10647 ( .A1(n8832), .A2(n11572), .ZN(n8295) );
  NOR2_X2 U10648 ( .A1(n11360), .A2(n10789), .ZN(n10779) );
  NAND2_X1 U10649 ( .A1(n10779), .A2(n10937), .ZN(n10946) );
  NAND2_X1 U10650 ( .A1(n8295), .A2(n10946), .ZN(n8814) );
  NAND2_X1 U10651 ( .A1(n11360), .A2(n10789), .ZN(n10290) );
  NAND2_X1 U10652 ( .A1(n8814), .A2(n10290), .ZN(n8805) );
  NAND2_X1 U10653 ( .A1(n13996), .A2(n8775), .ZN(n8807) );
  NOR2_X1 U10654 ( .A1(n8807), .A2(n13994), .ZN(n8296) );
  AOI211_X1 U10655 ( .C1(n8809), .C2(n13994), .A(n8805), .B(n8296), .ZN(n8819)
         );
  NAND2_X1 U10656 ( .A1(n8298), .A2(n8297), .ZN(n8364) );
  INV_X1 U10657 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n8299) );
  OR2_X1 U10658 ( .A1(n8364), .A2(n8299), .ZN(n8305) );
  INV_X1 U10659 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n8300) );
  INV_X1 U10660 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n8301) );
  NAND2_X1 U10661 ( .A1(n6587), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8302) );
  OR2_X1 U10662 ( .A1(n8683), .A2(n10009), .ZN(n8308) );
  NAND2_X1 U10663 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8306) );
  XNOR2_X1 U10664 ( .A(n8306), .B(P1_IR_REG_1__SCAN_IN), .ZN(n13904) );
  NAND2_X1 U10665 ( .A1(n10299), .A2(n14770), .ZN(n10794) );
  NAND2_X1 U10666 ( .A1(n6587), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8311) );
  INV_X1 U10667 ( .A(n6582), .ZN(n8309) );
  INV_X1 U10668 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n8312) );
  INV_X1 U10669 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10915) );
  NAND3_X2 U10670 ( .A1(n8315), .A2(n8314), .A3(n8313), .ZN(n10960) );
  INV_X1 U10671 ( .A(n10960), .ZN(n8320) );
  INV_X1 U10672 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n13900) );
  NAND2_X1 U10673 ( .A1(n8316), .A2(n7005), .ZN(n8318) );
  NAND2_X1 U10674 ( .A1(n8318), .A2(n8317), .ZN(n14309) );
  MUX2_X1 U10675 ( .A(n13900), .B(n14309), .S(n10064), .Z(n10953) );
  INV_X1 U10676 ( .A(n10953), .ZN(n8319) );
  NAND2_X1 U10677 ( .A1(n8320), .A2(n8319), .ZN(n10793) );
  NOR2_X1 U10678 ( .A1(n10793), .A2(n8544), .ZN(n8325) );
  NAND2_X1 U10679 ( .A1(n8325), .A2(n10781), .ZN(n8324) );
  OAI21_X1 U10680 ( .B1(n8319), .B2(n10779), .A(n8320), .ZN(n8322) );
  NAND2_X1 U10681 ( .A1(n8319), .A2(n10779), .ZN(n8321) );
  NAND4_X1 U10682 ( .A1(n8322), .A2(n10796), .A3(n8544), .A4(n8321), .ZN(n8323) );
  OAI211_X1 U10683 ( .C1(n8775), .C2(n10794), .A(n8324), .B(n8323), .ZN(n8339)
         );
  INV_X1 U10684 ( .A(n8325), .ZN(n8327) );
  OR2_X1 U10685 ( .A1(n10299), .A2(n8544), .ZN(n8326) );
  AOI21_X1 U10686 ( .B1(n8327), .B2(n8326), .A(n14770), .ZN(n8338) );
  NAND2_X1 U10687 ( .A1(n6588), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8334) );
  INV_X1 U10688 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n8328) );
  OR2_X1 U10689 ( .A1(n8364), .A2(n8328), .ZN(n8333) );
  INV_X1 U10690 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n8329) );
  INV_X1 U10691 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n8330) );
  OR2_X1 U10692 ( .A1(n6584), .A2(n8330), .ZN(n8331) );
  OR2_X1 U10693 ( .A1(n8683), .A2(n10007), .ZN(n8337) );
  INV_X1 U10694 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10006) );
  OR2_X1 U10695 ( .A1(n8335), .A2(n8592), .ZN(n8336) );
  XNOR2_X1 U10696 ( .A(n8336), .B(P1_IR_REG_2__SCAN_IN), .ZN(n14649) );
  OAI21_X1 U10697 ( .B1(n8339), .B2(n8338), .A(n10941), .ZN(n8357) );
  INV_X1 U10698 ( .A(n8340), .ZN(n8342) );
  INV_X1 U10699 ( .A(n10798), .ZN(n8341) );
  INV_X1 U10700 ( .A(n8343), .ZN(n8356) );
  INV_X1 U10701 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n14740) );
  OR2_X1 U10702 ( .A1(n8713), .A2(n14740), .ZN(n8349) );
  OR2_X1 U10703 ( .A1(n8364), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U10704 ( .A1(n8363), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8347) );
  INV_X1 U10705 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n8344) );
  OR2_X1 U10706 ( .A1(n6584), .A2(n8344), .ZN(n8346) );
  NAND4_X2 U10707 ( .A1(n8349), .A2(n8348), .A3(n8347), .A4(n8346), .ZN(n13897) );
  NAND2_X1 U10708 ( .A1(n8477), .A2(n10004), .ZN(n8355) );
  NOR2_X1 U10709 ( .A1(n8352), .A2(n8592), .ZN(n8350) );
  MUX2_X1 U10710 ( .A(n8592), .B(n8350), .S(P1_IR_REG_3__SCAN_IN), .Z(n8353)
         );
  INV_X1 U10711 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8351) );
  AND2_X1 U10712 ( .A1(n8352), .A2(n8351), .ZN(n8373) );
  NOR2_X1 U10713 ( .A1(n8353), .A2(n8373), .ZN(n13915) );
  NAND2_X1 U10714 ( .A1(n8612), .A2(n13915), .ZN(n8354) );
  OAI211_X2 U10715 ( .C1(n8767), .C2(n7054), .A(n8355), .B(n8354), .ZN(n14782)
         );
  XNOR2_X1 U10716 ( .A(n13897), .B(n14782), .ZN(n14733) );
  NAND3_X1 U10717 ( .A1(n8357), .A2(n8356), .A3(n14733), .ZN(n8362) );
  INV_X1 U10718 ( .A(n14782), .ZN(n8358) );
  AND2_X1 U10719 ( .A1(n13897), .A2(n8358), .ZN(n8359) );
  NOR2_X1 U10720 ( .A1(n13897), .A2(n8358), .ZN(n10799) );
  INV_X1 U10721 ( .A(n8360), .ZN(n8361) );
  NAND2_X1 U10722 ( .A1(n8362), .A2(n8361), .ZN(n8380) );
  NAND2_X1 U10723 ( .A1(n8363), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8372) );
  INV_X1 U10724 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10803) );
  OR2_X1 U10725 ( .A1(n8713), .A2(n10803), .ZN(n8371) );
  INV_X1 U10726 ( .A(n8383), .ZN(n8367) );
  INV_X1 U10727 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10768) );
  INV_X1 U10728 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n8365) );
  NAND2_X1 U10729 ( .A1(n10768), .A2(n8365), .ZN(n8366) );
  NAND2_X1 U10730 ( .A1(n8367), .A2(n8366), .ZN(n11250) );
  INV_X1 U10731 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n8368) );
  OR2_X1 U10732 ( .A1(n6584), .A2(n8368), .ZN(n8369) );
  INV_X1 U10733 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10015) );
  NAND2_X1 U10734 ( .A1(n10013), .A2(n8477), .ZN(n8376) );
  INV_X1 U10735 ( .A(n8373), .ZN(n8389) );
  NAND2_X1 U10736 ( .A1(n8389), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8374) );
  XNOR2_X1 U10737 ( .A(n8374), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10098) );
  NAND2_X1 U10738 ( .A1(n8612), .A2(n10098), .ZN(n8375) );
  OAI211_X1 U10739 ( .C1(n8767), .C2(n10015), .A(n8376), .B(n8375), .ZN(n14789) );
  MUX2_X1 U10740 ( .A(n13896), .B(n14789), .S(n8775), .Z(n8377) );
  INV_X1 U10741 ( .A(n8377), .ZN(n8379) );
  MUX2_X1 U10742 ( .A(n14789), .B(n13896), .S(n8775), .Z(n8378) );
  OAI21_X1 U10743 ( .B1(n8380), .B2(n8379), .A(n8378), .ZN(n8382) );
  NAND2_X1 U10744 ( .A1(n8380), .A2(n8379), .ZN(n8381) );
  NAND2_X1 U10745 ( .A1(n8382), .A2(n8381), .ZN(n8394) );
  NAND2_X1 U10746 ( .A1(n8770), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8388) );
  INV_X1 U10747 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10083) );
  OR2_X1 U10748 ( .A1(n8713), .A2(n10083), .ZN(n8387) );
  NAND2_X1 U10749 ( .A1(n8383), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n8398) );
  OAI21_X1 U10750 ( .B1(n8383), .B2(P1_REG3_REG_5__SCAN_IN), .A(n8398), .ZN(
        n14720) );
  OR2_X1 U10751 ( .A1(n8701), .A2(n14720), .ZN(n8386) );
  INV_X1 U10752 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n8384) );
  OR2_X1 U10753 ( .A1(n8740), .A2(n8384), .ZN(n8385) );
  NAND4_X1 U10754 ( .A1(n8388), .A2(n8387), .A3(n8386), .A4(n8385), .ZN(n13895) );
  NAND2_X1 U10755 ( .A1(n10038), .A2(n8477), .ZN(n8392) );
  NAND2_X1 U10756 ( .A1(n8405), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8390) );
  XNOR2_X1 U10757 ( .A(n8390), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10100) );
  AOI22_X1 U10758 ( .A1(n8613), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8612), .B2(
        n10100), .ZN(n8391) );
  NAND2_X1 U10759 ( .A1(n8392), .A2(n8391), .ZN(n14723) );
  MUX2_X1 U10760 ( .A(n13895), .B(n14723), .S(n8780), .Z(n8395) );
  MUX2_X1 U10761 ( .A(n13895), .B(n14723), .S(n8775), .Z(n8393) );
  INV_X1 U10762 ( .A(n8395), .ZN(n8396) );
  NAND2_X1 U10763 ( .A1(n8770), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8404) );
  INV_X1 U10764 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11125) );
  OR2_X1 U10765 ( .A1(n8713), .A2(n11125), .ZN(n8403) );
  INV_X1 U10766 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n8397) );
  AND2_X1 U10767 ( .A1(n8398), .A2(n8397), .ZN(n8399) );
  NOR2_X1 U10768 ( .A1(n8398), .A2(n8397), .ZN(n8419) );
  OR2_X1 U10769 ( .A1(n8399), .A2(n8419), .ZN(n13873) );
  OR2_X1 U10770 ( .A1(n8701), .A2(n13873), .ZN(n8402) );
  INV_X1 U10771 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n8400) );
  OR2_X1 U10772 ( .A1(n8740), .A2(n8400), .ZN(n8401) );
  NAND4_X1 U10773 ( .A1(n8404), .A2(n8403), .A3(n8402), .A4(n8401), .ZN(n13894) );
  NAND2_X1 U10774 ( .A1(n10045), .A2(n8477), .ZN(n8410) );
  INV_X1 U10775 ( .A(n8405), .ZN(n8407) );
  INV_X1 U10776 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8406) );
  NAND2_X1 U10777 ( .A1(n8407), .A2(n8406), .ZN(n8426) );
  NAND2_X1 U10778 ( .A1(n8426), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8408) );
  XNOR2_X1 U10779 ( .A(n8408), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10102) );
  AOI22_X1 U10780 ( .A1(n8613), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8612), .B2(
        n10102), .ZN(n8409) );
  NAND2_X1 U10781 ( .A1(n8410), .A2(n8409), .ZN(n13872) );
  MUX2_X1 U10782 ( .A(n13894), .B(n13872), .S(n8775), .Z(n8414) );
  MUX2_X1 U10783 ( .A(n13894), .B(n13872), .S(n8544), .Z(n8411) );
  NAND2_X1 U10784 ( .A1(n8412), .A2(n8411), .ZN(n8418) );
  INV_X1 U10785 ( .A(n8413), .ZN(n8416) );
  INV_X1 U10786 ( .A(n8414), .ZN(n8415) );
  NAND2_X1 U10787 ( .A1(n8416), .A2(n8415), .ZN(n8417) );
  NAND2_X1 U10788 ( .A1(n8418), .A2(n8417), .ZN(n8433) );
  NAND2_X1 U10789 ( .A1(n8770), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8425) );
  INV_X1 U10790 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10084) );
  OR2_X1 U10791 ( .A1(n8713), .A2(n10084), .ZN(n8424) );
  NAND2_X1 U10792 ( .A1(n8419), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8447) );
  OR2_X1 U10793 ( .A1(n8419), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8420) );
  NAND2_X1 U10794 ( .A1(n8447), .A2(n8420), .ZN(n11403) );
  OR2_X1 U10795 ( .A1(n8701), .A2(n11403), .ZN(n8423) );
  INV_X1 U10796 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n8421) );
  OR2_X1 U10797 ( .A1(n8740), .A2(n8421), .ZN(n8422) );
  NAND4_X1 U10798 ( .A1(n8425), .A2(n8424), .A3(n8423), .A4(n8422), .ZN(n13893) );
  NAND2_X1 U10799 ( .A1(n10057), .A2(n8766), .ZN(n8431) );
  INV_X1 U10800 ( .A(n8426), .ZN(n8428) );
  INV_X1 U10801 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8427) );
  NAND2_X1 U10802 ( .A1(n8428), .A2(n8427), .ZN(n8436) );
  NAND2_X1 U10803 ( .A1(n8436), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8429) );
  XNOR2_X1 U10804 ( .A(n8429), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10131) );
  AOI22_X1 U10805 ( .A1(n8613), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8612), .B2(
        n10131), .ZN(n8430) );
  MUX2_X1 U10806 ( .A(n13893), .B(n11390), .S(n8544), .Z(n8434) );
  MUX2_X1 U10807 ( .A(n13893), .B(n11390), .S(n8775), .Z(n8432) );
  INV_X1 U10808 ( .A(n8434), .ZN(n8435) );
  NAND2_X1 U10809 ( .A1(n10074), .A2(n8766), .ZN(n8444) );
  NAND2_X1 U10810 ( .A1(n8438), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8437) );
  MUX2_X1 U10811 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8437), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n8441) );
  INV_X1 U10812 ( .A(n8438), .ZN(n8440) );
  INV_X1 U10813 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U10814 ( .A1(n8440), .A2(n8439), .ZN(n8463) );
  NAND2_X1 U10815 ( .A1(n8441), .A2(n8463), .ZN(n10145) );
  INV_X1 U10816 ( .A(n10145), .ZN(n8442) );
  AOI22_X1 U10817 ( .A1(n8613), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8612), .B2(
        n8442), .ZN(n8443) );
  NAND2_X1 U10818 ( .A1(n8444), .A2(n8443), .ZN(n11506) );
  NAND2_X1 U10819 ( .A1(n8770), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8452) );
  INV_X1 U10820 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n8445) );
  OR2_X1 U10821 ( .A1(n8713), .A2(n8445), .ZN(n8451) );
  NAND2_X1 U10822 ( .A1(n8447), .A2(n8446), .ZN(n8448) );
  NAND2_X1 U10823 ( .A1(n8457), .A2(n8448), .ZN(n11518) );
  OR2_X1 U10824 ( .A1(n8701), .A2(n11518), .ZN(n8450) );
  INV_X1 U10825 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10125) );
  OR2_X1 U10826 ( .A1(n8740), .A2(n10125), .ZN(n8449) );
  NAND2_X1 U10827 ( .A1(n11506), .A2(n11600), .ZN(n8793) );
  OR2_X1 U10828 ( .A1(n11506), .A2(n11600), .ZN(n11315) );
  MUX2_X1 U10829 ( .A(n8793), .B(n11315), .S(n8775), .Z(n8453) );
  INV_X1 U10830 ( .A(n11600), .ZN(n11505) );
  NOR2_X1 U10831 ( .A1(n11506), .A2(n11505), .ZN(n11328) );
  MUX2_X1 U10832 ( .A(n11505), .B(n11506), .S(n8544), .Z(n8454) );
  OR2_X1 U10833 ( .A1(n11328), .A2(n8454), .ZN(n8455) );
  NAND2_X1 U10834 ( .A1(n8770), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8462) );
  INV_X1 U10835 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10132) );
  OR2_X1 U10836 ( .A1(n8713), .A2(n10132), .ZN(n8461) );
  INV_X1 U10837 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10122) );
  OR2_X1 U10838 ( .A1(n8740), .A2(n10122), .ZN(n8460) );
  AND2_X1 U10839 ( .A1(n8457), .A2(n13580), .ZN(n8458) );
  OR2_X1 U10840 ( .A1(n8458), .A2(n8471), .ZN(n14703) );
  OR2_X1 U10841 ( .A1(n8701), .A2(n14703), .ZN(n8459) );
  NAND2_X1 U10842 ( .A1(n10078), .A2(n8766), .ZN(n8467) );
  NAND2_X1 U10843 ( .A1(n8463), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8494) );
  INV_X1 U10844 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8464) );
  NAND2_X1 U10845 ( .A1(n8494), .A2(n8464), .ZN(n8478) );
  OR2_X1 U10846 ( .A1(n8494), .A2(n8464), .ZN(n8465) );
  AOI22_X1 U10847 ( .A1(n8613), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8612), .B2(
        n10189), .ZN(n8466) );
  MUX2_X1 U10848 ( .A(n11598), .B(n14825), .S(n8544), .Z(n8469) );
  INV_X1 U10849 ( .A(n11598), .ZN(n11650) );
  MUX2_X1 U10850 ( .A(n11650), .B(n14705), .S(n8775), .Z(n8468) );
  NAND2_X1 U10851 ( .A1(n8770), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8476) );
  INV_X1 U10852 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n8470) );
  OR2_X1 U10853 ( .A1(n8713), .A2(n8470), .ZN(n8475) );
  NOR2_X1 U10854 ( .A1(n8471), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8472) );
  OR2_X1 U10855 ( .A1(n8485), .A2(n8472), .ZN(n11645) );
  OR2_X1 U10856 ( .A1(n8701), .A2(n11645), .ZN(n8474) );
  INV_X1 U10857 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10188) );
  OR2_X1 U10858 ( .A1(n8740), .A2(n10188), .ZN(n8473) );
  NAND4_X1 U10859 ( .A1(n8476), .A2(n8475), .A3(n8474), .A4(n8473), .ZN(n13892) );
  NAND2_X1 U10860 ( .A1(n10157), .A2(n8766), .ZN(n8481) );
  NAND2_X1 U10861 ( .A1(n8478), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8479) );
  XNOR2_X1 U10862 ( .A(n8479), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10240) );
  AOI22_X1 U10863 ( .A1(n8613), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8612), 
        .B2(n10240), .ZN(n8480) );
  MUX2_X1 U10864 ( .A(n13892), .B(n14834), .S(n8775), .Z(n8483) );
  MUX2_X1 U10865 ( .A(n13892), .B(n14834), .S(n8544), .Z(n8482) );
  NAND2_X1 U10866 ( .A1(n6588), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8491) );
  NAND2_X1 U10867 ( .A1(n8485), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8506) );
  OR2_X1 U10868 ( .A1(n8485), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8486) );
  NAND2_X1 U10869 ( .A1(n8506), .A2(n8486), .ZN(n14540) );
  OR2_X1 U10870 ( .A1(n8701), .A2(n14540), .ZN(n8490) );
  INV_X1 U10871 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10243) );
  OR2_X1 U10872 ( .A1(n8740), .A2(n10243), .ZN(n8489) );
  INV_X1 U10873 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n8487) );
  OR2_X1 U10874 ( .A1(n6583), .A2(n8487), .ZN(n8488) );
  NAND4_X1 U10875 ( .A1(n8491), .A2(n8490), .A3(n8489), .A4(n8488), .ZN(n13891) );
  NAND2_X1 U10876 ( .A1(n10198), .A2(n8766), .ZN(n8497) );
  OR2_X1 U10877 ( .A1(n8492), .A2(n8592), .ZN(n8493) );
  NAND2_X1 U10878 ( .A1(n8494), .A2(n8493), .ZN(n8512) );
  INV_X1 U10879 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8495) );
  XNOR2_X1 U10880 ( .A(n8512), .B(n8495), .ZN(n10372) );
  AOI22_X1 U10881 ( .A1(n8613), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8612), 
        .B2(n10372), .ZN(n8496) );
  MUX2_X1 U10882 ( .A(n13891), .B(n14537), .S(n8780), .Z(n8501) );
  MUX2_X1 U10883 ( .A(n13891), .B(n14537), .S(n8775), .Z(n8498) );
  NAND2_X1 U10884 ( .A1(n8499), .A2(n8498), .ZN(n8505) );
  INV_X1 U10885 ( .A(n8500), .ZN(n8503) );
  INV_X1 U10886 ( .A(n8501), .ZN(n8502) );
  NAND2_X1 U10887 ( .A1(n8503), .A2(n8502), .ZN(n8504) );
  NAND2_X1 U10888 ( .A1(n8505), .A2(n8504), .ZN(n8517) );
  NAND2_X1 U10889 ( .A1(n8770), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8511) );
  INV_X1 U10890 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10362) );
  OR2_X1 U10891 ( .A1(n8713), .A2(n10362), .ZN(n8510) );
  NAND2_X1 U10892 ( .A1(n8506), .A2(n10368), .ZN(n8507) );
  NAND2_X1 U10893 ( .A1(n8532), .A2(n8507), .ZN(n11806) );
  OR2_X1 U10894 ( .A1(n8701), .A2(n11806), .ZN(n8509) );
  INV_X1 U10895 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10371) );
  OR2_X1 U10896 ( .A1(n8740), .A2(n10371), .ZN(n8508) );
  NAND4_X1 U10897 ( .A1(n8511), .A2(n8510), .A3(n8509), .A4(n8508), .ZN(n13890) );
  NAND2_X1 U10898 ( .A1(n10311), .A2(n8766), .ZN(n8515) );
  NAND2_X1 U10899 ( .A1(n8513), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8520) );
  XNOR2_X1 U10900 ( .A(n8520), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U10901 ( .A1(n8613), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n10607), 
        .B2(n8612), .ZN(n8514) );
  MUX2_X1 U10902 ( .A(n13890), .B(n11799), .S(n8775), .Z(n8518) );
  MUX2_X1 U10903 ( .A(n13890), .B(n11799), .S(n8780), .Z(n8516) );
  NAND2_X1 U10904 ( .A1(n10413), .A2(n8766), .ZN(n8524) );
  INV_X1 U10905 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8519) );
  NAND2_X1 U10906 ( .A1(n8520), .A2(n8519), .ZN(n8521) );
  NAND2_X1 U10907 ( .A1(n8521), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8539) );
  NAND2_X1 U10908 ( .A1(n8539), .A2(n13671), .ZN(n8541) );
  NAND2_X1 U10909 ( .A1(n8541), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8522) );
  AOI22_X1 U10910 ( .A1(n11281), .A2(n8612), .B1(n8613), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U10911 ( .A1(n8770), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8531) );
  AND2_X1 U10912 ( .A1(n8534), .A2(n8525), .ZN(n8526) );
  OR2_X1 U10913 ( .A1(n8526), .A2(n8549), .ZN(n14504) );
  OR2_X1 U10914 ( .A1(n14504), .A2(n8701), .ZN(n8530) );
  INV_X1 U10915 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8527) );
  OR2_X1 U10916 ( .A1(n8740), .A2(n8527), .ZN(n8529) );
  INV_X1 U10917 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11682) );
  OR2_X1 U10918 ( .A1(n8713), .A2(n11682), .ZN(n8528) );
  XNOR2_X1 U10919 ( .A(n14598), .B(n14544), .ZN(n11687) );
  NAND2_X1 U10920 ( .A1(n8770), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8538) );
  INV_X1 U10921 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11540) );
  OR2_X1 U10922 ( .A1(n8713), .A2(n11540), .ZN(n8537) );
  NAND2_X1 U10923 ( .A1(n8532), .A2(n13746), .ZN(n8533) );
  NAND2_X1 U10924 ( .A1(n8534), .A2(n8533), .ZN(n13845) );
  OR2_X1 U10925 ( .A1(n8701), .A2(n13845), .ZN(n8536) );
  INV_X1 U10926 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10606) );
  OR2_X1 U10927 ( .A1(n8740), .A2(n10606), .ZN(n8535) );
  NAND2_X1 U10928 ( .A1(n10318), .A2(n8766), .ZN(n8543) );
  OR2_X1 U10929 ( .A1(n8539), .A2(n13671), .ZN(n8540) );
  AOI22_X1 U10930 ( .A1(n10688), .A2(n8612), .B1(n8613), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n8542) );
  MUX2_X1 U10931 ( .A(n14494), .B(n11973), .S(n8780), .Z(n8559) );
  NAND2_X1 U10932 ( .A1(n11687), .A2(n8559), .ZN(n8557) );
  NAND2_X1 U10933 ( .A1(n10716), .A2(n8766), .ZN(n8548) );
  NAND2_X1 U10934 ( .A1(n8545), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8546) );
  XNOR2_X1 U10935 ( .A(n8546), .B(P1_IR_REG_15__SCAN_IN), .ZN(n14686) );
  AOI22_X1 U10936 ( .A1(n8613), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8612), 
        .B2(n14686), .ZN(n8547) );
  NAND2_X1 U10937 ( .A1(n6588), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8556) );
  NAND2_X1 U10938 ( .A1(n8549), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8573) );
  OR2_X1 U10939 ( .A1(n8549), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8550) );
  NAND2_X1 U10940 ( .A1(n8573), .A2(n8550), .ZN(n14574) );
  OR2_X1 U10941 ( .A1(n14574), .A2(n8701), .ZN(n8555) );
  INV_X1 U10942 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8551) );
  OR2_X1 U10943 ( .A1(n8740), .A2(n8551), .ZN(n8554) );
  INV_X1 U10944 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n8552) );
  OR2_X1 U10945 ( .A1(n6583), .A2(n8552), .ZN(n8553) );
  OR2_X1 U10946 ( .A1(n14598), .A2(n14556), .ZN(n11912) );
  NAND2_X1 U10947 ( .A1(n14592), .A2(n14493), .ZN(n8790) );
  NAND2_X1 U10948 ( .A1(n8558), .A2(n8790), .ZN(n8568) );
  INV_X1 U10949 ( .A(n8559), .ZN(n8560) );
  NAND2_X1 U10950 ( .A1(n8561), .A2(n8560), .ZN(n8566) );
  INV_X1 U10951 ( .A(n14494), .ZN(n11674) );
  NAND2_X1 U10952 ( .A1(n8790), .A2(n11674), .ZN(n8562) );
  MUX2_X1 U10953 ( .A(n11973), .B(n8562), .S(n8780), .Z(n8563) );
  NOR2_X1 U10954 ( .A1(n8563), .A2(n11686), .ZN(n8565) );
  NAND2_X1 U10955 ( .A1(n14598), .A2(n14556), .ZN(n11910) );
  AOI21_X1 U10956 ( .B1(n8790), .B2(n11910), .A(n8780), .ZN(n8564) );
  AOI21_X1 U10957 ( .B1(n8566), .B2(n8565), .A(n8564), .ZN(n8567) );
  NAND2_X1 U10958 ( .A1(n8568), .A2(n8567), .ZN(n8569) );
  INV_X1 U10959 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n8571) );
  NAND2_X1 U10960 ( .A1(n8363), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8570) );
  OAI21_X1 U10961 ( .B1(n6584), .B2(n8571), .A(n8570), .ZN(n8577) );
  INV_X1 U10962 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8572) );
  NAND2_X1 U10963 ( .A1(n8573), .A2(n8572), .ZN(n8574) );
  NAND2_X1 U10964 ( .A1(n8597), .A2(n8574), .ZN(n14514) );
  INV_X1 U10965 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11296) );
  OR2_X1 U10966 ( .A1(n8713), .A2(n11296), .ZN(n8575) );
  OAI21_X1 U10967 ( .B1(n8701), .B2(n14514), .A(n8575), .ZN(n8576) );
  NAND2_X1 U10968 ( .A1(n10772), .A2(n8766), .ZN(n8581) );
  NAND2_X1 U10969 ( .A1(n8578), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8579) );
  XNOR2_X1 U10970 ( .A(n8579), .B(P1_IR_REG_16__SCAN_IN), .ZN(n13937) );
  AOI22_X1 U10971 ( .A1(n8613), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8612), 
        .B2(n13937), .ZN(n8580) );
  MUX2_X1 U10972 ( .A(n14546), .B(n14184), .S(n8780), .Z(n8583) );
  MUX2_X1 U10973 ( .A(n14546), .B(n14184), .S(n8775), .Z(n8582) );
  INV_X1 U10974 ( .A(n8583), .ZN(n8584) );
  NOR2_X1 U10975 ( .A1(n8598), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8585) );
  OR2_X1 U10976 ( .A1(n8616), .A2(n8585), .ZN(n14149) );
  AOI22_X1 U10977 ( .A1(n6588), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n8770), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n8587) );
  INV_X1 U10978 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n13963) );
  OR2_X1 U10979 ( .A1(n8740), .A2(n13963), .ZN(n8586) );
  OAI211_X1 U10980 ( .C1(n14149), .C2(n8701), .A(n8587), .B(n8586), .ZN(n14159) );
  NAND2_X1 U10981 ( .A1(n11131), .A2(n8766), .ZN(n8591) );
  NAND2_X1 U10982 ( .A1(n8588), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8589) );
  XNOR2_X1 U10983 ( .A(n8589), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13976) );
  AOI22_X1 U10984 ( .A1(n8613), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8612), 
        .B2(n13976), .ZN(n8590) );
  MUX2_X1 U10985 ( .A(n14159), .B(n14265), .S(n8775), .Z(n8603) );
  NAND2_X1 U10986 ( .A1(n14265), .A2(n14159), .ZN(n11895) );
  NAND2_X1 U10987 ( .A1(n8603), .A2(n11895), .ZN(n8602) );
  NAND2_X1 U10988 ( .A1(n10892), .A2(n8766), .ZN(n8596) );
  OR2_X1 U10989 ( .A1(n8593), .A2(n8592), .ZN(n8594) );
  XNOR2_X1 U10990 ( .A(n8594), .B(P1_IR_REG_17__SCAN_IN), .ZN(n13961) );
  AOI22_X1 U10991 ( .A1(n8613), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8612), 
        .B2(n13961), .ZN(n8595) );
  AND2_X1 U10992 ( .A1(n8597), .A2(n13944), .ZN(n8599) );
  OR2_X1 U10993 ( .A1(n8599), .A2(n8598), .ZN(n14523) );
  AOI22_X1 U10994 ( .A1(n6588), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n8770), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n8601) );
  INV_X1 U10995 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n13938) );
  OR2_X1 U10996 ( .A1(n8740), .A2(n13938), .ZN(n8600) );
  OAI211_X2 U10997 ( .C1(n14523), .C2(n8701), .A(n8601), .B(n8600), .ZN(n14508) );
  XNOR2_X1 U10998 ( .A(n14575), .B(n14508), .ZN(n11916) );
  INV_X1 U10999 ( .A(n8603), .ZN(n8611) );
  OR2_X1 U11000 ( .A1(n14265), .A2(n14159), .ZN(n11894) );
  AND2_X1 U11001 ( .A1(n14508), .A2(n8775), .ZN(n8605) );
  NOR2_X1 U11002 ( .A1(n14508), .A2(n8775), .ZN(n8606) );
  MUX2_X1 U11003 ( .A(n8605), .B(n8606), .S(n14575), .Z(n8604) );
  OR2_X1 U11004 ( .A1(n11894), .A2(n8604), .ZN(n8610) );
  INV_X1 U11005 ( .A(n8605), .ZN(n8608) );
  NAND2_X1 U11006 ( .A1(n14575), .A2(n8606), .ZN(n8607) );
  OAI21_X1 U11007 ( .B1(n14575), .B2(n8608), .A(n8607), .ZN(n8609) );
  AOI22_X1 U11008 ( .A1(n8611), .A2(n8610), .B1(n7390), .B2(n8609), .ZN(n8620)
         );
  NAND2_X1 U11009 ( .A1(n11191), .A2(n8766), .ZN(n8615) );
  AOI22_X1 U11010 ( .A1(n8613), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10937), 
        .B2(n8612), .ZN(n8614) );
  NAND2_X1 U11011 ( .A1(n8616), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8627) );
  OR2_X1 U11012 ( .A1(n8616), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8617) );
  NAND2_X1 U11013 ( .A1(n8627), .A2(n8617), .ZN(n14137) );
  AOI22_X1 U11014 ( .A1(n6588), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n8770), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n8619) );
  INV_X1 U11015 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13973) );
  OR2_X1 U11016 ( .A1(n8740), .A2(n13973), .ZN(n8618) );
  XNOR2_X1 U11017 ( .A(n14260), .B(n14146), .ZN(n14132) );
  NAND2_X1 U11018 ( .A1(n8622), .A2(n8621), .ZN(n8626) );
  NAND2_X1 U11019 ( .A1(n14146), .A2(n8780), .ZN(n8624) );
  OR2_X1 U11020 ( .A1(n14146), .A2(n8780), .ZN(n8623) );
  MUX2_X1 U11021 ( .A(n8624), .B(n8623), .S(n14260), .Z(n8625) );
  INV_X1 U11022 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13834) );
  NAND2_X1 U11023 ( .A1(n8627), .A2(n13834), .ZN(n8629) );
  INV_X1 U11024 ( .A(n8641), .ZN(n8628) );
  NAND2_X1 U11025 ( .A1(n8629), .A2(n8628), .ZN(n13832) );
  OR2_X1 U11026 ( .A1(n13832), .A2(n8701), .ZN(n8635) );
  INV_X1 U11027 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n8632) );
  NAND2_X1 U11028 ( .A1(n8770), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8631) );
  NAND2_X1 U11029 ( .A1(n8363), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8630) );
  OAI211_X1 U11030 ( .C1(n8713), .C2(n8632), .A(n8631), .B(n8630), .ZN(n8633)
         );
  INV_X1 U11031 ( .A(n8633), .ZN(n8634) );
  NAND2_X1 U11032 ( .A1(n11260), .A2(n8766), .ZN(n8637) );
  OR2_X1 U11033 ( .A1(n8767), .A2(n7027), .ZN(n8636) );
  AND2_X2 U11034 ( .A1(n8637), .A2(n8636), .ZN(n14252) );
  MUX2_X1 U11035 ( .A(n13799), .B(n14252), .S(n8780), .Z(n8639) );
  MUX2_X1 U11036 ( .A(n14107), .B(n14125), .S(n8775), .Z(n8638) );
  NAND2_X1 U11037 ( .A1(n6588), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8645) );
  INV_X1 U11038 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8640) );
  OR2_X1 U11039 ( .A1(n8740), .A2(n8640), .ZN(n8644) );
  INV_X1 U11040 ( .A(n8659), .ZN(n8661) );
  OAI21_X1 U11041 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n8641), .A(n8661), .ZN(
        n14109) );
  OR2_X1 U11042 ( .A1(n8701), .A2(n14109), .ZN(n8643) );
  INV_X1 U11043 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n13690) );
  OR2_X1 U11044 ( .A1(n6584), .A2(n13690), .ZN(n8642) );
  NAND4_X1 U11045 ( .A1(n8645), .A2(n8644), .A3(n8643), .A4(n8642), .ZN(n13889) );
  OR2_X1 U11046 ( .A1(n11372), .A2(n8683), .ZN(n8647) );
  INV_X1 U11047 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11359) );
  OR2_X1 U11048 ( .A1(n8767), .A2(n11359), .ZN(n8646) );
  MUX2_X1 U11049 ( .A(n13889), .B(n14246), .S(n8775), .Z(n8651) );
  NAND2_X1 U11050 ( .A1(n8650), .A2(n8651), .ZN(n8649) );
  MUX2_X1 U11051 ( .A(n13889), .B(n14246), .S(n8780), .Z(n8648) );
  INV_X1 U11052 ( .A(n8651), .ZN(n8652) );
  NAND2_X1 U11053 ( .A1(n8653), .A2(n8652), .ZN(n8654) );
  NAND2_X1 U11054 ( .A1(n6588), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8667) );
  INV_X1 U11055 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n8658) );
  OR2_X1 U11056 ( .A1(n6583), .A2(n8658), .ZN(n8666) );
  INV_X1 U11057 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8660) );
  NAND2_X1 U11058 ( .A1(n8661), .A2(n8660), .ZN(n8662) );
  NAND2_X1 U11059 ( .A1(n8689), .A2(n8662), .ZN(n14096) );
  OR2_X1 U11060 ( .A1(n8701), .A2(n14096), .ZN(n8665) );
  INV_X1 U11061 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8663) );
  OR2_X1 U11062 ( .A1(n8740), .A2(n8663), .ZN(n8664) );
  MUX2_X1 U11063 ( .A(n14101), .B(n13788), .S(n8775), .Z(n8668) );
  INV_X1 U11064 ( .A(n8668), .ZN(n8669) );
  NAND2_X1 U11065 ( .A1(n6588), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8673) );
  INV_X1 U11066 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n13620) );
  OR2_X1 U11067 ( .A1(n6584), .A2(n13620), .ZN(n8672) );
  INV_X1 U11068 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8687) );
  XNOR2_X1 U11069 ( .A(n8689), .B(n8687), .ZN(n14081) );
  OR2_X1 U11070 ( .A1(n8701), .A2(n14081), .ZN(n8671) );
  INV_X1 U11071 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n13730) );
  OR2_X1 U11072 ( .A1(n8740), .A2(n13730), .ZN(n8670) );
  NAND4_X1 U11073 ( .A1(n8673), .A2(n8672), .A3(n8671), .A4(n8670), .ZN(n14059) );
  NAND2_X1 U11074 ( .A1(n11614), .A2(n8766), .ZN(n8675) );
  INV_X1 U11075 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11617) );
  OR2_X1 U11076 ( .A1(n8767), .A2(n11617), .ZN(n8674) );
  MUX2_X1 U11077 ( .A(n14059), .B(n14235), .S(n8775), .Z(n8679) );
  MUX2_X1 U11078 ( .A(n14235), .B(n14059), .S(n8775), .Z(n8676) );
  AOI21_X1 U11079 ( .B1(n8680), .B2(n8679), .A(n8677), .ZN(n8678) );
  INV_X1 U11080 ( .A(n8678), .ZN(n8682) );
  OR2_X1 U11081 ( .A1(n11697), .A2(n8683), .ZN(n8685) );
  INV_X1 U11082 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11694) );
  OR2_X1 U11083 ( .A1(n8767), .A2(n11694), .ZN(n8684) );
  NAND2_X1 U11084 ( .A1(n8770), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8695) );
  INV_X1 U11085 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14064) );
  OR2_X1 U11086 ( .A1(n8713), .A2(n14064), .ZN(n8694) );
  INV_X1 U11087 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8686) );
  OAI21_X1 U11088 ( .B1(n8689), .B2(n8687), .A(n8686), .ZN(n8691) );
  NAND2_X1 U11089 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n8688) );
  INV_X1 U11090 ( .A(n8699), .ZN(n8690) );
  NAND2_X1 U11091 ( .A1(n8691), .A2(n8690), .ZN(n14063) );
  OR2_X1 U11092 ( .A1(n8701), .A2(n14063), .ZN(n8693) );
  INV_X1 U11093 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n14231) );
  OR2_X1 U11094 ( .A1(n8740), .A2(n14231), .ZN(n8692) );
  NAND4_X1 U11095 ( .A1(n8695), .A2(n8694), .A3(n8693), .A4(n8692), .ZN(n13888) );
  MUX2_X1 U11096 ( .A(n14068), .B(n13888), .S(n8775), .Z(n8697) );
  MUX2_X1 U11097 ( .A(n13888), .B(n14068), .S(n8775), .Z(n8696) );
  NAND2_X1 U11098 ( .A1(n8770), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8706) );
  INV_X1 U11099 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n8698) );
  OR2_X1 U11100 ( .A1(n8713), .A2(n8698), .ZN(n8705) );
  NOR2_X1 U11101 ( .A1(n8699), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8700) );
  OR2_X1 U11102 ( .A1(n8714), .A2(n8700), .ZN(n14045) );
  OR2_X1 U11103 ( .A1(n8701), .A2(n14045), .ZN(n8704) );
  INV_X1 U11104 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n8702) );
  OR2_X1 U11105 ( .A1(n8740), .A2(n8702), .ZN(n8703) );
  NAND4_X1 U11106 ( .A1(n8706), .A2(n8705), .A3(n8704), .A4(n8703), .ZN(n14058) );
  NAND2_X1 U11107 ( .A1(n13772), .A2(n8766), .ZN(n8708) );
  INV_X1 U11108 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14302) );
  OR2_X1 U11109 ( .A1(n8767), .A2(n14302), .ZN(n8707) );
  MUX2_X1 U11110 ( .A(n14058), .B(n14221), .S(n8775), .Z(n8711) );
  MUX2_X1 U11111 ( .A(n14058), .B(n14221), .S(n8780), .Z(n8709) );
  NAND2_X1 U11112 ( .A1(n8363), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8719) );
  INV_X1 U11113 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n8712) );
  OR2_X1 U11114 ( .A1(n8713), .A2(n8712), .ZN(n8718) );
  INV_X1 U11115 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n13649) );
  OR2_X1 U11116 ( .A1(n6583), .A2(n13649), .ZN(n8717) );
  OR2_X1 U11117 ( .A1(n8714), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U11118 ( .A1(n8714), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8726) );
  NAND2_X1 U11119 ( .A1(n8715), .A2(n8726), .ZN(n14031) );
  OR2_X1 U11120 ( .A1(n8701), .A2(n14031), .ZN(n8716) );
  NAND4_X1 U11121 ( .A1(n8719), .A2(n8718), .A3(n8717), .A4(n8716), .ZN(n14012) );
  NAND2_X1 U11122 ( .A1(n14297), .A2(n8766), .ZN(n8721) );
  OR2_X1 U11123 ( .A1(n8767), .A2(n14299), .ZN(n8720) );
  MUX2_X1 U11124 ( .A(n14012), .B(n14214), .S(n8780), .Z(n8724) );
  MUX2_X1 U11125 ( .A(n14012), .B(n14214), .S(n8775), .Z(n8722) );
  INV_X1 U11126 ( .A(n8724), .ZN(n8725) );
  NAND2_X1 U11127 ( .A1(n6588), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8732) );
  INV_X1 U11128 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n13678) );
  OR2_X1 U11129 ( .A1(n6584), .A2(n13678), .ZN(n8731) );
  INV_X1 U11130 ( .A(n8726), .ZN(n8727) );
  NAND2_X1 U11131 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n8727), .ZN(n8751) );
  OAI21_X1 U11132 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(n8727), .A(n8751), .ZN(
        n14015) );
  OR2_X1 U11133 ( .A1(n8701), .A2(n14015), .ZN(n8730) );
  INV_X1 U11134 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8728) );
  OR2_X1 U11135 ( .A1(n8740), .A2(n8728), .ZN(n8729) );
  NAND2_X1 U11136 ( .A1(n14293), .A2(n8766), .ZN(n8734) );
  OR2_X1 U11137 ( .A1(n8767), .A2(n14296), .ZN(n8733) );
  MUX2_X1 U11138 ( .A(n13887), .B(n14020), .S(n8775), .Z(n8736) );
  MUX2_X1 U11139 ( .A(n14020), .B(n13887), .S(n8775), .Z(n8735) );
  INV_X1 U11140 ( .A(n8736), .ZN(n8737) );
  NAND2_X1 U11141 ( .A1(n6588), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8744) );
  INV_X1 U11142 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n13608) );
  OR2_X1 U11143 ( .A1(n6583), .A2(n13608), .ZN(n8743) );
  INV_X1 U11144 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8738) );
  XNOR2_X1 U11145 ( .A(n8751), .B(n8738), .ZN(n12086) );
  OR2_X1 U11146 ( .A1(n8701), .A2(n12086), .ZN(n8742) );
  INV_X1 U11147 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8739) );
  OR2_X1 U11148 ( .A1(n8740), .A2(n8739), .ZN(n8741) );
  NAND4_X1 U11149 ( .A1(n8744), .A2(n8743), .A3(n8742), .A4(n8741), .ZN(n14011) );
  NAND2_X1 U11150 ( .A1(n11876), .A2(n8766), .ZN(n8746) );
  OR2_X1 U11151 ( .A1(n8767), .A2(n11877), .ZN(n8745) );
  MUX2_X1 U11152 ( .A(n14011), .B(n14203), .S(n8780), .Z(n8748) );
  MUX2_X1 U11153 ( .A(n14011), .B(n14203), .S(n8775), .Z(n8747) );
  INV_X1 U11154 ( .A(n8748), .ZN(n8749) );
  NAND2_X1 U11155 ( .A1(n6588), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8757) );
  INV_X1 U11156 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8750) );
  OR2_X1 U11157 ( .A1(n6583), .A2(n8750), .ZN(n8756) );
  INV_X1 U11158 ( .A(n8751), .ZN(n8752) );
  NAND2_X1 U11159 ( .A1(n8752), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n11940) );
  OR2_X1 U11160 ( .A1(n8701), .A2(n11940), .ZN(n8755) );
  INV_X1 U11161 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8753) );
  OR2_X1 U11162 ( .A1(n8740), .A2(n8753), .ZN(n8754) );
  NAND4_X1 U11163 ( .A1(n8757), .A2(n8756), .A3(n8755), .A4(n8754), .ZN(n13886) );
  NAND2_X1 U11164 ( .A1(n11864), .A2(n8766), .ZN(n8759) );
  OR2_X1 U11165 ( .A1(n8767), .A2(n6778), .ZN(n8758) );
  MUX2_X1 U11166 ( .A(n13886), .B(n11937), .S(n8775), .Z(n8761) );
  MUX2_X1 U11167 ( .A(n13886), .B(n11937), .S(n8780), .Z(n8760) );
  NAND2_X1 U11168 ( .A1(n8763), .A2(n8762), .ZN(n8764) );
  NAND2_X1 U11169 ( .A1(n11874), .A2(n8766), .ZN(n8769) );
  INV_X1 U11170 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12313) );
  OR2_X1 U11171 ( .A1(n8767), .A2(n12313), .ZN(n8768) );
  INV_X1 U11172 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n13706) );
  NAND2_X1 U11173 ( .A1(n6588), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8772) );
  NAND2_X1 U11174 ( .A1(n8770), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8771) );
  OAI211_X1 U11175 ( .C1(n8740), .C2(n13706), .A(n8772), .B(n8771), .ZN(n13885) );
  OAI21_X1 U11176 ( .B1(n13994), .B2(n11261), .A(n13885), .ZN(n8773) );
  INV_X1 U11177 ( .A(n8773), .ZN(n8774) );
  MUX2_X1 U11178 ( .A(n13998), .B(n8774), .S(n8780), .Z(n8782) );
  NAND2_X1 U11179 ( .A1(n13994), .A2(n8775), .ZN(n8776) );
  OAI21_X1 U11180 ( .B1(n10790), .B2(n8777), .A(n8776), .ZN(n8778) );
  AND2_X1 U11181 ( .A1(n8778), .A2(n13885), .ZN(n8779) );
  AOI21_X1 U11182 ( .B1(n13998), .B2(n8780), .A(n8779), .ZN(n8781) );
  NAND2_X1 U11183 ( .A1(n8782), .A2(n8781), .ZN(n8784) );
  NOR2_X1 U11184 ( .A1(n8782), .A2(n8781), .ZN(n8783) );
  AOI21_X1 U11185 ( .B1(n8785), .B2(n8784), .A(n8783), .ZN(n8818) );
  XOR2_X1 U11186 ( .A(n13994), .B(n13996), .Z(n8815) );
  XNOR2_X1 U11187 ( .A(n13998), .B(n13885), .ZN(n8802) );
  INV_X1 U11188 ( .A(n14011), .ZN(n8786) );
  NAND2_X1 U11189 ( .A1(n14203), .A2(n8786), .ZN(n11934) );
  NAND2_X1 U11190 ( .A1(n11934), .A2(n8787), .ZN(n11909) );
  INV_X1 U11191 ( .A(n14058), .ZN(n13880) );
  XNOR2_X1 U11192 ( .A(n14221), .B(n13880), .ZN(n14041) );
  INV_X1 U11193 ( .A(n14012), .ZN(n8788) );
  NAND2_X1 U11194 ( .A1(n14214), .A2(n8788), .ZN(n11933) );
  OR2_X1 U11195 ( .A1(n14214), .A2(n8788), .ZN(n8789) );
  NAND2_X1 U11196 ( .A1(n11933), .A2(n8789), .ZN(n14023) );
  XNOR2_X1 U11197 ( .A(n14068), .B(n13888), .ZN(n11901) );
  XNOR2_X1 U11198 ( .A(n14101), .B(n13788), .ZN(n14088) );
  INV_X1 U11199 ( .A(n13889), .ZN(n11924) );
  XNOR2_X1 U11200 ( .A(n14246), .B(n11924), .ZN(n14113) );
  XNOR2_X1 U11201 ( .A(n14125), .B(n13799), .ZN(n14118) );
  NAND2_X1 U11202 ( .A1(n11894), .A2(n11895), .ZN(n14152) );
  NAND2_X1 U11203 ( .A1(n11915), .A2(n8790), .ZN(n14567) );
  XNOR2_X1 U11204 ( .A(n13847), .B(n14494), .ZN(n11536) );
  XNOR2_X1 U11205 ( .A(n11799), .B(n13890), .ZN(n11575) );
  XNOR2_X1 U11206 ( .A(n14705), .B(n11598), .ZN(n14698) );
  INV_X1 U11207 ( .A(n14733), .ZN(n10785) );
  XNOR2_X1 U11208 ( .A(n10266), .B(n10953), .ZN(n14761) );
  NOR4_X1 U11209 ( .A1(n10785), .A2(n14761), .A3(n10958), .A4(n10936), .ZN(
        n8791) );
  XNOR2_X1 U11210 ( .A(n13872), .B(n13894), .ZN(n11096) );
  XNOR2_X1 U11211 ( .A(n13895), .B(n14723), .ZN(n11107) );
  XNOR2_X1 U11212 ( .A(n13896), .B(n14789), .ZN(n11102) );
  NAND4_X1 U11213 ( .A1(n8791), .A2(n11096), .A3(n11107), .A4(n11102), .ZN(
        n8794) );
  INV_X1 U11214 ( .A(n13893), .ZN(n8792) );
  XNOR2_X1 U11215 ( .A(n11390), .B(n8792), .ZN(n11272) );
  NAND2_X1 U11216 ( .A1(n11315), .A2(n8793), .ZN(n11326) );
  NOR4_X1 U11217 ( .A1(n14698), .A2(n8794), .A3(n11272), .A4(n11326), .ZN(
        n8795) );
  XNOR2_X1 U11218 ( .A(n14834), .B(n13892), .ZN(n11318) );
  OR2_X1 U11219 ( .A1(n14537), .A2(n13891), .ZN(n11532) );
  NAND2_X1 U11220 ( .A1(n14537), .A2(n13891), .ZN(n11535) );
  NAND2_X1 U11221 ( .A1(n11532), .A2(n11535), .ZN(n11416) );
  NAND4_X1 U11222 ( .A1(n11575), .A2(n8795), .A3(n11318), .A4(n11416), .ZN(
        n8796) );
  NOR4_X1 U11223 ( .A1(n14567), .A2(n11686), .A3(n11536), .A4(n8796), .ZN(
        n8797) );
  XNOR2_X1 U11224 ( .A(n14184), .B(n14546), .ZN(n14171) );
  NAND4_X1 U11225 ( .A1(n14152), .A2(n8797), .A3(n11916), .A4(n14171), .ZN(
        n8798) );
  NOR4_X1 U11226 ( .A1(n14113), .A2(n14118), .A3(n14129), .A4(n8798), .ZN(
        n8799) );
  XNOR2_X1 U11227 ( .A(n14235), .B(n14059), .ZN(n14077) );
  NAND4_X1 U11228 ( .A1(n11901), .A2(n14088), .A3(n8799), .A4(n14077), .ZN(
        n8800) );
  NOR4_X1 U11229 ( .A1(n11909), .A2(n14041), .A3(n14023), .A4(n8800), .ZN(
        n8801) );
  XNOR2_X1 U11230 ( .A(n11937), .B(n13886), .ZN(n11935) );
  XNOR2_X1 U11231 ( .A(n14020), .B(n13887), .ZN(n14007) );
  NAND4_X1 U11232 ( .A1(n8802), .A2(n8801), .A3(n11935), .A4(n14007), .ZN(
        n8803) );
  NOR2_X1 U11233 ( .A1(n8815), .A2(n8803), .ZN(n8804) );
  XOR2_X1 U11234 ( .A(n13984), .B(n8804), .Z(n8813) );
  NOR3_X1 U11235 ( .A1(n14191), .A2(n13994), .A3(n8805), .ZN(n8808) );
  NOR3_X1 U11236 ( .A1(n8807), .A2(n13994), .A3(n8814), .ZN(n8806) );
  AOI21_X1 U11237 ( .B1(n8808), .B2(n8807), .A(n8806), .ZN(n8812) );
  XOR2_X1 U11238 ( .A(n8814), .B(n8809), .Z(n8810) );
  NAND4_X1 U11239 ( .A1(n8810), .A2(n14191), .A3(n13994), .A4(n10290), .ZN(
        n8811) );
  OAI211_X1 U11240 ( .C1(n8813), .C2(n10290), .A(n8812), .B(n8811), .ZN(n8817)
         );
  NOR3_X1 U11241 ( .A1(n8818), .A2(n8815), .A3(n8814), .ZN(n8816) );
  AOI211_X1 U11242 ( .C1(n8819), .C2(n8818), .A(n8817), .B(n8816), .ZN(n8839)
         );
  NAND2_X1 U11243 ( .A1(n6662), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8820) );
  INV_X1 U11244 ( .A(n10062), .ZN(n8821) );
  NAND2_X1 U11245 ( .A1(n8821), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11615) );
  NAND2_X1 U11246 ( .A1(n8825), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8827) );
  NAND2_X1 U11247 ( .A1(n8828), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8829) );
  MUX2_X1 U11248 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8829), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8830) );
  INV_X1 U11249 ( .A(n8832), .ZN(n10296) );
  NAND2_X1 U11250 ( .A1(n13984), .A2(n11261), .ZN(n8833) );
  NAND2_X1 U11251 ( .A1(n10296), .A2(n8833), .ZN(n10294) );
  AND2_X1 U11252 ( .A1(n10294), .A2(n10062), .ZN(n8834) );
  NAND2_X1 U11253 ( .A1(n10260), .A2(n8834), .ZN(n10753) );
  INV_X1 U11254 ( .A(n11878), .ZN(n14653) );
  INV_X1 U11255 ( .A(n14650), .ZN(n11938) );
  NAND2_X1 U11256 ( .A1(n11938), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14294) );
  NOR3_X1 U11257 ( .A1(n10753), .A2(n14555), .A3(n14294), .ZN(n8837) );
  OAI21_X1 U11258 ( .B1(n11615), .B2(n14307), .A(P1_B_REG_SCAN_IN), .ZN(n8836)
         );
  OR2_X1 U11259 ( .A1(n8837), .A2(n8836), .ZN(n8838) );
  OAI21_X1 U11260 ( .B1(n8839), .B2(n11615), .A(n8838), .ZN(P1_U3242) );
  INV_X1 U11261 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15031) );
  INV_X1 U11262 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15015) );
  INV_X1 U11263 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14696) );
  NOR2_X1 U11264 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14696), .ZN(n8869) );
  XOR2_X1 U11265 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n8868), .Z(n8923) );
  INV_X1 U11266 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n8866) );
  INV_X1 U11267 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n8864) );
  INV_X1 U11268 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n8862) );
  INV_X1 U11269 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n15155) );
  INV_X1 U11270 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n8888) );
  XNOR2_X1 U11271 ( .A(n8840), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n8883) );
  NOR2_X1 U11272 ( .A1(n8884), .A2(n8883), .ZN(n8842) );
  NOR2_X1 U11273 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n8881), .ZN(n8847) );
  NOR2_X1 U11274 ( .A1(n8845), .A2(n10731), .ZN(n8846) );
  INV_X1 U11275 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n8848) );
  NOR2_X1 U11276 ( .A1(n8849), .A2(n8848), .ZN(n8851) );
  NOR2_X1 U11277 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8897), .ZN(n8850) );
  NOR2_X1 U11278 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n13648), .ZN(n8853) );
  NOR2_X1 U11279 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n8854), .ZN(n8856) );
  XNOR2_X1 U11280 ( .A(n8854), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n8879) );
  NOR2_X1 U11281 ( .A1(n8879), .A2(n8880), .ZN(n8855) );
  XNOR2_X1 U11282 ( .A(n13653), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n8877) );
  NOR2_X1 U11283 ( .A1(n8878), .A2(n8877), .ZN(n8857) );
  XOR2_X1 U11284 ( .A(n13670), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n8909) );
  NAND2_X1 U11285 ( .A1(n8910), .A2(n8909), .ZN(n8858) );
  NAND2_X1 U11286 ( .A1(n8875), .A2(n8874), .ZN(n8860) );
  NOR2_X1 U11287 ( .A1(n8875), .A2(n8874), .ZN(n8859) );
  AOI21_X2 U11288 ( .B1(n15155), .B2(n8860), .A(n8859), .ZN(n8915) );
  XNOR2_X1 U11289 ( .A(n8862), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n8914) );
  NOR2_X1 U11290 ( .A1(n8915), .A2(n8914), .ZN(n8861) );
  XOR2_X1 U11291 ( .A(n8864), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n8916) );
  NAND2_X1 U11292 ( .A1(n8917), .A2(n8916), .ZN(n8863) );
  INV_X1 U11293 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U11294 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n8871), .ZN(n8865) );
  NAND2_X1 U11295 ( .A1(n8923), .A2(n8922), .ZN(n8867) );
  INV_X1 U11296 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14357) );
  OAI22_X1 U11297 ( .A1(n8869), .A2(n8925), .B1(P1_ADDR_REG_15__SCAN_IN), .B2(
        n14357), .ZN(n8928) );
  XNOR2_X1 U11298 ( .A(n14375), .B(P1_ADDR_REG_16__SCAN_IN), .ZN(n8870) );
  XOR2_X1 U11299 ( .A(n8928), .B(n8870), .Z(n14634) );
  INV_X1 U11300 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14991) );
  INV_X1 U11301 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14979) );
  XNOR2_X1 U11302 ( .A(n8871), .B(P1_ADDR_REG_13__SCAN_IN), .ZN(n8872) );
  INV_X1 U11303 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10338) );
  XOR2_X1 U11304 ( .A(n8875), .B(n8874), .Z(n8876) );
  XOR2_X1 U11305 ( .A(n15155), .B(n8876), .Z(n8912) );
  INV_X1 U11306 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14954) );
  XOR2_X1 U11307 ( .A(n8878), .B(n8877), .Z(n8908) );
  XOR2_X1 U11308 ( .A(n8880), .B(n8879), .Z(n15403) );
  INV_X1 U11309 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14927) );
  INV_X1 U11310 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14900) );
  OR2_X1 U11311 ( .A1(n14900), .A2(n8882), .ZN(n8896) );
  INV_X1 U11312 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n13749) );
  XNOR2_X1 U11313 ( .A(n8884), .B(n8883), .ZN(n14315) );
  XNOR2_X1 U11314 ( .A(n8886), .B(n8885), .ZN(n8889) );
  NAND2_X1 U11315 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n8889), .ZN(n8891) );
  AOI21_X1 U11316 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n8888), .A(n8887), .ZN(
        n15401) );
  INV_X1 U11317 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15400) );
  NOR2_X1 U11318 ( .A1(n15401), .A2(n15400), .ZN(n15410) );
  XOR2_X1 U11319 ( .A(n8889), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15409) );
  NAND2_X1 U11320 ( .A1(n15410), .A2(n15409), .ZN(n8890) );
  NAND2_X1 U11321 ( .A1(n8891), .A2(n8890), .ZN(n14316) );
  NAND2_X1 U11322 ( .A1(n14315), .A2(n14316), .ZN(n8892) );
  NOR2_X1 U11323 ( .A1(n14315), .A2(n14316), .ZN(n14314) );
  AOI21_X1 U11324 ( .B1(n13749), .B2(n8892), .A(n14314), .ZN(n15405) );
  INV_X1 U11325 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n13561) );
  XOR2_X1 U11326 ( .A(n13561), .B(n8893), .Z(n15406) );
  NOR2_X1 U11327 ( .A1(n15405), .A2(n15406), .ZN(n8894) );
  INV_X1 U11328 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15407) );
  NAND2_X1 U11329 ( .A1(n15405), .A2(n15406), .ZN(n15404) );
  OAI21_X1 U11330 ( .B1(n8894), .B2(n15407), .A(n15404), .ZN(n15396) );
  NAND2_X1 U11331 ( .A1(n8896), .A2(n8895), .ZN(n8899) );
  XNOR2_X1 U11332 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n8897), .ZN(n8898) );
  NAND2_X1 U11333 ( .A1(n8900), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n8904) );
  INV_X1 U11334 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n14914) );
  XOR2_X1 U11335 ( .A(n13648), .B(P3_ADDR_REG_6__SCAN_IN), .Z(n8902) );
  XOR2_X1 U11336 ( .A(n8902), .B(n8901), .Z(n14322) );
  NAND2_X1 U11337 ( .A1(n14323), .A2(n14322), .ZN(n8903) );
  NAND2_X1 U11338 ( .A1(n8904), .A2(n8903), .ZN(n8905) );
  XNOR2_X1 U11339 ( .A(n14927), .B(n8905), .ZN(n15402) );
  NAND2_X1 U11340 ( .A1(n15403), .A2(n15402), .ZN(n8907) );
  NAND2_X1 U11341 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n8905), .ZN(n8906) );
  XNOR2_X1 U11342 ( .A(n8910), .B(n8909), .ZN(n14331) );
  NAND2_X1 U11343 ( .A1(n14332), .A2(n14331), .ZN(n8911) );
  NOR2_X1 U11344 ( .A1(n14332), .A2(n14331), .ZN(n14330) );
  XOR2_X1 U11345 ( .A(n8915), .B(n8914), .Z(n14618) );
  XNOR2_X1 U11346 ( .A(n8917), .B(n8916), .ZN(n8919) );
  NOR2_X1 U11347 ( .A1(n8918), .A2(n8919), .ZN(n8921) );
  XNOR2_X1 U11348 ( .A(n8919), .B(n8918), .ZN(n14620) );
  XOR2_X1 U11349 ( .A(n8923), .B(n8922), .Z(n14626) );
  NAND2_X1 U11350 ( .A1(n14625), .A2(n14626), .ZN(n8924) );
  AOI21_X2 U11351 ( .B1(n14991), .B2(n8924), .A(n14624), .ZN(n14629) );
  XOR2_X1 U11352 ( .A(n14696), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n8926) );
  XOR2_X1 U11353 ( .A(n8926), .B(n8925), .Z(n14630) );
  INV_X1 U11354 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15002) );
  INV_X1 U11355 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14396) );
  NOR2_X1 U11356 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14375), .ZN(n8929) );
  INV_X1 U11357 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n8927) );
  OAI22_X1 U11358 ( .A1(n8929), .A2(n8928), .B1(P3_ADDR_REG_16__SCAN_IN), .B2(
        n8927), .ZN(n8931) );
  XOR2_X1 U11359 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n8931), .Z(n8932) );
  XOR2_X1 U11360 ( .A(n14396), .B(n8932), .Z(n14347) );
  NAND2_X1 U11361 ( .A1(n14348), .A2(n14347), .ZN(n8930) );
  NOR2_X1 U11362 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n8931), .ZN(n8934) );
  AND2_X1 U11363 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n8932), .ZN(n8933) );
  NOR2_X1 U11364 ( .A1(n8934), .A2(n8933), .ZN(n8938) );
  INV_X1 U11365 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n13691) );
  XNOR2_X1 U11366 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(n13691), .ZN(n8937) );
  XNOR2_X1 U11367 ( .A(n8938), .B(n8937), .ZN(n8936) );
  XNOR2_X1 U11368 ( .A(n8936), .B(n8935), .ZN(n14311) );
  NOR2_X1 U11369 ( .A1(n8938), .A2(n8937), .ZN(n8939) );
  AOI21_X1 U11370 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n13691), .A(n8939), .ZN(
        n8940) );
  INV_X1 U11371 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n12606) );
  INV_X1 U11372 ( .A(n8155), .ZN(n13088) );
  NAND3_X1 U11373 ( .A1(n10408), .A2(n9856), .A3(n10308), .ZN(n8942) );
  NAND2_X1 U11374 ( .A1(n8943), .A2(n8942), .ZN(n8946) );
  MUX2_X1 U11375 ( .A(n6745), .B(n10595), .S(n6589), .Z(n8945) );
  INV_X1 U11376 ( .A(n8156), .ZN(n13086) );
  MUX2_X1 U11377 ( .A(n13086), .B(n7573), .S(n9122), .Z(n8944) );
  OAI21_X1 U11378 ( .B1(n8946), .B2(n8945), .A(n8944), .ZN(n8948) );
  NAND2_X1 U11379 ( .A1(n8946), .A2(n8945), .ZN(n8947) );
  NAND2_X1 U11380 ( .A1(n8948), .A2(n8947), .ZN(n8951) );
  NAND2_X1 U11381 ( .A1(n8951), .A2(n8952), .ZN(n8950) );
  NAND2_X1 U11382 ( .A1(n8950), .A2(n8949), .ZN(n8956) );
  INV_X1 U11383 ( .A(n8951), .ZN(n8954) );
  INV_X1 U11384 ( .A(n8952), .ZN(n8953) );
  MUX2_X1 U11385 ( .A(n13084), .B(n9871), .S(n6589), .Z(n8958) );
  MUX2_X1 U11386 ( .A(n13084), .B(n9871), .S(n9122), .Z(n8957) );
  INV_X1 U11387 ( .A(n8958), .ZN(n8959) );
  MUX2_X1 U11388 ( .A(n13083), .B(n13022), .S(n9122), .Z(n8963) );
  NAND2_X1 U11389 ( .A1(n8962), .A2(n8963), .ZN(n8961) );
  MUX2_X1 U11390 ( .A(n13022), .B(n13083), .S(n9122), .Z(n8960) );
  NAND2_X1 U11391 ( .A1(n8961), .A2(n8960), .ZN(n8967) );
  INV_X1 U11392 ( .A(n8962), .ZN(n8965) );
  INV_X1 U11393 ( .A(n8963), .ZN(n8964) );
  NAND2_X1 U11394 ( .A1(n8965), .A2(n8964), .ZN(n8966) );
  NAND2_X1 U11395 ( .A1(n8967), .A2(n8966), .ZN(n8970) );
  MUX2_X1 U11396 ( .A(n13082), .B(n11242), .S(n6589), .Z(n8971) );
  NAND2_X1 U11397 ( .A1(n8970), .A2(n8971), .ZN(n8969) );
  MUX2_X1 U11398 ( .A(n13082), .B(n11242), .S(n9122), .Z(n8968) );
  NAND2_X1 U11399 ( .A1(n8969), .A2(n8968), .ZN(n8978) );
  MUX2_X1 U11400 ( .A(n13081), .B(n10869), .S(n9122), .Z(n8979) );
  NAND2_X1 U11401 ( .A1(n8974), .A2(n8979), .ZN(n8976) );
  MUX2_X1 U11402 ( .A(n13081), .B(n10869), .S(n6589), .Z(n8975) );
  NAND2_X1 U11403 ( .A1(n8976), .A2(n8975), .ZN(n8983) );
  AND2_X1 U11404 ( .A1(n8978), .A2(n8977), .ZN(n8981) );
  INV_X1 U11405 ( .A(n8979), .ZN(n8980) );
  NAND2_X1 U11406 ( .A1(n8981), .A2(n8980), .ZN(n8982) );
  MUX2_X1 U11407 ( .A(n13080), .B(n15057), .S(n6589), .Z(n8985) );
  MUX2_X1 U11408 ( .A(n13080), .B(n15057), .S(n9122), .Z(n8984) );
  MUX2_X1 U11409 ( .A(n13079), .B(n11052), .S(n9122), .Z(n8989) );
  NAND2_X1 U11410 ( .A1(n8988), .A2(n8989), .ZN(n8987) );
  MUX2_X1 U11411 ( .A(n13079), .B(n11052), .S(n6589), .Z(n8986) );
  NAND2_X1 U11412 ( .A1(n8987), .A2(n8986), .ZN(n8993) );
  INV_X1 U11413 ( .A(n8988), .ZN(n8991) );
  INV_X1 U11414 ( .A(n8989), .ZN(n8990) );
  NAND2_X1 U11415 ( .A1(n8991), .A2(n8990), .ZN(n8992) );
  MUX2_X1 U11416 ( .A(n13078), .B(n11339), .S(n6589), .Z(n8995) );
  MUX2_X1 U11417 ( .A(n13078), .B(n11339), .S(n9122), .Z(n8994) );
  INV_X1 U11418 ( .A(n8995), .ZN(n8996) );
  MUX2_X1 U11419 ( .A(n13077), .B(n11356), .S(n9122), .Z(n9000) );
  NAND2_X1 U11420 ( .A1(n8999), .A2(n9000), .ZN(n8998) );
  MUX2_X1 U11421 ( .A(n13077), .B(n11356), .S(n6589), .Z(n8997) );
  NAND2_X1 U11422 ( .A1(n8998), .A2(n8997), .ZN(n9004) );
  INV_X1 U11423 ( .A(n8999), .ZN(n9002) );
  INV_X1 U11424 ( .A(n9000), .ZN(n9001) );
  NAND2_X1 U11425 ( .A1(n9002), .A2(n9001), .ZN(n9003) );
  MUX2_X1 U11426 ( .A(n13076), .B(n11551), .S(n6589), .Z(n9006) );
  MUX2_X1 U11427 ( .A(n13076), .B(n11551), .S(n9122), .Z(n9005) );
  MUX2_X1 U11428 ( .A(n13075), .B(n14482), .S(n9122), .Z(n9010) );
  NAND2_X1 U11429 ( .A1(n9009), .A2(n9010), .ZN(n9008) );
  MUX2_X1 U11430 ( .A(n13075), .B(n14482), .S(n6589), .Z(n9007) );
  NAND2_X1 U11431 ( .A1(n9008), .A2(n9007), .ZN(n9014) );
  INV_X1 U11432 ( .A(n9009), .ZN(n9012) );
  INV_X1 U11433 ( .A(n9010), .ZN(n9011) );
  NAND2_X1 U11434 ( .A1(n9012), .A2(n9011), .ZN(n9013) );
  MUX2_X1 U11435 ( .A(n13074), .B(n11563), .S(n6589), .Z(n9016) );
  MUX2_X1 U11436 ( .A(n13074), .B(n11563), .S(n9122), .Z(n9015) );
  INV_X1 U11437 ( .A(n9016), .ZN(n9017) );
  MUX2_X1 U11438 ( .A(n13073), .B(n14461), .S(n9122), .Z(n9021) );
  NAND2_X1 U11439 ( .A1(n9020), .A2(n9021), .ZN(n9019) );
  MUX2_X1 U11440 ( .A(n13073), .B(n14461), .S(n6589), .Z(n9018) );
  NAND2_X1 U11441 ( .A1(n9019), .A2(n9018), .ZN(n9025) );
  INV_X1 U11442 ( .A(n9020), .ZN(n9023) );
  INV_X1 U11443 ( .A(n9021), .ZN(n9022) );
  NAND2_X1 U11444 ( .A1(n9023), .A2(n9022), .ZN(n9024) );
  MUX2_X1 U11445 ( .A(n13072), .B(n11841), .S(n6589), .Z(n9027) );
  MUX2_X1 U11446 ( .A(n13072), .B(n11841), .S(n9122), .Z(n9026) );
  MUX2_X1 U11447 ( .A(n13334), .B(n13437), .S(n6589), .Z(n9036) );
  MUX2_X1 U11448 ( .A(n11847), .B(n13445), .S(n9122), .Z(n9032) );
  MUX2_X1 U11449 ( .A(n13071), .B(n11829), .S(n6589), .Z(n9031) );
  AOI22_X1 U11450 ( .A1(n9036), .A2(n9154), .B1(n9032), .B2(n9031), .ZN(n9029)
         );
  NAND2_X1 U11451 ( .A1(n9030), .A2(n9029), .ZN(n9049) );
  INV_X1 U11452 ( .A(n9031), .ZN(n9034) );
  INV_X1 U11453 ( .A(n9032), .ZN(n9033) );
  NAND2_X1 U11454 ( .A1(n9034), .A2(n9033), .ZN(n9037) );
  NAND2_X1 U11455 ( .A1(n9035), .A2(n9037), .ZN(n9041) );
  INV_X1 U11456 ( .A(n9036), .ZN(n9040) );
  INV_X1 U11457 ( .A(n9037), .ZN(n9039) );
  AOI22_X1 U11458 ( .A1(n9041), .A2(n9040), .B1(n9039), .B2(n9038), .ZN(n9047)
         );
  MUX2_X1 U11459 ( .A(n13070), .B(n13429), .S(n6589), .Z(n9042) );
  AND2_X1 U11460 ( .A1(n9047), .A2(n9042), .ZN(n9044) );
  INV_X1 U11461 ( .A(n9042), .ZN(n9043) );
  MUX2_X1 U11462 ( .A(n13070), .B(n13429), .S(n9122), .Z(n9045) );
  INV_X1 U11463 ( .A(n9045), .ZN(n9046) );
  AND2_X1 U11464 ( .A1(n9047), .A2(n9046), .ZN(n9048) );
  NAND2_X1 U11465 ( .A1(n9049), .A2(n9048), .ZN(n9050) );
  MUX2_X1 U11466 ( .A(n13337), .B(n13426), .S(n6589), .Z(n9053) );
  MUX2_X1 U11467 ( .A(n13337), .B(n13426), .S(n9122), .Z(n9052) );
  INV_X1 U11468 ( .A(n9053), .ZN(n9054) );
  MUX2_X1 U11469 ( .A(n13069), .B(n13420), .S(n9122), .Z(n9058) );
  NAND2_X1 U11470 ( .A1(n9057), .A2(n9058), .ZN(n9056) );
  MUX2_X1 U11471 ( .A(n13069), .B(n13420), .S(n6589), .Z(n9055) );
  NAND2_X1 U11472 ( .A1(n9056), .A2(n9055), .ZN(n9062) );
  INV_X1 U11473 ( .A(n9057), .ZN(n9060) );
  INV_X1 U11474 ( .A(n9058), .ZN(n9059) );
  NAND2_X1 U11475 ( .A1(n9060), .A2(n9059), .ZN(n9061) );
  NAND2_X1 U11476 ( .A1(n9062), .A2(n9061), .ZN(n9065) );
  MUX2_X1 U11477 ( .A(n13272), .B(n13295), .S(n6589), .Z(n9066) );
  NAND2_X1 U11478 ( .A1(n9065), .A2(n9066), .ZN(n9064) );
  MUX2_X1 U11479 ( .A(n13272), .B(n13295), .S(n9122), .Z(n9063) );
  NAND2_X1 U11480 ( .A1(n9064), .A2(n9063), .ZN(n9070) );
  INV_X1 U11481 ( .A(n9065), .ZN(n9068) );
  INV_X1 U11482 ( .A(n9066), .ZN(n9067) );
  NAND2_X1 U11483 ( .A1(n9068), .A2(n9067), .ZN(n9069) );
  MUX2_X1 U11484 ( .A(n13068), .B(n13409), .S(n9122), .Z(n9072) );
  MUX2_X1 U11485 ( .A(n13068), .B(n13409), .S(n6589), .Z(n9071) );
  MUX2_X1 U11486 ( .A(n13271), .B(n13404), .S(n6589), .Z(n9076) );
  NAND2_X1 U11487 ( .A1(n9075), .A2(n9076), .ZN(n9074) );
  MUX2_X1 U11488 ( .A(n13271), .B(n13404), .S(n9122), .Z(n9073) );
  NAND2_X1 U11489 ( .A1(n9074), .A2(n9073), .ZN(n9080) );
  INV_X1 U11490 ( .A(n9075), .ZN(n9078) );
  INV_X1 U11491 ( .A(n9076), .ZN(n9077) );
  NAND2_X1 U11492 ( .A1(n9078), .A2(n9077), .ZN(n9079) );
  NAND2_X1 U11493 ( .A1(n9080), .A2(n9079), .ZN(n9083) );
  MUX2_X1 U11494 ( .A(n13067), .B(n13249), .S(n9122), .Z(n9084) );
  NAND2_X1 U11495 ( .A1(n9083), .A2(n9084), .ZN(n9082) );
  MUX2_X1 U11496 ( .A(n13249), .B(n13067), .S(n9122), .Z(n9081) );
  NAND2_X1 U11497 ( .A1(n9082), .A2(n9081), .ZN(n9088) );
  INV_X1 U11498 ( .A(n9083), .ZN(n9086) );
  INV_X1 U11499 ( .A(n9084), .ZN(n9085) );
  NAND2_X1 U11500 ( .A1(n9086), .A2(n9085), .ZN(n9087) );
  MUX2_X1 U11501 ( .A(n13066), .B(n13392), .S(n6589), .Z(n9090) );
  MUX2_X1 U11502 ( .A(n13066), .B(n13392), .S(n9122), .Z(n9089) );
  INV_X1 U11503 ( .A(n9090), .ZN(n9091) );
  MUX2_X1 U11504 ( .A(n13065), .B(n13387), .S(n9122), .Z(n9095) );
  NAND2_X1 U11505 ( .A1(n9094), .A2(n9095), .ZN(n9093) );
  MUX2_X1 U11506 ( .A(n13387), .B(n13065), .S(n9122), .Z(n9092) );
  NAND2_X1 U11507 ( .A1(n9093), .A2(n9092), .ZN(n9113) );
  INV_X1 U11508 ( .A(n9094), .ZN(n9097) );
  INV_X1 U11509 ( .A(n9095), .ZN(n9096) );
  NAND2_X1 U11510 ( .A1(n9097), .A2(n9096), .ZN(n9112) );
  NAND2_X1 U11511 ( .A1(n14285), .A2(n9118), .ZN(n9099) );
  INV_X1 U11512 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13477) );
  OR2_X1 U11513 ( .A1(n9119), .A2(n13477), .ZN(n9098) );
  INV_X1 U11514 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9104) );
  NAND2_X1 U11515 ( .A1(n9100), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9103) );
  NAND2_X1 U11516 ( .A1(n9101), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9102) );
  OAI211_X1 U11517 ( .C1(n9105), .C2(n9104), .A(n9103), .B(n9102), .ZN(n13168)
         );
  NAND2_X1 U11518 ( .A1(n13451), .A2(n13168), .ZN(n9106) );
  NAND2_X1 U11519 ( .A1(n9148), .A2(n9106), .ZN(n9178) );
  MUX2_X1 U11520 ( .A(n12120), .B(n11882), .S(n6589), .Z(n9130) );
  MUX2_X1 U11521 ( .A(n13062), .B(n7099), .S(n9122), .Z(n9129) );
  NAND2_X1 U11522 ( .A1(n9130), .A2(n9129), .ZN(n9135) );
  MUX2_X1 U11523 ( .A(n12969), .B(n13459), .S(n6589), .Z(n9132) );
  MUX2_X1 U11524 ( .A(n13063), .B(n7104), .S(n9122), .Z(n9131) );
  NAND2_X1 U11525 ( .A1(n9132), .A2(n9131), .ZN(n9107) );
  AND2_X1 U11526 ( .A1(n9135), .A2(n9107), .ZN(n9108) );
  NAND2_X1 U11527 ( .A1(n9178), .A2(n9108), .ZN(n9140) );
  MUX2_X1 U11528 ( .A(n13064), .B(n7105), .S(n9122), .Z(n9114) );
  MUX2_X1 U11529 ( .A(n13053), .B(n13202), .S(n6589), .Z(n9115) );
  NAND2_X1 U11530 ( .A1(n9110), .A2(n9109), .ZN(n9111) );
  AOI21_X1 U11531 ( .B1(n9113), .B2(n9112), .A(n9111), .ZN(n9145) );
  INV_X1 U11532 ( .A(n9114), .ZN(n9117) );
  INV_X1 U11533 ( .A(n9115), .ZN(n9116) );
  NAND2_X1 U11534 ( .A1(n9117), .A2(n9116), .ZN(n9139) );
  NAND2_X1 U11535 ( .A1(n11874), .A2(n9118), .ZN(n9121) );
  INV_X1 U11536 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12312) );
  OR2_X1 U11537 ( .A1(n9119), .A2(n12312), .ZN(n9120) );
  MUX2_X1 U11538 ( .A(n13061), .B(n13165), .S(n9122), .Z(n9142) );
  NAND2_X1 U11539 ( .A1(n13168), .A2(n9122), .ZN(n9146) );
  OAI211_X1 U11540 ( .C1(n9124), .C2(n9123), .A(n9179), .B(n9193), .ZN(n9125)
         );
  INV_X1 U11541 ( .A(n9125), .ZN(n9127) );
  INV_X1 U11542 ( .A(n13061), .ZN(n9126) );
  AOI21_X1 U11543 ( .B1(n9146), .B2(n9127), .A(n9126), .ZN(n9128) );
  AOI21_X1 U11544 ( .B1(n13165), .B2(n6589), .A(n9128), .ZN(n9141) );
  OAI22_X1 U11545 ( .A1(n9142), .A2(n9141), .B1(n9130), .B2(n9129), .ZN(n9137)
         );
  INV_X1 U11546 ( .A(n9131), .ZN(n9134) );
  INV_X1 U11547 ( .A(n9132), .ZN(n9133) );
  AND3_X1 U11548 ( .A1(n9135), .A2(n9134), .A3(n9133), .ZN(n9136) );
  OAI21_X1 U11549 ( .B1(n9137), .B2(n9136), .A(n9178), .ZN(n9138) );
  OAI21_X1 U11550 ( .B1(n9140), .B2(n9139), .A(n9138), .ZN(n9144) );
  NAND2_X1 U11551 ( .A1(n9142), .A2(n9141), .ZN(n9143) );
  OAI21_X1 U11552 ( .B1(n9145), .B2(n9144), .A(n9143), .ZN(n9185) );
  INV_X1 U11553 ( .A(n9146), .ZN(n9147) );
  AOI21_X1 U11554 ( .B1(n13451), .B2(n6589), .A(n9147), .ZN(n9149) );
  INV_X1 U11555 ( .A(n9191), .ZN(n9153) );
  OAI21_X1 U11556 ( .B1(n13161), .B2(n11373), .A(n9193), .ZN(n9150) );
  AOI21_X1 U11557 ( .B1(n9856), .B2(n11590), .A(n9150), .ZN(n9151) );
  INV_X1 U11558 ( .A(n9151), .ZN(n9152) );
  INV_X1 U11559 ( .A(n10165), .ZN(n9852) );
  AND2_X1 U11560 ( .A1(n9852), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9192) );
  NAND4_X1 U11561 ( .A1(n9185), .A2(n9153), .A3(n9152), .A4(n9192), .ZN(n9203)
         );
  XNOR2_X1 U11562 ( .A(n13165), .B(n13061), .ZN(n9176) );
  NAND2_X1 U11563 ( .A1(n9155), .A2(n9154), .ZN(n13363) );
  XNOR2_X1 U11564 ( .A(n11563), .B(n14442), .ZN(n11557) );
  NAND2_X1 U11565 ( .A1(n9156), .A2(n10408), .ZN(n11009) );
  NOR2_X1 U11566 ( .A1(n11009), .A2(n11262), .ZN(n9158) );
  NAND4_X1 U11567 ( .A1(n9158), .A2(n11076), .A3(n9994), .A4(n10583), .ZN(
        n9159) );
  NOR2_X1 U11568 ( .A1(n9159), .A2(n11026), .ZN(n9162) );
  NAND4_X1 U11569 ( .A1(n10982), .A2(n9162), .A3(n9161), .A4(n9160), .ZN(n9163) );
  OR4_X1 U11570 ( .A1(n11345), .A2(n11213), .A3(n11045), .A4(n9163), .ZN(n9164) );
  OR4_X1 U11571 ( .A1(n11557), .A2(n9164), .A3(n11459), .A4(n11487), .ZN(n9165) );
  NOR2_X1 U11572 ( .A1(n9166), .A2(n9165), .ZN(n9167) );
  NAND4_X1 U11573 ( .A1(n13363), .A2(n9167), .A3(n11764), .A4(n11758), .ZN(
        n9168) );
  NOR2_X1 U11574 ( .A1(n13332), .A2(n9168), .ZN(n9169) );
  XNOR2_X1 U11575 ( .A(n13426), .B(n13337), .ZN(n13317) );
  NAND4_X1 U11576 ( .A1(n13290), .A2(n9169), .A3(n13310), .A4(n13317), .ZN(
        n9170) );
  NOR2_X1 U11577 ( .A1(n13269), .A2(n9170), .ZN(n9171) );
  XNOR2_X1 U11578 ( .A(n13404), .B(n13271), .ZN(n13259) );
  NAND4_X1 U11579 ( .A1(n13230), .A2(n9171), .A3(n13259), .A4(n13246), .ZN(
        n9172) );
  NOR2_X1 U11580 ( .A1(n13215), .A2(n9172), .ZN(n9173) );
  AND2_X1 U11581 ( .A1(n13180), .A2(n9173), .ZN(n9175) );
  AND4_X1 U11582 ( .A1(n9176), .A2(n9175), .A3(n9174), .A4(n13206), .ZN(n9177)
         );
  AND2_X1 U11583 ( .A1(n9178), .A2(n9177), .ZN(n9186) );
  MUX2_X1 U11584 ( .A(n9179), .B(n9195), .S(n11262), .Z(n9190) );
  INV_X1 U11585 ( .A(n9190), .ZN(n9180) );
  AND2_X1 U11586 ( .A1(n9192), .A2(n13161), .ZN(n9189) );
  OAI21_X1 U11587 ( .B1(n9190), .B2(n11373), .A(n9189), .ZN(n9181) );
  INV_X1 U11588 ( .A(n9181), .ZN(n9182) );
  INV_X1 U11589 ( .A(n9186), .ZN(n9199) );
  NAND4_X1 U11590 ( .A1(n9199), .A2(n13161), .A3(n9192), .A4(n11373), .ZN(
        n9187) );
  AOI21_X1 U11591 ( .B1(n11262), .B2(n9153), .A(n9187), .ZN(n9188) );
  INV_X1 U11592 ( .A(n9188), .ZN(n9202) );
  NAND3_X1 U11593 ( .A1(n9192), .A2(n11373), .A3(n11192), .ZN(n9198) );
  NAND3_X1 U11594 ( .A1(n9191), .A2(n9190), .A3(n9189), .ZN(n9197) );
  INV_X1 U11595 ( .A(n9192), .ZN(n11611) );
  INV_X1 U11596 ( .A(n6740), .ZN(n10171) );
  INV_X1 U11597 ( .A(n9193), .ZN(n9979) );
  NAND4_X1 U11598 ( .A1(n15078), .A2(n10171), .A3(n9979), .A4(n13335), .ZN(
        n9194) );
  OAI211_X1 U11599 ( .C1(n9195), .C2(n11611), .A(n9194), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9196) );
  OAI211_X1 U11600 ( .C1(n9199), .C2(n9198), .A(n9197), .B(n9196), .ZN(n9200)
         );
  INV_X1 U11601 ( .A(n9200), .ZN(n9201) );
  NAND4_X1 U11602 ( .A1(n9203), .A2(n6657), .A3(n9202), .A4(n9201), .ZN(
        P2_U3328) );
  INV_X1 U11603 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9816) );
  NOR2_X1 U11604 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n9207) );
  NOR2_X1 U11605 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n9211) );
  NOR2_X1 U11606 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n9210) );
  NAND4_X1 U11607 ( .A1(n9211), .A2(n9210), .A3(n6874), .A4(n6875), .ZN(n9213)
         );
  NAND4_X1 U11608 ( .A1(n9571), .A2(n9539), .A3(n9496), .A4(n9535), .ZN(n9212)
         );
  NOR2_X1 U11609 ( .A1(n9213), .A2(n9212), .ZN(n9214) );
  NAND2_X1 U11610 ( .A1(n9219), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9220) );
  INV_X1 U11611 ( .A(SI_1_), .ZN(n10032) );
  OAI21_X1 U11612 ( .B1(n9225), .B2(n9224), .A(n9253), .ZN(n10031) );
  INV_X1 U11613 ( .A(n9738), .ZN(n9228) );
  NAND2_X1 U11614 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n9227) );
  NAND2_X1 U11615 ( .A1(n9228), .A2(n10435), .ZN(n9229) );
  NAND2_X1 U11616 ( .A1(n9230), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9233) );
  MUX2_X1 U11617 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9233), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n9234) );
  AND2_X2 U11618 ( .A1(n9234), .A2(n7205), .ZN(n9235) );
  INV_X2 U11619 ( .A(n9235), .ZN(n12959) );
  INV_X1 U11620 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10635) );
  AND2_X4 U11621 ( .A1(n11871), .A2(n9235), .ZN(n12302) );
  NAND2_X1 U11622 ( .A1(n12302), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9239) );
  INV_X1 U11623 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n12828) );
  OR2_X1 U11624 ( .A1(n9262), .A2(n12828), .ZN(n9238) );
  INV_X1 U11625 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n9236) );
  NAND2_X1 U11626 ( .A1(n12302), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9246) );
  INV_X1 U11627 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n9241) );
  INV_X1 U11628 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10656) );
  INV_X1 U11629 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n9242) );
  OR2_X1 U11630 ( .A1(n12304), .A2(n9242), .ZN(n9243) );
  XNOR2_X1 U11631 ( .A(n7005), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9247) );
  MUX2_X1 U11632 ( .A(n9247), .B(SI_0_), .S(n8655), .Z(n12963) );
  MUX2_X1 U11633 ( .A(P3_IR_REG_0__SCAN_IN), .B(n12963), .S(n9738), .Z(n10658)
         );
  NAND2_X1 U11634 ( .A1(n12817), .A2(n10658), .ZN(n12816) );
  NAND2_X1 U11635 ( .A1(n10827), .A2(n10876), .ZN(n15316) );
  NAND2_X1 U11636 ( .A1(n15318), .A2(n15316), .ZN(n9259) );
  NAND2_X1 U11637 ( .A1(n9279), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9252) );
  INV_X1 U11638 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10437) );
  INV_X1 U11639 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15311) );
  OR2_X1 U11640 ( .A1(n9262), .A2(n15311), .ZN(n9250) );
  INV_X1 U11641 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15332) );
  OR2_X1 U11642 ( .A1(n9304), .A2(n15332), .ZN(n9249) );
  NAND2_X1 U11643 ( .A1(n12319), .A2(n10027), .ZN(n9258) );
  XNOR2_X1 U11644 ( .A(n9269), .B(n9267), .ZN(n10028) );
  NAND2_X1 U11645 ( .A1(n12318), .A2(n10028), .ZN(n9257) );
  INV_X4 U11646 ( .A(n9738), .ZN(n10421) );
  INV_X1 U11647 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n13716) );
  XNOR2_X2 U11648 ( .A(n9255), .B(n13716), .ZN(n10631) );
  NAND2_X1 U11649 ( .A1(n10421), .A2(n10631), .ZN(n9256) );
  NAND2_X1 U11650 ( .A1(n12819), .A2(n15310), .ZN(n9260) );
  NAND2_X1 U11651 ( .A1(n9279), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9266) );
  INV_X1 U11652 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n9261) );
  OR2_X1 U11653 ( .A1(n9281), .A2(n9261), .ZN(n9265) );
  OR2_X1 U11654 ( .A1(n9262), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n9264) );
  INV_X1 U11655 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10927) );
  OR2_X1 U11656 ( .A1(n9304), .A2(n10927), .ZN(n9263) );
  INV_X1 U11657 ( .A(SI_3_), .ZN(n10029) );
  NAND2_X1 U11658 ( .A1(n12319), .A2(n10029), .ZN(n9276) );
  INV_X1 U11659 ( .A(n9267), .ZN(n9268) );
  NAND2_X1 U11660 ( .A1(n10003), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9270) );
  XNOR2_X1 U11661 ( .A(n7621), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n9288) );
  XNOR2_X1 U11662 ( .A(n9290), .B(n9288), .ZN(n10030) );
  NAND2_X1 U11663 ( .A1(n12318), .A2(n10030), .ZN(n9275) );
  INV_X1 U11664 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n9273) );
  NAND2_X1 U11665 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n9271), .ZN(n9272) );
  XNOR2_X1 U11666 ( .A(n9273), .B(n9272), .ZN(n10546) );
  NAND2_X1 U11667 ( .A1(n10421), .A2(n10546), .ZN(n9274) );
  INV_X1 U11668 ( .A(n10843), .ZN(n10928) );
  NAND2_X1 U11669 ( .A1(n15293), .A2(n10843), .ZN(n15286) );
  NAND2_X1 U11670 ( .A1(n9277), .A2(n10843), .ZN(n9278) );
  NAND2_X1 U11671 ( .A1(n10923), .A2(n9278), .ZN(n15291) );
  NAND2_X1 U11672 ( .A1(n9279), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9287) );
  INV_X1 U11673 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n9280) );
  OR2_X1 U11674 ( .A1(n9281), .A2(n9280), .ZN(n9286) );
  NOR2_X1 U11675 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9301) );
  AND2_X1 U11676 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9282) );
  NOR2_X1 U11677 ( .A1(n9301), .A2(n9282), .ZN(n15303) );
  OR2_X1 U11678 ( .A1(n9262), .A2(n15303), .ZN(n9285) );
  INV_X1 U11679 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n9283) );
  OR2_X1 U11680 ( .A1(n9304), .A2(n9283), .ZN(n9284) );
  INV_X1 U11681 ( .A(n9288), .ZN(n9289) );
  NAND2_X1 U11682 ( .A1(n9290), .A2(n9289), .ZN(n9292) );
  NAND2_X1 U11683 ( .A1(n7621), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9291) );
  XNOR2_X1 U11684 ( .A(n10014), .B(P2_DATAO_REG_4__SCAN_IN), .ZN(n9310) );
  XNOR2_X1 U11685 ( .A(n9312), .B(n9310), .ZN(n14318) );
  NAND2_X1 U11686 ( .A1(n12318), .A2(n14318), .ZN(n9298) );
  INV_X1 U11687 ( .A(SI_4_), .ZN(n9293) );
  NAND2_X1 U11688 ( .A1(n12319), .A2(n9293), .ZN(n9297) );
  NAND2_X1 U11689 ( .A1(n9315), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9295) );
  INV_X1 U11690 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n9294) );
  XNOR2_X1 U11691 ( .A(n9295), .B(n9294), .ZN(n14321) );
  NAND2_X1 U11692 ( .A1(n10421), .A2(n14321), .ZN(n9296) );
  NAND2_X1 U11693 ( .A1(n10841), .A2(n15302), .ZN(n12356) );
  INV_X1 U11694 ( .A(n15302), .ZN(n9299) );
  NAND2_X1 U11695 ( .A1(n12524), .A2(n9299), .ZN(n12355) );
  NAND2_X1 U11696 ( .A1(n12356), .A2(n12355), .ZN(n15290) );
  INV_X1 U11697 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9300) );
  NAND2_X1 U11698 ( .A1(n9301), .A2(n9300), .ZN(n9325) );
  OR2_X1 U11699 ( .A1(n9301), .A2(n9300), .ZN(n9302) );
  AND2_X1 U11700 ( .A1(n9325), .A2(n9302), .ZN(n11234) );
  OR2_X1 U11701 ( .A1(n9262), .A2(n11234), .ZN(n9309) );
  NAND2_X1 U11702 ( .A1(n12302), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n9308) );
  INV_X1 U11703 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n9303) );
  OR2_X1 U11704 ( .A1(n12304), .A2(n9303), .ZN(n9307) );
  INV_X1 U11705 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n9305) );
  OR2_X1 U11706 ( .A1(n9304), .A2(n9305), .ZN(n9306) );
  NAND4_X1 U11707 ( .A1(n9309), .A2(n9308), .A3(n9307), .A4(n9306), .ZN(n15276) );
  INV_X1 U11708 ( .A(SI_5_), .ZN(n10022) );
  NAND2_X1 U11709 ( .A1(n12319), .A2(n10022), .ZN(n9322) );
  INV_X1 U11710 ( .A(n9310), .ZN(n9311) );
  NAND2_X1 U11711 ( .A1(n10014), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9313) );
  XNOR2_X1 U11712 ( .A(n10041), .B(P1_DATAO_REG_5__SCAN_IN), .ZN(n9314) );
  XNOR2_X1 U11713 ( .A(n9334), .B(n9314), .ZN(n10023) );
  NAND2_X1 U11714 ( .A1(n12318), .A2(n10023), .ZN(n9321) );
  NOR2_X1 U11715 ( .A1(n9315), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n9318) );
  OR2_X1 U11716 ( .A1(n9318), .A2(n9231), .ZN(n9316) );
  MUX2_X1 U11717 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9316), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n9319) );
  NAND2_X1 U11718 ( .A1(n9318), .A2(n9317), .ZN(n9351) );
  NAND2_X1 U11719 ( .A1(n9319), .A2(n9351), .ZN(n10745) );
  NAND2_X1 U11720 ( .A1(n10421), .A2(n10745), .ZN(n9320) );
  XNOR2_X1 U11721 ( .A(n15276), .B(n11000), .ZN(n12358) );
  INV_X1 U11722 ( .A(n15276), .ZN(n15295) );
  INV_X1 U11723 ( .A(n11000), .ZN(n12360) );
  NAND2_X1 U11724 ( .A1(n15295), .A2(n12360), .ZN(n9324) );
  NAND2_X1 U11725 ( .A1(n9741), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9331) );
  INV_X1 U11726 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10554) );
  OR2_X1 U11727 ( .A1(n9281), .A2(n10554), .ZN(n9330) );
  NAND2_X1 U11728 ( .A1(n9325), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9326) );
  AND2_X1 U11729 ( .A1(n9341), .A2(n9326), .ZN(n15282) );
  OR2_X1 U11730 ( .A1(n9262), .A2(n15282), .ZN(n9329) );
  INV_X1 U11731 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n9327) );
  OR2_X1 U11732 ( .A1(n12304), .A2(n9327), .ZN(n9328) );
  INV_X1 U11733 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10040) );
  AND2_X1 U11734 ( .A1(n10040), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9333) );
  NAND2_X1 U11735 ( .A1(n10041), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n9332) );
  XNOR2_X1 U11736 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n9335) );
  XNOR2_X1 U11737 ( .A(n9349), .B(n9335), .ZN(n10019) );
  NAND2_X1 U11738 ( .A1(n12319), .A2(SI_6_), .ZN(n9338) );
  NAND2_X1 U11739 ( .A1(n9351), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9336) );
  NAND2_X1 U11740 ( .A1(n10421), .A2(n10674), .ZN(n9337) );
  OAI211_X1 U11741 ( .C1(n9603), .C2(n10019), .A(n9338), .B(n9337), .ZN(n15281) );
  NAND2_X1 U11742 ( .A1(n15260), .A2(n15281), .ZN(n12366) );
  INV_X1 U11743 ( .A(n15281), .ZN(n9339) );
  NAND2_X1 U11744 ( .A1(n12523), .A2(n9339), .ZN(n12367) );
  NAND2_X1 U11745 ( .A1(n9279), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9347) );
  INV_X1 U11746 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n9340) );
  OR2_X1 U11747 ( .A1(n9281), .A2(n9340), .ZN(n9346) );
  AND2_X1 U11748 ( .A1(n9341), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9342) );
  NOR2_X1 U11749 ( .A1(n9358), .A2(n9342), .ZN(n15261) );
  OR2_X1 U11750 ( .A1(n9262), .A2(n15261), .ZN(n9345) );
  INV_X1 U11751 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n9343) );
  OR2_X1 U11752 ( .A1(n9304), .A2(n9343), .ZN(n9344) );
  AND2_X1 U11753 ( .A1(n10048), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9348) );
  NAND2_X1 U11754 ( .A1(n10059), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9366) );
  INV_X1 U11755 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10061) );
  NAND2_X1 U11756 ( .A1(n10061), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n9350) );
  NAND2_X1 U11757 ( .A1(n9366), .A2(n9350), .ZN(n9367) );
  XNOR2_X1 U11758 ( .A(n9368), .B(n9367), .ZN(n10034) );
  NAND2_X1 U11759 ( .A1(n12318), .A2(n10034), .ZN(n9356) );
  INV_X1 U11760 ( .A(SI_7_), .ZN(n10035) );
  NAND2_X1 U11761 ( .A1(n12319), .A2(n10035), .ZN(n9355) );
  NAND2_X1 U11762 ( .A1(n9370), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9353) );
  INV_X1 U11763 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9352) );
  XNOR2_X1 U11764 ( .A(n9353), .B(n9352), .ZN(n10711) );
  NAND2_X1 U11765 ( .A1(n10421), .A2(n10711), .ZN(n9354) );
  NAND2_X1 U11766 ( .A1(n11309), .A2(n11203), .ZN(n12372) );
  INV_X1 U11767 ( .A(n11203), .ZN(n15264) );
  NAND2_X1 U11768 ( .A1(n15277), .A2(n15264), .ZN(n12373) );
  NAND2_X1 U11769 ( .A1(n12372), .A2(n12373), .ZN(n15256) );
  AND2_X1 U11770 ( .A1(n15277), .A2(n11203), .ZN(n9357) );
  NAND2_X1 U11771 ( .A1(n12302), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n9365) );
  NOR2_X1 U11772 ( .A1(n9358), .A2(n10681), .ZN(n9359) );
  OR2_X1 U11773 ( .A1(n9379), .A2(n9359), .ZN(n15252) );
  NAND2_X1 U11774 ( .A1(n9723), .A2(n15252), .ZN(n9364) );
  INV_X1 U11775 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n9360) );
  OR2_X1 U11776 ( .A1(n12304), .A2(n9360), .ZN(n9363) );
  INV_X1 U11777 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n9361) );
  OR2_X1 U11778 ( .A1(n9304), .A2(n9361), .ZN(n9362) );
  NAND4_X1 U11779 ( .A1(n9365), .A2(n9364), .A3(n9363), .A4(n9362), .ZN(n12522) );
  NAND2_X1 U11780 ( .A1(n10075), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9389) );
  NAND2_X1 U11781 ( .A1(n10235), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n9369) );
  NAND2_X1 U11782 ( .A1(n9389), .A2(n9369), .ZN(n9386) );
  XNOR2_X1 U11783 ( .A(n9388), .B(n9386), .ZN(n10024) );
  NAND2_X1 U11784 ( .A1(n12318), .A2(n10024), .ZN(n9374) );
  NAND2_X1 U11785 ( .A1(n12319), .A2(SI_8_), .ZN(n9373) );
  NAND2_X1 U11786 ( .A1(n9395), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9371) );
  XNOR2_X1 U11787 ( .A(n9371), .B(P3_IR_REG_8__SCAN_IN), .ZN(n12531) );
  NAND2_X1 U11788 ( .A1(n10421), .A2(n12531), .ZN(n9372) );
  XNOR2_X1 U11789 ( .A(n12522), .B(n15251), .ZN(n15246) );
  NAND2_X1 U11790 ( .A1(n15245), .A2(n15246), .ZN(n15244) );
  NAND2_X1 U11791 ( .A1(n15259), .A2(n15251), .ZN(n9375) );
  NAND2_X1 U11792 ( .A1(n15244), .A2(n9375), .ZN(n9376) );
  NAND2_X1 U11793 ( .A1(n9279), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9385) );
  INV_X1 U11794 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n9377) );
  OR2_X1 U11795 ( .A1(n9281), .A2(n9377), .ZN(n9384) );
  NAND2_X1 U11796 ( .A1(n9379), .A2(n9378), .ZN(n9402) );
  OR2_X1 U11797 ( .A1(n9379), .A2(n9378), .ZN(n9380) );
  AND2_X1 U11798 ( .A1(n9402), .A2(n9380), .ZN(n11478) );
  OR2_X1 U11799 ( .A1(n9262), .A2(n11478), .ZN(n9383) );
  INV_X1 U11800 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n9381) );
  OR2_X1 U11801 ( .A1(n9304), .A2(n9381), .ZN(n9382) );
  INV_X1 U11802 ( .A(n9386), .ZN(n9387) );
  NAND2_X1 U11803 ( .A1(n13553), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9409) );
  NAND2_X1 U11804 ( .A1(n10237), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9391) );
  AND2_X1 U11805 ( .A1(n9409), .A2(n9391), .ZN(n9392) );
  OR2_X1 U11806 ( .A1(n9393), .A2(n9392), .ZN(n9394) );
  NAND2_X1 U11807 ( .A1(n9410), .A2(n9394), .ZN(n10036) );
  NAND2_X1 U11808 ( .A1(n12318), .A2(n10036), .ZN(n9399) );
  INV_X1 U11809 ( .A(SI_9_), .ZN(n10037) );
  NAND2_X1 U11810 ( .A1(n12319), .A2(n10037), .ZN(n9398) );
  NOR2_X1 U11811 ( .A1(n9395), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9413) );
  OR2_X1 U11812 ( .A1(n9413), .A2(n9231), .ZN(n9396) );
  XNOR2_X1 U11813 ( .A(n9396), .B(n9412), .ZN(n15124) );
  NAND2_X1 U11814 ( .A1(n10421), .A2(n15124), .ZN(n9397) );
  NAND2_X1 U11815 ( .A1(n15233), .A2(n11480), .ZN(n12380) );
  INV_X1 U11816 ( .A(n11480), .ZN(n15369) );
  NAND2_X1 U11817 ( .A1(n15247), .A2(n15369), .ZN(n12381) );
  NAND2_X1 U11818 ( .A1(n15247), .A2(n11480), .ZN(n9401) );
  NAND2_X1 U11819 ( .A1(n12302), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9408) );
  INV_X1 U11820 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12548) );
  OR2_X1 U11821 ( .A1(n9304), .A2(n12548), .ZN(n9407) );
  NAND2_X1 U11822 ( .A1(n9402), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9403) );
  AND2_X1 U11823 ( .A1(n9432), .A2(n9403), .ZN(n11450) );
  OR2_X1 U11824 ( .A1(n9262), .A2(n11450), .ZN(n9406) );
  INV_X1 U11825 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n9404) );
  OR2_X1 U11826 ( .A1(n12304), .A2(n9404), .ZN(n9405) );
  NAND2_X1 U11827 ( .A1(n10161), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9421) );
  INV_X1 U11828 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10159) );
  NAND2_X1 U11829 ( .A1(n10159), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n9411) );
  XNOR2_X1 U11830 ( .A(n9420), .B(n9419), .ZN(n10021) );
  NAND2_X1 U11831 ( .A1(n10021), .A2(n12318), .ZN(n9416) );
  INV_X1 U11832 ( .A(SI_10_), .ZN(n10020) );
  NAND2_X1 U11833 ( .A1(n9413), .A2(n9412), .ZN(n9427) );
  NAND2_X1 U11834 ( .A1(n9427), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9414) );
  AOI22_X1 U11835 ( .A1(n12319), .A2(n10020), .B1(n10421), .B2(n12571), .ZN(
        n9415) );
  NAND2_X1 U11836 ( .A1(n14425), .A2(n11454), .ZN(n12384) );
  INV_X1 U11837 ( .A(n11454), .ZN(n15238) );
  NAND2_X1 U11838 ( .A1(n12521), .A2(n15238), .ZN(n12385) );
  NAND2_X1 U11839 ( .A1(n12384), .A2(n12385), .ZN(n15232) );
  NAND2_X1 U11840 ( .A1(n12521), .A2(n11454), .ZN(n9417) );
  NAND2_X1 U11841 ( .A1(n9418), .A2(n9417), .ZN(n14421) );
  NAND2_X1 U11842 ( .A1(n9422), .A2(n9421), .ZN(n9425) );
  NAND2_X1 U11843 ( .A1(n10199), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9440) );
  NAND2_X1 U11844 ( .A1(n10202), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9423) );
  NAND2_X1 U11845 ( .A1(n9425), .A2(n9424), .ZN(n9441) );
  OR2_X1 U11846 ( .A1(n9425), .A2(n9424), .ZN(n9426) );
  NAND2_X1 U11847 ( .A1(n9441), .A2(n9426), .ZN(n10043) );
  OAI21_X1 U11848 ( .B1(n9427), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9429) );
  INV_X1 U11849 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9428) );
  XNOR2_X1 U11850 ( .A(n9429), .B(n9428), .ZN(n15163) );
  OAI22_X1 U11851 ( .A1(n9430), .A2(SI_11_), .B1(n12574), .B2(n9738), .ZN(
        n9431) );
  AOI21_X1 U11852 ( .B1(n10043), .B2(n12318), .A(n9431), .ZN(n11719) );
  NAND2_X1 U11853 ( .A1(n9432), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9433) );
  AND2_X1 U11854 ( .A1(n9451), .A2(n9433), .ZN(n11715) );
  OR2_X1 U11855 ( .A1(n9262), .A2(n11715), .ZN(n9439) );
  NAND2_X1 U11856 ( .A1(n12302), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n9438) );
  INV_X1 U11857 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n9434) );
  OR2_X1 U11858 ( .A1(n12304), .A2(n9434), .ZN(n9437) );
  INV_X1 U11859 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n9435) );
  OR2_X1 U11860 ( .A1(n9304), .A2(n9435), .ZN(n9436) );
  NAND4_X1 U11861 ( .A1(n9439), .A2(n9438), .A3(n9437), .A4(n9436), .ZN(n12520) );
  INV_X1 U11862 ( .A(n12520), .ZN(n15234) );
  INV_X1 U11863 ( .A(n11719), .ZN(n14427) );
  NAND2_X1 U11864 ( .A1(n15234), .A2(n14427), .ZN(n11618) );
  NAND2_X1 U11865 ( .A1(n9441), .A2(n9440), .ZN(n9444) );
  NAND2_X1 U11866 ( .A1(n10312), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9458) );
  NAND2_X1 U11867 ( .A1(n10315), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n9442) );
  OR2_X1 U11868 ( .A1(n9444), .A2(n9443), .ZN(n9445) );
  NAND2_X1 U11869 ( .A1(n9459), .A2(n9445), .ZN(n10055) );
  OR2_X1 U11870 ( .A1(n10055), .A2(n9603), .ZN(n9449) );
  NAND2_X1 U11871 ( .A1(n9446), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9447) );
  XNOR2_X1 U11872 ( .A(n9447), .B(P3_IR_REG_12__SCAN_IN), .ZN(n12529) );
  AOI22_X1 U11873 ( .A1(n12319), .A2(SI_12_), .B1(n10421), .B2(n12529), .ZN(
        n9448) );
  NAND2_X1 U11874 ( .A1(n9449), .A2(n9448), .ZN(n11736) );
  NAND2_X1 U11875 ( .A1(n9279), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9456) );
  INV_X1 U11876 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n9450) );
  OR2_X1 U11877 ( .A1(n9281), .A2(n9450), .ZN(n9455) );
  AND2_X1 U11878 ( .A1(n9451), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9452) );
  NOR2_X1 U11879 ( .A1(n9469), .A2(n9452), .ZN(n11731) );
  OR2_X1 U11880 ( .A1(n9262), .A2(n11731), .ZN(n9454) );
  INV_X1 U11881 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11626) );
  OR2_X1 U11882 ( .A1(n9304), .A2(n11626), .ZN(n9453) );
  OR2_X1 U11883 ( .A1(n11736), .A2(n14426), .ZN(n12394) );
  NAND2_X1 U11884 ( .A1(n11736), .A2(n14426), .ZN(n12393) );
  NAND2_X1 U11885 ( .A1(n12394), .A2(n12393), .ZN(n11621) );
  AND2_X1 U11886 ( .A1(n11618), .A2(n11621), .ZN(n9457) );
  NAND2_X1 U11887 ( .A1(n9461), .A2(n10319), .ZN(n9462) );
  NAND2_X1 U11888 ( .A1(n9477), .A2(n9462), .ZN(n10077) );
  NAND2_X1 U11889 ( .A1(n10077), .A2(n12318), .ZN(n9467) );
  OR2_X1 U11890 ( .A1(n9463), .A2(n9231), .ZN(n9465) );
  XNOR2_X1 U11891 ( .A(n9465), .B(n9464), .ZN(n15199) );
  AOI22_X1 U11892 ( .A1(n12319), .A2(n13723), .B1(n10421), .B2(n15199), .ZN(
        n9466) );
  NAND2_X1 U11893 ( .A1(n9467), .A2(n9466), .ZN(n11816) );
  OR2_X1 U11894 ( .A1(n9469), .A2(n9468), .ZN(n9470) );
  NAND2_X1 U11895 ( .A1(n9469), .A2(n9468), .ZN(n9486) );
  AND2_X1 U11896 ( .A1(n9470), .A2(n9486), .ZN(n11668) );
  OR2_X1 U11897 ( .A1(n9262), .A2(n11668), .ZN(n9474) );
  NAND2_X1 U11898 ( .A1(n12302), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9473) );
  INV_X1 U11899 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n11779) );
  OR2_X1 U11900 ( .A1(n12304), .A2(n11779), .ZN(n9472) );
  INV_X1 U11901 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n15194) );
  OR2_X1 U11902 ( .A1(n9304), .A2(n15194), .ZN(n9471) );
  NAND4_X1 U11903 ( .A1(n9474), .A2(n9473), .A3(n9472), .A4(n9471), .ZN(n12518) );
  OR2_X1 U11904 ( .A1(n11816), .A2(n12518), .ZN(n12399) );
  NAND2_X1 U11905 ( .A1(n11816), .A2(n12518), .ZN(n12400) );
  NAND2_X1 U11906 ( .A1(n12399), .A2(n12400), .ZN(n12490) );
  INV_X1 U11907 ( .A(n12518), .ZN(n12127) );
  OR2_X1 U11908 ( .A1(n11816), .A2(n12127), .ZN(n9475) );
  NAND2_X1 U11909 ( .A1(n11663), .A2(n9475), .ZN(n11740) );
  NAND2_X1 U11910 ( .A1(n10414), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9493) );
  NAND2_X1 U11911 ( .A1(n10416), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9478) );
  OR2_X1 U11912 ( .A1(n9480), .A2(n9479), .ZN(n9481) );
  NAND2_X1 U11913 ( .A1(n9494), .A2(n9481), .ZN(n10162) );
  NAND2_X1 U11914 ( .A1(n10162), .A2(n12318), .ZN(n9485) );
  OR2_X1 U11915 ( .A1(n9482), .A2(n9231), .ZN(n9483) );
  XNOR2_X1 U11916 ( .A(n9483), .B(n9496), .ZN(n15217) );
  AOI22_X1 U11917 ( .A1(n12319), .A2(n10163), .B1(n10421), .B2(n15217), .ZN(
        n9484) );
  NAND2_X1 U11918 ( .A1(n9486), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9487) );
  AND2_X1 U11919 ( .A1(n9503), .A2(n9487), .ZN(n12179) );
  OR2_X1 U11920 ( .A1(n9262), .A2(n12179), .ZN(n9491) );
  NAND2_X1 U11921 ( .A1(n12302), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9490) );
  INV_X1 U11922 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12946) );
  OR2_X1 U11923 ( .A1(n12304), .A2(n12946), .ZN(n9489) );
  INV_X1 U11924 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n11744) );
  OR2_X1 U11925 ( .A1(n9304), .A2(n11744), .ZN(n9488) );
  NAND4_X1 U11926 ( .A1(n9491), .A2(n9490), .A3(n9489), .A4(n9488), .ZN(n12517) );
  OR2_X1 U11927 ( .A1(n12948), .A2(n12517), .ZN(n12405) );
  NAND2_X1 U11928 ( .A1(n12948), .A2(n12517), .ZN(n12404) );
  NAND2_X1 U11929 ( .A1(n12405), .A2(n12404), .ZN(n12489) );
  INV_X1 U11930 ( .A(n12517), .ZN(n12806) );
  OR2_X1 U11931 ( .A1(n12948), .A2(n12806), .ZN(n9492) );
  NAND2_X1 U11932 ( .A1(n10717), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9512) );
  NAND2_X1 U11933 ( .A1(n10719), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n9495) );
  XNOR2_X1 U11934 ( .A(n9511), .B(n9510), .ZN(n14324) );
  NAND2_X1 U11935 ( .A1(n14324), .A2(n12318), .ZN(n9502) );
  NAND2_X1 U11936 ( .A1(n9482), .A2(n9496), .ZN(n9497) );
  NAND2_X1 U11937 ( .A1(n9497), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9499) );
  INV_X1 U11938 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9498) );
  XNOR2_X1 U11939 ( .A(n9499), .B(n9498), .ZN(n14328) );
  AOI22_X1 U11940 ( .A1(n12319), .A2(n9500), .B1(n10421), .B2(n14328), .ZN(
        n9501) );
  NAND2_X1 U11941 ( .A1(n9279), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9508) );
  INV_X1 U11942 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12890) );
  OR2_X1 U11943 ( .A1(n9281), .A2(n12890), .ZN(n9507) );
  AND2_X1 U11944 ( .A1(n9503), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9504) );
  NOR2_X1 U11945 ( .A1(n9523), .A2(n9504), .ZN(n12290) );
  OR2_X1 U11946 ( .A1(n9262), .A2(n12290), .ZN(n9506) );
  INV_X1 U11947 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14352) );
  OR2_X1 U11948 ( .A1(n9304), .A2(n14352), .ZN(n9505) );
  NAND2_X1 U11949 ( .A1(n12944), .A2(n12175), .ZN(n9509) );
  NAND2_X1 U11950 ( .A1(n9511), .A2(n9510), .ZN(n9513) );
  NAND2_X1 U11951 ( .A1(n9513), .A2(n9512), .ZN(n9516) );
  NAND2_X1 U11952 ( .A1(n10773), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9532) );
  NAND2_X1 U11953 ( .A1(n10774), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n9514) );
  OR2_X1 U11954 ( .A1(n9516), .A2(n9515), .ZN(n9517) );
  NAND2_X1 U11955 ( .A1(n9533), .A2(n9517), .ZN(n10259) );
  OR2_X1 U11956 ( .A1(n10259), .A2(n9603), .ZN(n9521) );
  OR2_X1 U11957 ( .A1(n9536), .A2(n9231), .ZN(n9519) );
  XNOR2_X1 U11958 ( .A(n9519), .B(P3_IR_REG_16__SCAN_IN), .ZN(n14372) );
  AOI22_X1 U11959 ( .A1(n12319), .A2(SI_16_), .B1(n10421), .B2(n14372), .ZN(
        n9520) );
  NAND2_X1 U11960 ( .A1(n9521), .A2(n9520), .ZN(n12884) );
  NOR2_X1 U11961 ( .A1(n9523), .A2(n9522), .ZN(n9524) );
  OR2_X1 U11962 ( .A1(n9543), .A2(n9524), .ZN(n12799) );
  NAND2_X1 U11963 ( .A1(n9723), .A2(n12799), .ZN(n9529) );
  INV_X1 U11964 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12541) );
  OR2_X1 U11965 ( .A1(n9281), .A2(n12541), .ZN(n9528) );
  INV_X1 U11966 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n9525) );
  OR2_X1 U11967 ( .A1(n12304), .A2(n9525), .ZN(n9527) );
  OR2_X1 U11968 ( .A1(n9304), .A2(n12557), .ZN(n9526) );
  OR2_X1 U11969 ( .A1(n12884), .A2(n12807), .ZN(n12414) );
  NAND2_X1 U11970 ( .A1(n12884), .A2(n12807), .ZN(n12782) );
  NAND2_X1 U11971 ( .A1(n12414), .A2(n12782), .ZN(n12491) );
  NAND2_X1 U11972 ( .A1(n12790), .A2(n12491), .ZN(n9531) );
  NAND2_X1 U11973 ( .A1(n12884), .A2(n12516), .ZN(n9530) );
  NAND2_X1 U11974 ( .A1(n9531), .A2(n9530), .ZN(n12778) );
  NAND2_X1 U11975 ( .A1(n10893), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9551) );
  NAND2_X1 U11976 ( .A1(n13735), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n9534) );
  XNOR2_X1 U11977 ( .A(n9550), .B(n9549), .ZN(n10317) );
  NAND2_X1 U11978 ( .A1(n10317), .A2(n12318), .ZN(n9542) );
  NAND2_X1 U11979 ( .A1(n9538), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9537) );
  MUX2_X1 U11980 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9537), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n9540) );
  NAND2_X1 U11981 ( .A1(n9540), .A2(n9570), .ZN(n14397) );
  AOI22_X1 U11982 ( .A1(n12319), .A2(n10316), .B1(n10421), .B2(n14397), .ZN(
        n9541) );
  NAND2_X1 U11983 ( .A1(n12302), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9548) );
  OR2_X1 U11984 ( .A1(n9543), .A2(n12235), .ZN(n9544) );
  NAND2_X1 U11985 ( .A1(n9556), .A2(n9544), .ZN(n12785) );
  NAND2_X1 U11986 ( .A1(n9723), .A2(n12785), .ZN(n9547) );
  INV_X1 U11987 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12937) );
  OR2_X1 U11988 ( .A1(n12304), .A2(n12937), .ZN(n9546) );
  INV_X1 U11989 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14389) );
  OR2_X1 U11990 ( .A1(n9304), .A2(n14389), .ZN(n9545) );
  NAND4_X1 U11991 ( .A1(n9548), .A2(n9547), .A3(n9546), .A4(n9545), .ZN(n12792) );
  OR2_X1 U11992 ( .A1(n12939), .A2(n12792), .ZN(n12420) );
  NAND2_X1 U11993 ( .A1(n12939), .A2(n12792), .ZN(n12773) );
  NAND2_X1 U11994 ( .A1(n12420), .A2(n12773), .ZN(n12779) );
  INV_X1 U11995 ( .A(n12792), .ZN(n12228) );
  NAND2_X1 U11996 ( .A1(n11132), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9567) );
  NAND2_X1 U11997 ( .A1(n11135), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n9552) );
  NAND2_X1 U11998 ( .A1(n9567), .A2(n9552), .ZN(n9564) );
  XNOR2_X1 U11999 ( .A(n9566), .B(n9564), .ZN(n10403) );
  NAND2_X1 U12000 ( .A1(n10403), .A2(n12318), .ZN(n9555) );
  NAND2_X1 U12001 ( .A1(n9570), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9553) );
  XNOR2_X1 U12002 ( .A(n9553), .B(P3_IR_REG_18__SCAN_IN), .ZN(n14404) );
  AOI22_X1 U12003 ( .A1(n12319), .A2(SI_18_), .B1(n10421), .B2(n14404), .ZN(
        n9554) );
  NAND2_X1 U12004 ( .A1(n9555), .A2(n9554), .ZN(n12765) );
  NAND2_X1 U12005 ( .A1(n9556), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9557) );
  NAND2_X1 U12006 ( .A1(n9576), .A2(n9557), .ZN(n12766) );
  NAND2_X1 U12007 ( .A1(n12766), .A2(n9723), .ZN(n9561) );
  NAND2_X1 U12008 ( .A1(n9279), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9560) );
  NAND2_X1 U12009 ( .A1(n9741), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9559) );
  INV_X1 U12010 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12563) );
  OR2_X1 U12011 ( .A1(n9281), .A2(n12563), .ZN(n9558) );
  OR2_X1 U12012 ( .A1(n12765), .A2(n12781), .ZN(n12418) );
  NAND2_X1 U12013 ( .A1(n12765), .A2(n12781), .ZN(n12422) );
  OR2_X1 U12014 ( .A1(n12765), .A2(n12751), .ZN(n9563) );
  INV_X1 U12015 ( .A(n9564), .ZN(n9565) );
  NAND2_X1 U12016 ( .A1(n13560), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9584) );
  INV_X1 U12017 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11193) );
  NAND2_X1 U12018 ( .A1(n11193), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9569) );
  NAND2_X1 U12019 ( .A1(n9584), .A2(n9569), .ZN(n9581) );
  XNOR2_X1 U12020 ( .A(n9583), .B(n9581), .ZN(n10510) );
  NAND2_X1 U12021 ( .A1(n10510), .A2(n12318), .ZN(n9575) );
  NAND2_X1 U12022 ( .A1(n9730), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9573) );
  XNOR2_X2 U12023 ( .A(n9573), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12608) );
  AOI22_X1 U12024 ( .A1(n12319), .A2(SI_19_), .B1(n10421), .B2(n12608), .ZN(
        n9574) );
  NAND2_X1 U12025 ( .A1(n9575), .A2(n9574), .ZN(n12189) );
  AND2_X1 U12026 ( .A1(n9576), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9577) );
  OR2_X1 U12027 ( .A1(n9577), .A2(n9590), .ZN(n12756) );
  NAND2_X1 U12028 ( .A1(n12756), .A2(n9723), .ZN(n9580) );
  AOI22_X1 U12029 ( .A1(n9741), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n12302), 
        .B2(P3_REG1_REG_19__SCAN_IN), .ZN(n9579) );
  NAND2_X1 U12030 ( .A1(n9279), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9578) );
  OR2_X1 U12031 ( .A1(n12189), .A2(n12741), .ZN(n12429) );
  NAND2_X1 U12032 ( .A1(n12189), .A2(n12741), .ZN(n12430) );
  INV_X1 U12033 ( .A(n9581), .ZN(n9582) );
  NAND2_X1 U12034 ( .A1(n9586), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9587) );
  NAND2_X1 U12035 ( .A1(n9598), .A2(n9587), .ZN(n10752) );
  NAND2_X1 U12036 ( .A1(n12319), .A2(SI_20_), .ZN(n9588) );
  NOR2_X1 U12037 ( .A1(n9590), .A2(n12258), .ZN(n9591) );
  OR2_X1 U12038 ( .A1(n9607), .A2(n9591), .ZN(n12745) );
  NAND2_X1 U12039 ( .A1(n12745), .A2(n9723), .ZN(n9594) );
  AOI22_X1 U12040 ( .A1(n9741), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n12302), 
        .B2(P3_REG1_REG_20__SCAN_IN), .ZN(n9593) );
  NAND2_X1 U12041 ( .A1(n9279), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9592) );
  NAND2_X1 U12042 ( .A1(n12253), .A2(n12730), .ZN(n12435) );
  NAND2_X1 U12043 ( .A1(n12434), .A2(n12435), .ZN(n12744) );
  NAND2_X1 U12044 ( .A1(n12739), .A2(n12744), .ZN(n9596) );
  NAND2_X1 U12045 ( .A1(n12253), .A2(n12752), .ZN(n9595) );
  NAND2_X1 U12046 ( .A1(n11359), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9615) );
  NAND2_X1 U12047 ( .A1(n11374), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9599) );
  OR2_X1 U12048 ( .A1(n9601), .A2(n9600), .ZN(n9602) );
  NAND2_X1 U12049 ( .A1(n9616), .A2(n9602), .ZN(n10934) );
  NAND2_X1 U12050 ( .A1(n12319), .A2(SI_21_), .ZN(n9604) );
  INV_X1 U12051 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9606) );
  OR2_X1 U12052 ( .A1(n9607), .A2(n9606), .ZN(n9608) );
  NAND2_X1 U12053 ( .A1(n9619), .A2(n9608), .ZN(n12734) );
  INV_X1 U12054 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n9611) );
  NAND2_X1 U12055 ( .A1(n12302), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9610) );
  NAND2_X1 U12056 ( .A1(n9279), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n9609) );
  OAI211_X1 U12057 ( .C1(n9611), .C2(n9304), .A(n9610), .B(n9609), .ZN(n9612)
         );
  OR2_X1 U12058 ( .A1(n12209), .A2(n12742), .ZN(n12335) );
  NAND2_X1 U12059 ( .A1(n12209), .A2(n12742), .ZN(n12334) );
  OR2_X1 U12060 ( .A1(n12209), .A2(n12515), .ZN(n9614) );
  XNOR2_X1 U12061 ( .A(n11591), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n9629) );
  XNOR2_X1 U12062 ( .A(n9630), .B(n9629), .ZN(n11060) );
  NAND2_X1 U12063 ( .A1(n11060), .A2(n12318), .ZN(n9618) );
  NAND2_X1 U12064 ( .A1(n12319), .A2(SI_22_), .ZN(n9617) );
  NAND2_X1 U12065 ( .A1(n9619), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9620) );
  NAND2_X1 U12066 ( .A1(n9632), .A2(n9620), .ZN(n12721) );
  NAND2_X1 U12067 ( .A1(n12721), .A2(n9723), .ZN(n9626) );
  INV_X1 U12068 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n9623) );
  NAND2_X1 U12069 ( .A1(n9279), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n9622) );
  NAND2_X1 U12070 ( .A1(n12302), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9621) );
  OAI211_X1 U12071 ( .C1(n9623), .C2(n9304), .A(n9622), .B(n9621), .ZN(n9624)
         );
  INV_X1 U12072 ( .A(n9624), .ZN(n9625) );
  NAND2_X1 U12073 ( .A1(n12720), .A2(n12701), .ZN(n9627) );
  NAND2_X1 U12074 ( .A1(n11591), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9628) );
  XNOR2_X1 U12075 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n9641) );
  NAND2_X1 U12076 ( .A1(n12319), .A2(SI_23_), .ZN(n9631) );
  NAND2_X1 U12077 ( .A1(n9632), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9633) );
  NAND2_X1 U12078 ( .A1(n9647), .A2(n9633), .ZN(n12710) );
  NAND2_X1 U12079 ( .A1(n12710), .A2(n9723), .ZN(n9639) );
  INV_X1 U12080 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n9636) );
  NAND2_X1 U12081 ( .A1(n9279), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9635) );
  NAND2_X1 U12082 ( .A1(n12302), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9634) );
  OAI211_X1 U12083 ( .C1(n9636), .C2(n9304), .A(n9635), .B(n9634), .ZN(n9637)
         );
  INV_X1 U12084 ( .A(n9637), .ZN(n9638) );
  NAND2_X1 U12085 ( .A1(n12705), .A2(n12687), .ZN(n9640) );
  NAND2_X1 U12086 ( .A1(n12699), .A2(n9640), .ZN(n12665) );
  NAND2_X1 U12087 ( .A1(n9643), .A2(n13595), .ZN(n9644) );
  NAND2_X1 U12088 ( .A1(n9655), .A2(n9644), .ZN(n9656) );
  XNOR2_X1 U12089 ( .A(n9656), .B(n11694), .ZN(n11375) );
  NAND2_X1 U12090 ( .A1(n11375), .A2(n12318), .ZN(n9646) );
  NAND2_X1 U12091 ( .A1(n12319), .A2(SI_24_), .ZN(n9645) );
  INV_X1 U12092 ( .A(n9660), .ZN(n9649) );
  NAND2_X1 U12093 ( .A1(n9647), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9648) );
  NAND2_X1 U12094 ( .A1(n9649), .A2(n9648), .ZN(n12691) );
  NAND2_X1 U12095 ( .A1(n12691), .A2(n9723), .ZN(n9654) );
  INV_X1 U12096 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12692) );
  NAND2_X1 U12097 ( .A1(n9279), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9651) );
  NAND2_X1 U12098 ( .A1(n12302), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9650) );
  OAI211_X1 U12099 ( .C1(n12692), .C2(n9304), .A(n9651), .B(n9650), .ZN(n9652)
         );
  INV_X1 U12100 ( .A(n9652), .ZN(n9653) );
  XNOR2_X1 U12101 ( .A(n12849), .B(n12244), .ZN(n12686) );
  XNOR2_X1 U12102 ( .A(n13775), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n9657) );
  XNOR2_X1 U12103 ( .A(n9671), .B(n9657), .ZN(n11501) );
  NAND2_X1 U12104 ( .A1(n11501), .A2(n12318), .ZN(n9659) );
  NAND2_X1 U12105 ( .A1(n12319), .A2(SI_25_), .ZN(n9658) );
  NAND2_X1 U12106 ( .A1(n9660), .A2(n13624), .ZN(n9676) );
  OR2_X1 U12107 ( .A1(n9660), .A2(n13624), .ZN(n9661) );
  NAND2_X1 U12108 ( .A1(n9676), .A2(n9661), .ZN(n12675) );
  NAND2_X1 U12109 ( .A1(n12675), .A2(n9723), .ZN(n9667) );
  INV_X1 U12110 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n9664) );
  NAND2_X1 U12111 ( .A1(n9279), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9663) );
  NAND2_X1 U12112 ( .A1(n12302), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9662) );
  OAI211_X1 U12113 ( .C1(n9664), .C2(n9304), .A(n9663), .B(n9662), .ZN(n9665)
         );
  INV_X1 U12114 ( .A(n9665), .ZN(n9666) );
  XNOR2_X1 U12115 ( .A(n12845), .B(n12653), .ZN(n12669) );
  AND2_X1 U12116 ( .A1(n12686), .A2(n12669), .ZN(n9668) );
  INV_X1 U12117 ( .A(n12669), .ZN(n12673) );
  NAND2_X1 U12118 ( .A1(n12849), .A2(n12702), .ZN(n12666) );
  NAND2_X1 U12119 ( .A1(n12845), .A2(n12688), .ZN(n9669) );
  NAND2_X1 U12120 ( .A1(n12667), .A2(n9669), .ZN(n12651) );
  NAND2_X1 U12121 ( .A1(n13775), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9670) );
  NAND2_X1 U12122 ( .A1(n14302), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9672) );
  XNOR2_X1 U12123 ( .A(n9688), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n9673) );
  XNOR2_X1 U12124 ( .A(n9687), .B(n9673), .ZN(n11607) );
  NAND2_X1 U12125 ( .A1(n11607), .A2(n12318), .ZN(n9675) );
  NAND2_X1 U12126 ( .A1(n12319), .A2(SI_26_), .ZN(n9674) );
  NAND2_X1 U12127 ( .A1(n9676), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9677) );
  NAND2_X1 U12128 ( .A1(n9693), .A2(n9677), .ZN(n12658) );
  NAND2_X1 U12129 ( .A1(n12658), .A2(n9723), .ZN(n9682) );
  INV_X1 U12130 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12660) );
  NAND2_X1 U12131 ( .A1(n9279), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9679) );
  NAND2_X1 U12132 ( .A1(n12302), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9678) );
  OAI211_X1 U12133 ( .C1(n12660), .C2(n9304), .A(n9679), .B(n9678), .ZN(n9680)
         );
  INV_X1 U12134 ( .A(n9680), .ZN(n9681) );
  OR2_X1 U12135 ( .A1(n12840), .A2(n12670), .ZN(n9683) );
  NAND2_X1 U12136 ( .A1(n12840), .A2(n12670), .ZN(n9684) );
  AND2_X1 U12137 ( .A1(n14299), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9686) );
  NAND2_X1 U12138 ( .A1(n9688), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9689) );
  XNOR2_X1 U12139 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n9690) );
  XNOR2_X1 U12140 ( .A(n9704), .B(n9690), .ZN(n11632) );
  NAND2_X1 U12141 ( .A1(n11632), .A2(n12318), .ZN(n9692) );
  NAND2_X1 U12142 ( .A1(n12319), .A2(SI_27_), .ZN(n9691) );
  INV_X1 U12143 ( .A(n9710), .ZN(n9695) );
  NAND2_X1 U12144 ( .A1(n9693), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9694) );
  NAND2_X1 U12145 ( .A1(n9695), .A2(n9694), .ZN(n12644) );
  NAND2_X1 U12146 ( .A1(n12644), .A2(n9723), .ZN(n9701) );
  INV_X1 U12147 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n9698) );
  NAND2_X1 U12148 ( .A1(n9279), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9697) );
  NAND2_X1 U12149 ( .A1(n12302), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9696) );
  OAI211_X1 U12150 ( .C1(n9698), .C2(n9304), .A(n9697), .B(n9696), .ZN(n9699)
         );
  INV_X1 U12151 ( .A(n9699), .ZN(n9700) );
  NAND2_X1 U12152 ( .A1(n12836), .A2(n12654), .ZN(n12450) );
  OR2_X1 U12153 ( .A1(n12836), .A2(n12654), .ZN(n9702) );
  AND2_X2 U12154 ( .A1(n12450), .A2(n9702), .ZN(n12640) );
  INV_X1 U12155 ( .A(n12640), .ZN(n9703) );
  NAND2_X1 U12156 ( .A1(n14296), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9705) );
  XNOR2_X1 U12157 ( .A(n9719), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n9706) );
  XNOR2_X1 U12158 ( .A(n9716), .B(n9706), .ZN(n11722) );
  NAND2_X1 U12159 ( .A1(n11722), .A2(n12318), .ZN(n9708) );
  NAND2_X1 U12160 ( .A1(n12319), .A2(SI_28_), .ZN(n9707) );
  INV_X1 U12161 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n9709) );
  NOR2_X1 U12162 ( .A1(n9710), .A2(n9709), .ZN(n9711) );
  INV_X1 U12163 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13549) );
  NAND2_X1 U12164 ( .A1(n12302), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9713) );
  NAND2_X1 U12165 ( .A1(n9741), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9712) );
  OAI211_X1 U12166 ( .C1(n12304), .C2(n13549), .A(n9713), .B(n9712), .ZN(n9714) );
  AOI21_X2 U12167 ( .B1(n12626), .B2(n9723), .A(n9714), .ZN(n12637) );
  OR2_X1 U12168 ( .A1(n12836), .A2(n12514), .ZN(n9838) );
  AND2_X1 U12169 ( .A1(n12455), .A2(n9838), .ZN(n9715) );
  NAND2_X1 U12170 ( .A1(n9837), .A2(n7527), .ZN(n9729) );
  INV_X1 U12171 ( .A(n9716), .ZN(n9718) );
  NAND2_X1 U12172 ( .A1(n11877), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9717) );
  NAND2_X1 U12173 ( .A1(n9719), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9720) );
  XNOR2_X1 U12174 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n11866) );
  XNOR2_X1 U12175 ( .A(n11869), .B(n11866), .ZN(n12957) );
  NAND2_X1 U12176 ( .A1(n12957), .A2(n12318), .ZN(n9722) );
  NAND2_X1 U12177 ( .A1(n12319), .A2(SI_29_), .ZN(n9721) );
  NAND2_X1 U12178 ( .A1(n9722), .A2(n9721), .ZN(n9817) );
  NAND2_X1 U12179 ( .A1(n12618), .A2(n9723), .ZN(n12310) );
  INV_X1 U12180 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n9726) );
  NAND2_X1 U12181 ( .A1(n12302), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9725) );
  NAND2_X1 U12182 ( .A1(n9279), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9724) );
  OAI211_X1 U12183 ( .C1(n9304), .C2(n9726), .A(n9725), .B(n9724), .ZN(n9727)
         );
  INV_X1 U12184 ( .A(n9727), .ZN(n9728) );
  OR2_X1 U12185 ( .A1(n9817), .A2(n12205), .ZN(n12465) );
  NAND2_X1 U12186 ( .A1(n9817), .A2(n12205), .ZN(n12464) );
  NAND2_X1 U12187 ( .A1(n12465), .A2(n12464), .ZN(n12462) );
  XNOR2_X1 U12188 ( .A(n9729), .B(n12462), .ZN(n9748) );
  NAND2_X1 U12189 ( .A1(n12509), .A2(n12608), .ZN(n9821) );
  NAND2_X1 U12190 ( .A1(n9736), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9737) );
  NAND2_X1 U12191 ( .A1(n12340), .A2(n9820), .ZN(n12323) );
  INV_X1 U12192 ( .A(n12507), .ZN(n10420) );
  INV_X1 U12193 ( .A(n12589), .ZN(n12600) );
  NAND2_X1 U12194 ( .A1(n10420), .A2(n12600), .ZN(n10423) );
  NAND2_X1 U12195 ( .A1(n10423), .A2(n9738), .ZN(n10839) );
  INV_X1 U12196 ( .A(P3_B_REG_SCAN_IN), .ZN(n9739) );
  NOR2_X1 U12197 ( .A1(n12507), .A2(n9739), .ZN(n9740) );
  OR2_X1 U12198 ( .A1(n15294), .A2(n9740), .ZN(n12611) );
  INV_X1 U12199 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n13633) );
  NAND2_X1 U12200 ( .A1(n9279), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9743) );
  NAND2_X1 U12201 ( .A1(n9741), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9742) );
  OAI211_X1 U12202 ( .C1(n9281), .C2(n13633), .A(n9743), .B(n9742), .ZN(n9744)
         );
  INV_X1 U12203 ( .A(n9744), .ZN(n9745) );
  INV_X1 U12204 ( .A(n10658), .ZN(n10575) );
  NAND2_X1 U12205 ( .A1(n10825), .A2(n12341), .ZN(n15308) );
  NAND2_X1 U12206 ( .A1(n9749), .A2(n12344), .ZN(n10920) );
  NAND2_X1 U12207 ( .A1(n10920), .A2(n12480), .ZN(n15287) );
  AND2_X1 U12208 ( .A1(n15286), .A2(n12356), .ZN(n9752) );
  NAND2_X1 U12209 ( .A1(n11227), .A2(n12358), .ZN(n15270) );
  NAND2_X1 U12210 ( .A1(n15295), .A2(n11000), .ZN(n15271) );
  AND2_X1 U12211 ( .A1(n15271), .A2(n12366), .ZN(n9753) );
  INV_X1 U12212 ( .A(n12366), .ZN(n12363) );
  NAND2_X1 U12213 ( .A1(n15263), .A2(n15262), .ZN(n9754) );
  NAND2_X1 U12214 ( .A1(n9754), .A2(n12372), .ZN(n15243) );
  NAND2_X1 U12215 ( .A1(n15243), .A2(n15242), .ZN(n9756) );
  INV_X1 U12216 ( .A(n15251), .ZN(n9755) );
  NAND2_X1 U12217 ( .A1(n15259), .A2(n9755), .ZN(n12377) );
  INV_X1 U12218 ( .A(n12380), .ZN(n9757) );
  INV_X1 U12219 ( .A(n12385), .ZN(n9758) );
  NAND2_X1 U12220 ( .A1(n15234), .A2(n11719), .ZN(n12390) );
  NAND2_X1 U12221 ( .A1(n12520), .A2(n14427), .ZN(n12389) );
  NAND2_X1 U12222 ( .A1(n9759), .A2(n12390), .ZN(n11628) );
  INV_X1 U12223 ( .A(n11621), .ZN(n12485) );
  NAND2_X1 U12224 ( .A1(n11628), .A2(n12485), .ZN(n9760) );
  NAND2_X1 U12225 ( .A1(n9760), .A2(n12393), .ZN(n11667) );
  INV_X1 U12226 ( .A(n12399), .ZN(n9761) );
  NAND2_X1 U12227 ( .A1(n12944), .A2(n12791), .ZN(n12409) );
  INV_X1 U12228 ( .A(n12491), .ZN(n12798) );
  AND2_X1 U12229 ( .A1(n12808), .A2(n12798), .ZN(n9763) );
  AOI21_X2 U12230 ( .B1(n12809), .B2(n9763), .A(n6617), .ZN(n12796) );
  AND2_X1 U12231 ( .A1(n12782), .A2(n12420), .ZN(n12772) );
  AND2_X1 U12232 ( .A1(n12772), .A2(n12492), .ZN(n9764) );
  NAND2_X1 U12233 ( .A1(n12796), .A2(n9764), .ZN(n12771) );
  OR2_X1 U12234 ( .A1(n9562), .A2(n12773), .ZN(n12770) );
  AND2_X1 U12235 ( .A1(n12418), .A2(n12770), .ZN(n9765) );
  NAND2_X1 U12236 ( .A1(n12771), .A2(n9765), .ZN(n12755) );
  INV_X1 U12237 ( .A(n12755), .ZN(n9766) );
  NAND2_X1 U12238 ( .A1(n12733), .A2(n12334), .ZN(n9767) );
  NAND2_X1 U12239 ( .A1(n12720), .A2(n12731), .ZN(n12332) );
  INV_X1 U12240 ( .A(n12686), .ZN(n12681) );
  OR2_X1 U12241 ( .A1(n12717), .A2(n12705), .ZN(n12682) );
  AND2_X1 U12242 ( .A1(n12681), .A2(n12682), .ZN(n12327) );
  NAND2_X1 U12243 ( .A1(n12849), .A2(n12244), .ZN(n12325) );
  NAND2_X1 U12244 ( .A1(n12680), .A2(n12325), .ZN(n12674) );
  NAND2_X1 U12245 ( .A1(n12674), .A2(n12673), .ZN(n9768) );
  NAND2_X1 U12246 ( .A1(n12845), .A2(n12653), .ZN(n12328) );
  NAND2_X1 U12247 ( .A1(n12650), .A2(n12449), .ZN(n9769) );
  NAND2_X1 U12248 ( .A1(n12840), .A2(n12636), .ZN(n12457) );
  NAND2_X1 U12249 ( .A1(n9769), .A2(n12457), .ZN(n12641) );
  NAND2_X1 U12250 ( .A1(n12641), .A2(n12640), .ZN(n12643) );
  NAND2_X1 U12251 ( .A1(n12643), .A2(n12450), .ZN(n9770) );
  NAND2_X1 U12252 ( .A1(n12324), .A2(n12637), .ZN(n12453) );
  XOR2_X1 U12253 ( .A(n12462), .B(n12311), .Z(n12622) );
  OAI21_X1 U12254 ( .B1(n9809), .B2(n9820), .A(n12608), .ZN(n9771) );
  NAND2_X1 U12255 ( .A1(n9771), .A2(n10819), .ZN(n9773) );
  OAI21_X1 U12256 ( .B1(n9820), .B2(n12340), .A(n9809), .ZN(n9772) );
  NAND2_X1 U12257 ( .A1(n9773), .A2(n9772), .ZN(n10476) );
  INV_X1 U12258 ( .A(n12608), .ZN(n10513) );
  NAND2_X1 U12259 ( .A1(n10820), .A2(n10513), .ZN(n9822) );
  INV_X1 U12260 ( .A(n9822), .ZN(n12477) );
  AND2_X1 U12261 ( .A1(n15368), .A2(n12477), .ZN(n9774) );
  NAND2_X1 U12262 ( .A1(n10476), .A2(n9774), .ZN(n9775) );
  NAND2_X1 U12263 ( .A1(n6626), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9779) );
  MUX2_X1 U12264 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9779), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n9780) );
  NAND2_X1 U12265 ( .A1(n9781), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9782) );
  MUX2_X1 U12266 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9782), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9783) );
  INV_X1 U12267 ( .A(n9784), .ZN(n9785) );
  NAND2_X1 U12268 ( .A1(n9785), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9786) );
  MUX2_X1 U12269 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9786), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n9787) );
  NAND2_X1 U12270 ( .A1(n9787), .A2(n9781), .ZN(n11378) );
  INV_X1 U12271 ( .A(n11378), .ZN(n9788) );
  NAND2_X1 U12272 ( .A1(n9790), .A2(n9788), .ZN(n9789) );
  XNOR2_X1 U12273 ( .A(n11378), .B(P3_B_REG_SCAN_IN), .ZN(n9791) );
  INV_X1 U12274 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9793) );
  NAND2_X1 U12275 ( .A1(n10203), .A2(n9793), .ZN(n9795) );
  NAND2_X1 U12276 ( .A1(n11610), .A2(n11504), .ZN(n9794) );
  INV_X1 U12277 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9796) );
  NAND2_X1 U12278 ( .A1(n10647), .A2(n9797), .ZN(n9827) );
  NOR2_X1 U12279 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .ZN(
        n9801) );
  NOR4_X1 U12280 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_30__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n9800) );
  NOR4_X1 U12281 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n9799) );
  NOR4_X1 U12282 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n9798) );
  NAND4_X1 U12283 ( .A1(n9801), .A2(n9800), .A3(n9799), .A4(n9798), .ZN(n9807)
         );
  NOR4_X1 U12284 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n9805) );
  NOR4_X1 U12285 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n9804) );
  NOR4_X1 U12286 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9803) );
  NOR4_X1 U12287 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9802) );
  NAND4_X1 U12288 ( .A1(n9805), .A2(n9804), .A3(n9803), .A4(n9802), .ZN(n9806)
         );
  NAND2_X1 U12289 ( .A1(n9827), .A2(n9825), .ZN(n9808) );
  OAI22_X1 U12290 ( .A1(n15368), .A2(n9820), .B1(n12608), .B2(n9809), .ZN(
        n9810) );
  NAND2_X1 U12291 ( .A1(n9810), .A2(n9822), .ZN(n9811) );
  NAND2_X1 U12292 ( .A1(n9811), .A2(n12448), .ZN(n9812) );
  NAND2_X1 U12293 ( .A1(n9812), .A2(n10647), .ZN(n9815) );
  NAND2_X1 U12294 ( .A1(n12448), .A2(n9813), .ZN(n10649) );
  NAND2_X1 U12295 ( .A1(n10480), .A2(n10649), .ZN(n10648) );
  NAND2_X1 U12296 ( .A1(n10648), .A2(n12950), .ZN(n9814) );
  MUX2_X1 U12297 ( .A(n9816), .B(n9830), .S(n15395), .Z(n9819) );
  NAND2_X1 U12298 ( .A1(n9817), .A2(n10517), .ZN(n9818) );
  NAND2_X1 U12299 ( .A1(n9819), .A2(n9818), .ZN(P3_U3488) );
  INV_X1 U12300 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9831) );
  OR2_X1 U12301 ( .A1(n9821), .A2(n10817), .ZN(n10478) );
  OR2_X1 U12302 ( .A1(n12448), .A2(n9822), .ZN(n10514) );
  OAI21_X1 U12303 ( .B1(n10654), .B2(n10478), .A(n12508), .ZN(n9824) );
  AND2_X1 U12304 ( .A1(n9823), .A2(n9825), .ZN(n10492) );
  NAND2_X1 U12305 ( .A1(n9824), .A2(n10492), .ZN(n9829) );
  INV_X1 U12306 ( .A(n10654), .ZN(n10474) );
  INV_X1 U12307 ( .A(n9825), .ZN(n9826) );
  NAND3_X1 U12308 ( .A1(n10474), .A2(n10488), .A3(n10476), .ZN(n9828) );
  MUX2_X1 U12309 ( .A(n9831), .B(n9830), .S(n15379), .Z(n9834) );
  NAND2_X1 U12310 ( .A1(n9834), .A2(n9833), .ZN(P3_U3456) );
  NAND3_X1 U12311 ( .A1(n12643), .A2(n12455), .A3(n12450), .ZN(n9835) );
  NAND2_X1 U12312 ( .A1(n9836), .A2(n9835), .ZN(n12630) );
  INV_X1 U12313 ( .A(n9837), .ZN(n9840) );
  AOI21_X1 U12314 ( .B1(n12635), .B2(n9838), .A(n12455), .ZN(n9839) );
  NOR3_X1 U12315 ( .A1(n9840), .A2(n9839), .A3(n15299), .ZN(n9842) );
  OAI22_X1 U12316 ( .A1(n12654), .A2(n15292), .B1(n12205), .B2(n15294), .ZN(
        n9841) );
  AOI21_X1 U12317 ( .B1(n15366), .B2(n12630), .A(n12625), .ZN(n9847) );
  OR2_X1 U12318 ( .A1(n9847), .A2(n15392), .ZN(n9846) );
  INV_X1 U12319 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n9843) );
  INV_X1 U12320 ( .A(n9844), .ZN(n9845) );
  NAND2_X1 U12321 ( .A1(n9846), .A2(n9845), .ZN(P3_U3487) );
  OR2_X1 U12322 ( .A1(n9847), .A2(n15378), .ZN(n9850) );
  INV_X1 U12323 ( .A(n9848), .ZN(n9849) );
  NAND2_X1 U12324 ( .A1(n9850), .A2(n9849), .ZN(P3_U3455) );
  INV_X1 U12325 ( .A(n10170), .ZN(n9854) );
  INV_X4 U12326 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U12327 ( .A1(n10407), .A2(n14465), .ZN(n9855) );
  NAND2_X1 U12328 ( .A1(n9855), .A2(n9156), .ZN(n10409) );
  INV_X1 U12329 ( .A(n10409), .ZN(n9858) );
  NAND2_X1 U12330 ( .A1(n9858), .A2(n7536), .ZN(n10456) );
  NAND2_X1 U12331 ( .A1(n13086), .A2(n9942), .ZN(n9862) );
  INV_X1 U12332 ( .A(n9860), .ZN(n9861) );
  NAND2_X1 U12333 ( .A1(n9862), .A2(n9861), .ZN(n9863) );
  INV_X1 U12334 ( .A(n6579), .ZN(n9864) );
  INV_X1 U12335 ( .A(n9867), .ZN(n9865) );
  NAND2_X1 U12336 ( .A1(n9866), .A2(n9865), .ZN(n9870) );
  NAND2_X1 U12337 ( .A1(n9868), .A2(n9867), .ZN(n9869) );
  NAND2_X1 U12338 ( .A1(n13084), .A2(n9942), .ZN(n9872) );
  XNOR2_X1 U12339 ( .A(n9871), .B(n6580), .ZN(n9873) );
  XNOR2_X1 U12340 ( .A(n9872), .B(n9873), .ZN(n10520) );
  INV_X1 U12341 ( .A(n10520), .ZN(n9876) );
  INV_X1 U12342 ( .A(n9872), .ZN(n9875) );
  INV_X1 U12343 ( .A(n9873), .ZN(n9874) );
  XNOR2_X1 U12344 ( .A(n13022), .B(n6580), .ZN(n9878) );
  NAND2_X1 U12345 ( .A1(n9878), .A2(n9879), .ZN(n9883) );
  INV_X1 U12346 ( .A(n9878), .ZN(n9881) );
  INV_X1 U12347 ( .A(n9879), .ZN(n9880) );
  NAND2_X1 U12348 ( .A1(n9881), .A2(n9880), .ZN(n9882) );
  AND2_X1 U12349 ( .A1(n9883), .A2(n9882), .ZN(n13019) );
  NAND2_X1 U12350 ( .A1(n13020), .A2(n13019), .ZN(n13018) );
  XNOR2_X1 U12351 ( .A(n11242), .B(n6580), .ZN(n9884) );
  NAND2_X1 U12352 ( .A1(n13082), .A2(n9935), .ZN(n9885) );
  NAND2_X1 U12353 ( .A1(n9884), .A2(n9885), .ZN(n9889) );
  INV_X1 U12354 ( .A(n9884), .ZN(n9887) );
  INV_X1 U12355 ( .A(n9885), .ZN(n9886) );
  NAND2_X1 U12356 ( .A1(n9887), .A2(n9886), .ZN(n9888) );
  AND2_X1 U12357 ( .A1(n9889), .A2(n9888), .ZN(n10527) );
  NAND2_X1 U12358 ( .A1(n13081), .A2(n9935), .ZN(n9892) );
  XNOR2_X1 U12359 ( .A(n9891), .B(n9892), .ZN(n10566) );
  INV_X1 U12360 ( .A(n10566), .ZN(n9890) );
  INV_X1 U12361 ( .A(n9891), .ZN(n9894) );
  INV_X1 U12362 ( .A(n9892), .ZN(n9893) );
  NAND2_X1 U12363 ( .A1(n9894), .A2(n9893), .ZN(n9895) );
  XNOR2_X1 U12364 ( .A(n15057), .B(n12116), .ZN(n9898) );
  NAND2_X1 U12365 ( .A1(n13080), .A2(n9935), .ZN(n9896) );
  XNOR2_X1 U12366 ( .A(n9898), .B(n9896), .ZN(n10808) );
  INV_X1 U12367 ( .A(n9896), .ZN(n9897) );
  AND2_X1 U12368 ( .A1(n9898), .A2(n9897), .ZN(n9899) );
  XNOR2_X1 U12369 ( .A(n11052), .B(n6579), .ZN(n9900) );
  NAND2_X1 U12370 ( .A1(n13079), .A2(n9935), .ZN(n9901) );
  NAND2_X1 U12371 ( .A1(n9900), .A2(n9901), .ZN(n9905) );
  INV_X1 U12372 ( .A(n9900), .ZN(n9903) );
  INV_X1 U12373 ( .A(n9901), .ZN(n9902) );
  NAND2_X1 U12374 ( .A1(n9903), .A2(n9902), .ZN(n9904) );
  AND2_X1 U12375 ( .A1(n9905), .A2(n9904), .ZN(n10969) );
  NAND2_X1 U12376 ( .A1(n10970), .A2(n10969), .ZN(n10968) );
  XNOR2_X1 U12377 ( .A(n11339), .B(n6580), .ZN(n9906) );
  NAND2_X1 U12378 ( .A1(n13078), .A2(n9935), .ZN(n9907) );
  NAND2_X1 U12379 ( .A1(n9906), .A2(n9907), .ZN(n9911) );
  INV_X1 U12380 ( .A(n9906), .ZN(n9909) );
  INV_X1 U12381 ( .A(n9907), .ZN(n9908) );
  NAND2_X1 U12382 ( .A1(n9909), .A2(n9908), .ZN(n9910) );
  AND2_X1 U12383 ( .A1(n9911), .A2(n9910), .ZN(n11065) );
  XNOR2_X1 U12384 ( .A(n11356), .B(n6579), .ZN(n9912) );
  NAND2_X1 U12385 ( .A1(n13077), .A2(n9935), .ZN(n9913) );
  XNOR2_X1 U12386 ( .A(n9912), .B(n9913), .ZN(n11150) );
  INV_X1 U12387 ( .A(n9912), .ZN(n9915) );
  INV_X1 U12388 ( .A(n9913), .ZN(n9914) );
  NAND2_X1 U12389 ( .A1(n9915), .A2(n9914), .ZN(n9916) );
  XNOR2_X1 U12390 ( .A(n11551), .B(n6579), .ZN(n9917) );
  NAND2_X1 U12391 ( .A1(n13076), .A2(n9935), .ZN(n9918) );
  NAND2_X1 U12392 ( .A1(n9917), .A2(n9918), .ZN(n9923) );
  INV_X1 U12393 ( .A(n9917), .ZN(n9920) );
  INV_X1 U12394 ( .A(n9918), .ZN(n9919) );
  NAND2_X1 U12395 ( .A1(n9920), .A2(n9919), .ZN(n9921) );
  NAND2_X1 U12396 ( .A1(n9923), .A2(n9921), .ZN(n11363) );
  XNOR2_X1 U12397 ( .A(n14482), .B(n6580), .ZN(n9924) );
  NAND2_X1 U12398 ( .A1(n13075), .A2(n9935), .ZN(n9925) );
  NAND2_X1 U12399 ( .A1(n9924), .A2(n9925), .ZN(n9929) );
  INV_X1 U12400 ( .A(n9924), .ZN(n9927) );
  INV_X1 U12401 ( .A(n9925), .ZN(n9926) );
  NAND2_X1 U12402 ( .A1(n9927), .A2(n9926), .ZN(n9928) );
  AND2_X1 U12403 ( .A1(n9929), .A2(n9928), .ZN(n11381) );
  XNOR2_X1 U12404 ( .A(n11563), .B(n6579), .ZN(n9930) );
  NAND2_X1 U12405 ( .A1(n13074), .A2(n9935), .ZN(n9931) );
  XNOR2_X1 U12406 ( .A(n9930), .B(n9931), .ZN(n11436) );
  INV_X1 U12407 ( .A(n9930), .ZN(n9933) );
  INV_X1 U12408 ( .A(n9931), .ZN(n9932) );
  NAND2_X1 U12409 ( .A1(n9933), .A2(n9932), .ZN(n9934) );
  XNOR2_X1 U12410 ( .A(n14461), .B(n6580), .ZN(n9936) );
  NAND2_X1 U12411 ( .A1(n13073), .A2(n9935), .ZN(n9937) );
  NAND2_X1 U12412 ( .A1(n9936), .A2(n9937), .ZN(n9941) );
  INV_X1 U12413 ( .A(n9936), .ZN(n9939) );
  INV_X1 U12414 ( .A(n9937), .ZN(n9938) );
  NAND2_X1 U12415 ( .A1(n9939), .A2(n9938), .ZN(n9940) );
  AND2_X1 U12416 ( .A1(n9941), .A2(n9940), .ZN(n14447) );
  XOR2_X1 U12417 ( .A(n12116), .B(n11841), .Z(n9944) );
  NAND2_X1 U12418 ( .A1(n13072), .A2(n9935), .ZN(n11699) );
  XNOR2_X1 U12419 ( .A(n13445), .B(n12116), .ZN(n9946) );
  OR2_X1 U12420 ( .A1(n11847), .A2(n14465), .ZN(n9945) );
  NAND2_X1 U12421 ( .A1(n9946), .A2(n9945), .ZN(n9947) );
  OAI21_X1 U12422 ( .B1(n9946), .B2(n9945), .A(n9947), .ZN(n11824) );
  INV_X1 U12423 ( .A(n9947), .ZN(n9948) );
  XNOR2_X1 U12424 ( .A(n13437), .B(n6580), .ZN(n9950) );
  NAND2_X1 U12425 ( .A1(n13334), .A2(n9935), .ZN(n9949) );
  NAND2_X1 U12426 ( .A1(n9950), .A2(n9949), .ZN(n9951) );
  OAI21_X1 U12427 ( .B1(n9950), .B2(n9949), .A(n9951), .ZN(n11845) );
  INV_X1 U12428 ( .A(n9951), .ZN(n9952) );
  XNOR2_X1 U12429 ( .A(n13429), .B(n12116), .ZN(n9955) );
  NAND2_X1 U12430 ( .A1(n13070), .A2(n9935), .ZN(n9953) );
  XNOR2_X1 U12431 ( .A(n9955), .B(n9953), .ZN(n13041) );
  INV_X1 U12432 ( .A(n9953), .ZN(n9954) );
  AND2_X1 U12433 ( .A1(n13337), .A2(n9935), .ZN(n9957) );
  XNOR2_X1 U12434 ( .A(n13426), .B(n12116), .ZN(n9956) );
  NOR2_X1 U12435 ( .A1(n9956), .A2(n9957), .ZN(n9958) );
  AOI21_X1 U12436 ( .B1(n9957), .B2(n9956), .A(n9958), .ZN(n12984) );
  INV_X1 U12437 ( .A(n9958), .ZN(n9959) );
  XNOR2_X1 U12438 ( .A(n13420), .B(n12116), .ZN(n9961) );
  AND2_X1 U12439 ( .A1(n13069), .A2(n9935), .ZN(n9960) );
  NOR2_X1 U12440 ( .A1(n9961), .A2(n9960), .ZN(n13031) );
  NAND2_X1 U12441 ( .A1(n9961), .A2(n9960), .ZN(n13032) );
  XNOR2_X1 U12442 ( .A(n13295), .B(n12116), .ZN(n9962) );
  NAND2_X1 U12443 ( .A1(n13272), .A2(n9935), .ZN(n9963) );
  XNOR2_X1 U12444 ( .A(n9962), .B(n9963), .ZN(n12993) );
  NAND2_X1 U12445 ( .A1(n9962), .A2(n9964), .ZN(n9965) );
  XNOR2_X1 U12446 ( .A(n13409), .B(n12116), .ZN(n12090) );
  NAND2_X1 U12447 ( .A1(n13068), .A2(n9935), .ZN(n9968) );
  AND2_X1 U12448 ( .A1(n9987), .A2(n15074), .ZN(n9980) );
  INV_X1 U12449 ( .A(n9980), .ZN(n9970) );
  AOI211_X1 U12450 ( .C1(n9967), .C2(n9968), .A(n13059), .B(n12093), .ZN(n9984) );
  INV_X1 U12451 ( .A(n13409), .ZN(n13279) );
  INV_X1 U12452 ( .A(n11005), .ZN(n9969) );
  OR2_X1 U12453 ( .A1(n9969), .A2(n11262), .ZN(n9999) );
  OR2_X1 U12454 ( .A1(n9970), .A2(n9999), .ZN(n9972) );
  INV_X1 U12455 ( .A(n9973), .ZN(n9971) );
  NOR2_X1 U12456 ( .A1(n13279), .A2(n13017), .ZN(n9983) );
  OAI21_X1 U12457 ( .B1(n10383), .B2(n9974), .A(n9973), .ZN(n9977) );
  AND2_X1 U12458 ( .A1(n9975), .A2(n10381), .ZN(n9976) );
  NAND2_X1 U12459 ( .A1(n9977), .A2(n9976), .ZN(n10406) );
  OAI22_X1 U12460 ( .A1(n14453), .A2(n13276), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9978), .ZN(n9982) );
  NAND2_X1 U12461 ( .A1(n14450), .A2(n13336), .ZN(n13044) );
  NAND2_X1 U12462 ( .A1(n14450), .A2(n13335), .ZN(n13045) );
  OAI22_X1 U12463 ( .A1(n12094), .A2(n13044), .B1(n13045), .B2(n13036), .ZN(
        n9981) );
  INV_X1 U12464 ( .A(n9985), .ZN(n10481) );
  NAND2_X1 U12465 ( .A1(n9987), .A2(n9986), .ZN(n9988) );
  OAI211_X1 U12466 ( .C1(n11012), .C2(n10595), .A(n14465), .B(n11083), .ZN(
        n10466) );
  OR3_X1 U12467 ( .A1(n13358), .A2(n11192), .A3(n9989), .ZN(n13348) );
  INV_X1 U12468 ( .A(n9990), .ZN(n9991) );
  AOI21_X1 U12469 ( .B1(n9992), .B2(n9994), .A(n9991), .ZN(n10465) );
  OAI22_X1 U12470 ( .A1(n15061), .A2(n10466), .B1(n13348), .B2(n10465), .ZN(
        n10002) );
  OAI21_X1 U12471 ( .B1(n9995), .B2(n9994), .A(n9993), .ZN(n9997) );
  OAI22_X1 U12472 ( .A1(n10460), .A2(n14443), .B1(n8155), .B2(n14441), .ZN(
        n9996) );
  AOI21_X1 U12473 ( .B1(n9997), .B2(n14456), .A(n9996), .ZN(n9998) );
  OAI21_X1 U12474 ( .B1(n10465), .B2(n8198), .A(n9998), .ZN(n10467) );
  MUX2_X1 U12475 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10467), .S(n15055), .Z(
        n10001) );
  OAI22_X1 U12476 ( .A1(n13360), .A2(n10595), .B1(n10458), .B2(n15052), .ZN(
        n10000) );
  OR3_X1 U12477 ( .A1(n10002), .A2(n10001), .A3(n10000), .ZN(P2_U3264) );
  INV_X2 U12478 ( .A(n13769), .ZN(n13776) );
  INV_X2 U12479 ( .A(n6726), .ZN(n11134) );
  OAI222_X1 U12480 ( .A1(n13776), .A2(n10233), .B1(n11134), .B2(n10009), .C1(
        P2_U3088), .C2(n14868), .ZN(P2_U3326) );
  OAI222_X1 U12481 ( .A1(n13776), .A2(n10003), .B1(n11134), .B2(n10007), .C1(
        P2_U3088), .C2(n14879), .ZN(P2_U3325) );
  INV_X1 U12482 ( .A(n10004), .ZN(n10011) );
  OAI222_X1 U12483 ( .A1(n13776), .A2(n7621), .B1(n11134), .B2(n10011), .C1(
        P2_U3088), .C2(n13090), .ZN(P2_U3324) );
  INV_X1 U12484 ( .A(n14649), .ZN(n10082) );
  INV_X2 U12485 ( .A(n14292), .ZN(n14304) );
  OAI222_X1 U12486 ( .A1(n10082), .A2(P1_U3086), .B1(n14304), .B2(n10007), 
        .C1(n10006), .C2(n14298), .ZN(P1_U3353) );
  INV_X1 U12487 ( .A(n13904), .ZN(n10010) );
  OAI222_X1 U12488 ( .A1(n10010), .A2(P1_U3086), .B1(n14304), .B2(n10009), 
        .C1(n10008), .C2(n14298), .ZN(P1_U3354) );
  INV_X1 U12489 ( .A(n13915), .ZN(n10012) );
  OAI222_X1 U12490 ( .A1(n10012), .A2(P1_U3086), .B1(n14304), .B2(n10011), 
        .C1(n7054), .C2(n14298), .ZN(P1_U3352) );
  INV_X1 U12491 ( .A(n10013), .ZN(n10016) );
  OAI222_X1 U12492 ( .A1(n13776), .A2(n10014), .B1(n11134), .B2(n10016), .C1(
        P2_U3088), .C2(n10345), .ZN(P2_U3323) );
  INV_X1 U12493 ( .A(n10098), .ZN(n14672) );
  OAI222_X1 U12494 ( .A1(n14672), .A2(P1_U3086), .B1(n14304), .B2(n10016), 
        .C1(n10015), .C2(n14298), .ZN(P1_U3351) );
  INV_X2 U12495 ( .A(n14325), .ZN(n12961) );
  INV_X2 U12496 ( .A(n6727), .ZN(n12962) );
  INV_X1 U12497 ( .A(SI_6_), .ZN(n10018) );
  INV_X1 U12498 ( .A(n10674), .ZN(n10017) );
  OAI222_X1 U12499 ( .A1(n12961), .A2(n10019), .B1(n12962), .B2(n10018), .C1(
        P3_U3151), .C2(n10017), .ZN(P3_U3289) );
  OAI222_X1 U12500 ( .A1(n12571), .A2(P3_U3151), .B1(n12961), .B2(n10021), 
        .C1(n10020), .C2(n12962), .ZN(P3_U3285) );
  OAI222_X1 U12501 ( .A1(P3_U3151), .A2(n10745), .B1(n12961), .B2(n10023), 
        .C1(n10022), .C2(n12962), .ZN(P3_U3290) );
  INV_X1 U12502 ( .A(n10024), .ZN(n10026) );
  INV_X1 U12503 ( .A(SI_8_), .ZN(n10025) );
  OAI222_X1 U12504 ( .A1(n12564), .A2(P3_U3151), .B1(n12961), .B2(n10026), 
        .C1(n10025), .C2(n12962), .ZN(P3_U3287) );
  OAI222_X1 U12505 ( .A1(P3_U3151), .A2(n10546), .B1(n12961), .B2(n10030), 
        .C1(n10029), .C2(n12962), .ZN(P3_U3292) );
  INV_X1 U12506 ( .A(n10435), .ZN(n10646) );
  INV_X1 U12507 ( .A(n10031), .ZN(n10033) );
  OAI222_X1 U12508 ( .A1(n10646), .A2(P3_U3151), .B1(n12961), .B2(n10033), 
        .C1(n10032), .C2(n12962), .ZN(P3_U3294) );
  OAI222_X1 U12509 ( .A1(P3_U3151), .A2(n10711), .B1(n12962), .B2(n10035), 
        .C1(n12961), .C2(n10034), .ZN(P3_U3288) );
  OAI222_X1 U12510 ( .A1(P3_U3151), .A2(n15124), .B1(n12962), .B2(n10037), 
        .C1(n12961), .C2(n10036), .ZN(P3_U3286) );
  INV_X1 U12511 ( .A(n10038), .ZN(n10042) );
  INV_X1 U12512 ( .A(n13104), .ZN(n10039) );
  OAI222_X1 U12513 ( .A1(n13776), .A2(n10040), .B1(n11134), .B2(n10042), .C1(
        P2_U3088), .C2(n10039), .ZN(P2_U3322) );
  INV_X1 U12514 ( .A(n10100), .ZN(n10113) );
  OAI222_X1 U12515 ( .A1(n10113), .A2(P1_U3086), .B1(n14304), .B2(n10042), 
        .C1(n10041), .C2(n14298), .ZN(P1_U3350) );
  OAI222_X1 U12516 ( .A1(P3_U3151), .A2(n15163), .B1(n12962), .B2(n10044), 
        .C1(n12961), .C2(n10043), .ZN(P3_U3284) );
  INV_X1 U12517 ( .A(n10045), .ZN(n10049) );
  INV_X1 U12518 ( .A(n14907), .ZN(n10046) );
  OAI222_X1 U12519 ( .A1(n13776), .A2(n10047), .B1(n11134), .B2(n10049), .C1(
        P2_U3088), .C2(n10046), .ZN(P2_U3321) );
  INV_X1 U12520 ( .A(n10102), .ZN(n13921) );
  OAI222_X1 U12521 ( .A1(n13921), .A2(P1_U3086), .B1(n14304), .B2(n10049), 
        .C1(n10048), .C2(n14298), .ZN(P1_U3349) );
  INV_X1 U12522 ( .A(n14301), .ZN(n10050) );
  AND2_X1 U12523 ( .A1(n10051), .A2(n10050), .ZN(n10053) );
  NAND3_X1 U12524 ( .A1(n14305), .A2(P1_B_REG_SCAN_IN), .A3(n11695), .ZN(
        n10052) );
  INV_X1 U12525 ( .A(n10273), .ZN(n10287) );
  NAND2_X1 U12526 ( .A1(n10287), .A2(n10302), .ZN(n14760) );
  INV_X1 U12527 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10272) );
  AND2_X1 U12528 ( .A1(n14305), .A2(n14301), .ZN(n10271) );
  AOI22_X1 U12529 ( .A1(n14760), .A2(n10272), .B1(n10054), .B2(n10271), .ZN(
        P1_U3446) );
  OAI222_X1 U12530 ( .A1(P3_U3151), .A2(n15181), .B1(n12962), .B2(n10056), 
        .C1(n12961), .C2(n10055), .ZN(P3_U3283) );
  INV_X1 U12531 ( .A(n10057), .ZN(n10060) );
  INV_X1 U12532 ( .A(n10131), .ZN(n10058) );
  OAI222_X1 U12533 ( .A1(n14298), .A2(n10059), .B1(n14304), .B2(n10060), .C1(
        n10058), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U12534 ( .A(n10349), .ZN(n14923) );
  OAI222_X1 U12535 ( .A1(n13776), .A2(n10061), .B1(n11134), .B2(n10060), .C1(
        P2_U3088), .C2(n14923), .ZN(P2_U3320) );
  NAND2_X1 U12536 ( .A1(n10288), .A2(n11615), .ZN(n10067) );
  NAND2_X1 U12537 ( .A1(n10296), .A2(n10062), .ZN(n10063) );
  NAND2_X1 U12538 ( .A1(n10064), .A2(n10063), .ZN(n10065) );
  AND2_X1 U12539 ( .A1(n10067), .A2(n10065), .ZN(n14675) );
  INV_X1 U12540 ( .A(n10065), .ZN(n10066) );
  NAND2_X1 U12541 ( .A1(n10067), .A2(n10066), .ZN(n10086) );
  INV_X1 U12542 ( .A(n10086), .ZN(n10104) );
  NOR2_X1 U12543 ( .A1(n14650), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10068) );
  NOR2_X1 U12544 ( .A1(n11878), .A2(n10068), .ZN(n14657) );
  OAI21_X1 U12545 ( .B1(n11938), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14657), .ZN(
        n10069) );
  XNOR2_X1 U12546 ( .A(n10069), .B(P1_IR_REG_0__SCAN_IN), .ZN(n10070) );
  AOI22_X1 U12547 ( .A1(n10104), .A2(n10070), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10071) );
  OAI21_X1 U12548 ( .B1(n14695), .B2(n6842), .A(n10071), .ZN(P1_U3243) );
  NAND2_X1 U12549 ( .A1(n11695), .A2(n14301), .ZN(n10274) );
  OAI22_X1 U12550 ( .A1(n14759), .A2(P1_D_REG_0__SCAN_IN), .B1(n10072), .B2(
        n10274), .ZN(n10073) );
  INV_X1 U12551 ( .A(n10073), .ZN(P1_U3445) );
  INV_X1 U12552 ( .A(n10074), .ZN(n10076) );
  OAI222_X1 U12553 ( .A1(n10145), .A2(P1_U3086), .B1(n14304), .B2(n10076), 
        .C1(n10075), .C2(n14298), .ZN(P1_U3347) );
  INV_X1 U12554 ( .A(n10351), .ZN(n14936) );
  OAI222_X1 U12555 ( .A1(n13776), .A2(n10235), .B1(n11134), .B2(n10076), .C1(
        P2_U3088), .C2(n14936), .ZN(P2_U3319) );
  OAI222_X1 U12556 ( .A1(P3_U3151), .A2(n15199), .B1(n12962), .B2(n13723), 
        .C1(n12961), .C2(n10077), .ZN(P3_U3282) );
  INV_X1 U12557 ( .A(n10078), .ZN(n10079) );
  OAI222_X1 U12558 ( .A1(n13776), .A2(n10237), .B1(n11134), .B2(n10079), .C1(
        P2_U3088), .C2(n10354), .ZN(P2_U3318) );
  INV_X1 U12559 ( .A(n10189), .ZN(n10130) );
  OAI222_X1 U12560 ( .A1(n10130), .A2(P1_U3086), .B1(n14304), .B2(n10079), 
        .C1(n13553), .C2(n14298), .ZN(P1_U3346) );
  NOR2_X1 U12561 ( .A1(n14675), .A2(n14655), .ZN(P1_U3085) );
  INV_X1 U12562 ( .A(n14673), .ZN(n14687) );
  NAND2_X1 U12563 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11404) );
  OAI21_X1 U12564 ( .B1(n14695), .B2(n8880), .A(n11404), .ZN(n10092) );
  INV_X1 U12565 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10080) );
  MUX2_X1 U12566 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n10080), .S(n13904), .Z(
        n13901) );
  NAND3_X1 U12567 ( .A1(n13901), .A2(P1_REG2_REG_0__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n14637) );
  NAND2_X1 U12568 ( .A1(n13904), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n14636) );
  INV_X1 U12569 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10081) );
  MUX2_X1 U12570 ( .A(n10081), .B(P1_REG2_REG_2__SCAN_IN), .S(n14649), .Z(
        n14638) );
  AOI21_X1 U12571 ( .B1(n14637), .B2(n14636), .A(n14638), .ZN(n14640) );
  NOR2_X1 U12572 ( .A1(n10082), .A2(n10081), .ZN(n13912) );
  MUX2_X1 U12573 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n14740), .S(n13915), .Z(
        n13913) );
  OAI21_X1 U12574 ( .B1(n14640), .B2(n13912), .A(n13913), .ZN(n14666) );
  NAND2_X1 U12575 ( .A1(n13915), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14665) );
  MUX2_X1 U12576 ( .A(n10803), .B(P1_REG2_REG_4__SCAN_IN), .S(n10098), .Z(
        n14664) );
  AOI21_X1 U12577 ( .B1(n14666), .B2(n14665), .A(n14664), .ZN(n14663) );
  NOR2_X1 U12578 ( .A1(n14672), .A2(n10803), .ZN(n10117) );
  MUX2_X1 U12579 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10083), .S(n10100), .Z(
        n10116) );
  OAI21_X1 U12580 ( .B1(n14663), .B2(n10117), .A(n10116), .ZN(n13930) );
  NAND2_X1 U12581 ( .A1(n10100), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n13929) );
  MUX2_X1 U12582 ( .A(n11125), .B(P1_REG2_REG_6__SCAN_IN), .S(n10102), .Z(
        n13928) );
  AOI21_X1 U12583 ( .B1(n13930), .B2(n13929), .A(n13928), .ZN(n13927) );
  NOR2_X1 U12584 ( .A1(n13921), .A2(n11125), .ZN(n10088) );
  MUX2_X1 U12585 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10084), .S(n10131), .Z(
        n10087) );
  OAI21_X1 U12586 ( .B1(n13927), .B2(n10088), .A(n10087), .ZN(n10151) );
  INV_X1 U12587 ( .A(n10151), .ZN(n10090) );
  NAND2_X1 U12588 ( .A1(n14653), .A2(n11938), .ZN(n10085) );
  NOR3_X1 U12589 ( .A1(n13927), .A2(n10088), .A3(n10087), .ZN(n10089) );
  NOR3_X1 U12590 ( .A1(n10090), .A2(n14690), .A3(n10089), .ZN(n10091) );
  AOI211_X1 U12591 ( .C1(n14687), .C2(n10131), .A(n10092), .B(n10091), .ZN(
        n10108) );
  MUX2_X1 U12592 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n8421), .S(n10131), .Z(
        n10106) );
  NAND2_X1 U12593 ( .A1(n13915), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10096) );
  OR2_X1 U12594 ( .A1(n13915), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10093) );
  AND2_X1 U12595 ( .A1(n10096), .A2(n10093), .ZN(n13911) );
  MUX2_X1 U12596 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n8329), .S(n14649), .Z(
        n14641) );
  MUX2_X1 U12597 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n8300), .S(n13904), .Z(
        n13903) );
  AND2_X1 U12598 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13902) );
  NAND2_X1 U12599 ( .A1(n13903), .A2(n13902), .ZN(n14642) );
  NAND2_X1 U12600 ( .A1(n13904), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n14643) );
  NAND2_X1 U12601 ( .A1(n14642), .A2(n14643), .ZN(n10094) );
  NAND2_X1 U12602 ( .A1(n14641), .A2(n10094), .ZN(n14646) );
  NAND2_X1 U12603 ( .A1(n14649), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10095) );
  NAND2_X1 U12604 ( .A1(n14646), .A2(n10095), .ZN(n13910) );
  NAND2_X1 U12605 ( .A1(n13911), .A2(n13910), .ZN(n13909) );
  NAND2_X1 U12606 ( .A1(n13909), .A2(n10096), .ZN(n14661) );
  INV_X1 U12607 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10097) );
  XNOR2_X1 U12608 ( .A(n10098), .B(n10097), .ZN(n14662) );
  NAND2_X1 U12609 ( .A1(n14661), .A2(n14662), .ZN(n14660) );
  NAND2_X1 U12610 ( .A1(n10098), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10099) );
  NAND2_X1 U12611 ( .A1(n14660), .A2(n10099), .ZN(n10111) );
  MUX2_X1 U12612 ( .A(n8384), .B(P1_REG1_REG_5__SCAN_IN), .S(n10100), .Z(
        n10112) );
  OR2_X1 U12613 ( .A1(n10111), .A2(n10112), .ZN(n10109) );
  OR2_X1 U12614 ( .A1(n10100), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10101) );
  AND2_X1 U12615 ( .A1(n10109), .A2(n10101), .ZN(n13925) );
  MUX2_X1 U12616 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n8400), .S(n10102), .Z(
        n13926) );
  NAND2_X1 U12617 ( .A1(n13925), .A2(n13926), .ZN(n13924) );
  NAND2_X1 U12618 ( .A1(n10102), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10103) );
  NAND2_X1 U12619 ( .A1(n13924), .A2(n10103), .ZN(n10105) );
  NAND2_X1 U12620 ( .A1(n10105), .A2(n10106), .ZN(n10124) );
  OAI211_X1 U12621 ( .C1(n10106), .C2(n10105), .A(n14684), .B(n10124), .ZN(
        n10107) );
  NAND2_X1 U12622 ( .A1(n10108), .A2(n10107), .ZN(P1_U3250) );
  INV_X1 U12623 ( .A(n10109), .ZN(n10110) );
  AOI21_X1 U12624 ( .B1(n10112), .B2(n10111), .A(n10110), .ZN(n10121) );
  INV_X1 U12625 ( .A(n14684), .ZN(n13940) );
  NAND2_X1 U12626 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n11186) );
  INV_X1 U12627 ( .A(n11186), .ZN(n10115) );
  NOR2_X1 U12628 ( .A1(n14673), .A2(n10113), .ZN(n10114) );
  AOI211_X1 U12629 ( .C1(n14675), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n10115), .B(
        n10114), .ZN(n10120) );
  INV_X1 U12630 ( .A(n14690), .ZN(n14669) );
  OR3_X1 U12631 ( .A1(n14663), .A2(n10117), .A3(n10116), .ZN(n10118) );
  NAND3_X1 U12632 ( .A1(n14669), .A2(n13930), .A3(n10118), .ZN(n10119) );
  OAI211_X1 U12633 ( .C1(n10121), .C2(n13940), .A(n10120), .B(n10119), .ZN(
        P1_U3248) );
  MUX2_X1 U12634 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10122), .S(n10189), .Z(
        n10128) );
  NAND2_X1 U12635 ( .A1(n10131), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10123) );
  NAND2_X1 U12636 ( .A1(n10124), .A2(n10123), .ZN(n10143) );
  MUX2_X1 U12637 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10125), .S(n10145), .Z(
        n10144) );
  OR2_X1 U12638 ( .A1(n10143), .A2(n10144), .ZN(n10141) );
  NAND2_X1 U12639 ( .A1(n10145), .A2(n10125), .ZN(n10126) );
  NAND2_X1 U12640 ( .A1(n10141), .A2(n10126), .ZN(n10127) );
  NAND2_X1 U12641 ( .A1(n10127), .A2(n10128), .ZN(n10191) );
  OAI21_X1 U12642 ( .B1(n10128), .B2(n10127), .A(n10191), .ZN(n10139) );
  NOR2_X1 U12643 ( .A1(n13580), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11601) );
  AOI21_X1 U12644 ( .B1(n14675), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n11601), .ZN(
        n10129) );
  OAI21_X1 U12645 ( .B1(n10130), .B2(n14673), .A(n10129), .ZN(n10138) );
  NAND2_X1 U12646 ( .A1(n10131), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10150) );
  MUX2_X1 U12647 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n8445), .S(n10145), .Z(
        n10149) );
  AOI21_X1 U12648 ( .B1(n10151), .B2(n10150), .A(n10149), .ZN(n10148) );
  NOR2_X1 U12649 ( .A1(n10145), .A2(n8445), .ZN(n10134) );
  MUX2_X1 U12650 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10132), .S(n10189), .Z(
        n10133) );
  OAI21_X1 U12651 ( .B1(n10148), .B2(n10134), .A(n10133), .ZN(n10184) );
  INV_X1 U12652 ( .A(n10184), .ZN(n10136) );
  NOR3_X1 U12653 ( .A1(n10148), .A2(n10134), .A3(n10133), .ZN(n10135) );
  NOR3_X1 U12654 ( .A1(n10136), .A2(n10135), .A3(n14690), .ZN(n10137) );
  AOI211_X1 U12655 ( .C1(n14684), .C2(n10139), .A(n10138), .B(n10137), .ZN(
        n10140) );
  INV_X1 U12656 ( .A(n10140), .ZN(P1_U3252) );
  INV_X1 U12657 ( .A(n10141), .ZN(n10142) );
  AOI21_X1 U12658 ( .B1(n10144), .B2(n10143), .A(n10142), .ZN(n10156) );
  NAND2_X1 U12659 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11519) );
  INV_X1 U12660 ( .A(n11519), .ZN(n10147) );
  NOR2_X1 U12661 ( .A1(n14673), .A2(n10145), .ZN(n10146) );
  AOI211_X1 U12662 ( .C1(n14675), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10147), .B(
        n10146), .ZN(n10155) );
  INV_X1 U12663 ( .A(n10148), .ZN(n10153) );
  NAND3_X1 U12664 ( .A1(n10151), .A2(n10150), .A3(n10149), .ZN(n10152) );
  NAND3_X1 U12665 ( .A1(n10153), .A2(n14669), .A3(n10152), .ZN(n10154) );
  OAI211_X1 U12666 ( .C1(n10156), .C2(n13940), .A(n10155), .B(n10154), .ZN(
        P1_U3251) );
  INV_X1 U12667 ( .A(n10157), .ZN(n10160) );
  INV_X1 U12668 ( .A(n14964), .ZN(n10158) );
  OAI222_X1 U12669 ( .A1(n13776), .A2(n10159), .B1(n11134), .B2(n10160), .C1(
        P2_U3088), .C2(n10158), .ZN(P2_U3317) );
  INV_X1 U12670 ( .A(n10240), .ZN(n10246) );
  OAI222_X1 U12671 ( .A1(n14298), .A2(n10161), .B1(n14304), .B2(n10160), .C1(
        n10246), .C2(P1_U3086), .ZN(P1_U3345) );
  OAI222_X1 U12672 ( .A1(P3_U3151), .A2(n15217), .B1(n12962), .B2(n10163), 
        .C1(n12961), .C2(n10162), .ZN(P3_U3281) );
  NAND2_X1 U12673 ( .A1(n10960), .A2(n14655), .ZN(n10164) );
  OAI21_X1 U12674 ( .B1(n14655), .B2(n9223), .A(n10164), .ZN(P1_U3560) );
  NAND2_X1 U12675 ( .A1(n10166), .A2(n10165), .ZN(n10168) );
  NAND2_X1 U12676 ( .A1(n10168), .A2(n10167), .ZN(n10169) );
  NAND2_X1 U12677 ( .A1(n10170), .A2(n10169), .ZN(n10179) );
  NOR2_X1 U12678 ( .A1(n8145), .A2(P2_U3088), .ZN(n13481) );
  NAND2_X1 U12679 ( .A1(n10172), .A2(n10171), .ZN(n15018) );
  OAI22_X1 U12680 ( .A1(n15022), .A2(n10174), .B1(n10173), .B2(n15018), .ZN(
        n10178) );
  NAND2_X1 U12681 ( .A1(n15041), .A2(n10174), .ZN(n10176) );
  AND2_X1 U12682 ( .A1(n8145), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10175) );
  OAI211_X1 U12683 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n15018), .A(n10176), .B(
        n15046), .ZN(n10177) );
  MUX2_X1 U12684 ( .A(n10178), .B(n10177), .S(n13777), .Z(n10181) );
  INV_X1 U12685 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11006) );
  OAI22_X1 U12686 ( .A1(n15050), .A2(n15400), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11006), .ZN(n10180) );
  OR2_X1 U12687 ( .A1(n10181), .A2(n10180), .ZN(P2_U3214) );
  NAND2_X1 U12688 ( .A1(n10189), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10183) );
  MUX2_X1 U12689 ( .A(n8470), .B(P1_REG2_REG_10__SCAN_IN), .S(n10240), .Z(
        n10182) );
  AOI21_X1 U12690 ( .B1(n10184), .B2(n10183), .A(n10182), .ZN(n10252) );
  NAND3_X1 U12691 ( .A1(n10184), .A2(n10183), .A3(n10182), .ZN(n10185) );
  NAND2_X1 U12692 ( .A1(n10185), .A2(n14669), .ZN(n10197) );
  INV_X1 U12693 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n11646) );
  NOR2_X1 U12694 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11646), .ZN(n10187) );
  NOR2_X1 U12695 ( .A1(n14673), .A2(n10246), .ZN(n10186) );
  AOI211_X1 U12696 ( .C1(n14675), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n10187), 
        .B(n10186), .ZN(n10196) );
  MUX2_X1 U12697 ( .A(n10188), .B(P1_REG1_REG_10__SCAN_IN), .S(n10240), .Z(
        n10192) );
  OR2_X1 U12698 ( .A1(n10189), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10190) );
  NAND2_X1 U12699 ( .A1(n10191), .A2(n10190), .ZN(n10193) );
  AOI21_X1 U12700 ( .B1(n10192), .B2(n10193), .A(n13940), .ZN(n10194) );
  OR2_X1 U12701 ( .A1(n10193), .A2(n10192), .ZN(n10242) );
  NAND2_X1 U12702 ( .A1(n10194), .A2(n10242), .ZN(n10195) );
  OAI211_X1 U12703 ( .C1(n10252), .C2(n10197), .A(n10196), .B(n10195), .ZN(
        P1_U3253) );
  INV_X1 U12704 ( .A(n10198), .ZN(n10201) );
  INV_X1 U12705 ( .A(n10372), .ZN(n10365) );
  OAI222_X1 U12706 ( .A1(n14298), .A2(n10199), .B1(n14304), .B2(n10201), .C1(
        P1_U3086), .C2(n10365), .ZN(P1_U3344) );
  INV_X1 U12707 ( .A(n13122), .ZN(n10200) );
  OAI222_X1 U12708 ( .A1(n13776), .A2(n10202), .B1(n11134), .B2(n10201), .C1(
        P2_U3088), .C2(n10200), .ZN(P2_U3316) );
  CLKBUF_X1 U12709 ( .A(n10205), .Z(n10232) );
  INV_X1 U12710 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10204) );
  NOR2_X1 U12711 ( .A1(n10232), .A2(n10204), .ZN(P3_U3263) );
  INV_X1 U12712 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10206) );
  NOR2_X1 U12713 ( .A1(n10232), .A2(n10206), .ZN(P3_U3262) );
  INV_X1 U12714 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10207) );
  NOR2_X1 U12715 ( .A1(n10205), .A2(n10207), .ZN(P3_U3260) );
  INV_X1 U12716 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10208) );
  NOR2_X1 U12717 ( .A1(n10232), .A2(n10208), .ZN(P3_U3259) );
  INV_X1 U12718 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10209) );
  NOR2_X1 U12719 ( .A1(n10232), .A2(n10209), .ZN(P3_U3261) );
  INV_X1 U12720 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10210) );
  NOR2_X1 U12721 ( .A1(n10205), .A2(n10210), .ZN(P3_U3258) );
  INV_X1 U12722 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10211) );
  NOR2_X1 U12723 ( .A1(n10232), .A2(n10211), .ZN(P3_U3257) );
  INV_X1 U12724 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10212) );
  NOR2_X1 U12725 ( .A1(n10232), .A2(n10212), .ZN(P3_U3256) );
  INV_X1 U12726 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10213) );
  NOR2_X1 U12727 ( .A1(n10232), .A2(n10213), .ZN(P3_U3255) );
  INV_X1 U12728 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10214) );
  NOR2_X1 U12729 ( .A1(n10232), .A2(n10214), .ZN(P3_U3254) );
  INV_X1 U12730 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10215) );
  NOR2_X1 U12731 ( .A1(n10232), .A2(n10215), .ZN(P3_U3253) );
  INV_X1 U12732 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10216) );
  NOR2_X1 U12733 ( .A1(n10232), .A2(n10216), .ZN(P3_U3252) );
  INV_X1 U12734 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10217) );
  NOR2_X1 U12735 ( .A1(n10232), .A2(n10217), .ZN(P3_U3251) );
  INV_X1 U12736 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10218) );
  NOR2_X1 U12737 ( .A1(n10232), .A2(n10218), .ZN(P3_U3250) );
  INV_X1 U12738 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10219) );
  NOR2_X1 U12739 ( .A1(n10232), .A2(n10219), .ZN(P3_U3249) );
  INV_X1 U12740 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10220) );
  NOR2_X1 U12741 ( .A1(n10205), .A2(n10220), .ZN(P3_U3234) );
  INV_X1 U12742 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n13610) );
  NOR2_X1 U12743 ( .A1(n10205), .A2(n13610), .ZN(P3_U3235) );
  INV_X1 U12744 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10221) );
  NOR2_X1 U12745 ( .A1(n10205), .A2(n10221), .ZN(P3_U3236) );
  INV_X1 U12746 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10222) );
  NOR2_X1 U12747 ( .A1(n10205), .A2(n10222), .ZN(P3_U3237) );
  INV_X1 U12748 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n13651) );
  NOR2_X1 U12749 ( .A1(n10205), .A2(n13651), .ZN(P3_U3238) );
  INV_X1 U12750 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10223) );
  NOR2_X1 U12751 ( .A1(n10205), .A2(n10223), .ZN(P3_U3239) );
  INV_X1 U12752 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10224) );
  NOR2_X1 U12753 ( .A1(n10205), .A2(n10224), .ZN(P3_U3240) );
  INV_X1 U12754 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10225) );
  NOR2_X1 U12755 ( .A1(n10205), .A2(n10225), .ZN(P3_U3241) );
  INV_X1 U12756 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10226) );
  NOR2_X1 U12757 ( .A1(n10205), .A2(n10226), .ZN(P3_U3242) );
  INV_X1 U12758 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10227) );
  NOR2_X1 U12759 ( .A1(n10232), .A2(n10227), .ZN(P3_U3243) );
  INV_X1 U12760 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10228) );
  NOR2_X1 U12761 ( .A1(n10232), .A2(n10228), .ZN(P3_U3244) );
  INV_X1 U12762 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10229) );
  NOR2_X1 U12763 ( .A1(n10232), .A2(n10229), .ZN(P3_U3245) );
  INV_X1 U12764 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10230) );
  NOR2_X1 U12765 ( .A1(n10232), .A2(n10230), .ZN(P3_U3246) );
  INV_X1 U12766 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10231) );
  NOR2_X1 U12767 ( .A1(n10232), .A2(n10231), .ZN(P3_U3247) );
  INV_X1 U12768 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n13688) );
  NOR2_X1 U12769 ( .A1(n10232), .A2(n13688), .ZN(P3_U3248) );
  MUX2_X1 U12770 ( .A(n10233), .B(n10781), .S(n14655), .Z(n10234) );
  INV_X1 U12771 ( .A(n10234), .ZN(P1_U3561) );
  MUX2_X1 U12772 ( .A(n10235), .B(n11600), .S(n14655), .Z(n10236) );
  INV_X1 U12773 ( .A(n10236), .ZN(P1_U3568) );
  MUX2_X1 U12774 ( .A(n10237), .B(n11598), .S(n14655), .Z(n10238) );
  INV_X1 U12775 ( .A(n10238), .ZN(P1_U3569) );
  MUX2_X1 U12776 ( .A(n10319), .B(n14494), .S(n14655), .Z(n10239) );
  INV_X1 U12777 ( .A(n10239), .ZN(P1_U3573) );
  NAND2_X1 U12778 ( .A1(n10240), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10241) );
  AND2_X1 U12779 ( .A1(n10242), .A2(n10241), .ZN(n10245) );
  MUX2_X1 U12780 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10243), .S(n10372), .Z(
        n10244) );
  NAND2_X1 U12781 ( .A1(n10245), .A2(n10244), .ZN(n10374) );
  OAI21_X1 U12782 ( .B1(n10245), .B2(n10244), .A(n10374), .ZN(n10257) );
  NOR2_X1 U12783 ( .A1(n10246), .A2(n8470), .ZN(n10250) );
  INV_X1 U12784 ( .A(n10250), .ZN(n10248) );
  INV_X1 U12785 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10364) );
  MUX2_X1 U12786 ( .A(n10364), .B(P1_REG2_REG_11__SCAN_IN), .S(n10372), .Z(
        n10247) );
  NAND2_X1 U12787 ( .A1(n10248), .A2(n10247), .ZN(n10251) );
  MUX2_X1 U12788 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10364), .S(n10372), .Z(
        n10249) );
  OAI21_X1 U12789 ( .B1(n10252), .B2(n10250), .A(n10249), .ZN(n10363) );
  OAI211_X1 U12790 ( .C1(n10252), .C2(n10251), .A(n10363), .B(n14669), .ZN(
        n10255) );
  NAND2_X1 U12791 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14538)
         );
  INV_X1 U12792 ( .A(n14538), .ZN(n10253) );
  AOI21_X1 U12793 ( .B1(n14675), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n10253), 
        .ZN(n10254) );
  OAI211_X1 U12794 ( .C1(n10365), .C2(n14673), .A(n10255), .B(n10254), .ZN(
        n10256) );
  AOI21_X1 U12795 ( .B1(n14684), .B2(n10257), .A(n10256), .ZN(n10258) );
  INV_X1 U12796 ( .A(n10258), .ZN(P1_U3254) );
  INV_X1 U12797 ( .A(n14372), .ZN(n12590) );
  OAI222_X1 U12798 ( .A1(P3_U3151), .A2(n12590), .B1(n12962), .B2(n13582), 
        .C1(n12961), .C2(n10259), .ZN(P3_U3279) );
  INV_X1 U12799 ( .A(n10779), .ZN(n10388) );
  INV_X1 U12800 ( .A(n10260), .ZN(n10261) );
  NAND2_X1 U12801 ( .A1(n10788), .A2(n11360), .ZN(n10289) );
  OR2_X2 U12802 ( .A1(n10289), .A2(n10789), .ZN(n14745) );
  AOI21_X1 U12803 ( .B1(n6618), .B2(n10270), .A(n10390), .ZN(n14651) );
  OR2_X1 U12804 ( .A1(n10287), .A2(P1_D_REG_0__SCAN_IN), .ZN(n10275) );
  NOR2_X1 U12805 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .ZN(
        n10279) );
  NOR4_X1 U12806 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_30__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n10278) );
  NOR4_X1 U12807 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n10277) );
  NOR4_X1 U12808 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n10276) );
  NAND4_X1 U12809 ( .A1(n10279), .A2(n10278), .A3(n10277), .A4(n10276), .ZN(
        n10285) );
  NOR4_X1 U12810 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n10283) );
  NOR4_X1 U12811 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n10282) );
  NOR4_X1 U12812 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n10281) );
  NOR4_X1 U12813 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n10280) );
  NAND4_X1 U12814 ( .A1(n10283), .A2(n10282), .A3(n10281), .A4(n10280), .ZN(
        n10284) );
  NOR2_X1 U12815 ( .A1(n10285), .A2(n10284), .ZN(n10286) );
  OR2_X1 U12816 ( .A1(n10287), .A2(n10286), .ZN(n10295) );
  NAND3_X1 U12817 ( .A1(n11567), .A2(n11583), .A3(n10295), .ZN(n10297) );
  NOR2_X1 U12818 ( .A1(n10297), .A2(n10288), .ZN(n10301) );
  INV_X1 U12819 ( .A(n10289), .ZN(n14765) );
  NAND2_X1 U12820 ( .A1(n14765), .A2(n10937), .ZN(n10292) );
  INV_X1 U12821 ( .A(n10290), .ZN(n10291) );
  INV_X1 U12822 ( .A(n10300), .ZN(n14560) );
  NOR2_X1 U12823 ( .A1(n14833), .A2(n10296), .ZN(n10293) );
  AND2_X1 U12824 ( .A1(n10302), .A2(n10294), .ZN(n10298) );
  AND2_X1 U12825 ( .A1(n10298), .A2(n10295), .ZN(n11569) );
  AND2_X1 U12826 ( .A1(n11569), .A2(n11567), .ZN(n10778) );
  AND2_X1 U12827 ( .A1(n14517), .A2(n14177), .ZN(n14547) );
  INV_X1 U12828 ( .A(n11582), .ZN(n11570) );
  NAND2_X1 U12829 ( .A1(n10297), .A2(n11570), .ZN(n10755) );
  NAND2_X1 U12830 ( .A1(n10755), .A2(n10298), .ZN(n10506) );
  AOI22_X1 U12831 ( .A1(n14547), .A2(n10299), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n10506), .ZN(n10305) );
  NAND2_X1 U12832 ( .A1(n10301), .A2(n10300), .ZN(n10303) );
  NAND2_X1 U12833 ( .A1(n14536), .A2(n8319), .ZN(n10304) );
  OAI211_X1 U12834 ( .C1(n14651), .C2(n14532), .A(n10305), .B(n10304), .ZN(
        P1_U3232) );
  NAND2_X1 U12835 ( .A1(n8198), .A2(n13340), .ZN(n10307) );
  NOR2_X1 U12836 ( .A1(n6745), .A2(n14443), .ZN(n10306) );
  AOI21_X1 U12837 ( .B1(n11009), .B2(n10307), .A(n10306), .ZN(n11007) );
  INV_X1 U12838 ( .A(n10308), .ZN(n15097) );
  AOI22_X1 U12839 ( .A1(n11009), .A2(n15097), .B1(n11005), .B2(n10407), .ZN(
        n10309) );
  NAND2_X1 U12840 ( .A1(n11007), .A2(n10309), .ZN(n10385) );
  NAND2_X1 U12841 ( .A1(n15099), .A2(n10385), .ZN(n10310) );
  OAI21_X1 U12842 ( .B1(n15099), .B2(n7575), .A(n10310), .ZN(P2_U3430) );
  INV_X1 U12843 ( .A(n10607), .ZN(n10600) );
  INV_X1 U12844 ( .A(n10311), .ZN(n10314) );
  OAI222_X1 U12845 ( .A1(P1_U3086), .A2(n10600), .B1(n14304), .B2(n10314), 
        .C1(n10312), .C2(n14298), .ZN(P1_U3343) );
  INV_X1 U12846 ( .A(n13139), .ZN(n10313) );
  OAI222_X1 U12847 ( .A1(n13776), .A2(n10315), .B1(n11134), .B2(n10314), .C1(
        n10313), .C2(P2_U3088), .ZN(P2_U3315) );
  OAI222_X1 U12848 ( .A1(n14397), .A2(P3_U3151), .B1(n12961), .B2(n10317), 
        .C1(n10316), .C2(n12962), .ZN(P3_U3278) );
  INV_X1 U12849 ( .A(n10318), .ZN(n10320) );
  OAI222_X1 U12850 ( .A1(P2_U3088), .A2(n13141), .B1(n11134), .B2(n10320), 
        .C1(n10319), .C2(n13776), .ZN(P2_U3314) );
  INV_X1 U12851 ( .A(n10688), .ZN(n10694) );
  OAI222_X1 U12852 ( .A1(n14298), .A2(n10321), .B1(n14304), .B2(n10320), .C1(
        P1_U3086), .C2(n10694), .ZN(P1_U3342) );
  INV_X1 U12853 ( .A(n10354), .ZN(n14944) );
  INV_X1 U12854 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10322) );
  MUX2_X1 U12855 ( .A(n10322), .B(P2_REG2_REG_1__SCAN_IN), .S(n14868), .Z(
        n14862) );
  AND2_X1 U12856 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n13777), .ZN(n14861) );
  NAND2_X1 U12857 ( .A1(n14862), .A2(n14861), .ZN(n14860) );
  INV_X1 U12858 ( .A(n14868), .ZN(n10339) );
  NAND2_X1 U12859 ( .A1(n10339), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10323) );
  NAND2_X1 U12860 ( .A1(n14860), .A2(n10323), .ZN(n14874) );
  INV_X1 U12861 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10324) );
  MUX2_X1 U12862 ( .A(n10324), .B(P2_REG2_REG_2__SCAN_IN), .S(n14879), .Z(
        n14875) );
  NAND2_X1 U12863 ( .A1(n14874), .A2(n14875), .ZN(n14873) );
  OR2_X1 U12864 ( .A1(n14879), .A2(n10324), .ZN(n10325) );
  NAND2_X1 U12865 ( .A1(n14873), .A2(n10325), .ZN(n13093) );
  INV_X1 U12866 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10326) );
  MUX2_X1 U12867 ( .A(n10326), .B(P2_REG2_REG_3__SCAN_IN), .S(n13090), .Z(
        n13094) );
  NAND2_X1 U12868 ( .A1(n13093), .A2(n13094), .ZN(n13092) );
  OR2_X1 U12869 ( .A1(n13090), .A2(n10326), .ZN(n10327) );
  NAND2_X1 U12870 ( .A1(n13092), .A2(n10327), .ZN(n14888) );
  MUX2_X1 U12871 ( .A(n7639), .B(P2_REG2_REG_4__SCAN_IN), .S(n10345), .Z(
        n14889) );
  NAND2_X1 U12872 ( .A1(n14888), .A2(n14889), .ZN(n14887) );
  NAND2_X1 U12873 ( .A1(n14893), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10328) );
  NAND2_X1 U12874 ( .A1(n14887), .A2(n10328), .ZN(n13106) );
  MUX2_X1 U12875 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7647), .S(n13104), .Z(
        n13107) );
  NAND2_X1 U12876 ( .A1(n13106), .A2(n13107), .ZN(n13105) );
  NAND2_X1 U12877 ( .A1(n13104), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10329) );
  NAND2_X1 U12878 ( .A1(n13105), .A2(n10329), .ZN(n14902) );
  MUX2_X1 U12879 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11018), .S(n14907), .Z(
        n14903) );
  NAND2_X1 U12880 ( .A1(n14902), .A2(n14903), .ZN(n14901) );
  NAND2_X1 U12881 ( .A1(n14907), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10330) );
  NAND2_X1 U12882 ( .A1(n14901), .A2(n10330), .ZN(n14916) );
  XNOR2_X1 U12883 ( .A(n10349), .B(n15054), .ZN(n14917) );
  NAND2_X1 U12884 ( .A1(n14916), .A2(n14917), .ZN(n14915) );
  NAND2_X1 U12885 ( .A1(n10349), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10331) );
  NAND2_X1 U12886 ( .A1(n14915), .A2(n10331), .ZN(n14929) );
  MUX2_X1 U12887 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11051), .S(n10351), .Z(
        n14930) );
  NAND2_X1 U12888 ( .A1(n14929), .A2(n14930), .ZN(n14928) );
  NAND2_X1 U12889 ( .A1(n10351), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10332) );
  NAND2_X1 U12890 ( .A1(n14928), .A2(n10332), .ZN(n14941) );
  XNOR2_X1 U12891 ( .A(n10354), .B(n10333), .ZN(n14940) );
  OR2_X1 U12892 ( .A1(n14941), .A2(n14940), .ZN(n14943) );
  OAI21_X1 U12893 ( .B1(n14944), .B2(P2_REG2_REG_9__SCAN_IN), .A(n14943), .ZN(
        n14960) );
  XNOR2_X1 U12894 ( .A(n14964), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n14961) );
  NOR2_X1 U12895 ( .A1(n14960), .A2(n14961), .ZN(n14959) );
  AOI21_X1 U12896 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n14964), .A(n14959), 
        .ZN(n10336) );
  MUX2_X1 U12897 ( .A(n11495), .B(P2_REG2_REG_11__SCAN_IN), .S(n13122), .Z(
        n10334) );
  INV_X1 U12898 ( .A(n10334), .ZN(n10335) );
  NAND2_X1 U12899 ( .A1(n10336), .A2(n10335), .ZN(n13121) );
  OAI21_X1 U12900 ( .B1(n10336), .B2(n10335), .A(n13121), .ZN(n10360) );
  NAND2_X1 U12901 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n11365)
         );
  NAND2_X1 U12902 ( .A1(n15028), .A2(n13122), .ZN(n10337) );
  OAI211_X1 U12903 ( .C1(n15050), .C2(n10338), .A(n11365), .B(n10337), .ZN(
        n10359) );
  MUX2_X1 U12904 ( .A(n7558), .B(P2_REG1_REG_1__SCAN_IN), .S(n14868), .Z(
        n14865) );
  AND2_X1 U12905 ( .A1(n13777), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n14864) );
  NAND2_X1 U12906 ( .A1(n14865), .A2(n14864), .ZN(n14863) );
  NAND2_X1 U12907 ( .A1(n10339), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10340) );
  NAND2_X1 U12908 ( .A1(n14863), .A2(n10340), .ZN(n14877) );
  MUX2_X1 U12909 ( .A(n10341), .B(P2_REG1_REG_2__SCAN_IN), .S(n14879), .Z(
        n14878) );
  NAND2_X1 U12910 ( .A1(n14877), .A2(n14878), .ZN(n14876) );
  OR2_X1 U12911 ( .A1(n14879), .A2(n10341), .ZN(n10342) );
  NAND2_X1 U12912 ( .A1(n14876), .A2(n10342), .ZN(n13096) );
  MUX2_X1 U12913 ( .A(n10343), .B(P2_REG1_REG_3__SCAN_IN), .S(n13090), .Z(
        n13097) );
  NAND2_X1 U12914 ( .A1(n13096), .A2(n13097), .ZN(n13095) );
  OR2_X1 U12915 ( .A1(n13090), .A2(n10343), .ZN(n10344) );
  NAND2_X1 U12916 ( .A1(n13095), .A2(n10344), .ZN(n14891) );
  INV_X1 U12917 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n15101) );
  MUX2_X1 U12918 ( .A(n15101), .B(P2_REG1_REG_4__SCAN_IN), .S(n10345), .Z(
        n14892) );
  NAND2_X1 U12919 ( .A1(n14891), .A2(n14892), .ZN(n14890) );
  NAND2_X1 U12920 ( .A1(n14893), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10346) );
  NAND2_X1 U12921 ( .A1(n14890), .A2(n10346), .ZN(n13109) );
  INV_X1 U12922 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10907) );
  MUX2_X1 U12923 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10907), .S(n13104), .Z(
        n13110) );
  NAND2_X1 U12924 ( .A1(n13109), .A2(n13110), .ZN(n13108) );
  NAND2_X1 U12925 ( .A1(n13104), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10347) );
  NAND2_X1 U12926 ( .A1(n13108), .A2(n10347), .ZN(n14905) );
  INV_X1 U12927 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10870) );
  MUX2_X1 U12928 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10870), .S(n14907), .Z(
        n14906) );
  NAND2_X1 U12929 ( .A1(n14905), .A2(n14906), .ZN(n14904) );
  NAND2_X1 U12930 ( .A1(n14907), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10348) );
  NAND2_X1 U12931 ( .A1(n14904), .A2(n10348), .ZN(n14919) );
  MUX2_X1 U12932 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7704), .S(n10349), .Z(
        n14920) );
  NAND2_X1 U12933 ( .A1(n14919), .A2(n14920), .ZN(n14918) );
  NAND2_X1 U12934 ( .A1(n10349), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10350) );
  NAND2_X1 U12935 ( .A1(n14918), .A2(n10350), .ZN(n14932) );
  INV_X1 U12936 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n11159) );
  MUX2_X1 U12937 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n11159), .S(n10351), .Z(
        n14933) );
  NAND2_X1 U12938 ( .A1(n14932), .A2(n14933), .ZN(n14931) );
  NAND2_X1 U12939 ( .A1(n10351), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10352) );
  NAND2_X1 U12940 ( .A1(n14931), .A2(n10352), .ZN(n14947) );
  MUX2_X1 U12941 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10353), .S(n10354), .Z(
        n14946) );
  AOI21_X1 U12942 ( .B1(n10354), .B2(n10353), .A(n14949), .ZN(n14956) );
  MUX2_X1 U12943 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7758), .S(n14964), .Z(
        n14955) );
  AND2_X1 U12944 ( .A1(n14956), .A2(n14955), .ZN(n14957) );
  INV_X1 U12945 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10355) );
  MUX2_X1 U12946 ( .A(n10355), .B(P2_REG1_REG_11__SCAN_IN), .S(n13122), .Z(
        n10356) );
  NOR2_X1 U12947 ( .A1(n10357), .A2(n10356), .ZN(n13114) );
  AOI211_X1 U12948 ( .C1(n10357), .C2(n10356), .A(n15022), .B(n13114), .ZN(
        n10358) );
  AOI211_X1 U12949 ( .C1(n15035), .C2(n10360), .A(n10359), .B(n10358), .ZN(
        n10361) );
  INV_X1 U12950 ( .A(n10361), .ZN(P2_U3225) );
  MUX2_X1 U12951 ( .A(n10362), .B(P1_REG2_REG_12__SCAN_IN), .S(n10607), .Z(
        n10367) );
  OAI21_X1 U12952 ( .B1(n10365), .B2(n10364), .A(n10363), .ZN(n10366) );
  NOR2_X1 U12953 ( .A1(n10366), .A2(n10367), .ZN(n10599) );
  AOI21_X1 U12954 ( .B1(n10367), .B2(n10366), .A(n10599), .ZN(n10380) );
  INV_X1 U12955 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10369) );
  OAI22_X1 U12956 ( .A1(n14695), .A2(n10369), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10368), .ZN(n10370) );
  AOI21_X1 U12957 ( .B1(n10607), .B2(n14687), .A(n10370), .ZN(n10379) );
  MUX2_X1 U12958 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10371), .S(n10607), .Z(
        n10376) );
  OR2_X1 U12959 ( .A1(n10372), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10373) );
  NAND2_X1 U12960 ( .A1(n10374), .A2(n10373), .ZN(n10375) );
  NAND2_X1 U12961 ( .A1(n10375), .A2(n10376), .ZN(n10609) );
  OAI21_X1 U12962 ( .B1(n10376), .B2(n10375), .A(n10609), .ZN(n10377) );
  NAND2_X1 U12963 ( .A1(n10377), .A2(n14684), .ZN(n10378) );
  OAI211_X1 U12964 ( .C1(n10380), .C2(n14690), .A(n10379), .B(n10378), .ZN(
        P1_U3255) );
  NAND2_X1 U12965 ( .A1(n15078), .A2(n10381), .ZN(n10382) );
  NAND2_X1 U12966 ( .A1(n15105), .A2(n10385), .ZN(n10386) );
  OAI21_X1 U12967 ( .B1(n15105), .B2(n10174), .A(n10386), .ZN(P2_U3499) );
  NAND2_X1 U12968 ( .A1(n14307), .A2(n13984), .ZN(n10387) );
  NAND2_X2 U12969 ( .A1(n10388), .A2(n10387), .ZN(n11974) );
  INV_X1 U12970 ( .A(n11974), .ZN(n10389) );
  AOI21_X1 U12971 ( .B1(n6618), .B2(n11786), .A(n10390), .ZN(n10398) );
  INV_X1 U12972 ( .A(n14770), .ZN(n10392) );
  NAND2_X1 U12973 ( .A1(n10392), .A2(n10391), .ZN(n10393) );
  OAI21_X1 U12974 ( .B1(n10396), .B2(n10395), .A(n10496), .ZN(n10397) );
  NOR2_X1 U12975 ( .A1(n10398), .A2(n10397), .ZN(n10498) );
  AOI21_X1 U12976 ( .B1(n10398), .B2(n10397), .A(n10498), .ZN(n10402) );
  NOR2_X1 U12977 ( .A1(n14549), .A2(n14770), .ZN(n10400) );
  AND2_X1 U12978 ( .A1(n14517), .A2(n14178), .ZN(n14545) );
  INV_X1 U12979 ( .A(n14545), .ZN(n14525) );
  OAI22_X1 U12980 ( .A1(n8320), .A2(n14525), .B1(n14526), .B2(n7261), .ZN(
        n10399) );
  AOI211_X1 U12981 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n10506), .A(n10400), .B(
        n10399), .ZN(n10401) );
  OAI21_X1 U12982 ( .B1(n10402), .B2(n14532), .A(n10401), .ZN(P1_U3222) );
  INV_X1 U12983 ( .A(n14404), .ZN(n12597) );
  INV_X1 U12984 ( .A(n10403), .ZN(n10405) );
  INV_X1 U12985 ( .A(SI_18_), .ZN(n10404) );
  OAI222_X1 U12986 ( .A1(n12597), .A2(P3_U3151), .B1(n12961), .B2(n10405), 
        .C1(n10404), .C2(n12962), .ZN(P3_U3277) );
  NOR2_X1 U12987 ( .A1(n10406), .A2(P2_U3088), .ZN(n10459) );
  INV_X1 U12988 ( .A(n13044), .ZN(n13023) );
  AOI22_X1 U12989 ( .A1(n13023), .A2(n13086), .B1(n10407), .B2(n14451), .ZN(
        n10412) );
  NOR2_X1 U12990 ( .A1(n10408), .A2(n14465), .ZN(n10410) );
  OAI21_X1 U12991 ( .B1(n10410), .B2(n10409), .A(n14448), .ZN(n10411) );
  OAI211_X1 U12992 ( .C1(n10459), .C2(n11006), .A(n10412), .B(n10411), .ZN(
        P2_U3204) );
  INV_X1 U12993 ( .A(n11281), .ZN(n10697) );
  INV_X1 U12994 ( .A(n10413), .ZN(n10415) );
  OAI222_X1 U12995 ( .A1(n10697), .A2(P1_U3086), .B1(n14304), .B2(n10415), 
        .C1(n10414), .C2(n14298), .ZN(P1_U3341) );
  INV_X1 U12996 ( .A(n14988), .ZN(n13142) );
  OAI222_X1 U12997 ( .A1(n13776), .A2(n10416), .B1(n11134), .B2(n10415), .C1(
        P2_U3088), .C2(n13142), .ZN(P2_U3313) );
  MUX2_X1 U12998 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12589), .Z(n10534) );
  XNOR2_X1 U12999 ( .A(n10534), .B(n10546), .ZN(n10535) );
  XOR2_X1 U13000 ( .A(n10435), .B(n10417), .Z(n10642) );
  INV_X1 U13001 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10433) );
  MUX2_X1 U13002 ( .A(n10656), .B(n10433), .S(n12589), .Z(n15112) );
  NAND2_X1 U13003 ( .A1(n15112), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15109) );
  OAI22_X1 U13004 ( .A1(n10642), .A2(n15109), .B1(n10417), .B2(n10646), .ZN(
        n10627) );
  MUX2_X1 U13005 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12589), .Z(n10418) );
  XOR2_X1 U13006 ( .A(n10631), .B(n10418), .Z(n10626) );
  INV_X1 U13007 ( .A(n10631), .ZN(n10438) );
  INV_X1 U13008 ( .A(n10418), .ZN(n10419) );
  AOI22_X1 U13009 ( .A1(n10627), .A2(n10626), .B1(n10438), .B2(n10419), .ZN(
        n10536) );
  XOR2_X1 U13010 ( .A(n10535), .B(n10536), .Z(n10446) );
  NAND2_X1 U13011 ( .A1(n10654), .A2(n12512), .ZN(n10430) );
  AOI21_X1 U13012 ( .B1(n12473), .B2(n10422), .A(n10421), .ZN(n10429) );
  AND2_X1 U13013 ( .A1(n10430), .A2(n10429), .ZN(n10432) );
  MUX2_X1 U13014 ( .A(P3_U3897), .B(n10432), .S(n12507), .Z(n15149) );
  INV_X1 U13015 ( .A(n10423), .ZN(n10424) );
  NOR2_X1 U13016 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10656), .ZN(n15106) );
  INV_X1 U13017 ( .A(n15106), .ZN(n10425) );
  NAND2_X1 U13018 ( .A1(n10435), .A2(n10425), .ZN(n10426) );
  NAND2_X1 U13019 ( .A1(n10426), .A2(n7530), .ZN(n10636) );
  OR2_X1 U13020 ( .A1(n10636), .A2(n10635), .ZN(n10638) );
  XNOR2_X1 U13021 ( .A(n10631), .B(n15332), .ZN(n10617) );
  NAND2_X1 U13022 ( .A1(n10616), .A2(n10617), .ZN(n10615) );
  NAND2_X1 U13023 ( .A1(n10631), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10427) );
  NAND2_X1 U13024 ( .A1(n10615), .A2(n10427), .ZN(n10428) );
  XNOR2_X1 U13025 ( .A(n10540), .B(P3_REG2_REG_3__SCAN_IN), .ZN(n10443) );
  INV_X1 U13026 ( .A(n10429), .ZN(n10431) );
  INV_X1 U13027 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10929) );
  NOR2_X1 U13028 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10929), .ZN(n10842) );
  AOI21_X1 U13029 ( .B1(n15215), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10842), .ZN(
        n10442) );
  NAND2_X1 U13030 ( .A1(n10432), .A2(n12589), .ZN(n15108) );
  NOR2_X1 U13031 ( .A1(n10433), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15107) );
  INV_X1 U13032 ( .A(n15107), .ZN(n10436) );
  NOR2_X1 U13033 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10436), .ZN(n10434) );
  AOI21_X1 U13034 ( .B1(n10435), .B2(n10436), .A(n10434), .ZN(n10633) );
  NAND2_X1 U13035 ( .A1(n10633), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10632) );
  OAI21_X1 U13036 ( .B1(P3_IR_REG_1__SCAN_IN), .B2(n10436), .A(n10632), .ZN(
        n10619) );
  MUX2_X1 U13037 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n10437), .S(n10631), .Z(
        n10620) );
  NAND2_X1 U13038 ( .A1(n10619), .A2(n10620), .ZN(n10618) );
  OAI21_X1 U13039 ( .B1(n10438), .B2(n10437), .A(n10618), .ZN(n10547) );
  OAI21_X1 U13040 ( .B1(n10439), .B2(P3_REG1_REG_3__SCAN_IN), .A(n10548), .ZN(
        n10440) );
  NAND2_X1 U13041 ( .A1(n15220), .A2(n10440), .ZN(n10441) );
  OAI211_X1 U13042 ( .C1(n15228), .C2(n10443), .A(n10442), .B(n10441), .ZN(
        n10444) );
  AOI21_X1 U13043 ( .B1(n6765), .B2(n15149), .A(n10444), .ZN(n10445) );
  OAI21_X1 U13044 ( .B1(n10446), .B2(n15184), .A(n10445), .ZN(P3_U3185) );
  OAI21_X1 U13045 ( .B1(n10449), .B2(n10448), .A(n10447), .ZN(n10453) );
  OAI22_X1 U13046 ( .A1(n13017), .A2(n15080), .B1(n10459), .B2(n10450), .ZN(
        n10452) );
  OAI22_X1 U13047 ( .A1(n6745), .A2(n13045), .B1(n13044), .B2(n11077), .ZN(
        n10451) );
  AOI211_X1 U13048 ( .C1(n14448), .C2(n10453), .A(n10452), .B(n10451), .ZN(
        n10454) );
  INV_X1 U13049 ( .A(n10454), .ZN(P2_U3209) );
  OAI21_X1 U13050 ( .B1(n10457), .B2(n10456), .A(n10455), .ZN(n10463) );
  OAI22_X1 U13051 ( .A1(n13017), .A2(n10595), .B1(n10459), .B2(n10458), .ZN(
        n10462) );
  OAI22_X1 U13052 ( .A1(n8155), .A2(n13045), .B1(n13044), .B2(n10460), .ZN(
        n10461) );
  AOI211_X1 U13053 ( .C1(n14448), .C2(n10463), .A(n10462), .B(n10461), .ZN(
        n10464) );
  INV_X1 U13054 ( .A(n10464), .ZN(P2_U3194) );
  INV_X1 U13055 ( .A(n10465), .ZN(n10469) );
  INV_X1 U13056 ( .A(n10466), .ZN(n10468) );
  AOI211_X1 U13057 ( .C1(n15097), .C2(n10469), .A(n10468), .B(n10467), .ZN(
        n10598) );
  NAND2_X1 U13058 ( .A1(n15099), .A2(n14481), .ZN(n13468) );
  INV_X1 U13059 ( .A(n13468), .ZN(n13452) );
  AOI22_X1 U13060 ( .A1(n13452), .A2(n7573), .B1(n15098), .B2(
        P2_REG0_REG_1__SCAN_IN), .ZN(n10470) );
  OAI21_X1 U13061 ( .B1(n10598), .B2(n15098), .A(n10470), .ZN(P2_U3433) );
  AND2_X1 U13062 ( .A1(n12817), .A2(n10575), .ZN(n12338) );
  NOR2_X1 U13063 ( .A1(n12822), .A2(n12338), .ZN(n12479) );
  NAND3_X1 U13064 ( .A1(n10476), .A2(n10492), .A3(n15368), .ZN(n10473) );
  INV_X1 U13065 ( .A(n10478), .ZN(n10471) );
  NAND2_X1 U13066 ( .A1(n10471), .A2(n10488), .ZN(n10472) );
  NAND2_X1 U13067 ( .A1(n10473), .A2(n10472), .ZN(n10475) );
  INV_X1 U13068 ( .A(n10492), .ZN(n10477) );
  NAND2_X1 U13069 ( .A1(n10477), .A2(n10476), .ZN(n10482) );
  OR2_X1 U13070 ( .A1(n10478), .A2(n10488), .ZN(n10479) );
  NAND4_X1 U13071 ( .A1(n10482), .A2(n10481), .A3(n10480), .A4(n10479), .ZN(
        n10483) );
  NAND2_X1 U13072 ( .A1(n10483), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10485) );
  OR2_X1 U13073 ( .A1(n12508), .A2(n10488), .ZN(n10484) );
  AND2_X1 U13074 ( .A1(n10485), .A2(n10484), .ZN(n10816) );
  INV_X1 U13075 ( .A(n10816), .ZN(n10486) );
  NOR2_X1 U13076 ( .A1(n10486), .A2(n12951), .ZN(n10891) );
  INV_X1 U13077 ( .A(n10891), .ZN(n10487) );
  NAND2_X1 U13078 ( .A1(n10487), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10495) );
  INV_X1 U13079 ( .A(n10488), .ZN(n10489) );
  OR2_X1 U13080 ( .A1(n12508), .A2(n10489), .ZN(n10840) );
  INV_X1 U13081 ( .A(n10840), .ZN(n10490) );
  NAND2_X2 U13082 ( .A1(n10490), .A2(n10839), .ZN(n12293) );
  INV_X1 U13083 ( .A(n12293), .ZN(n12236) );
  NOR2_X1 U13084 ( .A1(n10492), .A2(n15313), .ZN(n10493) );
  AOI22_X1 U13085 ( .A1(n12236), .A2(n10491), .B1(n12282), .B2(n10658), .ZN(
        n10494) );
  OAI211_X1 U13086 ( .C1(n12479), .C2(n12285), .A(n10495), .B(n10494), .ZN(
        P3_U3172) );
  INV_X1 U13087 ( .A(n10496), .ZN(n10497) );
  OAI22_X1 U13088 ( .A1(n7261), .A2(n11597), .B1(n14776), .B2(n12036), .ZN(
        n10499) );
  XNOR2_X1 U13089 ( .A(n10499), .B(n11974), .ZN(n10758) );
  INV_X2 U13090 ( .A(n12034), .ZN(n12077) );
  NAND2_X1 U13091 ( .A1(n13898), .A2(n12077), .ZN(n10501) );
  NAND2_X1 U13092 ( .A1(n6812), .A2(n12078), .ZN(n10500) );
  NAND2_X1 U13093 ( .A1(n10501), .A2(n10500), .ZN(n10757) );
  XNOR2_X1 U13094 ( .A(n10758), .B(n10757), .ZN(n10502) );
  AOI21_X1 U13095 ( .B1(n10503), .B2(n10502), .A(n10761), .ZN(n10509) );
  OR2_X1 U13096 ( .A1(n10781), .A2(n14555), .ZN(n10505) );
  NAND2_X1 U13097 ( .A1(n13897), .A2(n14177), .ZN(n10504) );
  NAND2_X1 U13098 ( .A1(n10505), .A2(n10504), .ZN(n10942) );
  AOI22_X1 U13099 ( .A1(n14517), .A2(n10942), .B1(n10506), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10508) );
  NAND2_X1 U13100 ( .A1(n14536), .A2(n6812), .ZN(n10507) );
  OAI211_X1 U13101 ( .C1(n10509), .C2(n14532), .A(n10508), .B(n10507), .ZN(
        P1_U3237) );
  INV_X1 U13102 ( .A(n10510), .ZN(n10512) );
  INV_X1 U13103 ( .A(SI_19_), .ZN(n10511) );
  OAI222_X1 U13104 ( .A1(P3_U3151), .A2(n10513), .B1(n12961), .B2(n10512), 
        .C1(n10511), .C2(n12962), .ZN(P3_U3276) );
  INV_X1 U13105 ( .A(n10514), .ZN(n10515) );
  NOR3_X1 U13106 ( .A1(n12479), .A2(n10515), .A3(n15301), .ZN(n10516) );
  AOI21_X1 U13107 ( .B1(n15322), .B2(n10491), .A(n10516), .ZN(n10655) );
  INV_X1 U13108 ( .A(n12896), .ZN(n10517) );
  AOI22_X1 U13109 ( .A1(n10517), .A2(n10658), .B1(n15392), .B2(
        P3_REG1_REG_0__SCAN_IN), .ZN(n10518) );
  OAI21_X1 U13110 ( .B1(n10655), .B2(n15392), .A(n10518), .ZN(P3_U3459) );
  XNOR2_X1 U13111 ( .A(n10520), .B(n10519), .ZN(n10524) );
  INV_X1 U13112 ( .A(n13045), .ZN(n13027) );
  MUX2_X1 U13113 ( .A(n13014), .B(P2_U3088), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n10522) );
  OAI22_X1 U13114 ( .A1(n10528), .A2(n13044), .B1(n13017), .B2(n11855), .ZN(
        n10521) );
  AOI211_X1 U13115 ( .C1(n13027), .C2(n13085), .A(n10522), .B(n10521), .ZN(
        n10523) );
  OAI21_X1 U13116 ( .B1(n10524), .B2(n13059), .A(n10523), .ZN(P2_U3190) );
  OAI21_X1 U13117 ( .B1(n10527), .B2(n10526), .A(n10525), .ZN(n10532) );
  OAI22_X1 U13118 ( .A1(n10528), .A2(n13045), .B1(n13044), .B2(n10811), .ZN(
        n10531) );
  NAND2_X1 U13119 ( .A1(n14451), .A2(n11242), .ZN(n10529) );
  NAND2_X1 U13120 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n13101) );
  OAI211_X1 U13121 ( .C1(n14453), .C2(n11240), .A(n10529), .B(n13101), .ZN(
        n10530) );
  AOI211_X1 U13122 ( .C1(n10532), .C2(n14448), .A(n10531), .B(n10530), .ZN(
        n10533) );
  INV_X1 U13123 ( .A(n10533), .ZN(P2_U3199) );
  MUX2_X1 U13124 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12589), .Z(n10537) );
  INV_X1 U13125 ( .A(n14321), .ZN(n10550) );
  XNOR2_X1 U13126 ( .A(n10537), .B(n10550), .ZN(n10721) );
  INV_X1 U13127 ( .A(n10537), .ZN(n10538) );
  AOI22_X1 U13128 ( .A1(n10720), .A2(n10721), .B1(n10550), .B2(n10538), .ZN(
        n10737) );
  MUX2_X1 U13129 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12589), .Z(n10539) );
  XNOR2_X1 U13130 ( .A(n10539), .B(n10745), .ZN(n10738) );
  OAI22_X1 U13131 ( .A1(n10737), .A2(n10738), .B1(n10539), .B2(n10745), .ZN(
        n10664) );
  MUX2_X1 U13132 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12589), .Z(n10661) );
  XNOR2_X1 U13133 ( .A(n10661), .B(n10674), .ZN(n10663) );
  XNOR2_X1 U13134 ( .A(n10664), .B(n10663), .ZN(n10564) );
  INV_X1 U13135 ( .A(n10745), .ZN(n10552) );
  AOI22_X1 U13136 ( .A1(P3_REG2_REG_4__SCAN_IN), .A2(n10550), .B1(n14321), 
        .B2(n9283), .ZN(n10722) );
  INV_X1 U13137 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10669) );
  MUX2_X1 U13138 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n10669), .S(n10674), .Z(
        n10543) );
  NAND2_X1 U13139 ( .A1(n10544), .A2(n10543), .ZN(n10545) );
  AOI21_X1 U13140 ( .B1(n10671), .B2(n10545), .A(n15228), .ZN(n10563) );
  AOI22_X1 U13141 ( .A1(P3_REG1_REG_4__SCAN_IN), .A2(n14321), .B1(n10550), 
        .B2(n9280), .ZN(n10726) );
  NAND2_X1 U13142 ( .A1(n10547), .A2(n10546), .ZN(n10549) );
  NAND2_X1 U13143 ( .A1(n10549), .A2(n10548), .ZN(n10725) );
  NAND2_X1 U13144 ( .A1(n10726), .A2(n10725), .ZN(n10724) );
  NAND2_X1 U13145 ( .A1(n10745), .A2(n10551), .ZN(n10553) );
  NAND2_X1 U13146 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n10741), .ZN(n10740) );
  NAND2_X1 U13147 ( .A1(n10553), .A2(n10740), .ZN(n10556) );
  MUX2_X1 U13148 ( .A(n10554), .B(P3_REG1_REG_6__SCAN_IN), .S(n10674), .Z(
        n10555) );
  NAND2_X1 U13149 ( .A1(n10556), .A2(n10555), .ZN(n10673) );
  OAI21_X1 U13150 ( .B1(n10556), .B2(n10555), .A(n10673), .ZN(n10557) );
  INV_X1 U13151 ( .A(n10557), .ZN(n10561) );
  NAND2_X1 U13152 ( .A1(n15149), .A2(n10674), .ZN(n10560) );
  INV_X1 U13153 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10558) );
  NOR2_X1 U13154 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10558), .ZN(n11144) );
  AOI21_X1 U13155 ( .B1(n15215), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11144), .ZN(
        n10559) );
  OAI211_X1 U13156 ( .C1(n10561), .C2(n15108), .A(n10560), .B(n10559), .ZN(
        n10562) );
  AOI211_X1 U13157 ( .C1(n10564), .C2(n15222), .A(n10563), .B(n10562), .ZN(
        n10565) );
  INV_X1 U13158 ( .A(n10565), .ZN(P3_U3188) );
  XNOR2_X1 U13159 ( .A(n10567), .B(n10566), .ZN(n10574) );
  NAND2_X1 U13160 ( .A1(n13082), .A2(n13335), .ZN(n10569) );
  NAND2_X1 U13161 ( .A1(n13080), .A2(n13336), .ZN(n10568) );
  AND2_X1 U13162 ( .A1(n10569), .A2(n10568), .ZN(n10867) );
  INV_X1 U13163 ( .A(n10867), .ZN(n10570) );
  NAND2_X1 U13164 ( .A1(n14450), .A2(n10570), .ZN(n10571) );
  NAND2_X1 U13165 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n14912) );
  OAI211_X1 U13166 ( .C1(n14453), .C2(n11019), .A(n10571), .B(n14912), .ZN(
        n10572) );
  AOI21_X1 U13167 ( .B1(n10869), .B2(n14451), .A(n10572), .ZN(n10573) );
  OAI21_X1 U13168 ( .B1(n10574), .B2(n13059), .A(n10573), .ZN(P2_U3211) );
  OAI22_X1 U13169 ( .A1(n10575), .A2(n12949), .B1(n15379), .B2(n9242), .ZN(
        n10576) );
  INV_X1 U13170 ( .A(n10576), .ZN(n10577) );
  OAI21_X1 U13171 ( .B1(n10655), .B2(n15378), .A(n10577), .ZN(P3_U3390) );
  OR2_X1 U13172 ( .A1(n10579), .A2(n10578), .ZN(n10580) );
  NAND2_X1 U13173 ( .A1(n10581), .A2(n10580), .ZN(n11857) );
  OAI211_X1 U13174 ( .C1(n11086), .C2(n11855), .A(n14465), .B(n11039), .ZN(
        n11861) );
  INV_X1 U13175 ( .A(n11861), .ZN(n10589) );
  INV_X1 U13176 ( .A(n8198), .ZN(n13333) );
  NAND2_X1 U13177 ( .A1(n11857), .A2(n13333), .ZN(n10588) );
  OAI21_X1 U13178 ( .B1(n10584), .B2(n10583), .A(n10582), .ZN(n10585) );
  NAND2_X1 U13179 ( .A1(n10585), .A2(n14456), .ZN(n10587) );
  AOI22_X1 U13180 ( .A1(n13335), .A2(n13085), .B1(n13083), .B2(n13336), .ZN(
        n10586) );
  NAND3_X1 U13181 ( .A1(n10588), .A2(n10587), .A3(n10586), .ZN(n11854) );
  AOI211_X1 U13182 ( .C1(n15097), .C2(n11857), .A(n10589), .B(n11854), .ZN(
        n10594) );
  OAI22_X1 U13183 ( .A1(n13468), .A2(n11855), .B1(n15099), .B2(n7607), .ZN(
        n10590) );
  INV_X1 U13184 ( .A(n10590), .ZN(n10591) );
  OAI21_X1 U13185 ( .B1(n10594), .B2(n15098), .A(n10591), .ZN(P2_U3439) );
  OAI22_X1 U13186 ( .A1(n13418), .A2(n11855), .B1(n15105), .B2(n10343), .ZN(
        n10592) );
  INV_X1 U13187 ( .A(n10592), .ZN(n10593) );
  OAI21_X1 U13188 ( .B1(n10594), .B2(n15103), .A(n10593), .ZN(P2_U3502) );
  OAI22_X1 U13189 ( .A1(n13418), .A2(n10595), .B1(n15105), .B2(n7558), .ZN(
        n10596) );
  INV_X1 U13190 ( .A(n10596), .ZN(n10597) );
  OAI21_X1 U13191 ( .B1(n10598), .B2(n15103), .A(n10597), .ZN(P2_U3500) );
  AOI21_X1 U13192 ( .B1(n10362), .B2(n10600), .A(n10599), .ZN(n10602) );
  MUX2_X1 U13193 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n11540), .S(n10688), .Z(
        n10601) );
  NAND2_X1 U13194 ( .A1(n10602), .A2(n10601), .ZN(n10693) );
  OAI211_X1 U13195 ( .C1(n10602), .C2(n10601), .A(n10693), .B(n14669), .ZN(
        n10605) );
  NOR2_X1 U13196 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13746), .ZN(n10603) );
  AOI21_X1 U13197 ( .B1(n14675), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10603), 
        .ZN(n10604) );
  OAI211_X1 U13198 ( .C1(n14673), .C2(n10694), .A(n10605), .B(n10604), .ZN(
        n10614) );
  MUX2_X1 U13199 ( .A(n10606), .B(P1_REG1_REG_13__SCAN_IN), .S(n10688), .Z(
        n10612) );
  OR2_X1 U13200 ( .A1(n10607), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10608) );
  NAND2_X1 U13201 ( .A1(n10609), .A2(n10608), .ZN(n10611) );
  INV_X1 U13202 ( .A(n10690), .ZN(n10610) );
  AOI211_X1 U13203 ( .C1(n10612), .C2(n10611), .A(n13940), .B(n10610), .ZN(
        n10613) );
  OR2_X1 U13204 ( .A1(n10614), .A2(n10613), .ZN(P1_U3256) );
  INV_X1 U13205 ( .A(n15149), .ZN(n15218) );
  OAI21_X1 U13206 ( .B1(n10617), .B2(n10616), .A(n10615), .ZN(n10625) );
  OAI21_X1 U13207 ( .B1(n10620), .B2(n10619), .A(n10618), .ZN(n10621) );
  AND2_X1 U13208 ( .A1(n15220), .A2(n10621), .ZN(n10624) );
  INV_X1 U13209 ( .A(n15215), .ZN(n15156) );
  INV_X1 U13210 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10622) );
  OAI22_X1 U13211 ( .A1(n15156), .A2(n10622), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15311), .ZN(n10623) );
  AOI211_X1 U13212 ( .C1(n15151), .C2(n10625), .A(n10624), .B(n10623), .ZN(
        n10630) );
  XNOR2_X1 U13213 ( .A(n10627), .B(n10626), .ZN(n10628) );
  NAND2_X1 U13214 ( .A1(n10628), .A2(n15222), .ZN(n10629) );
  OAI211_X1 U13215 ( .C1(n15218), .C2(n10631), .A(n10630), .B(n10629), .ZN(
        P3_U3184) );
  OAI21_X1 U13216 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n10633), .A(n10632), .ZN(
        n10641) );
  INV_X1 U13217 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n10634) );
  OAI22_X1 U13218 ( .A1(n15156), .A2(n10634), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12828), .ZN(n10640) );
  NAND2_X1 U13219 ( .A1(n10636), .A2(n10635), .ZN(n10637) );
  AOI21_X1 U13220 ( .B1(n10638), .B2(n10637), .A(n15228), .ZN(n10639) );
  AOI211_X1 U13221 ( .C1(n15220), .C2(n10641), .A(n10640), .B(n10639), .ZN(
        n10645) );
  XNOR2_X1 U13222 ( .A(n10642), .B(n15109), .ZN(n10643) );
  NAND2_X1 U13223 ( .A1(n10643), .A2(n15222), .ZN(n10644) );
  OAI211_X1 U13224 ( .C1(n15218), .C2(n10646), .A(n10645), .B(n10644), .ZN(
        P3_U3183) );
  NAND2_X1 U13225 ( .A1(n10648), .A2(n10647), .ZN(n10651) );
  NAND2_X1 U13226 ( .A1(n10649), .A2(n12950), .ZN(n10650) );
  AND2_X1 U13227 ( .A1(n10651), .A2(n10650), .ZN(n10653) );
  NAND2_X1 U13228 ( .A1(n10653), .A2(n10652), .ZN(n10657) );
  INV_X1 U13229 ( .A(n15313), .ZN(n12476) );
  MUX2_X1 U13230 ( .A(n10656), .B(n10655), .S(n15330), .Z(n10660) );
  OR2_X1 U13231 ( .A1(n10657), .A2(n15313), .ZN(n11236) );
  INV_X1 U13232 ( .A(n12812), .ZN(n12695) );
  AOI22_X1 U13233 ( .A1(n12695), .A2(n10658), .B1(n15253), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10659) );
  NAND2_X1 U13234 ( .A1(n10660), .A2(n10659), .ZN(P3_U3233) );
  INV_X1 U13235 ( .A(n10661), .ZN(n10662) );
  AOI22_X1 U13236 ( .A1(n10664), .A2(n10663), .B1(n10674), .B2(n10662), .ZN(
        n10703) );
  MUX2_X1 U13237 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12589), .Z(n10665) );
  XNOR2_X1 U13238 ( .A(n10665), .B(n10711), .ZN(n10704) );
  OAI22_X1 U13239 ( .A1(n10703), .A2(n10704), .B1(n10665), .B2(n10711), .ZN(
        n10667) );
  MUX2_X1 U13240 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12589), .Z(n12565) );
  XNOR2_X1 U13241 ( .A(n12565), .B(n12531), .ZN(n10666) );
  NAND2_X1 U13242 ( .A1(n10667), .A2(n10666), .ZN(n12566) );
  OAI21_X1 U13243 ( .B1(n10667), .B2(n10666), .A(n12566), .ZN(n10668) );
  NAND2_X1 U13244 ( .A1(n10668), .A2(n15222), .ZN(n10687) );
  INV_X1 U13245 ( .A(n10711), .ZN(n10676) );
  OR2_X1 U13246 ( .A1(n10674), .A2(n10669), .ZN(n10670) );
  XOR2_X1 U13247 ( .A(n10711), .B(n10672), .Z(n10705) );
  AOI22_X1 U13248 ( .A1(n12531), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n9361), .B2(
        n12564), .ZN(n12544) );
  XNOR2_X1 U13249 ( .A(n12545), .B(n12544), .ZN(n10685) );
  INV_X1 U13250 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15389) );
  AOI22_X1 U13251 ( .A1(n12531), .A2(n15389), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n12564), .ZN(n10679) );
  NAND2_X1 U13252 ( .A1(n10711), .A2(n10675), .ZN(n10677) );
  XNOR2_X1 U13253 ( .A(n10676), .B(n10675), .ZN(n10707) );
  NAND2_X1 U13254 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n10707), .ZN(n10706) );
  NAND2_X1 U13255 ( .A1(n10677), .A2(n10706), .ZN(n10678) );
  NAND2_X1 U13256 ( .A1(n10679), .A2(n10678), .ZN(n12530) );
  OAI21_X1 U13257 ( .B1(n10679), .B2(n10678), .A(n12530), .ZN(n10680) );
  NAND2_X1 U13258 ( .A1(n10680), .A2(n15220), .ZN(n10683) );
  NOR2_X1 U13259 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10681), .ZN(n11307) );
  AOI21_X1 U13260 ( .B1(n15215), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11307), .ZN(
        n10682) );
  OAI211_X1 U13261 ( .C1(n15218), .C2(n12564), .A(n10683), .B(n10682), .ZN(
        n10684) );
  AOI21_X1 U13262 ( .B1(n10685), .B2(n15151), .A(n10684), .ZN(n10686) );
  NAND2_X1 U13263 ( .A1(n10687), .A2(n10686), .ZN(P3_U3190) );
  MUX2_X1 U13264 ( .A(n8527), .B(P1_REG1_REG_14__SCAN_IN), .S(n11281), .Z(
        n10692) );
  NAND2_X1 U13265 ( .A1(n10688), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10689) );
  NAND2_X1 U13266 ( .A1(n10690), .A2(n10689), .ZN(n10691) );
  NOR2_X1 U13267 ( .A1(n10691), .A2(n10692), .ZN(n11279) );
  AOI21_X1 U13268 ( .B1(n10692), .B2(n10691), .A(n11279), .ZN(n10702) );
  OAI21_X1 U13269 ( .B1(n11540), .B2(n10694), .A(n10693), .ZN(n10696) );
  MUX2_X1 U13270 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11682), .S(n11281), .Z(
        n10695) );
  NAND2_X1 U13271 ( .A1(n11281), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11292) );
  OAI211_X1 U13272 ( .C1(n11281), .C2(P1_REG2_REG_14__SCAN_IN), .A(n10696), 
        .B(n11292), .ZN(n11291) );
  OAI211_X1 U13273 ( .C1(n10696), .C2(n10695), .A(n11291), .B(n14669), .ZN(
        n10701) );
  NAND2_X1 U13274 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14502)
         );
  INV_X1 U13275 ( .A(n14502), .ZN(n10699) );
  NOR2_X1 U13276 ( .A1(n14673), .A2(n10697), .ZN(n10698) );
  AOI211_X1 U13277 ( .C1(n14675), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n10699), 
        .B(n10698), .ZN(n10700) );
  OAI211_X1 U13278 ( .C1(n10702), .C2(n13940), .A(n10701), .B(n10700), .ZN(
        P1_U3257) );
  XOR2_X1 U13279 ( .A(n10703), .B(n10704), .Z(n10715) );
  XOR2_X1 U13280 ( .A(P3_REG2_REG_7__SCAN_IN), .B(n10705), .Z(n10713) );
  OAI21_X1 U13281 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n10707), .A(n10706), .ZN(
        n10708) );
  NAND2_X1 U13282 ( .A1(n10708), .A2(n15220), .ZN(n10710) );
  AND2_X1 U13283 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11202) );
  AOI21_X1 U13284 ( .B1(n15215), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11202), .ZN(
        n10709) );
  OAI211_X1 U13285 ( .C1(n15218), .C2(n10711), .A(n10710), .B(n10709), .ZN(
        n10712) );
  AOI21_X1 U13286 ( .B1(n10713), .B2(n15151), .A(n10712), .ZN(n10714) );
  OAI21_X1 U13287 ( .B1(n10715), .B2(n15184), .A(n10714), .ZN(P3_U3189) );
  INV_X1 U13288 ( .A(n14686), .ZN(n11293) );
  INV_X1 U13289 ( .A(n10716), .ZN(n10718) );
  OAI222_X1 U13290 ( .A1(P1_U3086), .A2(n11293), .B1(n14304), .B2(n10718), 
        .C1(n10717), .C2(n14298), .ZN(P1_U3340) );
  INV_X1 U13291 ( .A(n14999), .ZN(n13145) );
  OAI222_X1 U13292 ( .A1(n13776), .A2(n10719), .B1(n11134), .B2(n10718), .C1(
        n13145), .C2(P2_U3088), .ZN(P2_U3312) );
  XOR2_X1 U13293 ( .A(n10720), .B(n10721), .Z(n10736) );
  XNOR2_X1 U13294 ( .A(n10723), .B(n10722), .ZN(n10734) );
  OAI21_X1 U13295 ( .B1(n10726), .B2(n10725), .A(n10724), .ZN(n10727) );
  NAND2_X1 U13296 ( .A1(n15220), .A2(n10727), .ZN(n10730) );
  INV_X1 U13297 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10728) );
  NOR2_X1 U13298 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10728), .ZN(n10855) );
  INV_X1 U13299 ( .A(n10855), .ZN(n10729) );
  OAI211_X1 U13300 ( .C1(n15156), .C2(n10731), .A(n10730), .B(n10729), .ZN(
        n10733) );
  NOR2_X1 U13301 ( .A1(n15218), .A2(n14321), .ZN(n10732) );
  AOI211_X1 U13302 ( .C1(n15151), .C2(n10734), .A(n10733), .B(n10732), .ZN(
        n10735) );
  OAI21_X1 U13303 ( .B1(n10736), .B2(n15184), .A(n10735), .ZN(P3_U3186) );
  XOR2_X1 U13304 ( .A(n10737), .B(n10738), .Z(n10750) );
  XOR2_X1 U13305 ( .A(P3_REG2_REG_5__SCAN_IN), .B(n10739), .Z(n10748) );
  OAI21_X1 U13306 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n10741), .A(n10740), .ZN(
        n10742) );
  NAND2_X1 U13307 ( .A1(n15220), .A2(n10742), .ZN(n10744) );
  NOR2_X1 U13308 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9300), .ZN(n10999) );
  INV_X1 U13309 ( .A(n10999), .ZN(n10743) );
  OAI211_X1 U13310 ( .C1(n15156), .C2(n8848), .A(n10744), .B(n10743), .ZN(
        n10747) );
  NOR2_X1 U13311 ( .A1(n15218), .A2(n10745), .ZN(n10746) );
  AOI211_X1 U13312 ( .C1(n15151), .C2(n10748), .A(n10747), .B(n10746), .ZN(
        n10749) );
  OAI21_X1 U13313 ( .B1(n10750), .B2(n15184), .A(n10749), .ZN(P3_U3187) );
  OAI222_X1 U13314 ( .A1(n12961), .A2(n10752), .B1(n12962), .B2(n10751), .C1(
        P3_U3151), .C2(n10820), .ZN(P3_U3275) );
  INV_X1 U13315 ( .A(n10753), .ZN(n10754) );
  NAND2_X1 U13316 ( .A1(n10755), .A2(n10754), .ZN(n10756) );
  INV_X1 U13317 ( .A(n10757), .ZN(n10760) );
  INV_X1 U13318 ( .A(n10758), .ZN(n10759) );
  NAND2_X1 U13319 ( .A1(n13897), .A2(n10391), .ZN(n10763) );
  NAND2_X1 U13320 ( .A1(n14782), .A2(n12079), .ZN(n10762) );
  NAND2_X1 U13321 ( .A1(n10763), .A2(n10762), .ZN(n10764) );
  XNOR2_X1 U13322 ( .A(n10764), .B(n11786), .ZN(n11166) );
  AND2_X1 U13323 ( .A1(n14782), .A2(n10391), .ZN(n10765) );
  AOI21_X1 U13324 ( .B1(n13897), .B2(n12077), .A(n10765), .ZN(n11167) );
  XNOR2_X1 U13325 ( .A(n11166), .B(n11167), .ZN(n10766) );
  OAI211_X1 U13326 ( .C1(n10767), .C2(n10766), .A(n11169), .B(n14551), .ZN(
        n10771) );
  INV_X1 U13327 ( .A(n14517), .ZN(n13835) );
  AOI22_X1 U13328 ( .A1(n14178), .A2(n13898), .B1(n13896), .B2(n14177), .ZN(
        n14731) );
  OAI22_X1 U13329 ( .A1(n13835), .A2(n14731), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10768), .ZN(n10769) );
  AOI21_X1 U13330 ( .B1(n14782), .B2(n14536), .A(n10769), .ZN(n10770) );
  OAI211_X1 U13331 ( .C1(n14554), .C2(P1_REG3_REG_3__SCAN_IN), .A(n10771), .B(
        n10770), .ZN(P1_U3218) );
  INV_X1 U13332 ( .A(n13937), .ZN(n13948) );
  INV_X1 U13333 ( .A(n10772), .ZN(n10775) );
  OAI222_X1 U13334 ( .A1(P1_U3086), .A2(n13948), .B1(n14304), .B2(n10775), 
        .C1(n10773), .C2(n14298), .ZN(P1_U3339) );
  INV_X1 U13335 ( .A(n15012), .ZN(n10776) );
  OAI222_X1 U13336 ( .A1(P2_U3088), .A2(n10776), .B1(n11134), .B2(n10775), 
        .C1(n10774), .C2(n13776), .ZN(P2_U3311) );
  INV_X1 U13337 ( .A(n11583), .ZN(n10777) );
  NAND2_X1 U13338 ( .A1(n10778), .A2(n10777), .ZN(n11941) );
  NAND2_X1 U13339 ( .A1(n10779), .A2(n14307), .ZN(n10780) );
  NAND2_X1 U13340 ( .A1(n11786), .A2(n10780), .ZN(n10938) );
  NAND2_X1 U13341 ( .A1(n10960), .A2(n8319), .ZN(n10952) );
  NAND2_X1 U13342 ( .A1(n10781), .A2(n14770), .ZN(n10782) );
  OR2_X1 U13343 ( .A1(n13898), .A2(n6812), .ZN(n10783) );
  NAND2_X1 U13344 ( .A1(n10784), .A2(n10783), .ZN(n14732) );
  NAND2_X1 U13345 ( .A1(n14732), .A2(n10785), .ZN(n10787) );
  OR2_X1 U13346 ( .A1(n13897), .A2(n14782), .ZN(n10786) );
  XNOR2_X1 U13347 ( .A(n11104), .B(n11102), .ZN(n14792) );
  OR2_X1 U13348 ( .A1(n10788), .A2(n13984), .ZN(n10792) );
  NAND2_X1 U13349 ( .A1(n10790), .A2(n10789), .ZN(n10791) );
  INV_X1 U13350 ( .A(n10793), .ZN(n10795) );
  NAND2_X1 U13351 ( .A1(n10795), .A2(n10794), .ZN(n10797) );
  NAND2_X1 U13352 ( .A1(n10797), .A2(n10796), .ZN(n10940) );
  NAND2_X1 U13353 ( .A1(n10941), .A2(n10940), .ZN(n10939) );
  NAND2_X1 U13354 ( .A1(n10939), .A2(n10798), .ZN(n14730) );
  NAND2_X1 U13355 ( .A1(n14730), .A2(n14733), .ZN(n14729) );
  INV_X1 U13356 ( .A(n10799), .ZN(n10800) );
  NAND2_X1 U13357 ( .A1(n10801), .A2(n11102), .ZN(n11093) );
  OAI21_X1 U13358 ( .B1(n10801), .B2(n11102), .A(n11093), .ZN(n10802) );
  AOI222_X1 U13359 ( .A1(n14738), .A2(n10802), .B1(n13895), .B2(n14177), .C1(
        n13897), .C2(n14178), .ZN(n14791) );
  MUX2_X1 U13360 ( .A(n10803), .B(n14791), .S(n14741), .Z(n10807) );
  NAND2_X1 U13361 ( .A1(n10955), .A2(n14776), .ZN(n14746) );
  INV_X1 U13362 ( .A(n14744), .ZN(n10804) );
  INV_X1 U13363 ( .A(n14789), .ZN(n11091) );
  AOI211_X1 U13364 ( .C1(n14789), .C2(n10804), .A(n14745), .B(n6723), .ZN(
        n14788) );
  OAI22_X1 U13365 ( .A1(n14337), .A2(n11091), .B1(n11250), .B2(n14739), .ZN(
        n10805) );
  AOI21_X1 U13366 ( .B1(n14788), .B2(n6575), .A(n10805), .ZN(n10806) );
  OAI211_X1 U13367 ( .C1(n14339), .C2(n14792), .A(n10807), .B(n10806), .ZN(
        P1_U3289) );
  XNOR2_X1 U13368 ( .A(n10809), .B(n10808), .ZN(n10815) );
  OAI22_X1 U13369 ( .A1(n10811), .A2(n14441), .B1(n10810), .B2(n14443), .ZN(
        n10984) );
  AOI22_X1 U13370 ( .A1(n14450), .A2(n10984), .B1(P2_REG3_REG_7__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10812) );
  OAI21_X1 U13371 ( .B1(n15053), .B2(n14453), .A(n10812), .ZN(n10813) );
  AOI21_X1 U13372 ( .B1(n15057), .B2(n14451), .A(n10813), .ZN(n10814) );
  OAI21_X1 U13373 ( .B1(n10815), .B2(n13059), .A(n10814), .ZN(P2_U3185) );
  INV_X1 U13374 ( .A(n10817), .ZN(n10818) );
  NAND2_X1 U13375 ( .A1(n12952), .A2(n10818), .ZN(n10823) );
  NAND2_X1 U13376 ( .A1(n10819), .A2(n12608), .ZN(n10821) );
  NAND2_X4 U13377 ( .A1(n10823), .A2(n10822), .ZN(n12200) );
  NAND2_X1 U13378 ( .A1(n12816), .A2(n12157), .ZN(n10824) );
  NAND2_X1 U13379 ( .A1(n10825), .A2(n10824), .ZN(n10829) );
  XNOR2_X1 U13380 ( .A(n12827), .B(n12200), .ZN(n10826) );
  NAND2_X1 U13381 ( .A1(n10827), .A2(n10826), .ZN(n10830) );
  NAND2_X1 U13382 ( .A1(n10880), .A2(n10830), .ZN(n10885) );
  XNOR2_X1 U13383 ( .A(n10832), .B(n12819), .ZN(n10886) );
  INV_X1 U13384 ( .A(n10832), .ZN(n10833) );
  NAND2_X1 U13385 ( .A1(n10833), .A2(n12819), .ZN(n10835) );
  AND2_X1 U13386 ( .A1(n10884), .A2(n10835), .ZN(n10838) );
  XNOR2_X1 U13387 ( .A(n10843), .B(n10834), .ZN(n10848) );
  XNOR2_X1 U13388 ( .A(n10848), .B(n15293), .ZN(n10837) );
  AND2_X1 U13389 ( .A1(n10837), .A2(n10835), .ZN(n10836) );
  OAI211_X1 U13390 ( .C1(n10838), .C2(n10837), .A(n12269), .B(n10850), .ZN(
        n10847) );
  AOI21_X1 U13391 ( .B1(n12282), .B2(n10843), .A(n10842), .ZN(n10844) );
  OAI21_X1 U13392 ( .B1(n12293), .B2(n10841), .A(n10844), .ZN(n10845) );
  AOI21_X1 U13393 ( .B1(n12291), .B2(n12525), .A(n10845), .ZN(n10846) );
  OAI211_X1 U13394 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12178), .A(n10847), .B(
        n10846), .ZN(P3_U3158) );
  NAND2_X1 U13395 ( .A1(n9277), .A2(n10848), .ZN(n10849) );
  XNOR2_X1 U13396 ( .A(n15302), .B(n12200), .ZN(n10851) );
  NAND2_X1 U13397 ( .A1(n10851), .A2(n10841), .ZN(n10994) );
  OAI21_X1 U13398 ( .B1(n10851), .B2(n10841), .A(n10994), .ZN(n10853) );
  INV_X1 U13399 ( .A(n10995), .ZN(n10852) );
  AOI21_X1 U13400 ( .B1(n10854), .B2(n10853), .A(n10852), .ZN(n10860) );
  AOI21_X1 U13401 ( .B1(n12282), .B2(n15302), .A(n10855), .ZN(n10856) );
  OAI21_X1 U13402 ( .B1(n12293), .B2(n15295), .A(n10856), .ZN(n10858) );
  NOR2_X1 U13403 ( .A1(n12178), .A2(n15303), .ZN(n10857) );
  AOI211_X1 U13404 ( .C1(n12291), .C2(n9277), .A(n10858), .B(n10857), .ZN(
        n10859) );
  OAI21_X1 U13405 ( .B1(n10860), .B2(n12285), .A(n10859), .ZN(P3_U3170) );
  OAI21_X1 U13406 ( .B1(n10862), .B2(n10866), .A(n10861), .ZN(n11015) );
  NAND2_X1 U13407 ( .A1(n10899), .A2(n10869), .ZN(n10863) );
  NAND2_X1 U13408 ( .A1(n10863), .A2(n14465), .ZN(n10864) );
  NOR2_X1 U13409 ( .A1(n10986), .A2(n10864), .ZN(n11022) );
  XNOR2_X1 U13410 ( .A(n10865), .B(n10866), .ZN(n10868) );
  OAI21_X1 U13411 ( .B1(n10868), .B2(n13340), .A(n10867), .ZN(n11016) );
  AOI211_X1 U13412 ( .C1(n14479), .C2(n11015), .A(n11022), .B(n11016), .ZN(
        n10875) );
  INV_X1 U13413 ( .A(n10869), .ZN(n11020) );
  OAI22_X1 U13414 ( .A1(n13418), .A2(n11020), .B1(n15105), .B2(n10870), .ZN(
        n10871) );
  INV_X1 U13415 ( .A(n10871), .ZN(n10872) );
  OAI21_X1 U13416 ( .B1(n10875), .B2(n15103), .A(n10872), .ZN(P2_U3505) );
  OAI22_X1 U13417 ( .A1(n13468), .A2(n11020), .B1(n15099), .B2(n7683), .ZN(
        n10873) );
  INV_X1 U13418 ( .A(n10873), .ZN(n10874) );
  OAI21_X1 U13419 ( .B1(n10875), .B2(n15098), .A(n10874), .ZN(P2_U3448) );
  OAI22_X1 U13420 ( .A1(n12293), .A2(n12819), .B1(n10876), .B2(n12298), .ZN(
        n10877) );
  AOI21_X1 U13421 ( .B1(n12291), .B2(n12817), .A(n10877), .ZN(n10883) );
  INV_X1 U13422 ( .A(n12822), .ZN(n10878) );
  NAND3_X1 U13423 ( .A1(n10878), .A2(n12823), .A3(n12200), .ZN(n10879) );
  NAND2_X1 U13424 ( .A1(n10881), .A2(n12269), .ZN(n10882) );
  OAI211_X1 U13425 ( .C1(n10891), .C2(n12828), .A(n10883), .B(n10882), .ZN(
        P3_U3162) );
  OAI21_X1 U13426 ( .B1(n10886), .B2(n10885), .A(n10884), .ZN(n10887) );
  NAND2_X1 U13427 ( .A1(n10887), .A2(n12269), .ZN(n10890) );
  OAI22_X1 U13428 ( .A1(n12293), .A2(n15293), .B1(n12298), .B2(n15310), .ZN(
        n10888) );
  AOI21_X1 U13429 ( .B1(n12291), .B2(n10491), .A(n10888), .ZN(n10889) );
  OAI211_X1 U13430 ( .C1(n10891), .C2(n15311), .A(n10890), .B(n10889), .ZN(
        P3_U3177) );
  INV_X1 U13431 ( .A(n13961), .ZN(n13957) );
  INV_X1 U13432 ( .A(n10892), .ZN(n10895) );
  OAI222_X1 U13433 ( .A1(P1_U3086), .A2(n13957), .B1(n14304), .B2(n10895), 
        .C1(n10893), .C2(n14298), .ZN(P1_U3338) );
  INV_X1 U13434 ( .A(n15027), .ZN(n10894) );
  OAI222_X1 U13435 ( .A1(n13776), .A2(n13735), .B1(n11134), .B2(n10895), .C1(
        n10894), .C2(P2_U3088), .ZN(P2_U3310) );
  OR2_X1 U13436 ( .A1(n10896), .A2(n10901), .ZN(n10897) );
  NAND2_X1 U13437 ( .A1(n10898), .A2(n10897), .ZN(n11248) );
  AOI21_X1 U13438 ( .B1(n11038), .B2(n11242), .A(n9935), .ZN(n10900) );
  NAND2_X1 U13439 ( .A1(n10900), .A2(n10899), .ZN(n11244) );
  INV_X1 U13440 ( .A(n11244), .ZN(n10906) );
  XNOR2_X1 U13441 ( .A(n10902), .B(n10901), .ZN(n10905) );
  NAND2_X1 U13442 ( .A1(n11248), .A2(n13333), .ZN(n10904) );
  AOI22_X1 U13443 ( .A1(n13335), .A2(n13083), .B1(n13081), .B2(n13336), .ZN(
        n10903) );
  OAI211_X1 U13444 ( .C1(n10905), .C2(n13340), .A(n10904), .B(n10903), .ZN(
        n11245) );
  AOI211_X1 U13445 ( .C1(n15097), .C2(n11248), .A(n10906), .B(n11245), .ZN(
        n10912) );
  OAI22_X1 U13446 ( .A1(n13418), .A2(n7085), .B1(n15105), .B2(n10907), .ZN(
        n10908) );
  INV_X1 U13447 ( .A(n10908), .ZN(n10909) );
  OAI21_X1 U13448 ( .B1(n10912), .B2(n15103), .A(n10909), .ZN(P2_U3504) );
  OAI22_X1 U13449 ( .A1(n13468), .A2(n7085), .B1(n15099), .B2(n7648), .ZN(
        n10910) );
  INV_X1 U13450 ( .A(n10910), .ZN(n10911) );
  OAI21_X1 U13451 ( .B1(n10912), .B2(n15098), .A(n10911), .ZN(P2_U3445) );
  INV_X1 U13452 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n10914) );
  NAND2_X1 U13453 ( .A1(n12702), .A2(P3_U3897), .ZN(n10913) );
  OAI21_X1 U13454 ( .B1(P3_U3897), .B2(n10914), .A(n10913), .ZN(P3_U3515) );
  AOI21_X1 U13455 ( .B1(n6575), .B2(n14765), .A(n14743), .ZN(n10919) );
  INV_X1 U13456 ( .A(n14177), .ZN(n14557) );
  NOR2_X1 U13457 ( .A1(n10781), .A2(n14557), .ZN(n14764) );
  INV_X1 U13458 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n13899) );
  OAI22_X1 U13459 ( .A1(n14741), .A2(n13899), .B1(n10915), .B2(n14739), .ZN(
        n10916) );
  AOI21_X1 U13460 ( .B1(n14764), .B2(n14741), .A(n10916), .ZN(n10918) );
  OAI21_X1 U13461 ( .B1(n14571), .B2(n14570), .A(n14761), .ZN(n10917) );
  OAI211_X1 U13462 ( .C1(n10919), .C2(n10953), .A(n10918), .B(n10917), .ZN(
        P1_U3293) );
  XNOR2_X1 U13463 ( .A(n10920), .B(n12480), .ZN(n15346) );
  INV_X1 U13464 ( .A(n15346), .ZN(n10932) );
  NAND2_X1 U13465 ( .A1(n15330), .A2(n15329), .ZN(n12698) );
  AOI21_X1 U13466 ( .B1(n10921), .B2(n12480), .A(n15299), .ZN(n10924) );
  OAI22_X1 U13467 ( .A1(n10841), .A2(n15294), .B1(n12819), .B2(n15292), .ZN(
        n10922) );
  AOI21_X1 U13468 ( .B1(n10924), .B2(n10923), .A(n10922), .ZN(n10926) );
  NAND2_X1 U13469 ( .A1(n15346), .A2(n15297), .ZN(n10925) );
  AND2_X1 U13470 ( .A1(n10926), .A2(n10925), .ZN(n15343) );
  MUX2_X1 U13471 ( .A(n10927), .B(n15343), .S(n15330), .Z(n10931) );
  NOR2_X1 U13472 ( .A1(n10928), .A2(n15368), .ZN(n15345) );
  AOI22_X1 U13473 ( .A1(n15305), .A2(n15345), .B1(n15253), .B2(n10929), .ZN(
        n10930) );
  OAI211_X1 U13474 ( .C1(n10932), .C2(n12698), .A(n10931), .B(n10930), .ZN(
        P3_U3230) );
  INV_X1 U13475 ( .A(SI_21_), .ZN(n10933) );
  OAI222_X1 U13476 ( .A1(n12961), .A2(n10934), .B1(n12962), .B2(n10933), .C1(
        P3_U3151), .C2(n10819), .ZN(P3_U3274) );
  XNOR2_X1 U13477 ( .A(n10936), .B(n10935), .ZN(n14778) );
  NAND2_X1 U13478 ( .A1(n14778), .A2(n14719), .ZN(n10945) );
  OAI21_X1 U13479 ( .B1(n10941), .B2(n10940), .A(n10939), .ZN(n10943) );
  AOI21_X1 U13480 ( .B1(n10943), .B2(n14738), .A(n10942), .ZN(n10944) );
  AND2_X1 U13481 ( .A1(n10945), .A2(n10944), .ZN(n14780) );
  OR2_X1 U13482 ( .A1(n14157), .A2(n10946), .ZN(n14071) );
  INV_X1 U13483 ( .A(n14071), .ZN(n14748) );
  OAI211_X1 U13484 ( .C1(n10955), .C2(n14776), .A(n14725), .B(n14746), .ZN(
        n14775) );
  INV_X1 U13485 ( .A(n14775), .ZN(n10947) );
  NAND2_X1 U13486 ( .A1(n6575), .A2(n10947), .ZN(n10949) );
  INV_X1 U13487 ( .A(n14739), .ZN(n14722) );
  AOI22_X1 U13488 ( .A1(n14157), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n14722), .ZN(n10948) );
  OAI211_X1 U13489 ( .C1(n14776), .C2(n14337), .A(n10949), .B(n10948), .ZN(
        n10950) );
  AOI21_X1 U13490 ( .B1(n14748), .B2(n14778), .A(n10950), .ZN(n10951) );
  OAI21_X1 U13491 ( .B1(n14157), .B2(n14780), .A(n10951), .ZN(P1_U3291) );
  XNOR2_X1 U13492 ( .A(n10958), .B(n10952), .ZN(n14774) );
  NOR2_X1 U13493 ( .A1(n14770), .A2(n10953), .ZN(n10954) );
  NOR2_X1 U13494 ( .A1(n10955), .A2(n10954), .ZN(n10959) );
  AND2_X1 U13495 ( .A1(n10959), .A2(n14725), .ZN(n14767) );
  NAND2_X1 U13496 ( .A1(n6575), .A2(n14767), .ZN(n10957) );
  AOI22_X1 U13497 ( .A1(n14157), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n14722), .ZN(n10956) );
  OAI211_X1 U13498 ( .C1(n14770), .C2(n14337), .A(n10957), .B(n10956), .ZN(
        n10966) );
  OAI21_X1 U13499 ( .B1(n10958), .B2(n8320), .A(n14738), .ZN(n10963) );
  XNOR2_X1 U13500 ( .A(n10959), .B(n10781), .ZN(n10961) );
  AOI21_X1 U13501 ( .B1(n10961), .B2(n14738), .A(n10960), .ZN(n10962) );
  AOI21_X1 U13502 ( .B1(n14555), .B2(n10963), .A(n10962), .ZN(n10964) );
  AOI21_X1 U13503 ( .B1(n14719), .B2(n14774), .A(n10964), .ZN(n14771) );
  NAND2_X1 U13504 ( .A1(n13898), .A2(n14177), .ZN(n14768) );
  AOI21_X1 U13505 ( .B1(n14771), .B2(n14768), .A(n14157), .ZN(n10965) );
  AOI211_X1 U13506 ( .C1(n14748), .C2(n14774), .A(n10966), .B(n10965), .ZN(
        n10967) );
  INV_X1 U13507 ( .A(n10967), .ZN(P1_U3292) );
  OAI21_X1 U13508 ( .B1(n10970), .B2(n10969), .A(n10968), .ZN(n10977) );
  INV_X1 U13509 ( .A(n11052), .ZN(n11162) );
  NOR2_X1 U13510 ( .A1(n13017), .A2(n11162), .ZN(n10976) );
  NAND2_X1 U13511 ( .A1(n13080), .A2(n13335), .ZN(n10972) );
  NAND2_X1 U13512 ( .A1(n13078), .A2(n13336), .ZN(n10971) );
  AND2_X1 U13513 ( .A1(n10972), .A2(n10971), .ZN(n11049) );
  INV_X1 U13514 ( .A(n11049), .ZN(n10973) );
  NAND2_X1 U13515 ( .A1(n14450), .A2(n10973), .ZN(n10974) );
  NAND2_X1 U13516 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n14938) );
  OAI211_X1 U13517 ( .C1(n14453), .C2(n11055), .A(n10974), .B(n14938), .ZN(
        n10975) );
  AOI211_X1 U13518 ( .C1(n10977), .C2(n14448), .A(n10976), .B(n10975), .ZN(
        n10978) );
  INV_X1 U13519 ( .A(n10978), .ZN(P2_U3193) );
  OAI21_X1 U13520 ( .B1(n10981), .B2(n10980), .A(n10979), .ZN(n15064) );
  INV_X1 U13521 ( .A(n15064), .ZN(n10987) );
  XNOR2_X1 U13522 ( .A(n10983), .B(n10982), .ZN(n10985) );
  AOI21_X1 U13523 ( .B1(n10985), .B2(n14456), .A(n10984), .ZN(n15066) );
  OAI211_X1 U13524 ( .C1(n10986), .C2(n10990), .A(n11053), .B(n14465), .ZN(
        n15060) );
  OAI211_X1 U13525 ( .C1(n10987), .C2(n13440), .A(n15066), .B(n15060), .ZN(
        n10992) );
  OAI22_X1 U13526 ( .A1(n13418), .A2(n10990), .B1(n15105), .B2(n7704), .ZN(
        n10988) );
  AOI21_X1 U13527 ( .B1(n10992), .B2(n15105), .A(n10988), .ZN(n10989) );
  INV_X1 U13528 ( .A(n10989), .ZN(P2_U3506) );
  INV_X1 U13529 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n13598) );
  OAI22_X1 U13530 ( .A1(n13468), .A2(n10990), .B1(n15099), .B2(n13598), .ZN(
        n10991) );
  AOI21_X1 U13531 ( .B1(n10992), .B2(n15099), .A(n10991), .ZN(n10993) );
  INV_X1 U13532 ( .A(n10993), .ZN(P2_U3451) );
  XNOR2_X1 U13533 ( .A(n11000), .B(n12200), .ZN(n11137) );
  XNOR2_X1 U13534 ( .A(n11137), .B(n15276), .ZN(n10997) );
  OAI21_X1 U13535 ( .B1(n10997), .B2(n10996), .A(n11139), .ZN(n10998) );
  NAND2_X1 U13536 ( .A1(n10998), .A2(n12269), .ZN(n11004) );
  AOI21_X1 U13537 ( .B1(n12282), .B2(n11000), .A(n10999), .ZN(n11001) );
  OAI21_X1 U13538 ( .B1(n12293), .B2(n15260), .A(n11001), .ZN(n11002) );
  AOI21_X1 U13539 ( .B1(n12291), .B2(n12524), .A(n11002), .ZN(n11003) );
  OAI211_X1 U13540 ( .C1(n11234), .C2(n12178), .A(n11004), .B(n11003), .ZN(
        P3_U3167) );
  AOI21_X1 U13541 ( .B1(n14467), .B2(n11005), .A(n15058), .ZN(n11013) );
  OAI22_X1 U13542 ( .A1(n13358), .A2(n11007), .B1(n11006), .B2(n15052), .ZN(
        n11008) );
  AOI21_X1 U13543 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n13358), .A(n11008), .ZN(
        n11011) );
  INV_X1 U13544 ( .A(n13348), .ZN(n11858) );
  NAND2_X1 U13545 ( .A1(n11858), .A2(n11009), .ZN(n11010) );
  OAI211_X1 U13546 ( .C1(n11013), .C2(n11012), .A(n11011), .B(n11010), .ZN(
        P2_U3265) );
  AND2_X1 U13547 ( .A1(n8198), .A2(n11192), .ZN(n11014) );
  INV_X1 U13548 ( .A(n11015), .ZN(n11025) );
  INV_X1 U13549 ( .A(n11016), .ZN(n11017) );
  MUX2_X1 U13550 ( .A(n11018), .B(n11017), .S(n15055), .Z(n11024) );
  OAI22_X1 U13551 ( .A1(n13360), .A2(n11020), .B1(n15052), .B2(n11019), .ZN(
        n11021) );
  AOI21_X1 U13552 ( .B1(n14467), .B2(n11022), .A(n11021), .ZN(n11023) );
  OAI211_X1 U13553 ( .C1(n13365), .C2(n11025), .A(n11024), .B(n11023), .ZN(
        P2_U3259) );
  OR2_X1 U13554 ( .A1(n11027), .A2(n11026), .ZN(n11028) );
  NAND2_X1 U13555 ( .A1(n11029), .A2(n11028), .ZN(n15089) );
  INV_X1 U13556 ( .A(n15089), .ZN(n11043) );
  NAND2_X1 U13557 ( .A1(n15089), .A2(n13333), .ZN(n11036) );
  OAI21_X1 U13558 ( .B1(n11032), .B2(n11031), .A(n11030), .ZN(n11033) );
  NAND2_X1 U13559 ( .A1(n11033), .A2(n14456), .ZN(n11035) );
  AOI22_X1 U13560 ( .A1(n13335), .A2(n13084), .B1(n13082), .B2(n13336), .ZN(
        n11034) );
  NAND3_X1 U13561 ( .A1(n11036), .A2(n11035), .A3(n11034), .ZN(n15087) );
  MUX2_X1 U13562 ( .A(n15087), .B(P2_REG2_REG_4__SCAN_IN), .S(n13358), .Z(
        n11037) );
  INV_X1 U13563 ( .A(n11037), .ZN(n11042) );
  AOI211_X1 U13564 ( .C1(n13022), .C2(n11039), .A(n9935), .B(n7086), .ZN(
        n15084) );
  OAI22_X1 U13565 ( .A1(n13360), .A2(n15086), .B1(n15052), .B2(n13024), .ZN(
        n11040) );
  AOI21_X1 U13566 ( .B1(n14467), .B2(n15084), .A(n11040), .ZN(n11041) );
  OAI211_X1 U13567 ( .C1(n11043), .C2(n13348), .A(n11042), .B(n11041), .ZN(
        P2_U3261) );
  OAI21_X1 U13568 ( .B1(n7534), .B2(n11045), .A(n11044), .ZN(n11158) );
  OAI211_X1 U13569 ( .C1(n11048), .C2(n11047), .A(n11046), .B(n14456), .ZN(
        n11050) );
  AND2_X1 U13570 ( .A1(n11050), .A2(n11049), .ZN(n11157) );
  MUX2_X1 U13571 ( .A(n11051), .B(n11157), .S(n15055), .Z(n11059) );
  AOI21_X1 U13572 ( .B1(n11053), .B2(n11052), .A(n9935), .ZN(n11054) );
  NAND2_X1 U13573 ( .A1(n11054), .A2(n11216), .ZN(n11156) );
  INV_X1 U13574 ( .A(n11156), .ZN(n11057) );
  OAI22_X1 U13575 ( .A1(n13360), .A2(n11162), .B1(n15052), .B2(n11055), .ZN(
        n11056) );
  AOI21_X1 U13576 ( .B1(n11057), .B2(n14467), .A(n11056), .ZN(n11058) );
  OAI211_X1 U13577 ( .C1(n13365), .C2(n11158), .A(n11059), .B(n11058), .ZN(
        P2_U3257) );
  INV_X1 U13578 ( .A(n11060), .ZN(n11062) );
  OAI22_X1 U13579 ( .A1(n12509), .A2(P3_U3151), .B1(SI_22_), .B2(n12962), .ZN(
        n11061) );
  AOI21_X1 U13580 ( .B1(n11062), .B2(n14325), .A(n11061), .ZN(P3_U3273) );
  INV_X1 U13581 ( .A(n11339), .ZN(n11222) );
  OAI21_X1 U13582 ( .B1(n11065), .B2(n11064), .A(n11063), .ZN(n11066) );
  NAND2_X1 U13583 ( .A1(n11066), .A2(n14448), .ZN(n11070) );
  INV_X1 U13584 ( .A(n11219), .ZN(n11068) );
  AOI22_X1 U13585 ( .A1(n13335), .A2(n13079), .B1(n13077), .B2(n13336), .ZN(
        n11214) );
  NAND2_X1 U13586 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14952) );
  OAI21_X1 U13587 ( .B1(n13012), .B2(n11214), .A(n14952), .ZN(n11067) );
  AOI21_X1 U13588 ( .B1(n11068), .B2(n13014), .A(n11067), .ZN(n11069) );
  OAI211_X1 U13589 ( .C1(n11222), .C2(n13017), .A(n11070), .B(n11069), .ZN(
        P2_U3203) );
  OAI21_X1 U13590 ( .B1(n11073), .B2(n11072), .A(n11071), .ZN(n15083) );
  INV_X1 U13591 ( .A(n15083), .ZN(n11087) );
  OAI21_X1 U13592 ( .B1(n11076), .B2(n11075), .A(n6576), .ZN(n11079) );
  OAI22_X1 U13593 ( .A1(n11077), .A2(n14443), .B1(n6745), .B2(n14441), .ZN(
        n11078) );
  AOI21_X1 U13594 ( .B1(n11079), .B2(n14456), .A(n11078), .ZN(n11080) );
  OAI21_X1 U13595 ( .B1(n11087), .B2(n8198), .A(n11080), .ZN(n15081) );
  INV_X1 U13596 ( .A(n15052), .ZN(n14460) );
  AOI22_X1 U13597 ( .A1(n13358), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n14460), .ZN(n11081) );
  OAI21_X1 U13598 ( .B1(n13360), .B2(n15080), .A(n11081), .ZN(n11089) );
  NAND2_X1 U13599 ( .A1(n11083), .A2(n11082), .ZN(n11084) );
  NAND2_X1 U13600 ( .A1(n11084), .A2(n14465), .ZN(n11085) );
  OR2_X1 U13601 ( .A1(n11086), .A2(n11085), .ZN(n15079) );
  OAI22_X1 U13602 ( .A1(n11087), .A2(n13348), .B1(n15061), .B2(n15079), .ZN(
        n11088) );
  AOI211_X1 U13603 ( .C1(n15055), .C2(n15081), .A(n11089), .B(n11088), .ZN(
        n11090) );
  INV_X1 U13604 ( .A(n11090), .ZN(P2_U3263) );
  OR2_X1 U13605 ( .A1(n13896), .A2(n11091), .ZN(n11092) );
  NAND2_X1 U13606 ( .A1(n11093), .A2(n11092), .ZN(n14715) );
  INV_X1 U13607 ( .A(n14723), .ZN(n14796) );
  NAND2_X1 U13608 ( .A1(n14796), .A2(n13895), .ZN(n11094) );
  OR2_X1 U13609 ( .A1(n13895), .A2(n14796), .ZN(n11095) );
  INV_X1 U13610 ( .A(n13894), .ZN(n11097) );
  OR2_X1 U13611 ( .A1(n13872), .A2(n11097), .ZN(n11098) );
  NAND2_X1 U13612 ( .A1(n11121), .A2(n11098), .ZN(n11271) );
  INV_X1 U13613 ( .A(n11390), .ZN(n14811) );
  XNOR2_X1 U13614 ( .A(n11314), .B(n11326), .ZN(n11101) );
  NAND2_X1 U13615 ( .A1(n13893), .A2(n14178), .ZN(n11099) );
  OAI21_X1 U13616 ( .B1(n11598), .B2(n14557), .A(n11099), .ZN(n11100) );
  AOI21_X1 U13617 ( .B1(n11101), .B2(n14738), .A(n11100), .ZN(n14821) );
  INV_X1 U13618 ( .A(n11102), .ZN(n11103) );
  NAND2_X1 U13619 ( .A1(n11104), .A2(n11103), .ZN(n11106) );
  OR2_X1 U13620 ( .A1(n13896), .A2(n14789), .ZN(n11105) );
  NAND2_X1 U13621 ( .A1(n11106), .A2(n11105), .ZN(n14713) );
  NAND2_X1 U13622 ( .A1(n14713), .A2(n14714), .ZN(n11109) );
  OR2_X1 U13623 ( .A1(n13895), .A2(n14723), .ZN(n11108) );
  OR2_X1 U13624 ( .A1(n13872), .A2(n13894), .ZN(n11110) );
  OR2_X1 U13625 ( .A1(n11390), .A2(n13893), .ZN(n11111) );
  NAND2_X1 U13626 ( .A1(n11112), .A2(n11111), .ZN(n11327) );
  XNOR2_X1 U13627 ( .A(n11327), .B(n11326), .ZN(n14819) );
  INV_X1 U13628 ( .A(n11506), .ZN(n14817) );
  NAND2_X1 U13629 ( .A1(n11265), .A2(n14817), .ZN(n14707) );
  OAI211_X1 U13630 ( .C1(n11265), .C2(n14817), .A(n14725), .B(n14707), .ZN(
        n14816) );
  OAI22_X1 U13631 ( .A1(n14741), .A2(n8445), .B1(n11518), .B2(n14739), .ZN(
        n11113) );
  AOI21_X1 U13632 ( .B1(n14743), .B2(n11506), .A(n11113), .ZN(n11114) );
  OAI21_X1 U13633 ( .B1(n14816), .B2(n14186), .A(n11114), .ZN(n11115) );
  AOI21_X1 U13634 ( .B1(n14819), .B2(n14570), .A(n11115), .ZN(n11116) );
  OAI21_X1 U13635 ( .B1(n14821), .B2(n14157), .A(n11116), .ZN(P1_U3285) );
  INV_X1 U13636 ( .A(n14806), .ZN(n11130) );
  AOI21_X1 U13637 ( .B1(n11118), .B2(n11117), .A(n14837), .ZN(n11122) );
  NAND2_X1 U13638 ( .A1(n13895), .A2(n14178), .ZN(n11120) );
  NAND2_X1 U13639 ( .A1(n13893), .A2(n14177), .ZN(n11119) );
  NAND2_X1 U13640 ( .A1(n11120), .A2(n11119), .ZN(n13871) );
  AOI21_X1 U13641 ( .B1(n11122), .B2(n11121), .A(n13871), .ZN(n11124) );
  NAND2_X1 U13642 ( .A1(n14806), .A2(n14719), .ZN(n11123) );
  AND2_X1 U13643 ( .A1(n11124), .A2(n11123), .ZN(n14808) );
  MUX2_X1 U13644 ( .A(n14808), .B(n11125), .S(n14157), .Z(n11129) );
  AOI21_X1 U13645 ( .B1(n14724), .B2(n13872), .A(n14745), .ZN(n11126) );
  AND2_X1 U13646 ( .A1(n11266), .A2(n11126), .ZN(n14802) );
  INV_X1 U13647 ( .A(n13872), .ZN(n14804) );
  OAI22_X1 U13648 ( .A1(n14337), .A2(n14804), .B1(n13873), .B2(n14739), .ZN(
        n11127) );
  AOI21_X1 U13649 ( .B1(n14802), .B2(n6575), .A(n11127), .ZN(n11128) );
  OAI211_X1 U13650 ( .C1(n11130), .C2(n14071), .A(n11129), .B(n11128), .ZN(
        P1_U3287) );
  INV_X1 U13651 ( .A(n13976), .ZN(n13969) );
  INV_X1 U13652 ( .A(n11131), .ZN(n11133) );
  OAI222_X1 U13653 ( .A1(P1_U3086), .A2(n13969), .B1(n14304), .B2(n11133), 
        .C1(n11132), .C2(n14298), .ZN(P1_U3337) );
  OAI222_X1 U13654 ( .A1(n13776), .A2(n11135), .B1(n11134), .B2(n11133), .C1(
        n15045), .C2(P2_U3088), .ZN(P2_U3309) );
  NAND2_X1 U13655 ( .A1(n12526), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11136) );
  OAI21_X1 U13656 ( .B1(n12205), .B2(n12526), .A(n11136), .ZN(P3_U3520) );
  NAND2_X1 U13657 ( .A1(n11137), .A2(n15295), .ZN(n11138) );
  XNOR2_X1 U13658 ( .A(n15281), .B(n12200), .ZN(n11198) );
  XNOR2_X1 U13659 ( .A(n11198), .B(n15260), .ZN(n11141) );
  AOI21_X1 U13660 ( .B1(n11140), .B2(n11141), .A(n12285), .ZN(n11143) );
  INV_X1 U13661 ( .A(n11141), .ZN(n11142) );
  NAND2_X1 U13662 ( .A1(n11143), .A2(n11201), .ZN(n11148) );
  AOI21_X1 U13663 ( .B1(n12282), .B2(n15281), .A(n11144), .ZN(n11145) );
  OAI21_X1 U13664 ( .B1(n12293), .B2(n11309), .A(n11145), .ZN(n11146) );
  AOI21_X1 U13665 ( .B1(n12291), .B2(n15276), .A(n11146), .ZN(n11147) );
  OAI211_X1 U13666 ( .C1(n15282), .C2(n12178), .A(n11148), .B(n11147), .ZN(
        P3_U3179) );
  NAND2_X1 U13667 ( .A1(n12526), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n11149) );
  OAI21_X1 U13668 ( .B1(n12466), .B2(n12526), .A(n11149), .ZN(P3_U3521) );
  XNOR2_X1 U13669 ( .A(n11151), .B(n11150), .ZN(n11155) );
  NAND2_X1 U13670 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n14965)
         );
  OAI21_X1 U13671 ( .B1(n14453), .B2(n11350), .A(n14965), .ZN(n11153) );
  OAI22_X1 U13672 ( .A1(n11346), .A2(n13045), .B1(n13044), .B2(n11383), .ZN(
        n11152) );
  AOI211_X1 U13673 ( .C1(n11356), .C2(n14451), .A(n11153), .B(n11152), .ZN(
        n11154) );
  OAI21_X1 U13674 ( .B1(n11155), .B2(n13059), .A(n11154), .ZN(P2_U3189) );
  OAI211_X1 U13675 ( .C1(n11158), .C2(n13440), .A(n11157), .B(n11156), .ZN(
        n11164) );
  OAI22_X1 U13676 ( .A1(n11162), .A2(n13418), .B1(n15105), .B2(n11159), .ZN(
        n11160) );
  AOI21_X1 U13677 ( .B1(n11164), .B2(n15105), .A(n11160), .ZN(n11161) );
  INV_X1 U13678 ( .A(n11161), .ZN(P2_U3507) );
  OAI22_X1 U13679 ( .A1(n13468), .A2(n11162), .B1(n15099), .B2(n7723), .ZN(
        n11163) );
  AOI21_X1 U13680 ( .B1(n11164), .B2(n15099), .A(n11163), .ZN(n11165) );
  INV_X1 U13681 ( .A(n11165), .ZN(P2_U3454) );
  INV_X1 U13682 ( .A(n11166), .ZN(n11168) );
  AOI22_X1 U13683 ( .A1(n13896), .A2(n12077), .B1(n12064), .B2(n14789), .ZN(
        n11171) );
  AOI22_X1 U13684 ( .A1(n13896), .A2(n6578), .B1(n12079), .B2(n14789), .ZN(
        n11170) );
  XOR2_X1 U13685 ( .A(n11786), .B(n11170), .Z(n11255) );
  INV_X1 U13686 ( .A(n11171), .ZN(n11172) );
  NAND2_X1 U13687 ( .A1(n13895), .A2(n6577), .ZN(n11176) );
  NAND2_X1 U13688 ( .A1(n14723), .A2(n12079), .ZN(n11175) );
  NAND2_X1 U13689 ( .A1(n11176), .A2(n11175), .ZN(n11177) );
  XNOR2_X1 U13690 ( .A(n11177), .B(n11974), .ZN(n11181) );
  NAND2_X1 U13691 ( .A1(n13895), .A2(n12077), .ZN(n11179) );
  NAND2_X1 U13692 ( .A1(n14723), .A2(n12064), .ZN(n11178) );
  NAND2_X1 U13693 ( .A1(n11179), .A2(n11178), .ZN(n11180) );
  NAND2_X1 U13694 ( .A1(n11181), .A2(n11180), .ZN(n11392) );
  NAND2_X1 U13695 ( .A1(n6724), .A2(n11392), .ZN(n11182) );
  XNOR2_X1 U13696 ( .A(n11393), .B(n11182), .ZN(n11189) );
  NAND2_X1 U13697 ( .A1(n13896), .A2(n14178), .ZN(n11184) );
  NAND2_X1 U13698 ( .A1(n13894), .A2(n14177), .ZN(n11183) );
  NAND2_X1 U13699 ( .A1(n11184), .A2(n11183), .ZN(n14718) );
  NAND2_X1 U13700 ( .A1(n14517), .A2(n14718), .ZN(n11185) );
  OAI211_X1 U13701 ( .C1(n14554), .C2(n14720), .A(n11186), .B(n11185), .ZN(
        n11187) );
  AOI21_X1 U13702 ( .B1(n14723), .B2(n14536), .A(n11187), .ZN(n11188) );
  OAI21_X1 U13703 ( .B1(n11189), .B2(n14532), .A(n11188), .ZN(P1_U3227) );
  NAND2_X1 U13704 ( .A1(n12526), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n11190) );
  OAI21_X1 U13705 ( .B1(n12637), .B2(n12526), .A(n11190), .ZN(P3_U3519) );
  INV_X1 U13706 ( .A(n11191), .ZN(n11194) );
  OAI222_X1 U13707 ( .A1(n13776), .A2(n11193), .B1(n11134), .B2(n11194), .C1(
        n11192), .C2(P2_U3088), .ZN(P2_U3308) );
  OAI222_X1 U13708 ( .A1(P1_U3086), .A2(n13984), .B1(n14304), .B2(n11194), 
        .C1(n13560), .C2(n14298), .ZN(P1_U3336) );
  INV_X1 U13709 ( .A(SI_23_), .ZN(n11197) );
  NAND2_X1 U13710 ( .A1(n11195), .A2(n14325), .ZN(n11196) );
  OAI211_X1 U13711 ( .C1(n11197), .C2(n12962), .A(n11196), .B(n12512), .ZN(
        P3_U3272) );
  INV_X1 U13712 ( .A(n11198), .ZN(n11199) );
  NAND2_X1 U13713 ( .A1(n12523), .A2(n11199), .ZN(n11200) );
  XNOR2_X1 U13714 ( .A(n11203), .B(n12157), .ZN(n11304) );
  XNOR2_X1 U13715 ( .A(n11304), .B(n11309), .ZN(n11302) );
  XNOR2_X1 U13716 ( .A(n11303), .B(n11302), .ZN(n11208) );
  AOI21_X1 U13717 ( .B1(n12282), .B2(n11203), .A(n11202), .ZN(n11204) );
  OAI21_X1 U13718 ( .B1(n12293), .B2(n15259), .A(n11204), .ZN(n11206) );
  NOR2_X1 U13719 ( .A1(n12178), .A2(n15261), .ZN(n11205) );
  AOI211_X1 U13720 ( .C1(n12291), .C2(n12523), .A(n11206), .B(n11205), .ZN(
        n11207) );
  OAI21_X1 U13721 ( .B1(n11208), .B2(n12285), .A(n11207), .ZN(P3_U3153) );
  XOR2_X1 U13722 ( .A(n11209), .B(n11213), .Z(n11335) );
  INV_X1 U13723 ( .A(n11335), .ZN(n11226) );
  INV_X1 U13724 ( .A(n11210), .ZN(n11211) );
  AOI21_X1 U13725 ( .B1(n11213), .B2(n11212), .A(n11211), .ZN(n11215) );
  OAI21_X1 U13726 ( .B1(n11215), .B2(n13340), .A(n11214), .ZN(n11333) );
  NAND2_X1 U13727 ( .A1(n11333), .A2(n15055), .ZN(n11225) );
  NAND2_X1 U13728 ( .A1(n11216), .A2(n11339), .ZN(n11217) );
  NAND2_X1 U13729 ( .A1(n11217), .A2(n14465), .ZN(n11218) );
  NOR2_X1 U13730 ( .A1(n11353), .A2(n11218), .ZN(n11334) );
  NOR2_X1 U13731 ( .A1(n15052), .A2(n11219), .ZN(n11220) );
  AOI21_X1 U13732 ( .B1(n13358), .B2(P2_REG2_REG_9__SCAN_IN), .A(n11220), .ZN(
        n11221) );
  OAI21_X1 U13733 ( .B1(n13360), .B2(n11222), .A(n11221), .ZN(n11223) );
  AOI21_X1 U13734 ( .B1(n11334), .B2(n14467), .A(n11223), .ZN(n11224) );
  OAI211_X1 U13735 ( .C1(n13365), .C2(n11226), .A(n11225), .B(n11224), .ZN(
        P2_U3256) );
  XNOR2_X1 U13736 ( .A(n11228), .B(n9323), .ZN(n15352) );
  OAI21_X1 U13737 ( .B1(n11230), .B2(n9323), .A(n11229), .ZN(n11232) );
  OAI22_X1 U13738 ( .A1(n10841), .A2(n15292), .B1(n15260), .B2(n15294), .ZN(
        n11231) );
  AOI21_X1 U13739 ( .B1(n11232), .B2(n15319), .A(n11231), .ZN(n11233) );
  OAI21_X1 U13740 ( .B1(n15327), .B2(n15352), .A(n11233), .ZN(n15353) );
  NAND2_X1 U13741 ( .A1(n15353), .A2(n15330), .ZN(n11239) );
  NOR2_X1 U13742 ( .A1(n12360), .A2(n15368), .ZN(n15354) );
  INV_X1 U13743 ( .A(n15354), .ZN(n11235) );
  OAI22_X1 U13744 ( .A1(n11236), .A2(n11235), .B1(n11234), .B2(n15312), .ZN(
        n11237) );
  AOI21_X1 U13745 ( .B1(n15333), .B2(P3_REG2_REG_5__SCAN_IN), .A(n11237), .ZN(
        n11238) );
  OAI211_X1 U13746 ( .C1(n15352), .C2(n12698), .A(n11239), .B(n11238), .ZN(
        P3_U3228) );
  INV_X1 U13747 ( .A(n11240), .ZN(n11241) );
  AOI22_X1 U13748 ( .A1(n15058), .A2(n11242), .B1(n14460), .B2(n11241), .ZN(
        n11243) );
  OAI21_X1 U13749 ( .B1(n15061), .B2(n11244), .A(n11243), .ZN(n11247) );
  MUX2_X1 U13750 ( .A(n11245), .B(P2_REG2_REG_5__SCAN_IN), .S(n13358), .Z(
        n11246) );
  AOI211_X1 U13751 ( .C1(n11858), .C2(n11248), .A(n11247), .B(n11246), .ZN(
        n11249) );
  INV_X1 U13752 ( .A(n11249), .ZN(P2_U3260) );
  NAND2_X1 U13753 ( .A1(n14545), .A2(n13897), .ZN(n11253) );
  NAND2_X1 U13754 ( .A1(n14547), .A2(n13895), .ZN(n11252) );
  NAND2_X1 U13755 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n14678) );
  OR2_X1 U13756 ( .A1(n14554), .A2(n11250), .ZN(n11251) );
  NAND4_X1 U13757 ( .A1(n11253), .A2(n11252), .A3(n14678), .A4(n11251), .ZN(
        n11258) );
  XNOR2_X1 U13758 ( .A(n11254), .B(n11255), .ZN(n11256) );
  NOR2_X1 U13759 ( .A1(n11256), .A2(n14532), .ZN(n11257) );
  AOI211_X1 U13760 ( .C1(n14789), .C2(n14536), .A(n11258), .B(n11257), .ZN(
        n11259) );
  INV_X1 U13761 ( .A(n11259), .ZN(P1_U3230) );
  INV_X1 U13762 ( .A(n11260), .ZN(n11263) );
  OAI222_X1 U13763 ( .A1(P1_U3086), .A2(n11261), .B1(n14304), .B2(n11263), 
        .C1(n7027), .C2(n14298), .ZN(P1_U3335) );
  OAI222_X1 U13764 ( .A1(n13776), .A2(n7319), .B1(n11134), .B2(n11263), .C1(
        n11262), .C2(P2_U3088), .ZN(P2_U3307) );
  XNOR2_X1 U13765 ( .A(n11264), .B(n11272), .ZN(n14814) );
  INV_X1 U13766 ( .A(n11265), .ZN(n11268) );
  AOI21_X1 U13767 ( .B1(n11266), .B2(n11390), .A(n14745), .ZN(n11267) );
  NAND2_X1 U13768 ( .A1(n11268), .A2(n11267), .ZN(n14810) );
  INV_X1 U13769 ( .A(n11403), .ZN(n11269) );
  AOI22_X1 U13770 ( .A1(n14743), .A2(n11390), .B1(n14722), .B2(n11269), .ZN(
        n11270) );
  OAI21_X1 U13771 ( .B1(n14810), .B2(n14186), .A(n11270), .ZN(n11277) );
  XOR2_X1 U13772 ( .A(n11271), .B(n11272), .Z(n11275) );
  AOI22_X1 U13773 ( .A1(n11505), .A2(n14177), .B1(n14178), .B2(n13894), .ZN(
        n11274) );
  NAND2_X1 U13774 ( .A1(n14814), .A2(n14719), .ZN(n11273) );
  OAI211_X1 U13775 ( .C1(n11275), .C2(n14837), .A(n11274), .B(n11273), .ZN(
        n14812) );
  MUX2_X1 U13776 ( .A(n14812), .B(P1_REG2_REG_7__SCAN_IN), .S(n14157), .Z(
        n11276) );
  AOI211_X1 U13777 ( .C1(n14814), .C2(n14748), .A(n11277), .B(n11276), .ZN(
        n11278) );
  INV_X1 U13778 ( .A(n11278), .ZN(P1_U3286) );
  INV_X1 U13779 ( .A(n11279), .ZN(n11280) );
  OAI21_X1 U13780 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n11281), .A(n11280), 
        .ZN(n11282) );
  NAND2_X1 U13781 ( .A1(n11293), .A2(n11282), .ZN(n11283) );
  XNOR2_X1 U13782 ( .A(n14686), .B(n11282), .ZN(n14683) );
  NAND2_X1 U13783 ( .A1(n14683), .A2(n8551), .ZN(n14682) );
  NAND2_X1 U13784 ( .A1(n11283), .A2(n14682), .ZN(n11286) );
  INV_X1 U13785 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14589) );
  NOR2_X1 U13786 ( .A1(n13937), .A2(n14589), .ZN(n11284) );
  AOI21_X1 U13787 ( .B1(n13937), .B2(n14589), .A(n11284), .ZN(n11285) );
  NOR2_X1 U13788 ( .A1(n11285), .A2(n11286), .ZN(n13936) );
  AOI211_X1 U13789 ( .C1(n11286), .C2(n11285), .A(n13936), .B(n13940), .ZN(
        n11290) );
  NAND2_X1 U13790 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14512)
         );
  INV_X1 U13791 ( .A(n14512), .ZN(n11287) );
  AOI21_X1 U13792 ( .B1(n14675), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11287), 
        .ZN(n11288) );
  OAI21_X1 U13793 ( .B1(n13948), .B2(n14673), .A(n11288), .ZN(n11289) );
  NOR2_X1 U13794 ( .A1(n11290), .A2(n11289), .ZN(n11301) );
  NAND2_X1 U13795 ( .A1(n11292), .A2(n11291), .ZN(n11294) );
  NOR2_X1 U13796 ( .A1(n14686), .A2(n11294), .ZN(n11295) );
  XOR2_X1 U13797 ( .A(n11294), .B(n11293), .Z(n14681) );
  NOR2_X1 U13798 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14681), .ZN(n14680) );
  NOR2_X1 U13799 ( .A1(n11295), .A2(n14680), .ZN(n11299) );
  NOR2_X1 U13800 ( .A1(n13948), .A2(n11296), .ZN(n11297) );
  AOI21_X1 U13801 ( .B1(n11296), .B2(n13948), .A(n11297), .ZN(n11298) );
  NAND2_X1 U13802 ( .A1(n11298), .A2(n11299), .ZN(n13947) );
  OAI211_X1 U13803 ( .C1(n11299), .C2(n11298), .A(n14669), .B(n13947), .ZN(
        n11300) );
  NAND2_X1 U13804 ( .A1(n11301), .A2(n11300), .ZN(P1_U3259) );
  NAND2_X1 U13805 ( .A1(n15277), .A2(n11304), .ZN(n11305) );
  XNOR2_X1 U13806 ( .A(n15251), .B(n12200), .ZN(n11425) );
  XNOR2_X1 U13807 ( .A(n11425), .B(n15259), .ZN(n11423) );
  XNOR2_X1 U13808 ( .A(n11424), .B(n11423), .ZN(n11312) );
  NOR2_X1 U13809 ( .A1(n12298), .A2(n15251), .ZN(n11306) );
  AOI211_X1 U13810 ( .C1(n12236), .C2(n15247), .A(n11307), .B(n11306), .ZN(
        n11308) );
  OAI21_X1 U13811 ( .B1(n11309), .B2(n12257), .A(n11308), .ZN(n11310) );
  AOI21_X1 U13812 ( .B1(n15252), .B2(n12295), .A(n11310), .ZN(n11311) );
  OAI21_X1 U13813 ( .B1(n11312), .B2(n12285), .A(n11311), .ZN(P3_U3161) );
  INV_X1 U13814 ( .A(n11326), .ZN(n11313) );
  OR2_X1 U13815 ( .A1(n14825), .A2(n11650), .ZN(n11316) );
  INV_X1 U13816 ( .A(n11317), .ZN(n11319) );
  INV_X1 U13817 ( .A(n11318), .ZN(n11412) );
  OR2_X2 U13818 ( .A1(n11317), .A2(n11412), .ZN(n11410) );
  OAI21_X1 U13819 ( .B1(n11319), .B2(n11318), .A(n11410), .ZN(n14838) );
  AOI211_X1 U13820 ( .C1(n14834), .C2(n14708), .A(n14745), .B(n11417), .ZN(
        n11320) );
  AOI21_X1 U13821 ( .B1(n14177), .B2(n13891), .A(n11320), .ZN(n14836) );
  INV_X1 U13822 ( .A(n14836), .ZN(n11325) );
  INV_X1 U13823 ( .A(n14834), .ZN(n11653) );
  NOR2_X1 U13824 ( .A1(n11598), .A2(n14555), .ZN(n14832) );
  INV_X1 U13825 ( .A(n14832), .ZN(n11321) );
  OAI22_X1 U13826 ( .A1(n14157), .A2(n11321), .B1(n11645), .B2(n14739), .ZN(
        n11322) );
  AOI21_X1 U13827 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n14157), .A(n11322), 
        .ZN(n11323) );
  OAI21_X1 U13828 ( .B1(n11653), .B2(n14337), .A(n11323), .ZN(n11324) );
  AOI21_X1 U13829 ( .B1(n11325), .B2(n6575), .A(n11324), .ZN(n11332) );
  INV_X1 U13830 ( .A(n11328), .ZN(n11329) );
  NAND2_X1 U13831 ( .A1(n14825), .A2(n11598), .ZN(n11330) );
  XNOR2_X1 U13832 ( .A(n11413), .B(n11412), .ZN(n14841) );
  NAND2_X1 U13833 ( .A1(n14841), .A2(n14570), .ZN(n11331) );
  OAI211_X1 U13834 ( .C1(n14838), .C2(n14189), .A(n11332), .B(n11331), .ZN(
        P1_U3283) );
  AOI211_X1 U13835 ( .C1(n14479), .C2(n11335), .A(n11334), .B(n11333), .ZN(
        n11341) );
  INV_X1 U13836 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11336) );
  NOR2_X1 U13837 ( .A1(n15099), .A2(n11336), .ZN(n11337) );
  AOI21_X1 U13838 ( .B1(n13452), .B2(n11339), .A(n11337), .ZN(n11338) );
  OAI21_X1 U13839 ( .B1(n11341), .B2(n15098), .A(n11338), .ZN(P2_U3457) );
  INV_X1 U13840 ( .A(n13418), .ZN(n13371) );
  AOI22_X1 U13841 ( .A1(n13371), .A2(n11339), .B1(n15103), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11340) );
  OAI21_X1 U13842 ( .B1(n11341), .B2(n15103), .A(n11340), .ZN(P2_U3508) );
  XNOR2_X1 U13843 ( .A(n11343), .B(n11345), .ZN(n15090) );
  XOR2_X1 U13844 ( .A(n11344), .B(n11345), .Z(n11348) );
  OAI22_X1 U13845 ( .A1(n11346), .A2(n14441), .B1(n11383), .B2(n14443), .ZN(
        n11347) );
  AOI21_X1 U13846 ( .B1(n11348), .B2(n14456), .A(n11347), .ZN(n11349) );
  OAI21_X1 U13847 ( .B1(n15090), .B2(n8198), .A(n11349), .ZN(n15094) );
  NAND2_X1 U13848 ( .A1(n15094), .A2(n15055), .ZN(n11358) );
  INV_X1 U13849 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11351) );
  OAI22_X1 U13850 ( .A1(n15055), .A2(n11351), .B1(n11350), .B2(n15052), .ZN(
        n11355) );
  INV_X1 U13851 ( .A(n11352), .ZN(n11493) );
  OAI211_X1 U13852 ( .C1(n15093), .C2(n11353), .A(n11493), .B(n14465), .ZN(
        n15091) );
  NOR2_X1 U13853 ( .A1(n15091), .A2(n15061), .ZN(n11354) );
  AOI211_X1 U13854 ( .C1(n15058), .C2(n11356), .A(n11355), .B(n11354), .ZN(
        n11357) );
  OAI211_X1 U13855 ( .C1(n15090), .C2(n13348), .A(n11358), .B(n11357), .ZN(
        P2_U3255) );
  OAI222_X1 U13856 ( .A1(n11360), .A2(P1_U3086), .B1(n14304), .B2(n11372), 
        .C1(n11359), .C2(n14298), .ZN(P1_U3334) );
  INV_X1 U13857 ( .A(n11361), .ZN(n11362) );
  AOI21_X1 U13858 ( .B1(n11364), .B2(n11363), .A(n11362), .ZN(n11371) );
  OAI21_X1 U13859 ( .B1(n14453), .B2(n11494), .A(n11365), .ZN(n11369) );
  OAI22_X1 U13860 ( .A1(n11367), .A2(n13045), .B1(n13044), .B2(n11366), .ZN(
        n11368) );
  AOI211_X1 U13861 ( .C1(n11551), .C2(n14451), .A(n11369), .B(n11368), .ZN(
        n11370) );
  OAI21_X1 U13862 ( .B1(n11371), .B2(n13059), .A(n11370), .ZN(P2_U3208) );
  OAI222_X1 U13863 ( .A1(n13776), .A2(n11374), .B1(P2_U3088), .B2(n11373), 
        .C1(n11134), .C2(n11372), .ZN(P2_U3306) );
  INV_X1 U13864 ( .A(n11375), .ZN(n11377) );
  INV_X1 U13865 ( .A(SI_24_), .ZN(n11376) );
  OAI222_X1 U13866 ( .A1(P3_U3151), .A2(n11378), .B1(n12961), .B2(n11377), 
        .C1(n11376), .C2(n12962), .ZN(P3_U3271) );
  INV_X1 U13867 ( .A(n14482), .ZN(n11388) );
  OAI21_X1 U13868 ( .B1(n11381), .B2(n11380), .A(n11379), .ZN(n11382) );
  NAND2_X1 U13869 ( .A1(n11382), .A2(n14448), .ZN(n11387) );
  INV_X1 U13870 ( .A(n11468), .ZN(n11385) );
  AND2_X1 U13871 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n13119) );
  OAI22_X1 U13872 ( .A1(n11383), .A2(n13045), .B1(n13044), .B2(n14442), .ZN(
        n11384) );
  AOI211_X1 U13873 ( .C1(n11385), .C2(n13014), .A(n13119), .B(n11384), .ZN(
        n11386) );
  OAI211_X1 U13874 ( .C1(n11388), .C2(n13017), .A(n11387), .B(n11386), .ZN(
        P2_U3196) );
  AND2_X1 U13875 ( .A1(n13893), .A2(n12077), .ZN(n11389) );
  AOI21_X1 U13876 ( .B1(n11390), .B2(n6578), .A(n11389), .ZN(n11509) );
  AOI22_X1 U13877 ( .A1(n11390), .A2(n12079), .B1(n12064), .B2(n13893), .ZN(
        n11391) );
  XNOR2_X1 U13878 ( .A(n11391), .B(n11786), .ZN(n11508) );
  XOR2_X1 U13879 ( .A(n11509), .B(n11508), .Z(n11402) );
  NAND2_X1 U13880 ( .A1(n13872), .A2(n12079), .ZN(n11395) );
  NAND2_X1 U13881 ( .A1(n13894), .A2(n6578), .ZN(n11394) );
  NAND2_X1 U13882 ( .A1(n11395), .A2(n11394), .ZN(n11396) );
  XNOR2_X1 U13883 ( .A(n11396), .B(n11974), .ZN(n11397) );
  AOI22_X1 U13884 ( .A1(n13872), .A2(n12064), .B1(n12077), .B2(n13894), .ZN(
        n11398) );
  XNOR2_X1 U13885 ( .A(n11397), .B(n11398), .ZN(n13869) );
  INV_X1 U13886 ( .A(n11398), .ZN(n11399) );
  NAND2_X1 U13887 ( .A1(n11397), .A2(n11399), .ZN(n11400) );
  OAI211_X1 U13888 ( .C1(n11402), .C2(n11401), .A(n7516), .B(n14551), .ZN(
        n11408) );
  NOR2_X1 U13889 ( .A1(n14554), .A2(n11403), .ZN(n11406) );
  OAI21_X1 U13890 ( .B1(n14526), .B2(n11600), .A(n11404), .ZN(n11405) );
  AOI211_X1 U13891 ( .C1(n14545), .C2(n13894), .A(n11406), .B(n11405), .ZN(
        n11407) );
  OAI211_X1 U13892 ( .C1(n14811), .C2(n14549), .A(n11408), .B(n11407), .ZN(
        P1_U3213) );
  INV_X1 U13893 ( .A(n13890), .ZN(n14527) );
  INV_X1 U13894 ( .A(n13892), .ZN(n14524) );
  OR2_X1 U13895 ( .A1(n14834), .A2(n14524), .ZN(n11409) );
  XNOR2_X1 U13896 ( .A(n11526), .B(n11416), .ZN(n11411) );
  OAI222_X1 U13897 ( .A1(n14557), .A2(n14527), .B1(n11411), .B2(n14837), .C1(
        n14555), .C2(n14524), .ZN(n14607) );
  INV_X1 U13898 ( .A(n14607), .ZN(n11422) );
  NAND2_X1 U13899 ( .A1(n11413), .A2(n11412), .ZN(n11415) );
  OR2_X1 U13900 ( .A1(n14834), .A2(n13892), .ZN(n11414) );
  XOR2_X1 U13901 ( .A(n11534), .B(n11416), .Z(n14609) );
  INV_X1 U13902 ( .A(n14537), .ZN(n14606) );
  OAI211_X1 U13903 ( .C1(n14606), .C2(n11417), .A(n6719), .B(n14725), .ZN(
        n14605) );
  OAI22_X1 U13904 ( .A1(n14741), .A2(n10364), .B1(n14540), .B2(n14739), .ZN(
        n11418) );
  AOI21_X1 U13905 ( .B1(n14537), .B2(n14743), .A(n11418), .ZN(n11419) );
  OAI21_X1 U13906 ( .B1(n14605), .B2(n14186), .A(n11419), .ZN(n11420) );
  AOI21_X1 U13907 ( .B1(n14609), .B2(n14570), .A(n11420), .ZN(n11421) );
  OAI21_X1 U13908 ( .B1(n11422), .B2(n14157), .A(n11421), .ZN(P1_U3282) );
  XNOR2_X1 U13909 ( .A(n11480), .B(n12200), .ZN(n11444) );
  XNOR2_X1 U13910 ( .A(n11444), .B(n15233), .ZN(n11430) );
  INV_X1 U13911 ( .A(n11448), .ZN(n11428) );
  AOI21_X1 U13912 ( .B1(n11430), .B2(n11429), .A(n11428), .ZN(n11435) );
  AND2_X1 U13913 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n15127) );
  AOI21_X1 U13914 ( .B1(n12282), .B2(n11480), .A(n15127), .ZN(n11431) );
  OAI21_X1 U13915 ( .B1(n12257), .B2(n15259), .A(n11431), .ZN(n11433) );
  NOR2_X1 U13916 ( .A1(n12178), .A2(n11478), .ZN(n11432) );
  AOI211_X1 U13917 ( .C1(n12236), .C2(n12521), .A(n11433), .B(n11432), .ZN(
        n11434) );
  OAI21_X1 U13918 ( .B1(n11435), .B2(n12285), .A(n11434), .ZN(P3_U3171) );
  XNOR2_X1 U13919 ( .A(n11437), .B(n11436), .ZN(n11443) );
  NAND2_X1 U13920 ( .A1(n13073), .A2(n13336), .ZN(n11439) );
  NAND2_X1 U13921 ( .A1(n13075), .A2(n13335), .ZN(n11438) );
  NAND2_X1 U13922 ( .A1(n11439), .A2(n11438), .ZN(n11555) );
  AOI22_X1 U13923 ( .A1(n14450), .A2(n11555), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11440) );
  OAI21_X1 U13924 ( .B1(n11561), .B2(n14453), .A(n11440), .ZN(n11441) );
  AOI21_X1 U13925 ( .B1(n11563), .B2(n14451), .A(n11441), .ZN(n11442) );
  OAI21_X1 U13926 ( .B1(n11443), .B2(n13059), .A(n11442), .ZN(P2_U3206) );
  XNOR2_X1 U13927 ( .A(n11454), .B(n12157), .ZN(n11707) );
  XNOR2_X1 U13928 ( .A(n11707), .B(n14425), .ZN(n11446) );
  NAND2_X1 U13929 ( .A1(n11444), .A2(n15233), .ZN(n11447) );
  AND2_X1 U13930 ( .A1(n11446), .A2(n11447), .ZN(n11445) );
  NAND2_X1 U13931 ( .A1(n11708), .A2(n12269), .ZN(n11457) );
  AOI21_X1 U13932 ( .B1(n11448), .B2(n11447), .A(n11446), .ZN(n11456) );
  INV_X1 U13933 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11449) );
  NOR2_X1 U13934 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11449), .ZN(n15137) );
  AOI21_X1 U13935 ( .B1(n12291), .B2(n15247), .A(n15137), .ZN(n11452) );
  INV_X1 U13936 ( .A(n11450), .ZN(n15239) );
  NAND2_X1 U13937 ( .A1(n12295), .A2(n15239), .ZN(n11451) );
  OAI211_X1 U13938 ( .C1(n15234), .C2(n12293), .A(n11452), .B(n11451), .ZN(
        n11453) );
  AOI21_X1 U13939 ( .B1(n11454), .B2(n12282), .A(n11453), .ZN(n11455) );
  OAI21_X1 U13940 ( .B1(n11457), .B2(n11456), .A(n11455), .ZN(P3_U3157) );
  XNOR2_X1 U13941 ( .A(n11458), .B(n11459), .ZN(n14486) );
  NAND2_X1 U13942 ( .A1(n14486), .A2(n13333), .ZN(n11466) );
  NAND2_X1 U13943 ( .A1(n11460), .A2(n11459), .ZN(n11461) );
  NAND3_X1 U13944 ( .A1(n11462), .A2(n14456), .A3(n11461), .ZN(n11464) );
  AOI22_X1 U13945 ( .A1(n13335), .A2(n13076), .B1(n13074), .B2(n13336), .ZN(
        n11463) );
  AND2_X1 U13946 ( .A1(n11464), .A2(n11463), .ZN(n11465) );
  AND2_X1 U13947 ( .A1(n11466), .A2(n11465), .ZN(n14488) );
  AOI21_X1 U13948 ( .B1(n11491), .B2(n14482), .A(n9935), .ZN(n11467) );
  NAND2_X1 U13949 ( .A1(n11467), .A2(n11559), .ZN(n14484) );
  OAI22_X1 U13950 ( .A1(n15055), .A2(n13120), .B1(n11468), .B2(n15052), .ZN(
        n11469) );
  AOI21_X1 U13951 ( .B1(n14482), .B2(n15058), .A(n11469), .ZN(n11470) );
  OAI21_X1 U13952 ( .B1(n14484), .B2(n15061), .A(n11470), .ZN(n11471) );
  AOI21_X1 U13953 ( .B1(n14486), .B2(n11858), .A(n11471), .ZN(n11472) );
  OAI21_X1 U13954 ( .B1(n14488), .B2(n13358), .A(n11472), .ZN(P2_U3253) );
  XOR2_X1 U13955 ( .A(n11473), .B(n12482), .Z(n15367) );
  OAI211_X1 U13956 ( .C1(n11475), .C2(n9400), .A(n15319), .B(n11474), .ZN(
        n11477) );
  AOI22_X1 U13957 ( .A1(n12521), .A2(n15322), .B1(n15323), .B2(n12522), .ZN(
        n11476) );
  OAI211_X1 U13958 ( .C1(n15327), .C2(n15367), .A(n11477), .B(n11476), .ZN(
        n15370) );
  NAND2_X1 U13959 ( .A1(n15370), .A2(n15330), .ZN(n11482) );
  OAI22_X1 U13960 ( .A1(n15330), .A2(n9381), .B1(n11478), .B2(n15312), .ZN(
        n11479) );
  AOI21_X1 U13961 ( .B1(n12695), .B2(n11480), .A(n11479), .ZN(n11481) );
  OAI211_X1 U13962 ( .C1(n15367), .C2(n12698), .A(n11482), .B(n11481), .ZN(
        P3_U3224) );
  XOR2_X1 U13963 ( .A(n11483), .B(n11487), .Z(n11547) );
  INV_X1 U13964 ( .A(n11547), .ZN(n11500) );
  INV_X1 U13965 ( .A(n6743), .ZN(n11485) );
  AOI21_X1 U13966 ( .B1(n11487), .B2(n11486), .A(n11485), .ZN(n11490) );
  NAND2_X1 U13967 ( .A1(n11547), .A2(n13333), .ZN(n11489) );
  AOI22_X1 U13968 ( .A1(n13335), .A2(n13077), .B1(n13075), .B2(n13336), .ZN(
        n11488) );
  OAI211_X1 U13969 ( .C1(n11490), .C2(n13340), .A(n11489), .B(n11488), .ZN(
        n11545) );
  NAND2_X1 U13970 ( .A1(n11545), .A2(n15055), .ZN(n11499) );
  INV_X1 U13971 ( .A(n11491), .ZN(n11492) );
  AOI211_X1 U13972 ( .C1(n11551), .C2(n11493), .A(n9942), .B(n11492), .ZN(
        n11546) );
  NOR2_X1 U13973 ( .A1(n11548), .A2(n13360), .ZN(n11497) );
  OAI22_X1 U13974 ( .A1(n15055), .A2(n11495), .B1(n11494), .B2(n15052), .ZN(
        n11496) );
  AOI211_X1 U13975 ( .C1(n11546), .C2(n14467), .A(n11497), .B(n11496), .ZN(
        n11498) );
  OAI211_X1 U13976 ( .C1(n11500), .C2(n13348), .A(n11499), .B(n11498), .ZN(
        P2_U3254) );
  INV_X1 U13977 ( .A(n11501), .ZN(n11503) );
  OAI222_X1 U13978 ( .A1(n11504), .A2(P3_U3151), .B1(n12961), .B2(n11503), 
        .C1(n11502), .C2(n12962), .ZN(P3_U3270) );
  AOI22_X1 U13979 ( .A1(n11506), .A2(n12064), .B1(n12077), .B2(n11505), .ZN(
        n11593) );
  AOI22_X1 U13980 ( .A1(n11506), .A2(n12079), .B1(n12064), .B2(n11505), .ZN(
        n11507) );
  XNOR2_X1 U13981 ( .A(n11507), .B(n11786), .ZN(n11592) );
  XOR2_X1 U13982 ( .A(n11593), .B(n11592), .Z(n11516) );
  INV_X1 U13983 ( .A(n11508), .ZN(n11511) );
  INV_X1 U13984 ( .A(n11509), .ZN(n11510) );
  NAND2_X1 U13985 ( .A1(n11511), .A2(n11510), .ZN(n11512) );
  OAI21_X1 U13986 ( .B1(n11516), .B2(n11515), .A(n11596), .ZN(n11517) );
  NAND2_X1 U13987 ( .A1(n11517), .A2(n14551), .ZN(n11523) );
  NOR2_X1 U13988 ( .A1(n14554), .A2(n11518), .ZN(n11521) );
  OAI21_X1 U13989 ( .B1(n14526), .B2(n11598), .A(n11519), .ZN(n11520) );
  AOI211_X1 U13990 ( .C1(n14545), .C2(n13893), .A(n11521), .B(n11520), .ZN(
        n11522) );
  OAI211_X1 U13991 ( .C1(n14817), .C2(n14549), .A(n11523), .B(n11522), .ZN(
        P1_U3221) );
  INV_X1 U13992 ( .A(n13891), .ZN(n11647) );
  NOR2_X1 U13993 ( .A1(n14537), .A2(n11647), .ZN(n11525) );
  NAND2_X1 U13994 ( .A1(n14537), .A2(n11647), .ZN(n11524) );
  INV_X1 U13995 ( .A(n11575), .ZN(n11573) );
  INV_X1 U13996 ( .A(n11536), .ZN(n11527) );
  OAI211_X1 U13997 ( .C1(n11528), .C2(n11527), .A(n11676), .B(n14738), .ZN(
        n11531) );
  NAND2_X1 U13998 ( .A1(n13890), .A2(n14178), .ZN(n11529) );
  OAI21_X1 U13999 ( .B1(n14556), .B2(n14557), .A(n11529), .ZN(n13843) );
  INV_X1 U14000 ( .A(n13843), .ZN(n11530) );
  AND2_X1 U14001 ( .A1(n11531), .A2(n11530), .ZN(n11658) );
  INV_X1 U14002 ( .A(n11532), .ZN(n11533) );
  OR2_X1 U14003 ( .A1(n11537), .A2(n11536), .ZN(n11538) );
  NAND2_X1 U14004 ( .A1(n11685), .A2(n11538), .ZN(n11656) );
  INV_X1 U14005 ( .A(n11799), .ZN(n14338) );
  AOI21_X1 U14006 ( .B1(n11579), .B2(n13847), .A(n14745), .ZN(n11539) );
  NAND2_X1 U14007 ( .A1(n11539), .A2(n11679), .ZN(n11654) );
  OAI22_X1 U14008 ( .A1(n14741), .A2(n11540), .B1(n13845), .B2(n14739), .ZN(
        n11541) );
  AOI21_X1 U14009 ( .B1(n13847), .B2(n14743), .A(n11541), .ZN(n11542) );
  OAI21_X1 U14010 ( .B1(n11654), .B2(n14186), .A(n11542), .ZN(n11543) );
  AOI21_X1 U14011 ( .B1(n11656), .B2(n14570), .A(n11543), .ZN(n11544) );
  OAI21_X1 U14012 ( .B1(n11658), .B2(n14157), .A(n11544), .ZN(P1_U3280) );
  AOI211_X1 U14013 ( .C1(n15097), .C2(n11547), .A(n11546), .B(n11545), .ZN(
        n11553) );
  OAI22_X1 U14014 ( .A1(n11548), .A2(n13468), .B1(n15099), .B2(n7786), .ZN(
        n11549) );
  INV_X1 U14015 ( .A(n11549), .ZN(n11550) );
  OAI21_X1 U14016 ( .B1(n11553), .B2(n15098), .A(n11550), .ZN(P2_U3463) );
  AOI22_X1 U14017 ( .A1(n11551), .A2(n13371), .B1(n15103), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11552) );
  OAI21_X1 U14018 ( .B1(n11553), .B2(n15103), .A(n11552), .ZN(P2_U3510) );
  XNOR2_X1 U14019 ( .A(n11554), .B(n11557), .ZN(n11556) );
  AOI21_X1 U14020 ( .B1(n11556), .B2(n14456), .A(n11555), .ZN(n14476) );
  XOR2_X1 U14021 ( .A(n11558), .B(n11557), .Z(n14480) );
  INV_X1 U14022 ( .A(n11559), .ZN(n11560) );
  OAI211_X1 U14023 ( .C1(n14477), .C2(n11560), .A(n7096), .B(n14465), .ZN(
        n14475) );
  INV_X1 U14024 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n13140) );
  OAI22_X1 U14025 ( .A1(n15055), .A2(n13140), .B1(n11561), .B2(n15052), .ZN(
        n11562) );
  AOI21_X1 U14026 ( .B1(n11563), .B2(n15058), .A(n11562), .ZN(n11564) );
  OAI21_X1 U14027 ( .B1(n14475), .B2(n15061), .A(n11564), .ZN(n11565) );
  AOI21_X1 U14028 ( .B1(n14480), .B2(n15063), .A(n11565), .ZN(n11566) );
  OAI21_X1 U14029 ( .B1(n13358), .B2(n14476), .A(n11566), .ZN(P2_U3252) );
  INV_X1 U14030 ( .A(n11567), .ZN(n11568) );
  AND2_X1 U14031 ( .A1(n11569), .A2(n11568), .ZN(n11585) );
  XNOR2_X1 U14032 ( .A(n11574), .B(n11573), .ZN(n14340) );
  XNOR2_X1 U14033 ( .A(n11576), .B(n11575), .ZN(n11578) );
  AOI22_X1 U14034 ( .A1(n11674), .A2(n14177), .B1(n14178), .B2(n13891), .ZN(
        n11807) );
  INV_X1 U14035 ( .A(n11807), .ZN(n11577) );
  AOI21_X1 U14036 ( .B1(n11578), .B2(n14738), .A(n11577), .ZN(n14345) );
  AOI211_X1 U14037 ( .C1(n11799), .C2(n6719), .A(n14745), .B(n6992), .ZN(
        n14343) );
  AOI21_X1 U14038 ( .B1(n11799), .B2(n14833), .A(n14343), .ZN(n11580) );
  OAI211_X1 U14039 ( .C1(n14793), .C2(n14340), .A(n14345), .B(n11580), .ZN(
        n11586) );
  NAND2_X1 U14040 ( .A1(n11586), .A2(n14858), .ZN(n11581) );
  OAI21_X1 U14041 ( .B1(n14858), .B2(n10371), .A(n11581), .ZN(P1_U3540) );
  NOR2_X1 U14042 ( .A1(n11583), .A2(n11582), .ZN(n11584) );
  INV_X1 U14043 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n13704) );
  NAND2_X1 U14044 ( .A1(n11586), .A2(n14844), .ZN(n11587) );
  OAI21_X1 U14045 ( .B1(n14844), .B2(n13704), .A(n11587), .ZN(P1_U3495) );
  INV_X1 U14046 ( .A(n11588), .ZN(n11589) );
  OAI222_X1 U14047 ( .A1(n13776), .A2(n11591), .B1(P2_U3088), .B2(n11590), 
        .C1(n11134), .C2(n11589), .ZN(P2_U3305) );
  INV_X1 U14048 ( .A(n11592), .ZN(n11595) );
  INV_X1 U14049 ( .A(n11593), .ZN(n11594) );
  OAI22_X1 U14050 ( .A1(n14825), .A2(n11597), .B1(n11598), .B2(n6586), .ZN(
        n11635) );
  OAI22_X1 U14051 ( .A1(n14825), .A2(n12036), .B1(n11598), .B2(n11597), .ZN(
        n11599) );
  XNOR2_X1 U14052 ( .A(n11599), .B(n11974), .ZN(n11634) );
  XOR2_X1 U14053 ( .A(n11635), .B(n11634), .Z(n11638) );
  XOR2_X1 U14054 ( .A(n11639), .B(n11638), .Z(n11606) );
  OAI22_X1 U14055 ( .A1(n14524), .A2(n14557), .B1(n11600), .B2(n14555), .ZN(
        n14701) );
  NAND2_X1 U14056 ( .A1(n14701), .A2(n14517), .ZN(n11603) );
  INV_X1 U14057 ( .A(n11601), .ZN(n11602) );
  OAI211_X1 U14058 ( .C1(n14554), .C2(n14703), .A(n11603), .B(n11602), .ZN(
        n11604) );
  AOI21_X1 U14059 ( .B1(n14705), .B2(n14536), .A(n11604), .ZN(n11605) );
  OAI21_X1 U14060 ( .B1(n11606), .B2(n14532), .A(n11605), .ZN(P1_U3231) );
  INV_X1 U14061 ( .A(n11607), .ZN(n11608) );
  OAI222_X1 U14062 ( .A1(n11610), .A2(P3_U3151), .B1(n12962), .B2(n11609), 
        .C1(n12961), .C2(n11608), .ZN(P3_U3269) );
  NAND2_X1 U14063 ( .A1(n11614), .A2(n6726), .ZN(n11612) );
  OAI211_X1 U14064 ( .C1(n11613), .C2(n13776), .A(n11612), .B(n11611), .ZN(
        P2_U3304) );
  NAND2_X1 U14065 ( .A1(n11614), .A2(n14292), .ZN(n11616) );
  OAI211_X1 U14066 ( .C1(n11617), .C2(n14298), .A(n11616), .B(n11615), .ZN(
        P1_U3332) );
  AND2_X1 U14067 ( .A1(n11619), .A2(n11618), .ZN(n11622) );
  OAI211_X1 U14068 ( .C1(n11622), .C2(n11621), .A(n11620), .B(n15319), .ZN(
        n11624) );
  AOI22_X1 U14069 ( .A1(n15322), .A2(n12518), .B1(n12520), .B2(n15323), .ZN(
        n11623) );
  NAND2_X1 U14070 ( .A1(n11624), .A2(n11623), .ZN(n14431) );
  INV_X1 U14071 ( .A(n14431), .ZN(n11631) );
  INV_X1 U14072 ( .A(n11736), .ZN(n11625) );
  NOR2_X1 U14073 ( .A1(n11625), .A2(n15368), .ZN(n14432) );
  OAI22_X1 U14074 ( .A1(n15330), .A2(n11626), .B1(n11731), .B2(n15312), .ZN(
        n11627) );
  AOI21_X1 U14075 ( .B1(n15305), .B2(n14432), .A(n11627), .ZN(n11630) );
  XNOR2_X1 U14076 ( .A(n11628), .B(n12485), .ZN(n14433) );
  OR2_X1 U14077 ( .A1(n15297), .A2(n15329), .ZN(n15250) );
  NAND2_X1 U14078 ( .A1(n14433), .A2(n15265), .ZN(n11629) );
  OAI211_X1 U14079 ( .C1(n11631), .C2(n15333), .A(n11630), .B(n11629), .ZN(
        P3_U3221) );
  INV_X1 U14080 ( .A(n11632), .ZN(n11633) );
  INV_X1 U14081 ( .A(SI_27_), .ZN(n13623) );
  OAI222_X1 U14082 ( .A1(P3_U3151), .A2(n12589), .B1(n12961), .B2(n11633), 
        .C1(n13623), .C2(n12962), .ZN(P3_U3268) );
  INV_X1 U14083 ( .A(n11634), .ZN(n11637) );
  INV_X1 U14084 ( .A(n11635), .ZN(n11636) );
  NAND2_X1 U14085 ( .A1(n14834), .A2(n12079), .ZN(n11641) );
  NAND2_X1 U14086 ( .A1(n13892), .A2(n12064), .ZN(n11640) );
  NAND2_X1 U14087 ( .A1(n11641), .A2(n11640), .ZN(n11642) );
  XNOR2_X1 U14088 ( .A(n11642), .B(n11974), .ZN(n11791) );
  AND2_X1 U14089 ( .A1(n13892), .A2(n12077), .ZN(n11643) );
  AOI21_X1 U14090 ( .B1(n14834), .B2(n12064), .A(n11643), .ZN(n11789) );
  XNOR2_X1 U14091 ( .A(n11791), .B(n11789), .ZN(n11644) );
  OAI211_X1 U14092 ( .C1(n6718), .C2(n11644), .A(n11793), .B(n14551), .ZN(
        n11652) );
  NOR2_X1 U14093 ( .A1(n14554), .A2(n11645), .ZN(n11649) );
  OAI22_X1 U14094 ( .A1(n14526), .A2(n11647), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11646), .ZN(n11648) );
  AOI211_X1 U14095 ( .C1(n14545), .C2(n11650), .A(n11649), .B(n11648), .ZN(
        n11651) );
  OAI211_X1 U14096 ( .C1(n11653), .C2(n14549), .A(n11652), .B(n11651), .ZN(
        P1_U3217) );
  OAI21_X1 U14097 ( .B1(n11973), .B2(n14824), .A(n11654), .ZN(n11655) );
  AOI21_X1 U14098 ( .B1(n11656), .B2(n14840), .A(n11655), .ZN(n11657) );
  AND2_X1 U14099 ( .A1(n11658), .A2(n11657), .ZN(n11660) );
  MUX2_X1 U14100 ( .A(n10606), .B(n11660), .S(n14858), .Z(n11659) );
  INV_X1 U14101 ( .A(n11659), .ZN(P1_U3541) );
  INV_X1 U14102 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11661) );
  MUX2_X1 U14103 ( .A(n11661), .B(n11660), .S(n14844), .Z(n11662) );
  INV_X1 U14104 ( .A(n11662), .ZN(P1_U3498) );
  OAI211_X1 U14105 ( .C1(n11664), .C2(n12490), .A(n11663), .B(n15319), .ZN(
        n11666) );
  AOI22_X1 U14106 ( .A1(n12519), .A2(n15323), .B1(n15322), .B2(n12517), .ZN(
        n11665) );
  NAND2_X1 U14107 ( .A1(n11666), .A2(n11665), .ZN(n11777) );
  INV_X1 U14108 ( .A(n11777), .ZN(n11672) );
  INV_X1 U14109 ( .A(n12490), .ZN(n12396) );
  XNOR2_X1 U14110 ( .A(n11667), .B(n12396), .ZN(n11778) );
  INV_X1 U14111 ( .A(n11668), .ZN(n11819) );
  AOI22_X1 U14112 ( .A1(n15333), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15253), 
        .B2(n11819), .ZN(n11669) );
  OAI21_X1 U14113 ( .B1(n11816), .B2(n12812), .A(n11669), .ZN(n11670) );
  AOI21_X1 U14114 ( .B1(n11778), .B2(n15265), .A(n11670), .ZN(n11671) );
  OAI21_X1 U14115 ( .B1(n11672), .B2(n15333), .A(n11671), .ZN(P3_U3220) );
  INV_X1 U14116 ( .A(n14504), .ZN(n11678) );
  OR2_X1 U14117 ( .A1(n14494), .A2(n14555), .ZN(n11673) );
  OAI21_X1 U14118 ( .B1(n14493), .B2(n14557), .A(n11673), .ZN(n14597) );
  NAND2_X1 U14119 ( .A1(n11973), .A2(n11674), .ZN(n11675) );
  NAND2_X1 U14120 ( .A1(n11676), .A2(n11675), .ZN(n11911) );
  XNOR2_X1 U14121 ( .A(n11911), .B(n11687), .ZN(n11677) );
  NOR2_X1 U14122 ( .A1(n11677), .A2(n14837), .ZN(n14604) );
  AOI211_X1 U14123 ( .C1(n14722), .C2(n11678), .A(n14597), .B(n14604), .ZN(
        n11693) );
  NOR2_X2 U14124 ( .A1(n11679), .A2(n14598), .ZN(n14564) );
  NAND2_X1 U14125 ( .A1(n11679), .A2(n14598), .ZN(n11680) );
  NAND2_X1 U14126 ( .A1(n11680), .A2(n14725), .ZN(n11681) );
  NOR2_X1 U14127 ( .A1(n14564), .A2(n11681), .ZN(n14599) );
  INV_X1 U14128 ( .A(n14598), .ZN(n11683) );
  OAI22_X1 U14129 ( .A1(n11683), .A2(n14337), .B1(n11682), .B2(n14741), .ZN(
        n11691) );
  NAND2_X1 U14130 ( .A1(n11973), .A2(n14494), .ZN(n11684) );
  NAND2_X1 U14131 ( .A1(n11685), .A2(n11684), .ZN(n11688) );
  NAND2_X1 U14132 ( .A1(n11688), .A2(n11687), .ZN(n11689) );
  NAND2_X1 U14133 ( .A1(n11889), .A2(n11689), .ZN(n14602) );
  NOR2_X1 U14134 ( .A1(n14602), .A2(n14339), .ZN(n11690) );
  AOI211_X1 U14135 ( .C1(n6575), .C2(n14599), .A(n11691), .B(n11690), .ZN(
        n11692) );
  OAI21_X1 U14136 ( .B1(n11693), .B2(n14157), .A(n11692), .ZN(P1_U3279) );
  OAI222_X1 U14137 ( .A1(n11695), .A2(P1_U3086), .B1(n14304), .B2(n11697), 
        .C1(n11694), .C2(n14298), .ZN(P1_U3331) );
  INV_X1 U14138 ( .A(n11696), .ZN(n11698) );
  OAI222_X1 U14139 ( .A1(P2_U3088), .A2(n11698), .B1(n11134), .B2(n11697), 
        .C1(n13595), .C2(n13776), .ZN(P2_U3303) );
  XNOR2_X1 U14140 ( .A(n11700), .B(n11699), .ZN(n11706) );
  OR2_X1 U14141 ( .A1(n11847), .A2(n14443), .ZN(n11702) );
  NAND2_X1 U14142 ( .A1(n13073), .A2(n13335), .ZN(n11701) );
  NAND2_X1 U14143 ( .A1(n11702), .A2(n11701), .ZN(n11760) );
  AOI22_X1 U14144 ( .A1(n14450), .A2(n11760), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11703) );
  OAI21_X1 U14145 ( .B1(n11753), .B2(n14453), .A(n11703), .ZN(n11704) );
  AOI21_X1 U14146 ( .B1(n11841), .B2(n14451), .A(n11704), .ZN(n11705) );
  OAI21_X1 U14147 ( .B1(n11706), .B2(n13059), .A(n11705), .ZN(P2_U3213) );
  XNOR2_X1 U14148 ( .A(n11719), .B(n12157), .ZN(n11709) );
  NAND2_X1 U14149 ( .A1(n11710), .A2(n11709), .ZN(n11711) );
  INV_X1 U14150 ( .A(n11714), .ZN(n11712) );
  NAND2_X1 U14151 ( .A1(n11712), .A2(n15234), .ZN(n11726) );
  INV_X1 U14152 ( .A(n11726), .ZN(n11713) );
  AOI21_X1 U14153 ( .B1(n12520), .B2(n11714), .A(n11713), .ZN(n11721) );
  AND2_X1 U14154 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n15161) );
  AOI21_X1 U14155 ( .B1(n12291), .B2(n12521), .A(n15161), .ZN(n11717) );
  INV_X1 U14156 ( .A(n11715), .ZN(n14428) );
  NAND2_X1 U14157 ( .A1(n12295), .A2(n14428), .ZN(n11716) );
  OAI211_X1 U14158 ( .C1(n14426), .C2(n12293), .A(n11717), .B(n11716), .ZN(
        n11718) );
  AOI21_X1 U14159 ( .B1(n11719), .B2(n12282), .A(n11718), .ZN(n11720) );
  OAI21_X1 U14160 ( .B1(n11721), .B2(n12285), .A(n11720), .ZN(P3_U3176) );
  INV_X1 U14161 ( .A(n11722), .ZN(n11724) );
  OAI222_X1 U14162 ( .A1(n12961), .A2(n11724), .B1(n12962), .B2(n11723), .C1(
        P3_U3151), .C2(n12507), .ZN(P3_U3267) );
  NAND2_X1 U14163 ( .A1(n11726), .A2(n11725), .ZN(n11813) );
  XNOR2_X1 U14164 ( .A(n11736), .B(n12200), .ZN(n11727) );
  AND2_X1 U14165 ( .A1(n11727), .A2(n14426), .ZN(n11812) );
  INV_X1 U14166 ( .A(n11812), .ZN(n11729) );
  INV_X1 U14167 ( .A(n11727), .ZN(n11728) );
  NAND2_X1 U14168 ( .A1(n11728), .A2(n12519), .ZN(n11811) );
  NAND2_X1 U14169 ( .A1(n11729), .A2(n11811), .ZN(n11730) );
  XNOR2_X1 U14170 ( .A(n11813), .B(n11730), .ZN(n11738) );
  INV_X1 U14171 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n13664) );
  NOR2_X1 U14172 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13664), .ZN(n15179) );
  AOI21_X1 U14173 ( .B1(n12291), .B2(n12520), .A(n15179), .ZN(n11734) );
  INV_X1 U14174 ( .A(n11731), .ZN(n11732) );
  NAND2_X1 U14175 ( .A1(n12295), .A2(n11732), .ZN(n11733) );
  OAI211_X1 U14176 ( .C1(n12127), .C2(n12293), .A(n11734), .B(n11733), .ZN(
        n11735) );
  AOI21_X1 U14177 ( .B1(n12282), .B2(n11736), .A(n11735), .ZN(n11737) );
  OAI21_X1 U14178 ( .B1(n11738), .B2(n12285), .A(n11737), .ZN(P3_U3164) );
  OAI211_X1 U14179 ( .C1(n11740), .C2(n12489), .A(n11739), .B(n15319), .ZN(
        n11742) );
  AOI22_X1 U14180 ( .A1(n12791), .A2(n15322), .B1(n15323), .B2(n12518), .ZN(
        n11741) );
  NAND2_X1 U14181 ( .A1(n11742), .A2(n11741), .ZN(n12892) );
  INV_X1 U14182 ( .A(n12892), .ZN(n11748) );
  XNOR2_X1 U14183 ( .A(n11743), .B(n12489), .ZN(n12893) );
  NOR2_X1 U14184 ( .A1(n12948), .A2(n12812), .ZN(n11746) );
  OAI22_X1 U14185 ( .A1(n15330), .A2(n11744), .B1(n12179), .B2(n15312), .ZN(
        n11745) );
  AOI211_X1 U14186 ( .C1(n12893), .C2(n15265), .A(n11746), .B(n11745), .ZN(
        n11747) );
  OAI21_X1 U14187 ( .B1(n11748), .B2(n15333), .A(n11747), .ZN(P3_U3219) );
  XNOR2_X1 U14188 ( .A(n11749), .B(n11750), .ZN(n11832) );
  NAND2_X1 U14189 ( .A1(n14464), .A2(n11841), .ZN(n11751) );
  NAND3_X1 U14190 ( .A1(n11752), .A2(n14465), .A3(n11751), .ZN(n11833) );
  OAI22_X1 U14191 ( .A1(n15055), .A2(n11754), .B1(n11753), .B2(n15052), .ZN(
        n11755) );
  AOI21_X1 U14192 ( .B1(n11841), .B2(n15058), .A(n11755), .ZN(n11756) );
  OAI21_X1 U14193 ( .B1(n11833), .B2(n15061), .A(n11756), .ZN(n11762) );
  XNOR2_X1 U14194 ( .A(n11757), .B(n11758), .ZN(n11759) );
  NAND2_X1 U14195 ( .A1(n11759), .A2(n14456), .ZN(n11836) );
  INV_X1 U14196 ( .A(n11760), .ZN(n11834) );
  AOI21_X1 U14197 ( .B1(n11836), .B2(n11834), .A(n13358), .ZN(n11761) );
  AOI211_X1 U14198 ( .C1(n11832), .C2(n15063), .A(n11762), .B(n11761), .ZN(
        n11763) );
  INV_X1 U14199 ( .A(n11763), .ZN(P2_U3250) );
  XNOR2_X1 U14200 ( .A(n11765), .B(n11764), .ZN(n11766) );
  NAND2_X1 U14201 ( .A1(n11766), .A2(n14456), .ZN(n11768) );
  AOI22_X1 U14202 ( .A1(n13334), .A2(n13336), .B1(n13072), .B2(n13335), .ZN(
        n11767) );
  NAND2_X1 U14203 ( .A1(n11768), .A2(n11767), .ZN(n13448) );
  AOI21_X1 U14204 ( .B1(n11825), .B2(n14460), .A(n13448), .ZN(n11776) );
  OAI211_X1 U14205 ( .C1(n13445), .C2(n11769), .A(n14465), .B(n13355), .ZN(
        n13444) );
  INV_X1 U14206 ( .A(n13444), .ZN(n11771) );
  INV_X1 U14207 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13148) );
  OAI22_X1 U14208 ( .A1(n13445), .A2(n13360), .B1(n15055), .B2(n13148), .ZN(
        n11770) );
  AOI21_X1 U14209 ( .B1(n11771), .B2(n14467), .A(n11770), .ZN(n11775) );
  OR2_X1 U14210 ( .A1(n11773), .A2(n11772), .ZN(n13443) );
  NAND3_X1 U14211 ( .A1(n13443), .A2(n13442), .A3(n15063), .ZN(n11774) );
  OAI211_X1 U14212 ( .C1(n11776), .C2(n13358), .A(n11775), .B(n11774), .ZN(
        P2_U3249) );
  AOI21_X1 U14213 ( .B1(n11778), .B2(n15366), .A(n11777), .ZN(n11781) );
  MUX2_X1 U14214 ( .A(n11779), .B(n11781), .S(n15379), .Z(n11780) );
  OAI21_X1 U14215 ( .B1(n12949), .B2(n11816), .A(n11780), .ZN(P3_U3429) );
  INV_X1 U14216 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n11782) );
  MUX2_X1 U14217 ( .A(n11782), .B(n11781), .S(n15395), .Z(n11783) );
  OAI21_X1 U14218 ( .B1(n12896), .B2(n11816), .A(n11783), .ZN(P3_U3472) );
  NAND2_X1 U14219 ( .A1(n14537), .A2(n12079), .ZN(n11785) );
  NAND2_X1 U14220 ( .A1(n13891), .A2(n12064), .ZN(n11784) );
  NAND2_X1 U14221 ( .A1(n11785), .A2(n11784), .ZN(n11787) );
  XNOR2_X1 U14222 ( .A(n11787), .B(n11786), .ZN(n11796) );
  AND2_X1 U14223 ( .A1(n13891), .A2(n12077), .ZN(n11788) );
  AOI21_X1 U14224 ( .B1(n14537), .B2(n6578), .A(n11788), .ZN(n11794) );
  XNOR2_X1 U14225 ( .A(n11796), .B(n11794), .ZN(n14528) );
  INV_X1 U14226 ( .A(n11789), .ZN(n11790) );
  NAND2_X1 U14227 ( .A1(n11791), .A2(n11790), .ZN(n14529) );
  INV_X1 U14228 ( .A(n11794), .ZN(n11795) );
  AND2_X1 U14229 ( .A1(n13890), .A2(n12077), .ZN(n11798) );
  AOI21_X1 U14230 ( .B1(n11799), .B2(n12064), .A(n11798), .ZN(n11968) );
  NAND2_X1 U14231 ( .A1(n11799), .A2(n12079), .ZN(n11801) );
  NAND2_X1 U14232 ( .A1(n13890), .A2(n12064), .ZN(n11800) );
  NAND2_X1 U14233 ( .A1(n11801), .A2(n11800), .ZN(n11802) );
  XNOR2_X1 U14234 ( .A(n11802), .B(n11974), .ZN(n11970) );
  XOR2_X1 U14235 ( .A(n11968), .B(n11970), .Z(n11804) );
  AOI21_X1 U14236 ( .B1(n11803), .B2(n11804), .A(n14532), .ZN(n11805) );
  NAND2_X1 U14237 ( .A1(n11805), .A2(n11972), .ZN(n11810) );
  INV_X1 U14238 ( .A(n11806), .ZN(n14335) );
  INV_X1 U14239 ( .A(n14554), .ZN(n13837) );
  OAI22_X1 U14240 ( .A1(n11807), .A2(n13835), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10368), .ZN(n11808) );
  AOI21_X1 U14241 ( .B1(n14335), .B2(n13837), .A(n11808), .ZN(n11809) );
  OAI211_X1 U14242 ( .C1(n14338), .C2(n14549), .A(n11810), .B(n11809), .ZN(
        P1_U3224) );
  XNOR2_X1 U14243 ( .A(n11816), .B(n12157), .ZN(n12129) );
  XNOR2_X1 U14244 ( .A(n12129), .B(n12518), .ZN(n11814) );
  XNOR2_X1 U14245 ( .A(n12128), .B(n11814), .ZN(n11821) );
  AND2_X1 U14246 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n15197) );
  AOI21_X1 U14247 ( .B1(n12291), .B2(n12519), .A(n15197), .ZN(n11815) );
  OAI21_X1 U14248 ( .B1(n12806), .B2(n12293), .A(n11815), .ZN(n11818) );
  NOR2_X1 U14249 ( .A1(n11816), .A2(n12298), .ZN(n11817) );
  AOI211_X1 U14250 ( .C1(n11819), .C2(n12295), .A(n11818), .B(n11817), .ZN(
        n11820) );
  OAI21_X1 U14251 ( .B1(n11821), .B2(n12285), .A(n11820), .ZN(P3_U3174) );
  AOI21_X1 U14252 ( .B1(n11824), .B2(n11823), .A(n11822), .ZN(n11831) );
  INV_X1 U14253 ( .A(n11825), .ZN(n11826) );
  NAND2_X1 U14254 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n15013)
         );
  OAI21_X1 U14255 ( .B1(n14453), .B2(n11826), .A(n15013), .ZN(n11828) );
  OAI22_X1 U14256 ( .A1(n14444), .A2(n13045), .B1(n13044), .B2(n13046), .ZN(
        n11827) );
  AOI211_X1 U14257 ( .C1(n11829), .C2(n14451), .A(n11828), .B(n11827), .ZN(
        n11830) );
  OAI21_X1 U14258 ( .B1(n11831), .B2(n13059), .A(n11830), .ZN(P2_U3198) );
  NAND2_X1 U14259 ( .A1(n11832), .A2(n14479), .ZN(n11835) );
  NAND4_X1 U14260 ( .A1(n11836), .A2(n11835), .A3(n11834), .A4(n11833), .ZN(
        n11839) );
  MUX2_X1 U14261 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n11839), .S(n15105), .Z(
        n11837) );
  AOI21_X1 U14262 ( .B1(n13371), .B2(n11841), .A(n11837), .ZN(n11838) );
  INV_X1 U14263 ( .A(n11838), .ZN(P2_U3514) );
  MUX2_X1 U14264 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n11839), .S(n15099), .Z(
        n11840) );
  AOI21_X1 U14265 ( .B1(n13452), .B2(n11841), .A(n11840), .ZN(n11842) );
  INV_X1 U14266 ( .A(n11842), .ZN(P2_U3475) );
  AOI21_X1 U14267 ( .B1(n11846), .B2(n11845), .A(n11844), .ZN(n11853) );
  NAND2_X1 U14268 ( .A1(n13070), .A2(n13336), .ZN(n11849) );
  OR2_X1 U14269 ( .A1(n11847), .A2(n14441), .ZN(n11848) );
  NAND2_X1 U14270 ( .A1(n11849), .A2(n11848), .ZN(n13351) );
  NAND2_X1 U14271 ( .A1(n14450), .A2(n13351), .ZN(n11850) );
  NAND2_X1 U14272 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n15029)
         );
  OAI211_X1 U14273 ( .C1(n14453), .C2(n13356), .A(n11850), .B(n15029), .ZN(
        n11851) );
  AOI21_X1 U14274 ( .B1(n13437), .B2(n14451), .A(n11851), .ZN(n11852) );
  OAI21_X1 U14275 ( .B1(n11853), .B2(n13059), .A(n11852), .ZN(P2_U3200) );
  MUX2_X1 U14276 ( .A(n11854), .B(P2_REG2_REG_3__SCAN_IN), .S(n13358), .Z(
        n11863) );
  OAI22_X1 U14277 ( .A1(n13360), .A2(n11855), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n15052), .ZN(n11856) );
  INV_X1 U14278 ( .A(n11856), .ZN(n11860) );
  NAND2_X1 U14279 ( .A1(n11858), .A2(n11857), .ZN(n11859) );
  OAI211_X1 U14280 ( .C1(n15061), .C2(n11861), .A(n11860), .B(n11859), .ZN(
        n11862) );
  OR2_X1 U14281 ( .A1(n11863), .A2(n11862), .ZN(P2_U3262) );
  INV_X1 U14282 ( .A(n11864), .ZN(n14291) );
  OAI222_X1 U14283 ( .A1(n11134), .A2(n14291), .B1(P2_U3088), .B2(n11865), 
        .C1(n11867), .C2(n13776), .ZN(P2_U3298) );
  INV_X1 U14284 ( .A(n11866), .ZN(n11868) );
  XNOR2_X1 U14285 ( .A(n12312), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n11870) );
  INV_X1 U14286 ( .A(n12299), .ZN(n11873) );
  INV_X1 U14287 ( .A(SI_30_), .ZN(n11872) );
  OAI222_X1 U14288 ( .A1(n12961), .A2(n11873), .B1(n12962), .B2(n11872), .C1(
        P3_U3151), .C2(n11871), .ZN(P3_U3265) );
  INV_X1 U14289 ( .A(n11874), .ZN(n11967) );
  OAI222_X1 U14290 ( .A1(n11134), .A2(n11967), .B1(P2_U3088), .B2(n11875), 
        .C1(n12312), .C2(n13776), .ZN(P2_U3297) );
  INV_X1 U14291 ( .A(n11876), .ZN(n13483) );
  OAI222_X1 U14292 ( .A1(P1_U3086), .A2(n11878), .B1(n14304), .B2(n13483), 
        .C1(n11877), .C2(n14298), .ZN(P1_U3327) );
  INV_X1 U14293 ( .A(n11879), .ZN(n11880) );
  AOI22_X1 U14294 ( .A1(n13358), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n11880), 
        .B2(n14460), .ZN(n11881) );
  OAI21_X1 U14295 ( .B1(n11882), .B2(n13360), .A(n11881), .ZN(n11884) );
  OAI21_X1 U14296 ( .B1(n11887), .B2(n13358), .A(n11886), .ZN(P2_U3236) );
  NAND2_X1 U14297 ( .A1(n14598), .A2(n14544), .ZN(n11888) );
  INV_X1 U14298 ( .A(n14493), .ZN(n14507) );
  INV_X1 U14299 ( .A(n14171), .ZN(n14174) );
  OR2_X1 U14300 ( .A1(n14184), .A2(n14546), .ZN(n11890) );
  NAND2_X1 U14301 ( .A1(n14173), .A2(n11890), .ZN(n14165) );
  NAND2_X1 U14302 ( .A1(n14575), .A2(n14508), .ZN(n11891) );
  NAND2_X1 U14303 ( .A1(n14165), .A2(n11891), .ZN(n11893) );
  OR2_X1 U14304 ( .A1(n14575), .A2(n14508), .ZN(n11892) );
  INV_X1 U14305 ( .A(n11894), .ZN(n11896) );
  INV_X1 U14306 ( .A(n14113), .ZN(n11923) );
  OR2_X1 U14307 ( .A1(n14246), .A2(n13889), .ZN(n11897) );
  INV_X1 U14308 ( .A(n14088), .ZN(n14091) );
  NAND2_X1 U14309 ( .A1(n14101), .A2(n13788), .ZN(n11898) );
  NAND2_X1 U14310 ( .A1(n14235), .A2(n14059), .ZN(n11900) );
  OR2_X1 U14311 ( .A1(n14068), .A2(n13888), .ZN(n11902) );
  NAND2_X1 U14312 ( .A1(n14221), .A2(n14058), .ZN(n11903) );
  INV_X1 U14313 ( .A(n14004), .ZN(n11905) );
  NAND2_X1 U14314 ( .A1(n11905), .A2(n11904), .ZN(n14006) );
  NAND2_X1 U14315 ( .A1(n14006), .A2(n11908), .ZN(n11955) );
  NOR2_X1 U14316 ( .A1(n11955), .A2(n11956), .ZN(n11954) );
  NAND2_X1 U14317 ( .A1(n11911), .A2(n11910), .ZN(n11913) );
  INV_X1 U14318 ( .A(n14567), .ZN(n11914) );
  INV_X1 U14319 ( .A(n14546), .ZN(n14558) );
  INV_X1 U14320 ( .A(n11916), .ZN(n14164) );
  INV_X1 U14321 ( .A(n14508), .ZN(n11917) );
  OR2_X1 U14322 ( .A1(n14575), .A2(n11917), .ZN(n11918) );
  NAND2_X1 U14323 ( .A1(n14144), .A2(n14152), .ZN(n11921) );
  INV_X1 U14324 ( .A(n14159), .ZN(n11919) );
  OR2_X1 U14325 ( .A1(n14265), .A2(n11919), .ZN(n11920) );
  INV_X1 U14326 ( .A(n14146), .ZN(n13863) );
  NAND2_X1 U14327 ( .A1(n14260), .A2(n13863), .ZN(n11922) );
  NAND2_X1 U14328 ( .A1(n14104), .A2(n11923), .ZN(n11926) );
  OR2_X1 U14329 ( .A1(n14246), .A2(n11924), .ZN(n11925) );
  INV_X1 U14330 ( .A(n13788), .ZN(n14106) );
  OR2_X1 U14331 ( .A1(n14101), .A2(n14106), .ZN(n11927) );
  NAND2_X1 U14332 ( .A1(n14078), .A2(n14077), .ZN(n14076) );
  INV_X1 U14333 ( .A(n14059), .ZN(n11928) );
  NAND2_X1 U14334 ( .A1(n14235), .A2(n11928), .ZN(n11929) );
  NAND2_X1 U14335 ( .A1(n14076), .A2(n11929), .ZN(n14055) );
  OR2_X2 U14336 ( .A1(n14055), .A2(n14054), .ZN(n14057) );
  INV_X1 U14337 ( .A(n13888), .ZN(n11930) );
  OR2_X1 U14338 ( .A1(n14068), .A2(n11930), .ZN(n11931) );
  NAND2_X1 U14339 ( .A1(n14221), .A2(n13880), .ZN(n11932) );
  INV_X1 U14340 ( .A(n14023), .ZN(n14027) );
  NAND2_X1 U14341 ( .A1(n14026), .A2(n14027), .ZN(n14025) );
  NOR2_X1 U14342 ( .A1(n11907), .A2(n13887), .ZN(n11948) );
  INV_X1 U14343 ( .A(n11937), .ZN(n14197) );
  INV_X1 U14344 ( .A(n14068), .ZN(n14228) );
  INV_X1 U14345 ( .A(n14592), .ZN(n14561) );
  NAND2_X1 U14346 ( .A1(n14252), .A2(n14135), .ZN(n14121) );
  NAND2_X1 U14347 ( .A1(n11907), .A2(n14035), .ZN(n14017) );
  NOR2_X2 U14348 ( .A1(n11937), .A2(n11960), .ZN(n13999) );
  NAND2_X1 U14349 ( .A1(n14199), .A2(n6575), .ZN(n11945) );
  NAND2_X1 U14350 ( .A1(n11938), .A2(P1_B_REG_SCAN_IN), .ZN(n11939) );
  AND2_X1 U14351 ( .A1(n14177), .A2(n11939), .ZN(n13993) );
  NAND2_X1 U14352 ( .A1(n13885), .A2(n13993), .ZN(n14196) );
  OAI22_X1 U14353 ( .A1(n11941), .A2(n14196), .B1(n11940), .B2(n14739), .ZN(
        n11943) );
  NAND2_X1 U14354 ( .A1(n14011), .A2(n14178), .ZN(n14195) );
  NOR2_X1 U14355 ( .A1(n14157), .A2(n14195), .ZN(n11942) );
  AOI211_X1 U14356 ( .C1(n14157), .C2(P1_REG2_REG_29__SCAN_IN), .A(n11943), 
        .B(n11942), .ZN(n11944) );
  OAI211_X1 U14357 ( .C1(n14197), .C2(n14337), .A(n11945), .B(n11944), .ZN(
        n11946) );
  AOI21_X1 U14358 ( .B1(n14200), .B2(n14571), .A(n11946), .ZN(n11947) );
  OAI21_X1 U14359 ( .B1(n14201), .B2(n14339), .A(n11947), .ZN(P1_U3356) );
  OR3_X1 U14360 ( .A1(n14010), .A2(n11956), .A3(n11948), .ZN(n11949) );
  NAND2_X1 U14361 ( .A1(n13886), .A2(n14177), .ZN(n11952) );
  AOI21_X1 U14362 ( .B1(n11956), .B2(n11955), .A(n11954), .ZN(n11957) );
  INV_X1 U14363 ( .A(n11957), .ZN(n14206) );
  NAND2_X1 U14364 ( .A1(n14157), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n11958) );
  OAI21_X1 U14365 ( .B1(n14739), .B2(n12086), .A(n11958), .ZN(n11959) );
  AOI21_X1 U14366 ( .B1(n14203), .B2(n14743), .A(n11959), .ZN(n11963) );
  AOI21_X1 U14367 ( .B1(n14017), .B2(n14203), .A(n14745), .ZN(n11961) );
  NAND2_X1 U14368 ( .A1(n14202), .A2(n6575), .ZN(n11962) );
  OAI211_X1 U14369 ( .C1(n14206), .C2(n14339), .A(n11963), .B(n11962), .ZN(
        n11964) );
  INV_X1 U14370 ( .A(n11964), .ZN(n11965) );
  OAI21_X1 U14371 ( .B1(n14205), .B2(n14157), .A(n11965), .ZN(P1_U3265) );
  OAI222_X1 U14372 ( .A1(n14304), .A2(n11967), .B1(n11966), .B2(P1_U3086), 
        .C1(n12313), .C2(n14298), .ZN(P1_U3325) );
  INV_X1 U14373 ( .A(n11968), .ZN(n11969) );
  NAND2_X1 U14374 ( .A1(n11970), .A2(n11969), .ZN(n11971) );
  NAND2_X1 U14375 ( .A1(n11972), .A2(n11971), .ZN(n13841) );
  OAI22_X1 U14376 ( .A1(n11973), .A2(n11597), .B1(n14494), .B2(n12034), .ZN(
        n11981) );
  OAI22_X1 U14377 ( .A1(n11973), .A2(n12036), .B1(n14494), .B2(n11597), .ZN(
        n11975) );
  XNOR2_X1 U14378 ( .A(n11975), .B(n11974), .ZN(n11980) );
  XOR2_X1 U14379 ( .A(n11981), .B(n11980), .Z(n13842) );
  NAND2_X1 U14380 ( .A1(n13841), .A2(n13842), .ZN(n13840) );
  NAND2_X1 U14381 ( .A1(n14598), .A2(n12079), .ZN(n11977) );
  NAND2_X1 U14382 ( .A1(n14544), .A2(n6578), .ZN(n11976) );
  NAND2_X1 U14383 ( .A1(n11977), .A2(n11976), .ZN(n11978) );
  XNOR2_X1 U14384 ( .A(n11978), .B(n10389), .ZN(n11986) );
  NOR2_X1 U14385 ( .A1(n14556), .A2(n12034), .ZN(n11979) );
  AOI21_X1 U14386 ( .B1(n14598), .B2(n12064), .A(n11979), .ZN(n11985) );
  XNOR2_X1 U14387 ( .A(n11986), .B(n11985), .ZN(n14495) );
  INV_X1 U14388 ( .A(n11980), .ZN(n11983) );
  INV_X1 U14389 ( .A(n11981), .ZN(n11982) );
  NOR2_X1 U14390 ( .A1(n11983), .A2(n11982), .ZN(n14496) );
  NOR2_X1 U14391 ( .A1(n14495), .A2(n14496), .ZN(n11984) );
  NAND2_X1 U14392 ( .A1(n13840), .A2(n11984), .ZN(n14498) );
  NAND2_X1 U14393 ( .A1(n11986), .A2(n11985), .ZN(n11987) );
  NAND2_X1 U14394 ( .A1(n14592), .A2(n12079), .ZN(n11989) );
  NAND2_X1 U14395 ( .A1(n14507), .A2(n6578), .ZN(n11988) );
  NAND2_X1 U14396 ( .A1(n11989), .A2(n11988), .ZN(n11990) );
  XNOR2_X1 U14397 ( .A(n11990), .B(n11974), .ZN(n11991) );
  AOI22_X1 U14398 ( .A1(n14592), .A2(n12064), .B1(n12077), .B2(n14507), .ZN(
        n14543) );
  INV_X1 U14399 ( .A(n11991), .ZN(n11992) );
  NAND2_X1 U14400 ( .A1(n11993), .A2(n11992), .ZN(n11994) );
  NAND2_X1 U14401 ( .A1(n14184), .A2(n12079), .ZN(n11996) );
  NAND2_X1 U14402 ( .A1(n14546), .A2(n6578), .ZN(n11995) );
  NAND2_X1 U14403 ( .A1(n11996), .A2(n11995), .ZN(n11997) );
  XNOR2_X1 U14404 ( .A(n11997), .B(n11786), .ZN(n11998) );
  AOI22_X1 U14405 ( .A1(n14184), .A2(n12064), .B1(n12077), .B2(n14546), .ZN(
        n11999) );
  XNOR2_X1 U14406 ( .A(n11998), .B(n11999), .ZN(n14506) );
  INV_X1 U14407 ( .A(n11998), .ZN(n12000) );
  NAND2_X1 U14408 ( .A1(n12000), .A2(n11999), .ZN(n12001) );
  NAND2_X1 U14409 ( .A1(n14575), .A2(n12079), .ZN(n12003) );
  NAND2_X1 U14410 ( .A1(n14508), .A2(n6578), .ZN(n12002) );
  NAND2_X1 U14411 ( .A1(n12003), .A2(n12002), .ZN(n12004) );
  XNOR2_X1 U14412 ( .A(n12004), .B(n11974), .ZN(n12005) );
  AOI22_X1 U14413 ( .A1(n14575), .A2(n12064), .B1(n12077), .B2(n14508), .ZN(
        n12006) );
  XNOR2_X1 U14414 ( .A(n12005), .B(n12006), .ZN(n14516) );
  INV_X1 U14415 ( .A(n12005), .ZN(n12007) );
  NAND2_X1 U14416 ( .A1(n12007), .A2(n12006), .ZN(n12008) );
  NAND2_X1 U14417 ( .A1(n12009), .A2(n12008), .ZN(n13860) );
  NAND2_X1 U14418 ( .A1(n14265), .A2(n12079), .ZN(n12011) );
  NAND2_X1 U14419 ( .A1(n14159), .A2(n6578), .ZN(n12010) );
  NAND2_X1 U14420 ( .A1(n12011), .A2(n12010), .ZN(n12012) );
  XNOR2_X1 U14421 ( .A(n12012), .B(n11974), .ZN(n12013) );
  AOI22_X1 U14422 ( .A1(n14265), .A2(n6578), .B1(n12077), .B2(n14159), .ZN(
        n12014) );
  XNOR2_X1 U14423 ( .A(n12013), .B(n12014), .ZN(n13861) );
  INV_X1 U14424 ( .A(n12013), .ZN(n12015) );
  NAND2_X1 U14425 ( .A1(n12015), .A2(n12014), .ZN(n12016) );
  AND2_X1 U14426 ( .A1(n14146), .A2(n12077), .ZN(n12017) );
  AOI21_X1 U14427 ( .B1(n14260), .B2(n12064), .A(n12017), .ZN(n12021) );
  NAND2_X1 U14428 ( .A1(n14260), .A2(n12079), .ZN(n12019) );
  NAND2_X1 U14429 ( .A1(n14146), .A2(n12064), .ZN(n12018) );
  NAND2_X1 U14430 ( .A1(n12019), .A2(n12018), .ZN(n12020) );
  XNOR2_X1 U14431 ( .A(n12020), .B(n11974), .ZN(n12023) );
  XOR2_X1 U14432 ( .A(n12021), .B(n12023), .Z(n13795) );
  INV_X1 U14433 ( .A(n12021), .ZN(n12022) );
  NAND2_X1 U14434 ( .A1(n12023), .A2(n12022), .ZN(n12024) );
  OAI22_X1 U14435 ( .A1(n14252), .A2(n11597), .B1(n13799), .B2(n12034), .ZN(
        n12026) );
  OAI22_X1 U14436 ( .A1(n14252), .A2(n12036), .B1(n13799), .B2(n11597), .ZN(
        n12025) );
  XNOR2_X1 U14437 ( .A(n12025), .B(n11974), .ZN(n12027) );
  XOR2_X1 U14438 ( .A(n12026), .B(n12027), .Z(n13830) );
  NAND2_X1 U14439 ( .A1(n12027), .A2(n12026), .ZN(n12028) );
  AOI22_X1 U14440 ( .A1(n14246), .A2(n12079), .B1(n6578), .B2(n13889), .ZN(
        n12029) );
  XNOR2_X1 U14441 ( .A(n12029), .B(n11974), .ZN(n12032) );
  AOI22_X1 U14442 ( .A1(n14246), .A2(n6578), .B1(n12077), .B2(n13889), .ZN(
        n12031) );
  XNOR2_X1 U14443 ( .A(n12032), .B(n12031), .ZN(n13808) );
  INV_X1 U14444 ( .A(n13808), .ZN(n12030) );
  NAND2_X1 U14445 ( .A1(n12032), .A2(n12031), .ZN(n12033) );
  NAND2_X1 U14446 ( .A1(n13805), .A2(n12033), .ZN(n13851) );
  OAI22_X1 U14447 ( .A1(n14101), .A2(n11597), .B1(n13788), .B2(n12034), .ZN(
        n12039) );
  OAI22_X1 U14448 ( .A1(n14101), .A2(n12036), .B1(n13788), .B2(n11597), .ZN(
        n12037) );
  XNOR2_X1 U14449 ( .A(n12037), .B(n11974), .ZN(n12038) );
  XOR2_X1 U14450 ( .A(n12039), .B(n12038), .Z(n13852) );
  INV_X1 U14451 ( .A(n12038), .ZN(n12041) );
  INV_X1 U14452 ( .A(n12039), .ZN(n12040) );
  NAND2_X1 U14453 ( .A1(n12041), .A2(n12040), .ZN(n12042) );
  NAND2_X1 U14454 ( .A1(n14235), .A2(n12079), .ZN(n12044) );
  NAND2_X1 U14455 ( .A1(n14059), .A2(n12064), .ZN(n12043) );
  NAND2_X1 U14456 ( .A1(n12044), .A2(n12043), .ZN(n12045) );
  XNOR2_X1 U14457 ( .A(n12045), .B(n11974), .ZN(n12046) );
  AOI22_X1 U14458 ( .A1(n14235), .A2(n6578), .B1(n12077), .B2(n14059), .ZN(
        n12047) );
  XNOR2_X1 U14459 ( .A(n12046), .B(n12047), .ZN(n13787) );
  INV_X1 U14460 ( .A(n12046), .ZN(n12048) );
  NAND2_X1 U14461 ( .A1(n14068), .A2(n12079), .ZN(n12050) );
  NAND2_X1 U14462 ( .A1(n13888), .A2(n6577), .ZN(n12049) );
  NAND2_X1 U14463 ( .A1(n12050), .A2(n12049), .ZN(n12051) );
  XNOR2_X1 U14464 ( .A(n12051), .B(n11974), .ZN(n12052) );
  AOI22_X1 U14465 ( .A1(n14068), .A2(n12064), .B1(n12077), .B2(n13888), .ZN(
        n12053) );
  XNOR2_X1 U14466 ( .A(n12052), .B(n12053), .ZN(n13823) );
  NAND2_X1 U14467 ( .A1(n13822), .A2(n13823), .ZN(n12056) );
  INV_X1 U14468 ( .A(n12052), .ZN(n12054) );
  NAND2_X1 U14469 ( .A1(n12054), .A2(n12053), .ZN(n12055) );
  NAND2_X1 U14470 ( .A1(n12056), .A2(n12055), .ZN(n13814) );
  NAND2_X1 U14471 ( .A1(n14221), .A2(n12079), .ZN(n12058) );
  NAND2_X1 U14472 ( .A1(n14058), .A2(n12064), .ZN(n12057) );
  NAND2_X1 U14473 ( .A1(n12058), .A2(n12057), .ZN(n12059) );
  XNOR2_X1 U14474 ( .A(n12059), .B(n11974), .ZN(n12060) );
  AOI22_X1 U14475 ( .A1(n14221), .A2(n6578), .B1(n12077), .B2(n14058), .ZN(
        n12061) );
  XNOR2_X1 U14476 ( .A(n12060), .B(n12061), .ZN(n13815) );
  INV_X1 U14477 ( .A(n12060), .ZN(n12062) );
  NAND2_X1 U14478 ( .A1(n12062), .A2(n12061), .ZN(n12063) );
  NAND2_X1 U14479 ( .A1(n14214), .A2(n12079), .ZN(n12066) );
  NAND2_X1 U14480 ( .A1(n14012), .A2(n12064), .ZN(n12065) );
  NAND2_X1 U14481 ( .A1(n12066), .A2(n12065), .ZN(n12067) );
  XNOR2_X1 U14482 ( .A(n12067), .B(n11974), .ZN(n12068) );
  AOI22_X1 U14483 ( .A1(n14214), .A2(n6577), .B1(n12077), .B2(n14012), .ZN(
        n12069) );
  XNOR2_X1 U14484 ( .A(n12068), .B(n12069), .ZN(n13879) );
  INV_X1 U14485 ( .A(n12068), .ZN(n12070) );
  NAND2_X1 U14486 ( .A1(n14020), .A2(n12079), .ZN(n12072) );
  NAND2_X1 U14487 ( .A1(n13887), .A2(n12064), .ZN(n12071) );
  NAND2_X1 U14488 ( .A1(n12072), .A2(n12071), .ZN(n12073) );
  XNOR2_X1 U14489 ( .A(n12073), .B(n11974), .ZN(n12074) );
  AOI22_X1 U14490 ( .A1(n14020), .A2(n6578), .B1(n12077), .B2(n13887), .ZN(
        n12075) );
  XNOR2_X1 U14491 ( .A(n12074), .B(n12075), .ZN(n13780) );
  INV_X1 U14492 ( .A(n12074), .ZN(n12076) );
  AOI22_X1 U14493 ( .A1(n14203), .A2(n6578), .B1(n12077), .B2(n14011), .ZN(
        n12082) );
  AOI22_X1 U14494 ( .A1(n14203), .A2(n12079), .B1(n6578), .B2(n14011), .ZN(
        n12080) );
  XNOR2_X1 U14495 ( .A(n12080), .B(n11974), .ZN(n12081) );
  XOR2_X1 U14496 ( .A(n12082), .B(n12081), .Z(n12083) );
  AOI22_X1 U14497 ( .A1(n14545), .A2(n13887), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12085) );
  NAND2_X1 U14498 ( .A1(n14547), .A2(n13886), .ZN(n12084) );
  OAI211_X1 U14499 ( .C1(n14554), .C2(n12086), .A(n12085), .B(n12084), .ZN(
        n12087) );
  AOI21_X1 U14500 ( .B1(n14203), .B2(n14536), .A(n12087), .ZN(n12088) );
  OAI21_X1 U14501 ( .B1(n12089), .B2(n14532), .A(n12088), .ZN(P1_U3220) );
  AND2_X1 U14502 ( .A1(n12091), .A2(n12090), .ZN(n12092) );
  NOR2_X2 U14503 ( .A1(n12093), .A2(n12092), .ZN(n12095) );
  XNOR2_X1 U14504 ( .A(n13404), .B(n12116), .ZN(n12096) );
  NOR2_X1 U14505 ( .A1(n12094), .A2(n14465), .ZN(n12977) );
  XNOR2_X1 U14506 ( .A(n13249), .B(n6580), .ZN(n12100) );
  NAND2_X1 U14507 ( .A1(n13067), .A2(n9935), .ZN(n12099) );
  NOR2_X1 U14508 ( .A1(n12100), .A2(n12099), .ZN(n12101) );
  AOI21_X1 U14509 ( .B1(n12100), .B2(n12099), .A(n12101), .ZN(n13009) );
  INV_X1 U14510 ( .A(n12101), .ZN(n12102) );
  NAND2_X1 U14511 ( .A1(n13008), .A2(n12102), .ZN(n12999) );
  XNOR2_X1 U14512 ( .A(n13392), .B(n6580), .ZN(n12104) );
  NAND2_X1 U14513 ( .A1(n13066), .A2(n9935), .ZN(n12103) );
  NOR2_X1 U14514 ( .A1(n12104), .A2(n12103), .ZN(n12105) );
  AOI21_X1 U14515 ( .B1(n12104), .B2(n12103), .A(n12105), .ZN(n13000) );
  XNOR2_X1 U14516 ( .A(n13387), .B(n12116), .ZN(n12108) );
  NAND2_X1 U14517 ( .A1(n13065), .A2(n9935), .ZN(n12106) );
  XNOR2_X1 U14518 ( .A(n12108), .B(n12106), .ZN(n13052) );
  INV_X1 U14519 ( .A(n12106), .ZN(n12107) );
  INV_X1 U14520 ( .A(n12965), .ZN(n12113) );
  XNOR2_X1 U14521 ( .A(n13202), .B(n6580), .ZN(n12111) );
  NOR2_X1 U14522 ( .A1(n13053), .A2(n14465), .ZN(n12110) );
  NAND2_X1 U14523 ( .A1(n12111), .A2(n12110), .ZN(n12114) );
  OAI21_X1 U14524 ( .B1(n12111), .B2(n12110), .A(n12114), .ZN(n12964) );
  INV_X1 U14525 ( .A(n12964), .ZN(n12112) );
  NAND2_X1 U14526 ( .A1(n12966), .A2(n12114), .ZN(n12119) );
  NAND2_X1 U14527 ( .A1(n13063), .A2(n9935), .ZN(n12115) );
  XOR2_X1 U14528 ( .A(n12116), .B(n12115), .Z(n12117) );
  XNOR2_X1 U14529 ( .A(n13459), .B(n12117), .ZN(n12118) );
  XNOR2_X1 U14530 ( .A(n12119), .B(n12118), .ZN(n12126) );
  OR2_X1 U14531 ( .A1(n12120), .A2(n14443), .ZN(n12122) );
  OR2_X1 U14532 ( .A1(n13053), .A2(n14441), .ZN(n12121) );
  NAND2_X1 U14533 ( .A1(n12122), .A2(n12121), .ZN(n13183) );
  AOI22_X1 U14534 ( .A1(n14450), .A2(n13183), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12123) );
  OAI21_X1 U14535 ( .B1(n13185), .B2(n14453), .A(n12123), .ZN(n12124) );
  AOI21_X1 U14536 ( .B1(n7104), .B2(n14451), .A(n12124), .ZN(n12125) );
  OAI21_X1 U14537 ( .B1(n12126), .B2(n13059), .A(n12125), .ZN(P2_U3192) );
  XNOR2_X1 U14538 ( .A(n12836), .B(n12200), .ZN(n12197) );
  XNOR2_X1 U14539 ( .A(n12197), .B(n12514), .ZN(n12198) );
  INV_X1 U14540 ( .A(n12129), .ZN(n12130) );
  XNOR2_X1 U14541 ( .A(n12948), .B(n12200), .ZN(n12171) );
  INV_X1 U14542 ( .A(n12171), .ZN(n12131) );
  NAND2_X1 U14543 ( .A1(n12131), .A2(n12806), .ZN(n12132) );
  XNOR2_X1 U14544 ( .A(n12944), .B(n12200), .ZN(n12134) );
  XNOR2_X1 U14545 ( .A(n12134), .B(n12791), .ZN(n12286) );
  INV_X1 U14546 ( .A(n12286), .ZN(n12133) );
  NAND2_X1 U14547 ( .A1(n12134), .A2(n12791), .ZN(n12135) );
  XNOR2_X1 U14548 ( .A(n12884), .B(n12200), .ZN(n12136) );
  XNOR2_X1 U14549 ( .A(n12136), .B(n12516), .ZN(n12225) );
  INV_X1 U14550 ( .A(n12136), .ZN(n12137) );
  NAND2_X1 U14551 ( .A1(n12137), .A2(n12516), .ZN(n12138) );
  NAND2_X1 U14552 ( .A1(n12224), .A2(n12138), .ZN(n12234) );
  XNOR2_X1 U14553 ( .A(n12939), .B(n12200), .ZN(n12139) );
  XNOR2_X1 U14554 ( .A(n12139), .B(n12228), .ZN(n12233) );
  NAND2_X1 U14555 ( .A1(n12234), .A2(n12233), .ZN(n12232) );
  NAND2_X1 U14556 ( .A1(n12139), .A2(n12792), .ZN(n12140) );
  NAND2_X1 U14557 ( .A1(n12232), .A2(n12140), .ZN(n12272) );
  XNOR2_X1 U14558 ( .A(n12765), .B(n12200), .ZN(n12141) );
  XNOR2_X1 U14559 ( .A(n12141), .B(n12751), .ZN(n12271) );
  NAND2_X1 U14560 ( .A1(n12272), .A2(n12271), .ZN(n12270) );
  INV_X1 U14561 ( .A(n12141), .ZN(n12142) );
  NAND2_X1 U14562 ( .A1(n12142), .A2(n12751), .ZN(n12143) );
  NAND2_X1 U14563 ( .A1(n12270), .A2(n12143), .ZN(n12192) );
  XNOR2_X1 U14564 ( .A(n12189), .B(n12200), .ZN(n12144) );
  XNOR2_X1 U14565 ( .A(n12144), .B(n12763), .ZN(n12191) );
  INV_X1 U14566 ( .A(n12144), .ZN(n12145) );
  NAND2_X1 U14567 ( .A1(n12145), .A2(n12763), .ZN(n12146) );
  XNOR2_X1 U14568 ( .A(n12253), .B(n12200), .ZN(n12147) );
  XNOR2_X1 U14569 ( .A(n12147), .B(n12752), .ZN(n12255) );
  INV_X1 U14570 ( .A(n12147), .ZN(n12148) );
  NAND2_X1 U14571 ( .A1(n12148), .A2(n12752), .ZN(n12149) );
  XNOR2_X1 U14572 ( .A(n12209), .B(n12200), .ZN(n12150) );
  XNOR2_X1 U14573 ( .A(n12150), .B(n12515), .ZN(n12211) );
  INV_X1 U14574 ( .A(n12150), .ZN(n12151) );
  NAND2_X1 U14575 ( .A1(n12151), .A2(n12515), .ZN(n12152) );
  XNOR2_X1 U14576 ( .A(n12720), .B(n12200), .ZN(n12153) );
  XNOR2_X2 U14577 ( .A(n12155), .B(n12153), .ZN(n12263) );
  INV_X1 U14578 ( .A(n12153), .ZN(n12154) );
  NOR2_X1 U14579 ( .A1(n12155), .A2(n12154), .ZN(n12156) );
  XNOR2_X1 U14580 ( .A(n12849), .B(n12200), .ZN(n12245) );
  XNOR2_X1 U14581 ( .A(n12705), .B(n12157), .ZN(n12241) );
  INV_X1 U14582 ( .A(n12241), .ZN(n12158) );
  OAI22_X1 U14583 ( .A1(n12245), .A2(n12244), .B1(n12717), .B2(n12158), .ZN(
        n12162) );
  OAI21_X1 U14584 ( .B1(n12241), .B2(n12687), .A(n12702), .ZN(n12160) );
  NOR2_X1 U14585 ( .A1(n12702), .A2(n12687), .ZN(n12159) );
  AOI22_X1 U14586 ( .A1(n12245), .A2(n12160), .B1(n12159), .B2(n12158), .ZN(
        n12161) );
  XNOR2_X1 U14587 ( .A(n12845), .B(n12200), .ZN(n12163) );
  XNOR2_X1 U14588 ( .A(n12163), .B(n12688), .ZN(n12218) );
  XNOR2_X1 U14589 ( .A(n12840), .B(n12200), .ZN(n12164) );
  XNOR2_X1 U14590 ( .A(n12164), .B(n12636), .ZN(n12278) );
  INV_X1 U14591 ( .A(n12164), .ZN(n12165) );
  XOR2_X1 U14592 ( .A(n12198), .B(n12199), .Z(n12170) );
  AOI22_X1 U14593 ( .A1(n12644), .A2(n12295), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12167) );
  NAND2_X1 U14594 ( .A1(n12670), .A2(n12291), .ZN(n12166) );
  OAI211_X1 U14595 ( .C1(n12637), .C2(n12293), .A(n12167), .B(n12166), .ZN(
        n12168) );
  AOI21_X1 U14596 ( .B1(n12836), .B2(n12282), .A(n12168), .ZN(n12169) );
  OAI21_X1 U14597 ( .B1(n12170), .B2(n12285), .A(n12169), .ZN(P3_U3154) );
  XNOR2_X1 U14598 ( .A(n12171), .B(n12806), .ZN(n12172) );
  XNOR2_X1 U14599 ( .A(n12173), .B(n12172), .ZN(n12183) );
  INV_X1 U14600 ( .A(n12948), .ZN(n12181) );
  INV_X1 U14601 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12174) );
  NOR2_X1 U14602 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12174), .ZN(n15214) );
  NOR2_X1 U14603 ( .A1(n12293), .A2(n12175), .ZN(n12176) );
  AOI211_X1 U14604 ( .C1(n12291), .C2(n12518), .A(n15214), .B(n12176), .ZN(
        n12177) );
  OAI21_X1 U14605 ( .B1(n12179), .B2(n12178), .A(n12177), .ZN(n12180) );
  AOI21_X1 U14606 ( .B1(n12181), .B2(n12282), .A(n12180), .ZN(n12182) );
  OAI21_X1 U14607 ( .B1(n12183), .B2(n12285), .A(n12182), .ZN(P3_U3155) );
  XNOR2_X1 U14608 ( .A(n12242), .B(n12241), .ZN(n12243) );
  XNOR2_X1 U14609 ( .A(n12243), .B(n12717), .ZN(n12188) );
  AOI22_X1 U14610 ( .A1(n12701), .A2(n12291), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12185) );
  NAND2_X1 U14611 ( .A1(n12710), .A2(n12295), .ZN(n12184) );
  OAI211_X1 U14612 ( .C1(n12244), .C2(n12293), .A(n12185), .B(n12184), .ZN(
        n12186) );
  AOI21_X1 U14613 ( .B1(n12705), .B2(n12282), .A(n12186), .ZN(n12187) );
  OAI21_X1 U14614 ( .B1(n12188), .B2(n12285), .A(n12187), .ZN(P3_U3156) );
  INV_X1 U14615 ( .A(n12189), .ZN(n12934) );
  OAI211_X1 U14616 ( .C1(n12192), .C2(n12191), .A(n12190), .B(n12269), .ZN(
        n12196) );
  NAND2_X1 U14617 ( .A1(n12291), .A2(n12751), .ZN(n12193) );
  NAND2_X1 U14618 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12605)
         );
  OAI211_X1 U14619 ( .C1(n12730), .C2(n12293), .A(n12193), .B(n12605), .ZN(
        n12194) );
  AOI21_X1 U14620 ( .B1(n12756), .B2(n12295), .A(n12194), .ZN(n12195) );
  OAI211_X1 U14621 ( .C1(n12934), .C2(n12298), .A(n12196), .B(n12195), .ZN(
        P3_U3159) );
  AOI22_X1 U14622 ( .A1(n12199), .A2(n12198), .B1(n12654), .B2(n12197), .ZN(
        n12202) );
  XNOR2_X1 U14623 ( .A(n12497), .B(n12200), .ZN(n12201) );
  XNOR2_X1 U14624 ( .A(n12202), .B(n12201), .ZN(n12208) );
  NAND2_X1 U14625 ( .A1(n12514), .A2(n12291), .ZN(n12204) );
  AOI22_X1 U14626 ( .A1(n12626), .A2(n12295), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12203) );
  OAI211_X1 U14627 ( .C1(n12205), .C2(n12293), .A(n12204), .B(n12203), .ZN(
        n12206) );
  AOI21_X1 U14628 ( .B1(n12324), .B2(n12282), .A(n12206), .ZN(n12207) );
  OAI21_X1 U14629 ( .B1(n12208), .B2(n12285), .A(n12207), .ZN(P3_U3160) );
  OAI211_X1 U14630 ( .C1(n12212), .C2(n12211), .A(n12210), .B(n12269), .ZN(
        n12216) );
  AOI22_X1 U14631 ( .A1(n12752), .A2(n12291), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12213) );
  OAI21_X1 U14632 ( .B1(n12731), .B2(n12293), .A(n12213), .ZN(n12214) );
  AOI21_X1 U14633 ( .B1(n12734), .B2(n12295), .A(n12214), .ZN(n12215) );
  OAI211_X1 U14634 ( .C1(n12926), .C2(n12298), .A(n12216), .B(n12215), .ZN(
        P3_U3163) );
  XOR2_X1 U14635 ( .A(n12218), .B(n12217), .Z(n12223) );
  AOI22_X1 U14636 ( .A1(n12702), .A2(n12291), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12220) );
  NAND2_X1 U14637 ( .A1(n12675), .A2(n12295), .ZN(n12219) );
  OAI211_X1 U14638 ( .C1(n12636), .C2(n12293), .A(n12220), .B(n12219), .ZN(
        n12221) );
  AOI21_X1 U14639 ( .B1(n12845), .B2(n12282), .A(n12221), .ZN(n12222) );
  OAI21_X1 U14640 ( .B1(n12223), .B2(n12285), .A(n12222), .ZN(P3_U3165) );
  INV_X1 U14641 ( .A(n12884), .ZN(n12801) );
  OAI211_X1 U14642 ( .C1(n12226), .C2(n12225), .A(n12224), .B(n12269), .ZN(
        n12231) );
  NAND2_X1 U14643 ( .A1(n12291), .A2(n12791), .ZN(n12227) );
  NAND2_X1 U14644 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n14373)
         );
  OAI211_X1 U14645 ( .C1(n12293), .C2(n12228), .A(n12227), .B(n14373), .ZN(
        n12229) );
  AOI21_X1 U14646 ( .B1(n12799), .B2(n12295), .A(n12229), .ZN(n12230) );
  OAI211_X1 U14647 ( .C1(n12801), .C2(n12298), .A(n12231), .B(n12230), .ZN(
        P3_U3166) );
  OAI211_X1 U14648 ( .C1(n12234), .C2(n12233), .A(n12232), .B(n12269), .ZN(
        n12240) );
  NOR2_X1 U14649 ( .A1(n12235), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14401) );
  AOI21_X1 U14650 ( .B1(n12236), .B2(n12751), .A(n14401), .ZN(n12237) );
  OAI21_X1 U14651 ( .B1(n12807), .B2(n12257), .A(n12237), .ZN(n12238) );
  AOI21_X1 U14652 ( .B1(n12785), .B2(n12295), .A(n12238), .ZN(n12239) );
  OAI211_X1 U14653 ( .C1(n12298), .C2(n12939), .A(n12240), .B(n12239), .ZN(
        P3_U3168) );
  OAI22_X1 U14654 ( .A1(n12243), .A2(n12687), .B1(n12242), .B2(n12241), .ZN(
        n12247) );
  XNOR2_X1 U14655 ( .A(n12245), .B(n12244), .ZN(n12246) );
  XNOR2_X1 U14656 ( .A(n12247), .B(n12246), .ZN(n12252) );
  AOI22_X1 U14657 ( .A1(n12687), .A2(n12291), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12249) );
  NAND2_X1 U14658 ( .A1(n12691), .A2(n12295), .ZN(n12248) );
  OAI211_X1 U14659 ( .C1(n12653), .C2(n12293), .A(n12249), .B(n12248), .ZN(
        n12250) );
  AOI21_X1 U14660 ( .B1(n12849), .B2(n12282), .A(n12250), .ZN(n12251) );
  OAI21_X1 U14661 ( .B1(n12252), .B2(n12285), .A(n12251), .ZN(P3_U3169) );
  OAI211_X1 U14662 ( .C1(n12256), .C2(n12255), .A(n12254), .B(n12269), .ZN(
        n12262) );
  NOR2_X1 U14663 ( .A1(n12257), .A2(n12741), .ZN(n12260) );
  OAI22_X1 U14664 ( .A1(n12742), .A2(n12293), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12258), .ZN(n12259) );
  AOI211_X1 U14665 ( .C1(n12745), .C2(n12295), .A(n12260), .B(n12259), .ZN(
        n12261) );
  OAI211_X1 U14666 ( .C1(n12930), .C2(n12298), .A(n12262), .B(n12261), .ZN(
        P3_U3173) );
  XNOR2_X1 U14667 ( .A(n12263), .B(n12701), .ZN(n12268) );
  AOI22_X1 U14668 ( .A1(n12515), .A2(n12291), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12265) );
  NAND2_X1 U14669 ( .A1(n12295), .A2(n12721), .ZN(n12264) );
  OAI211_X1 U14670 ( .C1(n12717), .C2(n12293), .A(n12265), .B(n12264), .ZN(
        n12266) );
  AOI21_X1 U14671 ( .B1(n12720), .B2(n12282), .A(n12266), .ZN(n12267) );
  OAI21_X1 U14672 ( .B1(n12268), .B2(n12285), .A(n12267), .ZN(P3_U3175) );
  INV_X1 U14673 ( .A(n12765), .ZN(n12277) );
  OAI211_X1 U14674 ( .C1(n12272), .C2(n12271), .A(n12270), .B(n12269), .ZN(
        n12276) );
  NAND2_X1 U14675 ( .A1(n12291), .A2(n12792), .ZN(n12273) );
  NAND2_X1 U14676 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n14417)
         );
  OAI211_X1 U14677 ( .C1(n12293), .C2(n12741), .A(n12273), .B(n14417), .ZN(
        n12274) );
  AOI21_X1 U14678 ( .B1(n12766), .B2(n12295), .A(n12274), .ZN(n12275) );
  OAI211_X1 U14679 ( .C1(n12277), .C2(n12298), .A(n12276), .B(n12275), .ZN(
        P3_U3178) );
  AOI22_X1 U14680 ( .A1(n12658), .A2(n12295), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12280) );
  NAND2_X1 U14681 ( .A1(n12688), .A2(n12291), .ZN(n12279) );
  OAI211_X1 U14682 ( .C1(n12654), .C2(n12293), .A(n12280), .B(n12279), .ZN(
        n12281) );
  AOI21_X1 U14683 ( .B1(n12840), .B2(n12282), .A(n12281), .ZN(n12283) );
  OAI21_X1 U14684 ( .B1(n12284), .B2(n12285), .A(n12283), .ZN(P3_U3180) );
  AOI21_X1 U14685 ( .B1(n12287), .B2(n12286), .A(n12285), .ZN(n12289) );
  NAND2_X1 U14686 ( .A1(n12289), .A2(n12288), .ZN(n12297) );
  INV_X1 U14687 ( .A(n12290), .ZN(n12810) );
  NAND2_X1 U14688 ( .A1(n12291), .A2(n12517), .ZN(n12292) );
  NAND2_X1 U14689 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n14355)
         );
  OAI211_X1 U14690 ( .C1(n12293), .C2(n12807), .A(n12292), .B(n14355), .ZN(
        n12294) );
  AOI21_X1 U14691 ( .B1(n12810), .B2(n12295), .A(n12294), .ZN(n12296) );
  OAI211_X1 U14692 ( .C1(n12298), .C2(n12944), .A(n12297), .B(n12296), .ZN(
        P3_U3181) );
  NAND2_X1 U14693 ( .A1(n12299), .A2(n12318), .ZN(n12301) );
  NAND2_X1 U14694 ( .A1(n12319), .A2(SI_30_), .ZN(n12300) );
  INV_X1 U14695 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12307) );
  NAND2_X1 U14696 ( .A1(n12302), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12306) );
  INV_X1 U14697 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12303) );
  OR2_X1 U14698 ( .A1(n12304), .A2(n12303), .ZN(n12305) );
  OAI211_X1 U14699 ( .C1(n12307), .C2(n9304), .A(n12306), .B(n12305), .ZN(
        n12308) );
  INV_X1 U14700 ( .A(n12308), .ZN(n12309) );
  NOR2_X1 U14701 ( .A1(n12901), .A2(n12466), .ZN(n12470) );
  NOR2_X1 U14702 ( .A1(n12312), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12314) );
  OAI22_X1 U14703 ( .A1(n12315), .A2(n12314), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n12313), .ZN(n12317) );
  XNOR2_X1 U14704 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12316) );
  XNOR2_X1 U14705 ( .A(n12317), .B(n12316), .ZN(n12953) );
  NAND2_X1 U14706 ( .A1(n12953), .A2(n12318), .ZN(n12321) );
  NAND2_X1 U14707 ( .A1(n12319), .A2(SI_31_), .ZN(n12320) );
  OR2_X1 U14708 ( .A1(n12324), .A2(n12637), .ZN(n12452) );
  INV_X1 U14709 ( .A(n12452), .ZN(n12456) );
  XNOR2_X1 U14710 ( .A(n12325), .B(n12473), .ZN(n12326) );
  NOR2_X1 U14711 ( .A1(n12327), .A2(n12326), .ZN(n12331) );
  OR2_X1 U14712 ( .A1(n12845), .A2(n12653), .ZN(n12329) );
  MUX2_X1 U14713 ( .A(n12329), .B(n12328), .S(n12448), .Z(n12330) );
  OAI21_X1 U14714 ( .B1(n12331), .B2(n12669), .A(n12330), .ZN(n12446) );
  NAND2_X1 U14715 ( .A1(n12449), .A2(n12457), .ZN(n12652) );
  INV_X1 U14716 ( .A(n12652), .ZN(n12649) );
  MUX2_X1 U14717 ( .A(n12332), .B(n12333), .S(n12473), .Z(n12441) );
  MUX2_X1 U14718 ( .A(n12335), .B(n12334), .S(n12473), .Z(n12439) );
  OAI21_X1 U14719 ( .B1(n12823), .B2(n12338), .A(n12341), .ZN(n12336) );
  MUX2_X1 U14720 ( .A(n12337), .B(n12336), .S(n12473), .Z(n12351) );
  INV_X1 U14721 ( .A(n12338), .ZN(n12339) );
  OAI22_X1 U14722 ( .A1(n12822), .A2(n12340), .B1(n12509), .B2(n12339), .ZN(
        n12342) );
  NAND2_X1 U14723 ( .A1(n12342), .A2(n12341), .ZN(n12343) );
  NAND2_X1 U14724 ( .A1(n12343), .A2(n15317), .ZN(n12350) );
  NAND2_X1 U14725 ( .A1(n15286), .A2(n12344), .ZN(n12347) );
  NAND2_X1 U14726 ( .A1(n12352), .A2(n12345), .ZN(n12346) );
  MUX2_X1 U14727 ( .A(n12347), .B(n12346), .S(n12473), .Z(n12348) );
  INV_X1 U14728 ( .A(n12348), .ZN(n12349) );
  OAI21_X1 U14729 ( .B1(n12351), .B2(n12350), .A(n12349), .ZN(n12354) );
  INV_X1 U14730 ( .A(n15290), .ZN(n15288) );
  MUX2_X1 U14731 ( .A(n15286), .B(n12352), .S(n12448), .Z(n12353) );
  NAND3_X1 U14732 ( .A1(n12354), .A2(n15288), .A3(n12353), .ZN(n12359) );
  MUX2_X1 U14733 ( .A(n12356), .B(n12355), .S(n12473), .Z(n12357) );
  NAND3_X1 U14734 ( .A1(n12359), .A2(n12358), .A3(n12357), .ZN(n12365) );
  NAND2_X1 U14735 ( .A1(n15276), .A2(n12360), .ZN(n12361) );
  NAND2_X1 U14736 ( .A1(n12367), .A2(n12361), .ZN(n12362) );
  NAND2_X1 U14737 ( .A1(n12362), .A2(n12448), .ZN(n12364) );
  AOI21_X1 U14738 ( .B1(n12365), .B2(n12364), .A(n12363), .ZN(n12371) );
  AOI21_X1 U14739 ( .B1(n12366), .B2(n15271), .A(n12448), .ZN(n12370) );
  INV_X1 U14740 ( .A(n12367), .ZN(n12368) );
  NAND2_X1 U14741 ( .A1(n12368), .A2(n12473), .ZN(n12369) );
  OAI211_X1 U14742 ( .C1(n12371), .C2(n12370), .A(n15262), .B(n12369), .ZN(
        n12375) );
  MUX2_X1 U14743 ( .A(n12373), .B(n12372), .S(n12473), .Z(n12374) );
  NAND3_X1 U14744 ( .A1(n12375), .A2(n15242), .A3(n12374), .ZN(n12379) );
  NAND2_X1 U14745 ( .A1(n12522), .A2(n15251), .ZN(n12376) );
  MUX2_X1 U14746 ( .A(n12377), .B(n12376), .S(n12473), .Z(n12378) );
  NAND3_X1 U14747 ( .A1(n12379), .A2(n12482), .A3(n12378), .ZN(n12383) );
  MUX2_X1 U14748 ( .A(n12381), .B(n12380), .S(n12473), .Z(n12382) );
  NAND2_X1 U14749 ( .A1(n12383), .A2(n12382), .ZN(n12388) );
  INV_X1 U14750 ( .A(n15232), .ZN(n12486) );
  MUX2_X1 U14751 ( .A(n12385), .B(n12384), .S(n12473), .Z(n12386) );
  NAND2_X1 U14752 ( .A1(n12386), .A2(n14422), .ZN(n12387) );
  AOI21_X1 U14753 ( .B1(n12388), .B2(n12486), .A(n12387), .ZN(n12398) );
  NAND2_X1 U14754 ( .A1(n12394), .A2(n12389), .ZN(n12392) );
  NAND2_X1 U14755 ( .A1(n12393), .A2(n12390), .ZN(n12391) );
  MUX2_X1 U14756 ( .A(n12392), .B(n12391), .S(n12448), .Z(n12397) );
  MUX2_X1 U14757 ( .A(n12394), .B(n12393), .S(n12473), .Z(n12395) );
  OAI211_X1 U14758 ( .C1(n12398), .C2(n12397), .A(n12396), .B(n12395), .ZN(
        n12403) );
  INV_X1 U14759 ( .A(n12489), .ZN(n12402) );
  MUX2_X1 U14760 ( .A(n12400), .B(n12399), .S(n12448), .Z(n12401) );
  NAND3_X1 U14761 ( .A1(n12403), .A2(n12402), .A3(n12401), .ZN(n12407) );
  MUX2_X1 U14762 ( .A(n12405), .B(n12404), .S(n12448), .Z(n12406) );
  NAND2_X1 U14763 ( .A1(n12407), .A2(n12406), .ZN(n12408) );
  NAND2_X1 U14764 ( .A1(n12408), .A2(n12808), .ZN(n12413) );
  NAND2_X1 U14765 ( .A1(n12414), .A2(n12409), .ZN(n12410) );
  NAND2_X1 U14766 ( .A1(n12410), .A2(n12448), .ZN(n12412) );
  INV_X1 U14767 ( .A(n12782), .ZN(n12411) );
  AOI21_X1 U14768 ( .B1(n12413), .B2(n12412), .A(n12411), .ZN(n12416) );
  AOI21_X1 U14769 ( .B1(n12782), .B2(n12794), .A(n12448), .ZN(n12415) );
  OAI22_X1 U14770 ( .A1(n12416), .A2(n12415), .B1(n12448), .B2(n12414), .ZN(
        n12417) );
  INV_X1 U14771 ( .A(n12779), .ZN(n12783) );
  NAND3_X1 U14772 ( .A1(n12417), .A2(n12783), .A3(n12492), .ZN(n12428) );
  INV_X1 U14773 ( .A(n12422), .ZN(n12419) );
  OAI211_X1 U14774 ( .C1(n12419), .C2(n12773), .A(n12429), .B(n12418), .ZN(
        n12425) );
  INV_X1 U14775 ( .A(n12420), .ZN(n12421) );
  NAND2_X1 U14776 ( .A1(n12492), .A2(n12421), .ZN(n12423) );
  NAND3_X1 U14777 ( .A1(n12423), .A2(n12422), .A3(n12430), .ZN(n12424) );
  MUX2_X1 U14778 ( .A(n12425), .B(n12424), .S(n12448), .Z(n12426) );
  INV_X1 U14779 ( .A(n12426), .ZN(n12427) );
  NAND2_X1 U14780 ( .A1(n12428), .A2(n12427), .ZN(n12433) );
  INV_X1 U14781 ( .A(n12744), .ZN(n12432) );
  MUX2_X1 U14782 ( .A(n12430), .B(n12429), .S(n12448), .Z(n12431) );
  NAND3_X1 U14783 ( .A1(n12433), .A2(n12432), .A3(n12431), .ZN(n12437) );
  MUX2_X1 U14784 ( .A(n12435), .B(n12434), .S(n12473), .Z(n12436) );
  NAND3_X1 U14785 ( .A1(n12437), .A2(n12732), .A3(n12436), .ZN(n12438) );
  NAND3_X1 U14786 ( .A1(n12718), .A2(n12439), .A3(n12438), .ZN(n12440) );
  NAND3_X1 U14787 ( .A1(n12706), .A2(n12441), .A3(n12440), .ZN(n12443) );
  NAND3_X1 U14788 ( .A1(n12705), .A2(n12717), .A3(n12473), .ZN(n12442) );
  AND2_X1 U14789 ( .A1(n12443), .A2(n12442), .ZN(n12444) );
  OR3_X1 U14790 ( .A1(n12669), .A2(n12686), .A3(n12444), .ZN(n12445) );
  NAND3_X1 U14791 ( .A1(n12446), .A2(n12649), .A3(n12445), .ZN(n12447) );
  INV_X1 U14792 ( .A(n12450), .ZN(n12451) );
  NAND2_X1 U14793 ( .A1(n12452), .A2(n12451), .ZN(n12454) );
  INV_X1 U14794 ( .A(n12457), .ZN(n12459) );
  OR3_X1 U14795 ( .A1(n12836), .A2(n12654), .A3(n12473), .ZN(n12458) );
  OAI21_X1 U14796 ( .B1(n12460), .B2(n12459), .A(n12458), .ZN(n12461) );
  AND2_X1 U14797 ( .A1(n12461), .A2(n12497), .ZN(n12463) );
  INV_X1 U14798 ( .A(n12462), .ZN(n12499) );
  MUX2_X1 U14799 ( .A(n12465), .B(n12464), .S(n12473), .Z(n12468) );
  XNOR2_X1 U14800 ( .A(n12901), .B(n12466), .ZN(n12501) );
  INV_X1 U14801 ( .A(n12501), .ZN(n12467) );
  INV_X1 U14802 ( .A(n12470), .ZN(n12471) );
  AND2_X1 U14803 ( .A1(n12897), .A2(n12612), .ZN(n12475) );
  INV_X1 U14804 ( .A(n12612), .ZN(n12513) );
  XOR2_X1 U14805 ( .A(n12513), .B(n12897), .Z(n12502) );
  NAND4_X1 U14806 ( .A1(n12480), .A2(n15272), .A3(n15262), .A4(n12479), .ZN(
        n12484) );
  INV_X1 U14807 ( .A(n12823), .ZN(n12481) );
  NAND4_X1 U14808 ( .A1(n12482), .A2(n12481), .A3(n15317), .A4(n15288), .ZN(
        n12483) );
  NOR4_X1 U14809 ( .A1(n15246), .A2(n12484), .A3(n12483), .A4(n9323), .ZN(
        n12487) );
  NAND4_X1 U14810 ( .A1(n12487), .A2(n12486), .A3(n14422), .A4(n12485), .ZN(
        n12488) );
  NOR4_X1 U14811 ( .A1(n12491), .A2(n12490), .A3(n12489), .A4(n12488), .ZN(
        n12493) );
  NAND4_X1 U14812 ( .A1(n12493), .A2(n12492), .A3(n12783), .A4(n12808), .ZN(
        n12494) );
  NOR3_X1 U14813 ( .A1(n12744), .A2(n7537), .A3(n12494), .ZN(n12495) );
  NAND4_X1 U14814 ( .A1(n12706), .A2(n12718), .A3(n12732), .A4(n12495), .ZN(
        n12496) );
  NOR4_X1 U14815 ( .A1(n12652), .A2(n12669), .A3(n12686), .A4(n12496), .ZN(
        n12498) );
  NAND4_X1 U14816 ( .A1(n12499), .A2(n12640), .A3(n12498), .A4(n12497), .ZN(
        n12500) );
  NOR3_X1 U14817 ( .A1(n12502), .A2(n12501), .A3(n12500), .ZN(n12503) );
  XNOR2_X1 U14818 ( .A(n12503), .B(n12608), .ZN(n12504) );
  NOR3_X1 U14819 ( .A1(n12508), .A2(n12600), .A3(n12507), .ZN(n12511) );
  OAI21_X1 U14820 ( .B1(n12512), .B2(n12509), .A(P3_B_REG_SCAN_IN), .ZN(n12510) );
  MUX2_X1 U14821 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12513), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14822 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12514), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14823 ( .A(n12670), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12526), .Z(
        P3_U3517) );
  MUX2_X1 U14824 ( .A(n12688), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12526), .Z(
        P3_U3516) );
  MUX2_X1 U14825 ( .A(n12687), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12526), .Z(
        P3_U3514) );
  MUX2_X1 U14826 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12701), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14827 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12515), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14828 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12752), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14829 ( .A(n12763), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12526), .Z(
        P3_U3510) );
  MUX2_X1 U14830 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12751), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14831 ( .A(n12792), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12526), .Z(
        P3_U3508) );
  MUX2_X1 U14832 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12516), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14833 ( .A(n12791), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12526), .Z(
        P3_U3506) );
  MUX2_X1 U14834 ( .A(n12517), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12526), .Z(
        P3_U3505) );
  MUX2_X1 U14835 ( .A(n12518), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12526), .Z(
        P3_U3504) );
  MUX2_X1 U14836 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12519), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14837 ( .A(n12520), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12526), .Z(
        P3_U3502) );
  MUX2_X1 U14838 ( .A(n12521), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12526), .Z(
        P3_U3501) );
  MUX2_X1 U14839 ( .A(n15247), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12526), .Z(
        P3_U3500) );
  MUX2_X1 U14840 ( .A(n12522), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12526), .Z(
        P3_U3499) );
  MUX2_X1 U14841 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n15277), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14842 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12523), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14843 ( .A(n15276), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12526), .Z(
        P3_U3496) );
  MUX2_X1 U14844 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12524), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14845 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n9277), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14846 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12525), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14847 ( .A(n10491), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12526), .Z(
        P3_U3492) );
  MUX2_X1 U14848 ( .A(n12817), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12526), .Z(
        P3_U3491) );
  AOI22_X1 U14849 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n12597), .B1(n14404), 
        .B2(n12563), .ZN(n14407) );
  AOI22_X1 U14850 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12590), .B1(n14372), 
        .B2(n12541), .ZN(n14371) );
  NAND2_X1 U14851 ( .A1(n15217), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12584) );
  INV_X1 U14852 ( .A(n15217), .ZN(n12527) );
  INV_X1 U14853 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12894) );
  NAND2_X1 U14854 ( .A1(n12527), .A2(n12894), .ZN(n12528) );
  AND2_X1 U14855 ( .A1(n12528), .A2(n12584), .ZN(n15213) );
  NAND2_X1 U14856 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n15181), .ZN(n12536) );
  AOI22_X1 U14857 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n15181), .B1(n12529), 
        .B2(n9450), .ZN(n15178) );
  INV_X1 U14858 ( .A(n12571), .ZN(n15150) );
  INV_X1 U14859 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15393) );
  OAI21_X1 U14860 ( .B1(n12531), .B2(n15389), .A(n12530), .ZN(n12532) );
  NAND2_X1 U14861 ( .A1(n15124), .A2(n12532), .ZN(n12533) );
  NAND2_X1 U14862 ( .A1(n12533), .A2(n15128), .ZN(n15136) );
  MUX2_X1 U14863 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n15393), .S(n12571), .Z(
        n15135) );
  NAND2_X1 U14864 ( .A1(n15136), .A2(n15135), .ZN(n15134) );
  OAI21_X1 U14865 ( .B1(n15150), .B2(n15393), .A(n15134), .ZN(n12534) );
  NAND2_X1 U14866 ( .A1(n15163), .A2(n12534), .ZN(n12535) );
  NAND2_X1 U14867 ( .A1(n12535), .A2(n15159), .ZN(n15177) );
  NAND2_X1 U14868 ( .A1(n15178), .A2(n15177), .ZN(n15176) );
  NAND2_X1 U14869 ( .A1(n15199), .A2(n12537), .ZN(n12538) );
  NAND2_X1 U14870 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n15196), .ZN(n15195) );
  NAND2_X1 U14871 ( .A1(n12538), .A2(n15195), .ZN(n15212) );
  NAND2_X1 U14872 ( .A1(n15213), .A2(n15212), .ZN(n15211) );
  NAND2_X1 U14873 ( .A1(n12584), .A2(n15211), .ZN(n12539) );
  NAND2_X1 U14874 ( .A1(n14328), .A2(n12539), .ZN(n12540) );
  XNOR2_X1 U14875 ( .A(n12554), .B(n12539), .ZN(n14354) );
  NAND2_X1 U14876 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n14354), .ZN(n14353) );
  NAND2_X1 U14877 ( .A1(n12540), .A2(n14353), .ZN(n14370) );
  NAND2_X1 U14878 ( .A1(n14371), .A2(n14370), .ZN(n14369) );
  OAI21_X1 U14879 ( .B1(n14372), .B2(n12541), .A(n14369), .ZN(n12542) );
  NAND2_X1 U14880 ( .A1(n14397), .A2(n12542), .ZN(n12543) );
  INV_X1 U14881 ( .A(n14397), .ZN(n12594) );
  XNOR2_X1 U14882 ( .A(n12542), .B(n12594), .ZN(n14391) );
  NAND2_X1 U14883 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14391), .ZN(n14390) );
  NAND2_X1 U14884 ( .A1(n12543), .A2(n14390), .ZN(n14406) );
  NAND2_X1 U14885 ( .A1(n14407), .A2(n14406), .ZN(n14405) );
  INV_X1 U14886 ( .A(n15124), .ZN(n12568) );
  XNOR2_X1 U14887 ( .A(n12546), .B(n12568), .ZN(n15118) );
  NOR2_X1 U14888 ( .A1(n12568), .A2(n12546), .ZN(n12547) );
  NOR2_X1 U14889 ( .A1(n15117), .A2(n12547), .ZN(n15139) );
  MUX2_X1 U14890 ( .A(n12548), .B(P3_REG2_REG_10__SCAN_IN), .S(n12571), .Z(
        n15140) );
  NAND2_X1 U14891 ( .A1(n12571), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n12549) );
  NOR2_X1 U14892 ( .A1(n12574), .A2(n12550), .ZN(n12551) );
  NOR2_X1 U14893 ( .A1(n9435), .A2(n15158), .ZN(n15157) );
  NAND2_X1 U14894 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n15181), .ZN(n12552) );
  OAI21_X1 U14895 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n15181), .A(n12552), 
        .ZN(n15174) );
  NOR2_X1 U14896 ( .A1(n15175), .A2(n15174), .ZN(n15173) );
  INV_X1 U14897 ( .A(n15199), .ZN(n12580) );
  XNOR2_X1 U14898 ( .A(n12553), .B(n12580), .ZN(n15193) );
  XNOR2_X1 U14899 ( .A(n15217), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n15210) );
  NOR2_X1 U14900 ( .A1(n12554), .A2(n12555), .ZN(n12556) );
  AOI22_X1 U14901 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n14372), .B1(n12590), 
        .B2(n12557), .ZN(n14367) );
  NOR2_X1 U14902 ( .A1(n12594), .A2(n12558), .ZN(n12559) );
  INV_X1 U14903 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12560) );
  AOI22_X1 U14904 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n14404), .B1(n12597), 
        .B2(n12560), .ZN(n14413) );
  INV_X1 U14905 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12561) );
  MUX2_X1 U14906 ( .A(P3_REG2_REG_19__SCAN_IN), .B(n12561), .S(n12608), .Z(
        n12601) );
  NAND2_X1 U14907 ( .A1(n12562), .A2(n15151), .ZN(n12609) );
  MUX2_X1 U14908 ( .A(n12560), .B(n12563), .S(n12589), .Z(n14409) );
  INV_X1 U14909 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12882) );
  MUX2_X1 U14910 ( .A(n14389), .B(n12882), .S(n12589), .Z(n12593) );
  NOR2_X1 U14911 ( .A1(n12593), .A2(n12594), .ZN(n12596) );
  MUX2_X1 U14912 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12589), .Z(n12573) );
  XNOR2_X1 U14913 ( .A(n12573), .B(n12574), .ZN(n15167) );
  MUX2_X1 U14914 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12589), .Z(n12572) );
  MUX2_X1 U14915 ( .A(n9381), .B(n9377), .S(n12589), .Z(n12569) );
  OR2_X1 U14916 ( .A1(n12569), .A2(n12568), .ZN(n15120) );
  OR2_X1 U14917 ( .A1(n12565), .A2(n12564), .ZN(n12567) );
  NAND2_X1 U14918 ( .A1(n12567), .A2(n12566), .ZN(n15123) );
  AND2_X1 U14919 ( .A1(n12569), .A2(n12568), .ZN(n15119) );
  XNOR2_X1 U14920 ( .A(n12572), .B(n12571), .ZN(n15145) );
  NOR2_X1 U14921 ( .A1(n15146), .A2(n15145), .ZN(n15144) );
  INV_X1 U14922 ( .A(n15144), .ZN(n12570) );
  INV_X1 U14923 ( .A(n12573), .ZN(n12575) );
  NAND2_X1 U14924 ( .A1(n12575), .A2(n12574), .ZN(n12576) );
  MUX2_X1 U14925 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12589), .Z(n12577) );
  XNOR2_X1 U14926 ( .A(n12577), .B(n15181), .ZN(n15186) );
  NAND2_X1 U14927 ( .A1(n12577), .A2(n15181), .ZN(n12578) );
  MUX2_X1 U14928 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12589), .Z(n12579) );
  XNOR2_X1 U14929 ( .A(n12579), .B(n12580), .ZN(n15203) );
  INV_X1 U14930 ( .A(n12579), .ZN(n12581) );
  NAND2_X1 U14931 ( .A1(n12581), .A2(n12580), .ZN(n12582) );
  INV_X1 U14932 ( .A(n15210), .ZN(n12583) );
  MUX2_X1 U14933 ( .A(n12583), .B(n15213), .S(n12589), .Z(n15224) );
  NAND2_X1 U14934 ( .A1(n15225), .A2(n15224), .ZN(n15223) );
  MUX2_X1 U14935 ( .A(n12585), .B(n12584), .S(n12589), .Z(n12586) );
  INV_X1 U14936 ( .A(n12587), .ZN(n12588) );
  XNOR2_X1 U14937 ( .A(n12587), .B(n14328), .ZN(n14361) );
  MUX2_X1 U14938 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12589), .Z(n14362) );
  NOR2_X1 U14939 ( .A1(n14361), .A2(n14362), .ZN(n14360) );
  MUX2_X1 U14940 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12589), .Z(n12591) );
  AND2_X1 U14941 ( .A1(n12591), .A2(n12590), .ZN(n14379) );
  INV_X1 U14942 ( .A(n12591), .ZN(n12592) );
  NAND2_X1 U14943 ( .A1(n12592), .A2(n14372), .ZN(n14378) );
  OAI21_X1 U14944 ( .B1(n14383), .B2(n14379), .A(n14378), .ZN(n14394) );
  AOI21_X1 U14945 ( .B1(n12594), .B2(n12593), .A(n12596), .ZN(n12595) );
  INV_X1 U14946 ( .A(n12595), .ZN(n14395) );
  NOR2_X1 U14947 ( .A1(n12596), .A2(n14393), .ZN(n12598) );
  NAND2_X1 U14948 ( .A1(n14409), .A2(n14410), .ZN(n14408) );
  NAND2_X1 U14949 ( .A1(n14404), .A2(n12598), .ZN(n12599) );
  NAND2_X1 U14950 ( .A1(n14408), .A2(n12599), .ZN(n12603) );
  MUX2_X1 U14951 ( .A(n6728), .B(n12601), .S(n12600), .Z(n12602) );
  XNOR2_X1 U14952 ( .A(n12603), .B(n12602), .ZN(n12604) );
  OAI21_X1 U14953 ( .B1(n15156), .B2(n12606), .A(n12605), .ZN(n12607) );
  OAI211_X1 U14954 ( .C1(n12610), .C2(n15108), .A(n12609), .B(n6698), .ZN(
        P3_U3201) );
  NAND2_X1 U14955 ( .A1(n12618), .A2(n15253), .ZN(n12613) );
  OR2_X1 U14956 ( .A1(n12612), .A2(n12611), .ZN(n12898) );
  AOI21_X1 U14957 ( .B1(n12613), .B2(n12898), .A(n15333), .ZN(n12615) );
  AOI21_X1 U14958 ( .B1(n15333), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12615), 
        .ZN(n12614) );
  OAI21_X1 U14959 ( .B1(n7195), .B2(n12812), .A(n12614), .ZN(P3_U3202) );
  AOI21_X1 U14960 ( .B1(n15333), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12615), 
        .ZN(n12616) );
  OAI21_X1 U14961 ( .B1(n12835), .B2(n12812), .A(n12616), .ZN(P3_U3203) );
  INV_X1 U14962 ( .A(n12617), .ZN(n12624) );
  AOI22_X1 U14963 ( .A1(n12618), .A2(n15253), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n15333), .ZN(n12619) );
  OAI21_X1 U14964 ( .B1(n12620), .B2(n12812), .A(n12619), .ZN(n12621) );
  AOI21_X1 U14965 ( .B1(n12622), .B2(n15265), .A(n12621), .ZN(n12623) );
  OAI21_X1 U14966 ( .B1(n12624), .B2(n15333), .A(n12623), .ZN(P3_U3204) );
  INV_X1 U14967 ( .A(n12625), .ZN(n12632) );
  AOI22_X1 U14968 ( .A1(n12626), .A2(n15253), .B1(n15333), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12627) );
  OAI21_X1 U14969 ( .B1(n12628), .B2(n12812), .A(n12627), .ZN(n12629) );
  AOI21_X1 U14970 ( .B1(n12630), .B2(n15265), .A(n12629), .ZN(n12631) );
  OAI21_X1 U14971 ( .B1(n12632), .B2(n15333), .A(n12631), .ZN(P3_U3205) );
  NAND2_X1 U14972 ( .A1(n12633), .A2(n12640), .ZN(n12634) );
  NAND2_X1 U14973 ( .A1(n12635), .A2(n12634), .ZN(n12639) );
  OAI22_X1 U14974 ( .A1(n12637), .A2(n15294), .B1(n12636), .B2(n15292), .ZN(
        n12638) );
  AOI21_X1 U14975 ( .B1(n12639), .B2(n15319), .A(n12638), .ZN(n12839) );
  OR2_X1 U14976 ( .A1(n12641), .A2(n12640), .ZN(n12642) );
  NAND2_X1 U14977 ( .A1(n12643), .A2(n12642), .ZN(n12837) );
  INV_X1 U14978 ( .A(n12836), .ZN(n12646) );
  AOI22_X1 U14979 ( .A1(n12644), .A2(n15253), .B1(n15333), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12645) );
  OAI21_X1 U14980 ( .B1(n12646), .B2(n12812), .A(n12645), .ZN(n12647) );
  AOI21_X1 U14981 ( .B1(n12837), .B2(n15265), .A(n12647), .ZN(n12648) );
  OAI21_X1 U14982 ( .B1(n12839), .B2(n15333), .A(n12648), .ZN(P3_U3206) );
  XNOR2_X1 U14983 ( .A(n12650), .B(n12649), .ZN(n12842) );
  INV_X1 U14984 ( .A(n12842), .ZN(n12664) );
  XNOR2_X1 U14985 ( .A(n12651), .B(n12652), .ZN(n12657) );
  OAI22_X1 U14986 ( .A1(n12654), .A2(n15294), .B1(n12653), .B2(n15292), .ZN(
        n12655) );
  AOI21_X1 U14987 ( .B1(n12842), .B2(n15297), .A(n12655), .ZN(n12656) );
  OAI21_X1 U14988 ( .B1(n12657), .B2(n15299), .A(n12656), .ZN(n12841) );
  NAND2_X1 U14989 ( .A1(n12841), .A2(n15330), .ZN(n12663) );
  NAND2_X1 U14990 ( .A1(n12658), .A2(n15253), .ZN(n12659) );
  OAI21_X1 U14991 ( .B1(n15330), .B2(n12660), .A(n12659), .ZN(n12661) );
  AOI21_X1 U14992 ( .B1(n12840), .B2(n12695), .A(n12661), .ZN(n12662) );
  OAI211_X1 U14993 ( .C1(n12664), .C2(n12698), .A(n12663), .B(n12662), .ZN(
        P3_U3207) );
  NAND2_X1 U14994 ( .A1(n12665), .A2(n12686), .ZN(n12685) );
  NAND2_X1 U14995 ( .A1(n12685), .A2(n12666), .ZN(n12668) );
  OAI211_X1 U14996 ( .C1(n12669), .C2(n12668), .A(n12667), .B(n15319), .ZN(
        n12672) );
  AOI22_X1 U14997 ( .A1(n15323), .A2(n12702), .B1(n12670), .B2(n15322), .ZN(
        n12671) );
  XNOR2_X1 U14998 ( .A(n12674), .B(n12673), .ZN(n12846) );
  INV_X1 U14999 ( .A(n12845), .ZN(n12677) );
  AOI22_X1 U15000 ( .A1(n12675), .A2(n15253), .B1(n15333), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12676) );
  OAI21_X1 U15001 ( .B1(n12677), .B2(n12812), .A(n12676), .ZN(n12678) );
  AOI21_X1 U15002 ( .B1(n12846), .B2(n15265), .A(n12678), .ZN(n12679) );
  OAI21_X1 U15003 ( .B1(n12848), .B2(n15333), .A(n12679), .ZN(P3_U3208) );
  INV_X1 U15004 ( .A(n12680), .ZN(n12684) );
  AOI21_X1 U15005 ( .B1(n12709), .B2(n12682), .A(n12681), .ZN(n12683) );
  OAI211_X1 U15006 ( .C1(n12665), .C2(n12686), .A(n12685), .B(n15319), .ZN(
        n12690) );
  AOI22_X1 U15007 ( .A1(n12688), .A2(n15322), .B1(n15323), .B2(n12687), .ZN(
        n12689) );
  OAI211_X1 U15008 ( .C1(n15327), .C2(n12850), .A(n12690), .B(n12689), .ZN(
        n12851) );
  NAND2_X1 U15009 ( .A1(n12851), .A2(n15330), .ZN(n12697) );
  INV_X1 U15010 ( .A(n12691), .ZN(n12693) );
  OAI22_X1 U15011 ( .A1(n12693), .A2(n15312), .B1(n15330), .B2(n12692), .ZN(
        n12694) );
  AOI21_X1 U15012 ( .B1(n12849), .B2(n12695), .A(n12694), .ZN(n12696) );
  OAI211_X1 U15013 ( .C1(n12850), .C2(n12698), .A(n12697), .B(n12696), .ZN(
        P3_U3209) );
  OAI211_X1 U15014 ( .C1(n12700), .C2(n7170), .A(n12699), .B(n15319), .ZN(
        n12704) );
  AOI22_X1 U15015 ( .A1(n12702), .A2(n15322), .B1(n15323), .B2(n12701), .ZN(
        n12703) );
  NAND2_X1 U15016 ( .A1(n12704), .A2(n12703), .ZN(n12855) );
  INV_X1 U15017 ( .A(n12705), .ZN(n12918) );
  OR2_X1 U15018 ( .A1(n12707), .A2(n12706), .ZN(n12708) );
  AND2_X1 U15019 ( .A1(n12709), .A2(n12708), .ZN(n12856) );
  NAND2_X1 U15020 ( .A1(n12856), .A2(n15265), .ZN(n12712) );
  AOI22_X1 U15021 ( .A1(n12710), .A2(n15253), .B1(n15333), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n12711) );
  OAI211_X1 U15022 ( .C1(n12918), .C2(n12812), .A(n12712), .B(n12711), .ZN(
        n12713) );
  AOI21_X1 U15023 ( .B1(n12855), .B2(n15330), .A(n12713), .ZN(n12714) );
  INV_X1 U15024 ( .A(n12714), .ZN(P3_U3210) );
  XNOR2_X1 U15025 ( .A(n12715), .B(n12718), .ZN(n12716) );
  OAI222_X1 U15026 ( .A1(n15294), .A2(n12717), .B1(n15292), .B2(n12742), .C1(
        n15299), .C2(n12716), .ZN(n12859) );
  INV_X1 U15027 ( .A(n12859), .ZN(n12725) );
  XOR2_X1 U15028 ( .A(n12719), .B(n12718), .Z(n12860) );
  INV_X1 U15029 ( .A(n12720), .ZN(n12922) );
  AOI22_X1 U15030 ( .A1(n15333), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n12721), 
        .B2(n15253), .ZN(n12722) );
  OAI21_X1 U15031 ( .B1(n12922), .B2(n12812), .A(n12722), .ZN(n12723) );
  AOI21_X1 U15032 ( .B1(n12860), .B2(n15265), .A(n12723), .ZN(n12724) );
  OAI21_X1 U15033 ( .B1(n12725), .B2(n15333), .A(n12724), .ZN(P3_U3211) );
  INV_X1 U15034 ( .A(n12726), .ZN(n12727) );
  AOI21_X1 U15035 ( .B1(n12732), .B2(n12728), .A(n12727), .ZN(n12729) );
  OAI222_X1 U15036 ( .A1(n15294), .A2(n12731), .B1(n15292), .B2(n12730), .C1(
        n15299), .C2(n12729), .ZN(n12863) );
  INV_X1 U15037 ( .A(n12863), .ZN(n12738) );
  XOR2_X1 U15038 ( .A(n12733), .B(n12732), .Z(n12864) );
  AOI22_X1 U15039 ( .A1(n15333), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15253), 
        .B2(n12734), .ZN(n12735) );
  OAI21_X1 U15040 ( .B1(n12926), .B2(n12812), .A(n12735), .ZN(n12736) );
  AOI21_X1 U15041 ( .B1(n12864), .B2(n15265), .A(n12736), .ZN(n12737) );
  OAI21_X1 U15042 ( .B1(n12738), .B2(n15333), .A(n12737), .ZN(P3_U3212) );
  XNOR2_X1 U15043 ( .A(n12739), .B(n12744), .ZN(n12740) );
  OAI222_X1 U15044 ( .A1(n15294), .A2(n12742), .B1(n15292), .B2(n12741), .C1(
        n12740), .C2(n15299), .ZN(n12867) );
  INV_X1 U15045 ( .A(n12867), .ZN(n12749) );
  AOI21_X1 U15046 ( .B1(n12744), .B2(n12743), .A(n6640), .ZN(n12868) );
  AOI22_X1 U15047 ( .A1(n15333), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15253), 
        .B2(n12745), .ZN(n12746) );
  OAI21_X1 U15048 ( .B1(n12930), .B2(n12812), .A(n12746), .ZN(n12747) );
  AOI21_X1 U15049 ( .B1(n12868), .B2(n15265), .A(n12747), .ZN(n12748) );
  OAI21_X1 U15050 ( .B1(n12749), .B2(n15333), .A(n12748), .ZN(P3_U3213) );
  OAI211_X1 U15051 ( .C1(n6716), .C2(n7537), .A(n15319), .B(n12750), .ZN(
        n12754) );
  AOI22_X1 U15052 ( .A1(n12752), .A2(n15322), .B1(n15323), .B2(n12751), .ZN(
        n12753) );
  NAND2_X1 U15053 ( .A1(n12754), .A2(n12753), .ZN(n12871) );
  INV_X1 U15054 ( .A(n12871), .ZN(n12760) );
  XNOR2_X1 U15055 ( .A(n12755), .B(n7537), .ZN(n12872) );
  AOI22_X1 U15056 ( .A1(n15333), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15253), 
        .B2(n12756), .ZN(n12757) );
  OAI21_X1 U15057 ( .B1(n12934), .B2(n12812), .A(n12757), .ZN(n12758) );
  AOI21_X1 U15058 ( .B1(n12872), .B2(n15265), .A(n12758), .ZN(n12759) );
  OAI21_X1 U15059 ( .B1(n12760), .B2(n15333), .A(n12759), .ZN(P3_U3214) );
  OAI21_X1 U15060 ( .B1(n12762), .B2(n9562), .A(n12761), .ZN(n12764) );
  AOI222_X1 U15061 ( .A1(n15319), .A2(n12764), .B1(n12792), .B2(n15323), .C1(
        n12763), .C2(n15322), .ZN(n12879) );
  NAND2_X1 U15062 ( .A1(n12765), .A2(n15301), .ZN(n12877) );
  INV_X1 U15063 ( .A(n12877), .ZN(n12769) );
  INV_X1 U15064 ( .A(n12766), .ZN(n12767) );
  OAI22_X1 U15065 ( .A1(n15330), .A2(n12560), .B1(n12767), .B2(n15312), .ZN(
        n12768) );
  AOI21_X1 U15066 ( .B1(n12769), .B2(n15305), .A(n12768), .ZN(n12777) );
  AND2_X1 U15067 ( .A1(n12771), .A2(n12770), .ZN(n12876) );
  NAND2_X1 U15068 ( .A1(n12796), .A2(n12772), .ZN(n12774) );
  AND2_X1 U15069 ( .A1(n12774), .A2(n12773), .ZN(n12775) );
  NAND2_X1 U15070 ( .A1(n12775), .A2(n9562), .ZN(n12875) );
  NAND3_X1 U15071 ( .A1(n12876), .A2(n12875), .A3(n15265), .ZN(n12776) );
  OAI211_X1 U15072 ( .C1(n12879), .C2(n15333), .A(n12777), .B(n12776), .ZN(
        P3_U3215) );
  XNOR2_X1 U15073 ( .A(n12778), .B(n12779), .ZN(n12780) );
  OAI222_X1 U15074 ( .A1(n15294), .A2(n12781), .B1(n15292), .B2(n12807), .C1(
        n12780), .C2(n15299), .ZN(n12880) );
  INV_X1 U15075 ( .A(n12880), .ZN(n12789) );
  NAND2_X1 U15076 ( .A1(n12796), .A2(n12782), .ZN(n12784) );
  XNOR2_X1 U15077 ( .A(n12784), .B(n12783), .ZN(n12881) );
  AOI22_X1 U15078 ( .A1(n15333), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15253), 
        .B2(n12785), .ZN(n12786) );
  OAI21_X1 U15079 ( .B1(n12939), .B2(n12812), .A(n12786), .ZN(n12787) );
  AOI21_X1 U15080 ( .B1(n12881), .B2(n15265), .A(n12787), .ZN(n12788) );
  OAI21_X1 U15081 ( .B1(n12789), .B2(n15333), .A(n12788), .ZN(P3_U3216) );
  XNOR2_X1 U15082 ( .A(n12790), .B(n12798), .ZN(n12793) );
  AOI222_X1 U15083 ( .A1(n15319), .A2(n12793), .B1(n12792), .B2(n15322), .C1(
        n12791), .C2(n15323), .ZN(n12887) );
  NAND2_X1 U15084 ( .A1(n12809), .A2(n12808), .ZN(n12795) );
  NAND2_X1 U15085 ( .A1(n12795), .A2(n12794), .ZN(n12797) );
  OAI21_X1 U15086 ( .B1(n12798), .B2(n12797), .A(n12796), .ZN(n12885) );
  AOI22_X1 U15087 ( .A1(n15333), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15253), 
        .B2(n12799), .ZN(n12800) );
  OAI21_X1 U15088 ( .B1(n12801), .B2(n12812), .A(n12800), .ZN(n12802) );
  AOI21_X1 U15089 ( .B1(n12885), .B2(n15265), .A(n12802), .ZN(n12803) );
  OAI21_X1 U15090 ( .B1(n12887), .B2(n15333), .A(n12803), .ZN(P3_U3217) );
  XOR2_X1 U15091 ( .A(n12808), .B(n12804), .Z(n12805) );
  OAI222_X1 U15092 ( .A1(n15294), .A2(n12807), .B1(n15292), .B2(n12806), .C1(
        n12805), .C2(n15299), .ZN(n12888) );
  INV_X1 U15093 ( .A(n12888), .ZN(n12815) );
  XNOR2_X1 U15094 ( .A(n12809), .B(n12808), .ZN(n12889) );
  AOI22_X1 U15095 ( .A1(n15333), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15253), 
        .B2(n12810), .ZN(n12811) );
  OAI21_X1 U15096 ( .B1(n12944), .B2(n12812), .A(n12811), .ZN(n12813) );
  AOI21_X1 U15097 ( .B1(n12889), .B2(n15265), .A(n12813), .ZN(n12814) );
  OAI21_X1 U15098 ( .B1(n12815), .B2(n15333), .A(n12814), .ZN(P3_U3218) );
  OAI21_X1 U15099 ( .B1(n12816), .B2(n12823), .A(n15318), .ZN(n12821) );
  NAND2_X1 U15100 ( .A1(n12817), .A2(n15323), .ZN(n12818) );
  OAI21_X1 U15101 ( .B1(n12819), .B2(n15294), .A(n12818), .ZN(n12820) );
  AOI21_X1 U15102 ( .B1(n12821), .B2(n15319), .A(n12820), .ZN(n12825) );
  XNOR2_X1 U15103 ( .A(n12823), .B(n12822), .ZN(n12826) );
  OR2_X1 U15104 ( .A1(n12826), .A2(n15327), .ZN(n12824) );
  AND2_X1 U15105 ( .A1(n12825), .A2(n12824), .ZN(n15335) );
  INV_X1 U15106 ( .A(n12826), .ZN(n15338) );
  NAND2_X1 U15107 ( .A1(n12827), .A2(n15301), .ZN(n15334) );
  OAI22_X1 U15108 ( .A1(n15312), .A2(n12828), .B1(n15313), .B2(n15334), .ZN(
        n12829) );
  AOI21_X1 U15109 ( .B1(n15338), .B2(n15329), .A(n12829), .ZN(n12830) );
  NAND2_X1 U15110 ( .A1(n15335), .A2(n12830), .ZN(n12831) );
  MUX2_X1 U15111 ( .A(n12831), .B(P3_REG2_REG_1__SCAN_IN), .S(n15333), .Z(
        P3_U3232) );
  NOR2_X1 U15112 ( .A1(n12898), .A2(n15392), .ZN(n12833) );
  AOI21_X1 U15113 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n15392), .A(n12833), 
        .ZN(n12832) );
  OAI21_X1 U15114 ( .B1(n7195), .B2(n12896), .A(n12832), .ZN(P3_U3490) );
  AOI21_X1 U15115 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(n15392), .A(n12833), 
        .ZN(n12834) );
  OAI21_X1 U15116 ( .B1(n12835), .B2(n12896), .A(n12834), .ZN(P3_U3489) );
  AOI22_X1 U15117 ( .A1(n12837), .A2(n15366), .B1(n15301), .B2(n12836), .ZN(
        n12838) );
  NAND2_X1 U15118 ( .A1(n12839), .A2(n12838), .ZN(n12905) );
  MUX2_X1 U15119 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n12905), .S(n15395), .Z(
        P3_U3486) );
  INV_X1 U15120 ( .A(n12840), .ZN(n12909) );
  INV_X1 U15121 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12843) );
  AOI21_X1 U15122 ( .B1(n15377), .B2(n12842), .A(n12841), .ZN(n12906) );
  MUX2_X1 U15123 ( .A(n12843), .B(n12906), .S(n15395), .Z(n12844) );
  OAI21_X1 U15124 ( .B1(n12909), .B2(n12896), .A(n12844), .ZN(P3_U3485) );
  AOI22_X1 U15125 ( .A1(n12846), .A2(n15366), .B1(n15301), .B2(n12845), .ZN(
        n12847) );
  NAND2_X1 U15126 ( .A1(n12848), .A2(n12847), .ZN(n12910) );
  MUX2_X1 U15127 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n12910), .S(n15395), .Z(
        P3_U3484) );
  INV_X1 U15128 ( .A(n12849), .ZN(n12914) );
  INV_X1 U15129 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12853) );
  INV_X1 U15130 ( .A(n12850), .ZN(n12852) );
  AOI21_X1 U15131 ( .B1(n15377), .B2(n12852), .A(n12851), .ZN(n12911) );
  MUX2_X1 U15132 ( .A(n12853), .B(n12911), .S(n15395), .Z(n12854) );
  OAI21_X1 U15133 ( .B1(n12914), .B2(n12896), .A(n12854), .ZN(P3_U3483) );
  INV_X1 U15134 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12857) );
  AOI21_X1 U15135 ( .B1(n12856), .B2(n15366), .A(n12855), .ZN(n12915) );
  MUX2_X1 U15136 ( .A(n12857), .B(n12915), .S(n15395), .Z(n12858) );
  OAI21_X1 U15137 ( .B1(n12918), .B2(n12896), .A(n12858), .ZN(P3_U3482) );
  INV_X1 U15138 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12861) );
  AOI21_X1 U15139 ( .B1(n15366), .B2(n12860), .A(n12859), .ZN(n12919) );
  MUX2_X1 U15140 ( .A(n12861), .B(n12919), .S(n15395), .Z(n12862) );
  OAI21_X1 U15141 ( .B1(n12922), .B2(n12896), .A(n12862), .ZN(P3_U3481) );
  INV_X1 U15142 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12865) );
  AOI21_X1 U15143 ( .B1(n15366), .B2(n12864), .A(n12863), .ZN(n12923) );
  MUX2_X1 U15144 ( .A(n12865), .B(n12923), .S(n15395), .Z(n12866) );
  OAI21_X1 U15145 ( .B1(n12926), .B2(n12896), .A(n12866), .ZN(P3_U3480) );
  INV_X1 U15146 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12869) );
  AOI21_X1 U15147 ( .B1(n12868), .B2(n15366), .A(n12867), .ZN(n12927) );
  MUX2_X1 U15148 ( .A(n12869), .B(n12927), .S(n15395), .Z(n12870) );
  OAI21_X1 U15149 ( .B1(n12930), .B2(n12896), .A(n12870), .ZN(P3_U3479) );
  INV_X1 U15150 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12873) );
  AOI21_X1 U15151 ( .B1(n15366), .B2(n12872), .A(n12871), .ZN(n12931) );
  MUX2_X1 U15152 ( .A(n12873), .B(n12931), .S(n15395), .Z(n12874) );
  OAI21_X1 U15153 ( .B1(n12934), .B2(n12896), .A(n12874), .ZN(P3_U3478) );
  NAND3_X1 U15154 ( .A1(n12876), .A2(n12875), .A3(n15366), .ZN(n12878) );
  NAND3_X1 U15155 ( .A1(n12879), .A2(n12878), .A3(n12877), .ZN(n12935) );
  MUX2_X1 U15156 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12935), .S(n15395), .Z(
        P3_U3477) );
  AOI21_X1 U15157 ( .B1(n12881), .B2(n15366), .A(n12880), .ZN(n12936) );
  MUX2_X1 U15158 ( .A(n12882), .B(n12936), .S(n15395), .Z(n12883) );
  OAI21_X1 U15159 ( .B1(n12896), .B2(n12939), .A(n12883), .ZN(P3_U3476) );
  AOI22_X1 U15160 ( .A1(n12885), .A2(n15366), .B1(n15301), .B2(n12884), .ZN(
        n12886) );
  NAND2_X1 U15161 ( .A1(n12887), .A2(n12886), .ZN(n12940) );
  MUX2_X1 U15162 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n12940), .S(n15395), .Z(
        P3_U3475) );
  AOI21_X1 U15163 ( .B1(n12889), .B2(n15366), .A(n12888), .ZN(n12941) );
  MUX2_X1 U15164 ( .A(n12890), .B(n12941), .S(n15395), .Z(n12891) );
  OAI21_X1 U15165 ( .B1(n12896), .B2(n12944), .A(n12891), .ZN(P3_U3474) );
  AOI21_X1 U15166 ( .B1(n15366), .B2(n12893), .A(n12892), .ZN(n12945) );
  MUX2_X1 U15167 ( .A(n12894), .B(n12945), .S(n15395), .Z(n12895) );
  OAI21_X1 U15168 ( .B1(n12896), .B2(n12948), .A(n12895), .ZN(P3_U3473) );
  NAND2_X1 U15169 ( .A1(n12897), .A2(n9832), .ZN(n12900) );
  INV_X1 U15170 ( .A(n12898), .ZN(n12899) );
  NAND2_X1 U15171 ( .A1(n12899), .A2(n15379), .ZN(n12902) );
  OAI211_X1 U15172 ( .C1(n12303), .C2(n15379), .A(n12900), .B(n12902), .ZN(
        P3_U3458) );
  INV_X1 U15173 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n12904) );
  NAND2_X1 U15174 ( .A1(n12901), .A2(n9832), .ZN(n12903) );
  OAI211_X1 U15175 ( .C1(n12904), .C2(n15379), .A(n12903), .B(n12902), .ZN(
        P3_U3457) );
  MUX2_X1 U15176 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n12905), .S(n15379), .Z(
        P3_U3454) );
  INV_X1 U15177 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12907) );
  MUX2_X1 U15178 ( .A(n12907), .B(n12906), .S(n15379), .Z(n12908) );
  OAI21_X1 U15179 ( .B1(n12909), .B2(n12949), .A(n12908), .ZN(P3_U3453) );
  MUX2_X1 U15180 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n12910), .S(n15379), .Z(
        P3_U3452) );
  INV_X1 U15181 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12912) );
  MUX2_X1 U15182 ( .A(n12912), .B(n12911), .S(n15379), .Z(n12913) );
  OAI21_X1 U15183 ( .B1(n12914), .B2(n12949), .A(n12913), .ZN(P3_U3451) );
  INV_X1 U15184 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12916) );
  MUX2_X1 U15185 ( .A(n12916), .B(n12915), .S(n15379), .Z(n12917) );
  OAI21_X1 U15186 ( .B1(n12918), .B2(n12949), .A(n12917), .ZN(P3_U3450) );
  INV_X1 U15187 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12920) );
  MUX2_X1 U15188 ( .A(n12920), .B(n12919), .S(n15379), .Z(n12921) );
  OAI21_X1 U15189 ( .B1(n12922), .B2(n12949), .A(n12921), .ZN(P3_U3449) );
  INV_X1 U15190 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12924) );
  MUX2_X1 U15191 ( .A(n12924), .B(n12923), .S(n15379), .Z(n12925) );
  OAI21_X1 U15192 ( .B1(n12926), .B2(n12949), .A(n12925), .ZN(P3_U3448) );
  INV_X1 U15193 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12928) );
  MUX2_X1 U15194 ( .A(n12928), .B(n12927), .S(n15379), .Z(n12929) );
  OAI21_X1 U15195 ( .B1(n12930), .B2(n12949), .A(n12929), .ZN(P3_U3447) );
  INV_X1 U15196 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12932) );
  MUX2_X1 U15197 ( .A(n12932), .B(n12931), .S(n15379), .Z(n12933) );
  OAI21_X1 U15198 ( .B1(n12934), .B2(n12949), .A(n12933), .ZN(P3_U3446) );
  MUX2_X1 U15199 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n12935), .S(n15379), .Z(
        P3_U3444) );
  MUX2_X1 U15200 ( .A(n12937), .B(n12936), .S(n15379), .Z(n12938) );
  OAI21_X1 U15201 ( .B1(n12949), .B2(n12939), .A(n12938), .ZN(P3_U3441) );
  MUX2_X1 U15202 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n12940), .S(n15379), .Z(
        P3_U3438) );
  INV_X1 U15203 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12942) );
  MUX2_X1 U15204 ( .A(n12942), .B(n12941), .S(n15379), .Z(n12943) );
  OAI21_X1 U15205 ( .B1(n12949), .B2(n12944), .A(n12943), .ZN(P3_U3435) );
  MUX2_X1 U15206 ( .A(n12946), .B(n12945), .S(n15379), .Z(n12947) );
  OAI21_X1 U15207 ( .B1(n12949), .B2(n12948), .A(n12947), .ZN(P3_U3432) );
  MUX2_X1 U15208 ( .A(n12950), .B(P3_D_REG_1__SCAN_IN), .S(n12951), .Z(
        P3_U3377) );
  MUX2_X1 U15209 ( .A(n12952), .B(P3_D_REG_0__SCAN_IN), .S(n12951), .Z(
        P3_U3376) );
  INV_X1 U15210 ( .A(n12953), .ZN(n12956) );
  NOR4_X1 U15211 ( .A1(n7205), .A2(P3_IR_REG_30__SCAN_IN), .A3(n9231), .A4(
        P3_U3151), .ZN(n12954) );
  AOI21_X1 U15212 ( .B1(n6727), .B2(SI_31_), .A(n12954), .ZN(n12955) );
  OAI21_X1 U15213 ( .B1(n12956), .B2(n12961), .A(n12955), .ZN(P3_U3264) );
  INV_X1 U15214 ( .A(n12957), .ZN(n12960) );
  OAI222_X1 U15215 ( .A1(n12962), .A2(n13652), .B1(n12961), .B2(n12960), .C1(
        n12959), .C2(P3_U3151), .ZN(P3_U3266) );
  MUX2_X1 U15216 ( .A(n12963), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  AOI21_X1 U15217 ( .B1(n12965), .B2(n12964), .A(n13059), .ZN(n12967) );
  NAND2_X1 U15218 ( .A1(n12967), .A2(n12966), .ZN(n12975) );
  INV_X1 U15219 ( .A(n12968), .ZN(n13200) );
  OR2_X1 U15220 ( .A1(n12969), .A2(n14443), .ZN(n12971) );
  NAND2_X1 U15221 ( .A1(n13065), .A2(n13335), .ZN(n12970) );
  AND2_X1 U15222 ( .A1(n12971), .A2(n12970), .ZN(n13195) );
  OAI22_X1 U15223 ( .A1(n13012), .A2(n13195), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12972), .ZN(n12973) );
  AOI21_X1 U15224 ( .B1(n13200), .B2(n13014), .A(n12973), .ZN(n12974) );
  OAI211_X1 U15225 ( .C1(n13202), .C2(n13017), .A(n12975), .B(n12974), .ZN(
        P2_U3186) );
  OAI211_X1 U15226 ( .C1(n12978), .C2(n12977), .A(n12976), .B(n14448), .ZN(
        n12982) );
  NOR2_X1 U15227 ( .A1(n14453), .A2(n13265), .ZN(n12980) );
  OAI22_X1 U15228 ( .A1(n13263), .A2(n13045), .B1(n13044), .B2(n13262), .ZN(
        n12979) );
  AOI211_X1 U15229 ( .C1(P2_REG3_REG_23__SCAN_IN), .C2(P2_U3088), .A(n12980), 
        .B(n12979), .ZN(n12981) );
  OAI211_X1 U15230 ( .C1(n7088), .C2(n13017), .A(n12982), .B(n12981), .ZN(
        P2_U3188) );
  OAI21_X1 U15231 ( .B1(n12985), .B2(n12984), .A(n12983), .ZN(n12986) );
  NAND2_X1 U15232 ( .A1(n12986), .A2(n14448), .ZN(n12991) );
  INV_X1 U15233 ( .A(n12987), .ZN(n13323) );
  AOI22_X1 U15234 ( .A1(n13069), .A2(n13336), .B1(n13335), .B2(n13070), .ZN(
        n13319) );
  OAI22_X1 U15235 ( .A1(n13012), .A2(n13319), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12988), .ZN(n12989) );
  AOI21_X1 U15236 ( .B1(n13323), .B2(n13014), .A(n12989), .ZN(n12990) );
  OAI211_X1 U15237 ( .C1(n8200), .C2(n13017), .A(n12991), .B(n12990), .ZN(
        P2_U3191) );
  OAI211_X1 U15238 ( .C1(n12994), .C2(n12993), .A(n12992), .B(n14448), .ZN(
        n12998) );
  AOI22_X1 U15239 ( .A1(n13069), .A2(n13335), .B1(n13336), .B2(n13068), .ZN(
        n13288) );
  INV_X1 U15240 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12995) );
  OAI22_X1 U15241 ( .A1(n13012), .A2(n13288), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12995), .ZN(n12996) );
  AOI21_X1 U15242 ( .B1(n13296), .B2(n13014), .A(n12996), .ZN(n12997) );
  OAI211_X1 U15243 ( .C1(n13469), .C2(n13017), .A(n12998), .B(n12997), .ZN(
        P2_U3195) );
  OAI21_X1 U15244 ( .B1(n12999), .B2(n13000), .A(n14448), .ZN(n13006) );
  OAI22_X1 U15245 ( .A1(n13262), .A2(n14441), .B1(n13001), .B2(n14443), .ZN(
        n13227) );
  AOI22_X1 U15246 ( .A1(n14450), .A2(n13227), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13002) );
  OAI21_X1 U15247 ( .B1(n13232), .B2(n14453), .A(n13002), .ZN(n13003) );
  AOI21_X1 U15248 ( .B1(n13392), .B2(n14451), .A(n13003), .ZN(n13004) );
  OAI21_X1 U15249 ( .B1(n13006), .B2(n13005), .A(n13004), .ZN(P2_U3197) );
  OAI211_X1 U15250 ( .C1(n13007), .C2(n13009), .A(n13008), .B(n14448), .ZN(
        n13016) );
  INV_X1 U15251 ( .A(n13010), .ZN(n13248) );
  AOI22_X1 U15252 ( .A1(n13335), .A2(n13271), .B1(n13066), .B2(n13336), .ZN(
        n13241) );
  INV_X1 U15253 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13011) );
  OAI22_X1 U15254 ( .A1(n13012), .A2(n13241), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13011), .ZN(n13013) );
  AOI21_X1 U15255 ( .B1(n13248), .B2(n13014), .A(n13013), .ZN(n13015) );
  OAI211_X1 U15256 ( .C1(n13397), .C2(n13017), .A(n13016), .B(n13015), .ZN(
        P2_U3201) );
  OAI21_X1 U15257 ( .B1(n13020), .B2(n13019), .A(n13018), .ZN(n13021) );
  NAND2_X1 U15258 ( .A1(n13021), .A2(n14448), .ZN(n13030) );
  AOI22_X1 U15259 ( .A1(n13023), .A2(n13082), .B1(n13022), .B2(n14451), .ZN(
        n13029) );
  NAND2_X1 U15260 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n14898) );
  INV_X1 U15261 ( .A(n14898), .ZN(n13026) );
  NOR2_X1 U15262 ( .A1(n14453), .A2(n13024), .ZN(n13025) );
  AOI211_X1 U15263 ( .C1(n13027), .C2(n13084), .A(n13026), .B(n13025), .ZN(
        n13028) );
  NAND3_X1 U15264 ( .A1(n13030), .A2(n13029), .A3(n13028), .ZN(P2_U3202) );
  INV_X1 U15265 ( .A(n13031), .ZN(n13033) );
  NAND2_X1 U15266 ( .A1(n13033), .A2(n13032), .ZN(n13034) );
  XNOR2_X1 U15267 ( .A(n13035), .B(n13034), .ZN(n13040) );
  OAI22_X1 U15268 ( .A1(n13036), .A2(n14443), .B1(n13043), .B2(n14441), .ZN(
        n13303) );
  AOI22_X1 U15269 ( .A1(n13303), .A2(n14450), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13037) );
  OAI21_X1 U15270 ( .B1(n13306), .B2(n14453), .A(n13037), .ZN(n13038) );
  AOI21_X1 U15271 ( .B1(n13420), .B2(n14451), .A(n13038), .ZN(n13039) );
  OAI21_X1 U15272 ( .B1(n13040), .B2(n13059), .A(n13039), .ZN(P2_U3205) );
  XNOR2_X1 U15273 ( .A(n13042), .B(n13041), .ZN(n13050) );
  NAND2_X1 U15274 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n15048)
         );
  OAI21_X1 U15275 ( .B1(n14453), .B2(n13342), .A(n15048), .ZN(n13048) );
  OAI22_X1 U15276 ( .A1(n13046), .A2(n13045), .B1(n13044), .B2(n13043), .ZN(
        n13047) );
  AOI211_X1 U15277 ( .C1(n13429), .C2(n14451), .A(n13048), .B(n13047), .ZN(
        n13049) );
  OAI21_X1 U15278 ( .B1(n13050), .B2(n13059), .A(n13049), .ZN(P2_U3210) );
  OR2_X1 U15279 ( .A1(n13053), .A2(n14443), .ZN(n13055) );
  NAND2_X1 U15280 ( .A1(n13066), .A2(n13335), .ZN(n13054) );
  NAND2_X1 U15281 ( .A1(n13055), .A2(n13054), .ZN(n13212) );
  AOI22_X1 U15282 ( .A1(n14450), .A2(n13212), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13056) );
  OAI21_X1 U15283 ( .B1(n13217), .B2(n14453), .A(n13056), .ZN(n13057) );
  AOI21_X1 U15284 ( .B1(n13387), .B2(n14451), .A(n13057), .ZN(n13058) );
  OAI21_X1 U15285 ( .B1(n13060), .B2(n13059), .A(n13058), .ZN(P2_U3212) );
  MUX2_X1 U15286 ( .A(n13168), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13087), .Z(
        P2_U3562) );
  MUX2_X1 U15287 ( .A(n13061), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13087), .Z(
        P2_U3561) );
  MUX2_X1 U15288 ( .A(n13062), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13087), .Z(
        P2_U3560) );
  MUX2_X1 U15289 ( .A(n13063), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13087), .Z(
        P2_U3559) );
  MUX2_X1 U15290 ( .A(n13064), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13087), .Z(
        P2_U3558) );
  MUX2_X1 U15291 ( .A(n13065), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13087), .Z(
        P2_U3557) );
  MUX2_X1 U15292 ( .A(n13066), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13087), .Z(
        P2_U3556) );
  MUX2_X1 U15293 ( .A(n13067), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13087), .Z(
        P2_U3555) );
  MUX2_X1 U15294 ( .A(n13271), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13087), .Z(
        P2_U3554) );
  MUX2_X1 U15295 ( .A(n13068), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13087), .Z(
        P2_U3553) );
  MUX2_X1 U15296 ( .A(n13272), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13087), .Z(
        P2_U3552) );
  MUX2_X1 U15297 ( .A(n13069), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13087), .Z(
        P2_U3551) );
  MUX2_X1 U15298 ( .A(n13337), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13087), .Z(
        P2_U3550) );
  MUX2_X1 U15299 ( .A(n13070), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13087), .Z(
        P2_U3549) );
  INV_X2 U15300 ( .A(P2_U3947), .ZN(n13087) );
  MUX2_X1 U15301 ( .A(n13334), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13087), .Z(
        P2_U3548) );
  MUX2_X1 U15302 ( .A(n13071), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13087), .Z(
        P2_U3547) );
  MUX2_X1 U15303 ( .A(n13072), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13087), .Z(
        P2_U3546) );
  MUX2_X1 U15304 ( .A(n13073), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13087), .Z(
        P2_U3545) );
  MUX2_X1 U15305 ( .A(n13074), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13087), .Z(
        P2_U3544) );
  MUX2_X1 U15306 ( .A(n13075), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13087), .Z(
        P2_U3543) );
  MUX2_X1 U15307 ( .A(n13076), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13087), .Z(
        P2_U3542) );
  MUX2_X1 U15308 ( .A(n13077), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13087), .Z(
        P2_U3541) );
  MUX2_X1 U15309 ( .A(n13078), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13087), .Z(
        P2_U3540) );
  MUX2_X1 U15310 ( .A(n13079), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13087), .Z(
        P2_U3539) );
  MUX2_X1 U15311 ( .A(n13080), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13087), .Z(
        P2_U3538) );
  MUX2_X1 U15312 ( .A(n13081), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13087), .Z(
        P2_U3537) );
  MUX2_X1 U15313 ( .A(n13082), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13087), .Z(
        P2_U3536) );
  MUX2_X1 U15314 ( .A(n13083), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13087), .Z(
        P2_U3535) );
  MUX2_X1 U15315 ( .A(n13084), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13087), .Z(
        P2_U3534) );
  MUX2_X1 U15316 ( .A(n13085), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13087), .Z(
        P2_U3533) );
  MUX2_X1 U15317 ( .A(n13086), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13087), .Z(
        P2_U3532) );
  MUX2_X1 U15318 ( .A(n13088), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13087), .Z(
        P2_U3531) );
  NAND2_X1 U15319 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n13089) );
  OAI21_X1 U15320 ( .B1(n15046), .B2(n13090), .A(n13089), .ZN(n13091) );
  AOI21_X1 U15321 ( .B1(n14872), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n13091), .ZN(
        n13100) );
  OAI211_X1 U15322 ( .C1(n13094), .C2(n13093), .A(n15035), .B(n13092), .ZN(
        n13099) );
  OAI211_X1 U15323 ( .C1(n13097), .C2(n13096), .A(n15041), .B(n13095), .ZN(
        n13098) );
  NAND3_X1 U15324 ( .A1(n13100), .A2(n13099), .A3(n13098), .ZN(P2_U3217) );
  INV_X1 U15325 ( .A(n13101), .ZN(n13103) );
  INV_X1 U15326 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15399) );
  NOR2_X1 U15327 ( .A1(n15050), .A2(n15399), .ZN(n13102) );
  AOI211_X1 U15328 ( .C1(n15028), .C2(n13104), .A(n13103), .B(n13102), .ZN(
        n13113) );
  OAI211_X1 U15329 ( .C1(n13107), .C2(n13106), .A(n15035), .B(n13105), .ZN(
        n13112) );
  OAI211_X1 U15330 ( .C1(n13110), .C2(n13109), .A(n15041), .B(n13108), .ZN(
        n13111) );
  NAND3_X1 U15331 ( .A1(n13113), .A2(n13112), .A3(n13111), .ZN(P2_U3219) );
  AOI21_X1 U15332 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n13122), .A(n13114), 
        .ZN(n13117) );
  MUX2_X1 U15333 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n13115), .S(n13139), .Z(
        n13116) );
  NAND2_X1 U15334 ( .A1(n13117), .A2(n13116), .ZN(n13130) );
  OAI21_X1 U15335 ( .B1(n13117), .B2(n13116), .A(n13130), .ZN(n13118) );
  NAND2_X1 U15336 ( .A1(n13118), .A2(n15041), .ZN(n13129) );
  AOI21_X1 U15337 ( .B1(n15028), .B2(n13139), .A(n13119), .ZN(n13128) );
  MUX2_X1 U15338 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n13120), .S(n13139), .Z(
        n13124) );
  OAI21_X1 U15339 ( .B1(n13122), .B2(P2_REG2_REG_11__SCAN_IN), .A(n13121), 
        .ZN(n13123) );
  NAND2_X1 U15340 ( .A1(n13123), .A2(n13124), .ZN(n13138) );
  OAI21_X1 U15341 ( .B1(n13124), .B2(n13123), .A(n13138), .ZN(n13125) );
  NAND2_X1 U15342 ( .A1(n13125), .A2(n15035), .ZN(n13127) );
  NAND2_X1 U15343 ( .A1(n14872), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n13126) );
  NAND4_X1 U15344 ( .A1(n13129), .A2(n13128), .A3(n13127), .A4(n13126), .ZN(
        P2_U3226) );
  INV_X1 U15345 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13638) );
  INV_X1 U15346 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n15037) );
  OAI21_X1 U15347 ( .B1(n13139), .B2(P2_REG1_REG_12__SCAN_IN), .A(n13130), 
        .ZN(n14972) );
  MUX2_X1 U15348 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n13131), .S(n13141), .Z(
        n14973) );
  NOR2_X1 U15349 ( .A1(n14972), .A2(n14973), .ZN(n14971) );
  MUX2_X1 U15350 ( .A(n13132), .B(P2_REG1_REG_14__SCAN_IN), .S(n14988), .Z(
        n14981) );
  NOR2_X1 U15351 ( .A1(n14982), .A2(n14981), .ZN(n14980) );
  NOR2_X1 U15352 ( .A1(n13133), .A2(n13145), .ZN(n13134) );
  XNOR2_X1 U15353 ( .A(n13145), .B(n13133), .ZN(n14996) );
  NOR2_X1 U15354 ( .A1(n14995), .A2(n14996), .ZN(n14994) );
  XNOR2_X1 U15355 ( .A(n15012), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15004) );
  NOR2_X1 U15356 ( .A1(n15005), .A2(n15004), .ZN(n15003) );
  AOI21_X1 U15357 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n15012), .A(n15003), 
        .ZN(n15024) );
  XNOR2_X1 U15358 ( .A(n15027), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15023) );
  NOR2_X1 U15359 ( .A1(n15024), .A2(n15023), .ZN(n15021) );
  XNOR2_X1 U15360 ( .A(n15045), .B(n13135), .ZN(n15038) );
  NOR2_X1 U15361 ( .A1(n15037), .A2(n15038), .ZN(n15039) );
  NOR2_X1 U15362 ( .A1(n13135), .A2(n15045), .ZN(n13136) );
  NOR2_X1 U15363 ( .A1(n15039), .A2(n13136), .ZN(n13137) );
  XOR2_X1 U15364 ( .A(n13137), .B(P2_REG1_REG_19__SCAN_IN), .Z(n13158) );
  OAI21_X1 U15365 ( .B1(n13139), .B2(P2_REG2_REG_12__SCAN_IN), .A(n13138), 
        .ZN(n14969) );
  XNOR2_X1 U15366 ( .A(n13141), .B(n13140), .ZN(n14970) );
  NOR2_X1 U15367 ( .A1(n14969), .A2(n14970), .ZN(n14968) );
  AOI21_X1 U15368 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n14976), .A(n14968), 
        .ZN(n13143) );
  NOR2_X1 U15369 ( .A1(n13143), .A2(n13142), .ZN(n13144) );
  INV_X1 U15370 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n14984) );
  XNOR2_X1 U15371 ( .A(n13143), .B(n13142), .ZN(n14985) );
  NOR2_X1 U15372 ( .A1(n14984), .A2(n14985), .ZN(n14983) );
  NOR2_X1 U15373 ( .A1(n13144), .A2(n14983), .ZN(n13146) );
  NOR2_X1 U15374 ( .A1(n13146), .A2(n13145), .ZN(n13147) );
  XNOR2_X1 U15375 ( .A(n13146), .B(n13145), .ZN(n14993) );
  NOR2_X1 U15376 ( .A1(n11754), .A2(n14993), .ZN(n14992) );
  NOR2_X1 U15377 ( .A1(n13147), .A2(n14992), .ZN(n15009) );
  MUX2_X1 U15378 ( .A(n13148), .B(P2_REG2_REG_16__SCAN_IN), .S(n15012), .Z(
        n15008) );
  OR2_X1 U15379 ( .A1(n15009), .A2(n15008), .ZN(n15006) );
  NAND2_X1 U15380 ( .A1(n15012), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13149) );
  NAND2_X1 U15381 ( .A1(n15006), .A2(n13149), .ZN(n15017) );
  OR2_X1 U15382 ( .A1(n15027), .A2(n13150), .ZN(n13152) );
  NAND2_X1 U15383 ( .A1(n15027), .A2(n13150), .ZN(n13151) );
  NAND2_X1 U15384 ( .A1(n13152), .A2(n13151), .ZN(n15016) );
  AOI21_X1 U15385 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n15027), .A(n15020), 
        .ZN(n13154) );
  INV_X1 U15386 ( .A(n13154), .ZN(n13153) );
  XNOR2_X1 U15387 ( .A(n15045), .B(n13153), .ZN(n15034) );
  INV_X1 U15388 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n15033) );
  NAND2_X1 U15389 ( .A1(n15034), .A2(n15033), .ZN(n15032) );
  NAND2_X1 U15390 ( .A1(n13154), .A2(n15045), .ZN(n13155) );
  NAND2_X1 U15391 ( .A1(n15032), .A2(n13155), .ZN(n13156) );
  XNOR2_X1 U15392 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13156), .ZN(n13160) );
  INV_X1 U15393 ( .A(n13160), .ZN(n13157) );
  OAI22_X1 U15394 ( .A1(n13158), .A2(n15022), .B1(n13157), .B2(n15018), .ZN(
        n13163) );
  AOI21_X1 U15395 ( .B1(n15041), .B2(n13158), .A(n15028), .ZN(n13159) );
  OAI21_X1 U15396 ( .B1(n13160), .B2(n15018), .A(n13159), .ZN(n13162) );
  NAND2_X1 U15397 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3088), .ZN(n13164)
         );
  NAND2_X1 U15398 ( .A1(n13457), .A2(n13172), .ZN(n13171) );
  XNOR2_X1 U15399 ( .A(n13171), .B(n13451), .ZN(n13166) );
  OR2_X1 U15400 ( .A1(n13166), .A2(n9935), .ZN(n13369) );
  NAND2_X1 U15401 ( .A1(n13168), .A2(n13167), .ZN(n13373) );
  NOR2_X1 U15402 ( .A1(n13358), .A2(n13373), .ZN(n13174) );
  AOI21_X1 U15403 ( .B1(n13358), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13174), 
        .ZN(n13170) );
  NAND2_X1 U15404 ( .A1(n13451), .A2(n15058), .ZN(n13169) );
  OAI211_X1 U15405 ( .C1(n13369), .C2(n15061), .A(n13170), .B(n13169), .ZN(
        P2_U3234) );
  OAI211_X1 U15406 ( .C1(n13457), .C2(n13172), .A(n14465), .B(n13171), .ZN(
        n13374) );
  NOR2_X1 U15407 ( .A1(n13457), .A2(n13360), .ZN(n13173) );
  AOI211_X1 U15408 ( .C1(n13358), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13174), 
        .B(n13173), .ZN(n13175) );
  OAI21_X1 U15409 ( .B1(n15061), .B2(n13374), .A(n13175), .ZN(P2_U3235) );
  OR2_X1 U15410 ( .A1(n13177), .A2(n13176), .ZN(n13178) );
  NOR2_X1 U15411 ( .A1(n13182), .A2(n13340), .ZN(n13184) );
  OAI21_X1 U15412 ( .B1(n13185), .B2(n15052), .A(n13379), .ZN(n13186) );
  NAND2_X1 U15413 ( .A1(n13186), .A2(n15055), .ZN(n13193) );
  OAI21_X1 U15414 ( .B1(n13459), .B2(n13199), .A(n14465), .ZN(n13187) );
  INV_X1 U15415 ( .A(n13378), .ZN(n13191) );
  INV_X1 U15416 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13189) );
  OAI22_X1 U15417 ( .A1(n13459), .A2(n13360), .B1(n15055), .B2(n13189), .ZN(
        n13190) );
  AOI21_X1 U15418 ( .B1(n13191), .B2(n14467), .A(n13190), .ZN(n13192) );
  OAI211_X1 U15419 ( .C1(n13365), .C2(n13380), .A(n13193), .B(n13192), .ZN(
        P2_U3237) );
  XNOR2_X1 U15420 ( .A(n13194), .B(n13206), .ZN(n13197) );
  INV_X1 U15421 ( .A(n13195), .ZN(n13196) );
  AOI21_X1 U15422 ( .B1(n13197), .B2(n14456), .A(n13196), .ZN(n13384) );
  OAI21_X1 U15423 ( .B1(n13202), .B2(n13221), .A(n14465), .ZN(n13198) );
  INV_X1 U15424 ( .A(n13383), .ZN(n13204) );
  AOI22_X1 U15425 ( .A1(n13358), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n13200), 
        .B2(n14460), .ZN(n13201) );
  OAI21_X1 U15426 ( .B1(n13202), .B2(n13360), .A(n13201), .ZN(n13203) );
  AOI21_X1 U15427 ( .B1(n13204), .B2(n14467), .A(n13203), .ZN(n13209) );
  NAND2_X1 U15428 ( .A1(n13207), .A2(n13206), .ZN(n13381) );
  NAND3_X1 U15429 ( .A1(n13205), .A2(n13381), .A3(n15063), .ZN(n13208) );
  OAI211_X1 U15430 ( .C1(n13384), .C2(n13358), .A(n13209), .B(n13208), .ZN(
        P2_U3238) );
  XNOR2_X1 U15431 ( .A(n13210), .B(n13211), .ZN(n13213) );
  AOI21_X1 U15432 ( .B1(n13213), .B2(n14456), .A(n13212), .ZN(n13389) );
  XNOR2_X1 U15433 ( .A(n13214), .B(n13215), .ZN(n13390) );
  NAND2_X1 U15434 ( .A1(n13358), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n13216) );
  OAI21_X1 U15435 ( .B1(n15052), .B2(n13217), .A(n13216), .ZN(n13218) );
  AOI21_X1 U15436 ( .B1(n13387), .B2(n15058), .A(n13218), .ZN(n13223) );
  NAND2_X1 U15437 ( .A1(n13387), .A2(n13234), .ZN(n13219) );
  NAND2_X1 U15438 ( .A1(n13219), .A2(n14465), .ZN(n13220) );
  NOR2_X1 U15439 ( .A1(n13221), .A2(n13220), .ZN(n13386) );
  NAND2_X1 U15440 ( .A1(n13386), .A2(n14467), .ZN(n13222) );
  OAI211_X1 U15441 ( .C1(n13390), .C2(n13365), .A(n13223), .B(n13222), .ZN(
        n13224) );
  INV_X1 U15442 ( .A(n13224), .ZN(n13225) );
  OAI21_X1 U15443 ( .B1(n13358), .B2(n13389), .A(n13225), .ZN(P2_U3239) );
  XNOR2_X1 U15444 ( .A(n13226), .B(n13230), .ZN(n13228) );
  AOI21_X1 U15445 ( .B1(n13228), .B2(n14456), .A(n13227), .ZN(n13394) );
  XOR2_X1 U15446 ( .A(n13230), .B(n13229), .Z(n13395) );
  NAND2_X1 U15447 ( .A1(n13358), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n13231) );
  OAI21_X1 U15448 ( .B1(n15052), .B2(n13232), .A(n13231), .ZN(n13233) );
  AOI21_X1 U15449 ( .B1(n13392), .B2(n15058), .A(n13233), .ZN(n13237) );
  AOI21_X1 U15450 ( .B1(n13392), .B2(n13247), .A(n9935), .ZN(n13235) );
  AND2_X1 U15451 ( .A1(n13235), .A2(n13234), .ZN(n13391) );
  NAND2_X1 U15452 ( .A1(n13391), .A2(n14467), .ZN(n13236) );
  OAI211_X1 U15453 ( .C1(n13395), .C2(n13365), .A(n13237), .B(n13236), .ZN(
        n13238) );
  INV_X1 U15454 ( .A(n13238), .ZN(n13239) );
  OAI21_X1 U15455 ( .B1(n13358), .B2(n13394), .A(n13239), .ZN(P2_U3240) );
  XOR2_X1 U15456 ( .A(n13240), .B(n13246), .Z(n13242) );
  OAI21_X1 U15457 ( .B1(n13242), .B2(n13340), .A(n13241), .ZN(n13398) );
  INV_X1 U15458 ( .A(n13398), .ZN(n13254) );
  INV_X1 U15459 ( .A(n13243), .ZN(n13244) );
  AOI21_X1 U15460 ( .B1(n13246), .B2(n13245), .A(n13244), .ZN(n13400) );
  OAI211_X1 U15461 ( .C1(n13397), .C2(n13256), .A(n14465), .B(n13247), .ZN(
        n13396) );
  AOI22_X1 U15462 ( .A1(n13358), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13248), 
        .B2(n14460), .ZN(n13251) );
  NAND2_X1 U15463 ( .A1(n13249), .A2(n15058), .ZN(n13250) );
  OAI211_X1 U15464 ( .C1(n13396), .C2(n15061), .A(n13251), .B(n13250), .ZN(
        n13252) );
  AOI21_X1 U15465 ( .B1(n13400), .B2(n15063), .A(n13252), .ZN(n13253) );
  OAI21_X1 U15466 ( .B1(n13358), .B2(n13254), .A(n13253), .ZN(P2_U3241) );
  XOR2_X1 U15467 ( .A(n13255), .B(n13259), .Z(n13407) );
  AOI211_X1 U15468 ( .C1(n13404), .C2(n13274), .A(n9935), .B(n13256), .ZN(
        n13402) );
  OAI22_X1 U15469 ( .A1(n7088), .A2(n13360), .B1(n15055), .B2(n13257), .ZN(
        n13258) );
  AOI21_X1 U15470 ( .B1(n13402), .B2(n14467), .A(n13258), .ZN(n13268) );
  XOR2_X1 U15471 ( .A(n13260), .B(n13259), .Z(n13261) );
  NAND2_X1 U15472 ( .A1(n13261), .A2(n14456), .ZN(n13405) );
  OAI22_X1 U15473 ( .A1(n13263), .A2(n14441), .B1(n13262), .B2(n14443), .ZN(
        n13403) );
  INV_X1 U15474 ( .A(n13403), .ZN(n13264) );
  OAI211_X1 U15475 ( .C1(n15052), .C2(n13265), .A(n13405), .B(n13264), .ZN(
        n13266) );
  NAND2_X1 U15476 ( .A1(n13266), .A2(n15055), .ZN(n13267) );
  OAI211_X1 U15477 ( .C1(n13407), .C2(n13365), .A(n13268), .B(n13267), .ZN(
        P2_U3242) );
  XNOR2_X1 U15478 ( .A(n13270), .B(n13269), .ZN(n13273) );
  AOI222_X1 U15479 ( .A1(n14456), .A2(n13273), .B1(n13272), .B2(n13335), .C1(
        n13271), .C2(n13336), .ZN(n13411) );
  INV_X1 U15480 ( .A(n13274), .ZN(n13275) );
  AOI211_X1 U15481 ( .C1(n13409), .C2(n13292), .A(n9942), .B(n13275), .ZN(
        n13408) );
  INV_X1 U15482 ( .A(n13276), .ZN(n13277) );
  AOI22_X1 U15483 ( .A1(n13358), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13277), 
        .B2(n14460), .ZN(n13278) );
  OAI21_X1 U15484 ( .B1(n13279), .B2(n13360), .A(n13278), .ZN(n13285) );
  NAND2_X1 U15485 ( .A1(n13281), .A2(n13280), .ZN(n13282) );
  NAND2_X1 U15486 ( .A1(n13283), .A2(n13282), .ZN(n13412) );
  NOR2_X1 U15487 ( .A1(n13412), .A2(n13365), .ZN(n13284) );
  AOI211_X1 U15488 ( .C1(n13408), .C2(n14467), .A(n13285), .B(n13284), .ZN(
        n13286) );
  OAI21_X1 U15489 ( .B1(n13358), .B2(n13411), .A(n13286), .ZN(P2_U3243) );
  XOR2_X1 U15490 ( .A(n13287), .B(n13290), .Z(n13289) );
  OAI21_X1 U15491 ( .B1(n13289), .B2(n13340), .A(n13288), .ZN(n13413) );
  INV_X1 U15492 ( .A(n13413), .ZN(n13301) );
  XNOR2_X1 U15493 ( .A(n13291), .B(n13290), .ZN(n13415) );
  INV_X1 U15494 ( .A(n13305), .ZN(n13294) );
  INV_X1 U15495 ( .A(n13292), .ZN(n13293) );
  AOI211_X1 U15496 ( .C1(n13295), .C2(n13294), .A(n9935), .B(n13293), .ZN(
        n13414) );
  NAND2_X1 U15497 ( .A1(n13414), .A2(n14467), .ZN(n13298) );
  AOI22_X1 U15498 ( .A1(n13358), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13296), 
        .B2(n14460), .ZN(n13297) );
  OAI211_X1 U15499 ( .C1(n13469), .C2(n13360), .A(n13298), .B(n13297), .ZN(
        n13299) );
  AOI21_X1 U15500 ( .B1(n13415), .B2(n15063), .A(n13299), .ZN(n13300) );
  OAI21_X1 U15501 ( .B1(n13301), .B2(n13358), .A(n13300), .ZN(P2_U3244) );
  XNOR2_X1 U15502 ( .A(n13302), .B(n13310), .ZN(n13304) );
  AOI21_X1 U15503 ( .B1(n13304), .B2(n14456), .A(n13303), .ZN(n13422) );
  AOI211_X1 U15504 ( .C1(n13420), .C2(n13321), .A(n9935), .B(n13305), .ZN(
        n13419) );
  INV_X1 U15505 ( .A(n13420), .ZN(n13309) );
  INV_X1 U15506 ( .A(n13306), .ZN(n13307) );
  AOI22_X1 U15507 ( .A1(n13358), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13307), 
        .B2(n14460), .ZN(n13308) );
  OAI21_X1 U15508 ( .B1(n13309), .B2(n13360), .A(n13308), .ZN(n13313) );
  XNOR2_X1 U15509 ( .A(n13311), .B(n13310), .ZN(n13423) );
  NOR2_X1 U15510 ( .A1(n13423), .A2(n13365), .ZN(n13312) );
  AOI211_X1 U15511 ( .C1(n13419), .C2(n14467), .A(n13313), .B(n13312), .ZN(
        n13314) );
  OAI21_X1 U15512 ( .B1(n13358), .B2(n13422), .A(n13314), .ZN(P2_U3245) );
  XNOR2_X1 U15513 ( .A(n13316), .B(n13317), .ZN(n13428) );
  XOR2_X1 U15514 ( .A(n13318), .B(n13317), .Z(n13320) );
  OAI21_X1 U15515 ( .B1(n13320), .B2(n13340), .A(n13319), .ZN(n13424) );
  NAND2_X1 U15516 ( .A1(n13424), .A2(n15055), .ZN(n13327) );
  INV_X1 U15517 ( .A(n13321), .ZN(n13322) );
  AOI211_X1 U15518 ( .C1(n13426), .C2(n7093), .A(n9935), .B(n13322), .ZN(
        n13425) );
  AOI22_X1 U15519 ( .A1(n13358), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13323), 
        .B2(n14460), .ZN(n13324) );
  OAI21_X1 U15520 ( .B1(n8200), .B2(n13360), .A(n13324), .ZN(n13325) );
  AOI21_X1 U15521 ( .B1(n13425), .B2(n14467), .A(n13325), .ZN(n13326) );
  OAI211_X1 U15522 ( .C1(n13365), .C2(n13428), .A(n13327), .B(n13326), .ZN(
        P2_U3246) );
  OR2_X1 U15523 ( .A1(n13328), .A2(n13332), .ZN(n13329) );
  NAND2_X1 U15524 ( .A1(n13330), .A2(n13329), .ZN(n13430) );
  INV_X1 U15525 ( .A(n13430), .ZN(n13349) );
  XNOR2_X1 U15526 ( .A(n13331), .B(n13332), .ZN(n13341) );
  NAND2_X1 U15527 ( .A1(n13430), .A2(n13333), .ZN(n13339) );
  AOI22_X1 U15528 ( .A1(n13337), .A2(n13336), .B1(n13335), .B2(n13334), .ZN(
        n13338) );
  OAI211_X1 U15529 ( .C1(n13341), .C2(n13340), .A(n13339), .B(n13338), .ZN(
        n13435) );
  NAND2_X1 U15530 ( .A1(n13435), .A2(n15055), .ZN(n13347) );
  OAI22_X1 U15531 ( .A1(n15055), .A2(n15033), .B1(n13342), .B2(n15052), .ZN(
        n13345) );
  AOI21_X1 U15532 ( .B1(n13429), .B2(n13353), .A(n9935), .ZN(n13343) );
  NAND2_X1 U15533 ( .A1(n13343), .A2(n7093), .ZN(n13431) );
  NOR2_X1 U15534 ( .A1(n13431), .A2(n15061), .ZN(n13344) );
  AOI211_X1 U15535 ( .C1(n15058), .C2(n13429), .A(n13345), .B(n13344), .ZN(
        n13346) );
  OAI211_X1 U15536 ( .C1(n13349), .C2(n13348), .A(n13347), .B(n13346), .ZN(
        P2_U3247) );
  XOR2_X1 U15537 ( .A(n13363), .B(n13350), .Z(n13352) );
  AOI21_X1 U15538 ( .B1(n13352), .B2(n14456), .A(n13351), .ZN(n13439) );
  INV_X1 U15539 ( .A(n13353), .ZN(n13354) );
  AOI211_X1 U15540 ( .C1(n13437), .C2(n13355), .A(n9935), .B(n13354), .ZN(
        n13436) );
  INV_X1 U15541 ( .A(n13437), .ZN(n13361) );
  INV_X1 U15542 ( .A(n13356), .ZN(n13357) );
  AOI22_X1 U15543 ( .A1(n13358), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13357), 
        .B2(n14460), .ZN(n13359) );
  OAI21_X1 U15544 ( .B1(n13361), .B2(n13360), .A(n13359), .ZN(n13367) );
  XOR2_X1 U15545 ( .A(n13364), .B(n13363), .Z(n13441) );
  NOR2_X1 U15546 ( .A1(n13441), .A2(n13365), .ZN(n13366) );
  AOI211_X1 U15547 ( .C1(n13436), .C2(n14467), .A(n13367), .B(n13366), .ZN(
        n13368) );
  OAI21_X1 U15548 ( .B1(n13358), .B2(n13439), .A(n13368), .ZN(P2_U3248) );
  NAND2_X1 U15549 ( .A1(n13369), .A2(n13373), .ZN(n13449) );
  MUX2_X1 U15550 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13449), .S(n15105), .Z(
        n13370) );
  AOI21_X1 U15551 ( .B1(n13371), .B2(n13451), .A(n13370), .ZN(n13372) );
  INV_X1 U15552 ( .A(n13372), .ZN(P2_U3530) );
  AND2_X1 U15553 ( .A1(n13374), .A2(n13373), .ZN(n13455) );
  MUX2_X1 U15554 ( .A(n13455), .B(n13375), .S(n15103), .Z(n13376) );
  OAI21_X1 U15555 ( .B1(n13457), .B2(n13418), .A(n13376), .ZN(P2_U3529) );
  MUX2_X1 U15556 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13377), .S(n15105), .Z(
        P2_U3528) );
  NAND3_X1 U15557 ( .A1(n13205), .A2(n14479), .A3(n13381), .ZN(n13385) );
  NAND2_X1 U15558 ( .A1(n7105), .A2(n14481), .ZN(n13382) );
  NAND4_X1 U15559 ( .A1(n13385), .A2(n13384), .A3(n13383), .A4(n13382), .ZN(
        n13460) );
  MUX2_X1 U15560 ( .A(n13460), .B(P2_REG1_REG_27__SCAN_IN), .S(n15103), .Z(
        P2_U3526) );
  AOI21_X1 U15561 ( .B1(n14481), .B2(n13387), .A(n13386), .ZN(n13388) );
  OAI211_X1 U15562 ( .C1(n13390), .C2(n13440), .A(n13389), .B(n13388), .ZN(
        n13461) );
  MUX2_X1 U15563 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13461), .S(n15105), .Z(
        P2_U3525) );
  AOI21_X1 U15564 ( .B1(n14481), .B2(n13392), .A(n13391), .ZN(n13393) );
  OAI211_X1 U15565 ( .C1(n13395), .C2(n13440), .A(n13394), .B(n13393), .ZN(
        n13462) );
  MUX2_X1 U15566 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13462), .S(n15105), .Z(
        P2_U3524) );
  INV_X1 U15567 ( .A(n14481), .ZN(n15092) );
  OAI21_X1 U15568 ( .B1(n13397), .B2(n15092), .A(n13396), .ZN(n13399) );
  AOI211_X1 U15569 ( .C1(n13400), .C2(n14479), .A(n13399), .B(n13398), .ZN(
        n13401) );
  INV_X1 U15570 ( .A(n13401), .ZN(n13463) );
  MUX2_X1 U15571 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13463), .S(n15105), .Z(
        P2_U3523) );
  AOI211_X1 U15572 ( .C1(n14481), .C2(n13404), .A(n13403), .B(n13402), .ZN(
        n13406) );
  OAI211_X1 U15573 ( .C1(n13407), .C2(n13440), .A(n13406), .B(n13405), .ZN(
        n13464) );
  MUX2_X1 U15574 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13464), .S(n15105), .Z(
        P2_U3522) );
  AOI21_X1 U15575 ( .B1(n14481), .B2(n13409), .A(n13408), .ZN(n13410) );
  OAI211_X1 U15576 ( .C1(n13440), .C2(n13412), .A(n13411), .B(n13410), .ZN(
        n13465) );
  MUX2_X1 U15577 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13465), .S(n15105), .Z(
        P2_U3521) );
  INV_X1 U15578 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13416) );
  AOI211_X1 U15579 ( .C1(n14479), .C2(n13415), .A(n13414), .B(n13413), .ZN(
        n13466) );
  MUX2_X1 U15580 ( .A(n13416), .B(n13466), .S(n15105), .Z(n13417) );
  OAI21_X1 U15581 ( .B1(n13469), .B2(n13418), .A(n13417), .ZN(P2_U3520) );
  AOI21_X1 U15582 ( .B1(n14481), .B2(n13420), .A(n13419), .ZN(n13421) );
  OAI211_X1 U15583 ( .C1(n13440), .C2(n13423), .A(n13422), .B(n13421), .ZN(
        n13470) );
  MUX2_X1 U15584 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13470), .S(n15105), .Z(
        P2_U3519) );
  AOI211_X1 U15585 ( .C1(n14481), .C2(n13426), .A(n13425), .B(n13424), .ZN(
        n13427) );
  OAI21_X1 U15586 ( .B1(n13440), .B2(n13428), .A(n13427), .ZN(n13471) );
  MUX2_X1 U15587 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13471), .S(n15105), .Z(
        P2_U3518) );
  INV_X1 U15588 ( .A(n13429), .ZN(n13433) );
  NAND2_X1 U15589 ( .A1(n13430), .A2(n15097), .ZN(n13432) );
  OAI211_X1 U15590 ( .C1(n13433), .C2(n15092), .A(n13432), .B(n13431), .ZN(
        n13434) );
  OR2_X1 U15591 ( .A1(n13435), .A2(n13434), .ZN(n13472) );
  MUX2_X1 U15592 ( .A(n13472), .B(P2_REG1_REG_18__SCAN_IN), .S(n15103), .Z(
        P2_U3517) );
  AOI21_X1 U15593 ( .B1(n14481), .B2(n13437), .A(n13436), .ZN(n13438) );
  OAI211_X1 U15594 ( .C1(n13441), .C2(n13440), .A(n13439), .B(n13438), .ZN(
        n13473) );
  MUX2_X1 U15595 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13473), .S(n15105), .Z(
        P2_U3516) );
  AND3_X1 U15596 ( .A1(n13442), .A2(n13443), .A3(n14479), .ZN(n13447) );
  OAI21_X1 U15597 ( .B1(n13445), .B2(n15092), .A(n13444), .ZN(n13446) );
  MUX2_X1 U15598 ( .A(n13474), .B(P2_REG1_REG_16__SCAN_IN), .S(n15103), .Z(
        P2_U3515) );
  MUX2_X1 U15599 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13449), .S(n15099), .Z(
        n13450) );
  AOI21_X1 U15600 ( .B1(n13452), .B2(n13451), .A(n13450), .ZN(n13453) );
  INV_X1 U15601 ( .A(n13453), .ZN(P2_U3498) );
  INV_X1 U15602 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13454) );
  MUX2_X1 U15603 ( .A(n13455), .B(n13454), .S(n15098), .Z(n13456) );
  OAI21_X1 U15604 ( .B1(n13457), .B2(n13468), .A(n13456), .ZN(P2_U3497) );
  MUX2_X1 U15605 ( .A(n13460), .B(P2_REG0_REG_27__SCAN_IN), .S(n15098), .Z(
        P2_U3494) );
  MUX2_X1 U15606 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13461), .S(n15099), .Z(
        P2_U3493) );
  MUX2_X1 U15607 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13462), .S(n15099), .Z(
        P2_U3492) );
  MUX2_X1 U15608 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13463), .S(n15099), .Z(
        P2_U3491) );
  MUX2_X1 U15609 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13464), .S(n15099), .Z(
        P2_U3490) );
  MUX2_X1 U15610 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13465), .S(n15099), .Z(
        P2_U3489) );
  MUX2_X1 U15611 ( .A(n13709), .B(n13466), .S(n15099), .Z(n13467) );
  OAI21_X1 U15612 ( .B1(n13469), .B2(n13468), .A(n13467), .ZN(P2_U3488) );
  MUX2_X1 U15613 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13470), .S(n15099), .Z(
        P2_U3487) );
  MUX2_X1 U15614 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13471), .S(n15099), .Z(
        P2_U3486) );
  MUX2_X1 U15615 ( .A(n13472), .B(P2_REG0_REG_18__SCAN_IN), .S(n15098), .Z(
        P2_U3484) );
  MUX2_X1 U15616 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13473), .S(n15099), .Z(
        P2_U3481) );
  MUX2_X1 U15617 ( .A(n13474), .B(P2_REG0_REG_16__SCAN_IN), .S(n15098), .Z(
        P2_U3478) );
  NAND3_X1 U15618 ( .A1(n13476), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13478) );
  OAI22_X1 U15619 ( .A1(n13475), .A2(n13478), .B1(n13477), .B2(n13776), .ZN(
        n13479) );
  AOI21_X1 U15620 ( .B1(n14285), .B2(n6726), .A(n13479), .ZN(n13480) );
  INV_X1 U15621 ( .A(n13480), .ZN(P2_U3296) );
  AOI21_X1 U15622 ( .B1(n13769), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13481), 
        .ZN(n13482) );
  OAI21_X1 U15623 ( .B1(n13483), .B2(n11134), .A(n13482), .ZN(P2_U3299) );
  INV_X1 U15624 ( .A(n14293), .ZN(n13485) );
  OAI222_X1 U15625 ( .A1(n13776), .A2(n13486), .B1(n11134), .B2(n13485), .C1(
        P2_U3088), .C2(n6740), .ZN(P2_U3300) );
  INV_X1 U15626 ( .A(keyinput107), .ZN(n13500) );
  NOR4_X1 U15627 ( .A1(keyinput9), .A2(keyinput55), .A3(keyinput38), .A4(
        keyinput51), .ZN(n13487) );
  NAND3_X1 U15628 ( .A1(keyinput18), .A2(keyinput19), .A3(n13487), .ZN(n13499)
         );
  INV_X1 U15629 ( .A(keyinput95), .ZN(n13488) );
  NAND4_X1 U15630 ( .A1(keyinput10), .A2(keyinput110), .A3(keyinput81), .A4(
        n13488), .ZN(n13489) );
  NOR3_X1 U15631 ( .A1(keyinput60), .A2(keyinput68), .A3(n13489), .ZN(n13497)
         );
  NOR4_X1 U15632 ( .A1(keyinput78), .A2(keyinput98), .A3(keyinput47), .A4(
        keyinput36), .ZN(n13490) );
  NAND3_X1 U15633 ( .A1(keyinput109), .A2(keyinput79), .A3(n13490), .ZN(n13495) );
  NOR2_X1 U15634 ( .A1(keyinput125), .A2(keyinput24), .ZN(n13491) );
  NAND3_X1 U15635 ( .A1(keyinput0), .A2(keyinput84), .A3(n13491), .ZN(n13494)
         );
  NOR2_X1 U15636 ( .A1(keyinput91), .A2(keyinput48), .ZN(n13492) );
  NAND3_X1 U15637 ( .A1(keyinput120), .A2(keyinput14), .A3(n13492), .ZN(n13493) );
  NOR4_X1 U15638 ( .A1(keyinput16), .A2(n13495), .A3(n13494), .A4(n13493), 
        .ZN(n13496) );
  NAND4_X1 U15639 ( .A1(keyinput88), .A2(keyinput40), .A3(n13497), .A4(n13496), 
        .ZN(n13498) );
  NOR4_X1 U15640 ( .A1(keyinput86), .A2(n13500), .A3(n13499), .A4(n13498), 
        .ZN(n13547) );
  NOR2_X1 U15641 ( .A1(keyinput67), .A2(keyinput96), .ZN(n13501) );
  NAND3_X1 U15642 ( .A1(keyinput97), .A2(keyinput56), .A3(n13501), .ZN(n13545)
         );
  NOR2_X1 U15643 ( .A1(keyinput115), .A2(keyinput32), .ZN(n13502) );
  NAND3_X1 U15644 ( .A1(keyinput74), .A2(keyinput37), .A3(n13502), .ZN(n13544)
         );
  NOR2_X1 U15645 ( .A1(keyinput75), .A2(keyinput92), .ZN(n13503) );
  NAND3_X1 U15646 ( .A1(keyinput25), .A2(keyinput1), .A3(n13503), .ZN(n13504)
         );
  NOR3_X1 U15647 ( .A1(keyinput114), .A2(keyinput123), .A3(n13504), .ZN(n13513) );
  NOR2_X1 U15648 ( .A1(keyinput116), .A2(keyinput52), .ZN(n13505) );
  NAND3_X1 U15649 ( .A1(keyinput118), .A2(keyinput29), .A3(n13505), .ZN(n13511) );
  INV_X1 U15650 ( .A(keyinput100), .ZN(n13506) );
  NAND4_X1 U15651 ( .A1(keyinput83), .A2(keyinput117), .A3(keyinput17), .A4(
        n13506), .ZN(n13510) );
  NOR2_X1 U15652 ( .A1(keyinput46), .A2(keyinput44), .ZN(n13507) );
  NAND3_X1 U15653 ( .A1(keyinput20), .A2(keyinput53), .A3(n13507), .ZN(n13509)
         );
  NAND4_X1 U15654 ( .A1(keyinput8), .A2(keyinput93), .A3(keyinput63), .A4(
        keyinput66), .ZN(n13508) );
  NOR4_X1 U15655 ( .A1(n13511), .A2(n13510), .A3(n13509), .A4(n13508), .ZN(
        n13512) );
  NAND4_X1 U15656 ( .A1(keyinput111), .A2(keyinput104), .A3(n13513), .A4(
        n13512), .ZN(n13543) );
  NAND2_X1 U15657 ( .A1(keyinput12), .A2(keyinput7), .ZN(n13514) );
  NOR3_X1 U15658 ( .A1(keyinput82), .A2(keyinput49), .A3(n13514), .ZN(n13541)
         );
  NOR4_X1 U15659 ( .A1(keyinput22), .A2(keyinput113), .A3(keyinput41), .A4(
        keyinput6), .ZN(n13540) );
  NOR2_X1 U15660 ( .A1(keyinput90), .A2(keyinput35), .ZN(n13515) );
  NAND3_X1 U15661 ( .A1(keyinput33), .A2(keyinput122), .A3(n13515), .ZN(n13516) );
  NOR3_X1 U15662 ( .A1(keyinput94), .A2(keyinput72), .A3(n13516), .ZN(n13524)
         );
  INV_X1 U15663 ( .A(keyinput5), .ZN(n13672) );
  NAND4_X1 U15664 ( .A1(keyinput57), .A2(keyinput43), .A3(keyinput13), .A4(
        n13672), .ZN(n13522) );
  NOR2_X1 U15665 ( .A1(keyinput39), .A2(keyinput65), .ZN(n13517) );
  NAND3_X1 U15666 ( .A1(keyinput2), .A2(keyinput121), .A3(n13517), .ZN(n13521)
         );
  NAND4_X1 U15667 ( .A1(keyinput126), .A2(keyinput21), .A3(keyinput70), .A4(
        keyinput99), .ZN(n13520) );
  NOR2_X1 U15668 ( .A1(keyinput77), .A2(keyinput28), .ZN(n13518) );
  NAND3_X1 U15669 ( .A1(keyinput23), .A2(keyinput61), .A3(n13518), .ZN(n13519)
         );
  NOR4_X1 U15670 ( .A1(n13522), .A2(n13521), .A3(n13520), .A4(n13519), .ZN(
        n13523) );
  AND4_X1 U15671 ( .A1(keyinput87), .A2(keyinput59), .A3(n13524), .A4(n13523), 
        .ZN(n13539) );
  NAND2_X1 U15672 ( .A1(keyinput119), .A2(keyinput15), .ZN(n13525) );
  NOR3_X1 U15673 ( .A1(keyinput34), .A2(keyinput64), .A3(n13525), .ZN(n13526)
         );
  NAND3_X1 U15674 ( .A1(keyinput11), .A2(keyinput112), .A3(n13526), .ZN(n13537) );
  NAND4_X1 U15675 ( .A1(keyinput85), .A2(keyinput73), .A3(keyinput76), .A4(
        keyinput30), .ZN(n13527) );
  NOR3_X1 U15676 ( .A1(keyinput50), .A2(keyinput108), .A3(n13527), .ZN(n13535)
         );
  OR4_X1 U15677 ( .A1(keyinput54), .A2(keyinput69), .A3(keyinput62), .A4(
        keyinput124), .ZN(n13533) );
  INV_X1 U15678 ( .A(keyinput45), .ZN(n13528) );
  NAND4_X1 U15679 ( .A1(keyinput80), .A2(keyinput27), .A3(keyinput102), .A4(
        n13528), .ZN(n13532) );
  NAND4_X1 U15680 ( .A1(keyinput103), .A2(keyinput89), .A3(keyinput71), .A4(
        keyinput3), .ZN(n13531) );
  NOR2_X1 U15681 ( .A1(keyinput26), .A2(keyinput105), .ZN(n13529) );
  NAND3_X1 U15682 ( .A1(keyinput106), .A2(keyinput31), .A3(n13529), .ZN(n13530) );
  NOR4_X1 U15683 ( .A1(n13533), .A2(n13532), .A3(n13531), .A4(n13530), .ZN(
        n13534) );
  NAND4_X1 U15684 ( .A1(keyinput4), .A2(keyinput58), .A3(n13535), .A4(n13534), 
        .ZN(n13536) );
  NOR4_X1 U15685 ( .A1(keyinput42), .A2(keyinput101), .A3(n13537), .A4(n13536), 
        .ZN(n13538) );
  NAND4_X1 U15686 ( .A1(n13541), .A2(n13540), .A3(n13539), .A4(n13538), .ZN(
        n13542) );
  NOR4_X1 U15687 ( .A1(n13545), .A2(n13544), .A3(n13543), .A4(n13542), .ZN(
        n13546) );
  AOI21_X1 U15688 ( .B1(n13547), .B2(n13546), .A(keyinput127), .ZN(n13767) );
  AOI22_X1 U15689 ( .A1(n7556), .A2(keyinput80), .B1(keyinput54), .B2(n13549), 
        .ZN(n13548) );
  OAI221_X1 U15690 ( .B1(n7556), .B2(keyinput80), .C1(n13549), .C2(keyinput54), 
        .A(n13548), .ZN(n13557) );
  INV_X1 U15691 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n14754) );
  INV_X1 U15692 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14614) );
  AOI22_X1 U15693 ( .A1(n14754), .A2(keyinput69), .B1(keyinput45), .B2(n14614), 
        .ZN(n13550) );
  OAI221_X1 U15694 ( .B1(n14754), .B2(keyinput69), .C1(n14614), .C2(keyinput45), .A(n13550), .ZN(n13556) );
  AOI22_X1 U15695 ( .A1(n15155), .A2(keyinput102), .B1(n12557), .B2(keyinput62), .ZN(n13551) );
  OAI221_X1 U15696 ( .B1(n15155), .B2(keyinput102), .C1(n12557), .C2(
        keyinput62), .A(n13551), .ZN(n13555) );
  AOI22_X1 U15697 ( .A1(n13553), .A2(keyinput124), .B1(keyinput11), .B2(n9340), 
        .ZN(n13552) );
  OAI221_X1 U15698 ( .B1(n13553), .B2(keyinput124), .C1(n9340), .C2(keyinput11), .A(n13552), .ZN(n13554) );
  NOR4_X1 U15699 ( .A1(n13557), .A2(n13556), .A3(n13555), .A4(n13554), .ZN(
        n13593) );
  AOI22_X1 U15700 ( .A1(n13120), .A2(keyinput112), .B1(keyinput42), .B2(n14914), .ZN(n13558) );
  OAI221_X1 U15701 ( .B1(n13120), .B2(keyinput112), .C1(n14914), .C2(
        keyinput42), .A(n13558), .ZN(n13568) );
  AOI22_X1 U15702 ( .A1(n13560), .A2(keyinput34), .B1(keyinput119), .B2(n9327), 
        .ZN(n13559) );
  OAI221_X1 U15703 ( .B1(n13560), .B2(keyinput34), .C1(n9327), .C2(keyinput119), .A(n13559), .ZN(n13567) );
  XOR2_X1 U15704 ( .A(n13561), .B(keyinput15), .Z(n13565) );
  XNOR2_X1 U15705 ( .A(SI_6_), .B(keyinput101), .ZN(n13564) );
  XNOR2_X1 U15706 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput64), .ZN(n13563)
         );
  XNOR2_X1 U15707 ( .A(P3_IR_REG_6__SCAN_IN), .B(keyinput4), .ZN(n13562) );
  NAND4_X1 U15708 ( .A1(n13565), .A2(n13564), .A3(n13563), .A4(n13562), .ZN(
        n13566) );
  NOR3_X1 U15709 ( .A1(n13568), .A2(n13567), .A3(n13566), .ZN(n13592) );
  INV_X1 U15710 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n14757) );
  INV_X1 U15711 ( .A(keyinput30), .ZN(n13570) );
  AOI22_X1 U15712 ( .A1(n14757), .A2(keyinput26), .B1(P3_DATAO_REG_7__SCAN_IN), 
        .B2(n13570), .ZN(n13569) );
  OAI221_X1 U15713 ( .B1(n14757), .B2(keyinput26), .C1(n13570), .C2(
        P3_DATAO_REG_7__SCAN_IN), .A(n13569), .ZN(n13578) );
  INV_X1 U15714 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n14752) );
  AOI22_X1 U15715 ( .A1(n15033), .A2(keyinput58), .B1(keyinput85), .B2(n14752), 
        .ZN(n13571) );
  OAI221_X1 U15716 ( .B1(n15033), .B2(keyinput58), .C1(n14752), .C2(keyinput85), .A(n13571), .ZN(n13577) );
  INV_X1 U15717 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n14753) );
  AOI22_X1 U15718 ( .A1(n10083), .A2(keyinput108), .B1(n14753), .B2(keyinput76), .ZN(n13572) );
  OAI221_X1 U15719 ( .B1(n10083), .B2(keyinput108), .C1(n14753), .C2(
        keyinput76), .A(n13572), .ZN(n13576) );
  XNOR2_X1 U15720 ( .A(P3_REG0_REG_19__SCAN_IN), .B(keyinput73), .ZN(n13574)
         );
  XNOR2_X1 U15721 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput50), .ZN(n13573) );
  NAND2_X1 U15722 ( .A1(n13574), .A2(n13573), .ZN(n13575) );
  NOR4_X1 U15723 ( .A1(n13578), .A2(n13577), .A3(n13576), .A4(n13575), .ZN(
        n13591) );
  AOI22_X1 U15724 ( .A1(n13580), .A2(keyinput3), .B1(keyinput31), .B2(n10122), 
        .ZN(n13579) );
  OAI221_X1 U15725 ( .B1(n13580), .B2(keyinput3), .C1(n10122), .C2(keyinput31), 
        .A(n13579), .ZN(n13589) );
  AOI22_X1 U15726 ( .A1(n13582), .A2(keyinput105), .B1(keyinput74), .B2(n9241), 
        .ZN(n13581) );
  OAI221_X1 U15727 ( .B1(n13582), .B2(keyinput105), .C1(n9241), .C2(keyinput74), .A(n13581), .ZN(n13588) );
  XOR2_X1 U15728 ( .A(n8124), .B(keyinput89), .Z(n13586) );
  XNOR2_X1 U15729 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput103), .ZN(n13585) );
  XNOR2_X1 U15730 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput106), .ZN(n13584)
         );
  XNOR2_X1 U15731 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput71), .ZN(n13583)
         );
  NAND4_X1 U15732 ( .A1(n13586), .A2(n13585), .A3(n13584), .A4(n13583), .ZN(
        n13587) );
  NOR3_X1 U15733 ( .A1(n13589), .A2(n13588), .A3(n13587), .ZN(n13590) );
  NAND4_X1 U15734 ( .A1(n13593), .A2(n13592), .A3(n13591), .A4(n13590), .ZN(
        n13765) );
  AOI22_X1 U15735 ( .A1(n13595), .A2(keyinput37), .B1(keyinput67), .B2(n8368), 
        .ZN(n13594) );
  OAI221_X1 U15736 ( .B1(n13595), .B2(keyinput37), .C1(n8368), .C2(keyinput67), 
        .A(n13594), .ZN(n13605) );
  INV_X1 U15737 ( .A(keyinput114), .ZN(n13597) );
  AOI22_X1 U15738 ( .A1(n13598), .A2(keyinput56), .B1(P3_DATAO_REG_20__SCAN_IN), .B2(n13597), .ZN(n13596) );
  OAI221_X1 U15739 ( .B1(n13598), .B2(keyinput56), .C1(n13597), .C2(
        P3_DATAO_REG_20__SCAN_IN), .A(n13596), .ZN(n13604) );
  XNOR2_X1 U15740 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput115), .ZN(n13602) );
  XNOR2_X1 U15741 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput32), .ZN(n13601)
         );
  XNOR2_X1 U15742 ( .A(P3_REG2_REG_0__SCAN_IN), .B(keyinput96), .ZN(n13600) );
  XNOR2_X1 U15743 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput97), .ZN(n13599)
         );
  NAND4_X1 U15744 ( .A1(n13602), .A2(n13601), .A3(n13600), .A4(n13599), .ZN(
        n13603) );
  NOR3_X1 U15745 ( .A1(n13605), .A2(n13604), .A3(n13603), .ZN(n13646) );
  INV_X1 U15746 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n14758) );
  AOI22_X1 U15747 ( .A1(n14758), .A2(keyinput123), .B1(n9303), .B2(keyinput111), .ZN(n13606) );
  OAI221_X1 U15748 ( .B1(n14758), .B2(keyinput123), .C1(n9303), .C2(
        keyinput111), .A(n13606), .ZN(n13616) );
  INV_X1 U15749 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15070) );
  AOI22_X1 U15750 ( .A1(n15070), .A2(keyinput104), .B1(keyinput75), .B2(n13608), .ZN(n13607) );
  OAI221_X1 U15751 ( .B1(n15070), .B2(keyinput104), .C1(n13608), .C2(
        keyinput75), .A(n13607), .ZN(n13615) );
  AOI22_X1 U15752 ( .A1(n13611), .A2(keyinput25), .B1(keyinput92), .B2(n13610), 
        .ZN(n13609) );
  OAI221_X1 U15753 ( .B1(n13611), .B2(keyinput25), .C1(n13610), .C2(keyinput92), .A(n13609), .ZN(n13614) );
  INV_X1 U15754 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14822) );
  INV_X1 U15755 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n15072) );
  AOI22_X1 U15756 ( .A1(n14822), .A2(keyinput1), .B1(n15072), .B2(keyinput100), 
        .ZN(n13612) );
  OAI221_X1 U15757 ( .B1(n14822), .B2(keyinput1), .C1(n15072), .C2(keyinput100), .A(n13612), .ZN(n13613) );
  NOR4_X1 U15758 ( .A1(n13616), .A2(n13615), .A3(n13614), .A4(n13613), .ZN(
        n13645) );
  INV_X1 U15759 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n13618) );
  AOI22_X1 U15760 ( .A1(n13618), .A2(keyinput83), .B1(n13257), .B2(keyinput117), .ZN(n13617) );
  OAI221_X1 U15761 ( .B1(n13618), .B2(keyinput83), .C1(n13257), .C2(
        keyinput117), .A(n13617), .ZN(n13628) );
  AOI22_X1 U15762 ( .A1(n14375), .A2(keyinput17), .B1(n13620), .B2(keyinput116), .ZN(n13619) );
  OAI221_X1 U15763 ( .B1(n14375), .B2(keyinput17), .C1(n13620), .C2(
        keyinput116), .A(n13619), .ZN(n13627) );
  AOI22_X1 U15764 ( .A1(n10343), .A2(keyinput118), .B1(keyinput52), .B2(n6852), 
        .ZN(n13621) );
  OAI221_X1 U15765 ( .B1(n10343), .B2(keyinput118), .C1(n6852), .C2(keyinput52), .A(n13621), .ZN(n13626) );
  AOI22_X1 U15766 ( .A1(n13624), .A2(keyinput29), .B1(n13623), .B2(keyinput8), 
        .ZN(n13622) );
  OAI221_X1 U15767 ( .B1(n13624), .B2(keyinput29), .C1(n13623), .C2(keyinput8), 
        .A(n13622), .ZN(n13625) );
  NOR4_X1 U15768 ( .A1(n13628), .A2(n13627), .A3(n13626), .A4(n13625), .ZN(
        n13644) );
  INV_X1 U15769 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n14755) );
  AOI22_X1 U15770 ( .A1(n14755), .A2(keyinput93), .B1(keyinput63), .B2(n13630), 
        .ZN(n13629) );
  OAI221_X1 U15771 ( .B1(n14755), .B2(keyinput93), .C1(n13630), .C2(keyinput63), .A(n13629), .ZN(n13642) );
  AOI22_X1 U15772 ( .A1(n13633), .A2(keyinput66), .B1(n13632), .B2(keyinput20), 
        .ZN(n13631) );
  OAI221_X1 U15773 ( .B1(n13633), .B2(keyinput66), .C1(n13632), .C2(keyinput20), .A(n13631), .ZN(n13641) );
  INV_X1 U15774 ( .A(keyinput46), .ZN(n13635) );
  AOI22_X1 U15775 ( .A1(n11006), .A2(keyinput53), .B1(P3_DATAO_REG_24__SCAN_IN), .B2(n13635), .ZN(n13634) );
  OAI221_X1 U15776 ( .B1(n11006), .B2(keyinput53), .C1(n13635), .C2(
        P3_DATAO_REG_24__SCAN_IN), .A(n13634), .ZN(n13640) );
  AOI22_X1 U15777 ( .A1(n13638), .A2(keyinput16), .B1(keyinput44), .B2(n13637), 
        .ZN(n13636) );
  OAI221_X1 U15778 ( .B1(n13638), .B2(keyinput16), .C1(n13637), .C2(keyinput44), .A(n13636), .ZN(n13639) );
  NOR4_X1 U15779 ( .A1(n13642), .A2(n13641), .A3(n13640), .A4(n13639), .ZN(
        n13643) );
  NAND4_X1 U15780 ( .A1(n13646), .A2(n13645), .A3(n13644), .A4(n13643), .ZN(
        n13764) );
  AOI22_X1 U15781 ( .A1(n13649), .A2(keyinput113), .B1(keyinput82), .B2(n13648), .ZN(n13647) );
  OAI221_X1 U15782 ( .B1(n13649), .B2(keyinput113), .C1(n13648), .C2(
        keyinput82), .A(n13647), .ZN(n13660) );
  INV_X1 U15783 ( .A(SI_29_), .ZN(n13652) );
  AOI22_X1 U15784 ( .A1(n13652), .A2(keyinput12), .B1(keyinput77), .B2(n13651), 
        .ZN(n13650) );
  OAI221_X1 U15785 ( .B1(n13652), .B2(keyinput12), .C1(n13651), .C2(keyinput77), .A(n13650), .ZN(n13659) );
  XOR2_X1 U15786 ( .A(n13653), .B(keyinput41), .Z(n13657) );
  XNOR2_X1 U15787 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput7), .ZN(n13656) );
  XNOR2_X1 U15788 ( .A(P1_REG1_REG_31__SCAN_IN), .B(keyinput49), .ZN(n13655)
         );
  XNOR2_X1 U15789 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput6), .ZN(n13654) );
  NAND4_X1 U15790 ( .A1(n13657), .A2(n13656), .A3(n13655), .A4(n13654), .ZN(
        n13658) );
  NOR3_X1 U15791 ( .A1(n13660), .A2(n13659), .A3(n13658), .ZN(n13702) );
  INV_X1 U15792 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14809) );
  AOI22_X1 U15793 ( .A1(n7648), .A2(keyinput65), .B1(keyinput39), .B2(n14809), 
        .ZN(n13661) );
  OAI221_X1 U15794 ( .B1(n7648), .B2(keyinput65), .C1(n14809), .C2(keyinput39), 
        .A(n13661), .ZN(n13668) );
  AOI22_X1 U15795 ( .A1(n13664), .A2(keyinput121), .B1(n13663), .B2(keyinput57), .ZN(n13662) );
  OAI221_X1 U15796 ( .B1(n13664), .B2(keyinput121), .C1(n13663), .C2(
        keyinput57), .A(n13662), .ZN(n13667) );
  XNOR2_X1 U15797 ( .A(n13665), .B(keyinput43), .ZN(n13666) );
  OR3_X1 U15798 ( .A1(n13668), .A2(n13667), .A3(n13666), .ZN(n13675) );
  AOI22_X1 U15799 ( .A1(n13671), .A2(keyinput13), .B1(keyinput22), .B2(n13670), 
        .ZN(n13669) );
  OAI221_X1 U15800 ( .B1(n13671), .B2(keyinput13), .C1(n13670), .C2(keyinput22), .A(n13669), .ZN(n13674) );
  XNOR2_X1 U15801 ( .A(n13672), .B(P3_DATAO_REG_16__SCAN_IN), .ZN(n13673) );
  NOR3_X1 U15802 ( .A1(n13675), .A2(n13674), .A3(n13673), .ZN(n13701) );
  AOI22_X1 U15803 ( .A1(n7723), .A2(keyinput59), .B1(keyinput90), .B2(n9450), 
        .ZN(n13676) );
  OAI221_X1 U15804 ( .B1(n7723), .B2(keyinput59), .C1(n9450), .C2(keyinput90), 
        .A(n13676), .ZN(n13686) );
  AOI22_X1 U15805 ( .A1(n13678), .A2(keyinput33), .B1(n10458), .B2(keyinput94), 
        .ZN(n13677) );
  OAI221_X1 U15806 ( .B1(n13678), .B2(keyinput33), .C1(n10458), .C2(keyinput94), .A(n13677), .ZN(n13685) );
  INV_X1 U15807 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n13679) );
  XOR2_X1 U15808 ( .A(n13679), .B(keyinput35), .Z(n13683) );
  XOR2_X1 U15809 ( .A(n8712), .B(keyinput72), .Z(n13682) );
  XNOR2_X1 U15810 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput27), .ZN(n13681) );
  XNOR2_X1 U15811 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput122), .ZN(n13680) );
  NAND4_X1 U15812 ( .A1(n13683), .A2(n13682), .A3(n13681), .A4(n13680), .ZN(
        n13684) );
  NOR3_X1 U15813 ( .A1(n13686), .A2(n13685), .A3(n13684), .ZN(n13700) );
  AOI22_X1 U15814 ( .A1(n13688), .A2(keyinput23), .B1(n7575), .B2(keyinput126), 
        .ZN(n13687) );
  OAI221_X1 U15815 ( .B1(n13688), .B2(keyinput23), .C1(n7575), .C2(keyinput126), .A(n13687), .ZN(n13698) );
  INV_X1 U15816 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n15069) );
  AOI22_X1 U15817 ( .A1(n15069), .A2(keyinput21), .B1(keyinput70), .B2(n13690), 
        .ZN(n13689) );
  OAI221_X1 U15818 ( .B1(n15069), .B2(keyinput21), .C1(n13690), .C2(keyinput70), .A(n13689), .ZN(n13697) );
  XOR2_X1 U15819 ( .A(n10341), .B(keyinput87), .Z(n13695) );
  XOR2_X1 U15820 ( .A(n13691), .B(keyinput99), .Z(n13694) );
  XNOR2_X1 U15821 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput61), .ZN(n13693) );
  XNOR2_X1 U15822 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput28), .ZN(n13692)
         );
  NAND4_X1 U15823 ( .A1(n13695), .A2(n13694), .A3(n13693), .A4(n13692), .ZN(
        n13696) );
  NOR3_X1 U15824 ( .A1(n13698), .A2(n13697), .A3(n13696), .ZN(n13699) );
  NAND4_X1 U15825 ( .A1(n13702), .A2(n13701), .A3(n13700), .A4(n13699), .ZN(
        n13763) );
  INV_X1 U15826 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n14756) );
  AOI22_X1 U15827 ( .A1(n14756), .A2(keyinput14), .B1(keyinput125), .B2(n13704), .ZN(n13703) );
  OAI221_X1 U15828 ( .B1(n14756), .B2(keyinput14), .C1(n13704), .C2(
        keyinput125), .A(n13703), .ZN(n13715) );
  AOI22_X1 U15829 ( .A1(n13707), .A2(keyinput0), .B1(keyinput24), .B2(n13706), 
        .ZN(n13705) );
  OAI221_X1 U15830 ( .B1(n13707), .B2(keyinput0), .C1(n13706), .C2(keyinput24), 
        .A(n13705), .ZN(n13714) );
  AOI22_X1 U15831 ( .A1(n13944), .A2(keyinput84), .B1(n13709), .B2(keyinput88), 
        .ZN(n13708) );
  OAI221_X1 U15832 ( .B1(n13944), .B2(keyinput84), .C1(n13709), .C2(keyinput88), .A(n13708), .ZN(n13713) );
  XNOR2_X1 U15833 ( .A(P3_IR_REG_27__SCAN_IN), .B(keyinput48), .ZN(n13711) );
  XNOR2_X1 U15834 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput120), .ZN(n13710) );
  NAND2_X1 U15835 ( .A1(n13711), .A2(n13710), .ZN(n13712) );
  NOR4_X1 U15836 ( .A1(n13715), .A2(n13714), .A3(n13713), .A4(n13712), .ZN(
        n13761) );
  XNOR2_X1 U15837 ( .A(n13716), .B(keyinput109), .ZN(n13718) );
  XNOR2_X1 U15838 ( .A(keyinput79), .B(n9300), .ZN(n13717) );
  NOR2_X1 U15839 ( .A1(n13718), .A2(n13717), .ZN(n13720) );
  XNOR2_X1 U15840 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput78), .ZN(n13719) );
  OAI211_X1 U15841 ( .C1(n14984), .C2(keyinput127), .A(n13720), .B(n13719), 
        .ZN(n13727) );
  INV_X1 U15842 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15068) );
  AOI22_X1 U15843 ( .A1(n15015), .A2(keyinput36), .B1(n15068), .B2(keyinput91), 
        .ZN(n13721) );
  OAI221_X1 U15844 ( .B1(n15015), .B2(keyinput36), .C1(n15068), .C2(keyinput91), .A(n13721), .ZN(n13726) );
  INV_X1 U15845 ( .A(P1_RD_REG_SCAN_IN), .ZN(n13724) );
  AOI22_X1 U15846 ( .A1(n7444), .A2(keyinput98), .B1(keyinput47), .B2(n13723), 
        .ZN(n13722) );
  OAI221_X1 U15847 ( .B1(n7444), .B2(keyinput98), .C1(n13723), .C2(keyinput47), 
        .A(n13722), .ZN(n13725) );
  NOR3_X1 U15848 ( .A1(n13727), .A2(n13726), .A3(n13725), .ZN(n13760) );
  INV_X1 U15849 ( .A(keyinput2), .ZN(n13729) );
  AOI22_X1 U15850 ( .A1(n13730), .A2(keyinput51), .B1(P3_DATAO_REG_29__SCAN_IN), .B2(n13729), .ZN(n13728) );
  OAI221_X1 U15851 ( .B1(n13730), .B2(keyinput51), .C1(n13729), .C2(
        P3_DATAO_REG_29__SCAN_IN), .A(n13728), .ZN(n13743) );
  INV_X1 U15852 ( .A(keyinput86), .ZN(n13733) );
  INV_X1 U15853 ( .A(keyinput18), .ZN(n13732) );
  AOI22_X1 U15854 ( .A1(n13733), .A2(P3_DATAO_REG_9__SCAN_IN), .B1(
        P3_DATAO_REG_15__SCAN_IN), .B2(n13732), .ZN(n13731) );
  OAI221_X1 U15855 ( .B1(n13733), .B2(P3_DATAO_REG_9__SCAN_IN), .C1(n13732), 
        .C2(P3_DATAO_REG_15__SCAN_IN), .A(n13731), .ZN(n13742) );
  INV_X1 U15856 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13736) );
  AOI22_X1 U15857 ( .A1(n13736), .A2(keyinput55), .B1(n13735), .B2(keyinput38), 
        .ZN(n13734) );
  OAI221_X1 U15858 ( .B1(n13736), .B2(keyinput55), .C1(n13735), .C2(keyinput38), .A(n13734), .ZN(n13741) );
  INV_X1 U15859 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n13737) );
  XOR2_X1 U15860 ( .A(n13737), .B(keyinput19), .Z(n13739) );
  XNOR2_X1 U15861 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput9), .ZN(n13738) );
  NAND2_X1 U15862 ( .A1(n13739), .A2(n13738), .ZN(n13740) );
  NOR4_X1 U15863 ( .A1(n13743), .A2(n13742), .A3(n13741), .A4(n13740), .ZN(
        n13759) );
  INV_X1 U15864 ( .A(keyinput10), .ZN(n13745) );
  AOI22_X1 U15865 ( .A1(n13746), .A2(keyinput60), .B1(P3_WR_REG_SCAN_IN), .B2(
        n13745), .ZN(n13744) );
  OAI221_X1 U15866 ( .B1(n13746), .B2(keyinput60), .C1(n13745), .C2(
        P3_WR_REG_SCAN_IN), .A(n13744), .ZN(n13757) );
  AOI22_X1 U15867 ( .A1(n13749), .A2(keyinput40), .B1(n13748), .B2(keyinput95), 
        .ZN(n13747) );
  OAI221_X1 U15868 ( .B1(n13749), .B2(keyinput40), .C1(n13748), .C2(keyinput95), .A(n13747), .ZN(n13756) );
  INV_X1 U15869 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13751) );
  AOI22_X1 U15870 ( .A1(n13751), .A2(keyinput81), .B1(n10669), .B2(keyinput107), .ZN(n13750) );
  OAI221_X1 U15871 ( .B1(n13751), .B2(keyinput81), .C1(n10669), .C2(
        keyinput107), .A(n13750), .ZN(n13755) );
  INV_X1 U15872 ( .A(keyinput110), .ZN(n13753) );
  AOI22_X1 U15873 ( .A1(n9361), .A2(keyinput68), .B1(P3_DATAO_REG_30__SCAN_IN), 
        .B2(n13753), .ZN(n13752) );
  OAI221_X1 U15874 ( .B1(n9361), .B2(keyinput68), .C1(n13753), .C2(
        P3_DATAO_REG_30__SCAN_IN), .A(n13752), .ZN(n13754) );
  NOR4_X1 U15875 ( .A1(n13757), .A2(n13756), .A3(n13755), .A4(n13754), .ZN(
        n13758) );
  NAND4_X1 U15876 ( .A1(n13761), .A2(n13760), .A3(n13759), .A4(n13758), .ZN(
        n13762) );
  NOR4_X1 U15877 ( .A1(n13765), .A2(n13764), .A3(n13763), .A4(n13762), .ZN(
        n13766) );
  OAI21_X1 U15878 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n13767), .A(n13766), 
        .ZN(n13771) );
  AOI222_X1 U15879 ( .A1(n14297), .A2(n6726), .B1(P1_DATAO_REG_26__SCAN_IN), 
        .B2(n13769), .C1(n13768), .C2(P2_STATE_REG_SCAN_IN), .ZN(n13770) );
  XOR2_X1 U15880 ( .A(n13771), .B(n13770), .Z(P2_U3301) );
  INV_X1 U15881 ( .A(n13772), .ZN(n14303) );
  INV_X1 U15882 ( .A(n13773), .ZN(n13774) );
  OAI222_X1 U15883 ( .A1(n13776), .A2(n13775), .B1(n11134), .B2(n14303), .C1(
        P2_U3088), .C2(n13774), .ZN(P2_U3302) );
  MUX2_X1 U15884 ( .A(n13778), .B(n13777), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3327) );
  XOR2_X1 U15885 ( .A(n13780), .B(n13779), .Z(n13785) );
  AOI22_X1 U15886 ( .A1(n14545), .A2(n14012), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13782) );
  NAND2_X1 U15887 ( .A1(n14547), .A2(n14011), .ZN(n13781) );
  OAI211_X1 U15888 ( .C1(n14554), .C2(n14015), .A(n13782), .B(n13781), .ZN(
        n13783) );
  AOI21_X1 U15889 ( .B1(n14020), .B2(n14536), .A(n13783), .ZN(n13784) );
  OAI21_X1 U15890 ( .B1(n13785), .B2(n14532), .A(n13784), .ZN(P1_U3214) );
  XOR2_X1 U15891 ( .A(n13787), .B(n13786), .Z(n13794) );
  OR2_X1 U15892 ( .A1(n13788), .A2(n14555), .ZN(n13790) );
  NAND2_X1 U15893 ( .A1(n13888), .A2(n14177), .ZN(n13789) );
  NAND2_X1 U15894 ( .A1(n13790), .A2(n13789), .ZN(n14234) );
  AOI22_X1 U15895 ( .A1(n14517), .A2(n14234), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13791) );
  OAI21_X1 U15896 ( .B1(n14081), .B2(n14554), .A(n13791), .ZN(n13792) );
  AOI21_X1 U15897 ( .B1(n14235), .B2(n14536), .A(n13792), .ZN(n13793) );
  OAI21_X1 U15898 ( .B1(n13794), .B2(n14532), .A(n13793), .ZN(P1_U3216) );
  INV_X1 U15899 ( .A(n14260), .ZN(n14141) );
  AOI21_X1 U15900 ( .B1(n13796), .B2(n13795), .A(n14532), .ZN(n13798) );
  NAND2_X1 U15901 ( .A1(n13798), .A2(n13797), .ZN(n13804) );
  OR2_X1 U15902 ( .A1(n13799), .A2(n14557), .ZN(n13801) );
  NAND2_X1 U15903 ( .A1(n14159), .A2(n14178), .ZN(n13800) );
  NAND2_X1 U15904 ( .A1(n13801), .A2(n13800), .ZN(n14259) );
  AND2_X1 U15905 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13987) );
  NOR2_X1 U15906 ( .A1(n14554), .A2(n14137), .ZN(n13802) );
  AOI211_X1 U15907 ( .C1(n14259), .C2(n14517), .A(n13987), .B(n13802), .ZN(
        n13803) );
  OAI211_X1 U15908 ( .C1(n14141), .C2(n14549), .A(n13804), .B(n13803), .ZN(
        P1_U3219) );
  INV_X1 U15909 ( .A(n13805), .ZN(n13806) );
  AOI21_X1 U15910 ( .B1(n13808), .B2(n13807), .A(n13806), .ZN(n13813) );
  AOI22_X1 U15911 ( .A1(n14547), .A2(n14106), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13810) );
  NAND2_X1 U15912 ( .A1(n14107), .A2(n14545), .ZN(n13809) );
  OAI211_X1 U15913 ( .C1(n14554), .C2(n14109), .A(n13810), .B(n13809), .ZN(
        n13811) );
  AOI21_X1 U15914 ( .B1(n14246), .B2(n14536), .A(n13811), .ZN(n13812) );
  OAI21_X1 U15915 ( .B1(n13813), .B2(n14532), .A(n13812), .ZN(P1_U3223) );
  XOR2_X1 U15916 ( .A(n13815), .B(n13814), .Z(n13821) );
  NAND2_X1 U15917 ( .A1(n13888), .A2(n14178), .ZN(n13817) );
  NAND2_X1 U15918 ( .A1(n14012), .A2(n14177), .ZN(n13816) );
  NAND2_X1 U15919 ( .A1(n13817), .A2(n13816), .ZN(n14220) );
  AOI22_X1 U15920 ( .A1(n14517), .A2(n14220), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13818) );
  OAI21_X1 U15921 ( .B1(n14045), .B2(n14554), .A(n13818), .ZN(n13819) );
  AOI21_X1 U15922 ( .B1(n14221), .B2(n14536), .A(n13819), .ZN(n13820) );
  OAI21_X1 U15923 ( .B1(n13821), .B2(n14532), .A(n13820), .ZN(P1_U3225) );
  XOR2_X1 U15924 ( .A(n13823), .B(n13822), .Z(n13828) );
  AOI22_X1 U15925 ( .A1(n14545), .A2(n14059), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13825) );
  NAND2_X1 U15926 ( .A1(n14547), .A2(n14058), .ZN(n13824) );
  OAI211_X1 U15927 ( .C1(n14554), .C2(n14063), .A(n13825), .B(n13824), .ZN(
        n13826) );
  AOI21_X1 U15928 ( .B1(n14068), .B2(n14536), .A(n13826), .ZN(n13827) );
  OAI21_X1 U15929 ( .B1(n13828), .B2(n14532), .A(n13827), .ZN(P1_U3229) );
  OAI211_X1 U15930 ( .C1(n13831), .C2(n13830), .A(n13829), .B(n14551), .ZN(
        n13839) );
  INV_X1 U15931 ( .A(n13832), .ZN(n14122) );
  AND2_X1 U15932 ( .A1(n13889), .A2(n14177), .ZN(n13833) );
  AOI21_X1 U15933 ( .B1(n14146), .B2(n14178), .A(n13833), .ZN(n14250) );
  OAI22_X1 U15934 ( .A1(n14250), .A2(n13835), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13834), .ZN(n13836) );
  AOI21_X1 U15935 ( .B1(n14122), .B2(n13837), .A(n13836), .ZN(n13838) );
  OAI211_X1 U15936 ( .C1(n14252), .C2(n14549), .A(n13839), .B(n13838), .ZN(
        P1_U3233) );
  OAI211_X1 U15937 ( .C1(n13842), .C2(n13841), .A(n13840), .B(n14551), .ZN(
        n13849) );
  AOI22_X1 U15938 ( .A1(n14517), .A2(n13843), .B1(P1_REG3_REG_13__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13844) );
  OAI21_X1 U15939 ( .B1(n13845), .B2(n14554), .A(n13844), .ZN(n13846) );
  AOI21_X1 U15940 ( .B1(n13847), .B2(n14536), .A(n13846), .ZN(n13848) );
  NAND2_X1 U15941 ( .A1(n13849), .A2(n13848), .ZN(P1_U3234) );
  OAI21_X1 U15942 ( .B1(n13852), .B2(n13851), .A(n13850), .ZN(n13858) );
  NOR2_X1 U15943 ( .A1(n14101), .A2(n14549), .ZN(n13857) );
  NAND2_X1 U15944 ( .A1(n13889), .A2(n14178), .ZN(n13854) );
  NAND2_X1 U15945 ( .A1(n14059), .A2(n14177), .ZN(n13853) );
  NAND2_X1 U15946 ( .A1(n13854), .A2(n13853), .ZN(n14240) );
  AOI22_X1 U15947 ( .A1(n14517), .A2(n14240), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13855) );
  OAI21_X1 U15948 ( .B1(n14096), .B2(n14554), .A(n13855), .ZN(n13856) );
  AOI211_X1 U15949 ( .C1(n13858), .C2(n14551), .A(n13857), .B(n13856), .ZN(
        n13859) );
  INV_X1 U15950 ( .A(n13859), .ZN(P1_U3235) );
  XOR2_X1 U15951 ( .A(n13860), .B(n13861), .Z(n13867) );
  NOR2_X1 U15952 ( .A1(n14554), .A2(n14149), .ZN(n13865) );
  NAND2_X1 U15953 ( .A1(n14545), .A2(n14508), .ZN(n13862) );
  NAND2_X1 U15954 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13954)
         );
  OAI211_X1 U15955 ( .C1(n14526), .C2(n13863), .A(n13862), .B(n13954), .ZN(
        n13864) );
  AOI211_X1 U15956 ( .C1(n14265), .C2(n14536), .A(n13865), .B(n13864), .ZN(
        n13866) );
  OAI21_X1 U15957 ( .B1(n13867), .B2(n14532), .A(n13866), .ZN(P1_U3238) );
  OAI211_X1 U15958 ( .C1(n13870), .C2(n13869), .A(n13868), .B(n14551), .ZN(
        n13877) );
  NOR2_X1 U15959 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8397), .ZN(n13923) );
  AOI21_X1 U15960 ( .B1(n14517), .B2(n13871), .A(n13923), .ZN(n13876) );
  NAND2_X1 U15961 ( .A1(n14536), .A2(n13872), .ZN(n13875) );
  OR2_X1 U15962 ( .A1(n14554), .A2(n13873), .ZN(n13874) );
  NAND4_X1 U15963 ( .A1(n13877), .A2(n13876), .A3(n13875), .A4(n13874), .ZN(
        P1_U3239) );
  XOR2_X1 U15964 ( .A(n13879), .B(n13878), .Z(n13884) );
  OAI22_X1 U15965 ( .A1(n13880), .A2(n14555), .B1(n11906), .B2(n14557), .ZN(
        n14028) );
  AOI22_X1 U15966 ( .A1(n14028), .A2(n14517), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13881) );
  OAI21_X1 U15967 ( .B1(n14031), .B2(n14554), .A(n13881), .ZN(n13882) );
  AOI21_X1 U15968 ( .B1(n14214), .B2(n14536), .A(n13882), .ZN(n13883) );
  OAI21_X1 U15969 ( .B1(n13884), .B2(n14532), .A(n13883), .ZN(P1_U3240) );
  MUX2_X1 U15970 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13994), .S(n14655), .Z(
        P1_U3591) );
  MUX2_X1 U15971 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13885), .S(n14655), .Z(
        P1_U3590) );
  MUX2_X1 U15972 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13886), .S(n14655), .Z(
        P1_U3589) );
  MUX2_X1 U15973 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14011), .S(n14655), .Z(
        P1_U3588) );
  MUX2_X1 U15974 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13887), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15975 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14012), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15976 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14058), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15977 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13888), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15978 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14059), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15979 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14106), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15980 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13889), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15981 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14107), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15982 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14146), .S(n14655), .Z(
        P1_U3579) );
  MUX2_X1 U15983 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14159), .S(n14655), .Z(
        P1_U3578) );
  MUX2_X1 U15984 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14508), .S(n14655), .Z(
        P1_U3577) );
  MUX2_X1 U15985 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14546), .S(n14655), .Z(
        P1_U3576) );
  MUX2_X1 U15986 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14507), .S(n14655), .Z(
        P1_U3575) );
  MUX2_X1 U15987 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14544), .S(n14655), .Z(
        P1_U3574) );
  MUX2_X1 U15988 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13890), .S(n14655), .Z(
        P1_U3572) );
  MUX2_X1 U15989 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13891), .S(n14655), .Z(
        P1_U3571) );
  MUX2_X1 U15990 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13892), .S(n14655), .Z(
        P1_U3570) );
  MUX2_X1 U15991 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13893), .S(n14655), .Z(
        P1_U3567) );
  MUX2_X1 U15992 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13894), .S(n14655), .Z(
        P1_U3566) );
  MUX2_X1 U15993 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13895), .S(n14655), .Z(
        P1_U3565) );
  MUX2_X1 U15994 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13896), .S(n14655), .Z(
        P1_U3564) );
  MUX2_X1 U15995 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13897), .S(n14655), .Z(
        P1_U3563) );
  MUX2_X1 U15996 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13898), .S(n14655), .Z(
        P1_U3562) );
  NOR2_X1 U15997 ( .A1(n13900), .A2(n13899), .ZN(n14652) );
  OAI211_X1 U15998 ( .C1(n14652), .C2(n13901), .A(n14669), .B(n14637), .ZN(
        n13908) );
  OAI211_X1 U15999 ( .C1(n13903), .C2(n13902), .A(n14684), .B(n14642), .ZN(
        n13907) );
  AOI22_X1 U16000 ( .A1(n14675), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13906) );
  NAND2_X1 U16001 ( .A1(n14687), .A2(n13904), .ZN(n13905) );
  NAND4_X1 U16002 ( .A1(n13908), .A2(n13907), .A3(n13906), .A4(n13905), .ZN(
        P1_U3244) );
  OAI211_X1 U16003 ( .C1(n13911), .C2(n13910), .A(n14684), .B(n13909), .ZN(
        n13920) );
  OR3_X1 U16004 ( .A1(n13913), .A2(n14640), .A3(n13912), .ZN(n13914) );
  NAND3_X1 U16005 ( .A1(n14669), .A2(n14666), .A3(n13914), .ZN(n13919) );
  NAND2_X1 U16006 ( .A1(n14687), .A2(n13915), .ZN(n13918) );
  NOR2_X1 U16007 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10768), .ZN(n13916) );
  AOI21_X1 U16008 ( .B1(n14675), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n13916), .ZN(
        n13917) );
  NAND4_X1 U16009 ( .A1(n13920), .A2(n13919), .A3(n13918), .A4(n13917), .ZN(
        P1_U3246) );
  NOR2_X1 U16010 ( .A1(n14673), .A2(n13921), .ZN(n13922) );
  AOI211_X1 U16011 ( .C1(n14675), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n13923), .B(
        n13922), .ZN(n13935) );
  OAI211_X1 U16012 ( .C1(n13926), .C2(n13925), .A(n14684), .B(n13924), .ZN(
        n13934) );
  INV_X1 U16013 ( .A(n13927), .ZN(n13932) );
  NAND3_X1 U16014 ( .A1(n13930), .A2(n13929), .A3(n13928), .ZN(n13931) );
  NAND3_X1 U16015 ( .A1(n14669), .A2(n13932), .A3(n13931), .ZN(n13933) );
  NAND3_X1 U16016 ( .A1(n13935), .A2(n13934), .A3(n13933), .ZN(P1_U3249) );
  AOI21_X1 U16017 ( .B1(n13937), .B2(P1_REG1_REG_16__SCAN_IN), .A(n13936), 
        .ZN(n13942) );
  NOR2_X1 U16018 ( .A1(n13961), .A2(n13938), .ZN(n13939) );
  AOI21_X1 U16019 ( .B1(n13961), .B2(n13938), .A(n13939), .ZN(n13941) );
  NOR2_X1 U16020 ( .A1(n13942), .A2(n13941), .ZN(n13960) );
  AOI211_X1 U16021 ( .C1(n13942), .C2(n13941), .A(n13960), .B(n13940), .ZN(
        n13943) );
  INV_X1 U16022 ( .A(n13943), .ZN(n13953) );
  NOR2_X1 U16023 ( .A1(n13944), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14520) );
  NOR2_X1 U16024 ( .A1(n14673), .A2(n13957), .ZN(n13945) );
  AOI211_X1 U16025 ( .C1(n14675), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n14520), 
        .B(n13945), .ZN(n13952) );
  INV_X1 U16026 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13958) );
  NOR2_X1 U16027 ( .A1(n13957), .A2(n13958), .ZN(n13946) );
  AOI21_X1 U16028 ( .B1(n13958), .B2(n13957), .A(n13946), .ZN(n13950) );
  OAI21_X1 U16029 ( .B1(n13948), .B2(n11296), .A(n13947), .ZN(n13949) );
  NAND2_X1 U16030 ( .A1(n13950), .A2(n13949), .ZN(n13956) );
  OAI211_X1 U16031 ( .C1(n13950), .C2(n13949), .A(n14669), .B(n13956), .ZN(
        n13951) );
  NAND3_X1 U16032 ( .A1(n13953), .A2(n13952), .A3(n13951), .ZN(P1_U3260) );
  OAI21_X1 U16033 ( .B1(n14695), .B2(n13691), .A(n13954), .ZN(n13955) );
  AOI21_X1 U16034 ( .B1(n13976), .B2(n14687), .A(n13955), .ZN(n13968) );
  OAI21_X1 U16035 ( .B1(n13958), .B2(n13957), .A(n13956), .ZN(n13975) );
  XNOR2_X1 U16036 ( .A(n13969), .B(n13975), .ZN(n13959) );
  NAND2_X1 U16037 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n13959), .ZN(n13978) );
  OAI211_X1 U16038 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n13959), .A(n14669), 
        .B(n13978), .ZN(n13967) );
  AOI21_X1 U16039 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n13961), .A(n13960), 
        .ZN(n13970) );
  XNOR2_X1 U16040 ( .A(n13969), .B(n13970), .ZN(n13962) );
  INV_X1 U16041 ( .A(n13962), .ZN(n13965) );
  NOR2_X1 U16042 ( .A1(n13963), .A2(n13962), .ZN(n13972) );
  INV_X1 U16043 ( .A(n13972), .ZN(n13964) );
  OAI211_X1 U16044 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n13965), .A(n14684), 
        .B(n13964), .ZN(n13966) );
  NAND3_X1 U16045 ( .A1(n13968), .A2(n13967), .A3(n13966), .ZN(P1_U3261) );
  NOR2_X1 U16046 ( .A1(n13970), .A2(n13969), .ZN(n13971) );
  NOR2_X1 U16047 ( .A1(n13972), .A2(n13971), .ZN(n13974) );
  XOR2_X1 U16048 ( .A(n13974), .B(n13973), .Z(n13983) );
  INV_X1 U16049 ( .A(n13983), .ZN(n13981) );
  NAND2_X1 U16050 ( .A1(n13976), .A2(n13975), .ZN(n13977) );
  NAND2_X1 U16051 ( .A1(n13978), .A2(n13977), .ZN(n13979) );
  XOR2_X1 U16052 ( .A(n13979), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13982) );
  OAI21_X1 U16053 ( .B1(n13982), .B2(n14690), .A(n14673), .ZN(n13980) );
  AOI21_X1 U16054 ( .B1(n13981), .B2(n14684), .A(n13980), .ZN(n13986) );
  AOI22_X1 U16055 ( .A1(n13983), .A2(n14684), .B1(n14669), .B2(n13982), .ZN(
        n13985) );
  MUX2_X1 U16056 ( .A(n13986), .B(n13985), .S(n13984), .Z(n13989) );
  INV_X1 U16057 ( .A(n13987), .ZN(n13988) );
  OAI211_X1 U16058 ( .C1(n7445), .C2(n14695), .A(n13989), .B(n13988), .ZN(
        P1_U3262) );
  NAND2_X1 U16059 ( .A1(n14194), .A2(n13999), .ZN(n13990) );
  XNOR2_X1 U16060 ( .A(n14191), .B(n13990), .ZN(n13991) );
  NAND2_X1 U16061 ( .A1(n13991), .A2(n14725), .ZN(n14190) );
  NOR2_X1 U16062 ( .A1(n14741), .A2(n13992), .ZN(n13995) );
  NAND2_X1 U16063 ( .A1(n13994), .A2(n13993), .ZN(n14192) );
  NOR2_X1 U16064 ( .A1(n14157), .A2(n14192), .ZN(n14002) );
  AOI211_X1 U16065 ( .C1(n13996), .C2(n14743), .A(n13995), .B(n14002), .ZN(
        n13997) );
  OAI21_X1 U16066 ( .B1(n14190), .B2(n14186), .A(n13997), .ZN(P1_U3263) );
  XNOR2_X1 U16067 ( .A(n13999), .B(n13998), .ZN(n14000) );
  NAND2_X1 U16068 ( .A1(n14000), .A2(n14725), .ZN(n14193) );
  NOR2_X1 U16069 ( .A1(n14194), .A2(n14337), .ZN(n14001) );
  AOI211_X1 U16070 ( .C1(n14157), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14002), 
        .B(n14001), .ZN(n14003) );
  OAI21_X1 U16071 ( .B1(n14186), .B2(n14193), .A(n14003), .ZN(P1_U3264) );
  NAND2_X1 U16072 ( .A1(n14004), .A2(n14007), .ZN(n14005) );
  NOR2_X1 U16073 ( .A1(n14008), .A2(n14007), .ZN(n14009) );
  OAI21_X1 U16074 ( .B1(n14010), .B2(n14009), .A(n14738), .ZN(n14014) );
  AOI22_X1 U16075 ( .A1(n14178), .A2(n14012), .B1(n14011), .B2(n14177), .ZN(
        n14013) );
  OAI211_X1 U16076 ( .C1(n14207), .C2(n14734), .A(n14014), .B(n14013), .ZN(
        n14212) );
  NAND2_X1 U16077 ( .A1(n14212), .A2(n14741), .ZN(n14022) );
  INV_X1 U16078 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14016) );
  OAI22_X1 U16079 ( .A1(n14741), .A2(n14016), .B1(n14015), .B2(n14739), .ZN(
        n14019) );
  OAI211_X1 U16080 ( .C1(n11907), .C2(n14035), .A(n14725), .B(n14017), .ZN(
        n14209) );
  NOR2_X1 U16081 ( .A1(n14209), .A2(n14186), .ZN(n14018) );
  AOI211_X1 U16082 ( .C1(n14743), .C2(n14020), .A(n14019), .B(n14018), .ZN(
        n14021) );
  OAI211_X1 U16083 ( .C1(n14207), .C2(n14071), .A(n14022), .B(n14021), .ZN(
        P1_U3266) );
  XNOR2_X1 U16084 ( .A(n14024), .B(n14023), .ZN(n14217) );
  OAI21_X1 U16085 ( .B1(n14027), .B2(n14026), .A(n14025), .ZN(n14029) );
  AOI21_X1 U16086 ( .B1(n14029), .B2(n14738), .A(n14028), .ZN(n14216) );
  NAND2_X1 U16087 ( .A1(n14157), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n14030) );
  OAI21_X1 U16088 ( .B1(n14739), .B2(n14031), .A(n14030), .ZN(n14032) );
  AOI21_X1 U16089 ( .B1(n14214), .B2(n14743), .A(n14032), .ZN(n14037) );
  NAND2_X1 U16090 ( .A1(n14214), .A2(n14043), .ZN(n14033) );
  NAND2_X1 U16091 ( .A1(n14033), .A2(n14725), .ZN(n14034) );
  NOR2_X1 U16092 ( .A1(n14035), .A2(n14034), .ZN(n14213) );
  NAND2_X1 U16093 ( .A1(n14213), .A2(n6575), .ZN(n14036) );
  OAI211_X1 U16094 ( .C1(n14216), .C2(n14157), .A(n14037), .B(n14036), .ZN(
        n14038) );
  INV_X1 U16095 ( .A(n14038), .ZN(n14039) );
  OAI21_X1 U16096 ( .B1(n14339), .B2(n14217), .A(n14039), .ZN(P1_U3267) );
  OAI21_X1 U16097 ( .B1(n6689), .B2(n14041), .A(n14040), .ZN(n14224) );
  XNOR2_X1 U16098 ( .A(n14042), .B(n14041), .ZN(n14218) );
  NAND2_X1 U16099 ( .A1(n14218), .A2(n14571), .ZN(n14051) );
  AOI21_X1 U16100 ( .B1(n14221), .B2(n14065), .A(n14745), .ZN(n14044) );
  AND2_X1 U16101 ( .A1(n14044), .A2(n14043), .ZN(n14219) );
  INV_X1 U16102 ( .A(n14220), .ZN(n14046) );
  OAI22_X1 U16103 ( .A1(n14157), .A2(n14046), .B1(n14045), .B2(n14739), .ZN(
        n14047) );
  AOI21_X1 U16104 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(n14157), .A(n14047), 
        .ZN(n14048) );
  OAI21_X1 U16105 ( .B1(n7000), .B2(n14337), .A(n14048), .ZN(n14049) );
  AOI21_X1 U16106 ( .B1(n14219), .B2(n6575), .A(n14049), .ZN(n14050) );
  OAI211_X1 U16107 ( .C1(n14224), .C2(n14339), .A(n14051), .B(n14050), .ZN(
        P1_U3268) );
  OAI21_X1 U16108 ( .B1(n14053), .B2(n14054), .A(n14052), .ZN(n14225) );
  INV_X1 U16109 ( .A(n14225), .ZN(n14072) );
  NAND2_X1 U16110 ( .A1(n14055), .A2(n14054), .ZN(n14056) );
  NAND3_X1 U16111 ( .A1(n14057), .A2(n14738), .A3(n14056), .ZN(n14062) );
  AOI22_X1 U16112 ( .A1(n14178), .A2(n14059), .B1(n14058), .B2(n14177), .ZN(
        n14061) );
  NAND2_X1 U16113 ( .A1(n14225), .A2(n14719), .ZN(n14060) );
  NAND3_X1 U16114 ( .A1(n14062), .A2(n14061), .A3(n14060), .ZN(n14230) );
  NAND2_X1 U16115 ( .A1(n14230), .A2(n14741), .ZN(n14070) );
  OAI22_X1 U16116 ( .A1(n14741), .A2(n14064), .B1(n14063), .B2(n14739), .ZN(
        n14067) );
  OAI211_X1 U16117 ( .C1(n14228), .C2(n6610), .A(n14725), .B(n14065), .ZN(
        n14226) );
  NOR2_X1 U16118 ( .A1(n14226), .A2(n14186), .ZN(n14066) );
  AOI211_X1 U16119 ( .C1(n14743), .C2(n14068), .A(n14067), .B(n14066), .ZN(
        n14069) );
  OAI211_X1 U16120 ( .C1(n14072), .C2(n14071), .A(n14070), .B(n14069), .ZN(
        P1_U3269) );
  NAND2_X1 U16121 ( .A1(n14073), .A2(n14077), .ZN(n14074) );
  NAND2_X1 U16122 ( .A1(n14075), .A2(n14074), .ZN(n14238) );
  OAI21_X1 U16123 ( .B1(n14078), .B2(n14077), .A(n14076), .ZN(n14079) );
  NAND2_X1 U16124 ( .A1(n14079), .A2(n14738), .ZN(n14237) );
  INV_X1 U16125 ( .A(n14234), .ZN(n14080) );
  OAI211_X1 U16126 ( .C1(n14739), .C2(n14081), .A(n14237), .B(n14080), .ZN(
        n14082) );
  NAND2_X1 U16127 ( .A1(n14082), .A2(n14741), .ZN(n14087) );
  AOI211_X1 U16128 ( .C1(n14235), .C2(n14093), .A(n14745), .B(n6610), .ZN(
        n14233) );
  INV_X1 U16129 ( .A(n14235), .ZN(n14084) );
  INV_X1 U16130 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14083) );
  OAI22_X1 U16131 ( .A1(n14084), .A2(n14337), .B1(n14083), .B2(n14741), .ZN(
        n14085) );
  AOI21_X1 U16132 ( .B1(n14233), .B2(n6575), .A(n14085), .ZN(n14086) );
  OAI211_X1 U16133 ( .C1(n14238), .C2(n14339), .A(n14087), .B(n14086), .ZN(
        P1_U3270) );
  XNOR2_X1 U16134 ( .A(n14089), .B(n14088), .ZN(n14244) );
  OAI21_X1 U16135 ( .B1(n14092), .B2(n14091), .A(n14090), .ZN(n14241) );
  INV_X1 U16136 ( .A(n14093), .ZN(n14094) );
  AOI211_X1 U16137 ( .C1(n7004), .C2(n14095), .A(n14745), .B(n14094), .ZN(
        n14239) );
  NAND2_X1 U16138 ( .A1(n14239), .A2(n6575), .ZN(n14100) );
  INV_X1 U16139 ( .A(n14240), .ZN(n14097) );
  OAI22_X1 U16140 ( .A1(n14157), .A2(n14097), .B1(n14096), .B2(n14739), .ZN(
        n14098) );
  AOI21_X1 U16141 ( .B1(P1_REG2_REG_22__SCAN_IN), .B2(n14157), .A(n14098), 
        .ZN(n14099) );
  OAI211_X1 U16142 ( .C1(n14337), .C2(n14101), .A(n14100), .B(n14099), .ZN(
        n14102) );
  AOI21_X1 U16143 ( .B1(n14570), .B2(n14241), .A(n14102), .ZN(n14103) );
  OAI21_X1 U16144 ( .B1(n14244), .B2(n14189), .A(n14103), .ZN(P1_U3271) );
  XNOR2_X1 U16145 ( .A(n14104), .B(n14113), .ZN(n14105) );
  AOI222_X1 U16146 ( .A1(n14107), .A2(n14178), .B1(n14106), .B2(n14177), .C1(
        n14738), .C2(n14105), .ZN(n14248) );
  AOI211_X1 U16147 ( .C1(n14246), .C2(n14121), .A(n14745), .B(n14108), .ZN(
        n14245) );
  INV_X1 U16148 ( .A(n14246), .ZN(n14112) );
  INV_X1 U16149 ( .A(n14109), .ZN(n14110) );
  AOI22_X1 U16150 ( .A1(n14157), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14110), 
        .B2(n14722), .ZN(n14111) );
  OAI21_X1 U16151 ( .B1(n14112), .B2(n14337), .A(n14111), .ZN(n14116) );
  XNOR2_X1 U16152 ( .A(n14114), .B(n14113), .ZN(n14249) );
  NOR2_X1 U16153 ( .A1(n14249), .A2(n14339), .ZN(n14115) );
  AOI211_X1 U16154 ( .C1(n14245), .C2(n6575), .A(n14116), .B(n14115), .ZN(
        n14117) );
  OAI21_X1 U16155 ( .B1(n14248), .B2(n14157), .A(n14117), .ZN(P1_U3272) );
  XNOR2_X1 U16156 ( .A(n14119), .B(n14118), .ZN(n14256) );
  AOI21_X1 U16157 ( .B1(n7305), .B2(n14120), .A(n6712), .ZN(n14254) );
  OAI211_X1 U16158 ( .C1(n14252), .C2(n14135), .A(n14725), .B(n14121), .ZN(
        n14251) );
  AOI22_X1 U16159 ( .A1(n14157), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14122), 
        .B2(n14722), .ZN(n14123) );
  OAI21_X1 U16160 ( .B1(n14250), .B2(n14157), .A(n14123), .ZN(n14124) );
  AOI21_X1 U16161 ( .B1(n14125), .B2(n14743), .A(n14124), .ZN(n14126) );
  OAI21_X1 U16162 ( .B1(n14251), .B2(n14186), .A(n14126), .ZN(n14127) );
  AOI21_X1 U16163 ( .B1(n14254), .B2(n14570), .A(n14127), .ZN(n14128) );
  OAI21_X1 U16164 ( .B1(n14256), .B2(n14189), .A(n14128), .ZN(P1_U3273) );
  XNOR2_X1 U16165 ( .A(n14130), .B(n14129), .ZN(n14263) );
  OAI21_X1 U16166 ( .B1(n6709), .B2(n14132), .A(n14131), .ZN(n14257) );
  NAND2_X1 U16167 ( .A1(n14260), .A2(n14147), .ZN(n14133) );
  NAND2_X1 U16168 ( .A1(n14133), .A2(n14725), .ZN(n14134) );
  NOR2_X1 U16169 ( .A1(n14135), .A2(n14134), .ZN(n14258) );
  NAND2_X1 U16170 ( .A1(n14258), .A2(n6575), .ZN(n14140) );
  NAND2_X1 U16171 ( .A1(n14157), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n14136) );
  OAI21_X1 U16172 ( .B1(n14739), .B2(n14137), .A(n14136), .ZN(n14138) );
  AOI21_X1 U16173 ( .B1(n14259), .B2(n14741), .A(n14138), .ZN(n14139) );
  OAI211_X1 U16174 ( .C1(n14141), .C2(n14337), .A(n14140), .B(n14139), .ZN(
        n14142) );
  AOI21_X1 U16175 ( .B1(n14257), .B2(n14571), .A(n14142), .ZN(n14143) );
  OAI21_X1 U16176 ( .B1(n14263), .B2(n14339), .A(n14143), .ZN(P1_U3274) );
  XOR2_X1 U16177 ( .A(n14144), .B(n14152), .Z(n14145) );
  AOI222_X1 U16178 ( .A1(n14508), .A2(n14178), .B1(n14146), .B2(n14177), .C1(
        n14738), .C2(n14145), .ZN(n14267) );
  INV_X1 U16179 ( .A(n14147), .ZN(n14148) );
  AOI211_X1 U16180 ( .C1(n14265), .C2(n6706), .A(n14745), .B(n14148), .ZN(
        n14264) );
  INV_X1 U16181 ( .A(n14149), .ZN(n14150) );
  AOI22_X1 U16182 ( .A1(n14157), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14150), 
        .B2(n14722), .ZN(n14151) );
  OAI21_X1 U16183 ( .B1(n11936), .B2(n14337), .A(n14151), .ZN(n14155) );
  XNOR2_X1 U16184 ( .A(n14153), .B(n14152), .ZN(n14268) );
  NOR2_X1 U16185 ( .A1(n14268), .A2(n14339), .ZN(n14154) );
  AOI211_X1 U16186 ( .C1(n14264), .C2(n6575), .A(n14155), .B(n14154), .ZN(
        n14156) );
  OAI21_X1 U16187 ( .B1(n14267), .B2(n14157), .A(n14156), .ZN(P1_U3275) );
  AOI21_X1 U16188 ( .B1(n14158), .B2(n14164), .A(n14837), .ZN(n14163) );
  NAND2_X1 U16189 ( .A1(n14159), .A2(n14177), .ZN(n14161) );
  NAND2_X1 U16190 ( .A1(n14546), .A2(n14178), .ZN(n14160) );
  NAND2_X1 U16191 ( .A1(n14161), .A2(n14160), .ZN(n14518) );
  AOI21_X1 U16192 ( .B1(n14163), .B2(n14162), .A(n14518), .ZN(n14581) );
  XNOR2_X1 U16193 ( .A(n14165), .B(n14164), .ZN(n14578) );
  AOI21_X1 U16194 ( .B1(n14176), .B2(n14575), .A(n14745), .ZN(n14166) );
  NAND2_X1 U16195 ( .A1(n14166), .A2(n6706), .ZN(n14577) );
  OAI22_X1 U16196 ( .A1(n14741), .A2(n13958), .B1(n14523), .B2(n14739), .ZN(
        n14167) );
  AOI21_X1 U16197 ( .B1(n14575), .B2(n14743), .A(n14167), .ZN(n14168) );
  OAI21_X1 U16198 ( .B1(n14577), .B2(n14186), .A(n14168), .ZN(n14169) );
  AOI21_X1 U16199 ( .B1(n14578), .B2(n14570), .A(n14169), .ZN(n14170) );
  OAI21_X1 U16200 ( .B1(n14581), .B2(n14157), .A(n14170), .ZN(P1_U3276) );
  XNOR2_X1 U16201 ( .A(n14172), .B(n14171), .ZN(n14585) );
  OAI21_X1 U16202 ( .B1(n14175), .B2(n14174), .A(n14173), .ZN(n14588) );
  OAI211_X1 U16203 ( .C1(n14565), .C2(n14584), .A(n14725), .B(n14176), .ZN(
        n14583) );
  NOR2_X1 U16204 ( .A1(n14741), .A2(n11296), .ZN(n14183) );
  NAND2_X1 U16205 ( .A1(n14508), .A2(n14177), .ZN(n14180) );
  NAND2_X1 U16206 ( .A1(n14507), .A2(n14178), .ZN(n14179) );
  AND2_X1 U16207 ( .A1(n14180), .A2(n14179), .ZN(n14582) );
  OAI22_X1 U16208 ( .A1(n14157), .A2(n14582), .B1(n14514), .B2(n14739), .ZN(
        n14182) );
  AOI211_X1 U16209 ( .C1(n14184), .C2(n14743), .A(n14183), .B(n14182), .ZN(
        n14185) );
  OAI21_X1 U16210 ( .B1(n14583), .B2(n14186), .A(n14185), .ZN(n14187) );
  AOI21_X1 U16211 ( .B1(n14588), .B2(n14570), .A(n14187), .ZN(n14188) );
  OAI21_X1 U16212 ( .B1(n14585), .B2(n14189), .A(n14188), .ZN(P1_U3277) );
  OAI211_X1 U16213 ( .C1(n14191), .C2(n14824), .A(n14190), .B(n14192), .ZN(
        n14269) );
  MUX2_X1 U16214 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14269), .S(n14858), .Z(
        P1_U3559) );
  OAI211_X1 U16215 ( .C1(n14194), .C2(n14824), .A(n14193), .B(n14192), .ZN(
        n14270) );
  MUX2_X1 U16216 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14270), .S(n14858), .Z(
        P1_U3558) );
  OAI211_X1 U16217 ( .C1(n14197), .C2(n14824), .A(n14196), .B(n14195), .ZN(
        n14198) );
  MUX2_X1 U16218 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14271), .S(n14858), .Z(
        P1_U3557) );
  AOI21_X1 U16219 ( .B1(n14203), .B2(n14833), .A(n14202), .ZN(n14204) );
  OAI211_X1 U16220 ( .C1(n14793), .C2(n14206), .A(n14205), .B(n14204), .ZN(
        n14272) );
  MUX2_X1 U16221 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14272), .S(n14858), .Z(
        P1_U3556) );
  INV_X1 U16222 ( .A(n14207), .ZN(n14208) );
  NAND2_X1 U16223 ( .A1(n14208), .A2(n14830), .ZN(n14210) );
  OAI211_X1 U16224 ( .C1(n11907), .C2(n14824), .A(n14210), .B(n14209), .ZN(
        n14211) );
  AOI21_X1 U16225 ( .B1(n14214), .B2(n14833), .A(n14213), .ZN(n14215) );
  OAI211_X1 U16226 ( .C1(n14793), .C2(n14217), .A(n14216), .B(n14215), .ZN(
        n14274) );
  MUX2_X1 U16227 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14274), .S(n14858), .Z(
        P1_U3554) );
  NAND2_X1 U16228 ( .A1(n14218), .A2(n14738), .ZN(n14223) );
  AOI211_X1 U16229 ( .C1(n14221), .C2(n14833), .A(n14220), .B(n14219), .ZN(
        n14222) );
  OAI211_X1 U16230 ( .C1(n14793), .C2(n14224), .A(n14223), .B(n14222), .ZN(
        n14275) );
  MUX2_X1 U16231 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14275), .S(n14858), .Z(
        P1_U3553) );
  NAND2_X1 U16232 ( .A1(n14225), .A2(n14830), .ZN(n14227) );
  OAI211_X1 U16233 ( .C1(n14228), .C2(n14824), .A(n14227), .B(n14226), .ZN(
        n14229) );
  NOR2_X1 U16234 ( .A1(n14230), .A2(n14229), .ZN(n14276) );
  MUX2_X1 U16235 ( .A(n14231), .B(n14276), .S(n14858), .Z(n14232) );
  INV_X1 U16236 ( .A(n14232), .ZN(P1_U3552) );
  AOI211_X1 U16237 ( .C1(n14235), .C2(n14833), .A(n14234), .B(n14233), .ZN(
        n14236) );
  OAI211_X1 U16238 ( .C1(n14793), .C2(n14238), .A(n14237), .B(n14236), .ZN(
        n14279) );
  MUX2_X1 U16239 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14279), .S(n14858), .Z(
        P1_U3551) );
  AOI211_X1 U16240 ( .C1(n7004), .C2(n14833), .A(n14240), .B(n14239), .ZN(
        n14243) );
  NAND2_X1 U16241 ( .A1(n14241), .A2(n14840), .ZN(n14242) );
  OAI211_X1 U16242 ( .C1(n14244), .C2(n14837), .A(n14243), .B(n14242), .ZN(
        n14280) );
  MUX2_X1 U16243 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14280), .S(n14858), .Z(
        P1_U3550) );
  AOI21_X1 U16244 ( .B1(n14246), .B2(n14833), .A(n14245), .ZN(n14247) );
  OAI211_X1 U16245 ( .C1(n14793), .C2(n14249), .A(n14248), .B(n14247), .ZN(
        n14281) );
  MUX2_X1 U16246 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14281), .S(n14858), .Z(
        P1_U3549) );
  OAI211_X1 U16247 ( .C1(n14252), .C2(n14824), .A(n14251), .B(n14250), .ZN(
        n14253) );
  AOI21_X1 U16248 ( .B1(n14254), .B2(n14840), .A(n14253), .ZN(n14255) );
  OAI21_X1 U16249 ( .B1(n14837), .B2(n14256), .A(n14255), .ZN(n14282) );
  MUX2_X1 U16250 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14282), .S(n14858), .Z(
        P1_U3548) );
  NAND2_X1 U16251 ( .A1(n14257), .A2(n14738), .ZN(n14262) );
  AOI211_X1 U16252 ( .C1(n14260), .C2(n14833), .A(n14259), .B(n14258), .ZN(
        n14261) );
  OAI211_X1 U16253 ( .C1(n14793), .C2(n14263), .A(n14262), .B(n14261), .ZN(
        n14283) );
  MUX2_X1 U16254 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14283), .S(n14858), .Z(
        P1_U3547) );
  AOI21_X1 U16255 ( .B1(n14265), .B2(n14833), .A(n14264), .ZN(n14266) );
  OAI211_X1 U16256 ( .C1(n14793), .C2(n14268), .A(n14267), .B(n14266), .ZN(
        n14284) );
  MUX2_X1 U16257 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14284), .S(n14858), .Z(
        P1_U3546) );
  MUX2_X1 U16258 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14269), .S(n14844), .Z(
        P1_U3527) );
  MUX2_X1 U16259 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14270), .S(n14844), .Z(
        P1_U3526) );
  MUX2_X1 U16260 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14272), .S(n14844), .Z(
        P1_U3524) );
  MUX2_X1 U16261 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14274), .S(n14844), .Z(
        P1_U3522) );
  MUX2_X1 U16262 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14275), .S(n14844), .Z(
        P1_U3521) );
  INV_X1 U16263 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n14277) );
  MUX2_X1 U16264 ( .A(n14277), .B(n14276), .S(n14844), .Z(n14278) );
  INV_X1 U16265 ( .A(n14278), .ZN(P1_U3520) );
  MUX2_X1 U16266 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14279), .S(n14844), .Z(
        P1_U3519) );
  MUX2_X1 U16267 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14280), .S(n14844), .Z(
        P1_U3518) );
  MUX2_X1 U16268 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14281), .S(n14844), .Z(
        P1_U3517) );
  MUX2_X1 U16269 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14282), .S(n14844), .Z(
        P1_U3516) );
  MUX2_X1 U16270 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14283), .S(n14844), .Z(
        P1_U3515) );
  MUX2_X1 U16271 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14284), .S(n14844), .Z(
        P1_U3513) );
  NAND2_X1 U16272 ( .A1(n14285), .A2(n14292), .ZN(n14289) );
  NAND2_X1 U16273 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_STATE_REG_SCAN_IN), 
        .ZN(n14286) );
  OR3_X1 U16274 ( .A1(n14287), .A2(P1_IR_REG_30__SCAN_IN), .A3(n14286), .ZN(
        n14288) );
  OAI211_X1 U16275 ( .C1(n14290), .C2(n14298), .A(n14289), .B(n14288), .ZN(
        P1_U3324) );
  OAI222_X1 U16276 ( .A1(n14304), .A2(n14291), .B1(n8290), .B2(P1_U3086), .C1(
        n6778), .C2(n14298), .ZN(P1_U3326) );
  NAND2_X1 U16277 ( .A1(n14293), .A2(n14292), .ZN(n14295) );
  OAI211_X1 U16278 ( .C1(n14296), .C2(n14298), .A(n14295), .B(n14294), .ZN(
        P1_U3328) );
  INV_X1 U16279 ( .A(n14297), .ZN(n14300) );
  OAI222_X1 U16280 ( .A1(n14301), .A2(P1_U3086), .B1(n14304), .B2(n14300), 
        .C1(n14299), .C2(n14298), .ZN(P1_U3329) );
  OAI222_X1 U16281 ( .A1(P1_U3086), .A2(n14305), .B1(n14304), .B2(n14303), 
        .C1(n14302), .C2(n14298), .ZN(P1_U3330) );
  MUX2_X1 U16282 ( .A(n14308), .B(n14307), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16283 ( .A(n14309), .ZN(n14310) );
  MUX2_X1 U16284 ( .A(n14310), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16285 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15051) );
  XOR2_X1 U16286 ( .A(n15051), .B(n14311), .Z(SUB_1596_U62) );
  AOI21_X1 U16287 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14312) );
  OAI21_X1 U16288 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14312), 
        .ZN(U28) );
  AOI21_X1 U16289 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14313) );
  OAI21_X1 U16290 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14313), 
        .ZN(U29) );
  AOI21_X1 U16291 ( .B1(n14316), .B2(n14315), .A(n14314), .ZN(n14317) );
  XOR2_X1 U16292 ( .A(n14317), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  INV_X1 U16293 ( .A(n14318), .ZN(n14319) );
  AOI22_X1 U16294 ( .A1(n14319), .A2(n14325), .B1(SI_4_), .B2(n6727), .ZN(
        n14320) );
  OAI21_X1 U16295 ( .B1(P3_U3151), .B2(n14321), .A(n14320), .ZN(P3_U3291) );
  XOR2_X1 U16296 ( .A(n14323), .B(n14322), .Z(SUB_1596_U57) );
  INV_X1 U16297 ( .A(n14324), .ZN(n14326) );
  AOI22_X1 U16298 ( .A1(n14326), .A2(n14325), .B1(SI_15_), .B2(n6727), .ZN(
        n14327) );
  OAI21_X1 U16299 ( .B1(P3_U3151), .B2(n14328), .A(n14327), .ZN(P3_U3280) );
  XOR2_X1 U16300 ( .A(n6852), .B(n14329), .Z(SUB_1596_U55) );
  AOI21_X1 U16301 ( .B1(n14332), .B2(n14331), .A(n14330), .ZN(n14333) );
  XOR2_X1 U16302 ( .A(n14333), .B(P2_ADDR_REG_9__SCAN_IN), .Z(SUB_1596_U54) );
  INV_X1 U16303 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14967) );
  XOR2_X1 U16304 ( .A(n14967), .B(n14334), .Z(SUB_1596_U70) );
  AOI22_X1 U16305 ( .A1(n14157), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n14335), 
        .B2(n14722), .ZN(n14336) );
  OAI21_X1 U16306 ( .B1(n14338), .B2(n14337), .A(n14336), .ZN(n14342) );
  NOR2_X1 U16307 ( .A1(n14340), .A2(n14339), .ZN(n14341) );
  AOI211_X1 U16308 ( .C1(n14343), .C2(n6575), .A(n14342), .B(n14341), .ZN(
        n14344) );
  OAI21_X1 U16309 ( .B1(n14157), .B2(n14345), .A(n14344), .ZN(P1_U3281) );
  AOI21_X1 U16310 ( .B1(n14348), .B2(n14347), .A(n14346), .ZN(n14349) );
  XOR2_X1 U16311 ( .A(n14349), .B(P2_ADDR_REG_17__SCAN_IN), .Z(SUB_1596_U63)
         );
  AOI21_X1 U16312 ( .B1(n14352), .B2(n14351), .A(n14350), .ZN(n14366) );
  OAI21_X1 U16313 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n14354), .A(n14353), 
        .ZN(n14359) );
  NAND2_X1 U16314 ( .A1(n15149), .A2(n12554), .ZN(n14356) );
  OAI211_X1 U16315 ( .C1(n14357), .C2(n15156), .A(n14356), .B(n14355), .ZN(
        n14358) );
  AOI21_X1 U16316 ( .B1(n14359), .B2(n15220), .A(n14358), .ZN(n14365) );
  AOI21_X1 U16317 ( .B1(n14362), .B2(n14361), .A(n14360), .ZN(n14363) );
  OR2_X1 U16318 ( .A1(n14363), .A2(n15184), .ZN(n14364) );
  OAI211_X1 U16319 ( .C1(n14366), .C2(n15228), .A(n14365), .B(n14364), .ZN(
        P3_U3197) );
  AOI21_X1 U16320 ( .B1(n14368), .B2(n14367), .A(n6638), .ZN(n14386) );
  OAI21_X1 U16321 ( .B1(n14371), .B2(n14370), .A(n14369), .ZN(n14377) );
  NAND2_X1 U16322 ( .A1(n15149), .A2(n14372), .ZN(n14374) );
  OAI211_X1 U16323 ( .C1(n14375), .C2(n15156), .A(n14374), .B(n14373), .ZN(
        n14376) );
  AOI21_X1 U16324 ( .B1(n14377), .B2(n15220), .A(n14376), .ZN(n14385) );
  INV_X1 U16325 ( .A(n14378), .ZN(n14380) );
  NOR2_X1 U16326 ( .A1(n14380), .A2(n14379), .ZN(n14382) );
  AOI21_X1 U16327 ( .B1(n14383), .B2(n14382), .A(n15184), .ZN(n14381) );
  OAI21_X1 U16328 ( .B1(n14383), .B2(n14382), .A(n14381), .ZN(n14384) );
  OAI211_X1 U16329 ( .C1(n14386), .C2(n15228), .A(n14385), .B(n14384), .ZN(
        P3_U3198) );
  AOI21_X1 U16330 ( .B1(n14389), .B2(n14388), .A(n14387), .ZN(n14403) );
  OAI21_X1 U16331 ( .B1(n14391), .B2(P3_REG1_REG_17__SCAN_IN), .A(n14390), 
        .ZN(n14392) );
  AND2_X1 U16332 ( .A1(n14392), .A2(n15220), .ZN(n14400) );
  AOI211_X1 U16333 ( .C1(n14395), .C2(n14394), .A(n15184), .B(n14393), .ZN(
        n14399) );
  OAI22_X1 U16334 ( .A1(n15218), .A2(n14397), .B1(n14396), .B2(n15156), .ZN(
        n14398) );
  NOR4_X1 U16335 ( .A1(n14401), .A2(n14400), .A3(n14399), .A4(n14398), .ZN(
        n14402) );
  OAI21_X1 U16336 ( .B1(n14403), .B2(n15228), .A(n14402), .ZN(P3_U3199) );
  AOI22_X1 U16337 ( .A1(n15149), .A2(n14404), .B1(n15215), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n14419) );
  OAI21_X1 U16338 ( .B1(n14407), .B2(n14406), .A(n14405), .ZN(n14412) );
  OAI21_X1 U16339 ( .B1(n14410), .B2(n14409), .A(n14408), .ZN(n14411) );
  AOI22_X1 U16340 ( .A1(n14412), .A2(n15220), .B1(n15222), .B2(n14411), .ZN(
        n14418) );
  OAI221_X1 U16341 ( .B1(n14415), .B2(n14414), .C1(n14415), .C2(n14413), .A(
        n15151), .ZN(n14416) );
  XNOR2_X1 U16342 ( .A(n14420), .B(n14422), .ZN(n14436) );
  XOR2_X1 U16343 ( .A(n14423), .B(n14422), .Z(n14424) );
  OAI222_X1 U16344 ( .A1(n15294), .A2(n14426), .B1(n15292), .B2(n14425), .C1(
        n14424), .C2(n15299), .ZN(n14434) );
  AOI21_X1 U16345 ( .B1(n14436), .B2(n15250), .A(n14434), .ZN(n14430) );
  NOR2_X1 U16346 ( .A1(n14427), .A2(n15368), .ZN(n14435) );
  AOI22_X1 U16347 ( .A1(n15305), .A2(n14435), .B1(n15253), .B2(n14428), .ZN(
        n14429) );
  OAI221_X1 U16348 ( .B1(n15333), .B2(n14430), .C1(n15330), .C2(n9435), .A(
        n14429), .ZN(P3_U3222) );
  AOI211_X1 U16349 ( .C1(n14433), .C2(n15366), .A(n14432), .B(n14431), .ZN(
        n14439) );
  AOI22_X1 U16350 ( .A1(n15395), .A2(n14439), .B1(n9450), .B2(n15392), .ZN(
        P3_U3471) );
  AOI211_X1 U16351 ( .C1(n14436), .C2(n15366), .A(n14435), .B(n14434), .ZN(
        n14440) );
  INV_X1 U16352 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14437) );
  AOI22_X1 U16353 ( .A1(n15395), .A2(n14440), .B1(n14437), .B2(n15392), .ZN(
        P3_U3470) );
  INV_X1 U16354 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14438) );
  AOI22_X1 U16355 ( .A1(n15379), .A2(n14439), .B1(n14438), .B2(n15378), .ZN(
        P3_U3426) );
  AOI22_X1 U16356 ( .A1(n15379), .A2(n14440), .B1(n9434), .B2(n15378), .ZN(
        P3_U3423) );
  OAI22_X1 U16357 ( .A1(n14444), .A2(n14443), .B1(n14442), .B2(n14441), .ZN(
        n14455) );
  OAI21_X1 U16358 ( .B1(n14447), .B2(n14446), .A(n14445), .ZN(n14449) );
  AOI222_X1 U16359 ( .A1(n14451), .A2(n14461), .B1(n14455), .B2(n14450), .C1(
        n14449), .C2(n14448), .ZN(n14452) );
  NAND2_X1 U16360 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14989)
         );
  OAI211_X1 U16361 ( .C1(n14453), .C2(n14458), .A(n14452), .B(n14989), .ZN(
        P2_U3187) );
  XNOR2_X1 U16362 ( .A(n14454), .B(n14462), .ZN(n14457) );
  AOI21_X1 U16363 ( .B1(n14457), .B2(n14456), .A(n14455), .ZN(n14471) );
  INV_X1 U16364 ( .A(n14458), .ZN(n14459) );
  AOI222_X1 U16365 ( .A1(n14461), .A2(n15058), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n13358), .C1(n14460), .C2(n14459), .ZN(n14469) );
  XNOR2_X1 U16366 ( .A(n14463), .B(n14462), .ZN(n14474) );
  OAI211_X1 U16367 ( .C1(n14472), .C2(n7094), .A(n14465), .B(n14464), .ZN(
        n14470) );
  INV_X1 U16368 ( .A(n14470), .ZN(n14466) );
  AOI22_X1 U16369 ( .A1(n14474), .A2(n15063), .B1(n14467), .B2(n14466), .ZN(
        n14468) );
  OAI211_X1 U16370 ( .C1(n13358), .C2(n14471), .A(n14469), .B(n14468), .ZN(
        P2_U3251) );
  OAI211_X1 U16371 ( .C1(n14472), .C2(n15092), .A(n14471), .B(n14470), .ZN(
        n14473) );
  AOI21_X1 U16372 ( .B1(n14479), .B2(n14474), .A(n14473), .ZN(n14489) );
  AOI22_X1 U16373 ( .A1(n15105), .A2(n14489), .B1(n13132), .B2(n15103), .ZN(
        P2_U3513) );
  OAI211_X1 U16374 ( .C1(n14477), .C2(n15092), .A(n14476), .B(n14475), .ZN(
        n14478) );
  AOI21_X1 U16375 ( .B1(n14480), .B2(n14479), .A(n14478), .ZN(n14490) );
  AOI22_X1 U16376 ( .A1(n15105), .A2(n14490), .B1(n13131), .B2(n15103), .ZN(
        P2_U3512) );
  NAND2_X1 U16377 ( .A1(n14482), .A2(n14481), .ZN(n14483) );
  NAND2_X1 U16378 ( .A1(n14484), .A2(n14483), .ZN(n14485) );
  AOI21_X1 U16379 ( .B1(n14486), .B2(n15097), .A(n14485), .ZN(n14487) );
  AND2_X1 U16380 ( .A1(n14488), .A2(n14487), .ZN(n14492) );
  AOI22_X1 U16381 ( .A1(n15105), .A2(n14492), .B1(n13115), .B2(n15103), .ZN(
        P2_U3511) );
  AOI22_X1 U16382 ( .A1(n15099), .A2(n14489), .B1(n7841), .B2(n15098), .ZN(
        P2_U3472) );
  AOI22_X1 U16383 ( .A1(n15099), .A2(n14490), .B1(n7825), .B2(n15098), .ZN(
        P2_U3469) );
  INV_X1 U16384 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14491) );
  AOI22_X1 U16385 ( .A1(n15099), .A2(n14492), .B1(n14491), .B2(n15098), .ZN(
        P2_U3466) );
  OAI22_X1 U16386 ( .A1(n14494), .A2(n14525), .B1(n14526), .B2(n14493), .ZN(
        n14501) );
  INV_X1 U16387 ( .A(n13840), .ZN(n14497) );
  OAI21_X1 U16388 ( .B1(n14497), .B2(n14496), .A(n14495), .ZN(n14499) );
  AOI21_X1 U16389 ( .B1(n14499), .B2(n14498), .A(n14532), .ZN(n14500) );
  AOI211_X1 U16390 ( .C1(n14598), .C2(n14536), .A(n14501), .B(n14500), .ZN(
        n14503) );
  OAI211_X1 U16391 ( .C1(n14554), .C2(n14504), .A(n14503), .B(n14502), .ZN(
        P1_U3215) );
  XNOR2_X1 U16392 ( .A(n14505), .B(n14506), .ZN(n14511) );
  AOI22_X1 U16393 ( .A1(n14547), .A2(n14508), .B1(n14545), .B2(n14507), .ZN(
        n14509) );
  OAI21_X1 U16394 ( .B1(n14584), .B2(n14549), .A(n14509), .ZN(n14510) );
  AOI21_X1 U16395 ( .B1(n14511), .B2(n14551), .A(n14510), .ZN(n14513) );
  OAI211_X1 U16396 ( .C1(n14554), .C2(n14514), .A(n14513), .B(n14512), .ZN(
        P1_U3226) );
  XNOR2_X1 U16397 ( .A(n14515), .B(n14516), .ZN(n14519) );
  AOI222_X1 U16398 ( .A1(n14536), .A2(n14575), .B1(n14551), .B2(n14519), .C1(
        n14518), .C2(n14517), .ZN(n14522) );
  INV_X1 U16399 ( .A(n14520), .ZN(n14521) );
  OAI211_X1 U16400 ( .C1(n14554), .C2(n14523), .A(n14522), .B(n14521), .ZN(
        P1_U3228) );
  OAI22_X1 U16401 ( .A1(n14527), .A2(n14526), .B1(n14525), .B2(n14524), .ZN(
        n14535) );
  AOI21_X1 U16402 ( .B1(n11793), .B2(n14529), .A(n14528), .ZN(n14530) );
  INV_X1 U16403 ( .A(n14530), .ZN(n14533) );
  AOI21_X1 U16404 ( .B1(n14533), .B2(n14531), .A(n14532), .ZN(n14534) );
  AOI211_X1 U16405 ( .C1(n14537), .C2(n14536), .A(n14535), .B(n14534), .ZN(
        n14539) );
  OAI211_X1 U16406 ( .C1(n14554), .C2(n14540), .A(n14539), .B(n14538), .ZN(
        P1_U3236) );
  OAI21_X1 U16407 ( .B1(n14543), .B2(n14542), .A(n14541), .ZN(n14552) );
  AOI22_X1 U16408 ( .A1(n14547), .A2(n14546), .B1(n14545), .B2(n14544), .ZN(
        n14548) );
  OAI21_X1 U16409 ( .B1(n14561), .B2(n14549), .A(n14548), .ZN(n14550) );
  AOI21_X1 U16410 ( .B1(n14552), .B2(n14551), .A(n14550), .ZN(n14553) );
  NAND2_X1 U16411 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14693)
         );
  OAI211_X1 U16412 ( .C1(n14554), .C2(n14574), .A(n14553), .B(n14693), .ZN(
        P1_U3241) );
  OAI22_X1 U16413 ( .A1(n14558), .A2(n14557), .B1(n14556), .B2(n14555), .ZN(
        n14591) );
  INV_X1 U16414 ( .A(n14591), .ZN(n14559) );
  OAI211_X1 U16415 ( .C1(n14561), .C2(n14560), .A(n14559), .B(n14741), .ZN(
        n14562) );
  OAI21_X1 U16416 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14741), .A(n14562), 
        .ZN(n14573) );
  XNOR2_X1 U16417 ( .A(n14563), .B(n14567), .ZN(n14596) );
  INV_X1 U16418 ( .A(n14564), .ZN(n14566) );
  AOI211_X1 U16419 ( .C1(n14592), .C2(n14566), .A(n14745), .B(n14565), .ZN(
        n14590) );
  XNOR2_X1 U16420 ( .A(n14568), .B(n14567), .ZN(n14594) );
  INV_X1 U16421 ( .A(n14594), .ZN(n14569) );
  AOI222_X1 U16422 ( .A1(n14596), .A2(n14571), .B1(n6575), .B2(n14590), .C1(
        n14570), .C2(n14569), .ZN(n14572) );
  OAI211_X1 U16423 ( .C1(n14739), .C2(n14574), .A(n14573), .B(n14572), .ZN(
        P1_U3278) );
  NAND2_X1 U16424 ( .A1(n14575), .A2(n14833), .ZN(n14576) );
  AND2_X1 U16425 ( .A1(n14577), .A2(n14576), .ZN(n14580) );
  NAND2_X1 U16426 ( .A1(n14578), .A2(n14840), .ZN(n14579) );
  AOI22_X1 U16427 ( .A1(n14858), .A2(n14611), .B1(n13938), .B2(n14856), .ZN(
        P1_U3545) );
  OAI211_X1 U16428 ( .C1(n14584), .C2(n14824), .A(n14583), .B(n14582), .ZN(
        n14587) );
  NOR2_X1 U16429 ( .A1(n14585), .A2(n14837), .ZN(n14586) );
  AOI211_X1 U16430 ( .C1(n14840), .C2(n14588), .A(n14587), .B(n14586), .ZN(
        n14612) );
  AOI22_X1 U16431 ( .A1(n14858), .A2(n14612), .B1(n14589), .B2(n14856), .ZN(
        P1_U3544) );
  AOI211_X1 U16432 ( .C1(n14592), .C2(n14833), .A(n14591), .B(n14590), .ZN(
        n14593) );
  OAI21_X1 U16433 ( .B1(n14594), .B2(n14793), .A(n14593), .ZN(n14595) );
  AOI21_X1 U16434 ( .B1(n14596), .B2(n14738), .A(n14595), .ZN(n14613) );
  AOI22_X1 U16435 ( .A1(n14858), .A2(n14613), .B1(n8551), .B2(n14856), .ZN(
        P1_U3543) );
  AOI21_X1 U16436 ( .B1(n14598), .B2(n14833), .A(n14597), .ZN(n14601) );
  INV_X1 U16437 ( .A(n14599), .ZN(n14600) );
  OAI211_X1 U16438 ( .C1(n14602), .C2(n14793), .A(n14601), .B(n14600), .ZN(
        n14603) );
  NOR2_X1 U16439 ( .A1(n14604), .A2(n14603), .ZN(n14615) );
  AOI22_X1 U16440 ( .A1(n14858), .A2(n14615), .B1(n8527), .B2(n14856), .ZN(
        P1_U3542) );
  OAI21_X1 U16441 ( .B1(n14606), .B2(n14824), .A(n14605), .ZN(n14608) );
  AOI211_X1 U16442 ( .C1(n14609), .C2(n14840), .A(n14608), .B(n14607), .ZN(
        n14616) );
  AOI22_X1 U16443 ( .A1(n14858), .A2(n14616), .B1(n10243), .B2(n14856), .ZN(
        P1_U3539) );
  INV_X1 U16444 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14610) );
  AOI22_X1 U16445 ( .A1(n14844), .A2(n14611), .B1(n14610), .B2(n14842), .ZN(
        P1_U3510) );
  AOI22_X1 U16446 ( .A1(n14844), .A2(n14612), .B1(n8571), .B2(n14842), .ZN(
        P1_U3507) );
  AOI22_X1 U16447 ( .A1(n14844), .A2(n14613), .B1(n8552), .B2(n14842), .ZN(
        P1_U3504) );
  AOI22_X1 U16448 ( .A1(n14844), .A2(n14615), .B1(n14614), .B2(n14842), .ZN(
        P1_U3501) );
  AOI22_X1 U16449 ( .A1(n14844), .A2(n14616), .B1(n8487), .B2(n14842), .ZN(
        P1_U3492) );
  AOI21_X1 U16450 ( .B1(n14618), .B2(n6708), .A(n14617), .ZN(n14619) );
  XOR2_X1 U16451 ( .A(n14619), .B(P2_ADDR_REG_11__SCAN_IN), .Z(SUB_1596_U69)
         );
  XNOR2_X1 U16452 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n14620), .ZN(SUB_1596_U68)
         );
  AOI21_X1 U16453 ( .B1(n14622), .B2(n14621), .A(n6715), .ZN(n14623) );
  XOR2_X1 U16454 ( .A(n14623), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  AOI21_X1 U16455 ( .B1(n14626), .B2(n14625), .A(n14624), .ZN(n14627) );
  XOR2_X1 U16456 ( .A(n14627), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  OAI21_X1 U16457 ( .B1(n14630), .B2(n14629), .A(n14628), .ZN(n14631) );
  XOR2_X1 U16458 ( .A(n14631), .B(n15002), .Z(SUB_1596_U65) );
  AOI21_X1 U16459 ( .B1(n14634), .B2(n14633), .A(n14632), .ZN(n14635) );
  XOR2_X1 U16460 ( .A(n14635), .B(P2_ADDR_REG_16__SCAN_IN), .Z(SUB_1596_U64)
         );
  AOI22_X1 U16461 ( .A1(n14675), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n14659) );
  AND3_X1 U16462 ( .A1(n14638), .A2(n14637), .A3(n14636), .ZN(n14639) );
  NOR3_X1 U16463 ( .A1(n14690), .A2(n14640), .A3(n14639), .ZN(n14648) );
  INV_X1 U16464 ( .A(n14641), .ZN(n14644) );
  NAND3_X1 U16465 ( .A1(n14644), .A2(n14643), .A3(n14642), .ZN(n14645) );
  AND3_X1 U16466 ( .A1(n14684), .A2(n14646), .A3(n14645), .ZN(n14647) );
  AOI211_X1 U16467 ( .C1(n14687), .C2(n14649), .A(n14648), .B(n14647), .ZN(
        n14658) );
  MUX2_X1 U16468 ( .A(n14652), .B(n14651), .S(n14650), .Z(n14654) );
  NAND2_X1 U16469 ( .A1(n14654), .A2(n14653), .ZN(n14656) );
  OAI211_X1 U16470 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n14657), .A(n14656), .B(
        n14655), .ZN(n14677) );
  NAND3_X1 U16471 ( .A1(n14659), .A2(n14658), .A3(n14677), .ZN(P1_U3245) );
  OAI211_X1 U16472 ( .C1(n14662), .C2(n14661), .A(n14684), .B(n14660), .ZN(
        n14671) );
  INV_X1 U16473 ( .A(n14663), .ZN(n14668) );
  NAND3_X1 U16474 ( .A1(n14666), .A2(n14665), .A3(n14664), .ZN(n14667) );
  NAND3_X1 U16475 ( .A1(n14669), .A2(n14668), .A3(n14667), .ZN(n14670) );
  OAI211_X1 U16476 ( .C1(n14673), .C2(n14672), .A(n14671), .B(n14670), .ZN(
        n14674) );
  INV_X1 U16477 ( .A(n14674), .ZN(n14679) );
  NAND2_X1 U16478 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n14675), .ZN(n14676) );
  NAND4_X1 U16479 ( .A1(n14679), .A2(n14678), .A3(n14677), .A4(n14676), .ZN(
        P1_U3247) );
  AOI21_X1 U16480 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14681), .A(n14680), 
        .ZN(n14691) );
  OAI21_X1 U16481 ( .B1(n14683), .B2(n8551), .A(n14682), .ZN(n14685) );
  NAND2_X1 U16482 ( .A1(n14685), .A2(n14684), .ZN(n14689) );
  NAND2_X1 U16483 ( .A1(n14687), .A2(n14686), .ZN(n14688) );
  OAI211_X1 U16484 ( .C1(n14691), .C2(n14690), .A(n14689), .B(n14688), .ZN(
        n14692) );
  INV_X1 U16485 ( .A(n14692), .ZN(n14694) );
  OAI211_X1 U16486 ( .C1(n14696), .C2(n14695), .A(n14694), .B(n14693), .ZN(
        P1_U3258) );
  XNOR2_X1 U16487 ( .A(n14697), .B(n14698), .ZN(n14702) );
  XOR2_X1 U16488 ( .A(n14699), .B(n14698), .Z(n14706) );
  NOR2_X1 U16489 ( .A1(n14706), .A2(n14734), .ZN(n14700) );
  AOI211_X1 U16490 ( .C1(n14702), .C2(n14738), .A(n14701), .B(n14700), .ZN(
        n14826) );
  INV_X1 U16491 ( .A(n14703), .ZN(n14704) );
  AOI222_X1 U16492 ( .A1(n14705), .A2(n14743), .B1(P1_REG2_REG_9__SCAN_IN), 
        .B2(n14157), .C1(n14722), .C2(n14704), .ZN(n14712) );
  INV_X1 U16493 ( .A(n14706), .ZN(n14829) );
  INV_X1 U16494 ( .A(n14707), .ZN(n14709) );
  OAI211_X1 U16495 ( .C1(n14709), .C2(n14825), .A(n14725), .B(n14708), .ZN(
        n14823) );
  INV_X1 U16496 ( .A(n14823), .ZN(n14710) );
  AOI22_X1 U16497 ( .A1(n14829), .A2(n14748), .B1(n6575), .B2(n14710), .ZN(
        n14711) );
  OAI211_X1 U16498 ( .C1(n14157), .C2(n14826), .A(n14712), .B(n14711), .ZN(
        P1_U3284) );
  XNOR2_X1 U16499 ( .A(n14713), .B(n14714), .ZN(n14800) );
  XNOR2_X1 U16500 ( .A(n14715), .B(n14714), .ZN(n14716) );
  NOR2_X1 U16501 ( .A1(n14716), .A2(n14837), .ZN(n14717) );
  AOI211_X1 U16502 ( .C1(n14719), .C2(n14800), .A(n14718), .B(n14717), .ZN(
        n14797) );
  INV_X1 U16503 ( .A(n14720), .ZN(n14721) );
  AOI222_X1 U16504 ( .A1(n14723), .A2(n14743), .B1(P1_REG2_REG_5__SCAN_IN), 
        .B2(n14157), .C1(n14722), .C2(n14721), .ZN(n14728) );
  OAI211_X1 U16505 ( .C1(n6723), .C2(n14796), .A(n14725), .B(n14724), .ZN(
        n14795) );
  INV_X1 U16506 ( .A(n14795), .ZN(n14726) );
  AOI22_X1 U16507 ( .A1(n14800), .A2(n14748), .B1(n6575), .B2(n14726), .ZN(
        n14727) );
  OAI211_X1 U16508 ( .C1(n14157), .C2(n14797), .A(n14728), .B(n14727), .ZN(
        P1_U3288) );
  OAI21_X1 U16509 ( .B1(n14730), .B2(n14733), .A(n14729), .ZN(n14737) );
  INV_X1 U16510 ( .A(n14731), .ZN(n14736) );
  XNOR2_X1 U16511 ( .A(n14732), .B(n14733), .ZN(n14785) );
  NOR2_X1 U16512 ( .A1(n14785), .A2(n14734), .ZN(n14735) );
  AOI211_X1 U16513 ( .C1(n14738), .C2(n14737), .A(n14736), .B(n14735), .ZN(
        n14784) );
  OAI22_X1 U16514 ( .A1(n14741), .A2(n14740), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14739), .ZN(n14742) );
  AOI21_X1 U16515 ( .B1(n14743), .B2(n14782), .A(n14742), .ZN(n14751) );
  INV_X1 U16516 ( .A(n14785), .ZN(n14749) );
  AOI211_X1 U16517 ( .C1(n14782), .C2(n14746), .A(n14745), .B(n14744), .ZN(
        n14781) );
  AOI22_X1 U16518 ( .A1(n14749), .A2(n14748), .B1(n14781), .B2(n6575), .ZN(
        n14750) );
  OAI211_X1 U16519 ( .C1(n14157), .C2(n14784), .A(n14751), .B(n14750), .ZN(
        P1_U3290) );
  AND2_X1 U16520 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14760), .ZN(P1_U3294) );
  NOR2_X1 U16521 ( .A1(n14759), .A2(n14752), .ZN(P1_U3295) );
  AND2_X1 U16522 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14760), .ZN(P1_U3296) );
  AND2_X1 U16523 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14760), .ZN(P1_U3297) );
  AND2_X1 U16524 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14760), .ZN(P1_U3298) );
  AND2_X1 U16525 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14760), .ZN(P1_U3299) );
  AND2_X1 U16526 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14760), .ZN(P1_U3300) );
  AND2_X1 U16527 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14760), .ZN(P1_U3301) );
  AND2_X1 U16528 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14760), .ZN(P1_U3302) );
  AND2_X1 U16529 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14760), .ZN(P1_U3303) );
  AND2_X1 U16530 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14760), .ZN(P1_U3304) );
  AND2_X1 U16531 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14760), .ZN(P1_U3305) );
  AND2_X1 U16532 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14760), .ZN(P1_U3306) );
  NOR2_X1 U16533 ( .A1(n14759), .A2(n14753), .ZN(P1_U3307) );
  NOR2_X1 U16534 ( .A1(n14759), .A2(n14754), .ZN(P1_U3308) );
  NOR2_X1 U16535 ( .A1(n14759), .A2(n14755), .ZN(P1_U3309) );
  AND2_X1 U16536 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14760), .ZN(P1_U3310) );
  NOR2_X1 U16537 ( .A1(n14759), .A2(n14756), .ZN(P1_U3311) );
  NOR2_X1 U16538 ( .A1(n14759), .A2(n14757), .ZN(P1_U3312) );
  AND2_X1 U16539 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14760), .ZN(P1_U3313) );
  AND2_X1 U16540 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14760), .ZN(P1_U3314) );
  AND2_X1 U16541 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14760), .ZN(P1_U3315) );
  NOR2_X1 U16542 ( .A1(n14759), .A2(n14758), .ZN(P1_U3316) );
  AND2_X1 U16543 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14760), .ZN(P1_U3317) );
  AND2_X1 U16544 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14760), .ZN(P1_U3318) );
  AND2_X1 U16545 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14760), .ZN(P1_U3319) );
  AND2_X1 U16546 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14760), .ZN(P1_U3320) );
  AND2_X1 U16547 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14760), .ZN(P1_U3321) );
  AND2_X1 U16548 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14760), .ZN(P1_U3322) );
  AND2_X1 U16549 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14760), .ZN(P1_U3323) );
  INV_X1 U16550 ( .A(n14761), .ZN(n14762) );
  AOI21_X1 U16551 ( .B1(n14793), .B2(n14837), .A(n14762), .ZN(n14763) );
  AOI211_X1 U16552 ( .C1(n14765), .C2(n8319), .A(n14764), .B(n14763), .ZN(
        n14845) );
  INV_X1 U16553 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n14766) );
  AOI22_X1 U16554 ( .A1(n14844), .A2(n14845), .B1(n14766), .B2(n14842), .ZN(
        P1_U3459) );
  INV_X1 U16555 ( .A(n14767), .ZN(n14769) );
  OAI211_X1 U16556 ( .C1(n14770), .C2(n14824), .A(n14769), .B(n14768), .ZN(
        n14773) );
  INV_X1 U16557 ( .A(n14771), .ZN(n14772) );
  AOI211_X1 U16558 ( .C1(n14830), .C2(n14774), .A(n14773), .B(n14772), .ZN(
        n14846) );
  AOI22_X1 U16559 ( .A1(n14844), .A2(n14846), .B1(n8301), .B2(n14842), .ZN(
        P1_U3462) );
  OAI21_X1 U16560 ( .B1(n14776), .B2(n14824), .A(n14775), .ZN(n14777) );
  AOI21_X1 U16561 ( .B1(n14778), .B2(n14830), .A(n14777), .ZN(n14779) );
  AND2_X1 U16562 ( .A1(n14780), .A2(n14779), .ZN(n14847) );
  AOI22_X1 U16563 ( .A1(n14844), .A2(n14847), .B1(n8330), .B2(n14842), .ZN(
        P1_U3465) );
  AOI21_X1 U16564 ( .B1(n14782), .B2(n14833), .A(n14781), .ZN(n14783) );
  OAI211_X1 U16565 ( .C1(n14786), .C2(n14785), .A(n14784), .B(n14783), .ZN(
        n14787) );
  INV_X1 U16566 ( .A(n14787), .ZN(n14849) );
  AOI22_X1 U16567 ( .A1(n14844), .A2(n14849), .B1(n8344), .B2(n14842), .ZN(
        P1_U3468) );
  AOI21_X1 U16568 ( .B1(n14789), .B2(n14833), .A(n14788), .ZN(n14790) );
  OAI211_X1 U16569 ( .C1(n14793), .C2(n14792), .A(n14791), .B(n14790), .ZN(
        n14794) );
  INV_X1 U16570 ( .A(n14794), .ZN(n14850) );
  AOI22_X1 U16571 ( .A1(n14844), .A2(n14850), .B1(n8368), .B2(n14842), .ZN(
        P1_U3471) );
  OAI21_X1 U16572 ( .B1(n14796), .B2(n14824), .A(n14795), .ZN(n14799) );
  INV_X1 U16573 ( .A(n14797), .ZN(n14798) );
  AOI211_X1 U16574 ( .C1(n14830), .C2(n14800), .A(n14799), .B(n14798), .ZN(
        n14851) );
  INV_X1 U16575 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14801) );
  AOI22_X1 U16576 ( .A1(n14844), .A2(n14851), .B1(n14801), .B2(n14842), .ZN(
        P1_U3474) );
  INV_X1 U16577 ( .A(n14802), .ZN(n14803) );
  OAI21_X1 U16578 ( .B1(n14804), .B2(n14824), .A(n14803), .ZN(n14805) );
  AOI21_X1 U16579 ( .B1(n14806), .B2(n14830), .A(n14805), .ZN(n14807) );
  AOI22_X1 U16580 ( .A1(n14844), .A2(n14852), .B1(n14809), .B2(n14842), .ZN(
        P1_U3477) );
  OAI21_X1 U16581 ( .B1(n14811), .B2(n14824), .A(n14810), .ZN(n14813) );
  AOI211_X1 U16582 ( .C1(n14830), .C2(n14814), .A(n14813), .B(n14812), .ZN(
        n14853) );
  INV_X1 U16583 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14815) );
  AOI22_X1 U16584 ( .A1(n14844), .A2(n14853), .B1(n14815), .B2(n14842), .ZN(
        P1_U3480) );
  OAI21_X1 U16585 ( .B1(n14817), .B2(n14824), .A(n14816), .ZN(n14818) );
  AOI21_X1 U16586 ( .B1(n14819), .B2(n14840), .A(n14818), .ZN(n14820) );
  AND2_X1 U16587 ( .A1(n14821), .A2(n14820), .ZN(n14854) );
  AOI22_X1 U16588 ( .A1(n14844), .A2(n14854), .B1(n14822), .B2(n14842), .ZN(
        P1_U3483) );
  OAI21_X1 U16589 ( .B1(n14825), .B2(n14824), .A(n14823), .ZN(n14828) );
  INV_X1 U16590 ( .A(n14826), .ZN(n14827) );
  AOI211_X1 U16591 ( .C1(n14830), .C2(n14829), .A(n14828), .B(n14827), .ZN(
        n14855) );
  INV_X1 U16592 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14831) );
  AOI22_X1 U16593 ( .A1(n14844), .A2(n14855), .B1(n14831), .B2(n14842), .ZN(
        P1_U3486) );
  AOI21_X1 U16594 ( .B1(n14834), .B2(n14833), .A(n14832), .ZN(n14835) );
  OAI211_X1 U16595 ( .C1(n14838), .C2(n14837), .A(n14836), .B(n14835), .ZN(
        n14839) );
  AOI21_X1 U16596 ( .B1(n14841), .B2(n14840), .A(n14839), .ZN(n14857) );
  INV_X1 U16597 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14843) );
  AOI22_X1 U16598 ( .A1(n14844), .A2(n14857), .B1(n14843), .B2(n14842), .ZN(
        P1_U3489) );
  AOI22_X1 U16599 ( .A1(n14858), .A2(n14845), .B1(n8312), .B2(n14856), .ZN(
        P1_U3528) );
  AOI22_X1 U16600 ( .A1(n14858), .A2(n14846), .B1(n8300), .B2(n14856), .ZN(
        P1_U3529) );
  AOI22_X1 U16601 ( .A1(n14858), .A2(n14847), .B1(n8329), .B2(n14856), .ZN(
        P1_U3530) );
  INV_X1 U16602 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n14848) );
  AOI22_X1 U16603 ( .A1(n14858), .A2(n14849), .B1(n14848), .B2(n14856), .ZN(
        P1_U3531) );
  AOI22_X1 U16604 ( .A1(n14858), .A2(n14850), .B1(n10097), .B2(n14856), .ZN(
        P1_U3532) );
  AOI22_X1 U16605 ( .A1(n14858), .A2(n14851), .B1(n8384), .B2(n14856), .ZN(
        P1_U3533) );
  AOI22_X1 U16606 ( .A1(n14858), .A2(n14852), .B1(n8400), .B2(n14856), .ZN(
        P1_U3534) );
  AOI22_X1 U16607 ( .A1(n14858), .A2(n14853), .B1(n8421), .B2(n14856), .ZN(
        P1_U3535) );
  AOI22_X1 U16608 ( .A1(n14858), .A2(n14854), .B1(n10125), .B2(n14856), .ZN(
        P1_U3536) );
  AOI22_X1 U16609 ( .A1(n14858), .A2(n14855), .B1(n10122), .B2(n14856), .ZN(
        P1_U3537) );
  AOI22_X1 U16610 ( .A1(n14858), .A2(n14857), .B1(n10188), .B2(n14856), .ZN(
        P1_U3538) );
  NOR2_X1 U16611 ( .A1(n14872), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16612 ( .A1(n14872), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n14871) );
  OAI211_X1 U16613 ( .C1(n14862), .C2(n14861), .A(n15035), .B(n14860), .ZN(
        n14867) );
  OAI211_X1 U16614 ( .C1(n14865), .C2(n14864), .A(n15041), .B(n14863), .ZN(
        n14866) );
  OAI211_X1 U16615 ( .C1(n15046), .C2(n14868), .A(n14867), .B(n14866), .ZN(
        n14869) );
  INV_X1 U16616 ( .A(n14869), .ZN(n14870) );
  NAND2_X1 U16617 ( .A1(n14871), .A2(n14870), .ZN(P2_U3215) );
  AOI22_X1 U16618 ( .A1(n14872), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14886) );
  OAI21_X1 U16619 ( .B1(n14875), .B2(n14874), .A(n14873), .ZN(n14883) );
  OAI211_X1 U16620 ( .C1(n14878), .C2(n14877), .A(n15041), .B(n14876), .ZN(
        n14882) );
  INV_X1 U16621 ( .A(n14879), .ZN(n14880) );
  NAND2_X1 U16622 ( .A1(n15028), .A2(n14880), .ZN(n14881) );
  OAI211_X1 U16623 ( .C1(n14883), .C2(n15018), .A(n14882), .B(n14881), .ZN(
        n14884) );
  INV_X1 U16624 ( .A(n14884), .ZN(n14885) );
  NAND2_X1 U16625 ( .A1(n14886), .A2(n14885), .ZN(P2_U3216) );
  OAI21_X1 U16626 ( .B1(n14889), .B2(n14888), .A(n14887), .ZN(n14896) );
  OAI211_X1 U16627 ( .C1(n14892), .C2(n14891), .A(n15041), .B(n14890), .ZN(
        n14895) );
  NAND2_X1 U16628 ( .A1(n15028), .A2(n14893), .ZN(n14894) );
  OAI211_X1 U16629 ( .C1(n15018), .C2(n14896), .A(n14895), .B(n14894), .ZN(
        n14897) );
  INV_X1 U16630 ( .A(n14897), .ZN(n14899) );
  OAI211_X1 U16631 ( .C1(n15050), .C2(n14900), .A(n14899), .B(n14898), .ZN(
        P2_U3218) );
  OAI21_X1 U16632 ( .B1(n14903), .B2(n14902), .A(n14901), .ZN(n14910) );
  OAI211_X1 U16633 ( .C1(n14906), .C2(n14905), .A(n15041), .B(n14904), .ZN(
        n14909) );
  NAND2_X1 U16634 ( .A1(n15028), .A2(n14907), .ZN(n14908) );
  OAI211_X1 U16635 ( .C1(n14910), .C2(n15018), .A(n14909), .B(n14908), .ZN(
        n14911) );
  INV_X1 U16636 ( .A(n14911), .ZN(n14913) );
  OAI211_X1 U16637 ( .C1(n15050), .C2(n14914), .A(n14913), .B(n14912), .ZN(
        P2_U3220) );
  OAI211_X1 U16638 ( .C1(n14917), .C2(n14916), .A(n15035), .B(n14915), .ZN(
        n14922) );
  OAI211_X1 U16639 ( .C1(n14920), .C2(n14919), .A(n15041), .B(n14918), .ZN(
        n14921) );
  OAI211_X1 U16640 ( .C1(n15046), .C2(n14923), .A(n14922), .B(n14921), .ZN(
        n14924) );
  INV_X1 U16641 ( .A(n14924), .ZN(n14926) );
  NAND2_X1 U16642 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n14925) );
  OAI211_X1 U16643 ( .C1(n14927), .C2(n15050), .A(n14926), .B(n14925), .ZN(
        P2_U3221) );
  OAI211_X1 U16644 ( .C1(n14930), .C2(n14929), .A(n15035), .B(n14928), .ZN(
        n14935) );
  OAI211_X1 U16645 ( .C1(n14933), .C2(n14932), .A(n15041), .B(n14931), .ZN(
        n14934) );
  OAI211_X1 U16646 ( .C1(n15046), .C2(n14936), .A(n14935), .B(n14934), .ZN(
        n14937) );
  INV_X1 U16647 ( .A(n14937), .ZN(n14939) );
  OAI211_X1 U16648 ( .C1(n6852), .C2(n15050), .A(n14939), .B(n14938), .ZN(
        P2_U3222) );
  NAND2_X1 U16649 ( .A1(n14941), .A2(n14940), .ZN(n14942) );
  NAND2_X1 U16650 ( .A1(n14943), .A2(n14942), .ZN(n14945) );
  AOI22_X1 U16651 ( .A1(n14945), .A2(n15035), .B1(n14944), .B2(n15028), .ZN(
        n14951) );
  AND2_X1 U16652 ( .A1(n14947), .A2(n14946), .ZN(n14948) );
  OAI21_X1 U16653 ( .B1(n14949), .B2(n14948), .A(n15041), .ZN(n14950) );
  AND2_X1 U16654 ( .A1(n14951), .A2(n14950), .ZN(n14953) );
  OAI211_X1 U16655 ( .C1(n14954), .C2(n15050), .A(n14953), .B(n14952), .ZN(
        P2_U3223) );
  OAI21_X1 U16656 ( .B1(n14956), .B2(n14955), .A(n15041), .ZN(n14958) );
  NOR2_X1 U16657 ( .A1(n14958), .A2(n14957), .ZN(n14963) );
  AOI211_X1 U16658 ( .C1(n14961), .C2(n14960), .A(n15018), .B(n14959), .ZN(
        n14962) );
  AOI211_X1 U16659 ( .C1(n15028), .C2(n14964), .A(n14963), .B(n14962), .ZN(
        n14966) );
  OAI211_X1 U16660 ( .C1(n14967), .C2(n15050), .A(n14966), .B(n14965), .ZN(
        P2_U3224) );
  AOI211_X1 U16661 ( .C1(n14970), .C2(n14969), .A(n15018), .B(n14968), .ZN(
        n14975) );
  AOI211_X1 U16662 ( .C1(n14973), .C2(n14972), .A(n15022), .B(n14971), .ZN(
        n14974) );
  AOI211_X1 U16663 ( .C1(n15028), .C2(n14976), .A(n14975), .B(n14974), .ZN(
        n14978) );
  NAND2_X1 U16664 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n14977)
         );
  OAI211_X1 U16665 ( .C1(n14979), .C2(n15050), .A(n14978), .B(n14977), .ZN(
        P2_U3227) );
  AOI211_X1 U16666 ( .C1(n14982), .C2(n14981), .A(n15022), .B(n14980), .ZN(
        n14987) );
  AOI211_X1 U16667 ( .C1(n14985), .C2(n14984), .A(n14983), .B(n15018), .ZN(
        n14986) );
  AOI211_X1 U16668 ( .C1(n15028), .C2(n14988), .A(n14987), .B(n14986), .ZN(
        n14990) );
  OAI211_X1 U16669 ( .C1(n14991), .C2(n15050), .A(n14990), .B(n14989), .ZN(
        P2_U3228) );
  AOI211_X1 U16670 ( .C1(n14993), .C2(n11754), .A(n14992), .B(n15018), .ZN(
        n14998) );
  AOI211_X1 U16671 ( .C1(n14996), .C2(n14995), .A(n14994), .B(n15022), .ZN(
        n14997) );
  AOI211_X1 U16672 ( .C1(n15028), .C2(n14999), .A(n14998), .B(n14997), .ZN(
        n15001) );
  NAND2_X1 U16673 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n15000)
         );
  OAI211_X1 U16674 ( .C1(n15002), .C2(n15050), .A(n15001), .B(n15000), .ZN(
        P2_U3229) );
  AOI211_X1 U16675 ( .C1(n15005), .C2(n15004), .A(n15022), .B(n15003), .ZN(
        n15011) );
  INV_X1 U16676 ( .A(n15006), .ZN(n15007) );
  AOI211_X1 U16677 ( .C1(n15009), .C2(n15008), .A(n15018), .B(n15007), .ZN(
        n15010) );
  AOI211_X1 U16678 ( .C1(n15028), .C2(n15012), .A(n15011), .B(n15010), .ZN(
        n15014) );
  OAI211_X1 U16679 ( .C1(n15015), .C2(n15050), .A(n15014), .B(n15013), .ZN(
        P2_U3230) );
  NOR2_X1 U16680 ( .A1(n15017), .A2(n15016), .ZN(n15019) );
  NOR3_X1 U16681 ( .A1(n15020), .A2(n15019), .A3(n15018), .ZN(n15026) );
  AOI211_X1 U16682 ( .C1(n15024), .C2(n15023), .A(n15022), .B(n15021), .ZN(
        n15025) );
  AOI211_X1 U16683 ( .C1(n15028), .C2(n15027), .A(n15026), .B(n15025), .ZN(
        n15030) );
  OAI211_X1 U16684 ( .C1(n15031), .C2(n15050), .A(n15030), .B(n15029), .ZN(
        P2_U3231) );
  OAI21_X1 U16685 ( .B1(n15034), .B2(n15033), .A(n15032), .ZN(n15036) );
  NAND2_X1 U16686 ( .A1(n15036), .A2(n15035), .ZN(n15044) );
  NAND2_X1 U16687 ( .A1(n15038), .A2(n15037), .ZN(n15042) );
  INV_X1 U16688 ( .A(n15039), .ZN(n15040) );
  NAND3_X1 U16689 ( .A1(n15042), .A2(n15041), .A3(n15040), .ZN(n15043) );
  OAI211_X1 U16690 ( .C1(n15046), .C2(n15045), .A(n15044), .B(n15043), .ZN(
        n15047) );
  INV_X1 U16691 ( .A(n15047), .ZN(n15049) );
  OAI211_X1 U16692 ( .C1(n15051), .C2(n15050), .A(n15049), .B(n15048), .ZN(
        P2_U3232) );
  OAI22_X1 U16693 ( .A1(n15055), .A2(n15054), .B1(n15053), .B2(n15052), .ZN(
        n15056) );
  AOI21_X1 U16694 ( .B1(n15058), .B2(n15057), .A(n15056), .ZN(n15059) );
  OAI21_X1 U16695 ( .B1(n15061), .B2(n15060), .A(n15059), .ZN(n15062) );
  AOI21_X1 U16696 ( .B1(n15064), .B2(n15063), .A(n15062), .ZN(n15065) );
  OAI21_X1 U16697 ( .B1(n13358), .B2(n15066), .A(n15065), .ZN(P2_U3258) );
  AND2_X1 U16698 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15071), .ZN(P2_U3266) );
  AND2_X1 U16699 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15071), .ZN(P2_U3267) );
  AND2_X1 U16700 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15071), .ZN(P2_U3268) );
  AND2_X1 U16701 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15071), .ZN(P2_U3269) );
  AND2_X1 U16702 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15071), .ZN(P2_U3270) );
  AND2_X1 U16703 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15071), .ZN(P2_U3271) );
  AND2_X1 U16704 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15071), .ZN(P2_U3272) );
  AND2_X1 U16705 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15071), .ZN(P2_U3273) );
  NOR2_X1 U16706 ( .A1(n15073), .A2(n15068), .ZN(P2_U3274) );
  NOR2_X1 U16707 ( .A1(n15073), .A2(n15069), .ZN(P2_U3275) );
  AND2_X1 U16708 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15071), .ZN(P2_U3276) );
  AND2_X1 U16709 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15071), .ZN(P2_U3277) );
  NOR2_X1 U16710 ( .A1(n15073), .A2(n15070), .ZN(P2_U3278) );
  AND2_X1 U16711 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15071), .ZN(P2_U3279) );
  AND2_X1 U16712 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15071), .ZN(P2_U3280) );
  AND2_X1 U16713 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15071), .ZN(P2_U3281) );
  AND2_X1 U16714 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15071), .ZN(P2_U3282) );
  AND2_X1 U16715 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15071), .ZN(P2_U3283) );
  AND2_X1 U16716 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15071), .ZN(P2_U3284) );
  AND2_X1 U16717 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15071), .ZN(P2_U3285) );
  AND2_X1 U16718 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15071), .ZN(P2_U3286) );
  AND2_X1 U16719 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15071), .ZN(P2_U3287) );
  AND2_X1 U16720 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15071), .ZN(P2_U3288) );
  AND2_X1 U16721 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15071), .ZN(P2_U3289) );
  AND2_X1 U16722 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15071), .ZN(P2_U3290) );
  AND2_X1 U16723 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15071), .ZN(P2_U3291) );
  AND2_X1 U16724 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15071), .ZN(P2_U3292) );
  AND2_X1 U16725 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15071), .ZN(P2_U3293) );
  AND2_X1 U16726 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15071), .ZN(P2_U3294) );
  NOR2_X1 U16727 ( .A1(n15073), .A2(n15072), .ZN(P2_U3295) );
  OAI22_X1 U16728 ( .A1(n15076), .A2(n15074), .B1(P2_D_REG_0__SCAN_IN), .B2(
        n15078), .ZN(n15075) );
  INV_X1 U16729 ( .A(n15075), .ZN(P2_U3416) );
  AOI22_X1 U16730 ( .A1(n15078), .A2(n15077), .B1(n8224), .B2(n15076), .ZN(
        P2_U3417) );
  OAI21_X1 U16731 ( .B1(n15080), .B2(n15092), .A(n15079), .ZN(n15082) );
  AOI211_X1 U16732 ( .C1(n15097), .C2(n15083), .A(n15082), .B(n15081), .ZN(
        n15100) );
  AOI22_X1 U16733 ( .A1(n15099), .A2(n15100), .B1(n7585), .B2(n15098), .ZN(
        P2_U3436) );
  INV_X1 U16734 ( .A(n15084), .ZN(n15085) );
  OAI21_X1 U16735 ( .B1(n15086), .B2(n15092), .A(n15085), .ZN(n15088) );
  AOI211_X1 U16736 ( .C1(n15097), .C2(n15089), .A(n15088), .B(n15087), .ZN(
        n15102) );
  AOI22_X1 U16737 ( .A1(n15099), .A2(n15102), .B1(n7641), .B2(n15098), .ZN(
        P2_U3442) );
  INV_X1 U16738 ( .A(n15090), .ZN(n15096) );
  OAI21_X1 U16739 ( .B1(n15093), .B2(n15092), .A(n15091), .ZN(n15095) );
  AOI211_X1 U16740 ( .C1(n15097), .C2(n15096), .A(n15095), .B(n15094), .ZN(
        n15104) );
  AOI22_X1 U16741 ( .A1(n15099), .A2(n15104), .B1(n7762), .B2(n15098), .ZN(
        P2_U3460) );
  AOI22_X1 U16742 ( .A1(n15105), .A2(n15100), .B1(n10341), .B2(n15103), .ZN(
        P2_U3501) );
  AOI22_X1 U16743 ( .A1(n15105), .A2(n15102), .B1(n15101), .B2(n15103), .ZN(
        P2_U3503) );
  AOI22_X1 U16744 ( .A1(n15105), .A2(n15104), .B1(n7758), .B2(n15103), .ZN(
        P2_U3509) );
  NOR2_X1 U16745 ( .A1(P3_U3897), .A2(n15215), .ZN(P3_U3150) );
  AOI22_X1 U16746 ( .A1(n15220), .A2(n15107), .B1(n15151), .B2(n15106), .ZN(
        n15116) );
  AOI22_X1 U16747 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n15215), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n15115) );
  NAND3_X1 U16748 ( .A1(n15228), .A2(n15108), .A3(n15184), .ZN(n15111) );
  INV_X1 U16749 ( .A(n15109), .ZN(n15110) );
  AOI22_X1 U16750 ( .A1(n15111), .A2(n15110), .B1(P3_IR_REG_0__SCAN_IN), .B2(
        n15149), .ZN(n15114) );
  OR3_X1 U16751 ( .A1(n15184), .A2(P3_IR_REG_0__SCAN_IN), .A3(n15112), .ZN(
        n15113) );
  NAND4_X1 U16752 ( .A1(n15116), .A2(n15115), .A3(n15114), .A4(n15113), .ZN(
        P3_U3182) );
  AOI21_X1 U16753 ( .B1(n9381), .B2(n15118), .A(n15117), .ZN(n15133) );
  INV_X1 U16754 ( .A(n15119), .ZN(n15121) );
  NAND2_X1 U16755 ( .A1(n15121), .A2(n15120), .ZN(n15122) );
  XNOR2_X1 U16756 ( .A(n15123), .B(n15122), .ZN(n15125) );
  OAI22_X1 U16757 ( .A1(n15125), .A2(n15184), .B1(n15124), .B2(n15218), .ZN(
        n15126) );
  AOI211_X1 U16758 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15215), .A(n15127), .B(
        n15126), .ZN(n15132) );
  OAI21_X1 U16759 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15129), .A(n15128), .ZN(
        n15130) );
  NAND2_X1 U16760 ( .A1(n15130), .A2(n15220), .ZN(n15131) );
  OAI211_X1 U16761 ( .C1(n15133), .C2(n15228), .A(n15132), .B(n15131), .ZN(
        P3_U3191) );
  OAI21_X1 U16762 ( .B1(n15136), .B2(n15135), .A(n15134), .ZN(n15138) );
  AOI21_X1 U16763 ( .B1(n15138), .B2(n15220), .A(n15137), .ZN(n15154) );
  INV_X1 U16764 ( .A(n15139), .ZN(n15143) );
  INV_X1 U16765 ( .A(n15140), .ZN(n15142) );
  OAI21_X1 U16766 ( .B1(n15143), .B2(n15142), .A(n15141), .ZN(n15152) );
  AOI21_X1 U16767 ( .B1(n15146), .B2(n15145), .A(n15144), .ZN(n15147) );
  INV_X1 U16768 ( .A(n15147), .ZN(n15148) );
  AOI222_X1 U16769 ( .A1(n15152), .A2(n15151), .B1(n15150), .B2(n15149), .C1(
        n15148), .C2(n15222), .ZN(n15153) );
  OAI211_X1 U16770 ( .C1(n15156), .C2(n15155), .A(n15154), .B(n15153), .ZN(
        P3_U3192) );
  AOI21_X1 U16771 ( .B1(n9435), .B2(n15158), .A(n15157), .ZN(n15172) );
  OAI21_X1 U16772 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n15160), .A(n15159), 
        .ZN(n15165) );
  AOI21_X1 U16773 ( .B1(n15215), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n15161), 
        .ZN(n15162) );
  OAI21_X1 U16774 ( .B1(n15218), .B2(n15163), .A(n15162), .ZN(n15164) );
  AOI21_X1 U16775 ( .B1(n15165), .B2(n15220), .A(n15164), .ZN(n15171) );
  OAI21_X1 U16776 ( .B1(n15168), .B2(n15167), .A(n15166), .ZN(n15169) );
  NAND2_X1 U16777 ( .A1(n15222), .A2(n15169), .ZN(n15170) );
  OAI211_X1 U16778 ( .C1(n15172), .C2(n15228), .A(n15171), .B(n15170), .ZN(
        P3_U3193) );
  AOI21_X1 U16779 ( .B1(n15175), .B2(n15174), .A(n15173), .ZN(n15191) );
  OAI21_X1 U16780 ( .B1(n15178), .B2(n15177), .A(n15176), .ZN(n15183) );
  AOI21_X1 U16781 ( .B1(n15215), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n15179), 
        .ZN(n15180) );
  OAI21_X1 U16782 ( .B1(n15218), .B2(n15181), .A(n15180), .ZN(n15182) );
  AOI21_X1 U16783 ( .B1(n15183), .B2(n15220), .A(n15182), .ZN(n15190) );
  AOI21_X1 U16784 ( .B1(n15186), .B2(n15185), .A(n15184), .ZN(n15188) );
  NAND2_X1 U16785 ( .A1(n15188), .A2(n15187), .ZN(n15189) );
  OAI211_X1 U16786 ( .C1(n15191), .C2(n15228), .A(n15190), .B(n15189), .ZN(
        P3_U3194) );
  AOI21_X1 U16787 ( .B1(n15194), .B2(n15193), .A(n15192), .ZN(n15208) );
  OAI21_X1 U16788 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n15196), .A(n15195), 
        .ZN(n15201) );
  AOI21_X1 U16789 ( .B1(n15215), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n15197), 
        .ZN(n15198) );
  OAI21_X1 U16790 ( .B1(n15218), .B2(n15199), .A(n15198), .ZN(n15200) );
  AOI21_X1 U16791 ( .B1(n15201), .B2(n15220), .A(n15200), .ZN(n15207) );
  OAI21_X1 U16792 ( .B1(n15204), .B2(n15203), .A(n15202), .ZN(n15205) );
  NAND2_X1 U16793 ( .A1(n15205), .A2(n15222), .ZN(n15206) );
  OAI211_X1 U16794 ( .C1(n15208), .C2(n15228), .A(n15207), .B(n15206), .ZN(
        P3_U3195) );
  AOI21_X1 U16795 ( .B1(n6717), .B2(n15210), .A(n15209), .ZN(n15229) );
  OAI21_X1 U16796 ( .B1(n15213), .B2(n15212), .A(n15211), .ZN(n15221) );
  AOI21_X1 U16797 ( .B1(n15215), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n15214), 
        .ZN(n15216) );
  OAI21_X1 U16798 ( .B1(n15218), .B2(n15217), .A(n15216), .ZN(n15219) );
  AOI21_X1 U16799 ( .B1(n15221), .B2(n15220), .A(n15219), .ZN(n15227) );
  OAI211_X1 U16800 ( .C1(n15225), .C2(n15224), .A(n15223), .B(n15222), .ZN(
        n15226) );
  OAI211_X1 U16801 ( .C1(n15229), .C2(n15228), .A(n15227), .B(n15226), .ZN(
        P3_U3196) );
  XNOR2_X1 U16802 ( .A(n15230), .B(n15232), .ZN(n15376) );
  XNOR2_X1 U16803 ( .A(n15231), .B(n15232), .ZN(n15237) );
  OAI22_X1 U16804 ( .A1(n15234), .A2(n15294), .B1(n15233), .B2(n15292), .ZN(
        n15235) );
  AOI21_X1 U16805 ( .B1(n15376), .B2(n15297), .A(n15235), .ZN(n15236) );
  OAI21_X1 U16806 ( .B1(n15237), .B2(n15299), .A(n15236), .ZN(n15374) );
  AOI21_X1 U16807 ( .B1(n15329), .B2(n15376), .A(n15374), .ZN(n15241) );
  NOR2_X1 U16808 ( .A1(n15238), .A2(n15368), .ZN(n15375) );
  AOI22_X1 U16809 ( .A1(n15305), .A2(n15375), .B1(n15253), .B2(n15239), .ZN(
        n15240) );
  OAI221_X1 U16810 ( .B1(n15333), .B2(n15241), .C1(n15330), .C2(n12548), .A(
        n15240), .ZN(P3_U3223) );
  XNOR2_X1 U16811 ( .A(n15243), .B(n15242), .ZN(n15365) );
  OAI21_X1 U16812 ( .B1(n15246), .B2(n15245), .A(n15244), .ZN(n15248) );
  AOI222_X1 U16813 ( .A1(n15319), .A2(n15248), .B1(n15277), .B2(n15323), .C1(
        n15247), .C2(n15322), .ZN(n15249) );
  INV_X1 U16814 ( .A(n15249), .ZN(n15363) );
  AOI21_X1 U16815 ( .B1(n15250), .B2(n15365), .A(n15363), .ZN(n15255) );
  NOR2_X1 U16816 ( .A1(n15251), .A2(n15368), .ZN(n15364) );
  AOI22_X1 U16817 ( .A1(n15305), .A2(n15364), .B1(n15253), .B2(n15252), .ZN(
        n15254) );
  OAI221_X1 U16818 ( .B1(n15333), .B2(n15255), .C1(n15330), .C2(n9361), .A(
        n15254), .ZN(P3_U3225) );
  XNOR2_X1 U16819 ( .A(n15257), .B(n15256), .ZN(n15258) );
  OAI222_X1 U16820 ( .A1(n15292), .A2(n15260), .B1(n15294), .B2(n15259), .C1(
        n15258), .C2(n15299), .ZN(n15359) );
  OAI22_X1 U16821 ( .A1(n15330), .A2(n9343), .B1(n15312), .B2(n15261), .ZN(
        n15268) );
  XNOR2_X1 U16822 ( .A(n15263), .B(n15262), .ZN(n15361) );
  NOR2_X1 U16823 ( .A1(n15264), .A2(n15368), .ZN(n15360) );
  AOI22_X1 U16824 ( .A1(n15361), .A2(n15265), .B1(n15305), .B2(n15360), .ZN(
        n15266) );
  INV_X1 U16825 ( .A(n15266), .ZN(n15267) );
  AOI211_X1 U16826 ( .C1(n15330), .C2(n15359), .A(n15268), .B(n15267), .ZN(
        n15269) );
  INV_X1 U16827 ( .A(n15269), .ZN(P3_U3226) );
  NAND2_X1 U16828 ( .A1(n15270), .A2(n15271), .ZN(n15273) );
  INV_X1 U16829 ( .A(n15272), .ZN(n15275) );
  XNOR2_X1 U16830 ( .A(n15273), .B(n15275), .ZN(n15280) );
  INV_X1 U16831 ( .A(n15280), .ZN(n15358) );
  OAI211_X1 U16832 ( .C1(n6721), .C2(n15275), .A(n15319), .B(n15274), .ZN(
        n15279) );
  AOI22_X1 U16833 ( .A1(n15277), .A2(n15322), .B1(n15323), .B2(n15276), .ZN(
        n15278) );
  OAI211_X1 U16834 ( .C1(n15327), .C2(n15280), .A(n15279), .B(n15278), .ZN(
        n15356) );
  AOI21_X1 U16835 ( .B1(n15329), .B2(n15358), .A(n15356), .ZN(n15285) );
  AND2_X1 U16836 ( .A1(n15281), .A2(n15301), .ZN(n15357) );
  NOR2_X1 U16837 ( .A1(n15312), .A2(n15282), .ZN(n15283) );
  AOI21_X1 U16838 ( .B1(n15305), .B2(n15357), .A(n15283), .ZN(n15284) );
  OAI221_X1 U16839 ( .B1(n15333), .B2(n15285), .C1(n15330), .C2(n10669), .A(
        n15284), .ZN(P3_U3227) );
  NAND2_X1 U16840 ( .A1(n15287), .A2(n15286), .ZN(n15289) );
  XNOR2_X1 U16841 ( .A(n15289), .B(n15288), .ZN(n15350) );
  XNOR2_X1 U16842 ( .A(n15291), .B(n15290), .ZN(n15300) );
  OAI22_X1 U16843 ( .A1(n15295), .A2(n15294), .B1(n15293), .B2(n15292), .ZN(
        n15296) );
  AOI21_X1 U16844 ( .B1(n15350), .B2(n15297), .A(n15296), .ZN(n15298) );
  OAI21_X1 U16845 ( .B1(n15300), .B2(n15299), .A(n15298), .ZN(n15348) );
  AOI21_X1 U16846 ( .B1(n15329), .B2(n15350), .A(n15348), .ZN(n15307) );
  AND2_X1 U16847 ( .A1(n15302), .A2(n15301), .ZN(n15349) );
  NOR2_X1 U16848 ( .A1(n15312), .A2(n15303), .ZN(n15304) );
  AOI21_X1 U16849 ( .B1(n15305), .B2(n15349), .A(n15304), .ZN(n15306) );
  OAI221_X1 U16850 ( .B1(n15333), .B2(n15307), .C1(n15330), .C2(n9283), .A(
        n15306), .ZN(P3_U3229) );
  XNOR2_X1 U16851 ( .A(n15309), .B(n15308), .ZN(n15326) );
  INV_X1 U16852 ( .A(n15326), .ZN(n15341) );
  NOR2_X1 U16853 ( .A1(n15310), .A2(n15368), .ZN(n15340) );
  INV_X1 U16854 ( .A(n15340), .ZN(n15314) );
  OAI22_X1 U16855 ( .A1(n15314), .A2(n15313), .B1(n15312), .B2(n15311), .ZN(
        n15328) );
  INV_X1 U16856 ( .A(n15315), .ZN(n15321) );
  AND3_X1 U16857 ( .A1(n15318), .A2(n15317), .A3(n15316), .ZN(n15320) );
  OAI21_X1 U16858 ( .B1(n15321), .B2(n15320), .A(n15319), .ZN(n15325) );
  AOI22_X1 U16859 ( .A1(n15323), .A2(n10491), .B1(n9277), .B2(n15322), .ZN(
        n15324) );
  OAI211_X1 U16860 ( .C1(n15327), .C2(n15326), .A(n15325), .B(n15324), .ZN(
        n15339) );
  AOI211_X1 U16861 ( .C1(n15329), .C2(n15341), .A(n15328), .B(n15339), .ZN(
        n15331) );
  AOI22_X1 U16862 ( .A1(n15333), .A2(n15332), .B1(n15331), .B2(n15330), .ZN(
        P3_U3231) );
  INV_X1 U16863 ( .A(n15334), .ZN(n15337) );
  INV_X1 U16864 ( .A(n15335), .ZN(n15336) );
  AOI211_X1 U16865 ( .C1(n15377), .C2(n15338), .A(n15337), .B(n15336), .ZN(
        n15381) );
  AOI22_X1 U16866 ( .A1(n15379), .A2(n15381), .B1(n9236), .B2(n15378), .ZN(
        P3_U3393) );
  AOI211_X1 U16867 ( .C1(n15341), .C2(n15377), .A(n15340), .B(n15339), .ZN(
        n15382) );
  INV_X1 U16868 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15342) );
  AOI22_X1 U16869 ( .A1(n15379), .A2(n15382), .B1(n15342), .B2(n15378), .ZN(
        P3_U3396) );
  INV_X1 U16870 ( .A(n15343), .ZN(n15344) );
  AOI211_X1 U16871 ( .C1(n15346), .C2(n15377), .A(n15345), .B(n15344), .ZN(
        n15383) );
  INV_X1 U16872 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15347) );
  AOI22_X1 U16873 ( .A1(n15379), .A2(n15383), .B1(n15347), .B2(n15378), .ZN(
        P3_U3399) );
  AOI211_X1 U16874 ( .C1(n15350), .C2(n15377), .A(n15349), .B(n15348), .ZN(
        n15384) );
  INV_X1 U16875 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15351) );
  AOI22_X1 U16876 ( .A1(n15379), .A2(n15384), .B1(n15351), .B2(n15378), .ZN(
        P3_U3402) );
  INV_X1 U16877 ( .A(n15352), .ZN(n15355) );
  AOI211_X1 U16878 ( .C1(n15355), .C2(n15377), .A(n15354), .B(n15353), .ZN(
        n15386) );
  AOI22_X1 U16879 ( .A1(n15379), .A2(n15386), .B1(n9303), .B2(n15378), .ZN(
        P3_U3405) );
  AOI211_X1 U16880 ( .C1(n15358), .C2(n15377), .A(n15357), .B(n15356), .ZN(
        n15387) );
  AOI22_X1 U16881 ( .A1(n15379), .A2(n15387), .B1(n9327), .B2(n15378), .ZN(
        P3_U3408) );
  AOI211_X1 U16882 ( .C1(n15361), .C2(n15366), .A(n15360), .B(n15359), .ZN(
        n15388) );
  INV_X1 U16883 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15362) );
  AOI22_X1 U16884 ( .A1(n15379), .A2(n15388), .B1(n15362), .B2(n15378), .ZN(
        P3_U3411) );
  AOI211_X1 U16885 ( .C1(n15366), .C2(n15365), .A(n15364), .B(n15363), .ZN(
        n15390) );
  AOI22_X1 U16886 ( .A1(n15379), .A2(n15390), .B1(n9360), .B2(n15378), .ZN(
        P3_U3414) );
  INV_X1 U16887 ( .A(n15367), .ZN(n15372) );
  NOR2_X1 U16888 ( .A1(n15369), .A2(n15368), .ZN(n15371) );
  AOI211_X1 U16889 ( .C1(n15372), .C2(n15377), .A(n15371), .B(n15370), .ZN(
        n15391) );
  INV_X1 U16890 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15373) );
  AOI22_X1 U16891 ( .A1(n15379), .A2(n15391), .B1(n15373), .B2(n15378), .ZN(
        P3_U3417) );
  AOI211_X1 U16892 ( .C1(n15377), .C2(n15376), .A(n15375), .B(n15374), .ZN(
        n15394) );
  AOI22_X1 U16893 ( .A1(n15379), .A2(n15394), .B1(n9404), .B2(n15378), .ZN(
        P3_U3420) );
  INV_X1 U16894 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15380) );
  AOI22_X1 U16895 ( .A1(n15395), .A2(n15381), .B1(n15380), .B2(n15392), .ZN(
        P3_U3460) );
  AOI22_X1 U16896 ( .A1(n15395), .A2(n15382), .B1(n10437), .B2(n15392), .ZN(
        P3_U3461) );
  AOI22_X1 U16897 ( .A1(n15395), .A2(n15383), .B1(n9261), .B2(n15392), .ZN(
        P3_U3462) );
  AOI22_X1 U16898 ( .A1(n15395), .A2(n15384), .B1(n9280), .B2(n15392), .ZN(
        P3_U3463) );
  INV_X1 U16899 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15385) );
  AOI22_X1 U16900 ( .A1(n15395), .A2(n15386), .B1(n15385), .B2(n15392), .ZN(
        P3_U3464) );
  AOI22_X1 U16901 ( .A1(n15395), .A2(n15387), .B1(n10554), .B2(n15392), .ZN(
        P3_U3465) );
  AOI22_X1 U16902 ( .A1(n15395), .A2(n15388), .B1(n9340), .B2(n15392), .ZN(
        P3_U3466) );
  AOI22_X1 U16903 ( .A1(n15395), .A2(n15390), .B1(n15389), .B2(n15392), .ZN(
        P3_U3467) );
  AOI22_X1 U16904 ( .A1(n15395), .A2(n15391), .B1(n9377), .B2(n15392), .ZN(
        P3_U3468) );
  AOI22_X1 U16905 ( .A1(n15395), .A2(n15394), .B1(n15393), .B2(n15392), .ZN(
        P3_U3469) );
  XOR2_X1 U16906 ( .A(n15397), .B(n15396), .Z(SUB_1596_U59) );
  XOR2_X1 U16907 ( .A(n15399), .B(n15398), .Z(SUB_1596_U58) );
  AOI21_X1 U16908 ( .B1(n15401), .B2(n15400), .A(n15410), .ZN(SUB_1596_U53) );
  XOR2_X1 U16909 ( .A(n15403), .B(n15402), .Z(SUB_1596_U56) );
  OAI21_X1 U16910 ( .B1(n15406), .B2(n15405), .A(n15404), .ZN(n15408) );
  XOR2_X1 U16911 ( .A(n15408), .B(n15407), .Z(SUB_1596_U60) );
  XOR2_X1 U16912 ( .A(n15410), .B(n15409), .Z(SUB_1596_U5) );
  INV_X2 U7674 ( .A(n10064), .ZN(n8612) );
  CLKBUF_X1 U7331 ( .A(n11484), .Z(n6743) );
  AND4_X1 U7357 ( .A1(n7546), .A2(n7545), .A3(n7544), .A4(n7547), .ZN(n7373)
         );
  CLKBUF_X1 U7414 ( .A(n7942), .Z(n7943) );
  CLKBUF_X1 U7765 ( .A(n8484), .Z(n6587) );
  CLKBUF_X1 U8435 ( .A(n7638), .Z(n8125) );
  CLKBUF_X2 U9197 ( .A(n7608), .Z(n9105) );
endmodule

