

module b21_C_AntiSAT_k_256_9 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, 
        keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, 
        keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, 
        keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, 
        keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, 
        keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, 
        keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, 
        keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, 
        keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, 
        keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, 
        keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, 
        keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, 
        keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, 
        keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, 
        keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, 
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, 
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, 
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, 
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, 
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, 
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, 
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, 
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, 
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, 
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249, 
        keyinput250, keyinput251, keyinput252, keyinput253, keyinput254, 
        keyinput255, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, 
        ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, 
        ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, 
        ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, 
        ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, 
        P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, 
        P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, 
        P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, 
        P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, 
        P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, 
        P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, 
        P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, 
        P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, 
        P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, 
        P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, 
        P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, 
        P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, 
        P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, 
        P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, 
        P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, 
        P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, 
        P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, 
        P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, 
        P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, 
        P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4478, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10469;

  XNOR2_X1 U4982 ( .A(n5698), .B(n5697), .ZN(n7746) );
  CLKBUF_X2 U4983 ( .A(n5961), .Z(n4478) );
  XNOR2_X2 U4984 ( .A(n5059), .B(n5058), .ZN(n6808) );
  INV_X1 U4985 ( .A(n5967), .ZN(n4894) );
  INV_X1 U4986 ( .A(n5968), .ZN(n6297) );
  INV_X1 U4987 ( .A(n6724), .ZN(n5936) );
  NAND2_X1 U4988 ( .A1(n5853), .A2(n9458), .ZN(n5140) );
  NAND2_X1 U4989 ( .A1(n6208), .A2(n6207), .ZN(n8977) );
  NAND2_X1 U4990 ( .A1(n6178), .A2(n6177), .ZN(n8994) );
  INV_X2 U4991 ( .A(n10193), .ZN(n9774) );
  NAND2_X2 U4992 ( .A1(n6388), .A2(n6391), .ZN(n7757) );
  OAI21_X2 U4993 ( .B1(n4953), .B2(n5771), .A(n4951), .ZN(n4954) );
  OAI21_X1 U4994 ( .B1(n8836), .B2(n4721), .A(n4718), .ZN(n8785) );
  OAI21_X2 U4995 ( .B1(n5547), .B2(n4840), .A(n4838), .ZN(n5596) );
  NAND2_X1 U4997 ( .A1(n6832), .A2(n6724), .ZN(n5961) );
  XNOR2_X2 U4998 ( .A(n5395), .B(n5391), .ZN(n6769) );
  OAI22_X2 U4999 ( .A1(n7756), .A2(n7755), .B1(n10372), .B2(n7754), .ZN(n7758)
         );
  NAND2_X2 U5000 ( .A1(n7710), .A2(n7709), .ZN(n7756) );
  XNOR2_X2 U5001 ( .A(n5675), .B(n5674), .ZN(n7656) );
  NAND2_X2 U5002 ( .A1(n5650), .A2(n5649), .ZN(n5675) );
  AOI21_X2 U5003 ( .B1(n10167), .B2(P1_REG2_REG_17__SCAN_IN), .A(n10162), .ZN(
        n9515) );
  INV_X1 U5004 ( .A(n5817), .ZN(n5793) );
  OAI21_X2 U5005 ( .B1(n6883), .B2(P1_REG2_REG_8__SCAN_IN), .A(n10081), .ZN(
        n10099) );
  OAI21_X2 U5006 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7506), .A(n7505), .ZN(
        n10111) );
  XNOR2_X2 U5007 ( .A(n5645), .B(n5646), .ZN(n7594) );
  CLKBUF_X1 U5008 ( .A(n8753), .Z(n8754) );
  NAND2_X1 U5009 ( .A1(n6199), .A2(n6198), .ZN(n8982) );
  NAND2_X1 U5010 ( .A1(n7970), .A2(n4896), .ZN(n8116) );
  INV_X1 U5011 ( .A(n10346), .ZN(n7279) );
  NAND2_X1 U5012 ( .A1(n6702), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8628) );
  CLKBUF_X3 U5013 ( .A(n8100), .Z(n5755) );
  NAND2_X2 U5014 ( .A1(n6476), .A2(n6475), .ZN(n7081) );
  AND4_X1 U5015 ( .A1(n5974), .A2(n5973), .A3(n5972), .A4(n5971), .ZN(n7460)
         );
  AND4_X1 U5016 ( .A1(n6001), .A2(n6000), .A3(n5999), .A4(n5998), .ZN(n6559)
         );
  BUF_X1 U5017 ( .A(n5140), .Z(n6777) );
  AOI21_X1 U5018 ( .B1(n6612), .B2(n7090), .A(n6329), .ZN(n6511) );
  NAND2_X1 U5019 ( .A1(n6275), .A2(n6449), .ZN(n8494) );
  OAI21_X1 U5020 ( .B1(n4972), .B2(n4969), .A(n4967), .ZN(n9659) );
  NAND2_X1 U5021 ( .A1(n5496), .A2(n5495), .ZN(n9157) );
  NAND2_X1 U5022 ( .A1(n9056), .A2(n9054), .ZN(n9059) );
  NAND2_X1 U5023 ( .A1(n6220), .A2(n6219), .ZN(n8972) );
  OAI21_X1 U5024 ( .B1(n7956), .B2(n7955), .A(n7954), .ZN(n8064) );
  NAND2_X1 U5025 ( .A1(n8900), .A2(n6163), .ZN(n8881) );
  NAND2_X1 U5026 ( .A1(n7794), .A2(n4667), .ZN(n4666) );
  NAND2_X1 U5027 ( .A1(n4958), .A2(n4520), .ZN(n7794) );
  OAI21_X1 U5028 ( .B1(n7960), .B2(n4768), .A(n4765), .ZN(n9765) );
  OAI21_X1 U5029 ( .B1(n7898), .B2(n7897), .A(n7896), .ZN(n7934) );
  NAND2_X1 U5030 ( .A1(n6189), .A2(n6188), .ZN(n8987) );
  NAND2_X1 U5031 ( .A1(n6590), .A2(n6589), .ZN(n7839) );
  NAND2_X1 U5032 ( .A1(n7879), .A2(n4521), .ZN(n7970) );
  OR2_X1 U5033 ( .A1(n8910), .A2(n9010), .ZN(n8908) );
  CLKBUF_X1 U5034 ( .A(n8998), .Z(n4584) );
  NOR3_X1 U5035 ( .A1(n7881), .A2(n4744), .A3(n9016), .ZN(n4743) );
  NAND2_X1 U5036 ( .A1(n6127), .A2(n6126), .ZN(n9016) );
  OR2_X1 U5037 ( .A1(n7877), .A2(n7889), .ZN(n6388) );
  NAND2_X1 U5038 ( .A1(n7634), .A2(n7565), .ZN(n7633) );
  NAND2_X1 U5039 ( .A1(n5150), .A2(n5149), .ZN(n7009) );
  OAI21_X1 U5040 ( .B1(n5423), .B2(n5422), .A(n5421), .ZN(n5446) );
  NAND2_X1 U5041 ( .A1(n5325), .A2(n5324), .ZN(n10236) );
  AND2_X1 U5042 ( .A1(n7218), .A2(n9214), .ZN(n9259) );
  NAND2_X1 U5043 ( .A1(n5288), .A2(n5287), .ZN(n4836) );
  AND2_X2 U5044 ( .A1(n7151), .A2(n7150), .ZN(n10255) );
  NAND2_X2 U5045 ( .A1(n7200), .A2(n8912), .ZN(n8915) );
  NAND4_X2 U5046 ( .A1(n5154), .A2(n5153), .A3(n5152), .A4(n5151), .ZN(n9477)
         );
  NAND4_X2 U5048 ( .A1(n5180), .A2(n5179), .A3(n5178), .A4(n5177), .ZN(n9476)
         );
  NAND4_X2 U5049 ( .A1(n5105), .A2(n5104), .A3(n5103), .A4(n5102), .ZN(n7153)
         );
  NAND2_X1 U5050 ( .A1(n5236), .A2(n5235), .ZN(n5268) );
  AOI21_X1 U5051 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n10069), .A(n6815), .ZN(
        n6816) );
  INV_X1 U5052 ( .A(n5175), .ZN(n8100) );
  AND3_X1 U5053 ( .A1(n5194), .A2(n5193), .A3(n5192), .ZN(n10210) );
  NAND4_X1 U5054 ( .A1(n5991), .A2(n5990), .A3(n5989), .A4(n5988), .ZN(n8645)
         );
  AND3_X1 U5055 ( .A1(n5166), .A2(n5165), .A3(n5164), .ZN(n7322) );
  AND4_X1 U5056 ( .A1(n5946), .A2(n5945), .A3(n5944), .A4(n5943), .ZN(n7298)
         );
  AND3_X1 U5057 ( .A1(n5965), .A2(n5964), .A3(n5963), .ZN(n7174) );
  NAND2_X1 U5058 ( .A1(n4963), .A2(n4964), .ZN(n5086) );
  INV_X1 U5059 ( .A(n8538), .ZN(n10338) );
  CLKBUF_X3 U5060 ( .A(n5954), .Z(n5967) );
  INV_X1 U5061 ( .A(n4478), .ZN(n6176) );
  OR2_X1 U5062 ( .A1(n5960), .A2(n6727), .ZN(n4594) );
  OR2_X1 U5063 ( .A1(n10056), .A2(n10057), .ZN(n10058) );
  NAND2_X2 U5064 ( .A1(n5140), .A2(n5936), .ZN(n9173) );
  AND2_X2 U5065 ( .A1(n6710), .A2(n10178), .ZN(n5817) );
  NAND2_X1 U5066 ( .A1(n9045), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U5067 ( .A1(n9453), .A2(n7467), .ZN(n10178) );
  AND2_X1 U5068 ( .A1(n5910), .A2(n4927), .ZN(n5913) );
  INV_X2 U5069 ( .A(n8014), .ZN(n4480) );
  INV_X2 U5070 ( .A(n8010), .ZN(n4481) );
  NAND4_X1 U5071 ( .A1(n5899), .A2(n5900), .A3(n4898), .A4(n5908), .ZN(n6512)
         );
  NAND2_X1 U5072 ( .A1(n4889), .A2(n4891), .ZN(n5057) );
  NOR2_X1 U5073 ( .A1(n5906), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n4898) );
  AND2_X1 U5074 ( .A1(n5940), .A2(n5939), .ZN(n9909) );
  AND4_X1 U5075 ( .A1(n5401), .A2(n5042), .A3(n5092), .A4(n5041), .ZN(n5043)
         );
  INV_X2 U5076 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U5077 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6519) );
  INV_X1 U5078 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6506) );
  BUF_X1 U5079 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n6791) );
  NOR2_X1 U5080 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5035) );
  INV_X1 U5081 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5238) );
  NOR2_X1 U5082 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6134) );
  INV_X1 U5083 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6002) );
  INV_X1 U5084 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5401) );
  INV_X1 U5085 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5092) );
  NOR2_X1 U5086 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5896) );
  INV_X2 U5087 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U5088 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4606) );
  OAI21_X2 U5089 ( .B1(n8134), .B2(n6300), .A(n6459), .ZN(n6313) );
  NOR2_X2 U5090 ( .A1(n4501), .A2(n5721), .ZN(n9087) );
  XNOR2_X2 U5091 ( .A(n5163), .B(n5162), .ZN(n9483) );
  AOI21_X2 U5092 ( .B1(n6105), .B2(n4515), .A(n4731), .ZN(n8901) );
  NAND2_X2 U5093 ( .A1(n4570), .A2(n7971), .ZN(n6105) );
  AND2_X4 U5094 ( .A1(n5114), .A2(n5817), .ZN(n5145) );
  NOR2_X4 U5095 ( .A1(n6029), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5900) );
  OAI21_X2 U5096 ( .B1(n8494), .B2(n8493), .A(n6455), .ZN(n8134) );
  OR3_X4 U5097 ( .A1(n7917), .A2(n7922), .A3(n5821), .ZN(n6710) );
  OAI222_X1 U5098 ( .A1(n4480), .A2(n7804), .B1(P1_U3084), .B2(n5821), .C1(
        n7776), .C2(n9896), .ZN(P1_U3329) );
  XNOR2_X2 U5099 ( .A(n5072), .B(n5071), .ZN(n5821) );
  INV_X2 U5100 ( .A(n5203), .ZN(n5856) );
  OR2_X1 U5101 ( .A1(n8966), .A2(n8789), .ZN(n8128) );
  OR2_X1 U5102 ( .A1(n8977), .A2(n8547), .ZN(n6435) );
  INV_X1 U5103 ( .A(n9903), .ZN(n5083) );
  AND2_X1 U5104 ( .A1(n5524), .A2(n5504), .ZN(n5522) );
  NAND2_X1 U5105 ( .A1(n5497), .A2(n5474), .ZN(n5498) );
  AND2_X1 U5106 ( .A1(n5086), .A2(n5083), .ZN(n5203) );
  NAND2_X1 U5107 ( .A1(n4989), .A2(n4987), .ZN(n9570) );
  NAND2_X1 U5108 ( .A1(n4988), .A2(n4525), .ZN(n4987) );
  NAND2_X1 U5109 ( .A1(n9296), .A2(n7402), .ZN(n9217) );
  AOI21_X1 U5110 ( .B1(n4845), .B2(n4847), .A(n4567), .ZN(n4843) );
  INV_X2 U5111 ( .A(n6649), .ZN(n6660) );
  NAND2_X1 U5112 ( .A1(n4632), .A2(n6467), .ZN(n4631) );
  INV_X1 U5113 ( .A(n6469), .ZN(n4632) );
  OR2_X1 U5114 ( .A1(n8716), .A2(n8495), .ZN(n6459) );
  OR2_X1 U5115 ( .A1(n8946), .A2(n8130), .ZN(n6450) );
  NAND2_X1 U5116 ( .A1(n8946), .A2(n8130), .ZN(n6455) );
  OR2_X1 U5117 ( .A1(n6252), .A2(n8627), .ZN(n6264) );
  OR2_X1 U5118 ( .A1(n9005), .A2(n8869), .ZN(n8864) );
  OR2_X1 U5119 ( .A1(n9972), .A2(n10386), .ZN(n4744) );
  NAND2_X1 U5120 ( .A1(n4935), .A2(n4483), .ZN(n4934) );
  AND2_X1 U5121 ( .A1(n4715), .A2(n7887), .ZN(n4712) );
  OR2_X1 U5122 ( .A1(n10386), .A2(n7976), .ZN(n6393) );
  NOR2_X1 U5123 ( .A1(n6020), .A2(n4727), .ZN(n4726) );
  INV_X1 U5124 ( .A(n6368), .ZN(n4727) );
  NAND2_X1 U5125 ( .A1(n4894), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6001) );
  OR2_X1 U5126 ( .A1(n4584), .A2(n9005), .ZN(n4747) );
  INV_X1 U5127 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U5128 ( .A1(n9131), .A2(n9133), .ZN(n4648) );
  NAND2_X1 U5129 ( .A1(n7247), .A2(n7248), .ZN(n5285) );
  OR2_X1 U5130 ( .A1(n9591), .A2(n5302), .ZN(n5764) );
  OR2_X1 U5131 ( .A1(n9786), .A2(n9556), .ZN(n9313) );
  OR2_X1 U5132 ( .A1(n9796), .A2(n9557), .ZN(n9423) );
  OR2_X1 U5133 ( .A1(n9802), .A2(n9611), .ZN(n9419) );
  AND2_X1 U5134 ( .A1(n9811), .A2(n9642), .ZN(n9251) );
  INV_X1 U5135 ( .A(n4970), .ZN(n4968) );
  OR2_X1 U5136 ( .A1(n9841), .A2(n9846), .ZN(n4692) );
  OR2_X1 U5137 ( .A1(n9948), .A2(n7816), .ZN(n9351) );
  NOR3_X1 U5138 ( .A1(n9740), .A2(n9833), .A3(n4691), .ZN(n9683) );
  NAND2_X1 U5139 ( .A1(n4871), .A2(n4870), .ZN(n5748) );
  AOI21_X1 U5140 ( .B1(n4496), .B2(n4876), .A(n4560), .ZN(n4870) );
  NAND2_X1 U5141 ( .A1(n5525), .A2(n5524), .ZN(n5547) );
  NAND2_X1 U5142 ( .A1(n4851), .A2(n4849), .ZN(n5525) );
  AOI21_X1 U5143 ( .B1(n4852), .B2(n4499), .A(n4850), .ZN(n4849) );
  AOI21_X1 U5144 ( .B1(n4867), .B2(n4865), .A(n4540), .ZN(n4864) );
  NAND2_X1 U5145 ( .A1(n5421), .A2(n5399), .ZN(n5422) );
  OR2_X1 U5146 ( .A1(n6192), .A2(n8594), .ZN(n6201) );
  AOI21_X1 U5147 ( .B1(n4807), .B2(n4811), .A(n4805), .ZN(n4804) );
  INV_X1 U5148 ( .A(n7702), .ZN(n4805) );
  INV_X1 U5149 ( .A(n4807), .ZN(n4806) );
  INV_X1 U5150 ( .A(n6312), .ZN(n6294) );
  NAND2_X1 U5152 ( .A1(n8487), .A2(n9049), .ZN(n5954) );
  OAI21_X1 U5153 ( .B1(n6082), .B2(n5889), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6164) );
  AOI21_X1 U5154 ( .B1(n4920), .B2(n4923), .A(n4532), .ZN(n4918) );
  AOI21_X1 U5155 ( .B1(n4907), .B2(n4906), .A(n4524), .ZN(n4905) );
  INV_X1 U5156 ( .A(n8811), .ZN(n4906) );
  NAND2_X1 U5157 ( .A1(n8128), .A2(n6238), .ZN(n8771) );
  NAND2_X1 U5158 ( .A1(n8801), .A2(n8811), .ZN(n4908) );
  AOI21_X1 U5159 ( .B1(n8865), .B2(n4910), .A(n8120), .ZN(n4909) );
  INV_X1 U5160 ( .A(n8118), .ZN(n4910) );
  NOR2_X1 U5161 ( .A1(n7971), .A2(n4897), .ZN(n4896) );
  INV_X1 U5162 ( .A(n7969), .ZN(n4897) );
  INV_X1 U5163 ( .A(n6088), .ZN(n6087) );
  NOR2_X1 U5164 ( .A1(n7572), .A2(n4900), .ZN(n4899) );
  INV_X1 U5165 ( .A(n7566), .ZN(n4900) );
  INV_X1 U5166 ( .A(n6832), .ZN(n6175) );
  NAND2_X1 U5167 ( .A1(n4543), .A2(n4574), .ZN(n7561) );
  INV_X1 U5168 ( .A(n7289), .ZN(n4574) );
  NAND2_X1 U5169 ( .A1(n4730), .A2(n6482), .ZN(n7274) );
  NAND2_X1 U5170 ( .A1(n7456), .A2(n6345), .ZN(n4730) );
  OR2_X1 U5171 ( .A1(n4478), .A2(n8328), .ZN(n5980) );
  NAND2_X1 U5172 ( .A1(n5140), .A2(n6724), .ZN(n5273) );
  NAND2_X1 U5174 ( .A1(n9169), .A2(n5368), .ZN(n4860) );
  NAND2_X1 U5175 ( .A1(n9553), .A2(n9552), .ZN(n9551) );
  NAND2_X1 U5176 ( .A1(n9802), .A2(n9611), .ZN(n9577) );
  OR2_X1 U5177 ( .A1(n9811), .A2(n9642), .ZN(n9250) );
  NAND2_X1 U5178 ( .A1(n9816), .A2(n9654), .ZN(n5001) );
  OR2_X1 U5179 ( .A1(n9816), .A2(n9654), .ZN(n8069) );
  AND2_X1 U5180 ( .A1(n9841), .A2(n9731), .ZN(n4974) );
  OR2_X1 U5181 ( .A1(n9853), .A2(n9770), .ZN(n9378) );
  NAND2_X1 U5182 ( .A1(n5007), .A2(n5005), .ZN(n9722) );
  NAND2_X1 U5183 ( .A1(n5006), .A2(n5016), .ZN(n5005) );
  INV_X1 U5184 ( .A(n5008), .ZN(n5006) );
  AND4_X1 U5185 ( .A1(n5487), .A2(n5486), .A3(n5485), .A4(n5484), .ZN(n9750)
         );
  AND2_X1 U5186 ( .A1(n5009), .A2(n5012), .ZN(n5008) );
  NAND2_X1 U5187 ( .A1(n7960), .A2(n9273), .ZN(n4770) );
  INV_X1 U5188 ( .A(n9173), .ZN(n5579) );
  AOI21_X1 U5189 ( .B1(n5079), .B2(n4962), .A(n4965), .ZN(n4964) );
  NOR2_X1 U5190 ( .A1(n9895), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n4962) );
  AND2_X1 U5191 ( .A1(n5699), .A2(n5679), .ZN(n5697) );
  NAND2_X1 U5192 ( .A1(n4848), .A2(n4852), .ZN(n5523) );
  OR2_X1 U5193 ( .A1(n5448), .A2(n4499), .ZN(n4848) );
  INV_X1 U5194 ( .A(n6777), .ZN(n6713) );
  NAND2_X1 U5195 ( .A1(n9787), .A2(n9735), .ZN(n4772) );
  NAND2_X1 U5196 ( .A1(n4578), .A2(n4577), .ZN(n9350) );
  NAND2_X1 U5197 ( .A1(n9341), .A2(n9406), .ZN(n4577) );
  INV_X1 U5198 ( .A(n4895), .ZN(n6346) );
  NAND2_X1 U5199 ( .A1(n4622), .A2(n4621), .ZN(n4620) );
  AND2_X1 U5200 ( .A1(n6388), .A2(n6382), .ZN(n4621) );
  NAND2_X1 U5201 ( .A1(n6386), .A2(n4623), .ZN(n4622) );
  NOR2_X1 U5202 ( .A1(n4624), .A2(n4717), .ZN(n4623) );
  NAND2_X1 U5203 ( .A1(n6415), .A2(n6414), .ZN(n4615) );
  INV_X1 U5204 ( .A(n9408), .ZN(n4576) );
  AND2_X1 U5205 ( .A1(n9661), .A2(n9399), .ZN(n4591) );
  OAI21_X1 U5206 ( .B1(n4610), .B2(n4609), .A(n6448), .ZN(n4608) );
  NAND2_X1 U5207 ( .A1(n6446), .A2(n8756), .ZN(n4609) );
  NOR2_X1 U5208 ( .A1(n4612), .A2(n4611), .ZN(n4610) );
  NOR2_X1 U5209 ( .A1(n6447), .A2(n8733), .ZN(n4607) );
  NOR2_X1 U5210 ( .A1(n9346), .A2(n4800), .ZN(n4799) );
  INV_X1 U5211 ( .A(n9343), .ZN(n4800) );
  NAND2_X1 U5212 ( .A1(n4841), .A2(n5570), .ZN(n4840) );
  NAND2_X1 U5213 ( .A1(n5546), .A2(n5545), .ZN(n4841) );
  NAND2_X1 U5214 ( .A1(n5341), .A2(n5028), .ZN(n5343) );
  NAND2_X1 U5215 ( .A1(n5320), .A2(n5319), .ZN(n5342) );
  NOR2_X1 U5216 ( .A1(P1_RD_REG_SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n5052) );
  NAND2_X1 U5217 ( .A1(n4887), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4893) );
  INV_X1 U5218 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4887) );
  NOR2_X1 U5219 ( .A1(n8957), .A2(n8557), .ZN(n6473) );
  AND2_X1 U5220 ( .A1(n8957), .A2(n8557), .ZN(n6472) );
  INV_X1 U5221 ( .A(n4722), .ZN(n4721) );
  AND2_X1 U5222 ( .A1(n4719), .A2(n6218), .ZN(n4718) );
  AND2_X1 U5223 ( .A1(n6206), .A2(n6423), .ZN(n4722) );
  OR2_X1 U5224 ( .A1(n8982), .A2(n8812), .ZN(n6429) );
  OR2_X1 U5225 ( .A1(n8994), .A2(n4747), .ZN(n4746) );
  NAND2_X1 U5226 ( .A1(n8891), .A2(n4915), .ZN(n4914) );
  INV_X1 U5227 ( .A(n4916), .ZN(n4915) );
  AOI21_X1 U5228 ( .B1(n4934), .B2(n8117), .A(n8927), .ZN(n4932) );
  INV_X1 U5229 ( .A(n8117), .ZN(n4930) );
  INV_X1 U5230 ( .A(n6121), .ZN(n4733) );
  OR2_X1 U5231 ( .A1(n8701), .A2(n7661), .ZN(n7089) );
  OR2_X1 U5232 ( .A1(n8972), .A2(n8977), .ZN(n4749) );
  AND2_X1 U5233 ( .A1(n7720), .A2(n10372), .ZN(n7762) );
  CLKBUF_X1 U5234 ( .A(n5900), .Z(n6035) );
  NAND2_X1 U5235 ( .A1(n5695), .A2(n9070), .ZN(n4642) );
  XNOR2_X1 U5236 ( .A(n5814), .B(n4671), .ZN(n5122) );
  NOR2_X1 U5237 ( .A1(n7828), .A2(n4668), .ZN(n4667) );
  INV_X1 U5238 ( .A(n5420), .ZN(n4668) );
  NOR2_X1 U5239 ( .A1(n9251), .A2(n5000), .ZN(n4999) );
  INV_X1 U5240 ( .A(n5001), .ZN(n5000) );
  NAND2_X1 U5241 ( .A1(n9635), .A2(n4685), .ZN(n4684) );
  OR2_X1 U5242 ( .A1(n9827), .A2(n9682), .ZN(n9399) );
  AND2_X1 U5243 ( .A1(n9689), .A2(n9701), .ZN(n9398) );
  NAND2_X1 U5244 ( .A1(n4762), .A2(n9253), .ZN(n4761) );
  INV_X1 U5245 ( .A(n4763), .ZN(n4762) );
  NOR2_X1 U5246 ( .A1(n8065), .A2(n5019), .ZN(n5015) );
  NAND2_X1 U5247 ( .A1(n4769), .A2(n4767), .ZN(n4766) );
  AND2_X1 U5248 ( .A1(n9275), .A2(n4530), .ZN(n4769) );
  OR2_X1 U5249 ( .A1(n9864), .A2(n9162), .ZN(n9761) );
  NOR2_X1 U5250 ( .A1(n7895), .A2(n9996), .ZN(n4678) );
  NAND2_X1 U5251 ( .A1(n9932), .A2(n4799), .ZN(n4798) );
  INV_X1 U5252 ( .A(n7779), .ZN(n5004) );
  OR2_X1 U5253 ( .A1(n9217), .A2(n4777), .ZN(n4782) );
  INV_X1 U5254 ( .A(n9218), .ZN(n4777) );
  NOR2_X1 U5255 ( .A1(n7404), .A2(n4783), .ZN(n4780) );
  NAND2_X1 U5256 ( .A1(n9302), .A2(n9258), .ZN(n7364) );
  NOR2_X1 U5257 ( .A1(n4764), .A2(n9255), .ZN(n4763) );
  INV_X1 U5258 ( .A(n9378), .ZN(n4764) );
  XNOR2_X1 U5259 ( .A(n7152), .B(n10185), .ZN(n9261) );
  NAND2_X1 U5260 ( .A1(n9261), .A2(n7154), .ZN(n7209) );
  OR2_X1 U5261 ( .A1(n6317), .A2(n6316), .ZN(n6321) );
  OR2_X1 U5262 ( .A1(n6319), .A2(n6318), .ZN(n6320) );
  XNOR2_X1 U5263 ( .A(n6319), .B(n6318), .ZN(n6317) );
  AND2_X1 U5264 ( .A1(n5777), .A2(n5752), .ZN(n5775) );
  NAND2_X1 U5265 ( .A1(n5623), .A2(n5622), .ZN(n4837) );
  NOR2_X1 U5266 ( .A1(n5469), .A2(n4857), .ZN(n4856) );
  INV_X1 U5267 ( .A(n5447), .ZN(n4857) );
  INV_X1 U5268 ( .A(n5465), .ZN(n5469) );
  XNOR2_X1 U5269 ( .A(n5466), .B(SI_14_), .ZN(n5465) );
  NAND2_X1 U5270 ( .A1(n5424), .A2(n8331), .ZN(n5447) );
  NAND2_X1 U5271 ( .A1(n5446), .A2(n5031), .ZN(n5448) );
  XNOR2_X1 U5272 ( .A(n5392), .B(SI_11_), .ZN(n5391) );
  NAND2_X1 U5273 ( .A1(n5345), .A2(n5344), .ZN(n5367) );
  NAND2_X1 U5274 ( .A1(n5343), .A2(n5342), .ZN(n5366) );
  XNOR2_X1 U5275 ( .A(n5289), .B(SI_7_), .ZN(n5286) );
  NAND2_X1 U5276 ( .A1(n5272), .A2(n5271), .ZN(n5288) );
  NOR2_X1 U5277 ( .A1(n6616), .A2(n8611), .ZN(n5033) );
  NAND2_X1 U5278 ( .A1(n7443), .A2(n6574), .ZN(n7586) );
  NAND2_X1 U5279 ( .A1(n6229), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6242) );
  INV_X1 U5280 ( .A(n7926), .ZN(n4829) );
  OR2_X1 U5281 ( .A1(n6608), .A2(n4828), .ZN(n4827) );
  INV_X1 U5282 ( .A(n6601), .ZN(n4828) );
  NAND2_X1 U5283 ( .A1(n7839), .A2(n7838), .ZN(n6595) );
  NAND2_X1 U5284 ( .A1(n6638), .A2(n6637), .ZN(n8581) );
  INV_X1 U5285 ( .A(n4823), .ZN(n4822) );
  OAI21_X1 U5286 ( .B1(n5033), .B2(n6617), .A(n4824), .ZN(n4823) );
  INV_X1 U5287 ( .A(n8527), .ZN(n4824) );
  AND2_X1 U5288 ( .A1(n4808), .A2(n4549), .ZN(n4807) );
  OR2_X1 U5289 ( .A1(n4809), .A2(n7662), .ZN(n4808) );
  INV_X1 U5290 ( .A(n7584), .ZN(n4812) );
  CLKBUF_X1 U5291 ( .A(n7586), .Z(n4583) );
  XNOR2_X1 U5292 ( .A(n8998), .B(n6660), .ZN(n6615) );
  AOI21_X1 U5293 ( .B1(n4493), .B2(n4631), .A(n4629), .ZN(n4628) );
  OR2_X1 U5294 ( .A1(n6466), .A2(n4630), .ZN(n4627) );
  INV_X1 U5295 ( .A(n4631), .ZN(n4630) );
  AND2_X1 U5296 ( .A1(n6285), .A2(n6284), .ZN(n8130) );
  AND2_X1 U5297 ( .A1(n6272), .A2(n6271), .ZN(n8626) );
  AND4_X1 U5298 ( .A1(n6133), .A2(n6132), .A3(n6131), .A4(n6130), .ZN(n8576)
         );
  AND4_X1 U5299 ( .A1(n6062), .A2(n6061), .A3(n6060), .A4(n6059), .ZN(n7754)
         );
  AND2_X1 U5300 ( .A1(n4696), .A2(n4695), .ZN(n9918) );
  OR2_X1 U5301 ( .A1(n6854), .A2(n6853), .ZN(n4703) );
  NAND2_X1 U5302 ( .A1(n4587), .A2(n4586), .ZN(n7118) );
  INV_X1 U5303 ( .A(n7065), .ZN(n4586) );
  NAND2_X1 U5304 ( .A1(n7867), .A2(n6128), .ZN(n8002) );
  OR2_X1 U5305 ( .A1(n8005), .A2(n8004), .ZN(n4699) );
  AND2_X1 U5306 ( .A1(n6459), .A2(n6460), .ZN(n8133) );
  NAND2_X1 U5307 ( .A1(n6450), .A2(n6455), .ZN(n8493) );
  NOR2_X1 U5308 ( .A1(n8747), .A2(n8756), .ZN(n4924) );
  AND2_X1 U5309 ( .A1(n6264), .A2(n6253), .ZN(n8743) );
  NOR2_X1 U5310 ( .A1(n6473), .A2(n6472), .ZN(n8747) );
  NOR2_X1 U5311 ( .A1(n4903), .A2(n8771), .ZN(n4902) );
  INV_X1 U5312 ( .A(n4905), .ZN(n4903) );
  NAND2_X1 U5313 ( .A1(n8823), .A2(n8812), .ZN(n4573) );
  NAND2_X1 U5314 ( .A1(n6435), .A2(n6434), .ZN(n8811) );
  NAND2_X1 U5315 ( .A1(n8836), .A2(n6197), .ZN(n4723) );
  NAND2_X1 U5316 ( .A1(n4723), .A2(n4722), .ZN(n8825) );
  OR2_X1 U5317 ( .A1(n6145), .A2(n6144), .ZN(n6157) );
  OR2_X1 U5318 ( .A1(n9015), .A2(n4914), .ZN(n8890) );
  AND4_X1 U5319 ( .A1(n6150), .A2(n6149), .A3(n6148), .A4(n6147), .ZN(n8885)
         );
  AND2_X1 U5320 ( .A1(n6407), .A2(n6406), .ZN(n8927) );
  NAND2_X1 U5321 ( .A1(n6105), .A2(n4504), .ZN(n9968) );
  OR2_X1 U5322 ( .A1(n4936), .A2(n4934), .ZN(n4933) );
  INV_X1 U5323 ( .A(n6391), .ZN(n4716) );
  OR2_X1 U5324 ( .A1(n7713), .A2(n7757), .ZN(n4713) );
  NAND2_X1 U5325 ( .A1(n7713), .A2(n7750), .ZN(n4714) );
  AND2_X1 U5326 ( .A1(n6382), .A2(n7750), .ZN(n7755) );
  AND4_X1 U5327 ( .A1(n6015), .A2(n6014), .A3(n6013), .A4(n6012), .ZN(n7573)
         );
  AND2_X1 U5328 ( .A1(n6370), .A2(n6371), .ZN(n7641) );
  NAND2_X1 U5329 ( .A1(n7274), .A2(n7292), .ZN(n6007) );
  OR2_X1 U5330 ( .A1(n4478), .A2(n8332), .ZN(n5964) );
  NAND2_X1 U5331 ( .A1(n8650), .A2(n8107), .ZN(n7300) );
  NAND2_X1 U5332 ( .A1(n6277), .A2(n6276), .ZN(n8946) );
  OR2_X1 U5333 ( .A1(n4478), .A2(n8013), .ZN(n6276) );
  NAND2_X1 U5334 ( .A1(n6261), .A2(n6260), .ZN(n8951) );
  OR2_X1 U5335 ( .A1(n4478), .A2(n7990), .ZN(n6260) );
  OR2_X1 U5336 ( .A1(n4478), .A2(n6721), .ZN(n5993) );
  AND2_X1 U5337 ( .A1(n5899), .A2(n5900), .ZN(n5903) );
  NAND2_X1 U5338 ( .A1(n4830), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U5339 ( .A1(n6164), .A2(n5890), .ZN(n4830) );
  NAND2_X1 U5340 ( .A1(n4606), .A2(n9910), .ZN(n5939) );
  AOI21_X1 U5341 ( .B1(n5567), .B2(n4940), .A(n4939), .ZN(n4938) );
  INV_X1 U5342 ( .A(n8047), .ZN(n4939) );
  NOR2_X1 U5343 ( .A1(n4955), .A2(n4522), .ZN(n4951) );
  OR2_X1 U5344 ( .A1(n5875), .A2(n5874), .ZN(n4955) );
  INV_X1 U5345 ( .A(n9086), .ZN(n4952) );
  NAND2_X1 U5346 ( .A1(n7649), .A2(n7648), .ZN(n4958) );
  NAND2_X1 U5347 ( .A1(n4484), .A2(n5695), .ZN(n4646) );
  AOI21_X1 U5348 ( .B1(n4648), .B2(n4484), .A(n5695), .ZN(n9113) );
  OR2_X1 U5349 ( .A1(n4641), .A2(n5671), .ZN(n4636) );
  INV_X1 U5350 ( .A(n4642), .ZN(n4641) );
  AND2_X1 U5351 ( .A1(n4644), .A2(n4640), .ZN(n4639) );
  NAND2_X1 U5352 ( .A1(n5696), .A2(n4645), .ZN(n4640) );
  INV_X1 U5353 ( .A(n9112), .ZN(n4644) );
  AND2_X1 U5354 ( .A1(n4642), .A2(n9133), .ZN(n4638) );
  INV_X1 U5355 ( .A(n5365), .ZN(n4661) );
  AND2_X1 U5356 ( .A1(n4663), .A2(n5340), .ZN(n4662) );
  NAND2_X1 U5357 ( .A1(n7697), .A2(n4943), .ZN(n4663) );
  NOR2_X1 U5358 ( .A1(n5365), .A2(n7697), .ZN(n4659) );
  NOR2_X1 U5359 ( .A1(n4949), .A2(n4946), .ZN(n4945) );
  NOR2_X1 U5360 ( .A1(n7421), .A2(n5314), .ZN(n4949) );
  INV_X1 U5361 ( .A(n7249), .ZN(n4946) );
  NAND2_X1 U5362 ( .A1(n5144), .A2(n4957), .ZN(n4956) );
  NAND2_X1 U5363 ( .A1(n7210), .A2(n5817), .ZN(n4957) );
  NOR2_X1 U5364 ( .A1(n5567), .A2(n4940), .ZN(n4941) );
  OR2_X1 U5365 ( .A1(n9102), .A2(n9105), .ZN(n9103) );
  AND4_X1 U5366 ( .A1(n5742), .A2(n5741), .A3(n5740), .A4(n5739), .ZN(n9469)
         );
  INV_X1 U5367 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n4961) );
  NAND2_X1 U5368 ( .A1(n4960), .A2(n4675), .ZN(n5049) );
  NOR2_X1 U5369 ( .A1(n4482), .A2(n5020), .ZN(n4675) );
  NAND2_X1 U5370 ( .A1(n4539), .A2(n5048), .ZN(n5020) );
  NOR2_X1 U5371 ( .A1(n9993), .A2(n4689), .ZN(n4687) );
  NAND2_X1 U5372 ( .A1(n4789), .A2(n4790), .ZN(n9555) );
  NOR2_X1 U5373 ( .A1(n9802), .A2(n9601), .ZN(n9587) );
  AND2_X1 U5374 ( .A1(n9419), .A2(n9577), .ZN(n9594) );
  NAND2_X1 U5375 ( .A1(n4509), .A2(n4996), .ZN(n4995) );
  INV_X1 U5376 ( .A(n9609), .ZN(n4996) );
  AND2_X1 U5377 ( .A1(n4509), .A2(n9250), .ZN(n4997) );
  AND4_X1 U5378 ( .A1(n5762), .A2(n5761), .A3(n5760), .A4(n5759), .ZN(n9611)
         );
  NAND2_X1 U5379 ( .A1(n4756), .A2(n4531), .ZN(n4755) );
  INV_X1 U5380 ( .A(n9808), .ZN(n9603) );
  OR2_X1 U5381 ( .A1(n9252), .A2(n9251), .ZN(n9624) );
  NAND2_X1 U5382 ( .A1(n9683), .A2(n8075), .ZN(n9668) );
  NAND2_X1 U5383 ( .A1(n4541), .A2(n4488), .ZN(n4970) );
  NAND2_X1 U5384 ( .A1(n9765), .A2(n9373), .ZN(n9748) );
  INV_X1 U5385 ( .A(n5013), .ZN(n5012) );
  OAI21_X1 U5386 ( .B1(n8065), .B2(n5014), .A(n5017), .ZN(n5013) );
  NAND2_X1 U5387 ( .A1(n5018), .A2(n8063), .ZN(n5014) );
  NAND2_X1 U5388 ( .A1(n8064), .A2(n5015), .ZN(n5010) );
  AND4_X1 U5389 ( .A1(n5514), .A2(n5513), .A3(n5512), .A4(n5511), .ZN(n9770)
         );
  AND2_X1 U5390 ( .A1(n5480), .A2(n5479), .ZN(n9759) );
  NAND2_X1 U5391 ( .A1(n4770), .A2(n4769), .ZN(n9762) );
  INV_X1 U5392 ( .A(n4795), .ZN(n4794) );
  NAND2_X1 U5393 ( .A1(n7810), .A2(n7809), .ZN(n7898) );
  OR2_X1 U5394 ( .A1(n7617), .A2(n9266), .ZN(n7780) );
  OR2_X1 U5395 ( .A1(n7619), .A2(n9264), .ZN(n7621) );
  OR2_X1 U5396 ( .A1(n9473), .A2(n7526), .ZN(n9335) );
  AOI21_X1 U5397 ( .B1(n4984), .B2(n7408), .A(n4527), .ZN(n4982) );
  NAND2_X1 U5398 ( .A1(n7494), .A2(n7526), .ZN(n7627) );
  INV_X1 U5399 ( .A(n7407), .ZN(n4986) );
  NAND2_X1 U5400 ( .A1(n7364), .A2(n9218), .ZN(n7403) );
  INV_X1 U5401 ( .A(n9772), .ZN(n9940) );
  AND2_X1 U5402 ( .A1(n7159), .A2(n9446), .ZN(n9938) );
  NAND2_X1 U5403 ( .A1(n10185), .A2(n7314), .ZN(n7395) );
  NOR2_X1 U5404 ( .A1(n7153), .A2(n7314), .ZN(n7157) );
  INV_X1 U5405 ( .A(n9591), .ZN(n9802) );
  AND2_X1 U5406 ( .A1(n7312), .A2(n7164), .ZN(n9994) );
  XNOR2_X1 U5407 ( .A(n6302), .B(n6301), .ZN(n8485) );
  NAND2_X1 U5408 ( .A1(n4844), .A2(n6290), .ZN(n6302) );
  NAND2_X1 U5409 ( .A1(n6287), .A2(n6286), .ZN(n4844) );
  NAND2_X1 U5410 ( .A1(n5801), .A2(n5800), .ZN(n6287) );
  NAND2_X1 U5411 ( .A1(n5799), .A2(n5798), .ZN(n5801) );
  NAND2_X1 U5412 ( .A1(n4872), .A2(n4873), .ZN(n5725) );
  OR2_X1 U5413 ( .A1(n5675), .A2(n4876), .ZN(n4872) );
  NAND2_X1 U5414 ( .A1(n4505), .A2(n5043), .ZN(n5044) );
  INV_X1 U5415 ( .A(n7639), .ZN(n10351) );
  AND4_X1 U5416 ( .A1(n6028), .A2(n6027), .A3(n6026), .A4(n6025), .ZN(n7644)
         );
  AND2_X1 U5417 ( .A1(n6216), .A2(n6215), .ZN(n8547) );
  NAND2_X1 U5418 ( .A1(n6832), .A2(n4739), .ZN(n4740) );
  OAI22_X1 U5419 ( .A1(n6725), .A2(n6724), .B1(n6719), .B2(n5936), .ZN(n4739)
         );
  AND3_X1 U5420 ( .A1(n6196), .A2(n6195), .A3(n6194), .ZN(n8548) );
  OAI21_X1 U5421 ( .B1(n8610), .B2(n4818), .A(n4815), .ZN(n8545) );
  AOI21_X1 U5422 ( .B1(n4820), .B2(n4817), .A(n4816), .ZN(n4815) );
  NAND2_X1 U5423 ( .A1(n4820), .A2(n4819), .ZN(n4818) );
  NOR2_X1 U5424 ( .A1(n6627), .A2(n6626), .ZN(n4816) );
  AND4_X1 U5425 ( .A1(n6077), .A2(n6076), .A3(n6075), .A4(n6074), .ZN(n7889)
         );
  NAND2_X1 U5426 ( .A1(n6086), .A2(n6085), .ZN(n10386) );
  OR2_X1 U5427 ( .A1(n4478), .A2(n7915), .ZN(n6239) );
  AND2_X1 U5428 ( .A1(n7024), .A2(n6552), .ZN(n7102) );
  NAND2_X1 U5429 ( .A1(n7102), .A2(n7101), .ZN(n7100) );
  NAND2_X1 U5430 ( .A1(n6154), .A2(n6153), .ZN(n9005) );
  INV_X1 U5431 ( .A(n8650), .ZN(n8109) );
  OR2_X1 U5432 ( .A1(n4478), .A2(n7502), .ZN(n6188) );
  AND4_X1 U5433 ( .A1(n6093), .A2(n6092), .A3(n6091), .A4(n6090), .ZN(n7976)
         );
  OR2_X1 U5434 ( .A1(n6738), .A2(n5960), .ZN(n6006) );
  OR2_X1 U5435 ( .A1(n4478), .A2(n6737), .ZN(n6005) );
  INV_X1 U5436 ( .A(n8130), .ZN(n8735) );
  OR2_X1 U5437 ( .A1(n6896), .A2(n6895), .ZN(n4701) );
  AND2_X1 U5438 ( .A1(n4703), .A2(n4702), .ZN(n6896) );
  NAND2_X1 U5439 ( .A1(n6898), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4702) );
  NOR2_X1 U5440 ( .A1(n6971), .A2(n6970), .ZN(n7063) );
  NOR2_X1 U5441 ( .A1(n6967), .A2(n4707), .ZN(n6971) );
  AND2_X1 U5442 ( .A1(n6968), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4707) );
  INV_X1 U5443 ( .A(n8702), .ZN(n4580) );
  XNOR2_X1 U5444 ( .A(n5905), .B(n5904), .ZN(n8701) );
  NAND2_X1 U5445 ( .A1(n4655), .A2(n4652), .ZN(n4651) );
  NAND2_X1 U5446 ( .A1(n5875), .A2(n4653), .ZN(n4652) );
  NAND2_X1 U5447 ( .A1(n4951), .A2(n4656), .ZN(n4655) );
  NOR2_X1 U5448 ( .A1(n4654), .A2(n9139), .ZN(n4653) );
  AND2_X1 U5449 ( .A1(n4951), .A2(n9152), .ZN(n4657) );
  NAND2_X1 U5450 ( .A1(n7746), .A2(n5368), .ZN(n5681) );
  AND2_X1 U5451 ( .A1(n5841), .A2(n9152), .ZN(n5871) );
  NAND2_X1 U5452 ( .A1(n5508), .A2(n5507), .ZN(n9853) );
  NAND2_X1 U5453 ( .A1(n5553), .A2(n5552), .ZN(n9841) );
  NAND2_X1 U5454 ( .A1(n9450), .A2(n9671), .ZN(n4886) );
  AOI21_X1 U5455 ( .B1(n9457), .B2(n7467), .A(n9465), .ZN(n4882) );
  NAND4_X1 U5456 ( .A1(n5210), .A2(n5209), .A3(n5208), .A4(n5207), .ZN(n9475)
         );
  NOR2_X1 U5457 ( .A1(n4776), .A2(n9772), .ZN(n4775) );
  AND2_X1 U5458 ( .A1(n9434), .A2(n9552), .ZN(n4975) );
  NOR2_X1 U5459 ( .A1(n9434), .A2(n4550), .ZN(n4978) );
  NAND2_X1 U5460 ( .A1(n9434), .A2(n4550), .ZN(n4979) );
  OR2_X1 U5461 ( .A1(n4771), .A2(n8097), .ZN(n4774) );
  AND2_X1 U5462 ( .A1(n9774), .A2(n7313), .ZN(n9735) );
  NOR2_X1 U5463 ( .A1(n10461), .A2(n10460), .ZN(n10459) );
  NOR2_X1 U5464 ( .A1(n10455), .A2(n10454), .ZN(n10453) );
  NAND2_X1 U5465 ( .A1(n7364), .A2(n4785), .ZN(n4784) );
  INV_X1 U5466 ( .A(n4782), .ZN(n4785) );
  INV_X1 U5467 ( .A(n6384), .ZN(n4624) );
  OR2_X1 U5468 ( .A1(n6380), .A2(n4547), .ZN(n6386) );
  NAND2_X1 U5469 ( .A1(n4619), .A2(n4617), .ZN(n6399) );
  NAND2_X1 U5470 ( .A1(n6383), .A2(n4618), .ZN(n4617) );
  NOR2_X1 U5471 ( .A1(n4615), .A2(n4616), .ZN(n4614) );
  INV_X1 U5472 ( .A(n6411), .ZN(n4616) );
  NOR2_X1 U5473 ( .A1(n4576), .A2(n9406), .ZN(n4575) );
  INV_X1 U5474 ( .A(n6443), .ZN(n4612) );
  NAND2_X1 U5475 ( .A1(n6442), .A2(n8771), .ZN(n4611) );
  INV_X1 U5476 ( .A(n4846), .ZN(n4845) );
  OAI21_X1 U5477 ( .B1(n6286), .B2(n4847), .A(n6301), .ZN(n4846) );
  INV_X1 U5478 ( .A(n6290), .ZN(n4847) );
  NAND2_X1 U5479 ( .A1(n4722), .A2(n4720), .ZN(n4719) );
  INV_X1 U5480 ( .A(n6197), .ZN(n4720) );
  INV_X1 U5481 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5883) );
  OAI21_X1 U5482 ( .B1(n4995), .B2(n4994), .A(n4538), .ZN(n4993) );
  INV_X1 U5483 ( .A(n8071), .ZN(n4994) );
  AND2_X1 U5484 ( .A1(n4879), .A2(n5697), .ZN(n4878) );
  NAND2_X1 U5485 ( .A1(n5674), .A2(n5673), .ZN(n4879) );
  INV_X1 U5486 ( .A(n5522), .ZN(n4850) );
  NOR2_X1 U5487 ( .A1(n4866), .A2(n4863), .ZN(n4862) );
  INV_X1 U5488 ( .A(n5342), .ZN(n4863) );
  INV_X1 U5489 ( .A(n4867), .ZN(n4866) );
  NOR2_X1 U5490 ( .A1(n5394), .A2(n4868), .ZN(n4867) );
  INV_X1 U5491 ( .A(n5367), .ZN(n4868) );
  INV_X1 U5492 ( .A(n5391), .ZN(n5394) );
  INV_X1 U5493 ( .A(n5030), .ZN(n4865) );
  NAND2_X1 U5494 ( .A1(n5292), .A2(n5291), .ZN(n5317) );
  OR2_X1 U5495 ( .A1(n6615), .A2(n4595), .ZN(n6613) );
  INV_X1 U5496 ( .A(n6614), .ZN(n4595) );
  NAND2_X1 U5497 ( .A1(n4813), .A2(n7584), .ZN(n4809) );
  OR2_X1 U5498 ( .A1(n6530), .A2(n6570), .ZN(n6540) );
  AOI21_X1 U5499 ( .B1(n8584), .B2(n8512), .A(n8582), .ZN(n6645) );
  AOI21_X1 U5500 ( .B1(n8584), .B2(n6639), .A(n8581), .ZN(n6641) );
  NOR2_X1 U5501 ( .A1(n4832), .A2(n4831), .ZN(n6570) );
  NOR2_X1 U5502 ( .A1(n6468), .A2(n6330), .ZN(n6497) );
  AOI211_X1 U5503 ( .C1(n4608), .C2(n4607), .A(n6453), .B(n6454), .ZN(n6458)
         );
  NAND2_X1 U5504 ( .A1(n7865), .A2(n4585), .ZN(n8000) );
  OR2_X1 U5505 ( .A1(n7866), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4585) );
  AOI21_X1 U5506 ( .B1(n4922), .B2(n4921), .A(n6273), .ZN(n4920) );
  INV_X1 U5507 ( .A(n4924), .ZN(n4921) );
  OR2_X1 U5508 ( .A1(n6221), .A2(n8511), .ZN(n6230) );
  NAND2_X1 U5509 ( .A1(n4913), .A2(n8865), .ZN(n4912) );
  INV_X1 U5510 ( .A(n4914), .ZN(n4913) );
  NOR2_X1 U5511 ( .A1(n4584), .A2(n8119), .ZN(n8120) );
  NOR2_X1 U5512 ( .A1(n7881), .A2(n10386), .ZN(n4745) );
  NAND2_X1 U5513 ( .A1(n4742), .A2(n7283), .ZN(n4741) );
  NAND2_X1 U5514 ( .A1(n4895), .A2(n6368), .ZN(n7285) );
  NOR2_X1 U5515 ( .A1(n7185), .A2(n7262), .ZN(n4742) );
  INV_X1 U5516 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6503) );
  INV_X1 U5517 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4605) );
  INV_X1 U5518 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4603) );
  INV_X1 U5519 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4604) );
  AND2_X1 U5520 ( .A1(n5683), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5703) );
  AND2_X1 U5521 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n5658), .ZN(n5683) );
  OR2_X1 U5522 ( .A1(n5806), .A2(n10192), .ZN(n5087) );
  NAND2_X1 U5523 ( .A1(n10046), .A2(n4507), .ZN(n10064) );
  NAND2_X1 U5524 ( .A1(n4572), .A2(n4571), .ZN(n5348) );
  INV_X1 U5525 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4571) );
  INV_X1 U5526 ( .A(n5298), .ZN(n4572) );
  NAND2_X1 U5527 ( .A1(n4791), .A2(n9423), .ZN(n4790) );
  INV_X1 U5528 ( .A(n8092), .ZN(n4791) );
  NOR2_X1 U5529 ( .A1(n4993), .A2(n4991), .ZN(n4990) );
  INV_X1 U5530 ( .A(n4999), .ZN(n4991) );
  INV_X1 U5531 ( .A(n4993), .ZN(n4988) );
  AND2_X1 U5532 ( .A1(n5703), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5732) );
  OR2_X1 U5533 ( .A1(n9821), .A2(n8087), .ZN(n9404) );
  NOR2_X1 U5534 ( .A1(n5627), .A2(n9078), .ZN(n5658) );
  OR2_X1 U5535 ( .A1(n9836), .A2(n4692), .ZN(n4691) );
  NAND2_X1 U5536 ( .A1(n9853), .A2(n9730), .ZN(n5016) );
  NAND2_X1 U5537 ( .A1(n4795), .A2(n4793), .ZN(n4792) );
  INV_X1 U5538 ( .A(n4799), .ZN(n4793) );
  NOR2_X1 U5539 ( .A1(n4797), .A2(n4796), .ZN(n4795) );
  INV_X1 U5540 ( .A(n4516), .ZN(n4796) );
  OR2_X1 U5541 ( .A1(n9475), .A2(n10217), .ZN(n9296) );
  NAND2_X1 U5542 ( .A1(n4787), .A2(n9238), .ZN(n4786) );
  OR2_X1 U5543 ( .A1(n4790), .A2(n9427), .ZN(n4787) );
  AND2_X1 U5544 ( .A1(n4512), .A2(n9426), .ZN(n4788) );
  OR2_X1 U5545 ( .A1(n7627), .A2(n7778), .ZN(n7787) );
  NOR2_X1 U5546 ( .A1(n7395), .A2(n7210), .ZN(n7396) );
  NOR2_X1 U5547 ( .A1(n9895), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4965) );
  AOI21_X1 U5548 ( .B1(n4878), .B2(n4875), .A(n4874), .ZN(n4873) );
  INV_X1 U5549 ( .A(n5699), .ZN(n4874) );
  INV_X1 U5550 ( .A(n5673), .ZN(n4875) );
  INV_X1 U5551 ( .A(n4878), .ZN(n4876) );
  NOR2_X1 U5552 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5038) );
  INV_X1 U5553 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5037) );
  INV_X1 U5554 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5042) );
  AND2_X1 U5555 ( .A1(n5624), .A2(n5605), .ZN(n5622) );
  INV_X1 U5556 ( .A(n4839), .ZN(n4838) );
  OAI21_X1 U5557 ( .B1(n4840), .B2(n5545), .A(n5573), .ZN(n4839) );
  INV_X1 U5558 ( .A(n5542), .ZN(n5546) );
  INV_X1 U5559 ( .A(n5468), .ZN(n4854) );
  INV_X1 U5560 ( .A(n4853), .ZN(n4852) );
  OAI21_X1 U5561 ( .B1(n4856), .B2(n4499), .A(n5497), .ZN(n4853) );
  NAND2_X1 U5562 ( .A1(n5318), .A2(n5317), .ZN(n5341) );
  NAND2_X1 U5563 ( .A1(n4836), .A2(n4834), .ZN(n5318) );
  NOR2_X1 U5564 ( .A1(n5316), .A2(n4835), .ZN(n4834) );
  INV_X1 U5565 ( .A(n5290), .ZN(n4835) );
  OAI21_X1 U5566 ( .B1(n6724), .B2(P1_DATAO_REG_5__SCAN_IN), .A(n4596), .ZN(
        n5233) );
  NAND2_X1 U5567 ( .A1(n6724), .A2(n6735), .ZN(n4596) );
  OAI21_X1 U5568 ( .B1(n6724), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n5187), .ZN(
        n5213) );
  OR2_X1 U5569 ( .A1(n6723), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5187) );
  OAI21_X1 U5570 ( .B1(n5052), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n4888), .ZN(
        n5053) );
  NAND2_X1 U5571 ( .A1(n4893), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4888) );
  NAND2_X1 U5572 ( .A1(n6595), .A2(n4503), .ZN(n7923) );
  INV_X1 U5573 ( .A(n4566), .ZN(n4813) );
  AND2_X1 U5574 ( .A1(n8111), .A2(n6532), .ZN(n8535) );
  INV_X1 U5575 ( .A(n8592), .ZN(n4819) );
  NOR2_X1 U5576 ( .A1(n4822), .A2(n8592), .ZN(n4817) );
  NAND2_X1 U5577 ( .A1(n6241), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6252) );
  XNOR2_X1 U5578 ( .A(n8773), .B(n6649), .ZN(n8584) );
  INV_X1 U5579 ( .A(n6623), .ZN(n4821) );
  INV_X1 U5580 ( .A(n6201), .ZN(n6200) );
  AND2_X1 U5581 ( .A1(n6828), .A2(n6709), .ZN(n6701) );
  NAND2_X1 U5582 ( .A1(n7923), .A2(n6601), .ZN(n8566) );
  NOR2_X1 U5583 ( .A1(n8941), .A2(n8032), .ZN(n6468) );
  AND2_X1 U5584 ( .A1(n6469), .A2(n6461), .ZN(n6496) );
  NOR2_X1 U5585 ( .A1(n6471), .A2(n6691), .ZN(n4626) );
  OAI21_X1 U5586 ( .B1(n9909), .B2(P2_REG2_REG_1__SCAN_IN), .A(n6844), .ZN(
        n9906) );
  OR2_X1 U5587 ( .A1(n7242), .A2(n7241), .ZN(n7550) );
  OR2_X1 U5588 ( .A1(n7554), .A2(n7553), .ZN(n4706) );
  AND2_X1 U5589 ( .A1(n4706), .A2(n4705), .ZN(n7605) );
  NAND2_X1 U5590 ( .A1(n7603), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4705) );
  NAND2_X1 U5591 ( .A1(n7605), .A2(n7604), .ZN(n7733) );
  NAND2_X1 U5592 ( .A1(n7733), .A2(n4704), .ZN(n7735) );
  OR2_X1 U5593 ( .A1(n7734), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4704) );
  XNOR2_X1 U5594 ( .A(n8000), .B(n7993), .ZN(n7867) );
  AOI21_X1 U5595 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n8678), .A(n8672), .ZN(
        n8674) );
  NOR2_X1 U5596 ( .A1(n8708), .A2(n8709), .ZN(n8707) );
  AND2_X1 U5597 ( .A1(n8714), .A2(n6279), .ZN(n8490) );
  NOR2_X1 U5598 ( .A1(n8725), .A2(n8946), .ZN(n8489) );
  OR2_X1 U5599 ( .A1(n8741), .A2(n8951), .ZN(n8725) );
  NAND2_X1 U5600 ( .A1(n4598), .A2(n4597), .ZN(n8741) );
  NAND2_X1 U5601 ( .A1(n8785), .A2(n6226), .ZN(n8787) );
  AND2_X1 U5602 ( .A1(n8987), .A2(n8853), .ZN(n8123) );
  NOR3_X1 U5603 ( .A1(n8908), .A2(n8987), .A3(n4746), .ZN(n8832) );
  AND2_X1 U5604 ( .A1(n6422), .A2(n8837), .ZN(n8848) );
  NAND2_X1 U5605 ( .A1(n6179), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6192) );
  INV_X1 U5606 ( .A(n6181), .ZN(n6179) );
  OR2_X1 U5607 ( .A1(n6169), .A2(n6168), .ZN(n6181) );
  NAND2_X1 U5608 ( .A1(n6166), .A2(n6165), .ZN(n8998) );
  NAND2_X1 U5609 ( .A1(n6156), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6169) );
  INV_X1 U5610 ( .A(n6157), .ZN(n6156) );
  AOI21_X1 U5611 ( .B1(n4932), .B2(n4930), .A(n4536), .ZN(n4929) );
  NAND2_X1 U5612 ( .A1(n4732), .A2(n6407), .ZN(n4731) );
  NAND2_X1 U5613 ( .A1(n8927), .A2(n4733), .ZN(n4732) );
  NAND2_X1 U5614 ( .A1(n8901), .A2(n8905), .ZN(n8900) );
  NOR2_X1 U5615 ( .A1(n8114), .A2(n4556), .ZN(n9977) );
  NAND2_X1 U5616 ( .A1(n6112), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6145) );
  OR2_X1 U5617 ( .A1(n6099), .A2(n7607), .ZN(n6113) );
  NAND2_X1 U5618 ( .A1(n4709), .A2(n4711), .ZN(n7975) );
  AOI21_X1 U5619 ( .B1(n4712), .B2(n7757), .A(n4710), .ZN(n4709) );
  INV_X1 U5620 ( .A(n6393), .ZN(n4710) );
  INV_X1 U5621 ( .A(n6071), .ZN(n6069) );
  OR2_X1 U5622 ( .A1(n6056), .A2(n6055), .ZN(n6071) );
  NAND2_X1 U5623 ( .A1(n6021), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6040) );
  INV_X1 U5624 ( .A(n6023), .ZN(n6021) );
  NAND2_X1 U5625 ( .A1(n7676), .A2(n7675), .ZN(n7710) );
  AND2_X1 U5626 ( .A1(n6385), .A2(n6381), .ZN(n7680) );
  OR2_X1 U5627 ( .A1(n7635), .A2(n7672), .ZN(n7688) );
  AND2_X1 U5628 ( .A1(n7572), .A2(n6371), .ZN(n4724) );
  AND2_X1 U5629 ( .A1(n4725), .A2(n6371), .ZN(n7571) );
  NAND2_X1 U5630 ( .A1(n7636), .A2(n10351), .ZN(n7635) );
  NAND2_X1 U5631 ( .A1(n5995), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6010) );
  NOR2_X1 U5632 ( .A1(n4741), .A2(n10346), .ZN(n7636) );
  INV_X1 U5633 ( .A(n4741), .ZN(n7453) );
  NOR2_X1 U5634 ( .A1(n5982), .A2(n4729), .ZN(n4728) );
  INV_X1 U5635 ( .A(n6349), .ZN(n4729) );
  INV_X1 U5636 ( .A(n4742), .ZN(n7454) );
  NAND2_X1 U5637 ( .A1(n10334), .A2(n10338), .ZN(n7302) );
  OR2_X1 U5638 ( .A1(n10357), .A2(n6682), .ZN(n7097) );
  NOR2_X1 U5639 ( .A1(n8140), .A2(n10381), .ZN(n4736) );
  NAND2_X1 U5640 ( .A1(n8138), .A2(n8137), .ZN(n4737) );
  XNOR2_X1 U5641 ( .A(n8134), .B(n8133), .ZN(n8135) );
  OR2_X1 U5642 ( .A1(n4478), .A2(n8321), .ZN(n6250) );
  NOR2_X1 U5643 ( .A1(n8908), .A2(n4747), .ZN(n8846) );
  INV_X1 U5644 ( .A(n10391), .ZN(n9020) );
  AND2_X1 U5645 ( .A1(n6677), .A2(n6672), .ZN(n10295) );
  NOR2_X1 U5646 ( .A1(n4928), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4927) );
  NAND2_X1 U5647 ( .A1(n5909), .A2(n5928), .ZN(n4928) );
  CLKBUF_X1 U5648 ( .A(n5975), .Z(n5976) );
  INV_X1 U5649 ( .A(n5874), .ZN(n4654) );
  AND2_X1 U5650 ( .A1(n5771), .A2(n9152), .ZN(n4656) );
  AND2_X1 U5651 ( .A1(n5490), .A2(n7829), .ZN(n4665) );
  XNOR2_X1 U5652 ( .A(n5517), .B(n5814), .ZN(n9094) );
  NAND2_X1 U5653 ( .A1(n7009), .A2(n7010), .ZN(n5174) );
  INV_X1 U5654 ( .A(n7421), .ZN(n4948) );
  AND2_X1 U5655 ( .A1(n5582), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5608) );
  AND2_X1 U5656 ( .A1(n5592), .A2(n5593), .ZN(n8054) );
  NOR2_X1 U5657 ( .A1(n5377), .A2(n5376), .ZN(n5406) );
  NOR2_X1 U5658 ( .A1(n5555), .A2(n5554), .ZN(n5582) );
  NAND2_X1 U5659 ( .A1(n5226), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5259) );
  AND3_X1 U5660 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U5661 ( .A1(n5757), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5785) );
  AND3_X1 U5662 ( .A1(n5840), .A2(n7147), .A3(n7309), .ZN(n6960) );
  INV_X1 U5663 ( .A(n5145), .ZN(n5811) );
  NAND2_X1 U5664 ( .A1(n4860), .A2(n4858), .ZN(n9451) );
  NOR2_X1 U5665 ( .A1(n9247), .A2(n4859), .ZN(n4858) );
  INV_X1 U5666 ( .A(n9170), .ZN(n4859) );
  AND2_X1 U5667 ( .A1(n9489), .A2(n6812), .ZN(n10031) );
  NAND2_X1 U5668 ( .A1(n4599), .A2(n10063), .ZN(n10067) );
  INV_X1 U5669 ( .A(n10064), .ZN(n4599) );
  NOR2_X1 U5670 ( .A1(n9511), .A2(n10137), .ZN(n10150) );
  AOI21_X1 U5671 ( .B1(n10153), .B2(P1_REG2_REG_16__SCAN_IN), .A(n10148), .ZN(
        n10164) );
  AOI21_X1 U5672 ( .B1(n9523), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9522), .ZN(
        n9524) );
  AND4_X1 U5673 ( .A1(n5861), .A2(n5860), .A3(n5859), .A4(n5858), .ZN(n9556)
         );
  AND4_X1 U5674 ( .A1(n5792), .A2(n5791), .A3(n5790), .A4(n5789), .ZN(n9557)
         );
  NAND2_X1 U5675 ( .A1(n9423), .A2(n9237), .ZN(n9579) );
  NAND2_X1 U5676 ( .A1(n4755), .A2(n4491), .ZN(n8091) );
  AND2_X1 U5677 ( .A1(n5732), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5757) );
  INV_X1 U5678 ( .A(n4684), .ZN(n4683) );
  OR2_X1 U5679 ( .A1(n9816), .A2(n8089), .ZN(n9622) );
  NOR3_X1 U5680 ( .A1(n9668), .A2(n9811), .A3(n4684), .ZN(n9616) );
  NAND2_X1 U5681 ( .A1(n4756), .A2(n8090), .ZN(n9636) );
  NOR2_X1 U5682 ( .A1(n9668), .A2(n4684), .ZN(n9631) );
  NAND2_X1 U5683 ( .A1(n9399), .A2(n9401), .ZN(n9660) );
  NAND2_X1 U5684 ( .A1(n4973), .A2(n8067), .ZN(n4969) );
  AOI21_X1 U5685 ( .B1(n8067), .B2(n4968), .A(n4529), .ZN(n4967) );
  OR2_X1 U5686 ( .A1(n9833), .A2(n9701), .ZN(n8067) );
  AOI21_X1 U5687 ( .B1(n4487), .B2(n9254), .A(n4759), .ZN(n4758) );
  INV_X1 U5688 ( .A(n9180), .ZN(n4759) );
  NOR2_X1 U5689 ( .A1(n9740), .A2(n4691), .ZN(n9693) );
  NOR2_X1 U5690 ( .A1(n9740), .A2(n4692), .ZN(n9708) );
  AND2_X1 U5691 ( .A1(n5482), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5509) );
  OR2_X1 U5692 ( .A1(n9758), .A2(n9853), .ZN(n9740) );
  INV_X1 U5693 ( .A(n4769), .ZN(n4768) );
  AND2_X1 U5694 ( .A1(n4766), .A2(n8080), .ZN(n4765) );
  NOR2_X1 U5695 ( .A1(n5455), .A2(n5454), .ZN(n5482) );
  AND2_X1 U5696 ( .A1(n9949), .A2(n4676), .ZN(n9760) );
  AND2_X1 U5697 ( .A1(n9067), .A2(n4497), .ZN(n4676) );
  NAND2_X1 U5698 ( .A1(n9949), .A2(n4678), .ZN(n7944) );
  NAND2_X1 U5699 ( .A1(n9949), .A2(n10003), .ZN(n7905) );
  NAND2_X1 U5700 ( .A1(n4798), .A2(n4795), .ZN(n7938) );
  NAND2_X1 U5701 ( .A1(n4798), .A2(n9181), .ZN(n7813) );
  AND2_X1 U5702 ( .A1(n9952), .A2(n9959), .ZN(n9949) );
  NOR2_X1 U5703 ( .A1(n7787), .A2(n10236), .ZN(n9952) );
  AOI21_X1 U5704 ( .B1(n4485), .B2(n9266), .A(n4534), .ZN(n5002) );
  OR2_X1 U5705 ( .A1(n5327), .A2(n5326), .ZN(n5352) );
  NAND2_X1 U5706 ( .A1(n9932), .A2(n9343), .ZN(n7811) );
  NOR2_X1 U5707 ( .A1(n5259), .A2(n5258), .ZN(n5303) );
  NOR2_X1 U5708 ( .A1(n7493), .A2(n7498), .ZN(n7494) );
  OAI21_X1 U5709 ( .B1(n7364), .B2(n4779), .A(n4778), .ZN(n7405) );
  NAND2_X1 U5710 ( .A1(n4680), .A2(n10217), .ZN(n7493) );
  INV_X1 U5711 ( .A(n9259), .ZN(n7217) );
  OR2_X1 U5712 ( .A1(n9173), .A2(n6726), .ZN(n5062) );
  AND2_X1 U5713 ( .A1(n9565), .A2(n9564), .ZN(n9792) );
  NAND2_X1 U5714 ( .A1(n4760), .A2(n9253), .ZN(n9713) );
  NAND2_X1 U5715 ( .A1(n8082), .A2(n4763), .ZN(n4760) );
  AND2_X1 U5716 ( .A1(n5301), .A2(n5300), .ZN(n10229) );
  AND2_X1 U5717 ( .A1(n5275), .A2(n5274), .ZN(n7526) );
  AND3_X1 U5718 ( .A1(n5243), .A2(n5242), .A3(n5241), .ZN(n10222) );
  XNOR2_X1 U5719 ( .A(n6324), .B(n6323), .ZN(n9169) );
  XNOR2_X1 U5720 ( .A(n6317), .B(SI_30_), .ZN(n9171) );
  INV_X1 U5721 ( .A(n5049), .ZN(n5078) );
  NAND2_X1 U5722 ( .A1(n5778), .A2(n5777), .ZN(n5799) );
  INV_X1 U5723 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5075) );
  NAND2_X1 U5724 ( .A1(n4855), .A2(n5468), .ZN(n5499) );
  NAND2_X1 U5725 ( .A1(n5448), .A2(n4856), .ZN(n4855) );
  NAND2_X1 U5726 ( .A1(n5448), .A2(n5447), .ZN(n5470) );
  NAND2_X1 U5727 ( .A1(n5366), .A2(n5030), .ZN(n4869) );
  INV_X1 U5728 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5296) );
  INV_X1 U5729 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4673) );
  INV_X1 U5730 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4674) );
  XNOR2_X1 U5731 ( .A(n5269), .B(SI_6_), .ZN(n5267) );
  XNOR2_X1 U5732 ( .A(n5233), .B(SI_5_), .ZN(n5231) );
  INV_X1 U5733 ( .A(n5057), .ZN(n6723) );
  AOI21_X1 U5734 ( .B1(n8743), .B2(n5969), .A(n6258), .ZN(n8557) );
  NAND2_X1 U5735 ( .A1(n6595), .A2(n6594), .ZN(n7925) );
  OR2_X1 U5736 ( .A1(n4478), .A2(n7749), .ZN(n6219) );
  OAI21_X1 U5737 ( .B1(n4583), .B2(n4813), .A(n7584), .ZN(n7663) );
  AND2_X1 U5738 ( .A1(n7020), .A2(n6547), .ZN(n8519) );
  OAI21_X1 U5739 ( .B1(n8610), .B2(n5033), .A(n4822), .ZN(n8525) );
  AOI21_X1 U5740 ( .B1(n8610), .B2(n6617), .A(n5033), .ZN(n8528) );
  AND4_X1 U5741 ( .A1(n6045), .A2(n6044), .A3(n6043), .A4(n6042), .ZN(n7664)
         );
  OR2_X1 U5742 ( .A1(n4478), .A2(n7595), .ZN(n6198) );
  AOI21_X1 U5743 ( .B1(n4804), .B2(n4806), .A(n4533), .ZN(n4802) );
  INV_X1 U5744 ( .A(n6650), .ZN(n8556) );
  NAND2_X1 U5745 ( .A1(n6141), .A2(n6140), .ZN(n9010) );
  INV_X1 U5746 ( .A(n4826), .ZN(n4825) );
  OAI21_X1 U5747 ( .B1(n4503), .B2(n4827), .A(n6607), .ZN(n4826) );
  OR2_X1 U5748 ( .A1(n4478), .A2(n7803), .ZN(n6227) );
  NAND2_X1 U5749 ( .A1(n4814), .A2(n4820), .ZN(n8593) );
  NAND2_X1 U5750 ( .A1(n8610), .A2(n4822), .ZN(n4814) );
  OR2_X1 U5751 ( .A1(n4478), .A2(n7659), .ZN(n6207) );
  NAND2_X1 U5752 ( .A1(n4803), .A2(n4807), .ZN(n7703) );
  NAND2_X1 U5753 ( .A1(n4583), .A2(n4810), .ZN(n4803) );
  INV_X1 U5754 ( .A(n7204), .ZN(n7125) );
  AND4_X1 U5755 ( .A1(n6162), .A2(n6161), .A3(n6160), .A4(n6159), .ZN(n8869)
         );
  NAND2_X1 U5756 ( .A1(n7100), .A2(n6558), .ZN(n7381) );
  AND2_X1 U5757 ( .A1(n6683), .A2(n8912), .ZN(n8634) );
  AND2_X1 U5758 ( .A1(n6698), .A2(n6697), .ZN(n8631) );
  INV_X1 U5759 ( .A(n8634), .ZN(n8618) );
  NAND2_X1 U5760 ( .A1(n4506), .A2(n6502), .ZN(n6510) );
  NAND2_X1 U5761 ( .A1(n6501), .A2(n6500), .ZN(n6502) );
  AND2_X1 U5762 ( .A1(n4628), .A2(n4626), .ZN(n4625) );
  INV_X1 U5763 ( .A(n8626), .ZN(n8637) );
  INV_X1 U5764 ( .A(n6559), .ZN(n8644) );
  NAND2_X1 U5765 ( .A1(n5925), .A2(n5924), .ZN(n8650) );
  INV_X1 U5766 ( .A(P2_U3966), .ZN(n8649) );
  NOR2_X1 U5767 ( .A1(n6845), .A2(n6846), .ZN(n4694) );
  AOI21_X1 U5768 ( .B1(n6848), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6925), .ZN(
        n6865) );
  NOR2_X1 U5769 ( .A1(n6864), .A2(n6865), .ZN(n6863) );
  AOI21_X1 U5770 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n6849), .A(n6863), .ZN(
        n6854) );
  INV_X1 U5771 ( .A(n4703), .ZN(n6893) );
  NAND2_X1 U5772 ( .A1(n6915), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4700) );
  NOR2_X1 U5773 ( .A1(n7063), .A2(n4552), .ZN(n7066) );
  INV_X1 U5774 ( .A(n7118), .ZN(n7117) );
  OAI21_X1 U5775 ( .B1(n7551), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7550), .ZN(
        n7554) );
  INV_X1 U5776 ( .A(n4706), .ZN(n7602) );
  INV_X1 U5777 ( .A(n4699), .ZN(n8651) );
  NOR2_X1 U5778 ( .A1(n8655), .A2(n8654), .ZN(n8672) );
  AND2_X1 U5779 ( .A1(n4699), .A2(n4698), .ZN(n8655) );
  NAND2_X1 U5780 ( .A1(n8652), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4698) );
  NOR2_X1 U5781 ( .A1(n8691), .A2(n4708), .ZN(n8675) );
  AND2_X1 U5782 ( .A1(n8674), .A2(n8673), .ZN(n4708) );
  OAI21_X1 U5783 ( .B1(n8705), .B2(n8706), .A(n8704), .ZN(n4582) );
  NAND2_X1 U5784 ( .A1(n6325), .A2(n6832), .ZN(n8941) );
  MUX2_X1 U5785 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9169), .S(n5936), .Z(n6325) );
  XNOR2_X1 U5786 ( .A(n8707), .B(n4738), .ZN(n8939) );
  INV_X1 U5787 ( .A(n8941), .ZN(n4738) );
  AOI21_X1 U5788 ( .B1(n9171), .B2(n6291), .A(n6305), .ZN(n8945) );
  NOR2_X1 U5789 ( .A1(n4478), .A2(n9051), .ZN(n6305) );
  AOI21_X1 U5790 ( .B1(n8488), .B2(n8493), .A(n8131), .ZN(n8132) );
  NAND2_X1 U5791 ( .A1(n6293), .A2(n6292), .ZN(n8716) );
  OR2_X1 U5792 ( .A1(n4478), .A2(n8486), .ZN(n6292) );
  INV_X1 U5793 ( .A(n4737), .ZN(n8720) );
  INV_X1 U5794 ( .A(n8946), .ZN(n8492) );
  NAND2_X1 U5795 ( .A1(n4919), .A2(n4922), .ZN(n8724) );
  NAND2_X1 U5796 ( .A1(n8754), .A2(n4924), .ZN(n4919) );
  AOI21_X1 U5797 ( .B1(n8754), .B2(n8129), .A(n4925), .ZN(n8740) );
  NAND2_X1 U5798 ( .A1(n4904), .A2(n4905), .ZN(n8770) );
  AND2_X1 U5799 ( .A1(n4908), .A2(n4513), .ZN(n8792) );
  AND2_X1 U5800 ( .A1(n4723), .A2(n6423), .ZN(n5032) );
  NAND2_X1 U5801 ( .A1(n8890), .A2(n8118), .ZN(n8863) );
  NOR2_X1 U5802 ( .A1(n8906), .A2(n8905), .ZN(n9015) );
  NAND2_X1 U5803 ( .A1(n9968), .A2(n6121), .ZN(n8926) );
  AND2_X1 U5804 ( .A1(n4933), .A2(n8117), .ZN(n8920) );
  INV_X1 U5805 ( .A(n4933), .ZN(n9973) );
  NAND2_X1 U5806 ( .A1(n7970), .A2(n7969), .ZN(n7972) );
  NAND2_X1 U5807 ( .A1(n4715), .A2(n4713), .ZN(n7888) );
  NAND2_X1 U5808 ( .A1(n6078), .A2(n4714), .ZN(n7752) );
  NAND2_X1 U5809 ( .A1(n7633), .A2(n7566), .ZN(n7567) );
  NAND2_X1 U5810 ( .A1(n6007), .A2(n6368), .ZN(n7642) );
  INV_X1 U5811 ( .A(n10283), .ZN(n8912) );
  NAND2_X1 U5812 ( .A1(n5966), .A2(n6349), .ZN(n7182) );
  AND2_X1 U5813 ( .A1(n8915), .A2(n10279), .ZN(n10288) );
  INV_X1 U5814 ( .A(n10284), .ZN(n8924) );
  INV_X1 U5815 ( .A(n10288), .ZN(n8938) );
  NAND2_X1 U5816 ( .A1(n5913), .A2(n5914), .ZN(n9045) );
  NAND2_X1 U5817 ( .A1(n6515), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U5818 ( .A1(n5891), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4833) );
  INV_X1 U5819 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6760) );
  INV_X1 U5820 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6748) );
  INV_X1 U5821 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6737) );
  NAND2_X1 U5822 ( .A1(n5939), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5948) );
  INV_X1 U5823 ( .A(n4643), .ZN(n9068) );
  AOI21_X1 U5824 ( .B1(n4486), .B2(n9105), .A(n4526), .ZN(n4669) );
  NAND2_X1 U5825 ( .A1(n4947), .A2(n5314), .ZN(n7420) );
  INV_X1 U5826 ( .A(n4950), .ZN(n4947) );
  NAND2_X1 U5827 ( .A1(n4950), .A2(n5313), .ZN(n7419) );
  INV_X1 U5828 ( .A(n10185), .ZN(n8039) );
  NAND2_X1 U5829 ( .A1(n5731), .A2(n5730), .ZN(n9808) );
  NAND2_X1 U5830 ( .A1(n5527), .A2(n5526), .ZN(n9846) );
  OAI21_X1 U5831 ( .B1(n5672), .B2(n4636), .A(n4639), .ZN(n4635) );
  INV_X1 U5832 ( .A(n10210), .ZN(n7476) );
  NAND2_X1 U5833 ( .A1(n7794), .A2(n5420), .ZN(n7832) );
  NAND2_X1 U5834 ( .A1(n4662), .A2(n4659), .ZN(n4658) );
  NAND2_X1 U5835 ( .A1(n9103), .A2(n4941), .ZN(n8045) );
  NAND2_X1 U5836 ( .A1(n4937), .A2(n5567), .ZN(n8044) );
  NAND2_X1 U5837 ( .A1(n9103), .A2(n5541), .ZN(n4937) );
  AND4_X1 U5838 ( .A1(n5411), .A2(n5410), .A3(n5409), .A4(n5408), .ZN(n7899)
         );
  AND4_X1 U5839 ( .A1(n5357), .A2(n5356), .A3(n5355), .A4(n5354), .ZN(n7816)
         );
  NAND2_X1 U5840 ( .A1(n5203), .A2(n4961), .ZN(n5151) );
  OR2_X1 U5841 ( .A1(n5175), .A2(n5127), .ZN(n5130) );
  OR2_X1 U5842 ( .A1(n5806), .A2(n5126), .ZN(n5131) );
  OR2_X1 U5843 ( .A1(n6710), .A2(n6752), .ZN(n9479) );
  NAND2_X1 U5844 ( .A1(n5203), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5102) );
  XNOR2_X1 U5845 ( .A(n4751), .B(n5048), .ZN(n9458) );
  OAI21_X1 U5846 ( .B1(n5068), .B2(n4753), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4751) );
  NAND2_X1 U5847 ( .A1(n4754), .A2(n4539), .ZN(n4753) );
  INV_X1 U5848 ( .A(n4482), .ZN(n4754) );
  NAND2_X1 U5849 ( .A1(n5803), .A2(n5802), .ZN(n9791) );
  AND2_X1 U5850 ( .A1(n5754), .A2(n5753), .ZN(n9591) );
  NAND2_X1 U5851 ( .A1(n4992), .A2(n4995), .ZN(n9586) );
  NAND2_X1 U5852 ( .A1(n4998), .A2(n4997), .ZN(n4992) );
  NAND2_X1 U5853 ( .A1(n4755), .A2(n9319), .ZN(n9608) );
  NAND2_X1 U5854 ( .A1(n4998), .A2(n9250), .ZN(n9600) );
  NAND2_X1 U5855 ( .A1(n8070), .A2(n5001), .ZN(n9615) );
  NAND2_X1 U5856 ( .A1(n5626), .A2(n5625), .ZN(n9827) );
  NAND2_X1 U5857 ( .A1(n4966), .A2(n4970), .ZN(n9677) );
  OR2_X1 U5858 ( .A1(n4972), .A2(n4971), .ZN(n4966) );
  NOR2_X1 U5859 ( .A1(n4553), .A2(n4974), .ZN(n9692) );
  NAND2_X1 U5860 ( .A1(n8082), .A2(n9378), .ZN(n9729) );
  NAND2_X1 U5861 ( .A1(n5010), .A2(n5012), .ZN(n9737) );
  NAND2_X1 U5862 ( .A1(n5011), .A2(n5018), .ZN(n9756) );
  OR2_X1 U5863 ( .A1(n8064), .A2(n8063), .ZN(n5011) );
  INV_X1 U5864 ( .A(n9759), .ZN(n9858) );
  AND2_X1 U5865 ( .A1(n4770), .A2(n4530), .ZN(n7961) );
  NAND2_X1 U5866 ( .A1(n5405), .A2(n5404), .ZN(n9996) );
  NAND2_X1 U5867 ( .A1(n5350), .A2(n5349), .ZN(n9948) );
  NAND2_X1 U5868 ( .A1(n7780), .A2(n7779), .ZN(n7807) );
  INV_X1 U5869 ( .A(n10229), .ZN(n7778) );
  AND2_X1 U5870 ( .A1(n4985), .A2(n4537), .ZN(n7485) );
  NAND2_X1 U5871 ( .A1(n4985), .A2(n4984), .ZN(n7484) );
  NAND2_X1 U5872 ( .A1(n4986), .A2(n9262), .ZN(n4985) );
  INV_X1 U5873 ( .A(n9742), .ZN(n9947) );
  NAND2_X1 U5874 ( .A1(n9774), .A2(n10183), .ZN(n9742) );
  INV_X1 U5875 ( .A(n9735), .ZN(n9550) );
  AOI211_X1 U5876 ( .C1(n9994), .C2(n9993), .A(n9992), .B(n9991), .ZN(n10011)
         );
  AOI21_X1 U5877 ( .B1(n8097), .B2(n9772), .A(n4776), .ZN(n9789) );
  XNOR2_X1 U5878 ( .A(n6287), .B(n6286), .ZN(n8015) );
  XNOR2_X1 U5879 ( .A(n5799), .B(n5798), .ZN(n7989) );
  NAND2_X1 U5880 ( .A1(n4960), .A2(n4959), .ZN(n5065) );
  NOR2_X1 U5881 ( .A1(n4482), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4959) );
  INV_X1 U5882 ( .A(n9462), .ZN(n9452) );
  INV_X1 U5883 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8352) );
  INV_X1 U5884 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6750) );
  INV_X1 U5885 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6736) );
  INV_X1 U5886 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6732) );
  NOR2_X1 U5887 ( .A1(n7855), .A2(n10438), .ZN(n10458) );
  NOR2_X1 U5888 ( .A1(n10458), .A2(n10457), .ZN(n10456) );
  AOI21_X1 U5889 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10456), .ZN(n10461) );
  NOR2_X1 U5890 ( .A1(n7858), .A2(n10453), .ZN(n10437) );
  AOI21_X1 U5891 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10435), .ZN(n10434) );
  NOR2_X1 U5892 ( .A1(n10434), .A2(n10433), .ZN(n10432) );
  INV_X1 U5893 ( .A(n4701), .ZN(n6911) );
  OAI211_X1 U5894 ( .C1(n8703), .C2(n8701), .A(n4581), .B(n4579), .ZN(P2_U3264) );
  INV_X1 U5895 ( .A(n4582), .ZN(n4581) );
  NAND2_X1 U5896 ( .A1(n4580), .A2(n8701), .ZN(n4579) );
  AOI21_X1 U5897 ( .B1(n4953), .B2(n4657), .A(n4651), .ZN(n4650) );
  NAND2_X1 U5898 ( .A1(n4954), .A2(n4555), .ZN(n5873) );
  OR2_X1 U5899 ( .A1(n9464), .A2(n9463), .ZN(n4880) );
  NAND2_X1 U5900 ( .A1(n4602), .A2(n4600), .ZN(P1_U3260) );
  AOI21_X1 U5901 ( .B1(n9535), .B2(n10180), .A(n4601), .ZN(n4600) );
  NAND2_X1 U5902 ( .A1(n9536), .A2(n9671), .ZN(n4602) );
  OAI21_X1 U5903 ( .B1(n10175), .B2(n4890), .A(n9537), .ZN(n4601) );
  NAND2_X1 U5904 ( .A1(n4772), .A2(n4498), .ZN(n4773) );
  AND2_X1 U5905 ( .A1(n9343), .A2(n9349), .ZN(n9266) );
  NAND2_X1 U5906 ( .A1(n5047), .A2(n5046), .ZN(n4482) );
  OR2_X1 U5907 ( .A1(n9022), .A2(n8115), .ZN(n4483) );
  INV_X2 U5908 ( .A(n6612), .ZN(n8108) );
  OR2_X1 U5909 ( .A1(n5672), .A2(n5671), .ZN(n4484) );
  AND2_X1 U5910 ( .A1(n9296), .A2(n9333), .ZN(n7408) );
  INV_X1 U5911 ( .A(n8966), .ZN(n8773) );
  NAND2_X1 U5912 ( .A1(n6228), .A2(n6227), .ZN(n8966) );
  NAND2_X1 U5913 ( .A1(n5681), .A2(n5680), .ZN(n9816) );
  NOR2_X1 U5914 ( .A1(n7806), .A2(n5004), .ZN(n4485) );
  OR2_X1 U5915 ( .A1(n4941), .A2(n4938), .ZN(n4486) );
  AND2_X1 U5916 ( .A1(n9712), .A2(n4761), .ZN(n4487) );
  INV_X1 U5917 ( .A(n5541), .ZN(n4940) );
  NAND2_X1 U5918 ( .A1(n9698), .A2(n9681), .ZN(n4488) );
  NAND2_X1 U5919 ( .A1(n5656), .A2(n5655), .ZN(n9821) );
  INV_X1 U5920 ( .A(n9821), .ZN(n4685) );
  OR3_X1 U5921 ( .A1(n4749), .A2(n8803), .A3(n8966), .ZN(n4489) );
  INV_X1 U5922 ( .A(n4923), .ZN(n4922) );
  OAI22_X1 U5923 ( .A1(n8747), .A2(n4926), .B1(n8734), .B2(n8957), .ZN(n4923)
         );
  AND2_X1 U5924 ( .A1(n9563), .A2(n9576), .ZN(n4490) );
  AND2_X1 U5925 ( .A1(n9319), .A2(n9415), .ZN(n4491) );
  NAND2_X1 U5926 ( .A1(n9622), .A2(n9409), .ZN(n9639) );
  INV_X1 U5927 ( .A(n9639), .ZN(n8090) );
  NAND2_X1 U5928 ( .A1(n9175), .A2(n9174), .ZN(n9993) );
  NOR3_X1 U5929 ( .A1(n4749), .A2(n8966), .A3(n8963), .ZN(n4492) );
  NAND2_X1 U5930 ( .A1(n4492), .A2(n4748), .ZN(n8760) );
  INV_X1 U5931 ( .A(n8760), .ZN(n4598) );
  OR2_X1 U5932 ( .A1(n6470), .A2(n4633), .ZN(n4493) );
  NOR2_X1 U5933 ( .A1(n8105), .A2(n4776), .ZN(n4494) );
  AND2_X1 U5934 ( .A1(n4979), .A2(n4981), .ZN(n4495) );
  AND2_X1 U5935 ( .A1(n4873), .A2(n5722), .ZN(n4496) );
  AND2_X1 U5936 ( .A1(n4678), .A2(n4677), .ZN(n4497) );
  NOR2_X1 U5937 ( .A1(n8105), .A2(n4565), .ZN(n4498) );
  NAND2_X1 U5938 ( .A1(n6097), .A2(n6096), .ZN(n8114) );
  INV_X2 U5939 ( .A(n5273), .ZN(n5368) );
  NAND2_X1 U5940 ( .A1(n4831), .A2(n6331), .ZN(n6467) );
  NAND2_X1 U5941 ( .A1(n8070), .A2(n4999), .ZN(n4998) );
  NAND2_X1 U5942 ( .A1(n8644), .A2(n7279), .ZN(n4895) );
  INV_X1 U5943 ( .A(n8701), .ZN(n4831) );
  OR2_X1 U5944 ( .A1(n9972), .A2(n8929), .ZN(n8117) );
  OR2_X1 U5945 ( .A1(n5498), .A2(n4854), .ZN(n4499) );
  NAND2_X2 U5946 ( .A1(n5086), .A2(n9903), .ZN(n5806) );
  AND2_X1 U5947 ( .A1(n4701), .A2(n4700), .ZN(n4500) );
  AND2_X1 U5948 ( .A1(n4637), .A2(n4634), .ZN(n4501) );
  NOR2_X1 U5949 ( .A1(n9917), .A2(n4694), .ZN(n4502) );
  NAND2_X1 U5950 ( .A1(n4908), .A2(n4907), .ZN(n8793) );
  INV_X1 U5951 ( .A(n6570), .ZN(n6612) );
  NAND2_X1 U5952 ( .A1(n5701), .A2(n5700), .ZN(n9811) );
  AND2_X1 U5953 ( .A1(n4829), .A2(n6594), .ZN(n4503) );
  XNOR2_X1 U5954 ( .A(n8951), .B(n8626), .ZN(n8733) );
  AND2_X1 U5955 ( .A1(n9975), .A2(n6401), .ZN(n4504) );
  AND4_X1 U5956 ( .A1(n5040), .A2(n5039), .A3(n5038), .A4(n5037), .ZN(n4505)
         );
  NAND2_X1 U5957 ( .A1(n4627), .A2(n4625), .ZN(n4506) );
  XNOR2_X1 U5958 ( .A(n8963), .B(n8777), .ZN(n8129) );
  INV_X1 U5959 ( .A(n8129), .ZN(n8756) );
  INV_X1 U5960 ( .A(n7757), .ZN(n6078) );
  OR2_X1 U5961 ( .A1(n10051), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4507) );
  INV_X1 U5962 ( .A(n7750), .ZN(n4717) );
  AND2_X1 U5963 ( .A1(n4589), .A2(n4588), .ZN(n4508) );
  NAND2_X1 U5964 ( .A1(n9603), .A2(n9469), .ZN(n4509) );
  AND2_X1 U5965 ( .A1(n9836), .A2(n9714), .ZN(n4510) );
  INV_X1 U5966 ( .A(n7697), .ZN(n4664) );
  INV_X2 U5967 ( .A(n7361), .ZN(n5814) );
  INV_X1 U5968 ( .A(n9070), .ZN(n4645) );
  NAND2_X1 U5969 ( .A1(n6110), .A2(n6109), .ZN(n9972) );
  OR3_X1 U5970 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4511) );
  OR2_X1 U5971 ( .A1(n8987), .A2(n8548), .ZN(n6423) );
  AND2_X1 U5972 ( .A1(n9594), .A2(n9423), .ZN(n4512) );
  NAND2_X1 U5973 ( .A1(n8807), .A2(n8547), .ZN(n4513) );
  NAND2_X1 U5974 ( .A1(n5374), .A2(n5373), .ZN(n7895) );
  AND2_X1 U5975 ( .A1(n9592), .A2(n8092), .ZN(n4514) );
  NAND2_X1 U5976 ( .A1(n5073), .A2(n5075), .ZN(n5068) );
  INV_X1 U5977 ( .A(n5068), .ZN(n4960) );
  AND2_X1 U5978 ( .A1(n4504), .A2(n8927), .ZN(n4515) );
  NAND2_X1 U5979 ( .A1(n7895), .A2(n7812), .ZN(n4516) );
  NOR2_X1 U5980 ( .A1(n9668), .A2(n4682), .ZN(n4681) );
  AND2_X1 U5981 ( .A1(n6402), .A2(n6401), .ZN(n7971) );
  AND2_X1 U5982 ( .A1(n6560), .A2(n6558), .ZN(n4517) );
  AND2_X1 U5983 ( .A1(n4643), .A2(n4645), .ZN(n4518) );
  AND2_X1 U5984 ( .A1(n5198), .A2(n5173), .ZN(n4519) );
  AND2_X1 U5985 ( .A1(n5419), .A2(n5390), .ZN(n4520) );
  AND2_X1 U5986 ( .A1(n7880), .A2(n7878), .ZN(n4521) );
  NOR2_X1 U5987 ( .A1(n5771), .A2(n4952), .ZN(n4522) );
  INV_X1 U5988 ( .A(n4811), .ZN(n4810) );
  OR2_X1 U5989 ( .A1(n7662), .A2(n4812), .ZN(n4811) );
  INV_X1 U5990 ( .A(n4943), .ZN(n4942) );
  NOR2_X1 U5991 ( .A1(n4948), .A2(n5313), .ZN(n4943) );
  AND2_X1 U5992 ( .A1(n5088), .A2(n5087), .ZN(n4523) );
  INV_X1 U5993 ( .A(n8982), .ZN(n8823) );
  NAND2_X1 U5994 ( .A1(n8500), .A2(n5083), .ZN(n5738) );
  AND2_X1 U5995 ( .A1(n8972), .A2(n8127), .ZN(n4524) );
  OR2_X1 U5996 ( .A1(n9808), .A2(n9469), .ZN(n9415) );
  NAND2_X1 U5997 ( .A1(n4997), .A2(n8071), .ZN(n4525) );
  AND2_X1 U5998 ( .A1(n6377), .A2(n6376), .ZN(n7572) );
  OR2_X1 U5999 ( .A1(n9016), .A2(n8576), .ZN(n6407) );
  AND2_X1 U6000 ( .A1(n4938), .A2(n5568), .ZN(n4526) );
  NOR2_X1 U6001 ( .A1(n9474), .A2(n7498), .ZN(n4527) );
  INV_X1 U6002 ( .A(n8963), .ZN(n8765) );
  NAND2_X1 U6003 ( .A1(n6240), .A2(n6239), .ZN(n8963) );
  OR2_X1 U6004 ( .A1(n4615), .A2(n8905), .ZN(n4528) );
  NOR2_X1 U6005 ( .A1(n9689), .A2(n9079), .ZN(n4529) );
  NAND2_X1 U6006 ( .A1(n9869), .A2(n9188), .ZN(n4530) );
  INV_X1 U6007 ( .A(n4926), .ZN(n4925) );
  AND2_X1 U6008 ( .A1(n8090), .A2(n9410), .ZN(n4531) );
  AND2_X1 U6009 ( .A1(n8729), .A2(n8626), .ZN(n4532) );
  AND2_X1 U6010 ( .A1(n6585), .A2(n6584), .ZN(n4533) );
  INV_X1 U6011 ( .A(n5019), .ZN(n5018) );
  NOR2_X1 U6012 ( .A1(n9067), .A2(n9162), .ZN(n5019) );
  NOR2_X1 U6013 ( .A1(n10236), .A2(n9937), .ZN(n4534) );
  OR2_X1 U6014 ( .A1(n5068), .A2(n4482), .ZN(n4535) );
  NOR2_X1 U6015 ( .A1(n5091), .A2(n5044), .ZN(n5073) );
  INV_X1 U6016 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5081) );
  NOR2_X1 U6017 ( .A1(n9016), .A2(n8902), .ZN(n4536) );
  INV_X1 U6018 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5063) );
  INV_X1 U6019 ( .A(n4689), .ZN(n4688) );
  NAND2_X1 U6020 ( .A1(n4490), .A2(n4690), .ZN(n4689) );
  INV_X1 U6021 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5911) );
  NAND2_X1 U6022 ( .A1(n9475), .A2(n7409), .ZN(n4537) );
  NAND2_X1 U6023 ( .A1(n9802), .A2(n9468), .ZN(n4538) );
  AND2_X1 U6024 ( .A1(n5063), .A2(n5066), .ZN(n4539) );
  AND3_X1 U6025 ( .A1(n5143), .A2(n5142), .A3(n5141), .ZN(n10205) );
  INV_X1 U6026 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6083) );
  AND2_X1 U6027 ( .A1(n5393), .A2(SI_11_), .ZN(n4540) );
  INV_X1 U6028 ( .A(n9181), .ZN(n4797) );
  OR2_X1 U6029 ( .A1(n4510), .A2(n4974), .ZN(n4541) );
  INV_X1 U6030 ( .A(n9816), .ZN(n9635) );
  INV_X1 U6031 ( .A(n4973), .ZN(n4971) );
  AND2_X1 U6032 ( .A1(n4488), .A2(n9706), .ZN(n4973) );
  AND2_X1 U6033 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n9895), .ZN(n4542) );
  OR2_X1 U6034 ( .A1(n9791), .A2(n9580), .ZN(n9426) );
  AND2_X1 U6035 ( .A1(n7285), .A2(n7290), .ZN(n4543) );
  AND2_X1 U6036 ( .A1(n5015), .A2(n5016), .ZN(n4544) );
  OR2_X1 U6037 ( .A1(n6832), .A2(n6845), .ZN(n4545) );
  NAND2_X1 U6038 ( .A1(n9313), .A2(n9432), .ZN(n9434) );
  AND2_X1 U6039 ( .A1(n6393), .A2(n6392), .ZN(n7887) );
  AND2_X1 U6040 ( .A1(n9378), .A2(n9377), .ZN(n9738) );
  INV_X1 U6041 ( .A(n9738), .ZN(n5009) );
  INV_X1 U6042 ( .A(n9864), .ZN(n9067) );
  NAND2_X1 U6043 ( .A1(n5452), .A2(n5451), .ZN(n9864) );
  AND2_X1 U6044 ( .A1(n4792), .A2(n9184), .ZN(n4546) );
  OR2_X1 U6045 ( .A1(n6379), .A2(n7711), .ZN(n4547) );
  AND2_X1 U6046 ( .A1(n6416), .A2(n4528), .ZN(n4548) );
  OR2_X1 U6047 ( .A1(n6582), .A2(n6581), .ZN(n4549) );
  AND2_X1 U6048 ( .A1(n8791), .A2(n4513), .ZN(n4907) );
  NAND2_X1 U6049 ( .A1(n5317), .A2(n5294), .ZN(n5316) );
  INV_X2 U6050 ( .A(n5115), .ZN(n5816) );
  AND2_X1 U6051 ( .A1(n9791), .A2(n8072), .ZN(n4550) );
  OR2_X1 U6052 ( .A1(n8908), .A2(n4746), .ZN(n4551) );
  NAND2_X1 U6053 ( .A1(n10180), .A2(n9452), .ZN(n9440) );
  INV_X1 U6054 ( .A(n9833), .ZN(n9689) );
  NAND2_X1 U6055 ( .A1(n5607), .A2(n5606), .ZN(n9833) );
  NAND2_X1 U6056 ( .A1(n5003), .A2(n5002), .ZN(n9928) );
  INV_X1 U6057 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5237) );
  AND2_X1 U6058 ( .A1(n7064), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4552) );
  AND2_X1 U6059 ( .A1(n9707), .A2(n9706), .ZN(n4553) );
  OR2_X1 U6060 ( .A1(n8908), .A2(n9005), .ZN(n4554) );
  NAND2_X1 U6061 ( .A1(n6251), .A2(n6250), .ZN(n8957) );
  INV_X1 U6062 ( .A(n8957), .ZN(n4597) );
  AND3_X1 U6063 ( .A1(n5866), .A2(n9152), .A3(n5865), .ZN(n4555) );
  NAND2_X1 U6064 ( .A1(n8074), .A2(n8073), .ZN(n9786) );
  INV_X1 U6065 ( .A(n9786), .ZN(n4690) );
  AND3_X1 U6066 ( .A1(n6205), .A2(n6204), .A3(n6203), .ZN(n8812) );
  AND3_X1 U6067 ( .A1(n5220), .A2(n5219), .A3(n5218), .ZN(n10217) );
  OR2_X1 U6068 ( .A1(n7881), .A2(n4744), .ZN(n4556) );
  NAND2_X1 U6069 ( .A1(n6105), .A2(n6401), .ZN(n4557) );
  INV_X1 U6070 ( .A(n9796), .ZN(n9576) );
  NAND2_X1 U6071 ( .A1(n5784), .A2(n5783), .ZN(n9796) );
  AND2_X1 U6072 ( .A1(n5010), .A2(n5008), .ZN(n4558) );
  INV_X1 U6073 ( .A(n4693), .ZN(n9723) );
  NOR2_X1 U6074 ( .A1(n9740), .A2(n9846), .ZN(n4693) );
  INV_X1 U6075 ( .A(n4686), .ZN(n9647) );
  NOR2_X1 U6076 ( .A1(n9668), .A2(n9821), .ZN(n4686) );
  NOR2_X1 U6077 ( .A1(n5427), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5449) );
  NAND3_X1 U6078 ( .A1(n5899), .A2(n5900), .A3(n4898), .ZN(n4559) );
  AND2_X1 U6079 ( .A1(n5724), .A2(SI_24_), .ZN(n4560) );
  AND2_X1 U6080 ( .A1(n4745), .A2(n9022), .ZN(n4561) );
  AND2_X1 U6081 ( .A1(n5646), .A2(n5624), .ZN(n4562) );
  AND2_X1 U6082 ( .A1(n5881), .A2(n5880), .ZN(n4563) );
  NAND2_X1 U6083 ( .A1(n5581), .A2(n5580), .ZN(n9836) );
  NOR2_X1 U6084 ( .A1(n9015), .A2(n4916), .ZN(n4564) );
  NOR2_X1 U6085 ( .A1(n4775), .A2(n10193), .ZN(n4565) );
  INV_X1 U6086 ( .A(n8104), .ZN(n4776) );
  NAND2_X1 U6087 ( .A1(n5285), .A2(n7249), .ZN(n4950) );
  INV_X1 U6088 ( .A(n9273), .ZN(n4767) );
  INV_X1 U6089 ( .A(n9866), .ZN(n4981) );
  NAND2_X1 U6090 ( .A1(n4725), .A2(n4724), .ZN(n7570) );
  AND2_X1 U6091 ( .A1(n9325), .A2(n4537), .ZN(n4984) );
  OAI21_X1 U6092 ( .B1(n4944), .B2(n4664), .A(n4662), .ZN(n7532) );
  NAND2_X1 U6093 ( .A1(n4944), .A2(n4942), .ZN(n7696) );
  INV_X1 U6094 ( .A(n9333), .ZN(n4783) );
  NAND2_X1 U6095 ( .A1(n5430), .A2(n5429), .ZN(n9869) );
  INV_X1 U6096 ( .A(n9869), .ZN(n4677) );
  INV_X1 U6097 ( .A(n9975), .ZN(n4935) );
  NAND2_X1 U6098 ( .A1(n4958), .A2(n5390), .ZN(n7793) );
  NAND2_X1 U6099 ( .A1(n5174), .A2(n4519), .ZN(n7057) );
  OR2_X1 U6100 ( .A1(n9474), .A2(n10222), .ZN(n9336) );
  INV_X1 U6101 ( .A(n9336), .ZN(n4781) );
  NAND2_X1 U6102 ( .A1(n5174), .A2(n5173), .ZN(n7055) );
  NAND2_X1 U6103 ( .A1(n9949), .A2(n4497), .ZN(n4679) );
  NAND2_X1 U6104 ( .A1(n6575), .A2(n6576), .ZN(n4566) );
  AND2_X1 U6105 ( .A1(n6304), .A2(n6303), .ZN(n4567) );
  AND2_X1 U6106 ( .A1(n7879), .A2(n7878), .ZN(n4568) );
  INV_X1 U6107 ( .A(n4832), .ZN(n9978) );
  AND3_X1 U6108 ( .A1(n5844), .A2(n6956), .A3(n6960), .ZN(n9152) );
  INV_X1 U6109 ( .A(n9671), .ZN(n10180) );
  BUF_X1 U6111 ( .A(n7152), .Z(n9480) );
  INV_X1 U6112 ( .A(n7152), .ZN(n4672) );
  INV_X1 U6113 ( .A(n4680), .ZN(n7473) );
  NOR2_X1 U6114 ( .A1(n7471), .A2(n7476), .ZN(n4680) );
  INV_X1 U6115 ( .A(n7504), .ZN(n4629) );
  INV_X1 U6116 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5097) );
  INV_X1 U6117 ( .A(n5086), .ZN(n8500) );
  INV_X1 U6118 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4890) );
  NAND2_X1 U6119 ( .A1(n4620), .A2(n6467), .ZN(n4619) );
  INV_X1 U6120 ( .A(n6467), .ZN(n4618) );
  NOR2_X2 U6121 ( .A1(n5898), .A2(n5897), .ZN(n5899) );
  NAND2_X1 U6122 ( .A1(n8757), .A2(n8756), .ZN(n8755) );
  INV_X1 U6123 ( .A(n7975), .ZN(n4570) );
  INV_X1 U6124 ( .A(n7088), .ZN(n5950) );
  NAND2_X1 U6125 ( .A1(n5966), .A2(n4728), .ZN(n7456) );
  AOI21_X1 U6126 ( .B1(n6327), .B2(n6496), .A(n6468), .ZN(n6328) );
  NAND2_X2 U6127 ( .A1(n5949), .A2(n4569), .ZN(n7204) );
  AND2_X1 U6128 ( .A1(n4594), .A2(n4545), .ZN(n4569) );
  INV_X1 U6129 ( .A(n4635), .ZN(n4634) );
  INV_X1 U6130 ( .A(n4954), .ZN(n5876) );
  NAND2_X1 U6131 ( .A1(n4837), .A2(n5624), .ZN(n5645) );
  AND2_X2 U6132 ( .A1(n9055), .A2(n5494), .ZN(n5493) );
  NAND2_X1 U6133 ( .A1(n7057), .A2(n5201), .ZN(n7329) );
  NOR2_X2 U6134 ( .A1(n5348), .A2(n5093), .ZN(n5400) );
  INV_X1 U6135 ( .A(n4648), .ZN(n4647) );
  NAND2_X1 U6136 ( .A1(n4670), .A2(n4669), .ZN(n8057) );
  NAND2_X2 U6137 ( .A1(n5644), .A2(n5643), .ZN(n5672) );
  NAND2_X1 U6138 ( .A1(n5136), .A2(n5135), .ZN(n5156) );
  NAND2_X1 U6140 ( .A1(n8126), .A2(n4573), .ZN(n8801) );
  INV_X1 U6142 ( .A(n7561), .ZN(n7562) );
  MUX2_X1 U6143 ( .A(n9355), .B(n9354), .S(n9406), .Z(n9366) );
  OAI21_X1 U6144 ( .B1(n9366), .B2(n9365), .A(n9364), .ZN(n9372) );
  OR2_X1 U6145 ( .A1(n9324), .A2(n9323), .ZN(n9327) );
  AOI211_X1 U6146 ( .C1(n9407), .C2(n9406), .A(n4575), .B(n9413), .ZN(n9417)
         );
  NAND3_X1 U6147 ( .A1(n9340), .A2(n9440), .A3(n9339), .ZN(n4578) );
  AOI21_X1 U6148 ( .B1(n8831), .B2(n8839), .A(n8123), .ZN(n8819) );
  NAND2_X1 U6149 ( .A1(n7158), .A2(n7157), .ZN(n7216) );
  NAND2_X1 U6150 ( .A1(n4901), .A2(n4907), .ZN(n4904) );
  NAND2_X1 U6151 ( .A1(n4883), .A2(n4882), .ZN(n4881) );
  NAND2_X1 U6152 ( .A1(n4931), .A2(n4929), .ZN(n8906) );
  NAND2_X1 U6153 ( .A1(n7757), .A2(n7758), .ZN(n7879) );
  AOI21_X1 U6154 ( .B1(n8722), .B2(n10391), .A(n4736), .ZN(n4735) );
  NOR2_X1 U6155 ( .A1(n4737), .A2(n4734), .ZN(n8143) );
  INV_X1 U6156 ( .A(n7066), .ZN(n4587) );
  NOR2_X1 U6157 ( .A1(n9919), .A2(n9918), .ZN(n9917) );
  XNOR2_X1 U6158 ( .A(n6635), .B(n6633), .ZN(n8602) );
  OAI21_X1 U6159 ( .B1(n5547), .B2(n5546), .A(n5545), .ZN(n5571) );
  NAND2_X2 U6160 ( .A1(n6067), .A2(n6066), .ZN(n7877) );
  NAND2_X1 U6161 ( .A1(n4869), .A2(n5367), .ZN(n5395) );
  INV_X1 U6162 ( .A(n4589), .ZN(n8690) );
  INV_X1 U6163 ( .A(n8691), .ZN(n4588) );
  NAND2_X1 U6164 ( .A1(n8675), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n4589) );
  NAND2_X1 U6165 ( .A1(n8002), .A2(n8003), .ZN(n8005) );
  NAND2_X1 U6166 ( .A1(n7120), .A2(n7121), .ZN(n7238) );
  MUX2_X1 U6167 ( .A(n9431), .B(n9430), .S(n9440), .Z(n9435) );
  NAND2_X1 U6168 ( .A1(n4590), .A2(n9401), .ZN(n9405) );
  NAND2_X1 U6169 ( .A1(n9400), .A2(n4591), .ZN(n4590) );
  NAND2_X1 U6170 ( .A1(n9449), .A2(n10180), .ZN(n4884) );
  NAND2_X1 U6171 ( .A1(n4592), .A2(n9438), .ZN(n9445) );
  NAND2_X1 U6172 ( .A1(n9436), .A2(n9437), .ZN(n4592) );
  NAND2_X1 U6173 ( .A1(n4784), .A2(n9333), .ZN(n9324) );
  NAND2_X1 U6174 ( .A1(n4881), .A2(n4880), .ZN(P1_U3240) );
  NAND2_X1 U6175 ( .A1(n5079), .A2(n5081), .ZN(n9894) );
  XNOR2_X1 U6176 ( .A(n5134), .B(n5056), .ZN(n5133) );
  NAND2_X1 U6177 ( .A1(n5108), .A2(n5055), .ZN(n5134) );
  OR2_X2 U6178 ( .A1(n9015), .A2(n4912), .ZN(n4911) );
  NAND2_X1 U6179 ( .A1(n7179), .A2(n7178), .ZN(n7288) );
  NAND2_X1 U6180 ( .A1(n8116), .A2(n4932), .ZN(n4931) );
  OAI21_X2 U6181 ( .B1(n6515), .B2(P2_IR_REG_27__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U6182 ( .A1(n8139), .A2(n4735), .ZN(n4734) );
  AOI21_X1 U6183 ( .B1(n8143), .B2(n10406), .A(n8142), .ZN(n8484) );
  NAND2_X1 U6184 ( .A1(n8600), .A2(n6636), .ZN(n6642) );
  NOR2_X1 U6185 ( .A1(n6641), .A2(n5027), .ZN(n6648) );
  NAND2_X1 U6186 ( .A1(n6648), .A2(n6647), .ZN(n6650) );
  NAND2_X1 U6187 ( .A1(n4892), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4891) );
  NAND2_X1 U6188 ( .A1(n5601), .A2(n5600), .ZN(n5623) );
  NAND2_X1 U6189 ( .A1(n8489), .A2(n8140), .ZN(n8708) );
  NAND2_X1 U6190 ( .A1(n4877), .A2(n5673), .ZN(n5698) );
  AOI21_X2 U6191 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n10114), .A(n10109), .ZN(
        n10124) );
  AOI21_X2 U6192 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n10102), .A(n10097), .ZN(
        n6885) );
  AOI21_X2 U6193 ( .B1(n10127), .B2(P1_REG2_REG_13__SCAN_IN), .A(n10122), .ZN(
        n9506) );
  INV_X1 U6194 ( .A(n5975), .ZN(n5885) );
  NAND4_X1 U6195 ( .A1(n4606), .A2(n4605), .A3(n4604), .A4(n4603), .ZN(n5975)
         );
  NAND3_X1 U6196 ( .A1(n6412), .A2(n6410), .A3(n4614), .ZN(n4613) );
  NAND2_X1 U6197 ( .A1(n4613), .A2(n4548), .ZN(n6421) );
  NAND2_X1 U6198 ( .A1(n4627), .A2(n4628), .ZN(n6500) );
  NOR2_X1 U6199 ( .A1(n6497), .A2(n4618), .ZN(n4633) );
  NAND2_X1 U6200 ( .A1(n9131), .A2(n4638), .ZN(n4637) );
  OR2_X2 U6201 ( .A1(n4647), .A2(n4646), .ZN(n4643) );
  NAND3_X1 U6202 ( .A1(n9141), .A2(n5875), .A3(n9152), .ZN(n4649) );
  NAND3_X1 U6203 ( .A1(n4649), .A2(n4650), .A3(n4563), .ZN(P1_U3212) );
  NAND3_X1 U6204 ( .A1(n4660), .A2(n5364), .A3(n4658), .ZN(n7649) );
  NAND3_X1 U6205 ( .A1(n4944), .A2(n4662), .A3(n4661), .ZN(n4660) );
  NAND2_X1 U6206 ( .A1(n4666), .A2(n7829), .ZN(n5489) );
  NAND2_X1 U6207 ( .A1(n4666), .A2(n4665), .ZN(n9056) );
  NAND2_X1 U6208 ( .A1(n9102), .A2(n4486), .ZN(n4670) );
  OAI22_X1 U6209 ( .A1(n5115), .A2(n4672), .B1(n10185), .B2(n5793), .ZN(n4671)
         );
  NAND2_X2 U6210 ( .A1(n5068), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5098) );
  NAND4_X1 U6211 ( .A1(n5238), .A2(n5237), .A3(n4674), .A4(n4673), .ZN(n5036)
         );
  INV_X1 U6212 ( .A(n4679), .ZN(n7957) );
  INV_X1 U6213 ( .A(n4681), .ZN(n9601) );
  NAND3_X1 U6214 ( .A1(n9621), .A2(n9603), .A3(n4683), .ZN(n4682) );
  AND2_X1 U6215 ( .A1(n9587), .A2(n4688), .ZN(n9544) );
  NAND2_X1 U6216 ( .A1(n9587), .A2(n4687), .ZN(n9543) );
  NAND2_X1 U6217 ( .A1(n9587), .A2(n4490), .ZN(n9564) );
  AND2_X1 U6218 ( .A1(n9587), .A2(n9576), .ZN(n9571) );
  AND3_X2 U6219 ( .A1(n5062), .A2(n5060), .A3(n5061), .ZN(n10185) );
  NAND2_X1 U6220 ( .A1(n7238), .A2(n7237), .ZN(n7242) );
  NAND2_X1 U6221 ( .A1(n7118), .A2(n7119), .ZN(n7120) );
  NAND2_X1 U6222 ( .A1(n6845), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4695) );
  NAND2_X1 U6223 ( .A1(n4697), .A2(n6846), .ZN(n4696) );
  INV_X1 U6224 ( .A(n6845), .ZN(n4697) );
  NAND2_X1 U6225 ( .A1(n7713), .A2(n4712), .ZN(n4711) );
  AOI21_X1 U6226 ( .B1(n6078), .B2(n4717), .A(n4716), .ZN(n4715) );
  NAND2_X1 U6227 ( .A1(n6007), .A2(n4726), .ZN(n4725) );
  NAND2_X1 U6228 ( .A1(n8648), .A2(n7125), .ZN(n6353) );
  NAND2_X2 U6229 ( .A1(n6832), .A2(n5936), .ZN(n5960) );
  NAND2_X2 U6230 ( .A1(n5021), .A2(n4740), .ZN(n8538) );
  NAND2_X1 U6231 ( .A1(n9022), .A2(n4743), .ZN(n8910) );
  INV_X1 U6232 ( .A(n4745), .ZN(n7982) );
  INV_X1 U6233 ( .A(n8803), .ZN(n4748) );
  NOR2_X1 U6234 ( .A1(n8803), .A2(n4749), .ZN(n8794) );
  NOR2_X1 U6235 ( .A1(n8803), .A2(n8977), .ZN(n4750) );
  INV_X1 U6236 ( .A(n4750), .ZN(n8802) );
  NAND2_X1 U6237 ( .A1(n7390), .A2(n7218), .ZN(n9302) );
  NAND2_X1 U6238 ( .A1(n9216), .A2(n9259), .ZN(n7390) );
  NAND2_X1 U6239 ( .A1(n7216), .A2(n7215), .ZN(n9216) );
  INV_X1 U6241 ( .A(n9638), .ZN(n4756) );
  NAND2_X1 U6242 ( .A1(n8082), .A2(n4487), .ZN(n4757) );
  NAND2_X1 U6243 ( .A1(n4757), .A2(n4758), .ZN(n9700) );
  NAND2_X1 U6244 ( .A1(n4772), .A2(n4494), .ZN(n4771) );
  NAND2_X1 U6245 ( .A1(n4774), .A2(n4773), .ZN(n8106) );
  AOI21_X1 U6246 ( .B1(n4780), .B2(n4782), .A(n4781), .ZN(n4778) );
  INV_X1 U6247 ( .A(n4780), .ZN(n4779) );
  AOI21_X1 U6248 ( .B1(n9593), .B2(n4788), .A(n4786), .ZN(n8093) );
  NAND2_X1 U6249 ( .A1(n9593), .A2(n4512), .ZN(n4789) );
  NAND2_X1 U6250 ( .A1(n9593), .A2(n9594), .ZN(n9592) );
  OAI21_X1 U6251 ( .B1(n9932), .B2(n4794), .A(n4546), .ZN(n7939) );
  OR2_X1 U6252 ( .A1(n6777), .A2(n6808), .ZN(n5060) );
  NAND2_X1 U6253 ( .A1(n7586), .A2(n4804), .ZN(n4801) );
  NAND2_X1 U6254 ( .A1(n4801), .A2(n4802), .ZN(n7769) );
  AOI21_X2 U6255 ( .B1(n4822), .B2(n5033), .A(n4821), .ZN(n4820) );
  NAND2_X1 U6256 ( .A1(n7100), .A2(n4517), .ZN(n7383) );
  OAI21_X2 U6257 ( .B1(n6595), .B2(n4827), .A(n4825), .ZN(n8024) );
  NAND2_X2 U6258 ( .A1(n7504), .A2(n6691), .ZN(n4832) );
  XNOR2_X2 U6259 ( .A(n4833), .B(n5892), .ZN(n7504) );
  NAND2_X1 U6260 ( .A1(n4836), .A2(n5290), .ZN(n5315) );
  NAND2_X1 U6261 ( .A1(n4837), .A2(n4562), .ZN(n5650) );
  INV_X1 U6262 ( .A(n5596), .ZN(n5599) );
  NAND2_X1 U6263 ( .A1(n6287), .A2(n4845), .ZN(n4842) );
  NAND2_X1 U6264 ( .A1(n4842), .A2(n4843), .ZN(n6319) );
  NAND2_X1 U6265 ( .A1(n5448), .A2(n4852), .ZN(n4851) );
  NAND2_X1 U6266 ( .A1(n4860), .A2(n9170), .ZN(n9783) );
  NAND2_X1 U6267 ( .A1(n5343), .A2(n4862), .ZN(n4861) );
  NAND2_X1 U6268 ( .A1(n4861), .A2(n4864), .ZN(n5423) );
  NAND2_X1 U6269 ( .A1(n5675), .A2(n4496), .ZN(n4871) );
  OR2_X1 U6270 ( .A1(n5675), .A2(n5674), .ZN(n4877) );
  NAND3_X1 U6271 ( .A1(n4886), .A2(n4885), .A3(n4884), .ZN(n4883) );
  NOR2_X2 U6272 ( .A1(n9455), .A2(n7467), .ZN(n4885) );
  NAND2_X1 U6273 ( .A1(n5052), .A2(n4890), .ZN(n4889) );
  INV_X1 U6274 ( .A(n4893), .ZN(n4892) );
  NAND2_X1 U6275 ( .A1(n4894), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U6276 ( .A1(n4894), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U6277 ( .A1(n4894), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U6278 ( .A1(n4894), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U6279 ( .A1(n4894), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U6280 ( .A1(n4894), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6133) );
  NAND2_X1 U6281 ( .A1(n4894), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6186) );
  NAND2_X1 U6282 ( .A1(n4894), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U6283 ( .A1(n4894), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6203) );
  NAND2_X1 U6284 ( .A1(n4894), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U6285 ( .A1(n4894), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U6286 ( .A1(n4894), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U6287 ( .A1(n4894), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U6288 ( .A1(n6365), .A2(n4895), .ZN(n6366) );
  NAND3_X1 U6289 ( .A1(n5899), .A2(n5900), .A3(n5902), .ZN(n5907) );
  NAND2_X1 U6290 ( .A1(n7633), .A2(n4899), .ZN(n7676) );
  INV_X1 U6291 ( .A(n8801), .ZN(n4901) );
  NAND2_X1 U6292 ( .A1(n4904), .A2(n4902), .ZN(n8768) );
  AND2_X2 U6293 ( .A1(n4911), .A2(n4909), .ZN(n8844) );
  AND2_X1 U6294 ( .A1(n9010), .A2(n8931), .ZN(n4916) );
  NAND2_X1 U6295 ( .A1(n8753), .A2(n4920), .ZN(n4917) );
  NAND2_X1 U6296 ( .A1(n4917), .A2(n4918), .ZN(n8488) );
  NAND2_X1 U6297 ( .A1(n8765), .A2(n8777), .ZN(n4926) );
  NAND2_X1 U6298 ( .A1(n5910), .A2(n5909), .ZN(n6515) );
  NAND2_X1 U6299 ( .A1(n8116), .A2(n4483), .ZN(n9974) );
  INV_X1 U6300 ( .A(n8116), .ZN(n4936) );
  NAND2_X1 U6301 ( .A1(n5285), .A2(n4945), .ZN(n4944) );
  NOR2_X1 U6302 ( .A1(n9087), .A2(n9086), .ZN(n9085) );
  INV_X1 U6303 ( .A(n9087), .ZN(n4953) );
  NOR2_X1 U6304 ( .A1(n9085), .A2(n5771), .ZN(n9141) );
  XNOR2_X1 U6305 ( .A(n4956), .B(n5814), .ZN(n5146) );
  NAND2_X1 U6306 ( .A1(n9894), .A2(n4542), .ZN(n4963) );
  INV_X1 U6307 ( .A(n9707), .ZN(n4972) );
  NAND2_X1 U6308 ( .A1(n9553), .A2(n4975), .ZN(n4976) );
  NAND3_X1 U6309 ( .A1(n4977), .A2(n4979), .A3(n4976), .ZN(n9790) );
  NAND3_X1 U6310 ( .A1(n4977), .A2(n4495), .A3(n4976), .ZN(n4980) );
  NAND2_X1 U6311 ( .A1(n9551), .A2(n4978), .ZN(n4977) );
  NAND3_X1 U6312 ( .A1(n9789), .A2(n9788), .A3(n4980), .ZN(n9877) );
  NAND2_X1 U6313 ( .A1(n7407), .A2(n4984), .ZN(n4983) );
  NAND2_X1 U6314 ( .A1(n4983), .A2(n4982), .ZN(n7410) );
  NAND2_X1 U6315 ( .A1(n8070), .A2(n4990), .ZN(n4989) );
  NAND2_X1 U6316 ( .A1(n7617), .A2(n4485), .ZN(n5003) );
  NAND2_X1 U6317 ( .A1(n8064), .A2(n4544), .ZN(n5007) );
  OR2_X1 U6318 ( .A1(n9858), .A2(n9470), .ZN(n5017) );
  AOI21_X1 U6319 ( .B1(n8503), .B2(n6690), .A(n5024), .ZN(n6694) );
  NAND2_X1 U6320 ( .A1(n8503), .A2(n8502), .ZN(n8501) );
  OR2_X1 U6321 ( .A1(n6635), .A2(n6634), .ZN(n6636) );
  INV_X1 U6322 ( .A(n8510), .ZN(n6646) );
  XNOR2_X1 U6323 ( .A(n5776), .B(n5775), .ZN(n7920) );
  INV_X1 U6324 ( .A(n6962), .ZN(n5113) );
  NAND2_X1 U6325 ( .A1(n5203), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U6326 ( .A1(n5113), .A2(n7361), .ZN(n5120) );
  NAND2_X1 U6327 ( .A1(n5122), .A2(n5121), .ZN(n8035) );
  NAND2_X1 U6328 ( .A1(n5120), .A2(n5119), .ZN(n5121) );
  OAI21_X1 U6329 ( .B1(n5748), .B2(n5747), .A(n5746), .ZN(n5776) );
  XNOR2_X1 U6330 ( .A(n5748), .B(n5747), .ZN(n7914) );
  NAND2_X1 U6331 ( .A1(n8081), .A2(n9377), .ZN(n8082) );
  NAND2_X1 U6332 ( .A1(n8091), .A2(n9414), .ZN(n9593) );
  NAND2_X1 U6333 ( .A1(n8083), .A2(n9396), .ZN(n9678) );
  OR2_X1 U6334 ( .A1(n5913), .A2(n6083), .ZN(n5915) );
  INV_X1 U6335 ( .A(n9678), .ZN(n8085) );
  OR2_X1 U6336 ( .A1(n5954), .A2(n5930), .ZN(n5935) );
  NAND2_X1 U6337 ( .A1(n5951), .A2(n5950), .ZN(n7085) );
  INV_X1 U6338 ( .A(n9261), .ZN(n7158) );
  NAND2_X1 U6339 ( .A1(n8085), .A2(n8084), .ZN(n9662) );
  INV_X1 U6340 ( .A(n5952), .ZN(n5969) );
  OR2_X1 U6341 ( .A1(n5952), .A2(n5931), .ZN(n5934) );
  OR2_X1 U6342 ( .A1(n5952), .A2(n5918), .ZN(n5922) );
  NAND2_X1 U6343 ( .A1(n5080), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5082) );
  NAND2_X1 U6344 ( .A1(n7153), .A2(n5795), .ZN(n5112) );
  OR2_X1 U6345 ( .A1(n6832), .A2(n6718), .ZN(n5021) );
  INV_X1 U6346 ( .A(n8824), .ZN(n6206) );
  NAND2_X1 U6347 ( .A1(n7211), .A2(n7210), .ZN(n7218) );
  OR2_X1 U6348 ( .A1(n8847), .A2(n8613), .ZN(n5022) );
  AND4_X1 U6349 ( .A1(n6002), .A2(n5884), .A3(n5883), .A4(n5882), .ZN(n5023)
         );
  NOR2_X1 U6350 ( .A1(n6689), .A2(n6688), .ZN(n5024) );
  AND2_X1 U6351 ( .A1(n9576), .A2(n9557), .ZN(n5025) );
  AND2_X1 U6352 ( .A1(n5475), .A2(n5094), .ZN(n5026) );
  AND2_X1 U6353 ( .A1(n6640), .A2(n8583), .ZN(n5027) );
  AND2_X1 U6354 ( .A1(n5342), .A2(n5322), .ZN(n5028) );
  OR2_X1 U6355 ( .A1(n8495), .A2(n8614), .ZN(n5029) );
  AND2_X1 U6356 ( .A1(n5367), .A2(n5347), .ZN(n5030) );
  AND2_X1 U6357 ( .A1(n5447), .A2(n5426), .ZN(n5031) );
  INV_X1 U6358 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n8328) );
  AND4_X1 U6359 ( .A1(n6174), .A2(n6173), .A3(n6172), .A4(n6171), .ZN(n8887)
         );
  INV_X1 U6360 ( .A(n8887), .ZN(n8119) );
  AND4_X1 U6361 ( .A1(n5810), .A2(n5809), .A3(n5808), .A4(n5807), .ZN(n9580)
         );
  INV_X4 U6362 ( .A(n6723), .ZN(n6724) );
  INV_X1 U6363 ( .A(n7641), .ZN(n7565) );
  INV_X1 U6364 ( .A(n9395), .ZN(n8084) );
  AND2_X1 U6365 ( .A1(n10187), .A2(n5843), .ZN(n9151) );
  INV_X1 U6366 ( .A(n9151), .ZN(n9165) );
  AND2_X1 U6367 ( .A1(n5774), .A2(n5773), .ZN(n5874) );
  AND2_X1 U6368 ( .A1(n8644), .A2(n10346), .ZN(n5034) );
  INV_X1 U6369 ( .A(n9266), .ZN(n7616) );
  INV_X1 U6370 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5041) );
  INV_X1 U6371 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U6372 ( .A1(n6497), .A2(n6465), .ZN(n6466) );
  INV_X1 U6373 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5902) );
  INV_X1 U6374 ( .A(n10205), .ZN(n7210) );
  INV_X1 U6375 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6047) );
  INV_X1 U6376 ( .A(n6010), .ZN(n6008) );
  INV_X1 U6377 ( .A(n6242), .ZN(n6241) );
  INV_X1 U6378 ( .A(n6230), .ZN(n6229) );
  INV_X1 U6379 ( .A(n6113), .ZN(n6112) );
  NAND2_X1 U6380 ( .A1(n6530), .A2(n8538), .ZN(n6475) );
  INV_X1 U6381 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6106) );
  INV_X1 U6382 ( .A(n7056), .ZN(n5198) );
  NOR2_X1 U6383 ( .A1(n5877), .A2(n5785), .ZN(n5805) );
  INV_X1 U6384 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5258) );
  INV_X1 U6385 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5048) );
  INV_X1 U6386 ( .A(n5286), .ZN(n5287) );
  NAND2_X1 U6387 ( .A1(n6008), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U6388 ( .A1(n6200), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U6389 ( .A1(n6087), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6099) );
  NOR2_X1 U6390 ( .A1(n7298), .A2(n6570), .ZN(n6536) );
  OR2_X1 U6391 ( .A1(n6278), .A2(n6703), .ZN(n8714) );
  OR2_X1 U6392 ( .A1(n6209), .A2(n8604), .ZN(n6221) );
  OR2_X1 U6393 ( .A1(n7233), .A2(n7232), .ZN(n7542) );
  NAND2_X1 U6394 ( .A1(n6069), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6088) );
  OR2_X1 U6395 ( .A1(n6040), .A2(n6039), .ZN(n6056) );
  NAND2_X1 U6396 ( .A1(n6356), .A2(n6476), .ZN(n7087) );
  INV_X1 U6397 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U6398 ( .A1(n9153), .A2(n9157), .ZN(n9093) );
  INV_X1 U6399 ( .A(n7796), .ZN(n5419) );
  OR2_X1 U6400 ( .A1(n5528), .A2(n8398), .ZN(n5555) );
  OR2_X1 U6401 ( .A1(n5432), .A2(n5431), .ZN(n5455) );
  INV_X1 U6402 ( .A(n9580), .ZN(n8072) );
  NAND2_X1 U6403 ( .A1(n5509), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5528) );
  OR2_X1 U6404 ( .A1(n5352), .A2(n6887), .ZN(n5377) );
  NAND2_X1 U6405 ( .A1(n5472), .A2(n5471), .ZN(n5497) );
  NAND2_X1 U6406 ( .A1(n5397), .A2(n5396), .ZN(n5421) );
  NAND2_X1 U6407 ( .A1(n8581), .A2(n6644), .ZN(n8510) );
  NOR2_X1 U6408 ( .A1(n7021), .A2(n6548), .ZN(n6549) );
  NOR2_X1 U6409 ( .A1(n6654), .A2(n6653), .ZN(n6655) );
  OR2_X1 U6410 ( .A1(n8504), .A2(n6266), .ZN(n6272) );
  INV_X1 U6411 ( .A(n8945), .ZN(n8709) );
  OR2_X1 U6412 ( .A1(n9005), .A2(n8903), .ZN(n8118) );
  INV_X1 U6413 ( .A(n7285), .ZN(n7292) );
  AND2_X1 U6414 ( .A1(n6334), .A2(n8880), .ZN(n8905) );
  NAND2_X1 U6415 ( .A1(n8109), .A2(n8107), .ZN(n7296) );
  NAND2_X1 U6416 ( .A1(n5608), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5627) );
  INV_X1 U6417 ( .A(n9767), .ZN(n9162) );
  OR2_X1 U6418 ( .A1(n9868), .A2(n9453), .ZN(n7149) );
  OR2_X1 U6419 ( .A1(n9440), .A2(n9456), .ZN(n9868) );
  INV_X1 U6420 ( .A(n8930), .ZN(n8886) );
  AND2_X1 U6421 ( .A1(n6834), .A2(n6833), .ZN(n10258) );
  AND2_X1 U6422 ( .A1(n10287), .A2(n9978), .ZN(n8936) );
  AND2_X1 U6423 ( .A1(n6523), .A2(n7078), .ZN(n8928) );
  AND2_X1 U6424 ( .A1(n8915), .A2(n10272), .ZN(n10284) );
  AND2_X1 U6425 ( .A1(n7096), .A2(n7095), .ZN(n7196) );
  NAND2_X1 U6426 ( .A1(n6701), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10294) );
  INV_X1 U6427 ( .A(n9141), .ZN(n9145) );
  AND2_X1 U6428 ( .A1(n5635), .A2(n5634), .ZN(n9682) );
  NAND2_X1 U6429 ( .A1(n9426), .A2(n9238), .ZN(n9552) );
  NAND2_X1 U6430 ( .A1(n9415), .A2(n9414), .ZN(n9609) );
  AOI22_X1 U6431 ( .A1(n9659), .A2(n9660), .B1(n9653), .B2(n9827), .ZN(n9646)
         );
  AND2_X1 U6432 ( .A1(n9392), .A2(n9396), .ZN(n9699) );
  AND2_X1 U6433 ( .A1(n9761), .A2(n9190), .ZN(n9275) );
  AND2_X1 U6434 ( .A1(n5853), .A2(n9446), .ZN(n9935) );
  NAND2_X1 U6435 ( .A1(n5842), .A2(n6956), .ZN(n10187) );
  AND2_X1 U6436 ( .A1(n9757), .A2(n9868), .ZN(n9866) );
  AND2_X1 U6437 ( .A1(n7743), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6740) );
  AND2_X1 U6438 ( .A1(n6710), .A2(n6740), .ZN(n6956) );
  OR2_X1 U6439 ( .A1(n6521), .A2(n7805), .ZN(n6828) );
  AND2_X1 U6440 ( .A1(n6706), .A2(n5029), .ZN(n6707) );
  OR2_X1 U6441 ( .A1(n8560), .A2(n8886), .ZN(n8614) );
  OR2_X1 U6442 ( .A1(n6526), .A2(n6525), .ZN(n6527) );
  AND2_X1 U6443 ( .A1(n6249), .A2(n6248), .ZN(n8777) );
  AND4_X1 U6444 ( .A1(n6104), .A2(n6103), .A3(n6102), .A4(n6101), .ZN(n8115)
         );
  INV_X1 U6445 ( .A(n7644), .ZN(n8642) );
  INV_X1 U6446 ( .A(n9921), .ZN(n10261) );
  INV_X1 U6447 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8706) );
  INV_X1 U6448 ( .A(n10395), .ZN(n10393) );
  CLKBUF_X1 U6449 ( .A(n10308), .Z(n10331) );
  INV_X1 U6450 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n8312) );
  INV_X1 U6451 ( .A(n9152), .ZN(n9139) );
  INV_X1 U6452 ( .A(n10041), .ZN(n10175) );
  AND2_X2 U6453 ( .A1(n7411), .A2(n10187), .ZN(n10193) );
  INV_X1 U6454 ( .A(n10255), .ZN(n10256) );
  NAND2_X1 U6455 ( .A1(n7310), .A2(n6994), .ZN(n10245) );
  INV_X1 U6456 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8288) );
  INV_X1 U6457 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8170) );
  XNOR2_X1 U6458 ( .A(n5268), .B(n5267), .ZN(n6738) );
  NOR2_X1 U6459 ( .A1(n10440), .A2(n10439), .ZN(n10438) );
  NOR2_X1 U6460 ( .A1(n10437), .A2(n10436), .ZN(n10435) );
  NOR2_X2 U6461 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5137) );
  NAND2_X1 U6462 ( .A1(n5137), .A2(n5035), .ZN(n5188) );
  NOR2_X2 U6463 ( .A1(n5188), .A2(n5036), .ZN(n5295) );
  NAND2_X1 U6464 ( .A1(n5295), .A2(n5296), .ZN(n5091) );
  NOR2_X1 U6465 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5040) );
  NOR2_X1 U6466 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5039) );
  INV_X1 U6467 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5045) );
  NAND2_X1 U6468 ( .A1(n5045), .A2(n5097), .ZN(n5069) );
  INV_X1 U6469 ( .A(n5069), .ZN(n5047) );
  NOR2_X1 U6470 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5046) );
  NAND2_X1 U6471 ( .A1(n5049), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5050) );
  INV_X1 U6472 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5077) );
  XNOR2_X1 U6473 ( .A(n5050), .B(n5077), .ZN(n5853) );
  INV_X1 U6474 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5051) );
  INV_X1 U6475 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6726) );
  NAND3_X1 U6476 ( .A1(n5053), .A2(P1_DATAO_REG_0__SCAN_IN), .A3(SI_0_), .ZN(
        n5055) );
  AND2_X1 U6477 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5054) );
  NAND2_X1 U6478 ( .A1(n5057), .A2(n5054), .ZN(n5108) );
  INV_X1 U6479 ( .A(SI_1_), .ZN(n5056) );
  MUX2_X1 U6480 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5057), .Z(n5132) );
  XNOR2_X1 U6481 ( .A(n5133), .B(n5132), .ZN(n6725) );
  OR2_X1 U6482 ( .A1(n5273), .A2(n6725), .ZN(n5061) );
  INV_X1 U6483 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U6484 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n6791), .ZN(n5058) );
  NAND2_X1 U6485 ( .A1(n4535), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5064) );
  XNOR2_X1 U6486 ( .A(n5064), .B(n5063), .ZN(n7917) );
  NAND2_X1 U6487 ( .A1(n5065), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5067) );
  INV_X1 U6488 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5066) );
  XNOR2_X1 U6489 ( .A(n5067), .B(n5066), .ZN(n7922) );
  NAND2_X1 U6490 ( .A1(n5069), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5070) );
  NAND2_X1 U6491 ( .A1(n5098), .A2(n5070), .ZN(n5820) );
  OAI21_X2 U6492 ( .B1(n5820), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5072) );
  INV_X1 U6493 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5071) );
  XNOR2_X1 U6494 ( .A(n5098), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9453) );
  INV_X1 U6495 ( .A(n5073), .ZN(n5074) );
  NAND2_X1 U6496 ( .A1(n5074), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5076) );
  XNOR2_X1 U6497 ( .A(n5076), .B(n5075), .ZN(n7467) );
  NAND2_X1 U6498 ( .A1(n5078), .A2(n5077), .ZN(n5080) );
  INV_X1 U6499 ( .A(n5080), .ZN(n5079) );
  INV_X1 U6500 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9895) );
  XNOR2_X2 U6501 ( .A(n5082), .B(n5081), .ZN(n9903) );
  NAND2_X1 U6502 ( .A1(n8101), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5085) );
  AND2_X1 U6503 ( .A1(n5085), .A2(n5084), .ZN(n5089) );
  NAND2_X1 U6504 ( .A1(n8500), .A2(n9903), .ZN(n5175) );
  NAND2_X1 U6505 ( .A1(n8100), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5088) );
  INV_X1 U6506 ( .A(n10178), .ZN(n5090) );
  AND2_X4 U6507 ( .A1(n6710), .A2(n5090), .ZN(n5795) );
  INV_X1 U6508 ( .A(n5795), .ZN(n5115) );
  BUF_X1 U6509 ( .A(n5091), .Z(n5298) );
  INV_X1 U6510 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5369) );
  NAND2_X1 U6511 ( .A1(n5369), .A2(n5092), .ZN(n5093) );
  NAND2_X1 U6512 ( .A1(n5400), .A2(n5401), .ZN(n5427) );
  INV_X1 U6513 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5475) );
  INV_X1 U6514 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U6515 ( .A1(n5449), .A2(n5026), .ZN(n5505) );
  OAI21_X2 U6516 ( .B1(n5505), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5549) );
  OAI21_X1 U6517 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6518 ( .A1(n5549), .A2(n5095), .ZN(n5096) );
  XNOR2_X2 U6519 ( .A(n5096), .B(P1_IR_REG_19__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U6520 ( .A1(n5098), .A2(n5097), .ZN(n5099) );
  NAND2_X1 U6521 ( .A1(n5099), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5100) );
  XNOR2_X1 U6522 ( .A(n5100), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9462) );
  NAND2_X1 U6523 ( .A1(n5578), .A2(n9462), .ZN(n5101) );
  AND2_X4 U6524 ( .A1(n5101), .A2(n10178), .ZN(n7361) );
  NAND2_X1 U6525 ( .A1(n8100), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5105) );
  INV_X1 U6526 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6775) );
  OR2_X1 U6527 ( .A1(n5738), .A2(n6775), .ZN(n5104) );
  INV_X1 U6528 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8337) );
  OR2_X1 U6529 ( .A1(n5806), .A2(n8337), .ZN(n5103) );
  INV_X1 U6530 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6965) );
  NAND2_X1 U6531 ( .A1(n6724), .A2(SI_0_), .ZN(n5107) );
  INV_X1 U6532 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U6533 ( .A1(n5107), .A2(n5106), .ZN(n5109) );
  AND2_X1 U6534 ( .A1(n5108), .A2(n5109), .ZN(n6716) );
  MUX2_X1 U6535 ( .A(n6791), .B(n6716), .S(n6777), .Z(n7165) );
  NOR2_X1 U6536 ( .A1(n6710), .A2(n6775), .ZN(n5110) );
  AOI21_X1 U6537 ( .B1(n7165), .B2(n5817), .A(n5110), .ZN(n5111) );
  NAND2_X1 U6538 ( .A1(n5112), .A2(n5111), .ZN(n6962) );
  NAND2_X1 U6539 ( .A1(n5578), .A2(n7467), .ZN(n7312) );
  OR2_X1 U6540 ( .A1(n7312), .A2(n9462), .ZN(n5114) );
  NAND2_X1 U6541 ( .A1(n7153), .A2(n5145), .ZN(n5118) );
  INV_X1 U6542 ( .A(n6791), .ZN(n6773) );
  NOR2_X1 U6543 ( .A1(n6710), .A2(n6773), .ZN(n5116) );
  AOI21_X1 U6544 ( .B1(n7165), .B2(n5816), .A(n5116), .ZN(n5117) );
  NAND2_X1 U6545 ( .A1(n5118), .A2(n5117), .ZN(n6961) );
  NAND2_X1 U6546 ( .A1(n6962), .A2(n6961), .ZN(n5119) );
  AOI22_X1 U6547 ( .A1(n9480), .A2(n5145), .B1(n8039), .B2(n5816), .ZN(n8037)
         );
  NAND2_X1 U6548 ( .A1(n8035), .A2(n8037), .ZN(n5125) );
  INV_X1 U6549 ( .A(n5121), .ZN(n5124) );
  INV_X1 U6550 ( .A(n5122), .ZN(n5123) );
  NAND2_X1 U6551 ( .A1(n5124), .A2(n5123), .ZN(n8036) );
  NAND2_X1 U6552 ( .A1(n5125), .A2(n8036), .ZN(n7000) );
  INV_X1 U6553 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5126) );
  INV_X1 U6554 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5127) );
  NAND2_X1 U6555 ( .A1(n5203), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U6556 ( .A1(n8101), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5128) );
  NAND4_X2 U6557 ( .A1(n5131), .A2(n5130), .A3(n5129), .A4(n5128), .ZN(n9478)
         );
  NAND2_X1 U6558 ( .A1(n9478), .A2(n5795), .ZN(n5144) );
  NAND2_X1 U6559 ( .A1(n5133), .A2(n5132), .ZN(n5136) );
  NAND2_X1 U6560 ( .A1(n5134), .A2(SI_1_), .ZN(n5135) );
  INV_X1 U6561 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6720) );
  INV_X1 U6562 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6728) );
  MUX2_X1 U6563 ( .A(n6720), .B(n6728), .S(n5057), .Z(n5157) );
  XNOR2_X1 U6564 ( .A(n5157), .B(SI_2_), .ZN(n5155) );
  XNOR2_X1 U6565 ( .A(n5156), .B(n5155), .ZN(n6727) );
  OR2_X1 U6566 ( .A1(n5273), .A2(n6727), .ZN(n5143) );
  OR2_X1 U6567 ( .A1(n9173), .A2(n6728), .ZN(n5142) );
  OR2_X1 U6568 ( .A1(n5137), .A2(n5051), .ZN(n5139) );
  INV_X1 U6569 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U6570 ( .A1(n5139), .A2(n5138), .ZN(n5161) );
  OAI21_X1 U6571 ( .B1(n5139), .B2(n5138), .A(n5161), .ZN(n7044) );
  OR2_X1 U6572 ( .A1(n5140), .A2(n7044), .ZN(n5141) );
  AOI22_X1 U6573 ( .A1(n9478), .A2(n5145), .B1(n7210), .B2(n5816), .ZN(n5147)
         );
  XNOR2_X1 U6574 ( .A(n5146), .B(n5147), .ZN(n7001) );
  NAND2_X1 U6575 ( .A1(n7000), .A2(n7001), .ZN(n5150) );
  INV_X1 U6576 ( .A(n5146), .ZN(n5148) );
  NAND2_X1 U6577 ( .A1(n5148), .A2(n5147), .ZN(n5149) );
  NAND2_X1 U6578 ( .A1(n5755), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5154) );
  INV_X1 U6579 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6797) );
  OR2_X1 U6580 ( .A1(n5738), .A2(n6797), .ZN(n5153) );
  INV_X1 U6581 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6811) );
  OR2_X1 U6582 ( .A1(n5806), .A2(n6811), .ZN(n5152) );
  NAND2_X1 U6583 ( .A1(n9477), .A2(n5795), .ZN(n5168) );
  INV_X1 U6584 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8332) );
  INV_X1 U6585 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6730) );
  MUX2_X1 U6586 ( .A(n8332), .B(n6730), .S(n5057), .Z(n5183) );
  XNOR2_X1 U6587 ( .A(n5183), .B(SI_3_), .ZN(n5181) );
  NAND2_X1 U6588 ( .A1(n5156), .A2(n5155), .ZN(n5160) );
  INV_X1 U6589 ( .A(n5157), .ZN(n5158) );
  NAND2_X1 U6590 ( .A1(n5158), .A2(SI_2_), .ZN(n5159) );
  NAND2_X1 U6591 ( .A1(n5160), .A2(n5159), .ZN(n5182) );
  XNOR2_X1 U6592 ( .A(n5182), .B(n5181), .ZN(n6729) );
  OR2_X1 U6593 ( .A1(n5273), .A2(n6729), .ZN(n5166) );
  OR2_X1 U6594 ( .A1(n9173), .A2(n6730), .ZN(n5165) );
  NAND2_X1 U6595 ( .A1(n5161), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5163) );
  INV_X1 U6596 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5162) );
  OR2_X1 U6597 ( .A1(n6777), .A2(n9483), .ZN(n5164) );
  OR2_X1 U6598 ( .A1(n7322), .A2(n5793), .ZN(n5167) );
  NAND2_X1 U6599 ( .A1(n5168), .A2(n5167), .ZN(n5169) );
  XNOR2_X1 U6600 ( .A(n5169), .B(n5814), .ZN(n5170) );
  INV_X1 U6601 ( .A(n7322), .ZN(n7356) );
  AOI22_X1 U6602 ( .A1(n9477), .A2(n5145), .B1(n7356), .B2(n5816), .ZN(n5171)
         );
  XNOR2_X1 U6603 ( .A(n5170), .B(n5171), .ZN(n7010) );
  INV_X1 U6604 ( .A(n5170), .ZN(n5172) );
  NAND2_X1 U6605 ( .A1(n5172), .A2(n5171), .ZN(n5173) );
  INV_X2 U6606 ( .A(n5738), .ZN(n8101) );
  NAND2_X1 U6607 ( .A1(n8101), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5180) );
  INV_X1 U6608 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5176) );
  OR2_X1 U6609 ( .A1(n5175), .A2(n5176), .ZN(n5179) );
  XNOR2_X1 U6610 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7474) );
  OR2_X1 U6611 ( .A1(n5856), .A2(n7474), .ZN(n5178) );
  INV_X1 U6612 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6813) );
  OR2_X1 U6613 ( .A1(n5806), .A2(n6813), .ZN(n5177) );
  NAND2_X1 U6614 ( .A1(n9476), .A2(n5795), .ZN(n5196) );
  NAND2_X1 U6615 ( .A1(n5182), .A2(n5181), .ZN(n5186) );
  INV_X1 U6616 ( .A(n5183), .ZN(n5184) );
  NAND2_X1 U6617 ( .A1(n5184), .A2(SI_3_), .ZN(n5185) );
  NAND2_X1 U6618 ( .A1(n5186), .A2(n5185), .ZN(n5212) );
  XNOR2_X1 U6619 ( .A(n5213), .B(SI_4_), .ZN(n5211) );
  XNOR2_X1 U6620 ( .A(n5211), .B(n5212), .ZN(n6731) );
  OR2_X1 U6621 ( .A1(n5273), .A2(n6731), .ZN(n5194) );
  OR2_X1 U6622 ( .A1(n9173), .A2(n6732), .ZN(n5193) );
  NOR2_X1 U6623 ( .A1(n5188), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5239) );
  INV_X1 U6624 ( .A(n5239), .ZN(n5191) );
  NAND2_X1 U6625 ( .A1(n5188), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5189) );
  MUX2_X1 U6626 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5189), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5190) );
  NAND2_X1 U6627 ( .A1(n5191), .A2(n5190), .ZN(n10032) );
  OR2_X1 U6628 ( .A1(n6777), .A2(n10032), .ZN(n5192) );
  OR2_X1 U6629 ( .A1(n10210), .A2(n5793), .ZN(n5195) );
  NAND2_X1 U6630 ( .A1(n5196), .A2(n5195), .ZN(n5197) );
  XNOR2_X1 U6631 ( .A(n5197), .B(n7361), .ZN(n5200) );
  AOI22_X1 U6632 ( .A1(n9476), .A2(n5145), .B1(n7476), .B2(n5816), .ZN(n5199)
         );
  XNOR2_X1 U6633 ( .A(n5200), .B(n5199), .ZN(n7056) );
  OR2_X1 U6634 ( .A1(n5200), .A2(n5199), .ZN(n5201) );
  AOI21_X1 U6635 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5202) );
  NOR2_X1 U6636 ( .A1(n5202), .A2(n5226), .ZN(n7369) );
  NAND2_X1 U6637 ( .A1(n5203), .A2(n7369), .ZN(n5210) );
  INV_X1 U6638 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5204) );
  OR2_X1 U6639 ( .A1(n5738), .A2(n5204), .ZN(n5209) );
  INV_X1 U6640 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5205) );
  OR2_X1 U6641 ( .A1(n5175), .A2(n5205), .ZN(n5208) );
  INV_X1 U6642 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5206) );
  OR2_X1 U6643 ( .A1(n5806), .A2(n5206), .ZN(n5207) );
  NAND2_X1 U6644 ( .A1(n9475), .A2(n5795), .ZN(n5222) );
  NAND2_X1 U6645 ( .A1(n5212), .A2(n5211), .ZN(n5216) );
  INV_X1 U6646 ( .A(n5213), .ZN(n5214) );
  NAND2_X1 U6647 ( .A1(n5214), .A2(SI_4_), .ZN(n5215) );
  NAND2_X1 U6648 ( .A1(n5216), .A2(n5215), .ZN(n5232) );
  INV_X1 U6649 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6721) );
  INV_X1 U6650 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6735) );
  XNOR2_X1 U6651 ( .A(n5232), .B(n5231), .ZN(n6734) );
  OR2_X1 U6652 ( .A1(n5273), .A2(n6734), .ZN(n5220) );
  OR2_X1 U6653 ( .A1(n9173), .A2(n6735), .ZN(n5219) );
  OR2_X1 U6654 ( .A1(n5239), .A2(n5051), .ZN(n5217) );
  XNOR2_X1 U6655 ( .A(n5217), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10051) );
  INV_X1 U6656 ( .A(n10051), .ZN(n6733) );
  OR2_X1 U6657 ( .A1(n6777), .A2(n6733), .ZN(n5218) );
  OR2_X1 U6658 ( .A1(n10217), .A2(n5793), .ZN(n5221) );
  NAND2_X1 U6659 ( .A1(n5222), .A2(n5221), .ZN(n5223) );
  XNOR2_X1 U6660 ( .A(n5223), .B(n7361), .ZN(n7330) );
  NAND2_X1 U6661 ( .A1(n9475), .A2(n5145), .ZN(n5225) );
  OR2_X1 U6662 ( .A1(n10217), .A2(n5302), .ZN(n5224) );
  AND2_X1 U6663 ( .A1(n5225), .A2(n5224), .ZN(n7332) );
  NAND2_X1 U6664 ( .A1(n5755), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5230) );
  INV_X1 U6665 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6801) );
  OR2_X1 U6666 ( .A1(n5738), .A2(n6801), .ZN(n5229) );
  OAI21_X1 U6667 ( .B1(n5226), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5259), .ZN(
        n7491) );
  OR2_X1 U6668 ( .A1(n5856), .A2(n7491), .ZN(n5228) );
  INV_X1 U6669 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7492) );
  OR2_X1 U6670 ( .A1(n5806), .A2(n7492), .ZN(n5227) );
  NAND4_X1 U6671 ( .A1(n5230), .A2(n5229), .A3(n5228), .A4(n5227), .ZN(n9474)
         );
  NAND2_X1 U6672 ( .A1(n9474), .A2(n5795), .ZN(n5245) );
  NAND2_X1 U6673 ( .A1(n5232), .A2(n5231), .ZN(n5236) );
  INV_X1 U6674 ( .A(n5233), .ZN(n5234) );
  NAND2_X1 U6675 ( .A1(n5234), .A2(SI_5_), .ZN(n5235) );
  MUX2_X1 U6676 ( .A(n6737), .B(n6736), .S(n6724), .Z(n5269) );
  OR2_X1 U6677 ( .A1(n5273), .A2(n6738), .ZN(n5243) );
  OR2_X1 U6678 ( .A1(n9173), .A2(n6736), .ZN(n5242) );
  NAND2_X1 U6679 ( .A1(n5239), .A2(n5238), .ZN(n5265) );
  NAND2_X1 U6680 ( .A1(n5265), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5240) );
  XNOR2_X1 U6681 ( .A(n5237), .B(n5240), .ZN(n6806) );
  OR2_X1 U6682 ( .A1(n6777), .A2(n6806), .ZN(n5241) );
  OR2_X1 U6683 ( .A1(n10222), .A2(n5793), .ZN(n5244) );
  NAND2_X1 U6684 ( .A1(n5245), .A2(n5244), .ZN(n5246) );
  XNOR2_X1 U6685 ( .A(n5246), .B(n7361), .ZN(n7432) );
  NAND2_X1 U6686 ( .A1(n9474), .A2(n5145), .ZN(n5248) );
  INV_X1 U6687 ( .A(n5795), .ZN(n5302) );
  OR2_X1 U6688 ( .A1(n10222), .A2(n5302), .ZN(n5247) );
  AND2_X1 U6689 ( .A1(n5248), .A2(n5247), .ZN(n5250) );
  AOI22_X1 U6690 ( .A1(n7330), .A2(n7332), .B1(n7432), .B2(n5250), .ZN(n5249)
         );
  NAND2_X1 U6691 ( .A1(n7329), .A2(n5249), .ZN(n5256) );
  OAI21_X1 U6692 ( .B1(n7330), .B2(n7332), .A(n5250), .ZN(n5254) );
  INV_X1 U6693 ( .A(n7432), .ZN(n5253) );
  INV_X1 U6694 ( .A(n7332), .ZN(n5251) );
  INV_X1 U6695 ( .A(n5250), .ZN(n7431) );
  AND2_X1 U6696 ( .A1(n5251), .A2(n7431), .ZN(n5252) );
  INV_X1 U6697 ( .A(n7330), .ZN(n7430) );
  AOI22_X1 U6698 ( .A1(n5254), .A2(n5253), .B1(n5252), .B2(n7430), .ZN(n5255)
         );
  NAND2_X1 U6699 ( .A1(n5256), .A2(n5255), .ZN(n7247) );
  NAND2_X1 U6700 ( .A1(n5755), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5264) );
  INV_X1 U6701 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5257) );
  OR2_X1 U6702 ( .A1(n4593), .A2(n5257), .ZN(n5263) );
  AND2_X1 U6703 ( .A1(n5259), .A2(n5258), .ZN(n5260) );
  OR2_X1 U6704 ( .A1(n5260), .A2(n5303), .ZN(n7412) );
  OR2_X1 U6705 ( .A1(n5856), .A2(n7412), .ZN(n5262) );
  INV_X1 U6706 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7413) );
  OR2_X1 U6707 ( .A1(n5806), .A2(n7413), .ZN(n5261) );
  NAND4_X1 U6708 ( .A1(n5264), .A2(n5263), .A3(n5262), .A4(n5261), .ZN(n9473)
         );
  NAND2_X1 U6709 ( .A1(n9473), .A2(n5795), .ZN(n5277) );
  OAI21_X1 U6710 ( .B1(n5265), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5266) );
  XNOR2_X1 U6711 ( .A(n5266), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6881) );
  AOI22_X1 U6712 ( .A1(n5579), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6713), .B2(
        n6881), .ZN(n5275) );
  NAND2_X1 U6713 ( .A1(n5268), .A2(n5267), .ZN(n5272) );
  INV_X1 U6714 ( .A(n5269), .ZN(n5270) );
  NAND2_X1 U6715 ( .A1(n5270), .A2(SI_6_), .ZN(n5271) );
  MUX2_X1 U6716 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6724), .Z(n5289) );
  XNOR2_X1 U6717 ( .A(n5288), .B(n5286), .ZN(n6743) );
  NAND2_X1 U6718 ( .A1(n6743), .A2(n5368), .ZN(n5274) );
  OR2_X1 U6719 ( .A1(n7526), .A2(n5793), .ZN(n5276) );
  NAND2_X1 U6720 ( .A1(n5277), .A2(n5276), .ZN(n5278) );
  XNOR2_X1 U6721 ( .A(n5278), .B(n7361), .ZN(n5281) );
  NAND2_X1 U6722 ( .A1(n9473), .A2(n5145), .ZN(n5280) );
  OR2_X1 U6723 ( .A1(n7526), .A2(n5302), .ZN(n5279) );
  AND2_X1 U6724 ( .A1(n5280), .A2(n5279), .ZN(n5282) );
  NAND2_X1 U6725 ( .A1(n5281), .A2(n5282), .ZN(n7248) );
  INV_X1 U6726 ( .A(n5281), .ZN(n5284) );
  INV_X1 U6727 ( .A(n5282), .ZN(n5283) );
  NAND2_X1 U6728 ( .A1(n5284), .A2(n5283), .ZN(n7249) );
  NAND2_X1 U6729 ( .A1(n5289), .A2(SI_7_), .ZN(n5290) );
  MUX2_X1 U6730 ( .A(n6748), .B(n6750), .S(n6724), .Z(n5292) );
  INV_X1 U6731 ( .A(SI_8_), .ZN(n5291) );
  INV_X1 U6732 ( .A(n5292), .ZN(n5293) );
  NAND2_X1 U6733 ( .A1(n5293), .A2(SI_8_), .ZN(n5294) );
  XNOR2_X1 U6734 ( .A(n5315), .B(n5316), .ZN(n6747) );
  NAND2_X1 U6735 ( .A1(n6747), .A2(n5368), .ZN(n5301) );
  OR2_X1 U6736 ( .A1(n5295), .A2(n5051), .ZN(n5297) );
  MUX2_X1 U6737 ( .A(n5297), .B(P1_IR_REG_31__SCAN_IN), .S(n5296), .Z(n5299)
         );
  NAND2_X1 U6738 ( .A1(n5299), .A2(n5298), .ZN(n10084) );
  INV_X1 U6739 ( .A(n10084), .ZN(n6883) );
  AOI22_X1 U6740 ( .A1(n5579), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6713), .B2(
        n6883), .ZN(n5300) );
  OR2_X1 U6741 ( .A1(n10229), .A2(n5302), .ZN(n5310) );
  NAND2_X1 U6742 ( .A1(n5755), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5308) );
  INV_X1 U6743 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6873) );
  OR2_X1 U6744 ( .A1(n4593), .A2(n6873), .ZN(n5307) );
  NAND2_X1 U6745 ( .A1(n5303), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5327) );
  OR2_X1 U6746 ( .A1(n5303), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6747 ( .A1(n5327), .A2(n5304), .ZN(n7625) );
  OR2_X1 U6748 ( .A1(n5856), .A2(n7625), .ZN(n5306) );
  INV_X1 U6749 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7626) );
  OR2_X1 U6750 ( .A1(n5806), .A2(n7626), .ZN(n5305) );
  NAND4_X1 U6751 ( .A1(n5308), .A2(n5307), .A3(n5306), .A4(n5305), .ZN(n9472)
         );
  NAND2_X1 U6752 ( .A1(n9472), .A2(n5145), .ZN(n5309) );
  NAND2_X1 U6753 ( .A1(n5310), .A2(n5309), .ZN(n5313) );
  NAND2_X1 U6754 ( .A1(n9472), .A2(n5795), .ZN(n5311) );
  OAI21_X1 U6755 ( .B1(n10229), .B2(n5793), .A(n5311), .ZN(n5312) );
  XNOR2_X1 U6756 ( .A(n5312), .B(n7361), .ZN(n7421) );
  INV_X1 U6757 ( .A(n5313), .ZN(n5314) );
  MUX2_X1 U6758 ( .A(n6760), .B(n8352), .S(n6724), .Z(n5320) );
  INV_X1 U6759 ( .A(SI_9_), .ZN(n5319) );
  INV_X1 U6760 ( .A(n5320), .ZN(n5321) );
  NAND2_X1 U6761 ( .A1(n5321), .A2(SI_9_), .ZN(n5322) );
  XNOR2_X1 U6762 ( .A(n5341), .B(n5028), .ZN(n6758) );
  NAND2_X1 U6763 ( .A1(n6758), .A2(n5368), .ZN(n5325) );
  NAND2_X1 U6764 ( .A1(n5298), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5323) );
  XNOR2_X1 U6765 ( .A(n5323), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10102) );
  AOI22_X1 U6766 ( .A1(n5579), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6713), .B2(
        n10102), .ZN(n5324) );
  NAND2_X1 U6767 ( .A1(n10236), .A2(n5817), .ZN(n5334) );
  NAND2_X1 U6768 ( .A1(n5755), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5332) );
  INV_X1 U6769 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6770 ( .A1(n5327), .A2(n5326), .ZN(n5328) );
  NAND2_X1 U6771 ( .A1(n5352), .A2(n5328), .ZN(n7785) );
  OR2_X1 U6772 ( .A1(n5856), .A2(n7785), .ZN(n5331) );
  INV_X1 U6773 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7786) );
  OR2_X1 U6774 ( .A1(n5806), .A2(n7786), .ZN(n5330) );
  INV_X1 U6775 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6874) );
  OR2_X1 U6776 ( .A1(n4593), .A2(n6874), .ZN(n5329) );
  NAND4_X1 U6777 ( .A1(n5332), .A2(n5331), .A3(n5330), .A4(n5329), .ZN(n9937)
         );
  NAND2_X1 U6778 ( .A1(n9937), .A2(n5795), .ZN(n5333) );
  NAND2_X1 U6779 ( .A1(n5334), .A2(n5333), .ZN(n5335) );
  XNOR2_X1 U6780 ( .A(n5335), .B(n5814), .ZN(n5337) );
  AND2_X1 U6781 ( .A1(n9937), .A2(n5145), .ZN(n5336) );
  AOI21_X1 U6782 ( .B1(n10236), .B2(n5795), .A(n5336), .ZN(n5338) );
  XNOR2_X1 U6783 ( .A(n5337), .B(n5338), .ZN(n7697) );
  INV_X1 U6784 ( .A(n5337), .ZN(n5339) );
  NAND2_X1 U6785 ( .A1(n5339), .A2(n5338), .ZN(n5340) );
  INV_X1 U6786 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6789) );
  MUX2_X1 U6787 ( .A(n6789), .B(n8170), .S(n6724), .Z(n5345) );
  INV_X1 U6788 ( .A(SI_10_), .ZN(n5344) );
  INV_X1 U6789 ( .A(n5345), .ZN(n5346) );
  NAND2_X1 U6790 ( .A1(n5346), .A2(SI_10_), .ZN(n5347) );
  XNOR2_X1 U6791 ( .A(n5366), .B(n5030), .ZN(n6762) );
  NAND2_X1 U6792 ( .A1(n6762), .A2(n5368), .ZN(n5350) );
  NAND2_X1 U6793 ( .A1(n5348), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5370) );
  XNOR2_X1 U6794 ( .A(n5370), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6945) );
  AOI22_X1 U6795 ( .A1(n5579), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6713), .B2(
        n6945), .ZN(n5349) );
  NAND2_X1 U6796 ( .A1(n9948), .A2(n5817), .ZN(n5359) );
  NAND2_X1 U6797 ( .A1(n5755), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5357) );
  INV_X1 U6798 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5351) );
  OR2_X1 U6799 ( .A1(n5806), .A2(n5351), .ZN(n5356) );
  INV_X1 U6800 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6887) );
  NAND2_X1 U6801 ( .A1(n5352), .A2(n6887), .ZN(n5353) );
  NAND2_X1 U6802 ( .A1(n5377), .A2(n5353), .ZN(n9944) );
  OR2_X1 U6803 ( .A1(n5856), .A2(n9944), .ZN(n5355) );
  INV_X1 U6804 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6876) );
  OR2_X1 U6805 ( .A1(n4593), .A2(n6876), .ZN(n5354) );
  OR2_X1 U6806 ( .A1(n7816), .A2(n5302), .ZN(n5358) );
  NAND2_X1 U6807 ( .A1(n5359), .A2(n5358), .ZN(n5360) );
  XNOR2_X1 U6808 ( .A(n5360), .B(n7361), .ZN(n7534) );
  NOR2_X1 U6809 ( .A1(n7816), .A2(n5811), .ZN(n5361) );
  AOI21_X1 U6810 ( .B1(n9948), .B2(n5795), .A(n5361), .ZN(n7533) );
  AND2_X1 U6811 ( .A1(n7534), .A2(n7533), .ZN(n5365) );
  INV_X1 U6812 ( .A(n7534), .ZN(n5363) );
  INV_X1 U6813 ( .A(n7533), .ZN(n5362) );
  NAND2_X1 U6814 ( .A1(n5363), .A2(n5362), .ZN(n5364) );
  INV_X1 U6815 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6770) );
  MUX2_X1 U6816 ( .A(n8312), .B(n6770), .S(n6724), .Z(n5392) );
  NAND2_X1 U6817 ( .A1(n6769), .A2(n5368), .ZN(n5374) );
  NAND2_X1 U6818 ( .A1(n5370), .A2(n5369), .ZN(n5371) );
  NAND2_X1 U6819 ( .A1(n5371), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5372) );
  XNOR2_X1 U6820 ( .A(n5372), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7506) );
  AOI22_X1 U6821 ( .A1(n5579), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6713), .B2(
        n7506), .ZN(n5373) );
  NAND2_X1 U6822 ( .A1(n7895), .A2(n5817), .ZN(n5384) );
  NAND2_X1 U6823 ( .A1(n8101), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5382) );
  INV_X1 U6824 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5375) );
  OR2_X1 U6825 ( .A1(n5175), .A2(n5375), .ZN(n5381) );
  INV_X1 U6826 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7823) );
  OR2_X1 U6827 ( .A1(n5806), .A2(n7823), .ZN(n5380) );
  INV_X1 U6828 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5376) );
  AND2_X1 U6829 ( .A1(n5377), .A2(n5376), .ZN(n5378) );
  OR2_X1 U6830 ( .A1(n5378), .A2(n5406), .ZN(n7822) );
  OR2_X1 U6831 ( .A1(n5856), .A2(n7822), .ZN(n5379) );
  NAND4_X1 U6832 ( .A1(n5382), .A2(n5381), .A3(n5380), .A4(n5379), .ZN(n9936)
         );
  NAND2_X1 U6833 ( .A1(n9936), .A2(n5795), .ZN(n5383) );
  NAND2_X1 U6834 ( .A1(n5384), .A2(n5383), .ZN(n5385) );
  XNOR2_X1 U6835 ( .A(n5385), .B(n5814), .ZN(n5389) );
  AND2_X1 U6836 ( .A1(n9936), .A2(n5145), .ZN(n5386) );
  AOI21_X1 U6837 ( .B1(n7895), .B2(n5795), .A(n5386), .ZN(n5387) );
  XNOR2_X1 U6838 ( .A(n5389), .B(n5387), .ZN(n7648) );
  INV_X1 U6839 ( .A(n5387), .ZN(n5388) );
  NAND2_X1 U6840 ( .A1(n5389), .A2(n5388), .ZN(n5390) );
  INV_X1 U6841 ( .A(n5392), .ZN(n5393) );
  INV_X1 U6842 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6825) );
  INV_X1 U6843 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6827) );
  MUX2_X1 U6844 ( .A(n6825), .B(n6827), .S(n6724), .Z(n5397) );
  INV_X1 U6845 ( .A(SI_12_), .ZN(n5396) );
  INV_X1 U6846 ( .A(n5397), .ZN(n5398) );
  NAND2_X1 U6847 ( .A1(n5398), .A2(SI_12_), .ZN(n5399) );
  XNOR2_X1 U6848 ( .A(n5423), .B(n5422), .ZN(n6824) );
  NAND2_X1 U6849 ( .A1(n6824), .A2(n5368), .ZN(n5405) );
  OR2_X1 U6850 ( .A1(n5400), .A2(n5051), .ZN(n5402) );
  MUX2_X1 U6851 ( .A(n5402), .B(P1_IR_REG_31__SCAN_IN), .S(n5401), .Z(n5403)
         );
  AND2_X1 U6852 ( .A1(n5403), .A2(n5427), .ZN(n10114) );
  AOI22_X1 U6853 ( .A1(n5579), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6713), .B2(
        n10114), .ZN(n5404) );
  NAND2_X1 U6854 ( .A1(n9996), .A2(n5817), .ZN(n5413) );
  NAND2_X1 U6855 ( .A1(n5755), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5411) );
  INV_X1 U6856 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7908) );
  OR2_X1 U6857 ( .A1(n5806), .A2(n7908), .ZN(n5410) );
  NAND2_X1 U6858 ( .A1(n5406), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5432) );
  OR2_X1 U6859 ( .A1(n5406), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U6860 ( .A1(n5432), .A2(n5407), .ZN(n7907) );
  OR2_X1 U6861 ( .A1(n5856), .A2(n7907), .ZN(n5409) );
  INV_X1 U6862 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7510) );
  OR2_X1 U6863 ( .A1(n4593), .A2(n7510), .ZN(n5408) );
  OR2_X1 U6864 ( .A1(n7899), .A2(n5302), .ZN(n5412) );
  NAND2_X1 U6865 ( .A1(n5413), .A2(n5412), .ZN(n5414) );
  XNOR2_X1 U6866 ( .A(n5414), .B(n7361), .ZN(n5417) );
  NOR2_X1 U6867 ( .A1(n7899), .A2(n5811), .ZN(n5415) );
  AOI21_X1 U6868 ( .B1(n9996), .B2(n5795), .A(n5415), .ZN(n5416) );
  NAND2_X1 U6869 ( .A1(n5417), .A2(n5416), .ZN(n5420) );
  OR2_X1 U6870 ( .A1(n5417), .A2(n5416), .ZN(n5418) );
  NAND2_X1 U6871 ( .A1(n5420), .A2(n5418), .ZN(n7796) );
  INV_X1 U6872 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6936) );
  MUX2_X1 U6873 ( .A(n6936), .B(n8288), .S(n6724), .Z(n5424) );
  INV_X1 U6874 ( .A(SI_13_), .ZN(n8331) );
  INV_X1 U6875 ( .A(n5424), .ZN(n5425) );
  NAND2_X1 U6876 ( .A1(n5425), .A2(SI_13_), .ZN(n5426) );
  XNOR2_X1 U6877 ( .A(n5446), .B(n5031), .ZN(n6892) );
  NAND2_X1 U6878 ( .A1(n6892), .A2(n5368), .ZN(n5430) );
  NAND2_X1 U6879 ( .A1(n5427), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5428) );
  XNOR2_X1 U6880 ( .A(n5428), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10127) );
  AOI22_X1 U6881 ( .A1(n5579), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6713), .B2(
        n10127), .ZN(n5429) );
  NAND2_X1 U6882 ( .A1(n9869), .A2(n5817), .ZN(n5439) );
  NAND2_X1 U6883 ( .A1(n5755), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5437) );
  INV_X1 U6884 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7513) );
  OR2_X1 U6885 ( .A1(n4593), .A2(n7513), .ZN(n5436) );
  INV_X1 U6886 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6887 ( .A1(n5432), .A2(n5431), .ZN(n5433) );
  NAND2_X1 U6888 ( .A1(n5455), .A2(n5433), .ZN(n7946) );
  OR2_X1 U6889 ( .A1(n5856), .A2(n7946), .ZN(n5435) );
  INV_X1 U6890 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7947) );
  OR2_X1 U6891 ( .A1(n5806), .A2(n7947), .ZN(n5434) );
  NAND4_X1 U6892 ( .A1(n5437), .A2(n5436), .A3(n5435), .A4(n5434), .ZN(n9471)
         );
  NAND2_X1 U6893 ( .A1(n9471), .A2(n5816), .ZN(n5438) );
  NAND2_X1 U6894 ( .A1(n5439), .A2(n5438), .ZN(n5440) );
  XNOR2_X1 U6895 ( .A(n5440), .B(n7361), .ZN(n5442) );
  AND2_X1 U6896 ( .A1(n9471), .A2(n5145), .ZN(n5441) );
  AOI21_X1 U6897 ( .B1(n9869), .B2(n5816), .A(n5441), .ZN(n5443) );
  AND2_X1 U6898 ( .A1(n5442), .A2(n5443), .ZN(n7828) );
  INV_X1 U6899 ( .A(n5442), .ZN(n5445) );
  INV_X1 U6900 ( .A(n5443), .ZN(n5444) );
  NAND2_X1 U6901 ( .A1(n5445), .A2(n5444), .ZN(n7829) );
  INV_X1 U6902 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6954) );
  INV_X1 U6903 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6953) );
  MUX2_X1 U6904 ( .A(n6954), .B(n6953), .S(n6724), .Z(n5466) );
  XNOR2_X1 U6905 ( .A(n5470), .B(n5465), .ZN(n6952) );
  NAND2_X1 U6906 ( .A1(n6952), .A2(n5368), .ZN(n5452) );
  INV_X1 U6907 ( .A(n5449), .ZN(n5450) );
  NAND2_X1 U6908 ( .A1(n5450), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5476) );
  XNOR2_X1 U6909 ( .A(n5476), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7518) );
  AOI22_X1 U6910 ( .A1(n5579), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6713), .B2(
        n7518), .ZN(n5451) );
  NAND2_X1 U6911 ( .A1(n9864), .A2(n5817), .ZN(n5462) );
  NAND2_X1 U6912 ( .A1(n5755), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5460) );
  INV_X1 U6913 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n5453) );
  OR2_X1 U6914 ( .A1(n5806), .A2(n5453), .ZN(n5459) );
  INV_X1 U6915 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5454) );
  AND2_X1 U6916 ( .A1(n5455), .A2(n5454), .ZN(n5456) );
  OR2_X1 U6917 ( .A1(n5456), .A2(n5482), .ZN(n9062) );
  OR2_X1 U6918 ( .A1(n5856), .A2(n9062), .ZN(n5458) );
  INV_X1 U6919 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9496) );
  OR2_X1 U6920 ( .A1(n4593), .A2(n9496), .ZN(n5457) );
  NAND4_X1 U6921 ( .A1(n5460), .A2(n5459), .A3(n5458), .A4(n5457), .ZN(n9767)
         );
  NAND2_X1 U6922 ( .A1(n9767), .A2(n5816), .ZN(n5461) );
  NAND2_X1 U6923 ( .A1(n5462), .A2(n5461), .ZN(n5463) );
  XNOR2_X1 U6924 ( .A(n5463), .B(n7361), .ZN(n5490) );
  INV_X1 U6925 ( .A(n5490), .ZN(n5464) );
  NAND2_X2 U6926 ( .A1(n5489), .A2(n5464), .ZN(n9055) );
  INV_X1 U6927 ( .A(n5466), .ZN(n5467) );
  NAND2_X1 U6928 ( .A1(n5467), .A2(SI_14_), .ZN(n5468) );
  INV_X1 U6929 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7017) );
  INV_X1 U6930 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7019) );
  MUX2_X1 U6931 ( .A(n7017), .B(n7019), .S(n6724), .Z(n5472) );
  INV_X1 U6932 ( .A(SI_15_), .ZN(n5471) );
  INV_X1 U6933 ( .A(n5472), .ZN(n5473) );
  NAND2_X1 U6934 ( .A1(n5473), .A2(SI_15_), .ZN(n5474) );
  XNOR2_X1 U6935 ( .A(n5499), .B(n5498), .ZN(n7016) );
  NAND2_X1 U6936 ( .A1(n7016), .A2(n5368), .ZN(n5480) );
  NAND2_X1 U6937 ( .A1(n5476), .A2(n5475), .ZN(n5477) );
  NAND2_X1 U6938 ( .A1(n5477), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5478) );
  XNOR2_X1 U6939 ( .A(n5478), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10141) );
  AOI22_X1 U6940 ( .A1(n5579), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6713), .B2(
        n10141), .ZN(n5479) );
  NAND2_X1 U6941 ( .A1(n5755), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5487) );
  INV_X1 U6942 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5481) );
  OR2_X1 U6943 ( .A1(n5738), .A2(n5481), .ZN(n5486) );
  NOR2_X1 U6944 ( .A1(n5482), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5483) );
  OR2_X1 U6945 ( .A1(n5509), .A2(n5483), .ZN(n9777) );
  OR2_X1 U6946 ( .A1(n5856), .A2(n9777), .ZN(n5485) );
  INV_X1 U6947 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9778) );
  OR2_X1 U6948 ( .A1(n5806), .A2(n9778), .ZN(n5484) );
  OAI22_X1 U6949 ( .A1(n9759), .A2(n5793), .B1(n9750), .B2(n5302), .ZN(n5488)
         );
  XNOR2_X1 U6950 ( .A(n5488), .B(n7361), .ZN(n5494) );
  NAND2_X1 U6951 ( .A1(n9864), .A2(n5795), .ZN(n5492) );
  NAND2_X1 U6952 ( .A1(n9767), .A2(n5145), .ZN(n5491) );
  NAND2_X1 U6953 ( .A1(n5492), .A2(n5491), .ZN(n9054) );
  NAND2_X1 U6954 ( .A1(n5493), .A2(n9059), .ZN(n9156) );
  OAI22_X1 U6955 ( .A1(n9759), .A2(n5302), .B1(n9750), .B2(n5811), .ZN(n9155)
         );
  NAND2_X1 U6956 ( .A1(n9156), .A2(n9155), .ZN(n9153) );
  NAND2_X1 U6957 ( .A1(n9059), .A2(n9055), .ZN(n5496) );
  INV_X1 U6958 ( .A(n5494), .ZN(n5495) );
  INV_X1 U6959 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7032) );
  INV_X1 U6960 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5500) );
  MUX2_X1 U6961 ( .A(n7032), .B(n5500), .S(n6724), .Z(n5502) );
  INV_X1 U6962 ( .A(SI_16_), .ZN(n5501) );
  NAND2_X1 U6963 ( .A1(n5502), .A2(n5501), .ZN(n5524) );
  INV_X1 U6964 ( .A(n5502), .ZN(n5503) );
  NAND2_X1 U6965 ( .A1(n5503), .A2(SI_16_), .ZN(n5504) );
  XNOR2_X1 U6966 ( .A(n5523), .B(n5522), .ZN(n7006) );
  NAND2_X1 U6967 ( .A1(n7006), .A2(n5368), .ZN(n5508) );
  NAND2_X1 U6968 ( .A1(n5505), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5506) );
  XNOR2_X1 U6969 ( .A(n5506), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10153) );
  AOI22_X1 U6970 ( .A1(n5579), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6713), .B2(
        n10153), .ZN(n5507) );
  NAND2_X1 U6971 ( .A1(n9853), .A2(n5817), .ZN(n5516) );
  NAND2_X1 U6972 ( .A1(n5755), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5514) );
  INV_X1 U6973 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9745) );
  OR2_X1 U6974 ( .A1(n5806), .A2(n9745), .ZN(n5513) );
  OR2_X1 U6975 ( .A1(n5509), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U6976 ( .A1(n5528), .A2(n5510), .ZN(n9744) );
  OR2_X1 U6977 ( .A1(n5856), .A2(n9744), .ZN(n5512) );
  INV_X1 U6978 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9499) );
  OR2_X1 U6979 ( .A1(n4593), .A2(n9499), .ZN(n5511) );
  OR2_X1 U6980 ( .A1(n9770), .A2(n5302), .ZN(n5515) );
  NAND2_X1 U6981 ( .A1(n5516), .A2(n5515), .ZN(n5517) );
  NAND2_X1 U6982 ( .A1(n9853), .A2(n5795), .ZN(n5519) );
  OR2_X1 U6983 ( .A1(n9770), .A2(n5811), .ZN(n5518) );
  NAND2_X1 U6984 ( .A1(n5519), .A2(n5518), .ZN(n9095) );
  OAI21_X1 U6985 ( .B1(n9093), .B2(n9094), .A(n9095), .ZN(n5521) );
  NAND2_X1 U6986 ( .A1(n9093), .A2(n9094), .ZN(n5520) );
  NAND2_X1 U6987 ( .A1(n5521), .A2(n5520), .ZN(n9102) );
  INV_X1 U6988 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7139) );
  INV_X1 U6989 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7109) );
  MUX2_X1 U6990 ( .A(n7139), .B(n7109), .S(n6724), .Z(n5543) );
  XNOR2_X1 U6991 ( .A(n5543), .B(SI_17_), .ZN(n5542) );
  XNOR2_X1 U6992 ( .A(n5547), .B(n5542), .ZN(n7108) );
  NAND2_X1 U6993 ( .A1(n7108), .A2(n5368), .ZN(n5527) );
  XNOR2_X1 U6994 ( .A(n5549), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U6995 ( .A1(n5579), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6713), .B2(
        n10167), .ZN(n5526) );
  NAND2_X1 U6996 ( .A1(n9846), .A2(n5817), .ZN(n5536) );
  NAND2_X1 U6997 ( .A1(n5755), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5534) );
  INV_X1 U6998 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9501) );
  OR2_X1 U6999 ( .A1(n5738), .A2(n9501), .ZN(n5533) );
  INV_X1 U7000 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8398) );
  NAND2_X1 U7001 ( .A1(n5528), .A2(n8398), .ZN(n5529) );
  NAND2_X1 U7002 ( .A1(n5555), .A2(n5529), .ZN(n9724) );
  OR2_X1 U7003 ( .A1(n5856), .A2(n9724), .ZN(n5532) );
  INV_X1 U7004 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5530) );
  OR2_X1 U7005 ( .A1(n5806), .A2(n5530), .ZN(n5531) );
  NAND4_X1 U7006 ( .A1(n5534), .A2(n5533), .A3(n5532), .A4(n5531), .ZN(n9715)
         );
  NAND2_X1 U7007 ( .A1(n9715), .A2(n5795), .ZN(n5535) );
  NAND2_X1 U7008 ( .A1(n5536), .A2(n5535), .ZN(n5537) );
  XNOR2_X1 U7009 ( .A(n5537), .B(n7361), .ZN(n5540) );
  AND2_X1 U7010 ( .A1(n9715), .A2(n5145), .ZN(n5538) );
  AOI21_X1 U7011 ( .B1(n9846), .B2(n5795), .A(n5538), .ZN(n5539) );
  XNOR2_X1 U7012 ( .A(n5540), .B(n5539), .ZN(n9105) );
  NAND2_X1 U7013 ( .A1(n5540), .A2(n5539), .ZN(n5541) );
  INV_X1 U7014 ( .A(n5543), .ZN(n5544) );
  NAND2_X1 U7015 ( .A1(n5544), .A2(SI_17_), .ZN(n5545) );
  MUX2_X1 U7016 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6724), .Z(n5572) );
  XNOR2_X1 U7017 ( .A(n5572), .B(SI_18_), .ZN(n5569) );
  XNOR2_X1 U7018 ( .A(n5571), .B(n5569), .ZN(n7270) );
  NAND2_X1 U7019 ( .A1(n7270), .A2(n5368), .ZN(n5553) );
  INV_X1 U7020 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U7021 ( .A1(n5549), .A2(n5548), .ZN(n5550) );
  NAND2_X1 U7022 ( .A1(n5550), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5551) );
  XNOR2_X1 U7023 ( .A(n5551), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9523) );
  AOI22_X1 U7024 ( .A1(n5579), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6713), .B2(
        n9523), .ZN(n5552) );
  NAND2_X1 U7025 ( .A1(n9841), .A2(n5817), .ZN(n5563) );
  INV_X1 U7026 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5554) );
  AND2_X1 U7027 ( .A1(n5555), .A2(n5554), .ZN(n5556) );
  OR2_X1 U7028 ( .A1(n5556), .A2(n5582), .ZN(n9717) );
  INV_X1 U7029 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9709) );
  OR2_X1 U7030 ( .A1(n5806), .A2(n9709), .ZN(n5557) );
  OAI21_X1 U7031 ( .B1(n9717), .B2(n5856), .A(n5557), .ZN(n5561) );
  NAND2_X1 U7032 ( .A1(n5755), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5559) );
  INV_X1 U7033 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9526) );
  OR2_X1 U7034 ( .A1(n5738), .A2(n9526), .ZN(n5558) );
  NAND2_X1 U7035 ( .A1(n5559), .A2(n5558), .ZN(n5560) );
  NOR2_X1 U7036 ( .A1(n5561), .A2(n5560), .ZN(n9106) );
  OR2_X1 U7037 ( .A1(n9106), .A2(n5302), .ZN(n5562) );
  NAND2_X1 U7038 ( .A1(n5563), .A2(n5562), .ZN(n5564) );
  XNOR2_X1 U7039 ( .A(n5564), .B(n7361), .ZN(n5567) );
  NAND2_X1 U7040 ( .A1(n9841), .A2(n5795), .ZN(n5566) );
  OR2_X1 U7041 ( .A1(n9106), .A2(n5811), .ZN(n5565) );
  NAND2_X1 U7042 ( .A1(n5566), .A2(n5565), .ZN(n8047) );
  INV_X1 U7043 ( .A(n5567), .ZN(n5568) );
  INV_X1 U7044 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U7045 ( .A1(n5572), .A2(SI_18_), .ZN(n5573) );
  INV_X1 U7046 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7353) );
  INV_X1 U7047 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7355) );
  MUX2_X1 U7048 ( .A(n7353), .B(n7355), .S(n6724), .Z(n5575) );
  INV_X1 U7049 ( .A(SI_19_), .ZN(n5574) );
  NAND2_X1 U7050 ( .A1(n5575), .A2(n5574), .ZN(n5600) );
  INV_X1 U7051 ( .A(n5575), .ZN(n5576) );
  NAND2_X1 U7052 ( .A1(n5576), .A2(SI_19_), .ZN(n5577) );
  NAND2_X1 U7053 ( .A1(n5600), .A2(n5577), .ZN(n5597) );
  XNOR2_X1 U7054 ( .A(n5596), .B(n5597), .ZN(n7352) );
  NAND2_X1 U7055 ( .A1(n7352), .A2(n5368), .ZN(n5581) );
  AOI22_X1 U7056 ( .A1(n5579), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6713), .B2(
        n10180), .ZN(n5580) );
  NAND2_X1 U7057 ( .A1(n9836), .A2(n5817), .ZN(n5588) );
  NOR2_X1 U7058 ( .A1(n5582), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5583) );
  OR2_X1 U7059 ( .A1(n5608), .A2(n5583), .ZN(n9695) );
  AOI22_X1 U7060 ( .A1(n8101), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n5755), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5586) );
  INV_X1 U7061 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n5584) );
  OR2_X1 U7062 ( .A1(n5806), .A2(n5584), .ZN(n5585) );
  OAI211_X1 U7063 ( .C1(n9695), .C2(n5856), .A(n5586), .B(n5585), .ZN(n9714)
         );
  NAND2_X1 U7064 ( .A1(n9714), .A2(n5795), .ZN(n5587) );
  NAND2_X1 U7065 ( .A1(n5588), .A2(n5587), .ZN(n5589) );
  XNOR2_X1 U7066 ( .A(n5589), .B(n5814), .ZN(n5592) );
  NAND2_X1 U7067 ( .A1(n9836), .A2(n5795), .ZN(n5591) );
  NAND2_X1 U7068 ( .A1(n9714), .A2(n5145), .ZN(n5590) );
  NAND2_X1 U7069 ( .A1(n5591), .A2(n5590), .ZN(n5593) );
  INV_X1 U7070 ( .A(n5592), .ZN(n5595) );
  INV_X1 U7071 ( .A(n5593), .ZN(n5594) );
  NAND2_X1 U7072 ( .A1(n5595), .A2(n5594), .ZN(n8053) );
  OAI21_X1 U7073 ( .B1(n8057), .B2(n8054), .A(n8053), .ZN(n9122) );
  INV_X1 U7074 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U7075 ( .A1(n5599), .A2(n5598), .ZN(n5601) );
  INV_X1 U7076 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7502) );
  INV_X1 U7077 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7466) );
  MUX2_X1 U7078 ( .A(n7502), .B(n7466), .S(n6724), .Z(n5603) );
  INV_X1 U7079 ( .A(SI_20_), .ZN(n5602) );
  NAND2_X1 U7080 ( .A1(n5603), .A2(n5602), .ZN(n5624) );
  INV_X1 U7081 ( .A(n5603), .ZN(n5604) );
  NAND2_X1 U7082 ( .A1(n5604), .A2(SI_20_), .ZN(n5605) );
  XNOR2_X1 U7083 ( .A(n5623), .B(n5622), .ZN(n7465) );
  NAND2_X1 U7084 ( .A1(n7465), .A2(n5368), .ZN(n5607) );
  OR2_X1 U7085 ( .A1(n9173), .A2(n7466), .ZN(n5606) );
  NAND2_X1 U7086 ( .A1(n9833), .A2(n5817), .ZN(n5613) );
  OR2_X1 U7087 ( .A1(n5608), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U7088 ( .A1(n5627), .A2(n5609), .ZN(n9685) );
  AOI22_X1 U7089 ( .A1(n8101), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n5755), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n5611) );
  INV_X1 U7090 ( .A(n5806), .ZN(n5629) );
  NAND2_X1 U7091 ( .A1(n5629), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5610) );
  OAI211_X1 U7092 ( .C1(n9685), .C2(n5856), .A(n5611), .B(n5610), .ZN(n9701)
         );
  NAND2_X1 U7093 ( .A1(n9701), .A2(n5795), .ZN(n5612) );
  NAND2_X1 U7094 ( .A1(n5613), .A2(n5612), .ZN(n5614) );
  XNOR2_X1 U7095 ( .A(n5614), .B(n5814), .ZN(n5617) );
  NAND2_X1 U7096 ( .A1(n9833), .A2(n5795), .ZN(n5616) );
  NAND2_X1 U7097 ( .A1(n9701), .A2(n5145), .ZN(n5615) );
  NAND2_X1 U7098 ( .A1(n5616), .A2(n5615), .ZN(n5618) );
  NAND2_X1 U7099 ( .A1(n5617), .A2(n5618), .ZN(n9123) );
  NAND2_X1 U7100 ( .A1(n9122), .A2(n9123), .ZN(n5621) );
  INV_X1 U7101 ( .A(n5617), .ZN(n5620) );
  INV_X1 U7102 ( .A(n5618), .ZN(n5619) );
  NAND2_X1 U7103 ( .A1(n5620), .A2(n5619), .ZN(n9124) );
  NAND2_X1 U7104 ( .A1(n5621), .A2(n9124), .ZN(n9076) );
  INV_X1 U7105 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7595) );
  INV_X1 U7106 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8162) );
  MUX2_X1 U7107 ( .A(n7595), .B(n8162), .S(n6724), .Z(n5647) );
  XNOR2_X1 U7108 ( .A(n5647), .B(SI_21_), .ZN(n5646) );
  NAND2_X1 U7109 ( .A1(n7594), .A2(n5368), .ZN(n5626) );
  OR2_X1 U7110 ( .A1(n9173), .A2(n8162), .ZN(n5625) );
  NAND2_X1 U7111 ( .A1(n9827), .A2(n5817), .ZN(n5637) );
  INV_X1 U7112 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9078) );
  NAND2_X1 U7113 ( .A1(n5627), .A2(n9078), .ZN(n5628) );
  INV_X1 U7114 ( .A(n5658), .ZN(n5659) );
  NAND2_X1 U7115 ( .A1(n5628), .A2(n5659), .ZN(n9673) );
  OR2_X1 U7116 ( .A1(n9673), .A2(n5856), .ZN(n5635) );
  INV_X1 U7117 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U7118 ( .A1(n5755), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U7119 ( .A1(n5629), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5630) );
  OAI211_X1 U7120 ( .C1(n4593), .C2(n5632), .A(n5631), .B(n5630), .ZN(n5633)
         );
  INV_X1 U7121 ( .A(n5633), .ZN(n5634) );
  OR2_X1 U7122 ( .A1(n9682), .A2(n5302), .ZN(n5636) );
  NAND2_X1 U7123 ( .A1(n5637), .A2(n5636), .ZN(n5638) );
  XNOR2_X1 U7124 ( .A(n5638), .B(n5814), .ZN(n5640) );
  NOR2_X1 U7125 ( .A1(n9682), .A2(n5811), .ZN(n5639) );
  AOI21_X1 U7126 ( .B1(n9827), .B2(n5816), .A(n5639), .ZN(n5641) );
  XNOR2_X1 U7127 ( .A(n5640), .B(n5641), .ZN(n9077) );
  NAND2_X1 U7128 ( .A1(n9076), .A2(n9077), .ZN(n5644) );
  INV_X1 U7129 ( .A(n5640), .ZN(n5642) );
  NAND2_X1 U7130 ( .A1(n5642), .A2(n5641), .ZN(n5643) );
  INV_X1 U7131 ( .A(n5647), .ZN(n5648) );
  NAND2_X1 U7132 ( .A1(n5648), .A2(SI_21_), .ZN(n5649) );
  INV_X1 U7133 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7659) );
  INV_X1 U7134 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7658) );
  MUX2_X1 U7135 ( .A(n7659), .B(n7658), .S(n6724), .Z(n5652) );
  INV_X1 U7136 ( .A(SI_22_), .ZN(n5651) );
  NAND2_X1 U7137 ( .A1(n5652), .A2(n5651), .ZN(n5673) );
  INV_X1 U7138 ( .A(n5652), .ZN(n5653) );
  NAND2_X1 U7139 ( .A1(n5653), .A2(SI_22_), .ZN(n5654) );
  NAND2_X1 U7140 ( .A1(n5673), .A2(n5654), .ZN(n5674) );
  NAND2_X1 U7141 ( .A1(n7656), .A2(n5368), .ZN(n5656) );
  OR2_X1 U7142 ( .A1(n9173), .A2(n7658), .ZN(n5655) );
  NAND2_X1 U7143 ( .A1(n8101), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5666) );
  INV_X1 U7144 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n5657) );
  OR2_X1 U7145 ( .A1(n5175), .A2(n5657), .ZN(n5665) );
  INV_X1 U7146 ( .A(n5683), .ZN(n5685) );
  INV_X1 U7147 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U7148 ( .A1(n5660), .A2(n5659), .ZN(n5661) );
  NAND2_X1 U7149 ( .A1(n5685), .A2(n5661), .ZN(n9648) );
  OR2_X1 U7150 ( .A1(n5856), .A2(n9648), .ZN(n5664) );
  INV_X1 U7151 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n5662) );
  OR2_X1 U7152 ( .A1(n5806), .A2(n5662), .ZN(n5663) );
  NAND4_X1 U7153 ( .A1(n5666), .A2(n5665), .A3(n5664), .A4(n5663), .ZN(n9666)
         );
  AND2_X1 U7154 ( .A1(n9666), .A2(n5145), .ZN(n5667) );
  AOI21_X1 U7155 ( .B1(n9821), .B2(n5816), .A(n5667), .ZN(n5671) );
  NAND2_X1 U7156 ( .A1(n5672), .A2(n5671), .ZN(n9131) );
  NAND2_X1 U7157 ( .A1(n9821), .A2(n5817), .ZN(n5669) );
  NAND2_X1 U7158 ( .A1(n9666), .A2(n5795), .ZN(n5668) );
  NAND2_X1 U7159 ( .A1(n5669), .A2(n5668), .ZN(n5670) );
  XNOR2_X1 U7160 ( .A(n5670), .B(n5814), .ZN(n9133) );
  INV_X1 U7161 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7749) );
  INV_X1 U7162 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7745) );
  MUX2_X1 U7163 ( .A(n7749), .B(n7745), .S(n6724), .Z(n5677) );
  INV_X1 U7164 ( .A(SI_23_), .ZN(n5676) );
  NAND2_X1 U7165 ( .A1(n5677), .A2(n5676), .ZN(n5699) );
  INV_X1 U7166 ( .A(n5677), .ZN(n5678) );
  NAND2_X1 U7167 ( .A1(n5678), .A2(SI_23_), .ZN(n5679) );
  OR2_X1 U7168 ( .A1(n9173), .A2(n7745), .ZN(n5680) );
  NAND2_X1 U7169 ( .A1(n9816), .A2(n5817), .ZN(n5693) );
  NAND2_X1 U7170 ( .A1(n5755), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5691) );
  INV_X1 U7171 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5682) );
  OR2_X1 U7172 ( .A1(n4593), .A2(n5682), .ZN(n5690) );
  INV_X1 U7173 ( .A(n5703), .ZN(n5704) );
  INV_X1 U7174 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U7175 ( .A1(n5685), .A2(n5684), .ZN(n5686) );
  NAND2_X1 U7176 ( .A1(n5704), .A2(n5686), .ZN(n9632) );
  OR2_X1 U7177 ( .A1(n5856), .A2(n9632), .ZN(n5689) );
  INV_X1 U7178 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5687) );
  OR2_X1 U7179 ( .A1(n5806), .A2(n5687), .ZN(n5688) );
  NAND4_X1 U7180 ( .A1(n5691), .A2(n5690), .A3(n5689), .A4(n5688), .ZN(n9654)
         );
  NAND2_X1 U7181 ( .A1(n9654), .A2(n5795), .ZN(n5692) );
  NAND2_X1 U7182 ( .A1(n5693), .A2(n5692), .ZN(n5694) );
  XNOR2_X1 U7183 ( .A(n5694), .B(n5814), .ZN(n5696) );
  INV_X1 U7184 ( .A(n5696), .ZN(n5695) );
  AOI22_X1 U7185 ( .A1(n9816), .A2(n5795), .B1(n5145), .B2(n9654), .ZN(n9070)
         );
  INV_X1 U7186 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7803) );
  INV_X1 U7187 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7776) );
  MUX2_X1 U7188 ( .A(n7803), .B(n7776), .S(n6724), .Z(n5723) );
  XNOR2_X1 U7189 ( .A(n5723), .B(SI_24_), .ZN(n5722) );
  XNOR2_X1 U7190 ( .A(n5725), .B(n5722), .ZN(n7775) );
  NAND2_X1 U7191 ( .A1(n7775), .A2(n5368), .ZN(n5701) );
  OR2_X1 U7192 ( .A1(n9173), .A2(n7776), .ZN(n5700) );
  NAND2_X1 U7193 ( .A1(n9811), .A2(n5817), .ZN(n5712) );
  NAND2_X1 U7194 ( .A1(n8101), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5710) );
  INV_X1 U7195 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n5702) );
  OR2_X1 U7196 ( .A1(n5175), .A2(n5702), .ZN(n5709) );
  INV_X1 U7197 ( .A(n5732), .ZN(n5734) );
  INV_X1 U7198 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9116) );
  NAND2_X1 U7199 ( .A1(n5704), .A2(n9116), .ZN(n5705) );
  NAND2_X1 U7200 ( .A1(n5734), .A2(n5705), .ZN(n9618) );
  OR2_X1 U7201 ( .A1(n5856), .A2(n9618), .ZN(n5708) );
  INV_X1 U7202 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n5706) );
  OR2_X1 U7203 ( .A1(n5806), .A2(n5706), .ZN(n5707) );
  NAND4_X1 U7204 ( .A1(n5710), .A2(n5709), .A3(n5708), .A4(n5707), .ZN(n9642)
         );
  NAND2_X1 U7205 ( .A1(n9642), .A2(n5795), .ZN(n5711) );
  NAND2_X1 U7206 ( .A1(n5712), .A2(n5711), .ZN(n5713) );
  XNOR2_X1 U7207 ( .A(n5713), .B(n7361), .ZN(n5715) );
  AND2_X1 U7208 ( .A1(n9642), .A2(n5145), .ZN(n5714) );
  AOI21_X1 U7209 ( .B1(n9811), .B2(n5816), .A(n5714), .ZN(n5716) );
  NAND2_X1 U7210 ( .A1(n5715), .A2(n5716), .ZN(n5720) );
  INV_X1 U7211 ( .A(n5715), .ZN(n5718) );
  INV_X1 U7212 ( .A(n5716), .ZN(n5717) );
  NAND2_X1 U7213 ( .A1(n5718), .A2(n5717), .ZN(n5719) );
  NAND2_X1 U7214 ( .A1(n5720), .A2(n5719), .ZN(n9112) );
  INV_X1 U7215 ( .A(n5720), .ZN(n5721) );
  INV_X1 U7216 ( .A(n5723), .ZN(n5724) );
  INV_X1 U7217 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7915) );
  INV_X1 U7218 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7919) );
  MUX2_X1 U7219 ( .A(n7915), .B(n7919), .S(n6724), .Z(n5727) );
  INV_X1 U7220 ( .A(SI_25_), .ZN(n5726) );
  NAND2_X1 U7221 ( .A1(n5727), .A2(n5726), .ZN(n5746) );
  INV_X1 U7222 ( .A(n5727), .ZN(n5728) );
  NAND2_X1 U7223 ( .A1(n5728), .A2(SI_25_), .ZN(n5729) );
  NAND2_X1 U7224 ( .A1(n5746), .A2(n5729), .ZN(n5747) );
  NAND2_X1 U7225 ( .A1(n7914), .A2(n5368), .ZN(n5731) );
  OR2_X1 U7226 ( .A1(n9173), .A2(n7919), .ZN(n5730) );
  NAND2_X1 U7227 ( .A1(n5755), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5742) );
  INV_X1 U7228 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9605) );
  OR2_X1 U7229 ( .A1(n5806), .A2(n9605), .ZN(n5741) );
  INV_X1 U7230 ( .A(n5757), .ZN(n5736) );
  INV_X1 U7231 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U7232 ( .A1(n5734), .A2(n5733), .ZN(n5735) );
  NAND2_X1 U7233 ( .A1(n5736), .A2(n5735), .ZN(n9604) );
  OR2_X1 U7234 ( .A1(n5856), .A2(n9604), .ZN(n5740) );
  INV_X1 U7235 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5737) );
  OR2_X1 U7236 ( .A1(n5738), .A2(n5737), .ZN(n5739) );
  OAI22_X1 U7237 ( .A1(n9603), .A2(n5302), .B1(n9469), .B2(n5811), .ZN(n5767)
         );
  NAND2_X1 U7238 ( .A1(n9808), .A2(n5817), .ZN(n5744) );
  OR2_X1 U7239 ( .A1(n9469), .A2(n5302), .ZN(n5743) );
  NAND2_X1 U7240 ( .A1(n5744), .A2(n5743), .ZN(n5745) );
  XNOR2_X1 U7241 ( .A(n5745), .B(n7361), .ZN(n5766) );
  XOR2_X1 U7242 ( .A(n5767), .B(n5766), .Z(n9086) );
  INV_X1 U7243 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8321) );
  INV_X1 U7244 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7921) );
  MUX2_X1 U7245 ( .A(n8321), .B(n7921), .S(n6724), .Z(n5750) );
  INV_X1 U7246 ( .A(SI_26_), .ZN(n5749) );
  NAND2_X1 U7247 ( .A1(n5750), .A2(n5749), .ZN(n5777) );
  INV_X1 U7248 ( .A(n5750), .ZN(n5751) );
  NAND2_X1 U7249 ( .A1(n5751), .A2(SI_26_), .ZN(n5752) );
  NAND2_X1 U7250 ( .A1(n7920), .A2(n5368), .ZN(n5754) );
  OR2_X1 U7251 ( .A1(n9173), .A2(n7921), .ZN(n5753) );
  NAND2_X1 U7252 ( .A1(n5755), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5762) );
  INV_X1 U7253 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5756) );
  OR2_X1 U7254 ( .A1(n4593), .A2(n5756), .ZN(n5761) );
  OAI21_X1 U7255 ( .B1(n5757), .B2(P1_REG3_REG_26__SCAN_IN), .A(n5785), .ZN(
        n9588) );
  OR2_X1 U7256 ( .A1(n5856), .A2(n9588), .ZN(n5760) );
  INV_X1 U7257 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5758) );
  OR2_X1 U7258 ( .A1(n5806), .A2(n5758), .ZN(n5759) );
  OR2_X1 U7259 ( .A1(n9611), .A2(n5811), .ZN(n5763) );
  NAND2_X1 U7260 ( .A1(n5764), .A2(n5763), .ZN(n5773) );
  OAI22_X1 U7261 ( .A1(n9591), .A2(n5793), .B1(n9611), .B2(n5302), .ZN(n5765)
         );
  XNOR2_X1 U7262 ( .A(n5765), .B(n7361), .ZN(n5772) );
  XOR2_X1 U7263 ( .A(n5773), .B(n5772), .Z(n9142) );
  INV_X1 U7264 ( .A(n9142), .ZN(n5770) );
  INV_X1 U7265 ( .A(n5766), .ZN(n5768) );
  NOR2_X1 U7266 ( .A1(n5768), .A2(n5767), .ZN(n9143) );
  INV_X1 U7267 ( .A(n9143), .ZN(n5769) );
  NAND2_X1 U7268 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  INV_X1 U7269 ( .A(n5772), .ZN(n5774) );
  NAND2_X1 U7270 ( .A1(n5776), .A2(n5775), .ZN(n5778) );
  INV_X1 U7271 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7990) );
  INV_X1 U7272 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7968) );
  MUX2_X1 U7273 ( .A(n7990), .B(n7968), .S(n6724), .Z(n5780) );
  INV_X1 U7274 ( .A(SI_27_), .ZN(n5779) );
  NAND2_X1 U7275 ( .A1(n5780), .A2(n5779), .ZN(n5800) );
  INV_X1 U7276 ( .A(n5780), .ZN(n5781) );
  NAND2_X1 U7277 ( .A1(n5781), .A2(SI_27_), .ZN(n5782) );
  AND2_X1 U7278 ( .A1(n5800), .A2(n5782), .ZN(n5798) );
  NAND2_X1 U7279 ( .A1(n7989), .A2(n5368), .ZN(n5784) );
  OR2_X1 U7280 ( .A1(n9173), .A2(n7968), .ZN(n5783) );
  NAND2_X1 U7281 ( .A1(n5755), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5792) );
  INV_X1 U7282 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8389) );
  OR2_X1 U7283 ( .A1(n4593), .A2(n8389), .ZN(n5791) );
  INV_X1 U7284 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U7285 ( .A1(n5785), .A2(n5877), .ZN(n5787) );
  INV_X1 U7286 ( .A(n5805), .ZN(n5786) );
  NAND2_X1 U7287 ( .A1(n5787), .A2(n5786), .ZN(n9573) );
  OR2_X1 U7288 ( .A1(n5856), .A2(n9573), .ZN(n5790) );
  INV_X1 U7289 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5788) );
  OR2_X1 U7290 ( .A1(n5806), .A2(n5788), .ZN(n5789) );
  OAI22_X1 U7291 ( .A1(n9576), .A2(n5793), .B1(n9557), .B2(n5302), .ZN(n5794)
         );
  XNOR2_X1 U7292 ( .A(n5794), .B(n7361), .ZN(n5797) );
  INV_X1 U7293 ( .A(n9557), .ZN(n9595) );
  AOI22_X1 U7294 ( .A1(n9796), .A2(n5795), .B1(n5145), .B2(n9595), .ZN(n5796)
         );
  NAND2_X1 U7295 ( .A1(n5797), .A2(n5796), .ZN(n5865) );
  OAI21_X1 U7296 ( .B1(n5797), .B2(n5796), .A(n5865), .ZN(n5875) );
  MUX2_X1 U7297 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6724), .Z(n6288) );
  INV_X1 U7298 ( .A(SI_28_), .ZN(n8388) );
  XNOR2_X1 U7299 ( .A(n6288), .B(n8388), .ZN(n6286) );
  NAND2_X1 U7300 ( .A1(n8015), .A2(n5368), .ZN(n5803) );
  INV_X1 U7301 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8017) );
  OR2_X1 U7302 ( .A1(n9173), .A2(n8017), .ZN(n5802) );
  NAND2_X1 U7303 ( .A1(n9791), .A2(n5795), .ZN(n5813) );
  NAND2_X1 U7304 ( .A1(n8101), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5810) );
  INV_X1 U7305 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5804) );
  OR2_X1 U7306 ( .A1(n5175), .A2(n5804), .ZN(n5809) );
  NAND2_X1 U7307 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(n5805), .ZN(n8076) );
  OAI21_X1 U7308 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(n5805), .A(n8076), .ZN(
        n9560) );
  OR2_X1 U7309 ( .A1(n5856), .A2(n9560), .ZN(n5808) );
  INV_X1 U7310 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9561) );
  OR2_X1 U7311 ( .A1(n5806), .A2(n9561), .ZN(n5807) );
  OR2_X1 U7312 ( .A1(n9580), .A2(n5811), .ZN(n5812) );
  NAND2_X1 U7313 ( .A1(n5813), .A2(n5812), .ZN(n5815) );
  XNOR2_X1 U7314 ( .A(n5815), .B(n5814), .ZN(n5819) );
  AOI22_X1 U7315 ( .A1(n9791), .A2(n5817), .B1(n5816), .B2(n8072), .ZN(n5818)
         );
  XNOR2_X1 U7316 ( .A(n5819), .B(n5818), .ZN(n5841) );
  INV_X1 U7317 ( .A(n5841), .ZN(n5866) );
  INV_X1 U7318 ( .A(n9453), .ZN(n9290) );
  AND2_X1 U7319 ( .A1(n9452), .A2(n9290), .ZN(n7164) );
  AND2_X1 U7320 ( .A1(n9462), .A2(n9453), .ZN(n9446) );
  NOR2_X1 U7321 ( .A1(n9994), .A2(n9446), .ZN(n5844) );
  XNOR2_X1 U7322 ( .A(n5820), .B(P1_IR_REG_23__SCAN_IN), .ZN(n7743) );
  INV_X1 U7323 ( .A(n5821), .ZN(n5823) );
  INV_X1 U7324 ( .A(P1_B_REG_SCAN_IN), .ZN(n5822) );
  NAND2_X1 U7325 ( .A1(n5823), .A2(n5822), .ZN(n5826) );
  NAND3_X1 U7326 ( .A1(n5821), .A2(P1_B_REG_SCAN_IN), .A3(n7917), .ZN(n5825)
         );
  INV_X1 U7327 ( .A(n7922), .ZN(n5824) );
  NAND3_X1 U7328 ( .A1(n5826), .A2(n5825), .A3(n5824), .ZN(n6739) );
  NOR4_X1 U7329 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n5835) );
  NOR4_X1 U7330 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5834) );
  INV_X1 U7331 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10200) );
  INV_X1 U7332 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10202) );
  INV_X1 U7333 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10195) );
  INV_X1 U7334 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10199) );
  NAND4_X1 U7335 ( .A1(n10200), .A2(n10202), .A3(n10195), .A4(n10199), .ZN(
        n5832) );
  NOR4_X1 U7336 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5830) );
  NOR4_X1 U7337 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5829) );
  NOR4_X1 U7338 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n5828) );
  NOR4_X1 U7339 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5827) );
  NAND4_X1 U7340 ( .A1(n5830), .A2(n5829), .A3(n5828), .A4(n5827), .ZN(n5831)
         );
  NOR4_X1 U7341 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        n5832), .A4(n5831), .ZN(n5833) );
  AND3_X1 U7342 ( .A1(n5835), .A2(n5834), .A3(n5833), .ZN(n5836) );
  NOR2_X1 U7343 ( .A1(n6739), .A2(n5836), .ZN(n6991) );
  INV_X1 U7344 ( .A(n6991), .ZN(n5840) );
  OR2_X1 U7345 ( .A1(n6739), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U7346 ( .A1(n5821), .A2(n7922), .ZN(n5837) );
  AND2_X1 U7347 ( .A1(n5838), .A2(n5837), .ZN(n7147) );
  OR2_X1 U7348 ( .A1(n6739), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U7349 ( .A1(n7922), .A2(n7917), .ZN(n6751) );
  NAND2_X1 U7350 ( .A1(n5839), .A2(n6751), .ZN(n7146) );
  INV_X1 U7351 ( .A(n7146), .ZN(n7309) );
  INV_X1 U7352 ( .A(n7467), .ZN(n9456) );
  INV_X1 U7353 ( .A(n7149), .ZN(n5842) );
  INV_X1 U7354 ( .A(n6960), .ZN(n5852) );
  AND2_X1 U7355 ( .A1(n7164), .A2(n9456), .ZN(n10183) );
  NAND2_X1 U7356 ( .A1(n6956), .A2(n10183), .ZN(n5849) );
  OR2_X1 U7357 ( .A1(n5852), .A2(n5849), .ZN(n5843) );
  INV_X1 U7358 ( .A(n5844), .ZN(n5846) );
  NAND2_X1 U7359 ( .A1(n7312), .A2(n9446), .ZN(n6957) );
  AND3_X1 U7360 ( .A1(n6957), .A2(n7743), .A3(n6710), .ZN(n5845) );
  OAI21_X1 U7361 ( .B1(n6960), .B2(n5846), .A(n5845), .ZN(n5847) );
  NAND2_X1 U7362 ( .A1(n5847), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5851) );
  NOR2_X1 U7363 ( .A1(n9452), .A2(n10178), .ZN(n5848) );
  AND2_X1 U7364 ( .A1(n9671), .A2(n5848), .ZN(n7360) );
  NAND2_X1 U7365 ( .A1(n7360), .A2(n6956), .ZN(n9461) );
  NAND2_X1 U7366 ( .A1(n9461), .A2(n5849), .ZN(n5850) );
  NAND2_X1 U7367 ( .A1(n5852), .A2(n5850), .ZN(n6958) );
  AND2_X2 U7368 ( .A1(n5851), .A2(n6958), .ZN(n9158) );
  OR2_X1 U7369 ( .A1(n5852), .A2(n9461), .ZN(n5862) );
  INV_X1 U7370 ( .A(n5862), .ZN(n5854) );
  INV_X1 U7371 ( .A(n5853), .ZN(n7159) );
  NAND2_X1 U7372 ( .A1(n5854), .A2(n7159), .ZN(n9161) );
  INV_X1 U7373 ( .A(n9161), .ZN(n9134) );
  AOI22_X1 U7374 ( .A1(n9595), .A2(n9134), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n5864) );
  NAND2_X1 U7375 ( .A1(n8101), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5861) );
  INV_X1 U7376 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5855) );
  OR2_X1 U7377 ( .A1(n5175), .A2(n5855), .ZN(n5860) );
  OR2_X1 U7378 ( .A1(n5856), .A2(n8076), .ZN(n5859) );
  INV_X1 U7379 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n5857) );
  OR2_X1 U7380 ( .A1(n5806), .A2(n5857), .ZN(n5858) );
  INV_X1 U7381 ( .A(n9556), .ZN(n9467) );
  NAND2_X1 U7382 ( .A1(n9467), .A2(n10469), .ZN(n5863) );
  OAI211_X1 U7383 ( .C1(n9158), .C2(n9560), .A(n5864), .B(n5863), .ZN(n5868)
         );
  NOR3_X1 U7384 ( .A1(n5866), .A2(n9139), .A3(n5865), .ZN(n5867) );
  AOI211_X1 U7385 ( .C1(n9791), .C2(n9165), .A(n5868), .B(n5867), .ZN(n5869)
         );
  INV_X1 U7386 ( .A(n5869), .ZN(n5870) );
  AOI21_X1 U7387 ( .B1(n5876), .B2(n5871), .A(n5870), .ZN(n5872) );
  NAND2_X1 U7388 ( .A1(n5873), .A2(n5872), .ZN(P1_U3218) );
  NAND2_X1 U7389 ( .A1(n9796), .A2(n9165), .ZN(n5881) );
  OAI22_X1 U7390 ( .A1(n9611), .A2(n9161), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5877), .ZN(n5879) );
  NOR2_X1 U7391 ( .A1(n9158), .A2(n9573), .ZN(n5878) );
  AOI211_X1 U7392 ( .C1(n10469), .C2(n8072), .A(n5879), .B(n5878), .ZN(n5880)
         );
  NAND2_X1 U7393 ( .A1(n5885), .A2(n5023), .ZN(n6029) );
  NAND2_X1 U7394 ( .A1(n5900), .A2(n6047), .ZN(n6082) );
  NOR2_X1 U7395 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5888) );
  NOR2_X1 U7396 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5887) );
  NOR2_X1 U7397 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5886) );
  NAND4_X1 U7398 ( .A1(n5896), .A2(n5888), .A3(n5887), .A4(n5886), .ZN(n5889)
         );
  INV_X1 U7399 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5890) );
  INV_X1 U7400 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U7401 ( .A1(n5905), .A2(n5904), .ZN(n5891) );
  INV_X1 U7402 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5892) );
  NOR2_X1 U7403 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5895) );
  NOR2_X1 U7404 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5894) );
  NOR2_X1 U7405 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5893) );
  NAND4_X1 U7406 ( .A1(n5896), .A2(n5895), .A3(n5894), .A4(n5893), .ZN(n5898)
         );
  NAND3_X1 U7407 ( .A1(n6134), .A2(n6106), .A3(n6047), .ZN(n5897) );
  OR2_X1 U7408 ( .A1(n5903), .A2(n6083), .ZN(n5901) );
  XNOR2_X1 U7409 ( .A(n5901), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6682) );
  NAND2_X1 U7410 ( .A1(n5907), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6504) );
  XNOR2_X1 U7411 ( .A(n6504), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6524) );
  OR2_X1 U7412 ( .A1(n6682), .A2(n6524), .ZN(n10333) );
  INV_X1 U7413 ( .A(n10333), .ZN(n6691) );
  INV_X1 U7414 ( .A(n6682), .ZN(n7597) );
  OR2_X1 U7415 ( .A1(n7504), .A2(n7597), .ZN(n7090) );
  NAND3_X1 U7416 ( .A1(n6506), .A2(n6503), .A3(n6519), .ZN(n5906) );
  INV_X1 U7417 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5908) );
  INV_X1 U7418 ( .A(n6512), .ZN(n5910) );
  INV_X1 U7419 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5914) );
  XNOR2_X2 U7420 ( .A(n5912), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5919) );
  XNOR2_X2 U7421 ( .A(n5915), .B(n5914), .ZN(n8487) );
  AND2_X2 U7422 ( .A1(n5919), .A2(n8487), .ZN(n5968) );
  NAND2_X1 U7423 ( .A1(n5968), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5925) );
  OR2_X2 U7424 ( .A1(n5919), .A2(n8487), .ZN(n5953) );
  INV_X1 U7425 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5916) );
  OR2_X1 U7426 ( .A1(n5953), .A2(n5916), .ZN(n5923) );
  INV_X1 U7427 ( .A(n8487), .ZN(n5917) );
  NAND2_X1 U7428 ( .A1(n5919), .A2(n5917), .ZN(n5952) );
  INV_X1 U7429 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5918) );
  INV_X1 U7430 ( .A(n5919), .ZN(n9049) );
  INV_X1 U7431 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5920) );
  OR2_X1 U7432 ( .A1(n5954), .A2(n5920), .ZN(n5921) );
  AND3_X1 U7433 ( .A1(n5923), .A2(n5922), .A3(n5921), .ZN(n5924) );
  NAND2_X1 U7434 ( .A1(n5936), .A2(SI_0_), .ZN(n5926) );
  XNOR2_X1 U7435 ( .A(n5926), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9053) );
  XNOR2_X2 U7436 ( .A(n5927), .B(n5911), .ZN(n6522) );
  INV_X1 U7437 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5928) );
  XNOR2_X2 U7438 ( .A(n5929), .B(n5928), .ZN(n8029) );
  NAND2_X4 U7439 ( .A1(n6522), .A2(n8029), .ZN(n6832) );
  MUX2_X1 U7440 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9053), .S(n6832), .Z(n8107) );
  INV_X1 U7441 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5930) );
  INV_X1 U7442 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7443 ( .A1(n5968), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5933) );
  INV_X1 U7444 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6837) );
  OR2_X1 U7445 ( .A1(n5953), .A2(n6837), .ZN(n5932) );
  AND4_X2 U7446 ( .A1(n5935), .A2(n5934), .A3(n5933), .A4(n5932), .ZN(n6530)
         );
  INV_X1 U7447 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6719) );
  NAND2_X1 U7448 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5938) );
  INV_X1 U7449 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5937) );
  MUX2_X1 U7450 ( .A(n5938), .B(P2_IR_REG_31__SCAN_IN), .S(n5937), .Z(n5940)
         );
  INV_X1 U7451 ( .A(n9909), .ZN(n6718) );
  NAND2_X1 U7452 ( .A1(n7296), .A2(n6475), .ZN(n6356) );
  INV_X1 U7453 ( .A(n6530), .ZN(n5941) );
  NAND2_X1 U7454 ( .A1(n5941), .A2(n10338), .ZN(n6476) );
  INV_X1 U7455 ( .A(n7087), .ZN(n5951) );
  NAND2_X1 U7456 ( .A1(n5968), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5946) );
  INV_X1 U7457 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7201) );
  OR2_X1 U7458 ( .A1(n5952), .A2(n7201), .ZN(n5945) );
  INV_X1 U7459 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6836) );
  OR2_X1 U7460 ( .A1(n5953), .A2(n6836), .ZN(n5944) );
  INV_X1 U7461 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5942) );
  OR2_X1 U7462 ( .A1(n5954), .A2(n5942), .ZN(n5943) );
  INV_X1 U7463 ( .A(n7298), .ZN(n8648) );
  INV_X1 U7464 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5947) );
  XNOR2_X1 U7465 ( .A(n5948), .B(n5947), .ZN(n6845) );
  OR2_X1 U7466 ( .A1(n5961), .A2(n6720), .ZN(n5949) );
  NAND2_X1 U7467 ( .A1(n7298), .A2(n7204), .ZN(n6357) );
  NAND2_X2 U7468 ( .A1(n6353), .A2(n6357), .ZN(n7088) );
  NAND2_X1 U7469 ( .A1(n7085), .A2(n6357), .ZN(n7131) );
  NAND2_X1 U7470 ( .A1(n5968), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5959) );
  OR2_X1 U7471 ( .A1(n5952), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5958) );
  INV_X1 U7472 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6835) );
  OR2_X1 U7473 ( .A1(n5953), .A2(n6835), .ZN(n5957) );
  INV_X1 U7474 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5955) );
  OR2_X1 U7475 ( .A1(n5967), .A2(n5955), .ZN(n5956) );
  NAND4_X1 U7476 ( .A1(n5959), .A2(n5958), .A3(n5957), .A4(n5956), .ZN(n8647)
         );
  OR2_X1 U7477 ( .A1(n5960), .A2(n6729), .ZN(n5965) );
  NAND2_X1 U7478 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4511), .ZN(n5962) );
  XNOR2_X1 U7479 ( .A(n5962), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6848) );
  INV_X1 U7480 ( .A(n6848), .ZN(n6933) );
  OR2_X1 U7481 ( .A1(n6832), .A2(n6933), .ZN(n5963) );
  XNOR2_X1 U7482 ( .A(n8647), .B(n7174), .ZN(n7128) );
  INV_X1 U7483 ( .A(n7128), .ZN(n7130) );
  NAND2_X1 U7484 ( .A1(n7131), .A2(n7130), .ZN(n5966) );
  INV_X1 U7485 ( .A(n8647), .ZN(n7175) );
  INV_X1 U7486 ( .A(n7174), .ZN(n10285) );
  NAND2_X1 U7487 ( .A1(n7175), .A2(n10285), .ZN(n6349) );
  INV_X1 U7488 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6843) );
  OR2_X1 U7489 ( .A1(n6297), .A2(n6843), .ZN(n5973) );
  INV_X2 U7490 ( .A(n5969), .ZN(n6266) );
  XNOR2_X1 U7491 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7260) );
  OR2_X1 U7492 ( .A1(n6266), .A2(n7260), .ZN(n5972) );
  INV_X1 U7493 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5970) );
  OR2_X1 U7494 ( .A1(n6312), .A2(n5970), .ZN(n5971) );
  NOR2_X1 U7495 ( .A1(n5976), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n6003) );
  INV_X1 U7496 ( .A(n6003), .ZN(n5979) );
  NAND2_X1 U7497 ( .A1(n5976), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5977) );
  MUX2_X1 U7498 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5977), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5978) );
  NAND2_X1 U7499 ( .A1(n5979), .A2(n5978), .ZN(n6869) );
  OR2_X1 U7500 ( .A1(n5960), .A2(n6731), .ZN(n5981) );
  OAI211_X1 U7501 ( .C1(n6832), .C2(n6869), .A(n5981), .B(n5980), .ZN(n7262)
         );
  NAND2_X1 U7502 ( .A1(n7460), .A2(n7262), .ZN(n6477) );
  INV_X1 U7503 ( .A(n6477), .ZN(n5982) );
  INV_X1 U7504 ( .A(n7460), .ZN(n8646) );
  INV_X1 U7505 ( .A(n7262), .ZN(n7282) );
  NAND2_X1 U7506 ( .A1(n8646), .A2(n7282), .ZN(n7455) );
  NAND2_X1 U7507 ( .A1(n5968), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5991) );
  INV_X1 U7508 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5983) );
  OR2_X1 U7509 ( .A1(n5967), .A2(n5983), .ZN(n5990) );
  NAND3_X1 U7510 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5996) );
  INV_X1 U7511 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U7512 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5984) );
  NAND2_X1 U7513 ( .A1(n5985), .A2(n5984), .ZN(n5986) );
  NAND2_X1 U7514 ( .A1(n5996), .A2(n5986), .ZN(n7103) );
  OR2_X1 U7515 ( .A1(n6266), .A2(n7103), .ZN(n5989) );
  INV_X1 U7516 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5987) );
  OR2_X1 U7517 ( .A1(n5953), .A2(n5987), .ZN(n5988) );
  OR2_X1 U7518 ( .A1(n6003), .A2(n6083), .ZN(n5992) );
  XNOR2_X1 U7519 ( .A(n5992), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6898) );
  INV_X1 U7520 ( .A(n6898), .ZN(n6722) );
  OR2_X1 U7521 ( .A1(n5960), .A2(n6734), .ZN(n5994) );
  OAI211_X1 U7522 ( .C1(n6832), .C2(n6722), .A(n5994), .B(n5993), .ZN(n10271)
         );
  INV_X1 U7523 ( .A(n10271), .ZN(n7283) );
  NAND2_X1 U7524 ( .A1(n8645), .A2(n7283), .ZN(n6481) );
  AND2_X1 U7525 ( .A1(n7455), .A2(n6481), .ZN(n6345) );
  INV_X1 U7526 ( .A(n8645), .ZN(n7284) );
  NAND2_X1 U7527 ( .A1(n7284), .A2(n10271), .ZN(n6482) );
  INV_X1 U7528 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6894) );
  OR2_X1 U7529 ( .A1(n6297), .A2(n6894), .ZN(n6000) );
  INV_X1 U7530 ( .A(n5996), .ZN(n5995) );
  INV_X1 U7531 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6897) );
  NAND2_X1 U7532 ( .A1(n5996), .A2(n6897), .ZN(n5997) );
  NAND2_X1 U7533 ( .A1(n6010), .A2(n5997), .ZN(n7379) );
  OR2_X1 U7534 ( .A1(n6266), .A2(n7379), .ZN(n5999) );
  INV_X1 U7535 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6903) );
  OR2_X1 U7536 ( .A1(n5953), .A2(n6903), .ZN(n5998) );
  NAND2_X1 U7537 ( .A1(n6003), .A2(n6002), .ZN(n6016) );
  NAND2_X1 U7538 ( .A1(n6016), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6004) );
  XNOR2_X1 U7539 ( .A(n6004), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6915) );
  INV_X1 U7540 ( .A(n6915), .ZN(n6908) );
  OAI211_X1 U7541 ( .C1(n6832), .C2(n6908), .A(n6006), .B(n6005), .ZN(n10346)
         );
  NAND2_X1 U7542 ( .A1(n6559), .A2(n10346), .ZN(n6368) );
  INV_X1 U7543 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6912) );
  OR2_X1 U7544 ( .A1(n6297), .A2(n6912), .ZN(n6014) );
  INV_X1 U7545 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7546 ( .A1(n6010), .A2(n6009), .ZN(n6011) );
  NAND2_X1 U7547 ( .A1(n6023), .A2(n6011), .ZN(n7637) );
  OR2_X1 U7548 ( .A1(n6266), .A2(n7637), .ZN(n6013) );
  INV_X1 U7549 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6918) );
  OR2_X1 U7550 ( .A1(n5953), .A2(n6918), .ZN(n6012) );
  OAI21_X1 U7551 ( .B1(n6016), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6017) );
  XNOR2_X1 U7552 ( .A(n6017), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6968) );
  AOI22_X1 U7553 ( .A1(n6176), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6175), .B2(
        n6968), .ZN(n6019) );
  INV_X2 U7554 ( .A(n5960), .ZN(n6291) );
  NAND2_X1 U7555 ( .A1(n6743), .A2(n6291), .ZN(n6018) );
  NAND2_X1 U7556 ( .A1(n6019), .A2(n6018), .ZN(n7639) );
  NAND2_X1 U7557 ( .A1(n7573), .A2(n7639), .ZN(n6370) );
  INV_X1 U7558 ( .A(n6370), .ZN(n6020) );
  INV_X1 U7559 ( .A(n7573), .ZN(n8643) );
  NAND2_X1 U7560 ( .A1(n8643), .A2(n10351), .ZN(n6371) );
  INV_X1 U7561 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7578) );
  OR2_X1 U7562 ( .A1(n6297), .A2(n7578), .ZN(n6027) );
  INV_X1 U7563 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U7564 ( .A1(n6023), .A2(n6022), .ZN(n6024) );
  NAND2_X1 U7565 ( .A1(n6040), .A2(n6024), .ZN(n7577) );
  OR2_X1 U7566 ( .A1(n6266), .A2(n7577), .ZN(n6026) );
  INV_X1 U7567 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6975) );
  OR2_X1 U7568 ( .A1(n6312), .A2(n6975), .ZN(n6025) );
  NAND2_X1 U7569 ( .A1(n6747), .A2(n6291), .ZN(n6034) );
  NAND2_X1 U7570 ( .A1(n6029), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6030) );
  MUX2_X1 U7571 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6030), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n6031) );
  INV_X1 U7572 ( .A(n6031), .ZN(n6032) );
  NOR2_X1 U7573 ( .A1(n6032), .A2(n6035), .ZN(n7064) );
  AOI22_X1 U7574 ( .A1(n6176), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6175), .B2(
        n7064), .ZN(n6033) );
  NAND2_X1 U7575 ( .A1(n6034), .A2(n6033), .ZN(n7672) );
  NAND2_X1 U7576 ( .A1(n7644), .A2(n7672), .ZN(n6377) );
  INV_X1 U7577 ( .A(n7672), .ZN(n10359) );
  NAND2_X1 U7578 ( .A1(n10359), .A2(n8642), .ZN(n6376) );
  NAND2_X1 U7579 ( .A1(n7570), .A2(n6377), .ZN(n6046) );
  NAND2_X1 U7580 ( .A1(n6758), .A2(n6291), .ZN(n6037) );
  OR2_X1 U7581 ( .A1(n6035), .A2(n6083), .ZN(n6048) );
  XNOR2_X1 U7582 ( .A(n6048), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7112) );
  AOI22_X1 U7583 ( .A1(n6176), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6175), .B2(
        n7112), .ZN(n6036) );
  NAND2_X1 U7584 ( .A1(n6037), .A2(n6036), .ZN(n7708) );
  NAND2_X1 U7585 ( .A1(n5968), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6045) );
  INV_X1 U7586 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6038) );
  OR2_X1 U7587 ( .A1(n5967), .A2(n6038), .ZN(n6044) );
  INV_X1 U7588 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7589 ( .A1(n6040), .A2(n6039), .ZN(n6041) );
  NAND2_X1 U7590 ( .A1(n6056), .A2(n6041), .ZN(n7686) );
  OR2_X1 U7591 ( .A1(n6266), .A2(n7686), .ZN(n6043) );
  INV_X1 U7592 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7070) );
  OR2_X1 U7593 ( .A1(n5953), .A2(n7070), .ZN(n6042) );
  OR2_X1 U7594 ( .A1(n7708), .A2(n7664), .ZN(n6385) );
  NAND2_X1 U7595 ( .A1(n7708), .A2(n7664), .ZN(n6381) );
  NAND2_X1 U7596 ( .A1(n6046), .A2(n7680), .ZN(n7682) );
  NAND2_X1 U7597 ( .A1(n7682), .A2(n6381), .ZN(n6063) );
  NAND2_X1 U7598 ( .A1(n6762), .A2(n6291), .ZN(n6054) );
  NAND2_X1 U7599 ( .A1(n6048), .A2(n6047), .ZN(n6049) );
  NAND2_X1 U7600 ( .A1(n6049), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6051) );
  INV_X1 U7601 ( .A(n6051), .ZN(n6050) );
  NAND2_X1 U7602 ( .A1(n6050), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n6052) );
  INV_X1 U7603 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7604 ( .A1(n6051), .A2(n6079), .ZN(n6064) );
  AND2_X1 U7605 ( .A1(n6052), .A2(n6064), .ZN(n7236) );
  AOI22_X1 U7606 ( .A1(n6176), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6175), .B2(
        n7236), .ZN(n6053) );
  NAND2_X1 U7607 ( .A1(n6054), .A2(n6053), .ZN(n7724) );
  INV_X1 U7608 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7719) );
  OR2_X1 U7609 ( .A1(n6297), .A2(n7719), .ZN(n6061) );
  INV_X1 U7610 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7611 ( .A1(n6056), .A2(n6055), .ZN(n6057) );
  NAND2_X1 U7612 ( .A1(n6071), .A2(n6057), .ZN(n7718) );
  OR2_X1 U7613 ( .A1(n6266), .A2(n7718), .ZN(n6060) );
  INV_X1 U7614 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6058) );
  OR2_X1 U7615 ( .A1(n6312), .A2(n6058), .ZN(n6059) );
  OR2_X1 U7616 ( .A1(n7724), .A2(n7754), .ZN(n6382) );
  NAND2_X1 U7617 ( .A1(n7724), .A2(n7754), .ZN(n7750) );
  NAND2_X1 U7618 ( .A1(n6063), .A2(n7755), .ZN(n7713) );
  NAND2_X1 U7619 ( .A1(n6769), .A2(n6291), .ZN(n6067) );
  NAND2_X1 U7620 ( .A1(n6064), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6065) );
  XNOR2_X1 U7621 ( .A(n6065), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7551) );
  AOI22_X1 U7622 ( .A1(n6176), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6175), .B2(
        n7551), .ZN(n6066) );
  NAND2_X1 U7623 ( .A1(n5968), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6077) );
  INV_X1 U7624 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n6068) );
  OR2_X1 U7625 ( .A1(n5967), .A2(n6068), .ZN(n6076) );
  INV_X1 U7626 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7627 ( .A1(n6071), .A2(n6070), .ZN(n6072) );
  NAND2_X1 U7628 ( .A1(n6088), .A2(n6072), .ZN(n7760) );
  OR2_X1 U7629 ( .A1(n6266), .A2(n7760), .ZN(n6075) );
  INV_X1 U7630 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6073) );
  OR2_X1 U7631 ( .A1(n5953), .A2(n6073), .ZN(n6074) );
  NAND2_X1 U7632 ( .A1(n7877), .A2(n7889), .ZN(n6391) );
  NAND2_X1 U7633 ( .A1(n6824), .A2(n6291), .ZN(n6086) );
  INV_X1 U7634 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7635 ( .A1(n6080), .A2(n6079), .ZN(n6081) );
  NOR2_X1 U7636 ( .A1(n6082), .A2(n6081), .ZN(n6095) );
  OR2_X1 U7637 ( .A1(n6095), .A2(n6083), .ZN(n6084) );
  XNOR2_X1 U7638 ( .A(n6084), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7603) );
  AOI22_X1 U7639 ( .A1(n6176), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6175), .B2(
        n7603), .ZN(n6085) );
  INV_X1 U7640 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7884) );
  OR2_X1 U7641 ( .A1(n6297), .A2(n7884), .ZN(n6092) );
  INV_X1 U7642 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7544) );
  OR2_X1 U7643 ( .A1(n6312), .A2(n7544), .ZN(n6091) );
  INV_X1 U7644 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U7645 ( .A1(n6088), .A2(n7770), .ZN(n6089) );
  NAND2_X1 U7646 ( .A1(n6099), .A2(n6089), .ZN(n7883) );
  OR2_X1 U7647 ( .A1(n6266), .A2(n7883), .ZN(n6090) );
  NAND2_X1 U7648 ( .A1(n10386), .A2(n7976), .ZN(n6392) );
  NAND2_X1 U7649 ( .A1(n6892), .A2(n6291), .ZN(n6097) );
  INV_X1 U7650 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7651 ( .A1(n6095), .A2(n6094), .ZN(n6136) );
  NAND2_X1 U7652 ( .A1(n6136), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6107) );
  XNOR2_X1 U7653 ( .A(n6107), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7734) );
  AOI22_X1 U7654 ( .A1(n6176), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6175), .B2(
        n7734), .ZN(n6096) );
  INV_X1 U7655 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n6098) );
  OR2_X1 U7656 ( .A1(n5967), .A2(n6098), .ZN(n6104) );
  INV_X1 U7657 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7981) );
  OR2_X1 U7658 ( .A1(n6297), .A2(n7981), .ZN(n6103) );
  INV_X1 U7659 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7607) );
  NAND2_X1 U7660 ( .A1(n6099), .A2(n7607), .ZN(n6100) );
  NAND2_X1 U7661 ( .A1(n6113), .A2(n6100), .ZN(n7980) );
  OR2_X1 U7662 ( .A1(n6266), .A2(n7980), .ZN(n6102) );
  INV_X1 U7663 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7728) );
  OR2_X1 U7664 ( .A1(n5953), .A2(n7728), .ZN(n6101) );
  OR2_X1 U7665 ( .A1(n8114), .A2(n8115), .ZN(n6402) );
  NAND2_X1 U7666 ( .A1(n8114), .A2(n8115), .ZN(n6401) );
  INV_X1 U7667 ( .A(n7971), .ZN(n7974) );
  NAND2_X1 U7668 ( .A1(n6952), .A2(n6291), .ZN(n6110) );
  NAND2_X1 U7669 ( .A1(n6107), .A2(n6106), .ZN(n6108) );
  NAND2_X1 U7670 ( .A1(n6108), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6123) );
  XNOR2_X1 U7671 ( .A(n6123), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7866) );
  AOI22_X1 U7672 ( .A1(n6176), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6175), .B2(
        n7866), .ZN(n6109) );
  NAND2_X1 U7673 ( .A1(n5968), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6119) );
  INV_X1 U7674 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6111) );
  OR2_X1 U7675 ( .A1(n6312), .A2(n6111), .ZN(n6118) );
  INV_X1 U7676 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8290) );
  NAND2_X1 U7677 ( .A1(n6113), .A2(n8290), .ZN(n6114) );
  NAND2_X1 U7678 ( .A1(n6145), .A2(n6114), .ZN(n9970) );
  OR2_X1 U7679 ( .A1(n6266), .A2(n9970), .ZN(n6117) );
  INV_X1 U7680 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n6115) );
  OR2_X1 U7681 ( .A1(n5967), .A2(n6115), .ZN(n6116) );
  NAND4_X1 U7682 ( .A1(n6119), .A2(n6118), .A3(n6117), .A4(n6116), .ZN(n8929)
         );
  NAND2_X1 U7683 ( .A1(n9972), .A2(n8929), .ZN(n6120) );
  NAND2_X1 U7684 ( .A1(n8117), .A2(n6120), .ZN(n9975) );
  INV_X1 U7685 ( .A(n8929), .ZN(n8018) );
  OR2_X1 U7686 ( .A1(n9972), .A2(n8018), .ZN(n6121) );
  NAND2_X1 U7687 ( .A1(n7016), .A2(n6291), .ZN(n6127) );
  INV_X1 U7688 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U7689 ( .A1(n6123), .A2(n6122), .ZN(n6124) );
  NAND2_X1 U7690 ( .A1(n6124), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6125) );
  XNOR2_X1 U7691 ( .A(n6125), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7993) );
  AOI22_X1 U7692 ( .A1(n6176), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6175), .B2(
        n7993), .ZN(n6126) );
  INV_X1 U7693 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6143) );
  XNOR2_X1 U7694 ( .A(n6145), .B(n6143), .ZN(n8921) );
  OR2_X1 U7695 ( .A1(n6266), .A2(n8921), .ZN(n6132) );
  INV_X1 U7696 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n6128) );
  OR2_X1 U7697 ( .A1(n6297), .A2(n6128), .ZN(n6131) );
  INV_X1 U7698 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6129) );
  OR2_X1 U7699 ( .A1(n5953), .A2(n6129), .ZN(n6130) );
  NAND2_X1 U7700 ( .A1(n9016), .A2(n8576), .ZN(n6406) );
  INV_X1 U7701 ( .A(n6407), .ZN(n6337) );
  NAND2_X1 U7702 ( .A1(n7006), .A2(n6291), .ZN(n6141) );
  INV_X1 U7703 ( .A(n6134), .ZN(n6135) );
  OR3_X1 U7704 ( .A1(n6136), .A2(P2_IR_REG_13__SCAN_IN), .A3(n6135), .ZN(n6138) );
  NAND2_X1 U7705 ( .A1(n6138), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6137) );
  MUX2_X1 U7706 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6137), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6139) );
  OR2_X1 U7707 ( .A1(n6138), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n6151) );
  AND2_X1 U7708 ( .A1(n6139), .A2(n6151), .ZN(n8652) );
  AOI22_X1 U7709 ( .A1(n6176), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6175), .B2(
        n8652), .ZN(n6140) );
  NAND2_X1 U7710 ( .A1(n5968), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6150) );
  INV_X1 U7711 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8657) );
  OR2_X1 U7712 ( .A1(n5953), .A2(n8657), .ZN(n6149) );
  INV_X1 U7713 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6142) );
  OAI21_X1 U7714 ( .B1(n6145), .B2(n6143), .A(n6142), .ZN(n6146) );
  NAND2_X1 U7715 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n6144) );
  NAND2_X1 U7716 ( .A1(n6146), .A2(n6157), .ZN(n8913) );
  OR2_X1 U7717 ( .A1(n6266), .A2(n8913), .ZN(n6148) );
  INV_X1 U7718 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8329) );
  OR2_X1 U7719 ( .A1(n5967), .A2(n8329), .ZN(n6147) );
  OR2_X1 U7720 ( .A1(n9010), .A2(n8885), .ZN(n6334) );
  NAND2_X1 U7721 ( .A1(n9010), .A2(n8885), .ZN(n8880) );
  NAND2_X1 U7722 ( .A1(n7108), .A2(n6291), .ZN(n6154) );
  NAND2_X1 U7723 ( .A1(n6151), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6152) );
  XNOR2_X1 U7724 ( .A(n6152), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8678) );
  AOI22_X1 U7725 ( .A1(n6176), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6175), .B2(
        n8678), .ZN(n6153) );
  NAND2_X1 U7726 ( .A1(n5968), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6162) );
  INV_X1 U7727 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n6155) );
  OR2_X1 U7728 ( .A1(n5967), .A2(n6155), .ZN(n6161) );
  INV_X1 U7729 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8665) );
  NAND2_X1 U7730 ( .A1(n6157), .A2(n8665), .ZN(n6158) );
  NAND2_X1 U7731 ( .A1(n6169), .A2(n6158), .ZN(n8894) );
  OR2_X1 U7732 ( .A1(n6266), .A2(n8894), .ZN(n6160) );
  INV_X1 U7733 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8656) );
  OR2_X1 U7734 ( .A1(n6312), .A2(n8656), .ZN(n6159) );
  NAND2_X1 U7735 ( .A1(n9005), .A2(n8869), .ZN(n6414) );
  NAND2_X1 U7736 ( .A1(n8864), .A2(n6414), .ZN(n8891) );
  INV_X1 U7737 ( .A(n8880), .ZN(n6336) );
  NOR2_X1 U7738 ( .A1(n8891), .A2(n6336), .ZN(n6163) );
  NAND2_X1 U7739 ( .A1(n7270), .A2(n6291), .ZN(n6166) );
  XNOR2_X1 U7740 ( .A(n6164), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8679) );
  AOI22_X1 U7741 ( .A1(n6176), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6175), .B2(
        n8679), .ZN(n6165) );
  NAND2_X1 U7742 ( .A1(n6294), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6174) );
  INV_X1 U7743 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n6167) );
  OR2_X1 U7744 ( .A1(n5967), .A2(n6167), .ZN(n6173) );
  INV_X1 U7745 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8873) );
  OR2_X1 U7746 ( .A1(n6297), .A2(n8873), .ZN(n6172) );
  INV_X1 U7747 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7748 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  NAND2_X1 U7749 ( .A1(n6181), .A2(n6170), .ZN(n8872) );
  OR2_X1 U7750 ( .A1(n6266), .A2(n8872), .ZN(n6171) );
  OR2_X1 U7751 ( .A1(n4584), .A2(n8887), .ZN(n6474) );
  AND2_X1 U7752 ( .A1(n6474), .A2(n8864), .ZN(n6338) );
  NAND2_X1 U7753 ( .A1(n8881), .A2(n6338), .ZN(n8851) );
  NAND2_X1 U7754 ( .A1(n4584), .A2(n8887), .ZN(n8849) );
  NAND2_X1 U7755 ( .A1(n8851), .A2(n8849), .ZN(n6187) );
  NAND2_X1 U7756 ( .A1(n7352), .A2(n6291), .ZN(n6178) );
  AOI22_X1 U7757 ( .A1(n6176), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n4831), .B2(
        n6175), .ZN(n6177) );
  INV_X1 U7758 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8858) );
  OR2_X1 U7759 ( .A1(n6297), .A2(n8858), .ZN(n6185) );
  INV_X1 U7760 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8694) );
  OR2_X1 U7761 ( .A1(n5953), .A2(n8694), .ZN(n6184) );
  INV_X1 U7762 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7763 ( .A1(n6181), .A2(n6180), .ZN(n6182) );
  NAND2_X1 U7764 ( .A1(n6192), .A2(n6182), .ZN(n8857) );
  OR2_X1 U7765 ( .A1(n6266), .A2(n8857), .ZN(n6183) );
  NAND4_X1 U7766 ( .A1(n6186), .A2(n6185), .A3(n6184), .A4(n6183), .ZN(n8867)
         );
  INV_X1 U7767 ( .A(n8867), .ZN(n8613) );
  OR2_X1 U7768 ( .A1(n8994), .A2(n8613), .ZN(n6422) );
  NAND2_X1 U7769 ( .A1(n8994), .A2(n8613), .ZN(n8837) );
  NAND2_X1 U7770 ( .A1(n6187), .A2(n8848), .ZN(n8836) );
  NAND2_X1 U7771 ( .A1(n7465), .A2(n6291), .ZN(n6189) );
  NAND2_X1 U7772 ( .A1(n5968), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7773 ( .A1(n6294), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6190) );
  AND2_X1 U7774 ( .A1(n6191), .A2(n6190), .ZN(n6196) );
  INV_X1 U7775 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U7776 ( .A1(n6192), .A2(n8594), .ZN(n6193) );
  AND2_X1 U7777 ( .A1(n6201), .A2(n6193), .ZN(n8833) );
  NAND2_X1 U7778 ( .A1(n8833), .A2(n5969), .ZN(n6195) );
  NAND2_X1 U7779 ( .A1(n8987), .A2(n8548), .ZN(n6424) );
  NAND2_X1 U7780 ( .A1(n6423), .A2(n6424), .ZN(n8839) );
  INV_X1 U7781 ( .A(n8837), .ZN(n6420) );
  NOR2_X1 U7782 ( .A1(n8839), .A2(n6420), .ZN(n6197) );
  NAND2_X1 U7783 ( .A1(n7594), .A2(n6291), .ZN(n6199) );
  INV_X1 U7784 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U7785 ( .A1(n6201), .A2(n8546), .ZN(n6202) );
  NAND2_X1 U7786 ( .A1(n6209), .A2(n6202), .ZN(n8820) );
  OR2_X1 U7787 ( .A1(n8820), .A2(n6266), .ZN(n6205) );
  AOI22_X1 U7788 ( .A1(n6294), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n5968), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U7789 ( .A1(n8982), .A2(n8812), .ZN(n8808) );
  NAND2_X1 U7790 ( .A1(n6429), .A2(n8808), .ZN(n8824) );
  NAND2_X1 U7791 ( .A1(n7656), .A2(n6291), .ZN(n6208) );
  INV_X1 U7792 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U7793 ( .A1(n6209), .A2(n8604), .ZN(n6210) );
  NAND2_X1 U7794 ( .A1(n6221), .A2(n6210), .ZN(n8804) );
  OR2_X1 U7795 ( .A1(n8804), .A2(n6266), .ZN(n6216) );
  INV_X1 U7796 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6213) );
  NAND2_X1 U7797 ( .A1(n5968), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6211) );
  OAI211_X1 U7798 ( .C1(n6213), .C2(n6312), .A(n6212), .B(n6211), .ZN(n6214)
         );
  INV_X1 U7799 ( .A(n6214), .ZN(n6215) );
  NAND2_X1 U7800 ( .A1(n8977), .A2(n8547), .ZN(n6434) );
  INV_X1 U7801 ( .A(n8808), .ZN(n6217) );
  NOR2_X1 U7802 ( .A1(n8811), .A2(n6217), .ZN(n6218) );
  NAND2_X1 U7803 ( .A1(n7746), .A2(n6291), .ZN(n6220) );
  INV_X1 U7804 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8511) );
  NAND2_X1 U7805 ( .A1(n6221), .A2(n8511), .ZN(n6222) );
  AND2_X1 U7806 ( .A1(n6230), .A2(n6222), .ZN(n8795) );
  INV_X1 U7807 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U7808 ( .A1(n6294), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U7809 ( .A1(n5968), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6223) );
  OAI211_X1 U7810 ( .C1(n5967), .C2(n8200), .A(n6224), .B(n6223), .ZN(n6225)
         );
  AOI21_X1 U7811 ( .B1(n8795), .B2(n5969), .A(n6225), .ZN(n8813) );
  OR2_X1 U7812 ( .A1(n8972), .A2(n8813), .ZN(n6441) );
  NAND2_X1 U7813 ( .A1(n8972), .A2(n8813), .ZN(n6440) );
  NAND2_X1 U7814 ( .A1(n6441), .A2(n6440), .ZN(n8791) );
  INV_X1 U7815 ( .A(n6435), .ZN(n8786) );
  NOR2_X1 U7816 ( .A1(n8791), .A2(n8786), .ZN(n6226) );
  NAND2_X1 U7817 ( .A1(n8787), .A2(n6440), .ZN(n8776) );
  NAND2_X1 U7818 ( .A1(n7775), .A2(n6291), .ZN(n6228) );
  INV_X1 U7819 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8587) );
  NAND2_X1 U7820 ( .A1(n6230), .A2(n8587), .ZN(n6231) );
  NAND2_X1 U7821 ( .A1(n6242), .A2(n6231), .ZN(n8781) );
  OR2_X1 U7822 ( .A1(n8781), .A2(n6266), .ZN(n6237) );
  INV_X1 U7823 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U7824 ( .A1(n5968), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6233) );
  NAND2_X1 U7825 ( .A1(n6294), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6232) );
  OAI211_X1 U7826 ( .C1(n6234), .C2(n5967), .A(n6233), .B(n6232), .ZN(n6235)
         );
  INV_X1 U7827 ( .A(n6235), .ZN(n6236) );
  NAND2_X1 U7828 ( .A1(n6237), .A2(n6236), .ZN(n8789) );
  NAND2_X1 U7829 ( .A1(n8966), .A2(n8789), .ZN(n6238) );
  INV_X1 U7830 ( .A(n8771), .ZN(n8775) );
  OR2_X2 U7831 ( .A1(n8776), .A2(n8775), .ZN(n8779) );
  INV_X1 U7832 ( .A(n8789), .ZN(n8512) );
  OR2_X1 U7833 ( .A1(n8966), .A2(n8512), .ZN(n6444) );
  NAND2_X1 U7834 ( .A1(n8779), .A2(n6444), .ZN(n8757) );
  NAND2_X1 U7835 ( .A1(n7914), .A2(n6291), .ZN(n6240) );
  INV_X1 U7836 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U7837 ( .A1(n6242), .A2(n8561), .ZN(n6243) );
  NAND2_X1 U7838 ( .A1(n6252), .A2(n6243), .ZN(n8761) );
  OR2_X1 U7839 ( .A1(n8761), .A2(n6266), .ZN(n6249) );
  INV_X1 U7840 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U7841 ( .A1(n5968), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6244) );
  OAI211_X1 U7842 ( .C1(n6246), .C2(n6312), .A(n6245), .B(n6244), .ZN(n6247)
         );
  INV_X1 U7843 ( .A(n6247), .ZN(n6248) );
  NAND2_X1 U7844 ( .A1(n7920), .A2(n6291), .ZN(n6251) );
  INV_X1 U7845 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U7846 ( .A1(n6252), .A2(n8627), .ZN(n6253) );
  INV_X1 U7847 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n6257) );
  NAND2_X1 U7848 ( .A1(n6294), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6256) );
  INV_X1 U7849 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n6254) );
  OR2_X1 U7850 ( .A1(n5967), .A2(n6254), .ZN(n6255) );
  OAI211_X1 U7851 ( .C1(n6297), .C2(n6257), .A(n6256), .B(n6255), .ZN(n6258)
         );
  INV_X1 U7852 ( .A(n6473), .ZN(n6259) );
  OR2_X1 U7853 ( .A1(n8963), .A2(n8777), .ZN(n8745) );
  AND2_X1 U7854 ( .A1(n6259), .A2(n8745), .ZN(n6333) );
  NAND2_X1 U7855 ( .A1(n8755), .A2(n6333), .ZN(n8731) );
  NAND2_X1 U7856 ( .A1(n7989), .A2(n6291), .ZN(n6261) );
  INV_X1 U7857 ( .A(n6264), .ZN(n6262) );
  NAND2_X1 U7858 ( .A1(n6262), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6278) );
  INV_X1 U7859 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6263) );
  NAND2_X1 U7860 ( .A1(n6264), .A2(n6263), .ZN(n6265) );
  NAND2_X1 U7861 ( .A1(n6278), .A2(n6265), .ZN(n8504) );
  INV_X1 U7862 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U7863 ( .A1(n5968), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U7864 ( .A1(n6294), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6267) );
  OAI211_X1 U7865 ( .C1(n5967), .C2(n6269), .A(n6268), .B(n6267), .ZN(n6270)
         );
  INV_X1 U7866 ( .A(n6270), .ZN(n6271) );
  INV_X1 U7867 ( .A(n8733), .ZN(n6273) );
  INV_X1 U7868 ( .A(n6472), .ZN(n8730) );
  AND2_X1 U7869 ( .A1(n6273), .A2(n8730), .ZN(n6274) );
  NAND2_X1 U7870 ( .A1(n8731), .A2(n6274), .ZN(n6275) );
  OR2_X1 U7871 ( .A1(n8951), .A2(n8626), .ZN(n6449) );
  NAND2_X1 U7872 ( .A1(n8015), .A2(n6291), .ZN(n6277) );
  INV_X1 U7873 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8013) );
  INV_X1 U7874 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U7875 ( .A1(n6278), .A2(n6703), .ZN(n6279) );
  NAND2_X1 U7876 ( .A1(n8490), .A2(n5969), .ZN(n6285) );
  INV_X1 U7877 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6282) );
  NAND2_X1 U7878 ( .A1(n6294), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6280) );
  OAI211_X1 U7879 ( .C1(n6297), .C2(n6282), .A(n6281), .B(n6280), .ZN(n6283)
         );
  INV_X1 U7880 ( .A(n6283), .ZN(n6284) );
  INV_X1 U7881 ( .A(n6288), .ZN(n6289) );
  NAND2_X1 U7882 ( .A1(n6289), .A2(n8388), .ZN(n6290) );
  INV_X1 U7883 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8486) );
  INV_X1 U7884 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9902) );
  MUX2_X1 U7885 ( .A(n8486), .B(n9902), .S(n6724), .Z(n6304) );
  XNOR2_X1 U7886 ( .A(n6304), .B(SI_29_), .ZN(n6301) );
  NAND2_X1 U7887 ( .A1(n8485), .A2(n6291), .ZN(n6293) );
  INV_X1 U7888 ( .A(n8714), .ZN(n6299) );
  INV_X1 U7889 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U7890 ( .A1(n6294), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6296) );
  INV_X1 U7891 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8201) );
  OR2_X1 U7892 ( .A1(n5967), .A2(n8201), .ZN(n6295) );
  OAI211_X1 U7893 ( .C1(n6297), .C2(n8713), .A(n6296), .B(n6295), .ZN(n6298)
         );
  AOI21_X1 U7894 ( .B1(n6299), .B2(n5969), .A(n6298), .ZN(n8495) );
  NAND2_X1 U7895 ( .A1(n8716), .A2(n8495), .ZN(n6460) );
  INV_X1 U7896 ( .A(n8133), .ZN(n6300) );
  INV_X1 U7897 ( .A(n6313), .ZN(n6315) );
  INV_X1 U7898 ( .A(SI_29_), .ZN(n6303) );
  INV_X1 U7899 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9051) );
  INV_X1 U7900 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9172) );
  MUX2_X1 U7901 ( .A(n9051), .B(n9172), .S(n6724), .Z(n6318) );
  INV_X1 U7902 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U7903 ( .A1(n5968), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6307) );
  OAI211_X1 U7904 ( .C1(n6312), .C2(n8198), .A(n6307), .B(n6306), .ZN(n8635)
         );
  AND2_X1 U7905 ( .A1(n8945), .A2(n8635), .ZN(n6330) );
  INV_X1 U7906 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U7907 ( .A1(n5968), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6310) );
  INV_X1 U7908 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6308) );
  OR2_X1 U7909 ( .A1(n5967), .A2(n6308), .ZN(n6309) );
  OAI211_X1 U7910 ( .C1(n6312), .C2(n6311), .A(n6310), .B(n6309), .ZN(n8032)
         );
  OAI22_X1 U7911 ( .A1(n6313), .A2(n6330), .B1(n7597), .B2(n8032), .ZN(n6314)
         );
  OAI21_X1 U7912 ( .B1(n6315), .B2(n8709), .A(n6314), .ZN(n6327) );
  INV_X1 U7913 ( .A(SI_30_), .ZN(n6316) );
  NAND2_X1 U7914 ( .A1(n6321), .A2(n6320), .ZN(n6324) );
  MUX2_X1 U7915 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6724), .Z(n6322) );
  XNOR2_X1 U7916 ( .A(n6322), .B(SI_31_), .ZN(n6323) );
  NAND2_X1 U7917 ( .A1(n8941), .A2(n8032), .ZN(n6469) );
  INV_X1 U7918 ( .A(n8635), .ZN(n6326) );
  NAND2_X1 U7919 ( .A1(n8709), .A2(n6326), .ZN(n6461) );
  XNOR2_X1 U7920 ( .A(n6328), .B(n4831), .ZN(n6329) );
  NOR2_X1 U7921 ( .A1(n6524), .A2(n7597), .ZN(n6331) );
  AOI21_X1 U7922 ( .B1(n8777), .B2(n8963), .A(n6472), .ZN(n6332) );
  MUX2_X1 U7923 ( .A(n6333), .B(n6332), .S(n6467), .Z(n6448) );
  NAND2_X1 U7924 ( .A1(n8864), .A2(n6334), .ZN(n6335) );
  MUX2_X1 U7925 ( .A(n6336), .B(n6335), .S(n4618), .Z(n6413) );
  OAI211_X1 U7926 ( .C1(n6413), .C2(n6406), .A(n8849), .B(n6414), .ZN(n6341)
         );
  NAND2_X1 U7927 ( .A1(n6414), .A2(n6337), .ZN(n6339) );
  OAI21_X1 U7928 ( .B1(n6413), .B2(n6339), .A(n6338), .ZN(n6340) );
  MUX2_X1 U7929 ( .A(n6341), .B(n6340), .S(n6467), .Z(n6342) );
  INV_X1 U7930 ( .A(n6342), .ZN(n6416) );
  NAND2_X1 U7931 ( .A1(n6391), .A2(n7750), .ZN(n6383) );
  AND2_X1 U7932 ( .A1(n6482), .A2(n6477), .ZN(n6343) );
  MUX2_X1 U7933 ( .A(n6345), .B(n6343), .S(n4618), .Z(n6361) );
  INV_X1 U7934 ( .A(n6361), .ZN(n6344) );
  NAND2_X1 U7935 ( .A1(n6344), .A2(n6481), .ZN(n6348) );
  OAI21_X1 U7936 ( .B1(n7175), .B2(n10285), .A(n6345), .ZN(n6347) );
  AOI21_X1 U7937 ( .B1(n6348), .B2(n6347), .A(n6346), .ZN(n6367) );
  NAND2_X1 U7938 ( .A1(n6477), .A2(n6349), .ZN(n6351) );
  NAND2_X1 U7939 ( .A1(n6368), .A2(n6482), .ZN(n6350) );
  AOI21_X1 U7940 ( .B1(n6361), .B2(n6351), .A(n6350), .ZN(n6364) );
  INV_X1 U7941 ( .A(n8107), .ZN(n10334) );
  NAND2_X1 U7942 ( .A1(n8650), .A2(n10334), .ZN(n6478) );
  NAND2_X1 U7943 ( .A1(n6476), .A2(n6478), .ZN(n6352) );
  NAND3_X1 U7944 ( .A1(n6357), .A2(n6475), .A3(n6352), .ZN(n6354) );
  NAND2_X1 U7945 ( .A1(n6354), .A2(n6353), .ZN(n6360) );
  AND2_X1 U7946 ( .A1(n6478), .A2(n6682), .ZN(n6355) );
  OAI211_X1 U7947 ( .C1(n6356), .C2(n6355), .A(n6353), .B(n6476), .ZN(n6358)
         );
  NAND2_X1 U7948 ( .A1(n6358), .A2(n6357), .ZN(n6359) );
  MUX2_X1 U7949 ( .A(n6360), .B(n6359), .S(n6467), .Z(n6362) );
  NAND3_X1 U7950 ( .A1(n6362), .A2(n6361), .A3(n7130), .ZN(n6363) );
  OAI21_X1 U7951 ( .B1(n4618), .B2(n6364), .A(n6363), .ZN(n6365) );
  OAI21_X1 U7952 ( .B1(n6367), .B2(n6467), .A(n6366), .ZN(n6375) );
  OR2_X1 U7953 ( .A1(n6368), .A2(n6467), .ZN(n6369) );
  AND2_X1 U7954 ( .A1(n7641), .A2(n6369), .ZN(n6374) );
  MUX2_X1 U7955 ( .A(n6371), .B(n6370), .S(n6467), .Z(n6372) );
  NAND2_X1 U7956 ( .A1(n6372), .A2(n7572), .ZN(n6373) );
  AOI21_X1 U7957 ( .B1(n6375), .B2(n6374), .A(n6373), .ZN(n6380) );
  INV_X1 U7958 ( .A(n6381), .ZN(n7711) );
  NAND2_X1 U7959 ( .A1(n6385), .A2(n6376), .ZN(n6378) );
  INV_X1 U7960 ( .A(n6377), .ZN(n7679) );
  MUX2_X1 U7961 ( .A(n6378), .B(n7679), .S(n4618), .Z(n6379) );
  OR2_X1 U7962 ( .A1(n6381), .A2(n4618), .ZN(n6384) );
  NAND4_X1 U7963 ( .A1(n6386), .A2(n7755), .A3(n6385), .A4(n6384), .ZN(n6387)
         );
  NAND2_X1 U7964 ( .A1(n6387), .A2(n7887), .ZN(n6398) );
  INV_X1 U7965 ( .A(n6388), .ZN(n6389) );
  NAND2_X1 U7966 ( .A1(n6392), .A2(n6389), .ZN(n6390) );
  AND2_X1 U7967 ( .A1(n6390), .A2(n6393), .ZN(n6396) );
  NAND2_X1 U7968 ( .A1(n6392), .A2(n6391), .ZN(n6394) );
  NAND2_X1 U7969 ( .A1(n6394), .A2(n6393), .ZN(n6395) );
  MUX2_X1 U7970 ( .A(n6396), .B(n6395), .S(n6467), .Z(n6397) );
  OAI21_X1 U7971 ( .B1(n6399), .B2(n6398), .A(n6397), .ZN(n6400) );
  NAND2_X1 U7972 ( .A1(n6400), .A2(n7971), .ZN(n6404) );
  MUX2_X1 U7973 ( .A(n6402), .B(n6401), .S(n6467), .Z(n6403) );
  NAND2_X1 U7974 ( .A1(n6404), .A2(n6403), .ZN(n6409) );
  INV_X1 U7975 ( .A(n9972), .ZN(n9985) );
  MUX2_X1 U7976 ( .A(n8018), .B(n9985), .S(n4618), .Z(n6408) );
  MUX2_X1 U7977 ( .A(n8929), .B(n9972), .S(n6467), .Z(n6405) );
  OAI21_X1 U7978 ( .B1(n6409), .B2(n6408), .A(n6405), .ZN(n6412) );
  MUX2_X1 U7979 ( .A(n6407), .B(n6406), .S(n6467), .Z(n6411) );
  NAND2_X1 U7980 ( .A1(n6409), .A2(n6408), .ZN(n6410) );
  INV_X1 U7981 ( .A(n6413), .ZN(n6415) );
  NAND2_X1 U7982 ( .A1(n6421), .A2(n8849), .ZN(n6417) );
  NAND2_X1 U7983 ( .A1(n6417), .A2(n6422), .ZN(n6418) );
  NAND3_X1 U7984 ( .A1(n6418), .A2(n6424), .A3(n8837), .ZN(n6419) );
  NAND3_X1 U7985 ( .A1(n6419), .A2(n6429), .A3(n6423), .ZN(n6428) );
  AOI21_X1 U7986 ( .B1(n6421), .B2(n6474), .A(n6420), .ZN(n6426) );
  NAND2_X1 U7987 ( .A1(n6423), .A2(n6422), .ZN(n6425) );
  OAI211_X1 U7988 ( .C1(n6426), .C2(n6425), .A(n8808), .B(n6424), .ZN(n6427)
         );
  MUX2_X1 U7989 ( .A(n6428), .B(n6427), .S(n4618), .Z(n6433) );
  NAND2_X1 U7990 ( .A1(n6435), .A2(n6429), .ZN(n6430) );
  NAND2_X1 U7991 ( .A1(n6430), .A2(n4618), .ZN(n6432) );
  INV_X1 U7992 ( .A(n6434), .ZN(n6431) );
  AOI21_X1 U7993 ( .B1(n6433), .B2(n6432), .A(n6431), .ZN(n6439) );
  AOI21_X1 U7994 ( .B1(n6434), .B2(n8808), .A(n4618), .ZN(n6438) );
  NOR2_X1 U7995 ( .A1(n6435), .A2(n4618), .ZN(n6436) );
  NOR2_X1 U7996 ( .A1(n8791), .A2(n6436), .ZN(n6437) );
  OAI21_X1 U7997 ( .B1(n6439), .B2(n6438), .A(n6437), .ZN(n6443) );
  MUX2_X1 U7998 ( .A(n6441), .B(n6440), .S(n6467), .Z(n6442) );
  NAND2_X1 U7999 ( .A1(n8966), .A2(n8512), .ZN(n6445) );
  MUX2_X1 U8000 ( .A(n6445), .B(n6444), .S(n6467), .Z(n6446) );
  MUX2_X1 U8001 ( .A(n6472), .B(n6473), .S(n6467), .Z(n6447) );
  INV_X1 U8002 ( .A(n6455), .ZN(n6454) );
  NAND2_X1 U8003 ( .A1(n6450), .A2(n6449), .ZN(n6452) );
  INV_X1 U8004 ( .A(n8951), .ZN(n8729) );
  NOR2_X1 U8005 ( .A1(n8729), .A2(n8637), .ZN(n6451) );
  MUX2_X1 U8006 ( .A(n6452), .B(n6451), .S(n6467), .Z(n6453) );
  NAND2_X1 U8007 ( .A1(n8492), .A2(n6467), .ZN(n6456) );
  AOI22_X1 U8008 ( .A1(n6456), .A2(n6455), .B1(n8130), .B2(n6467), .ZN(n6457)
         );
  OAI21_X1 U8009 ( .B1(n6458), .B2(n6457), .A(n8133), .ZN(n6464) );
  MUX2_X1 U8010 ( .A(n6460), .B(n6459), .S(n6467), .Z(n6463) );
  INV_X1 U8011 ( .A(n6461), .ZN(n6462) );
  AOI21_X1 U8012 ( .B1(n6464), .B2(n6463), .A(n6462), .ZN(n6465) );
  NOR3_X1 U8013 ( .A1(n6496), .A2(n6468), .A3(n6467), .ZN(n6470) );
  INV_X1 U8014 ( .A(n6524), .ZN(n7661) );
  INV_X1 U8015 ( .A(n7089), .ZN(n6471) );
  INV_X1 U8016 ( .A(n8791), .ZN(n6493) );
  NAND2_X1 U8017 ( .A1(n6474), .A2(n8849), .ZN(n8865) );
  INV_X1 U8018 ( .A(n8905), .ZN(n6489) );
  NOR2_X1 U8019 ( .A1(n7088), .A2(n7081), .ZN(n6480) );
  NAND2_X1 U8020 ( .A1(n6477), .A2(n7455), .ZN(n7178) );
  INV_X1 U8021 ( .A(n7178), .ZN(n7181) );
  NAND2_X1 U8022 ( .A1(n7296), .A2(n6478), .ZN(n10337) );
  NOR2_X1 U8023 ( .A1(n10337), .A2(n7504), .ZN(n6479) );
  NAND4_X1 U8024 ( .A1(n6480), .A2(n7181), .A3(n6479), .A4(n7130), .ZN(n6483)
         );
  NAND2_X1 U8025 ( .A1(n6482), .A2(n6481), .ZN(n7458) );
  NOR3_X1 U8026 ( .A1(n6483), .A2(n7285), .A3(n7458), .ZN(n6484) );
  NAND4_X1 U8027 ( .A1(n6484), .A2(n7680), .A3(n7572), .A4(n7641), .ZN(n6486)
         );
  INV_X1 U8028 ( .A(n7755), .ZN(n6485) );
  NOR4_X1 U8029 ( .A1(n7880), .A2(n7757), .A3(n6486), .A4(n6485), .ZN(n6487)
         );
  NAND4_X1 U8030 ( .A1(n8927), .A2(n7971), .A3(n6487), .A4(n9975), .ZN(n6488)
         );
  NOR4_X1 U8031 ( .A1(n8865), .A2(n8891), .A3(n6489), .A4(n6488), .ZN(n6490)
         );
  NAND2_X1 U8032 ( .A1(n6490), .A2(n8848), .ZN(n6491) );
  NOR4_X1 U8033 ( .A1(n8811), .A2(n8824), .A3(n8839), .A4(n6491), .ZN(n6492)
         );
  NAND4_X1 U8034 ( .A1(n8747), .A2(n6493), .A3(n6492), .A4(n8771), .ZN(n6494)
         );
  NOR4_X1 U8035 ( .A1(n8493), .A2(n6494), .A3(n8733), .A4(n8129), .ZN(n6495)
         );
  NAND4_X1 U8036 ( .A1(n6497), .A2(n6496), .A3(n8133), .A4(n6495), .ZN(n6498)
         );
  XNOR2_X1 U8037 ( .A(n6498), .B(n8701), .ZN(n6499) );
  OAI22_X1 U8038 ( .A1(n6499), .A2(n6682), .B1(n4629), .B2(n7089), .ZN(n6501)
         );
  NAND2_X1 U8039 ( .A1(n6504), .A2(n6503), .ZN(n6505) );
  NAND2_X1 U8040 ( .A1(n6505), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6507) );
  NAND2_X1 U8041 ( .A1(n6507), .A2(n6506), .ZN(n6518) );
  OR2_X1 U8042 ( .A1(n6507), .A2(n6506), .ZN(n6508) );
  NAND2_X1 U8043 ( .A1(n6518), .A2(n6508), .ZN(n6709) );
  OR2_X1 U8044 ( .A1(n6709), .A2(P2_U3152), .ZN(n7747) );
  INV_X1 U8045 ( .A(n7747), .ZN(n6509) );
  OAI21_X1 U8046 ( .B1(n6511), .B2(n6510), .A(n6509), .ZN(n6528) );
  NAND2_X1 U8047 ( .A1(n6512), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6513) );
  MUX2_X1 U8048 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6513), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6514) );
  AND2_X1 U8049 ( .A1(n6515), .A2(n6514), .ZN(n6677) );
  NAND2_X1 U8050 ( .A1(n4559), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6516) );
  MUX2_X1 U8051 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6516), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6517) );
  NAND2_X1 U8052 ( .A1(n6517), .A2(n6512), .ZN(n7916) );
  INV_X1 U8053 ( .A(n7916), .ZN(n6678) );
  NAND2_X1 U8054 ( .A1(n6677), .A2(n6678), .ZN(n6521) );
  NAND2_X1 U8055 ( .A1(n6518), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6520) );
  XNOR2_X1 U8056 ( .A(n6520), .B(n6519), .ZN(n7805) );
  INV_X1 U8057 ( .A(n6522), .ZN(n6523) );
  AND2_X1 U8058 ( .A1(n6524), .A2(n6682), .ZN(n7078) );
  INV_X1 U8059 ( .A(n8928), .ZN(n8884) );
  NAND2_X1 U8060 ( .A1(n7504), .A2(n8701), .ZN(n6699) );
  NOR4_X1 U8061 ( .A1(n10294), .A2(n8884), .A3(n8029), .A4(n6699), .ZN(n6526)
         );
  OAI21_X1 U8062 ( .B1(n7747), .B2(n6524), .A(P2_B_REG_SCAN_IN), .ZN(n6525) );
  NAND2_X1 U8063 ( .A1(n6528), .A2(n6527), .ZN(P2_U3244) );
  NAND2_X1 U8064 ( .A1(n7504), .A2(n6682), .ZN(n7197) );
  NAND3_X1 U8065 ( .A1(n7089), .A2(n7597), .A3(n10333), .ZN(n6529) );
  NAND2_X4 U8066 ( .A1(n7197), .A2(n6529), .ZN(n6649) );
  NAND2_X1 U8067 ( .A1(n8789), .A2(n6612), .ZN(n6639) );
  XNOR2_X1 U8068 ( .A(n8538), .B(n6649), .ZN(n6538) );
  XNOR2_X1 U8069 ( .A(n6540), .B(n6538), .ZN(n8534) );
  INV_X1 U8070 ( .A(n7300), .ZN(n6531) );
  NAND2_X1 U8071 ( .A1(n6531), .A2(n6612), .ZN(n8111) );
  OR2_X1 U8072 ( .A1(n8107), .A2(n6649), .ZN(n6532) );
  NAND2_X1 U8073 ( .A1(n8534), .A2(n8535), .ZN(n8533) );
  INV_X1 U8074 ( .A(n6536), .ZN(n6534) );
  XNOR2_X1 U8075 ( .A(n7204), .B(n6649), .ZN(n6535) );
  INV_X1 U8076 ( .A(n6535), .ZN(n6533) );
  NAND2_X1 U8077 ( .A1(n6534), .A2(n6533), .ZN(n6537) );
  NAND2_X1 U8078 ( .A1(n6536), .A2(n6535), .ZN(n6542) );
  AND2_X1 U8079 ( .A1(n6537), .A2(n6542), .ZN(n6984) );
  INV_X1 U8080 ( .A(n6538), .ZN(n6539) );
  NAND2_X1 U8081 ( .A1(n6540), .A2(n6539), .ZN(n6982) );
  AND2_X1 U8082 ( .A1(n6984), .A2(n6982), .ZN(n6541) );
  NAND2_X1 U8083 ( .A1(n8533), .A2(n6541), .ZN(n6983) );
  NAND2_X1 U8084 ( .A1(n6983), .A2(n6542), .ZN(n8520) );
  AND2_X1 U8085 ( .A1(n8647), .A2(n6612), .ZN(n6543) );
  XNOR2_X1 U8086 ( .A(n7174), .B(n6660), .ZN(n6544) );
  NAND2_X1 U8087 ( .A1(n6543), .A2(n6544), .ZN(n7020) );
  INV_X1 U8088 ( .A(n6543), .ZN(n6546) );
  INV_X1 U8089 ( .A(n6544), .ZN(n6545) );
  NAND2_X1 U8090 ( .A1(n6546), .A2(n6545), .ZN(n6547) );
  NAND2_X1 U8091 ( .A1(n8520), .A2(n8519), .ZN(n8518) );
  OR2_X1 U8092 ( .A1(n7460), .A2(n6570), .ZN(n6551) );
  XNOR2_X1 U8093 ( .A(n7262), .B(n6660), .ZN(n6550) );
  XNOR2_X1 U8094 ( .A(n6551), .B(n6550), .ZN(n7021) );
  INV_X1 U8095 ( .A(n7020), .ZN(n6548) );
  NAND2_X1 U8096 ( .A1(n8518), .A2(n6549), .ZN(n7024) );
  NAND2_X1 U8097 ( .A1(n6551), .A2(n6550), .ZN(n6552) );
  AND2_X1 U8098 ( .A1(n8645), .A2(n6612), .ZN(n6553) );
  XNOR2_X1 U8099 ( .A(n10271), .B(n6649), .ZN(n6554) );
  NAND2_X1 U8100 ( .A1(n6553), .A2(n6554), .ZN(n6558) );
  INV_X1 U8101 ( .A(n6553), .ZN(n6556) );
  INV_X1 U8102 ( .A(n6554), .ZN(n6555) );
  NAND2_X1 U8103 ( .A1(n6556), .A2(n6555), .ZN(n6557) );
  AND2_X1 U8104 ( .A1(n6558), .A2(n6557), .ZN(n7101) );
  OR2_X1 U8105 ( .A1(n6559), .A2(n8108), .ZN(n6562) );
  XNOR2_X1 U8106 ( .A(n10346), .B(n6660), .ZN(n6561) );
  XNOR2_X1 U8107 ( .A(n6562), .B(n6561), .ZN(n7380) );
  INV_X1 U8108 ( .A(n7380), .ZN(n6560) );
  NAND2_X1 U8109 ( .A1(n6562), .A2(n6561), .ZN(n6563) );
  AND2_X1 U8110 ( .A1(n7383), .A2(n6563), .ZN(n7346) );
  NOR2_X1 U8111 ( .A1(n7573), .A2(n8108), .ZN(n6564) );
  XNOR2_X1 U8112 ( .A(n7639), .B(n6649), .ZN(n6565) );
  NAND2_X1 U8113 ( .A1(n6564), .A2(n6565), .ZN(n6569) );
  INV_X1 U8114 ( .A(n6564), .ZN(n6567) );
  INV_X1 U8115 ( .A(n6565), .ZN(n6566) );
  NAND2_X1 U8116 ( .A1(n6567), .A2(n6566), .ZN(n6568) );
  AND2_X1 U8117 ( .A1(n6569), .A2(n6568), .ZN(n7345) );
  NAND2_X1 U8118 ( .A1(n7346), .A2(n7345), .ZN(n7344) );
  NAND2_X1 U8119 ( .A1(n7344), .A2(n6569), .ZN(n7445) );
  XNOR2_X1 U8120 ( .A(n7672), .B(n6649), .ZN(n6572) );
  OR2_X1 U8121 ( .A1(n7644), .A2(n8108), .ZN(n6571) );
  XNOR2_X1 U8122 ( .A(n6572), .B(n6571), .ZN(n7444) );
  NAND2_X1 U8123 ( .A1(n7445), .A2(n7444), .ZN(n7443) );
  INV_X1 U8124 ( .A(n6571), .ZN(n6573) );
  NAND2_X1 U8125 ( .A1(n6573), .A2(n6572), .ZN(n6574) );
  XNOR2_X1 U8126 ( .A(n7708), .B(n6649), .ZN(n6575) );
  NOR2_X1 U8127 ( .A1(n7664), .A2(n8108), .ZN(n6576) );
  INV_X1 U8128 ( .A(n6575), .ZN(n6578) );
  INV_X1 U8129 ( .A(n6576), .ZN(n6577) );
  NAND2_X1 U8130 ( .A1(n6578), .A2(n6577), .ZN(n7584) );
  XNOR2_X1 U8131 ( .A(n7724), .B(n6649), .ZN(n6579) );
  NOR2_X1 U8132 ( .A1(n7754), .A2(n8108), .ZN(n6580) );
  XNOR2_X1 U8133 ( .A(n6579), .B(n6580), .ZN(n7662) );
  INV_X1 U8134 ( .A(n6579), .ZN(n6582) );
  INV_X1 U8135 ( .A(n6580), .ZN(n6581) );
  XNOR2_X1 U8136 ( .A(n7877), .B(n6660), .ZN(n6583) );
  NOR2_X1 U8137 ( .A1(n7889), .A2(n8108), .ZN(n6584) );
  XNOR2_X1 U8138 ( .A(n6583), .B(n6584), .ZN(n7702) );
  INV_X1 U8139 ( .A(n6583), .ZN(n6585) );
  XNOR2_X1 U8140 ( .A(n10386), .B(n6660), .ZN(n6586) );
  NOR2_X1 U8141 ( .A1(n7976), .A2(n8108), .ZN(n6587) );
  XNOR2_X1 U8142 ( .A(n6586), .B(n6587), .ZN(n7768) );
  NAND2_X1 U8143 ( .A1(n7769), .A2(n7768), .ZN(n6590) );
  INV_X1 U8144 ( .A(n6586), .ZN(n6588) );
  NAND2_X1 U8145 ( .A1(n6588), .A2(n6587), .ZN(n6589) );
  XNOR2_X1 U8146 ( .A(n8114), .B(n6660), .ZN(n6591) );
  NOR2_X1 U8147 ( .A1(n8115), .A2(n8108), .ZN(n6592) );
  XNOR2_X1 U8148 ( .A(n6591), .B(n6592), .ZN(n7838) );
  INV_X1 U8149 ( .A(n6591), .ZN(n6593) );
  NAND2_X1 U8150 ( .A1(n6593), .A2(n6592), .ZN(n6594) );
  XNOR2_X1 U8151 ( .A(n9972), .B(n6660), .ZN(n6596) );
  NAND2_X1 U8152 ( .A1(n8929), .A2(n6612), .ZN(n6597) );
  NAND2_X1 U8153 ( .A1(n6596), .A2(n6597), .ZN(n6601) );
  INV_X1 U8154 ( .A(n6596), .ZN(n6599) );
  INV_X1 U8155 ( .A(n6597), .ZN(n6598) );
  NAND2_X1 U8156 ( .A1(n6599), .A2(n6598), .ZN(n6600) );
  NAND2_X1 U8157 ( .A1(n6601), .A2(n6600), .ZN(n7926) );
  NOR2_X1 U8158 ( .A1(n8576), .A2(n8108), .ZN(n8569) );
  XNOR2_X1 U8159 ( .A(n9016), .B(n6649), .ZN(n8567) );
  XNOR2_X1 U8160 ( .A(n9010), .B(n6660), .ZN(n6602) );
  OR2_X1 U8161 ( .A1(n8885), .A2(n8108), .ZN(n6603) );
  NAND2_X1 U8162 ( .A1(n6602), .A2(n6603), .ZN(n8572) );
  OAI21_X1 U8163 ( .B1(n8569), .B2(n8567), .A(n8572), .ZN(n6608) );
  NAND3_X1 U8164 ( .A1(n8572), .A2(n8569), .A3(n8567), .ZN(n6606) );
  INV_X1 U8165 ( .A(n6602), .ZN(n6605) );
  INV_X1 U8166 ( .A(n6603), .ZN(n6604) );
  NAND2_X1 U8167 ( .A1(n6605), .A2(n6604), .ZN(n8571) );
  AND2_X1 U8168 ( .A1(n6606), .A2(n8571), .ZN(n6607) );
  XNOR2_X1 U8169 ( .A(n9005), .B(n6660), .ZN(n6609) );
  NOR2_X1 U8170 ( .A1(n8869), .A2(n8108), .ZN(n6610) );
  XNOR2_X1 U8171 ( .A(n6609), .B(n6610), .ZN(n8023) );
  NAND2_X1 U8172 ( .A1(n8024), .A2(n8023), .ZN(n8610) );
  INV_X1 U8173 ( .A(n6609), .ZN(n6611) );
  NAND2_X1 U8174 ( .A1(n6611), .A2(n6610), .ZN(n8609) );
  NOR2_X1 U8175 ( .A1(n8887), .A2(n8108), .ZN(n6614) );
  AND2_X1 U8176 ( .A1(n8609), .A2(n6613), .ZN(n6617) );
  INV_X1 U8177 ( .A(n6613), .ZN(n6616) );
  XNOR2_X1 U8178 ( .A(n6615), .B(n6614), .ZN(n8611) );
  XNOR2_X1 U8179 ( .A(n8994), .B(n6660), .ZN(n6618) );
  NAND2_X1 U8180 ( .A1(n8867), .A2(n6612), .ZN(n6619) );
  NAND2_X1 U8181 ( .A1(n6618), .A2(n6619), .ZN(n6623) );
  INV_X1 U8182 ( .A(n6618), .ZN(n6621) );
  INV_X1 U8183 ( .A(n6619), .ZN(n6620) );
  NAND2_X1 U8184 ( .A1(n6621), .A2(n6620), .ZN(n6622) );
  NAND2_X1 U8185 ( .A1(n6623), .A2(n6622), .ZN(n8527) );
  XNOR2_X1 U8186 ( .A(n8987), .B(n6649), .ZN(n6624) );
  NOR2_X1 U8187 ( .A1(n8548), .A2(n8108), .ZN(n6625) );
  XNOR2_X1 U8188 ( .A(n6624), .B(n6625), .ZN(n8592) );
  INV_X1 U8189 ( .A(n6624), .ZN(n6627) );
  INV_X1 U8190 ( .A(n6625), .ZN(n6626) );
  XNOR2_X1 U8191 ( .A(n8823), .B(n6649), .ZN(n6628) );
  NOR2_X1 U8192 ( .A1(n8812), .A2(n8108), .ZN(n6629) );
  XNOR2_X1 U8193 ( .A(n6628), .B(n6629), .ZN(n8544) );
  NAND2_X1 U8194 ( .A1(n8545), .A2(n8544), .ZN(n6632) );
  INV_X1 U8195 ( .A(n6628), .ZN(n6630) );
  NAND2_X1 U8196 ( .A1(n6630), .A2(n6629), .ZN(n6631) );
  NAND2_X1 U8197 ( .A1(n6632), .A2(n6631), .ZN(n6635) );
  XNOR2_X1 U8198 ( .A(n8977), .B(n6660), .ZN(n6633) );
  INV_X1 U8199 ( .A(n8547), .ZN(n8826) );
  NAND2_X1 U8200 ( .A1(n8826), .A2(n6612), .ZN(n8601) );
  NAND2_X1 U8201 ( .A1(n8602), .A2(n8601), .ZN(n8600) );
  INV_X1 U8202 ( .A(n6633), .ZN(n6634) );
  INV_X1 U8203 ( .A(n6642), .ZN(n6638) );
  XNOR2_X1 U8204 ( .A(n8972), .B(n6649), .ZN(n6637) );
  INV_X1 U8205 ( .A(n6637), .ZN(n6643) );
  INV_X1 U8206 ( .A(n8584), .ZN(n6640) );
  INV_X1 U8207 ( .A(n6639), .ZN(n8583) );
  NAND2_X1 U8208 ( .A1(n6643), .A2(n6642), .ZN(n6644) );
  OR2_X1 U8209 ( .A1(n8813), .A2(n8108), .ZN(n8582) );
  NAND2_X1 U8210 ( .A1(n6646), .A2(n6645), .ZN(n6647) );
  XNOR2_X1 U8211 ( .A(n8963), .B(n6649), .ZN(n8554) );
  INV_X1 U8212 ( .A(n8554), .ZN(n6652) );
  NOR2_X1 U8213 ( .A1(n8777), .A2(n8108), .ZN(n8553) );
  AOI21_X1 U8214 ( .B1(n6650), .B2(n8554), .A(n8553), .ZN(n6651) );
  AOI21_X2 U8215 ( .B1(n8556), .B2(n6652), .A(n6651), .ZN(n8625) );
  XNOR2_X1 U8216 ( .A(n8957), .B(n6660), .ZN(n6654) );
  OR2_X1 U8217 ( .A1(n8557), .A2(n8108), .ZN(n6653) );
  AOI21_X1 U8218 ( .B1(n6654), .B2(n6653), .A(n6655), .ZN(n8624) );
  NAND2_X1 U8219 ( .A1(n8625), .A2(n8624), .ZN(n8623) );
  INV_X1 U8220 ( .A(n6655), .ZN(n6656) );
  NAND2_X2 U8221 ( .A1(n8623), .A2(n6656), .ZN(n8503) );
  XNOR2_X1 U8222 ( .A(n8951), .B(n6660), .ZN(n6658) );
  NAND2_X1 U8223 ( .A1(n8637), .A2(n6612), .ZN(n6657) );
  NOR2_X1 U8224 ( .A1(n6658), .A2(n6657), .ZN(n6659) );
  AOI21_X1 U8225 ( .B1(n6658), .B2(n6657), .A(n6659), .ZN(n8502) );
  INV_X1 U8226 ( .A(n6659), .ZN(n6688) );
  NAND2_X1 U8227 ( .A1(n8501), .A2(n6688), .ZN(n6696) );
  NOR2_X1 U8228 ( .A1(n8130), .A2(n8108), .ZN(n6661) );
  XNOR2_X1 U8229 ( .A(n6661), .B(n6660), .ZN(n6686) );
  NOR4_X1 U8230 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6670) );
  INV_X1 U8231 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10302) );
  INV_X1 U8232 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10299) );
  INV_X1 U8233 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10313) );
  INV_X1 U8234 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10321) );
  NAND4_X1 U8235 ( .A1(n10302), .A2(n10299), .A3(n10313), .A4(n10321), .ZN(
        n6667) );
  NOR4_X1 U8236 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6665) );
  NOR4_X1 U8237 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6664) );
  NOR4_X1 U8238 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n6663) );
  NOR4_X1 U8239 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6662) );
  NAND4_X1 U8240 ( .A1(n6665), .A2(n6664), .A3(n6663), .A4(n6662), .ZN(n6666)
         );
  NOR4_X1 U8241 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n6667), .A4(n6666), .ZN(n6669) );
  NOR4_X1 U8242 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6668) );
  NAND3_X1 U8243 ( .A1(n6670), .A2(n6669), .A3(n6668), .ZN(n6673) );
  XNOR2_X1 U8244 ( .A(n7805), .B(P2_B_REG_SCAN_IN), .ZN(n6671) );
  NAND2_X1 U8245 ( .A1(n7916), .A2(n6671), .ZN(n6672) );
  NAND2_X1 U8246 ( .A1(n6673), .A2(n10295), .ZN(n7095) );
  INV_X1 U8247 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6674) );
  NAND2_X1 U8248 ( .A1(n10295), .A2(n6674), .ZN(n6675) );
  INV_X1 U8249 ( .A(n6677), .ZN(n7953) );
  NAND2_X1 U8250 ( .A1(n7953), .A2(n7805), .ZN(n10327) );
  NAND2_X1 U8251 ( .A1(n6675), .A2(n10327), .ZN(n7141) );
  INV_X1 U8252 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6676) );
  NAND2_X1 U8253 ( .A1(n10295), .A2(n6676), .ZN(n6679) );
  OR2_X1 U8254 ( .A1(n6678), .A2(n6677), .ZN(n10330) );
  NAND2_X1 U8255 ( .A1(n6679), .A2(n10330), .ZN(n7193) );
  NOR2_X1 U8256 ( .A1(n7141), .A2(n7193), .ZN(n6680) );
  NAND2_X1 U8257 ( .A1(n7095), .A2(n6680), .ZN(n6700) );
  NOR2_X1 U8258 ( .A1(n6700), .A2(n10294), .ZN(n6698) );
  NOR2_X1 U8259 ( .A1(n7504), .A2(n10333), .ZN(n10272) );
  NAND2_X1 U8260 ( .A1(n6698), .A2(n10272), .ZN(n6683) );
  AND2_X1 U8261 ( .A1(n4831), .A2(n7661), .ZN(n6681) );
  NAND2_X1 U8262 ( .A1(n7504), .A2(n6681), .ZN(n10357) );
  NOR2_X2 U8263 ( .A1(n10294), .A2(n7097), .ZN(n10283) );
  NOR3_X1 U8264 ( .A1(n8492), .A2(n8618), .A3(n6686), .ZN(n6684) );
  AOI21_X1 U8265 ( .B1(n8492), .B2(n6686), .A(n6684), .ZN(n6695) );
  NAND3_X1 U8266 ( .A1(n8946), .A2(n8634), .A3(n6686), .ZN(n6685) );
  OAI21_X1 U8267 ( .B1(n8946), .B2(n6686), .A(n6685), .ZN(n6687) );
  AND2_X1 U8268 ( .A1(n8502), .A2(n6687), .ZN(n6690) );
  INV_X1 U8269 ( .A(n6687), .ZN(n6689) );
  NAND2_X1 U8270 ( .A1(n6699), .A2(n6691), .ZN(n10381) );
  INV_X1 U8271 ( .A(n7078), .ZN(n6755) );
  AND2_X1 U8272 ( .A1(n10381), .A2(n6755), .ZN(n6692) );
  NAND2_X1 U8273 ( .A1(n6698), .A2(n6692), .ZN(n8620) );
  OAI21_X1 U8274 ( .B1(n8492), .B2(n8634), .A(n8620), .ZN(n6693) );
  OAI211_X1 U8275 ( .C1(n6696), .C2(n6695), .A(n6694), .B(n6693), .ZN(n6708)
         );
  INV_X1 U8276 ( .A(n6699), .ZN(n6697) );
  AND2_X1 U8277 ( .A1(n8631), .A2(n8928), .ZN(n8539) );
  INV_X1 U8278 ( .A(n8490), .ZN(n6704) );
  AND2_X1 U8279 ( .A1(n6699), .A2(n7078), .ZN(n7094) );
  AOI21_X1 U8280 ( .B1(n6700), .B2(n7097), .A(n7094), .ZN(n6987) );
  NAND2_X1 U8281 ( .A1(n6987), .A2(n6701), .ZN(n6702) );
  OAI22_X1 U8282 ( .A1(n6704), .A2(n8628), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6703), .ZN(n6705) );
  AOI21_X1 U8283 ( .B1(n8539), .B2(n8637), .A(n6705), .ZN(n6706) );
  INV_X1 U8284 ( .A(n8631), .ZN(n8560) );
  AND2_X1 U8285 ( .A1(n6522), .A2(n7078), .ZN(n8930) );
  NAND2_X1 U8286 ( .A1(n6708), .A2(n6707), .ZN(P2_U3222) );
  INV_X1 U8287 ( .A(n6740), .ZN(n6752) );
  INV_X2 U8288 ( .A(n9479), .ZN(P1_U4006) );
  NAND2_X1 U8289 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6709), .ZN(n10329) );
  NOR2_X4 U8290 ( .A1(n6828), .A2(n10329), .ZN(P2_U3966) );
  INV_X1 U8291 ( .A(n6710), .ZN(n6711) );
  NAND2_X1 U8292 ( .A1(n6711), .A2(n7743), .ZN(n7039) );
  NAND2_X1 U8293 ( .A1(n9446), .A2(n7743), .ZN(n6712) );
  NAND2_X1 U8294 ( .A1(n7039), .A2(n6712), .ZN(n6818) );
  OR2_X1 U8295 ( .A1(n6818), .A2(n6713), .ZN(n6714) );
  NAND2_X1 U8296 ( .A1(n6714), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8297 ( .A(n6716), .ZN(n6717) );
  NAND2_X1 U8298 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6791), .ZN(n7040) );
  OAI21_X1 U8299 ( .B1(n6717), .B2(P1_STATE_REG_SCAN_IN), .A(n7040), .ZN(
        P1_U3353) );
  AND2_X1 U8300 ( .A1(n6724), .A2(P2_U3152), .ZN(n9047) );
  INV_X2 U8301 ( .A(n9047), .ZN(n9050) );
  AND2_X1 U8302 ( .A1(n6723), .A2(P2_U3152), .ZN(n8010) );
  OAI222_X1 U8303 ( .A1(n9050), .A2(n6719), .B1(n4481), .B2(n6725), .C1(n6718), 
        .C2(P2_U3152), .ZN(P2_U3357) );
  OAI222_X1 U8304 ( .A1(n9050), .A2(n6720), .B1(n4481), .B2(n6727), .C1(n6845), 
        .C2(P2_U3152), .ZN(P2_U3356) );
  OAI222_X1 U8305 ( .A1(n6933), .A2(P2_U3152), .B1(n4481), .B2(n6729), .C1(
        n8332), .C2(n9050), .ZN(P2_U3355) );
  OAI222_X1 U8306 ( .A1(n6869), .A2(P2_U3152), .B1(n4481), .B2(n6731), .C1(
        n8328), .C2(n9050), .ZN(P2_U3354) );
  OAI222_X1 U8307 ( .A1(n6722), .A2(P2_U3152), .B1(n4481), .B2(n6734), .C1(
        n6721), .C2(n9050), .ZN(P2_U3353) );
  NAND2_X1 U8308 ( .A1(n6723), .A2(P1_U3084), .ZN(n9901) );
  AND2_X1 U8309 ( .A1(n6724), .A2(P1_U3084), .ZN(n8014) );
  OAI222_X1 U8310 ( .A1(n9901), .A2(n6726), .B1(n4480), .B2(n6725), .C1(
        P1_U3084), .C2(n6808), .ZN(P1_U3352) );
  INV_X1 U8311 ( .A(n9901), .ZN(n7007) );
  INV_X1 U8312 ( .A(n7007), .ZN(n9896) );
  OAI222_X1 U8313 ( .A1(n9896), .A2(n6728), .B1(n4480), .B2(n6727), .C1(
        P1_U3084), .C2(n7044), .ZN(P1_U3351) );
  OAI222_X1 U8314 ( .A1(n9896), .A2(n6730), .B1(n4480), .B2(n6729), .C1(
        P1_U3084), .C2(n9483), .ZN(P1_U3350) );
  OAI222_X1 U8315 ( .A1(n9896), .A2(n6732), .B1(n4480), .B2(n6731), .C1(
        P1_U3084), .C2(n10032), .ZN(P1_U3349) );
  OAI222_X1 U8316 ( .A1(n9896), .A2(n6735), .B1(n4480), .B2(n6734), .C1(
        P1_U3084), .C2(n6733), .ZN(P1_U3348) );
  OAI222_X1 U8317 ( .A1(n9896), .A2(n6736), .B1(n4480), .B2(n6738), .C1(
        P1_U3084), .C2(n6806), .ZN(P1_U3347) );
  OAI222_X1 U8318 ( .A1(n6908), .A2(P2_U3152), .B1(n4481), .B2(n6738), .C1(
        n6737), .C2(n9050), .ZN(P2_U3352) );
  NAND2_X1 U8319 ( .A1(n6956), .A2(n6739), .ZN(n10201) );
  INV_X1 U8320 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6742) );
  AND2_X1 U8321 ( .A1(n6740), .A2(n7922), .ZN(n6741) );
  AOI22_X1 U8322 ( .A1(n10201), .A2(n6742), .B1(n6741), .B2(n5821), .ZN(
        P1_U3440) );
  INV_X1 U8323 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6744) );
  INV_X1 U8324 ( .A(n6743), .ZN(n6746) );
  INV_X1 U8325 ( .A(n6881), .ZN(n6872) );
  OAI222_X1 U8326 ( .A1(n9896), .A2(n6744), .B1(n4480), .B2(n6746), .C1(
        P1_U3084), .C2(n6872), .ZN(P1_U3346) );
  INV_X1 U8327 ( .A(n6968), .ZN(n6974) );
  INV_X1 U8328 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6745) );
  OAI222_X1 U8329 ( .A1(n6974), .A2(P2_U3152), .B1(n4481), .B2(n6746), .C1(
        n6745), .C2(n9050), .ZN(P2_U3351) );
  INV_X1 U8330 ( .A(n7064), .ZN(n7069) );
  INV_X1 U8331 ( .A(n6747), .ZN(n6749) );
  OAI222_X1 U8332 ( .A1(n7069), .A2(P2_U3152), .B1(n4481), .B2(n6749), .C1(
        n6748), .C2(n9050), .ZN(P2_U3350) );
  OAI222_X1 U8333 ( .A1(n9896), .A2(n6750), .B1(n4480), .B2(n6749), .C1(
        P1_U3084), .C2(n10084), .ZN(P1_U3345) );
  INV_X1 U8334 ( .A(n10201), .ZN(n10203) );
  OAI22_X1 U8335 ( .A1(n10203), .A2(P1_D_REG_1__SCAN_IN), .B1(n6752), .B2(
        n6751), .ZN(n6753) );
  INV_X1 U8336 ( .A(n6753), .ZN(P1_U3441) );
  OR2_X1 U8337 ( .A1(n6832), .A2(n7747), .ZN(n6754) );
  NAND2_X1 U8338 ( .A1(n10294), .A2(n6754), .ZN(n6757) );
  NAND2_X1 U8339 ( .A1(n6832), .A2(n6755), .ZN(n6756) );
  NAND2_X1 U8340 ( .A1(n6757), .A2(n6756), .ZN(n8705) );
  INV_X1 U8341 ( .A(n8705), .ZN(n10260) );
  NOR2_X1 U8342 ( .A1(n10260), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8343 ( .A(n6758), .ZN(n6761) );
  INV_X1 U8344 ( .A(n10102), .ZN(n6759) );
  OAI222_X1 U8345 ( .A1(n4480), .A2(n6761), .B1(n6759), .B2(P1_U3084), .C1(
        n8352), .C2(n9896), .ZN(P1_U3344) );
  INV_X1 U8346 ( .A(n7112), .ZN(n7075) );
  OAI222_X1 U8347 ( .A1(P2_U3152), .A2(n7075), .B1(n4481), .B2(n6761), .C1(
        n6760), .C2(n9050), .ZN(P2_U3349) );
  INV_X1 U8348 ( .A(n6762), .ZN(n6766) );
  AOI22_X1 U8349 ( .A1(n7236), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n9047), .ZN(n6763) );
  OAI21_X1 U8350 ( .B1(n6766), .B2(n4481), .A(n6763), .ZN(P2_U3348) );
  INV_X1 U8351 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U8352 ( .A1(n7153), .A2(P1_U4006), .ZN(n6764) );
  OAI21_X1 U8353 ( .B1(P1_U4006), .B2(n6765), .A(n6764), .ZN(P1_U3555) );
  INV_X1 U8354 ( .A(n6945), .ZN(n6939) );
  OAI222_X1 U8355 ( .A1(n4480), .A2(n6766), .B1(n6939), .B2(P1_U3084), .C1(
        n8170), .C2(n9896), .ZN(P1_U3343) );
  INV_X1 U8356 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6768) );
  NAND2_X1 U8357 ( .A1(n8032), .A2(P2_U3966), .ZN(n6767) );
  OAI21_X1 U8358 ( .B1(P2_U3966), .B2(n6768), .A(n6767), .ZN(P2_U3583) );
  INV_X1 U8359 ( .A(n6769), .ZN(n6771) );
  INV_X1 U8360 ( .A(n7506), .ZN(n7509) );
  OAI222_X1 U8361 ( .A1(n4480), .A2(n6771), .B1(n7509), .B2(P1_U3084), .C1(
        n6770), .C2(n9896), .ZN(P1_U3342) );
  INV_X1 U8362 ( .A(n7551), .ZN(n7543) );
  OAI222_X1 U8363 ( .A1(P2_U3152), .A2(n7543), .B1(n4481), .B2(n6771), .C1(
        n8312), .C2(n9050), .ZN(P2_U3347) );
  INV_X1 U8364 ( .A(n7039), .ZN(n6772) );
  NOR2_X1 U8365 ( .A1(P1_U3083), .A2(n6772), .ZN(n10041) );
  OR2_X1 U8366 ( .A1(n5853), .A2(P1_U3084), .ZN(n9459) );
  NOR2_X1 U8367 ( .A1(n6818), .A2(n9459), .ZN(n6805) );
  NAND2_X1 U8368 ( .A1(n6805), .A2(n9458), .ZN(n10131) );
  NOR3_X1 U8369 ( .A1(n10131), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n6773), .ZN(
        n6774) );
  AOI21_X1 U8370 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .A(n6774), .ZN(
        n6781) );
  NAND2_X1 U8371 ( .A1(n6791), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7034) );
  INV_X1 U8372 ( .A(n7034), .ZN(n10016) );
  OAI22_X1 U8373 ( .A1(n9458), .A2(n10016), .B1(n6791), .B2(n6775), .ZN(n6779)
         );
  NAND2_X1 U8374 ( .A1(n6805), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6776) );
  OAI211_X1 U8375 ( .C1(n7040), .C2(n6818), .A(n10131), .B(n6776), .ZN(n6778)
         );
  OAI211_X1 U8376 ( .C1(n5853), .C2(n6779), .A(n6778), .B(n6777), .ZN(n6780)
         );
  OAI211_X1 U8377 ( .C1(n10175), .C2(n10413), .A(n6781), .B(n6780), .ZN(
        P1_U3241) );
  MUX2_X1 U8378 ( .A(n6825), .B(n7899), .S(P1_U4006), .Z(n6782) );
  INV_X1 U8379 ( .A(n6782), .ZN(P1_U3567) );
  INV_X1 U8380 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6787) );
  INV_X1 U8381 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6785) );
  NAND2_X1 U8382 ( .A1(n5755), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6784) );
  INV_X1 U8383 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9538) );
  OR2_X1 U8384 ( .A1(n5806), .A2(n9538), .ZN(n6783) );
  OAI211_X1 U8385 ( .C1(n4593), .C2(n6785), .A(n6784), .B(n6783), .ZN(n9540)
         );
  NAND2_X1 U8386 ( .A1(n9540), .A2(P1_U4006), .ZN(n6786) );
  OAI21_X1 U8387 ( .B1(P1_U4006), .B2(n6787), .A(n6786), .ZN(P1_U3586) );
  NAND2_X1 U8388 ( .A1(n8649), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n6788) );
  OAI21_X1 U8389 ( .B1(n8115), .B2(n8649), .A(n6788), .ZN(P2_U3565) );
  MUX2_X1 U8390 ( .A(n6789), .B(n7816), .S(P1_U4006), .Z(n6790) );
  INV_X1 U8391 ( .A(n6790), .ZN(P1_U3565) );
  INV_X1 U8392 ( .A(n6806), .ZN(n10069) );
  NOR2_X1 U8393 ( .A1(n10069), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6802) );
  INV_X1 U8394 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6792) );
  MUX2_X1 U8395 ( .A(n6792), .B(P1_REG1_REG_1__SCAN_IN), .S(n6808), .Z(n10025)
         );
  AND2_X1 U8396 ( .A1(n6791), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10026) );
  NAND2_X1 U8397 ( .A1(n10025), .A2(n10026), .ZN(n10024) );
  OR2_X1 U8398 ( .A1(n6808), .A2(n6792), .ZN(n7045) );
  NAND2_X1 U8399 ( .A1(n10024), .A2(n7045), .ZN(n6794) );
  MUX2_X1 U8400 ( .A(n10248), .B(P1_REG1_REG_2__SCAN_IN), .S(n7044), .Z(n6793)
         );
  NAND2_X1 U8401 ( .A1(n6794), .A2(n6793), .ZN(n9485) );
  INV_X1 U8402 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10248) );
  OR2_X1 U8403 ( .A1(n7044), .A2(n10248), .ZN(n9484) );
  NAND2_X1 U8404 ( .A1(n9485), .A2(n9484), .ZN(n6796) );
  MUX2_X1 U8405 ( .A(n6797), .B(P1_REG1_REG_3__SCAN_IN), .S(n9483), .Z(n6795)
         );
  NAND2_X1 U8406 ( .A1(n6796), .A2(n6795), .ZN(n9488) );
  OR2_X1 U8407 ( .A1(n9483), .A2(n6797), .ZN(n6798) );
  AND2_X1 U8408 ( .A1(n9488), .A2(n6798), .ZN(n10037) );
  INV_X1 U8409 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10250) );
  MUX2_X1 U8410 ( .A(n10250), .B(P1_REG1_REG_4__SCAN_IN), .S(n10032), .Z(
        n10036) );
  NAND2_X1 U8411 ( .A1(n10037), .A2(n10036), .ZN(n10035) );
  NAND2_X1 U8412 ( .A1(n10032), .A2(n10250), .ZN(n6799) );
  NAND2_X1 U8413 ( .A1(n10035), .A2(n6799), .ZN(n10056) );
  MUX2_X1 U8414 ( .A(n5204), .B(P1_REG1_REG_5__SCAN_IN), .S(n10051), .Z(n10057) );
  NAND2_X1 U8415 ( .A1(n10051), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6800) );
  NAND2_X1 U8416 ( .A1(n10058), .A2(n6800), .ZN(n10075) );
  MUX2_X1 U8417 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6801), .S(n6806), .Z(n10076)
         );
  NOR2_X1 U8418 ( .A1(n10075), .A2(n10076), .ZN(n10074) );
  NOR2_X1 U8419 ( .A1(n6802), .A2(n10074), .ZN(n6804) );
  AOI22_X1 U8420 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6872), .B1(n6881), .B2(
        n5257), .ZN(n6803) );
  NOR2_X1 U8421 ( .A1(n6804), .A2(n6803), .ZN(n6871) );
  AOI21_X1 U8422 ( .B1(n6804), .B2(n6803), .A(n6871), .ZN(n6823) );
  INV_X1 U8423 ( .A(n9458), .ZN(n8098) );
  NAND2_X1 U8424 ( .A1(n6805), .A2(n8098), .ZN(n10161) );
  INV_X1 U8425 ( .A(n10161), .ZN(n10088) );
  AOI22_X1 U8426 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6881), .B1(n6872), .B2(
        n7413), .ZN(n6817) );
  XNOR2_X1 U8427 ( .A(n6806), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n10063) );
  NOR2_X1 U8428 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n10051), .ZN(n6807) );
  AOI21_X1 U8429 ( .B1(n10051), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6807), .ZN(
        n10047) );
  MUX2_X1 U8430 ( .A(n5126), .B(P1_REG2_REG_2__SCAN_IN), .S(n7044), .Z(n7043)
         );
  INV_X1 U8431 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10192) );
  MUX2_X1 U8432 ( .A(n10192), .B(P1_REG2_REG_1__SCAN_IN), .S(n6808), .Z(n10017) );
  NAND2_X1 U8433 ( .A1(n10017), .A2(n10016), .ZN(n10015) );
  INV_X1 U8434 ( .A(n6808), .ZN(n10019) );
  NAND2_X1 U8435 ( .A1(n10019), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6809) );
  NAND2_X1 U8436 ( .A1(n10015), .A2(n6809), .ZN(n7042) );
  NAND2_X1 U8437 ( .A1(n7043), .A2(n7042), .ZN(n7041) );
  INV_X1 U8438 ( .A(n7044), .ZN(n7050) );
  NAND2_X1 U8439 ( .A1(n7050), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U8440 ( .A1(n7041), .A2(n6810), .ZN(n9490) );
  MUX2_X1 U8441 ( .A(n6811), .B(P1_REG2_REG_3__SCAN_IN), .S(n9483), .Z(n9491)
         );
  NAND2_X1 U8442 ( .A1(n9490), .A2(n9491), .ZN(n9489) );
  OR2_X1 U8443 ( .A1(n9483), .A2(n6811), .ZN(n6812) );
  MUX2_X1 U8444 ( .A(n6813), .B(P1_REG2_REG_4__SCAN_IN), .S(n10032), .Z(n10030) );
  NAND2_X1 U8445 ( .A1(n10031), .A2(n10030), .ZN(n10029) );
  NAND2_X1 U8446 ( .A1(n10032), .A2(n6813), .ZN(n6814) );
  NAND2_X1 U8447 ( .A1(n10029), .A2(n6814), .ZN(n10048) );
  NAND2_X1 U8448 ( .A1(n10047), .A2(n10048), .ZN(n10046) );
  INV_X1 U8449 ( .A(n10067), .ZN(n6815) );
  NAND2_X1 U8450 ( .A1(n6817), .A2(n6816), .ZN(n6880) );
  OAI21_X1 U8451 ( .B1(n6817), .B2(n6816), .A(n6880), .ZN(n6821) );
  INV_X1 U8452 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n8193) );
  NAND2_X1 U8453 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7251) );
  OR2_X1 U8454 ( .A1(n9458), .A2(P1_U3084), .ZN(n7966) );
  OR2_X1 U8455 ( .A1(n6818), .A2(n7966), .ZN(n9533) );
  NOR2_X2 U8456 ( .A1(n9533), .A2(n7159), .ZN(n10168) );
  NAND2_X1 U8457 ( .A1(n10168), .A2(n6881), .ZN(n6819) );
  OAI211_X1 U8458 ( .C1(n10175), .C2(n8193), .A(n7251), .B(n6819), .ZN(n6820)
         );
  AOI21_X1 U8459 ( .B1(n10088), .B2(n6821), .A(n6820), .ZN(n6822) );
  OAI21_X1 U8460 ( .B1(n6823), .B2(n10131), .A(n6822), .ZN(P1_U3248) );
  INV_X1 U8461 ( .A(n7603), .ZN(n7599) );
  INV_X1 U8462 ( .A(n6824), .ZN(n6826) );
  OAI222_X1 U8463 ( .A1(n7599), .A2(P2_U3152), .B1(n4481), .B2(n6826), .C1(
        n6825), .C2(n9050), .ZN(P2_U3346) );
  INV_X1 U8464 ( .A(n10114), .ZN(n7511) );
  OAI222_X1 U8465 ( .A1(n9896), .A2(n6827), .B1(n4480), .B2(n6826), .C1(
        P1_U3084), .C2(n7511), .ZN(P1_U3341) );
  OR2_X1 U8466 ( .A1(n6522), .A2(P2_U3152), .ZN(n8011) );
  OAI21_X1 U8467 ( .B1(n8011), .B2(n6828), .A(n7747), .ZN(n6829) );
  INV_X1 U8468 ( .A(n6829), .ZN(n6830) );
  OAI21_X1 U8469 ( .B1(n10294), .B2(n7078), .A(n6830), .ZN(n6834) );
  NAND2_X1 U8470 ( .A1(n6834), .A2(n6832), .ZN(n6831) );
  NAND2_X1 U8471 ( .A1(n6831), .A2(n8649), .ZN(n6852) );
  AND2_X1 U8472 ( .A1(n6852), .A2(n6522), .ZN(n9921) );
  AND2_X1 U8473 ( .A1(n6832), .A2(n8029), .ZN(n6833) );
  INV_X1 U8474 ( .A(n10258), .ZN(n10262) );
  INV_X1 U8475 ( .A(n6869), .ZN(n6849) );
  NAND2_X1 U8476 ( .A1(n6848), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6839) );
  MUX2_X1 U8477 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6835), .S(n6848), .Z(n6929)
         );
  MUX2_X1 U8478 ( .A(n6836), .B(P2_REG1_REG_2__SCAN_IN), .S(n6845), .Z(n9923)
         );
  NAND2_X1 U8479 ( .A1(n9909), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6838) );
  MUX2_X1 U8480 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6837), .S(n9909), .Z(n9912)
         );
  NAND3_X1 U8481 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n9912), .ZN(n9911) );
  NAND2_X1 U8482 ( .A1(n6838), .A2(n9911), .ZN(n9924) );
  NAND2_X1 U8483 ( .A1(n9923), .A2(n9924), .ZN(n9922) );
  OAI21_X1 U8484 ( .B1(n6845), .B2(n6836), .A(n9922), .ZN(n6930) );
  NAND2_X1 U8485 ( .A1(n6929), .A2(n6930), .ZN(n6928) );
  AND2_X1 U8486 ( .A1(n6839), .A2(n6928), .ZN(n6860) );
  MUX2_X1 U8487 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n5970), .S(n6869), .Z(n6859)
         );
  NOR2_X1 U8488 ( .A1(n6860), .A2(n6859), .ZN(n6858) );
  AOI21_X1 U8489 ( .B1(n6849), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6858), .ZN(
        n6900) );
  MUX2_X1 U8490 ( .A(n5987), .B(P2_REG1_REG_5__SCAN_IN), .S(n6898), .Z(n6899)
         );
  XNOR2_X1 U8491 ( .A(n6900), .B(n6899), .ZN(n6842) );
  NOR2_X1 U8492 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5985), .ZN(n6840) );
  AOI21_X1 U8493 ( .B1(n10260), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6840), .ZN(
        n6841) );
  OAI21_X1 U8494 ( .B1(n10262), .B2(n6842), .A(n6841), .ZN(n6856) );
  MUX2_X1 U8495 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6843), .S(n6869), .Z(n6864)
         );
  NAND2_X1 U8496 ( .A1(n9909), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6844) );
  NAND2_X1 U8497 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9907) );
  NOR2_X1 U8498 ( .A1(n9906), .A2(n9907), .ZN(n9905) );
  AOI21_X1 U8499 ( .B1(n9909), .B2(P2_REG2_REG_1__SCAN_IN), .A(n9905), .ZN(
        n9919) );
  INV_X1 U8500 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6846) );
  NAND2_X1 U8501 ( .A1(n6848), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6847) );
  OAI21_X1 U8502 ( .B1(n6848), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6847), .ZN(
        n6926) );
  NOR2_X1 U8503 ( .A1(n4502), .A2(n6926), .ZN(n6925) );
  NAND2_X1 U8504 ( .A1(n6898), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6850) );
  OAI21_X1 U8505 ( .B1(n6898), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6850), .ZN(
        n6853) );
  NOR2_X1 U8506 ( .A1(n6522), .A2(n8029), .ZN(n6851) );
  NAND2_X1 U8507 ( .A1(n6852), .A2(n6851), .ZN(n10263) );
  AOI211_X1 U8508 ( .C1(n6854), .C2(n6853), .A(n6893), .B(n10263), .ZN(n6855)
         );
  AOI211_X1 U8509 ( .C1(n9921), .C2(n6898), .A(n6856), .B(n6855), .ZN(n6857)
         );
  INV_X1 U8510 ( .A(n6857), .ZN(P2_U3250) );
  AND2_X1 U8511 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6862) );
  AOI211_X1 U8512 ( .C1(n6860), .C2(n6859), .A(n6858), .B(n10262), .ZN(n6861)
         );
  AOI211_X1 U8513 ( .C1(n10260), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6862), .B(
        n6861), .ZN(n6868) );
  AOI211_X1 U8514 ( .C1(n6865), .C2(n6864), .A(n6863), .B(n10263), .ZN(n6866)
         );
  INV_X1 U8515 ( .A(n6866), .ZN(n6867) );
  OAI211_X1 U8516 ( .C1(n10261), .C2(n6869), .A(n6868), .B(n6867), .ZN(
        P2_U3249) );
  NAND2_X1 U8517 ( .A1(n8649), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6870) );
  OAI21_X1 U8518 ( .B1(n8813), .B2(n8649), .A(n6870), .ZN(P2_U3575) );
  NOR2_X1 U8519 ( .A1(n10102), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6875) );
  AOI21_X1 U8520 ( .B1(n5257), .B2(n6872), .A(n6871), .ZN(n10092) );
  MUX2_X1 U8521 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6873), .S(n10084), .Z(n10091) );
  NOR2_X1 U8522 ( .A1(n10092), .A2(n10091), .ZN(n10090) );
  AOI21_X1 U8523 ( .B1(n6873), .B2(n10084), .A(n10090), .ZN(n10105) );
  MUX2_X1 U8524 ( .A(n6874), .B(P1_REG1_REG_9__SCAN_IN), .S(n10102), .Z(n10104) );
  NOR2_X1 U8525 ( .A1(n10105), .A2(n10104), .ZN(n10103) );
  NOR2_X1 U8526 ( .A1(n6875), .A2(n10103), .ZN(n6878) );
  MUX2_X1 U8527 ( .A(n6876), .B(P1_REG1_REG_10__SCAN_IN), .S(n6945), .Z(n6877)
         );
  NOR2_X1 U8528 ( .A1(n6878), .A2(n6877), .ZN(n6938) );
  AOI21_X1 U8529 ( .B1(n6878), .B2(n6877), .A(n6938), .ZN(n6891) );
  NAND2_X1 U8530 ( .A1(n10102), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6879) );
  OAI21_X1 U8531 ( .B1(n10102), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6879), .ZN(
        n10098) );
  OAI21_X1 U8532 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6881), .A(n6880), .ZN(
        n10083) );
  MUX2_X1 U8533 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n7626), .S(n10084), .Z(n6882)
         );
  INV_X1 U8534 ( .A(n6882), .ZN(n10082) );
  NAND2_X1 U8535 ( .A1(n10083), .A2(n10082), .ZN(n10081) );
  NOR2_X1 U8536 ( .A1(n10098), .A2(n10099), .ZN(n10097) );
  AOI22_X1 U8537 ( .A1(n6945), .A2(n5351), .B1(P1_REG2_REG_10__SCAN_IN), .B2(
        n6939), .ZN(n6884) );
  NOR2_X1 U8538 ( .A1(n6885), .A2(n6884), .ZN(n6944) );
  AOI211_X1 U8539 ( .C1(n6885), .C2(n6884), .A(n6944), .B(n10161), .ZN(n6886)
         );
  INV_X1 U8540 ( .A(n6886), .ZN(n6890) );
  NOR2_X1 U8541 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6887), .ZN(n7537) );
  INV_X1 U8542 ( .A(n10168), .ZN(n10085) );
  NOR2_X1 U8543 ( .A1(n10085), .A2(n6939), .ZN(n6888) );
  AOI211_X1 U8544 ( .C1(n10041), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n7537), .B(
        n6888), .ZN(n6889) );
  OAI211_X1 U8545 ( .C1(n6891), .C2(n10131), .A(n6890), .B(n6889), .ZN(
        P1_U3251) );
  INV_X1 U8546 ( .A(n6892), .ZN(n6937) );
  INV_X1 U8547 ( .A(n10127), .ZN(n7512) );
  OAI222_X1 U8548 ( .A1(n4480), .A2(n6937), .B1(n7512), .B2(P1_U3084), .C1(
        n8288), .C2(n9896), .ZN(P1_U3340) );
  MUX2_X1 U8549 ( .A(n6894), .B(P2_REG2_REG_6__SCAN_IN), .S(n6915), .Z(n6895)
         );
  AOI211_X1 U8550 ( .C1(n6896), .C2(n6895), .A(n6911), .B(n10263), .ZN(n6910)
         );
  NOR2_X1 U8551 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6897), .ZN(n7376) );
  AOI21_X1 U8552 ( .B1(n10260), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7376), .ZN(
        n6907) );
  NAND2_X1 U8553 ( .A1(n6898), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6902) );
  OR2_X1 U8554 ( .A1(n6900), .A2(n6899), .ZN(n6901) );
  NAND2_X1 U8555 ( .A1(n6902), .A2(n6901), .ZN(n6905) );
  MUX2_X1 U8556 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6903), .S(n6915), .Z(n6904)
         );
  NAND2_X1 U8557 ( .A1(n6904), .A2(n6905), .ZN(n6916) );
  OAI211_X1 U8558 ( .C1(n6905), .C2(n6904), .A(n10258), .B(n6916), .ZN(n6906)
         );
  OAI211_X1 U8559 ( .C1(n10261), .C2(n6908), .A(n6907), .B(n6906), .ZN(n6909)
         );
  OR2_X1 U8560 ( .A1(n6910), .A2(n6909), .ZN(P2_U3251) );
  MUX2_X1 U8561 ( .A(n6912), .B(P2_REG2_REG_7__SCAN_IN), .S(n6968), .Z(n6913)
         );
  NOR2_X1 U8562 ( .A1(n4500), .A2(n6913), .ZN(n6967) );
  AOI211_X1 U8563 ( .C1(n4500), .C2(n6913), .A(n6967), .B(n10263), .ZN(n6924)
         );
  NOR2_X1 U8564 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6009), .ZN(n6914) );
  AOI21_X1 U8565 ( .B1(n10260), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6914), .ZN(
        n6922) );
  NAND2_X1 U8566 ( .A1(n6915), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6917) );
  NAND2_X1 U8567 ( .A1(n6917), .A2(n6916), .ZN(n6920) );
  MUX2_X1 U8568 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6918), .S(n6968), .Z(n6919)
         );
  NAND2_X1 U8569 ( .A1(n6919), .A2(n6920), .ZN(n6973) );
  OAI211_X1 U8570 ( .C1(n6920), .C2(n6919), .A(n10258), .B(n6973), .ZN(n6921)
         );
  OAI211_X1 U8571 ( .C1(n10261), .C2(n6974), .A(n6922), .B(n6921), .ZN(n6923)
         );
  OR2_X1 U8572 ( .A1(n6924), .A2(n6923), .ZN(P2_U3252) );
  AOI211_X1 U8573 ( .C1(n4502), .C2(n6926), .A(n6925), .B(n10263), .ZN(n6935)
         );
  INV_X1 U8574 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10282) );
  NOR2_X1 U8575 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10282), .ZN(n6927) );
  AOI21_X1 U8576 ( .B1(n10260), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6927), .ZN(
        n6932) );
  OAI211_X1 U8577 ( .C1(n6930), .C2(n6929), .A(n10258), .B(n6928), .ZN(n6931)
         );
  OAI211_X1 U8578 ( .C1(n10261), .C2(n6933), .A(n6932), .B(n6931), .ZN(n6934)
         );
  OR2_X1 U8579 ( .A1(n6935), .A2(n6934), .ZN(P2_U3248) );
  INV_X1 U8580 ( .A(n7734), .ZN(n7729) );
  OAI222_X1 U8581 ( .A1(P2_U3152), .A2(n7729), .B1(n4481), .B2(n6937), .C1(
        n6936), .C2(n9050), .ZN(P2_U3345) );
  AOI21_X1 U8582 ( .B1(n6939), .B2(n6876), .A(n6938), .ZN(n6941) );
  INV_X1 U8583 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10009) );
  AOI22_X1 U8584 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n7509), .B1(n7506), .B2(
        n10009), .ZN(n6940) );
  NOR2_X1 U8585 ( .A1(n6941), .A2(n6940), .ZN(n7508) );
  AOI21_X1 U8586 ( .B1(n6941), .B2(n6940), .A(n7508), .ZN(n6951) );
  NOR2_X1 U8587 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5376), .ZN(n7651) );
  NOR2_X1 U8588 ( .A1(n10085), .A2(n7509), .ZN(n6942) );
  AOI211_X1 U8589 ( .C1(n10041), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n7651), .B(
        n6942), .ZN(n6950) );
  NOR2_X1 U8590 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7506), .ZN(n6943) );
  AOI21_X1 U8591 ( .B1(n7506), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6943), .ZN(
        n6947) );
  AOI21_X1 U8592 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n6945), .A(n6944), .ZN(
        n6946) );
  NAND2_X1 U8593 ( .A1(n6947), .A2(n6946), .ZN(n7505) );
  OAI21_X1 U8594 ( .B1(n6947), .B2(n6946), .A(n7505), .ZN(n6948) );
  NAND2_X1 U8595 ( .A1(n6948), .A2(n10088), .ZN(n6949) );
  OAI211_X1 U8596 ( .C1(n6951), .C2(n10131), .A(n6950), .B(n6949), .ZN(
        P1_U3252) );
  INV_X1 U8597 ( .A(n6952), .ZN(n6955) );
  INV_X1 U8598 ( .A(n7518), .ZN(n9505) );
  OAI222_X1 U8599 ( .A1(n4480), .A2(n6955), .B1(n9505), .B2(P1_U3084), .C1(
        n6953), .C2(n9896), .ZN(P1_U3339) );
  INV_X1 U8600 ( .A(n7866), .ZN(n7873) );
  OAI222_X1 U8601 ( .A1(P2_U3152), .A2(n7873), .B1(n4481), .B2(n6955), .C1(
        n6954), .C2(n9050), .ZN(P2_U3344) );
  NAND2_X1 U8602 ( .A1(n6957), .A2(n6956), .ZN(n6992) );
  INV_X1 U8603 ( .A(n6992), .ZN(n6959) );
  OAI211_X1 U8604 ( .C1(n6960), .C2(n9994), .A(n6959), .B(n6958), .ZN(n8040)
         );
  INV_X1 U8605 ( .A(n8040), .ZN(n6966) );
  XOR2_X1 U8606 ( .A(n6962), .B(n6961), .Z(n7035) );
  NAND2_X1 U8607 ( .A1(n7035), .A2(n9152), .ZN(n6964) );
  AOI22_X1 U8608 ( .A1(n9165), .A2(n7165), .B1(n10469), .B2(n9480), .ZN(n6963)
         );
  OAI211_X1 U8609 ( .C1(n6966), .C2(n6965), .A(n6964), .B(n6963), .ZN(P1_U3230) );
  MUX2_X1 U8610 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7578), .S(n7064), .Z(n6969)
         );
  INV_X1 U8611 ( .A(n6969), .ZN(n6970) );
  AOI211_X1 U8612 ( .C1(n6971), .C2(n6970), .A(n7063), .B(n10263), .ZN(n6981)
         );
  NAND2_X1 U8613 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7447) );
  INV_X1 U8614 ( .A(n7447), .ZN(n6972) );
  AOI21_X1 U8615 ( .B1(n10260), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6972), .ZN(
        n6979) );
  OAI21_X1 U8616 ( .B1(n6974), .B2(n6918), .A(n6973), .ZN(n6977) );
  MUX2_X1 U8617 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6975), .S(n7064), .Z(n6976)
         );
  NAND2_X1 U8618 ( .A1(n6976), .A2(n6977), .ZN(n7068) );
  OAI211_X1 U8619 ( .C1(n6977), .C2(n6976), .A(n10258), .B(n7068), .ZN(n6978)
         );
  OAI211_X1 U8620 ( .C1(n10261), .C2(n7069), .A(n6979), .B(n6978), .ZN(n6980)
         );
  OR2_X1 U8621 ( .A1(n6981), .A2(n6980), .ZN(P2_U3253) );
  AND2_X1 U8622 ( .A1(n8533), .A2(n6982), .ZN(n6985) );
  INV_X1 U8623 ( .A(n8620), .ZN(n8622) );
  OAI211_X1 U8624 ( .C1(n6985), .C2(n6984), .A(n6983), .B(n8622), .ZN(n6990)
         );
  AOI22_X1 U8625 ( .A1(n5941), .A2(n8928), .B1(n8930), .B2(n8647), .ZN(n7091)
         );
  INV_X1 U8626 ( .A(n7091), .ZN(n6988) );
  INV_X1 U8627 ( .A(n10294), .ZN(n6986) );
  NAND2_X1 U8628 ( .A1(n6987), .A2(n6986), .ZN(n8537) );
  AOI22_X1 U8629 ( .A1(n6988), .A2(n8631), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n8537), .ZN(n6989) );
  OAI211_X1 U8630 ( .C1(n7125), .C2(n8634), .A(n6990), .B(n6989), .ZN(P2_U3239) );
  NOR2_X1 U8631 ( .A1(n6992), .A2(n6991), .ZN(n7151) );
  INV_X1 U8632 ( .A(n7147), .ZN(n6993) );
  AND2_X1 U8633 ( .A1(n7151), .A2(n6993), .ZN(n7310) );
  AND2_X1 U8634 ( .A1(n7149), .A2(n7146), .ZN(n6994) );
  INV_X2 U8635 ( .A(n10245), .ZN(n10247) );
  INV_X1 U8636 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6999) );
  INV_X1 U8637 ( .A(n7165), .ZN(n7314) );
  INV_X1 U8638 ( .A(n7164), .ZN(n7311) );
  AND2_X1 U8639 ( .A1(n7153), .A2(n7314), .ZN(n9210) );
  NOR2_X1 U8640 ( .A1(n7157), .A2(n9210), .ZN(n9260) );
  INV_X1 U8641 ( .A(n7360), .ZN(n6995) );
  NAND2_X1 U8642 ( .A1(n6995), .A2(n7311), .ZN(n6996) );
  INV_X1 U8643 ( .A(n9935), .ZN(n9769) );
  OAI22_X1 U8644 ( .A1(n9260), .A2(n6996), .B1(n4672), .B2(n9769), .ZN(n7308)
         );
  INV_X1 U8645 ( .A(n7308), .ZN(n6997) );
  OAI21_X1 U8646 ( .B1(n7314), .B2(n7311), .A(n6997), .ZN(n9875) );
  NAND2_X1 U8647 ( .A1(n9875), .A2(n10247), .ZN(n6998) );
  OAI21_X1 U8648 ( .B1(n10247), .B2(n6999), .A(n6998), .ZN(P1_U3454) );
  XOR2_X1 U8649 ( .A(n7001), .B(n7000), .Z(n7004) );
  AOI22_X1 U8650 ( .A1(n9165), .A2(n7210), .B1(n9134), .B2(n9480), .ZN(n7003)
         );
  AOI22_X1 U8651 ( .A1(n10469), .A2(n9477), .B1(n8040), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7002) );
  OAI211_X1 U8652 ( .C1(n7004), .C2(n9139), .A(n7003), .B(n7002), .ZN(P1_U3235) );
  NAND2_X1 U8653 ( .A1(n8649), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7005) );
  OAI21_X1 U8654 ( .B1(n8777), .B2(n8649), .A(n7005), .ZN(P2_U3577) );
  INV_X1 U8655 ( .A(n7006), .ZN(n7031) );
  AOI22_X1 U8656 ( .A1(n10153), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n7007), .ZN(n7008) );
  OAI21_X1 U8657 ( .B1(n7031), .B2(n4480), .A(n7008), .ZN(P1_U3337) );
  XNOR2_X1 U8658 ( .A(n7009), .B(n7010), .ZN(n7011) );
  NAND2_X1 U8659 ( .A1(n7011), .A2(n9152), .ZN(n7015) );
  NAND2_X1 U8660 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9481) );
  INV_X1 U8661 ( .A(n9481), .ZN(n7013) );
  INV_X1 U8662 ( .A(n10469), .ZN(n9117) );
  INV_X1 U8663 ( .A(n9476), .ZN(n7335) );
  OAI22_X1 U8664 ( .A1(n9117), .A2(n7335), .B1(n7211), .B2(n9161), .ZN(n7012)
         );
  AOI211_X1 U8665 ( .C1(n7356), .C2(n9165), .A(n7013), .B(n7012), .ZN(n7014)
         );
  OAI211_X1 U8666 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9158), .A(n7015), .B(
        n7014), .ZN(P1_U3216) );
  INV_X1 U8667 ( .A(n7993), .ZN(n8001) );
  INV_X1 U8668 ( .A(n7016), .ZN(n7018) );
  OAI222_X1 U8669 ( .A1(n8001), .A2(P2_U3152), .B1(n4481), .B2(n7018), .C1(
        n7017), .C2(n9050), .ZN(P2_U3343) );
  INV_X1 U8670 ( .A(n10141), .ZN(n9510) );
  OAI222_X1 U8671 ( .A1(n9896), .A2(n7019), .B1(n4480), .B2(n7018), .C1(
        P1_U3084), .C2(n9510), .ZN(P1_U3338) );
  NAND2_X1 U8672 ( .A1(n8518), .A2(n7020), .ZN(n7022) );
  NAND2_X1 U8673 ( .A1(n7022), .A2(n7021), .ZN(n7023) );
  AOI21_X1 U8674 ( .B1(n7024), .B2(n7023), .A(n8620), .ZN(n7030) );
  NAND2_X1 U8675 ( .A1(n8645), .A2(n8930), .ZN(n7026) );
  NAND2_X1 U8676 ( .A1(n8647), .A2(n8928), .ZN(n7025) );
  NAND2_X1 U8677 ( .A1(n7026), .A2(n7025), .ZN(n7183) );
  AOI22_X1 U8678 ( .A1(n7183), .A2(n8631), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n7028) );
  OR2_X1 U8679 ( .A1(n8628), .A2(n7260), .ZN(n7027) );
  OAI211_X1 U8680 ( .C1(n7282), .C2(n8634), .A(n7028), .B(n7027), .ZN(n7029)
         );
  OR2_X1 U8681 ( .A1(n7030), .A2(n7029), .ZN(P2_U3232) );
  INV_X1 U8682 ( .A(n8652), .ZN(n8658) );
  OAI222_X1 U8683 ( .A1(n9050), .A2(n7032), .B1(n4481), .B2(n7031), .C1(
        P2_U3152), .C2(n8658), .ZN(P2_U3342) );
  INV_X1 U8684 ( .A(n7040), .ZN(n7033) );
  OAI22_X1 U8685 ( .A1(n5853), .A2(n7034), .B1(P1_REG2_REG_0__SCAN_IN), .B2(
        n7033), .ZN(n7037) );
  NOR2_X1 U8686 ( .A1(n7035), .A2(n5853), .ZN(n7036) );
  MUX2_X1 U8687 ( .A(n7037), .B(n7036), .S(n9458), .Z(n7038) );
  AOI211_X1 U8688 ( .C1(n7040), .C2(n9459), .A(n7039), .B(n7038), .ZN(n10042)
         );
  AND2_X1 U8689 ( .A1(n10041), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n7054) );
  OAI21_X1 U8690 ( .B1(n7043), .B2(n7042), .A(n7041), .ZN(n7049) );
  MUX2_X1 U8691 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10248), .S(n7044), .Z(n7046)
         );
  NAND3_X1 U8692 ( .A1(n7046), .A2(n10024), .A3(n7045), .ZN(n7047) );
  NAND2_X1 U8693 ( .A1(n9485), .A2(n7047), .ZN(n7048) );
  OAI22_X1 U8694 ( .A1(n10161), .A2(n7049), .B1(n10131), .B2(n7048), .ZN(n7053) );
  INV_X1 U8695 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7394) );
  NAND2_X1 U8696 ( .A1(n10168), .A2(n7050), .ZN(n7051) );
  OAI21_X1 U8697 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7394), .A(n7051), .ZN(n7052) );
  OR4_X1 U8698 ( .A1(n10042), .A2(n7054), .A3(n7053), .A4(n7052), .ZN(P1_U3243) );
  AOI21_X1 U8699 ( .B1(n7055), .B2(n7056), .A(n9139), .ZN(n7058) );
  NAND2_X1 U8700 ( .A1(n7058), .A2(n7057), .ZN(n7062) );
  AND2_X1 U8701 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10040) );
  INV_X1 U8702 ( .A(n9475), .ZN(n7436) );
  INV_X1 U8703 ( .A(n9477), .ZN(n7059) );
  OAI22_X1 U8704 ( .A1(n9117), .A2(n7436), .B1(n7059), .B2(n9161), .ZN(n7060)
         );
  AOI211_X1 U8705 ( .C1(n7476), .C2(n9165), .A(n10040), .B(n7060), .ZN(n7061)
         );
  OAI211_X1 U8706 ( .C1(n9158), .C2(n7474), .A(n7062), .B(n7061), .ZN(P1_U3228) );
  NAND2_X1 U8707 ( .A1(n7112), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7119) );
  OAI21_X1 U8708 ( .B1(n7112), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7119), .ZN(
        n7065) );
  AOI211_X1 U8709 ( .C1(n7066), .C2(n7065), .A(n7117), .B(n10263), .ZN(n7077)
         );
  NAND2_X1 U8710 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7589) );
  INV_X1 U8711 ( .A(n7589), .ZN(n7067) );
  AOI21_X1 U8712 ( .B1(n10260), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7067), .ZN(
        n7074) );
  OAI21_X1 U8713 ( .B1(n7069), .B2(n6975), .A(n7068), .ZN(n7072) );
  MUX2_X1 U8714 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7070), .S(n7112), .Z(n7071)
         );
  NAND2_X1 U8715 ( .A1(n7071), .A2(n7072), .ZN(n7110) );
  OAI211_X1 U8716 ( .C1(n7072), .C2(n7071), .A(n10258), .B(n7110), .ZN(n7073)
         );
  OAI211_X1 U8717 ( .C1(n10261), .C2(n7075), .A(n7074), .B(n7073), .ZN(n7076)
         );
  OR2_X1 U8718 ( .A1(n7077), .A2(n7076), .ZN(P2_U3254) );
  AOI21_X1 U8719 ( .B1(n7504), .B2(n7078), .A(n4831), .ZN(n7080) );
  NAND2_X1 U8720 ( .A1(n7197), .A2(n7661), .ZN(n7079) );
  NAND2_X1 U8721 ( .A1(n7080), .A2(n7079), .ZN(n8845) );
  NAND2_X1 U8722 ( .A1(n8845), .A2(n10357), .ZN(n10391) );
  NAND2_X1 U8723 ( .A1(n7081), .A2(n7300), .ZN(n7299) );
  NAND2_X1 U8724 ( .A1(n6530), .A2(n10338), .ZN(n7082) );
  NAND2_X1 U8725 ( .A1(n7299), .A2(n7082), .ZN(n7083) );
  NAND2_X1 U8726 ( .A1(n7083), .A2(n7088), .ZN(n7127) );
  OAI21_X1 U8727 ( .B1(n7083), .B2(n7088), .A(n7127), .ZN(n7192) );
  NOR2_X1 U8728 ( .A1(n7302), .A2(n7204), .ZN(n7133) );
  INV_X1 U8729 ( .A(n7133), .ZN(n7135) );
  AOI21_X1 U8730 ( .B1(n7302), .B2(n7204), .A(n4832), .ZN(n7084) );
  NAND2_X1 U8731 ( .A1(n7135), .A2(n7084), .ZN(n7202) );
  OAI21_X1 U8732 ( .B1(n7125), .B2(n10381), .A(n7202), .ZN(n7093) );
  INV_X1 U8733 ( .A(n7085), .ZN(n7086) );
  AOI21_X1 U8734 ( .B1(n7088), .B2(n7087), .A(n7086), .ZN(n7092) );
  NAND2_X1 U8735 ( .A1(n7090), .A2(n7089), .ZN(n8933) );
  INV_X1 U8736 ( .A(n8933), .ZN(n9966) );
  OAI21_X1 U8737 ( .B1(n7092), .B2(n9966), .A(n7091), .ZN(n7198) );
  AOI211_X1 U8738 ( .C1(n10391), .C2(n7192), .A(n7093), .B(n7198), .ZN(n7172)
         );
  NOR2_X1 U8739 ( .A1(n10294), .A2(n7094), .ZN(n7096) );
  NAND2_X1 U8740 ( .A1(n7193), .A2(n7097), .ZN(n7142) );
  NOR2_X1 U8741 ( .A1(n7142), .A2(n7141), .ZN(n7098) );
  NAND2_X1 U8742 ( .A1(n7196), .A2(n7098), .ZN(n10404) );
  NAND2_X1 U8743 ( .A1(n10404), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7099) );
  OAI21_X1 U8744 ( .B1(n7172), .B2(n10404), .A(n7099), .ZN(P2_U3522) );
  OAI211_X1 U8745 ( .C1(n7102), .C2(n7101), .A(n7100), .B(n8622), .ZN(n7107)
         );
  INV_X1 U8746 ( .A(n7103), .ZN(n10273) );
  INV_X1 U8747 ( .A(n8628), .ZN(n8505) );
  OAI22_X1 U8748 ( .A1(n8634), .A2(n7283), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5985), .ZN(n7105) );
  INV_X1 U8749 ( .A(n8539), .ZN(n8615) );
  OAI22_X1 U8750 ( .A1(n8615), .A2(n7460), .B1(n6559), .B2(n8614), .ZN(n7104)
         );
  AOI211_X1 U8751 ( .C1(n10273), .C2(n8505), .A(n7105), .B(n7104), .ZN(n7106)
         );
  NAND2_X1 U8752 ( .A1(n7107), .A2(n7106), .ZN(P2_U3229) );
  INV_X1 U8753 ( .A(n7108), .ZN(n7140) );
  INV_X1 U8754 ( .A(n10167), .ZN(n9502) );
  OAI222_X1 U8755 ( .A1(n4480), .A2(n7140), .B1(n9502), .B2(P1_U3084), .C1(
        n7109), .C2(n9896), .ZN(P1_U3336) );
  INV_X1 U8756 ( .A(n7236), .ZN(n7124) );
  NAND2_X1 U8757 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7666) );
  INV_X1 U8758 ( .A(n7666), .ZN(n7116) );
  INV_X1 U8759 ( .A(n7110), .ZN(n7111) );
  AOI21_X1 U8760 ( .B1(n7112), .B2(P2_REG1_REG_9__SCAN_IN), .A(n7111), .ZN(
        n7114) );
  MUX2_X1 U8761 ( .A(n6058), .B(P2_REG1_REG_10__SCAN_IN), .S(n7236), .Z(n7113)
         );
  NOR2_X1 U8762 ( .A1(n7113), .A2(n7114), .ZN(n7230) );
  AOI211_X1 U8763 ( .C1(n7114), .C2(n7113), .A(n7230), .B(n10262), .ZN(n7115)
         );
  AOI211_X1 U8764 ( .C1(n10260), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7116), .B(
        n7115), .ZN(n7123) );
  XNOR2_X1 U8765 ( .A(n7236), .B(n7719), .ZN(n7121) );
  INV_X1 U8766 ( .A(n10263), .ZN(n10259) );
  OAI211_X1 U8767 ( .C1(n7121), .C2(n7120), .A(n10259), .B(n7238), .ZN(n7122)
         );
  OAI211_X1 U8768 ( .C1(n10261), .C2(n7124), .A(n7123), .B(n7122), .ZN(
        P2_U3255) );
  INV_X2 U8769 ( .A(n10404), .ZN(n10406) );
  NAND2_X1 U8770 ( .A1(n7298), .A2(n7125), .ZN(n7126) );
  NAND2_X1 U8771 ( .A1(n7127), .A2(n7126), .ZN(n7129) );
  NAND2_X1 U8772 ( .A1(n7129), .A2(n7128), .ZN(n7177) );
  OAI21_X1 U8773 ( .B1(n7129), .B2(n7128), .A(n7177), .ZN(n10289) );
  INV_X1 U8774 ( .A(n10289), .ZN(n7137) );
  XNOR2_X1 U8775 ( .A(n7131), .B(n7130), .ZN(n7132) );
  OAI22_X1 U8776 ( .A1(n7460), .A2(n8886), .B1(n7298), .B2(n8884), .ZN(n8521)
         );
  AOI21_X1 U8777 ( .B1(n7132), .B2(n8933), .A(n8521), .ZN(n10292) );
  INV_X1 U8778 ( .A(n10381), .ZN(n10385) );
  NAND2_X1 U8779 ( .A1(n7133), .A2(n7174), .ZN(n7185) );
  INV_X1 U8780 ( .A(n7185), .ZN(n7134) );
  AOI211_X1 U8781 ( .C1(n10285), .C2(n7135), .A(n4832), .B(n7134), .ZN(n10286)
         );
  AOI21_X1 U8782 ( .B1(n10385), .B2(n10285), .A(n10286), .ZN(n7136) );
  OAI211_X1 U8783 ( .C1(n7137), .C2(n9020), .A(n10292), .B(n7136), .ZN(n7144)
         );
  NAND2_X1 U8784 ( .A1(n7144), .A2(n10406), .ZN(n7138) );
  OAI21_X1 U8785 ( .B1(n10406), .B2(n6835), .A(n7138), .ZN(P2_U3523) );
  INV_X1 U8786 ( .A(n8678), .ZN(n8668) );
  OAI222_X1 U8787 ( .A1(P2_U3152), .A2(n8668), .B1(n4481), .B2(n7140), .C1(
        n7139), .C2(n9050), .ZN(P2_U3341) );
  INV_X1 U8788 ( .A(n7141), .ZN(n7194) );
  NOR2_X1 U8789 ( .A1(n7194), .A2(n7142), .ZN(n7143) );
  AND2_X2 U8790 ( .A1(n7196), .A2(n7143), .ZN(n10395) );
  NAND2_X1 U8791 ( .A1(n7144), .A2(n10395), .ZN(n7145) );
  OAI21_X1 U8792 ( .B1(n10395), .B2(n5955), .A(n7145), .ZN(P2_U3460) );
  AND2_X1 U8793 ( .A1(n7147), .A2(n7146), .ZN(n7148) );
  AND2_X1 U8794 ( .A1(n7149), .A2(n7148), .ZN(n7150) );
  AND2_X1 U8795 ( .A1(n7153), .A2(n7165), .ZN(n7154) );
  OAI21_X1 U8796 ( .B1(n9261), .B2(n7154), .A(n7209), .ZN(n10179) );
  NAND2_X1 U8797 ( .A1(n10180), .A2(n9462), .ZN(n7156) );
  NAND2_X1 U8798 ( .A1(n9453), .A2(n9456), .ZN(n7155) );
  NAND2_X1 U8799 ( .A1(n7156), .A2(n7155), .ZN(n9772) );
  OAI21_X1 U8800 ( .B1(n7158), .B2(n7157), .A(n7216), .ZN(n7163) );
  INV_X1 U8801 ( .A(n7153), .ZN(n7160) );
  INV_X1 U8802 ( .A(n9938), .ZN(n9751) );
  OAI22_X1 U8803 ( .A1(n7160), .A2(n9751), .B1(n7211), .B2(n9769), .ZN(n7162)
         );
  OR3_X1 U8804 ( .A1(n7361), .A2(n7360), .A3(n10180), .ZN(n9757) );
  NOR2_X1 U8805 ( .A1(n10179), .A2(n9757), .ZN(n7161) );
  AOI211_X1 U8806 ( .C1(n9772), .C2(n7163), .A(n7162), .B(n7161), .ZN(n10177)
         );
  OR2_X1 U8807 ( .A1(n7314), .A2(n10185), .ZN(n7166) );
  AND2_X1 U8808 ( .A1(n7164), .A2(n7467), .ZN(n9950) );
  AND3_X1 U8809 ( .A1(n7166), .A2(n9950), .A3(n7395), .ZN(n10182) );
  AOI21_X1 U8810 ( .B1(n9994), .B2(n8039), .A(n10182), .ZN(n7167) );
  OAI211_X1 U8811 ( .C1(n9868), .C2(n10179), .A(n10177), .B(n7167), .ZN(n7169)
         );
  NAND2_X1 U8812 ( .A1(n7169), .A2(n10255), .ZN(n7168) );
  OAI21_X1 U8813 ( .B1(n10255), .B2(n6792), .A(n7168), .ZN(P1_U3524) );
  INV_X1 U8814 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7171) );
  NAND2_X1 U8815 ( .A1(n7169), .A2(n10247), .ZN(n7170) );
  OAI21_X1 U8816 ( .B1(n10247), .B2(n7171), .A(n7170), .ZN(P1_U3457) );
  OR2_X1 U8817 ( .A1(n7172), .A2(n10393), .ZN(n7173) );
  OAI21_X1 U8818 ( .B1(n10395), .B2(n5942), .A(n7173), .ZN(P2_U3457) );
  NAND2_X1 U8819 ( .A1(n7175), .A2(n7174), .ZN(n7176) );
  NAND2_X1 U8820 ( .A1(n7177), .A2(n7176), .ZN(n7179) );
  OAI21_X1 U8821 ( .B1(n7179), .B2(n7178), .A(n7288), .ZN(n7180) );
  INV_X1 U8822 ( .A(n7180), .ZN(n7266) );
  XNOR2_X1 U8823 ( .A(n7182), .B(n7181), .ZN(n7184) );
  AOI21_X1 U8824 ( .B1(n7184), .B2(n8933), .A(n7183), .ZN(n7269) );
  AOI21_X1 U8825 ( .B1(n7185), .B2(n7262), .A(n4832), .ZN(n7186) );
  AND2_X1 U8826 ( .A1(n7186), .A2(n7454), .ZN(n7263) );
  AOI21_X1 U8827 ( .B1(n10385), .B2(n7262), .A(n7263), .ZN(n7187) );
  OAI211_X1 U8828 ( .C1(n7266), .C2(n9020), .A(n7269), .B(n7187), .ZN(n7189)
         );
  NAND2_X1 U8829 ( .A1(n7189), .A2(n10406), .ZN(n7188) );
  OAI21_X1 U8830 ( .B1(n10406), .B2(n5970), .A(n7188), .ZN(P2_U3524) );
  INV_X1 U8831 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7191) );
  NAND2_X1 U8832 ( .A1(n7189), .A2(n10395), .ZN(n7190) );
  OAI21_X1 U8833 ( .B1(n10395), .B2(n7191), .A(n7190), .ZN(P2_U3463) );
  INV_X1 U8834 ( .A(n7192), .ZN(n7207) );
  NOR2_X1 U8835 ( .A1(n7194), .A2(n7193), .ZN(n7195) );
  NAND2_X1 U8836 ( .A1(n7196), .A2(n7195), .ZN(n7200) );
  OR2_X1 U8837 ( .A1(n7197), .A2(n8701), .ZN(n7569) );
  NAND2_X1 U8838 ( .A1(n8845), .A2(n7569), .ZN(n10279) );
  INV_X1 U8839 ( .A(n7198), .ZN(n7199) );
  MUX2_X1 U8840 ( .A(n6846), .B(n7199), .S(n8915), .Z(n7206) );
  NOR2_X1 U8841 ( .A1(n7200), .A2(n4831), .ZN(n10287) );
  INV_X1 U8842 ( .A(n10287), .ZN(n7763) );
  OAI22_X1 U8843 ( .A1(n7763), .A2(n7202), .B1(n7201), .B2(n8912), .ZN(n7203)
         );
  AOI21_X1 U8844 ( .B1(n10284), .B2(n7204), .A(n7203), .ZN(n7205) );
  OAI211_X1 U8845 ( .C1(n7207), .C2(n8938), .A(n7206), .B(n7205), .ZN(P2_U3294) );
  NAND2_X1 U8846 ( .A1(n9480), .A2(n8039), .ZN(n7208) );
  NAND2_X1 U8847 ( .A1(n7209), .A2(n7208), .ZN(n7389) );
  INV_X1 U8848 ( .A(n7389), .ZN(n7212) );
  INV_X1 U8849 ( .A(n9478), .ZN(n7211) );
  NAND2_X1 U8850 ( .A1(n9478), .A2(n10205), .ZN(n9214) );
  NAND2_X1 U8851 ( .A1(n7212), .A2(n7217), .ZN(n7387) );
  OR2_X1 U8852 ( .A1(n9478), .A2(n7210), .ZN(n7213) );
  NAND2_X1 U8853 ( .A1(n7387), .A2(n7213), .ZN(n7214) );
  OR2_X1 U8854 ( .A1(n9477), .A2(n7322), .ZN(n9218) );
  NAND2_X1 U8855 ( .A1(n9477), .A2(n7322), .ZN(n9219) );
  NAND2_X1 U8856 ( .A1(n9218), .A2(n9219), .ZN(n7363) );
  NAND2_X1 U8857 ( .A1(n7214), .A2(n7363), .ZN(n7358) );
  OAI21_X1 U8858 ( .B1(n7214), .B2(n7363), .A(n7358), .ZN(n7326) );
  INV_X1 U8859 ( .A(n7326), .ZN(n7225) );
  OR2_X1 U8860 ( .A1(n9480), .A2(n10185), .ZN(n7215) );
  XNOR2_X1 U8861 ( .A(n9302), .B(n7363), .ZN(n7221) );
  INV_X1 U8862 ( .A(n9757), .ZN(n9943) );
  NAND2_X1 U8863 ( .A1(n7326), .A2(n9943), .ZN(n7220) );
  AOI22_X1 U8864 ( .A1(n9935), .A2(n9476), .B1(n9478), .B2(n9938), .ZN(n7219)
         );
  OAI211_X1 U8865 ( .C1(n9940), .C2(n7221), .A(n7220), .B(n7219), .ZN(n7318)
         );
  INV_X1 U8866 ( .A(n7318), .ZN(n7224) );
  NAND2_X1 U8867 ( .A1(n7396), .A2(n7322), .ZN(n7471) );
  OR2_X1 U8868 ( .A1(n7396), .A2(n7322), .ZN(n7222) );
  AND2_X1 U8869 ( .A1(n7471), .A2(n7222), .ZN(n7321) );
  AOI22_X1 U8870 ( .A1(n7321), .A2(n9950), .B1(n9994), .B2(n7356), .ZN(n7223)
         );
  OAI211_X1 U8871 ( .C1(n7225), .C2(n9868), .A(n7224), .B(n7223), .ZN(n7227)
         );
  NAND2_X1 U8872 ( .A1(n7227), .A2(n10255), .ZN(n7226) );
  OAI21_X1 U8873 ( .B1(n10255), .B2(n6797), .A(n7226), .ZN(P1_U3526) );
  INV_X1 U8874 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7229) );
  NAND2_X1 U8875 ( .A1(n7227), .A2(n10247), .ZN(n7228) );
  OAI21_X1 U8876 ( .B1(n10247), .B2(n7229), .A(n7228), .ZN(P1_U3463) );
  NOR2_X1 U8877 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6070), .ZN(n7235) );
  AOI21_X1 U8878 ( .B1(n7236), .B2(P2_REG1_REG_10__SCAN_IN), .A(n7230), .ZN(
        n7233) );
  MUX2_X1 U8879 ( .A(n6073), .B(P2_REG1_REG_11__SCAN_IN), .S(n7551), .Z(n7232)
         );
  INV_X1 U8880 ( .A(n7542), .ZN(n7231) );
  AOI211_X1 U8881 ( .C1(n7233), .C2(n7232), .A(n7231), .B(n10262), .ZN(n7234)
         );
  AOI211_X1 U8882 ( .C1(n10260), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n7235), .B(
        n7234), .ZN(n7246) );
  NAND2_X1 U8883 ( .A1(n7236), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7237) );
  NAND2_X1 U8884 ( .A1(n7551), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7240) );
  OR2_X1 U8885 ( .A1(n7551), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7239) );
  NAND2_X1 U8886 ( .A1(n7240), .A2(n7239), .ZN(n7241) );
  INV_X1 U8887 ( .A(n7550), .ZN(n7244) );
  AND2_X1 U8888 ( .A1(n7242), .A2(n7241), .ZN(n7243) );
  OAI21_X1 U8889 ( .B1(n7244), .B2(n7243), .A(n10259), .ZN(n7245) );
  OAI211_X1 U8890 ( .C1(n10261), .C2(n7543), .A(n7246), .B(n7245), .ZN(
        P2_U3256) );
  NAND2_X1 U8891 ( .A1(n7249), .A2(n7248), .ZN(n7250) );
  XNOR2_X1 U8892 ( .A(n7247), .B(n7250), .ZN(n7258) );
  NOR2_X1 U8893 ( .A1(n9151), .A2(n7526), .ZN(n7257) );
  INV_X1 U8894 ( .A(n7251), .ZN(n7252) );
  AOI21_X1 U8895 ( .B1(n10469), .B2(n9472), .A(n7252), .ZN(n7255) );
  INV_X1 U8896 ( .A(n9474), .ZN(n7253) );
  OR2_X1 U8897 ( .A1(n9161), .A2(n7253), .ZN(n7254) );
  OAI211_X1 U8898 ( .C1(n9158), .C2(n7412), .A(n7255), .B(n7254), .ZN(n7256)
         );
  AOI211_X1 U8899 ( .C1(n7258), .C2(n9152), .A(n7257), .B(n7256), .ZN(n7259)
         );
  INV_X1 U8900 ( .A(n7259), .ZN(P1_U3211) );
  INV_X2 U8901 ( .A(n8915), .ZN(n10293) );
  OAI22_X1 U8902 ( .A1(n8915), .A2(n6843), .B1(n7260), .B2(n8912), .ZN(n7261)
         );
  AOI21_X1 U8903 ( .B1(n10284), .B2(n7262), .A(n7261), .ZN(n7265) );
  NAND2_X1 U8904 ( .A1(n7263), .A2(n10287), .ZN(n7264) );
  OAI211_X1 U8905 ( .C1(n7266), .C2(n8938), .A(n7265), .B(n7264), .ZN(n7267)
         );
  INV_X1 U8906 ( .A(n7267), .ZN(n7268) );
  OAI21_X1 U8907 ( .B1(n10293), .B2(n7269), .A(n7268), .ZN(P2_U3292) );
  INV_X1 U8908 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7271) );
  INV_X1 U8909 ( .A(n7270), .ZN(n7272) );
  INV_X1 U8910 ( .A(n8679), .ZN(n8673) );
  OAI222_X1 U8911 ( .A1(n9050), .A2(n7271), .B1(n4481), .B2(n7272), .C1(n8673), 
        .C2(P2_U3152), .ZN(P2_U3340) );
  INV_X1 U8912 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7273) );
  INV_X1 U8913 ( .A(n9523), .ZN(n9527) );
  OAI222_X1 U8914 ( .A1(n9896), .A2(n7273), .B1(n4480), .B2(n7272), .C1(
        P1_U3084), .C2(n9527), .ZN(P1_U3335) );
  XNOR2_X1 U8915 ( .A(n7274), .B(n7292), .ZN(n7277) );
  OR2_X1 U8916 ( .A1(n7573), .A2(n8886), .ZN(n7276) );
  NAND2_X1 U8917 ( .A1(n8645), .A2(n8928), .ZN(n7275) );
  NAND2_X1 U8918 ( .A1(n7276), .A2(n7275), .ZN(n7375) );
  AOI21_X1 U8919 ( .B1(n7277), .B2(n8933), .A(n7375), .ZN(n10349) );
  OAI21_X1 U8920 ( .B1(n7453), .B2(n7279), .A(n9978), .ZN(n7278) );
  NOR2_X1 U8921 ( .A1(n7278), .A2(n7636), .ZN(n10345) );
  NOR2_X1 U8922 ( .A1(n8924), .A2(n7279), .ZN(n7281) );
  OAI22_X1 U8923 ( .A1(n8915), .A2(n6894), .B1(n7379), .B2(n8912), .ZN(n7280)
         );
  AOI211_X1 U8924 ( .C1(n10345), .C2(n10287), .A(n7281), .B(n7280), .ZN(n7295)
         );
  NAND2_X1 U8925 ( .A1(n7460), .A2(n7282), .ZN(n7287) );
  NAND2_X1 U8926 ( .A1(n7284), .A2(n7283), .ZN(n7290) );
  AND2_X1 U8927 ( .A1(n7287), .A2(n4543), .ZN(n7286) );
  NAND2_X1 U8928 ( .A1(n7288), .A2(n7286), .ZN(n7564) );
  NAND2_X1 U8929 ( .A1(n8645), .A2(n10271), .ZN(n7289) );
  AND2_X1 U8930 ( .A1(n7564), .A2(n7561), .ZN(n10344) );
  NAND2_X1 U8931 ( .A1(n7288), .A2(n7287), .ZN(n7452) );
  NAND2_X1 U8932 ( .A1(n7452), .A2(n7289), .ZN(n7291) );
  NAND2_X1 U8933 ( .A1(n7291), .A2(n7290), .ZN(n7293) );
  NAND2_X1 U8934 ( .A1(n7293), .A2(n7292), .ZN(n10343) );
  NAND3_X1 U8935 ( .A1(n10344), .A2(n10343), .A3(n10288), .ZN(n7294) );
  OAI211_X1 U8936 ( .C1(n10349), .C2(n10293), .A(n7295), .B(n7294), .ZN(
        P2_U3290) );
  XOR2_X1 U8937 ( .A(n7081), .B(n7296), .Z(n7297) );
  OAI222_X1 U8938 ( .A1(n8886), .A2(n7298), .B1(n8884), .B2(n8109), .C1(n9966), 
        .C2(n7297), .ZN(n10340) );
  AOI21_X1 U8939 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n10283), .A(n10340), .ZN(
        n7307) );
  OAI21_X1 U8940 ( .B1(n7081), .B2(n7300), .A(n7299), .ZN(n10342) );
  NOR2_X1 U8941 ( .A1(n8924), .A2(n10338), .ZN(n7305) );
  INV_X1 U8942 ( .A(n8936), .ZN(n7984) );
  NAND2_X1 U8943 ( .A1(n8538), .A2(n8107), .ZN(n7301) );
  NAND2_X1 U8944 ( .A1(n7302), .A2(n7301), .ZN(n10339) );
  INV_X1 U8945 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7303) );
  OAI22_X1 U8946 ( .A1(n7984), .A2(n10339), .B1(n7303), .B2(n8915), .ZN(n7304)
         );
  AOI211_X1 U8947 ( .C1(n10288), .C2(n10342), .A(n7305), .B(n7304), .ZN(n7306)
         );
  OAI21_X1 U8948 ( .B1(n7307), .B2(n10293), .A(n7306), .ZN(P2_U3295) );
  INV_X1 U8949 ( .A(n10187), .ZN(n9946) );
  AOI21_X1 U8950 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n9946), .A(n7308), .ZN(
        n7317) );
  NAND2_X1 U8951 ( .A1(n7310), .A2(n7309), .ZN(n7411) );
  NOR2_X1 U8952 ( .A1(n7312), .A2(n7311), .ZN(n7313) );
  AOI21_X1 U8953 ( .B1(n9550), .B2(n9742), .A(n7314), .ZN(n7315) );
  AOI21_X1 U8954 ( .B1(n10193), .B2(P1_REG2_REG_0__SCAN_IN), .A(n7315), .ZN(
        n7316) );
  OAI21_X1 U8955 ( .B1(n7317), .B2(n10193), .A(n7316), .ZN(P1_U3291) );
  MUX2_X1 U8956 ( .A(n7318), .B(P1_REG2_REG_3__SCAN_IN), .S(n10193), .Z(n7319)
         );
  INV_X1 U8957 ( .A(n7319), .ZN(n7328) );
  NOR2_X1 U8958 ( .A1(n9671), .A2(n10178), .ZN(n7320) );
  NAND2_X1 U8959 ( .A1(n9774), .A2(n7320), .ZN(n9782) );
  INV_X1 U8960 ( .A(n9782), .ZN(n9955) );
  NAND2_X1 U8961 ( .A1(n9735), .A2(n7321), .ZN(n7324) );
  OR2_X1 U8962 ( .A1(n9742), .A2(n7322), .ZN(n7323) );
  OAI211_X1 U8963 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n10187), .A(n7324), .B(
        n7323), .ZN(n7325) );
  AOI21_X1 U8964 ( .B1(n7326), .B2(n9955), .A(n7325), .ZN(n7327) );
  NAND2_X1 U8965 ( .A1(n7328), .A2(n7327), .ZN(P1_U3288) );
  XNOR2_X1 U8966 ( .A(n7329), .B(n7330), .ZN(n7331) );
  NAND2_X1 U8967 ( .A1(n7331), .A2(n7332), .ZN(n7429) );
  OAI21_X1 U8968 ( .B1(n7332), .B2(n7331), .A(n7429), .ZN(n7333) );
  NAND2_X1 U8969 ( .A1(n7333), .A2(n9152), .ZN(n7339) );
  INV_X1 U8970 ( .A(n9158), .ZN(n7337) );
  AND2_X1 U8971 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10050) );
  AOI21_X1 U8972 ( .B1(n10469), .B2(n9474), .A(n10050), .ZN(n7334) );
  OAI21_X1 U8973 ( .B1(n7335), .B2(n9161), .A(n7334), .ZN(n7336) );
  AOI21_X1 U8974 ( .B1(n7369), .B2(n7337), .A(n7336), .ZN(n7338) );
  OAI211_X1 U8975 ( .C1(n10217), .C2(n9151), .A(n7339), .B(n7338), .ZN(
        P1_U3225) );
  INV_X1 U8976 ( .A(n10337), .ZN(n7343) );
  OAI22_X1 U8977 ( .A1(n7343), .A2(n9966), .B1(n6530), .B2(n8886), .ZN(n10335)
         );
  AOI21_X1 U8978 ( .B1(n7984), .B2(n8924), .A(n10334), .ZN(n7340) );
  AOI21_X1 U8979 ( .B1(n8915), .B2(n10335), .A(n7340), .ZN(n7342) );
  AOI22_X1 U8980 ( .A1(n10293), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(n10283), .ZN(n7341) );
  OAI211_X1 U8981 ( .C1(n7343), .C2(n8938), .A(n7342), .B(n7341), .ZN(P2_U3296) );
  OAI211_X1 U8982 ( .C1(n7346), .C2(n7345), .A(n7344), .B(n8622), .ZN(n7351)
         );
  NAND2_X1 U8983 ( .A1(n8539), .A2(n8644), .ZN(n7347) );
  OAI21_X1 U8984 ( .B1(n8628), .B2(n7637), .A(n7347), .ZN(n7349) );
  OAI22_X1 U8985 ( .A1(n8614), .A2(n7644), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6009), .ZN(n7348) );
  NOR2_X1 U8986 ( .A1(n7349), .A2(n7348), .ZN(n7350) );
  OAI211_X1 U8987 ( .C1(n10351), .C2(n8634), .A(n7351), .B(n7350), .ZN(
        P2_U3215) );
  INV_X1 U8988 ( .A(n7352), .ZN(n7354) );
  OAI222_X1 U8989 ( .A1(n8701), .A2(P2_U3152), .B1(n4481), .B2(n7354), .C1(
        n7353), .C2(n9050), .ZN(P2_U3339) );
  OAI222_X1 U8990 ( .A1(n9901), .A2(n7355), .B1(n4480), .B2(n7354), .C1(
        P1_U3084), .C2(n9671), .ZN(P1_U3334) );
  OR2_X1 U8991 ( .A1(n9477), .A2(n7356), .ZN(n7357) );
  NAND2_X1 U8992 ( .A1(n7358), .A2(n7357), .ZN(n7468) );
  OR2_X1 U8993 ( .A1(n9476), .A2(n10210), .ZN(n7402) );
  NAND2_X1 U8994 ( .A1(n9476), .A2(n10210), .ZN(n9330) );
  NAND2_X1 U8995 ( .A1(n7402), .A2(n9330), .ZN(n9256) );
  NAND2_X1 U8996 ( .A1(n7468), .A2(n9256), .ZN(n7470) );
  OR2_X1 U8997 ( .A1(n9476), .A2(n7476), .ZN(n7359) );
  NAND2_X1 U8998 ( .A1(n7470), .A2(n7359), .ZN(n7407) );
  NAND2_X1 U8999 ( .A1(n9475), .A2(n10217), .ZN(n9333) );
  INV_X1 U9000 ( .A(n7408), .ZN(n9262) );
  XNOR2_X1 U9001 ( .A(n7407), .B(n9262), .ZN(n10221) );
  INV_X1 U9002 ( .A(n10221), .ZN(n7374) );
  NOR2_X1 U9003 ( .A1(n7361), .A2(n7360), .ZN(n7362) );
  NAND2_X1 U9004 ( .A1(n9774), .A2(n7362), .ZN(n9755) );
  INV_X1 U9005 ( .A(n10217), .ZN(n7409) );
  OAI211_X1 U9006 ( .C1(n4680), .C2(n10217), .A(n9950), .B(n7493), .ZN(n10216)
         );
  INV_X1 U9007 ( .A(n7363), .ZN(n9258) );
  INV_X1 U9008 ( .A(n7403), .ZN(n7365) );
  INV_X1 U9009 ( .A(n9330), .ZN(n9297) );
  AOI21_X1 U9010 ( .B1(n7365), .B2(n7402), .A(n9297), .ZN(n7366) );
  NAND2_X1 U9011 ( .A1(n7366), .A2(n7408), .ZN(n7486) );
  OAI21_X1 U9012 ( .B1(n7408), .B2(n7366), .A(n7486), .ZN(n7367) );
  AOI22_X1 U9013 ( .A1(n7367), .A2(n9772), .B1(n9938), .B2(n9476), .ZN(n10218)
         );
  NAND2_X1 U9014 ( .A1(n9474), .A2(n9935), .ZN(n10215) );
  INV_X1 U9015 ( .A(n10215), .ZN(n7368) );
  AOI21_X1 U9016 ( .B1(n9946), .B2(n7369), .A(n7368), .ZN(n7370) );
  OAI211_X1 U9017 ( .C1(n10180), .C2(n10216), .A(n10218), .B(n7370), .ZN(n7372) );
  OAI22_X1 U9018 ( .A1(n9742), .A2(n10217), .B1(n5206), .B2(n9774), .ZN(n7371)
         );
  AOI21_X1 U9019 ( .B1(n7372), .B2(n9774), .A(n7371), .ZN(n7373) );
  OAI21_X1 U9020 ( .B1(n7374), .B2(n9755), .A(n7373), .ZN(P1_U3286) );
  NAND2_X1 U9021 ( .A1(n7375), .A2(n8631), .ZN(n7378) );
  INV_X1 U9022 ( .A(n7376), .ZN(n7377) );
  OAI211_X1 U9023 ( .C1(n8628), .C2(n7379), .A(n7378), .B(n7377), .ZN(n7385)
         );
  NAND2_X1 U9024 ( .A1(n7381), .A2(n7380), .ZN(n7382) );
  AOI21_X1 U9025 ( .B1(n7383), .B2(n7382), .A(n8620), .ZN(n7384) );
  AOI211_X1 U9026 ( .C1(n10346), .C2(n8618), .A(n7385), .B(n7384), .ZN(n7386)
         );
  INV_X1 U9027 ( .A(n7386), .ZN(P2_U3241) );
  INV_X1 U9028 ( .A(n7387), .ZN(n7388) );
  AOI21_X1 U9029 ( .B1(n9259), .B2(n7389), .A(n7388), .ZN(n10204) );
  AOI22_X1 U9030 ( .A1(n9935), .A2(n9477), .B1(n9480), .B2(n9938), .ZN(n7393)
         );
  OAI21_X1 U9031 ( .B1(n9259), .B2(n9216), .A(n7390), .ZN(n7391) );
  NAND2_X1 U9032 ( .A1(n7391), .A2(n9772), .ZN(n7392) );
  OAI211_X1 U9033 ( .C1(n10204), .C2(n9757), .A(n7393), .B(n7392), .ZN(n10207)
         );
  NAND2_X1 U9034 ( .A1(n10207), .A2(n9774), .ZN(n7401) );
  OAI22_X1 U9035 ( .A1(n10187), .A2(n7394), .B1(n5126), .B2(n9774), .ZN(n7399)
         );
  AND2_X1 U9036 ( .A1(n7210), .A2(n7395), .ZN(n7397) );
  OR2_X1 U9037 ( .A1(n7397), .A2(n7396), .ZN(n10206) );
  NOR2_X1 U9038 ( .A1(n9550), .A2(n10206), .ZN(n7398) );
  AOI211_X1 U9039 ( .C1(n9947), .C2(n7210), .A(n7399), .B(n7398), .ZN(n7400)
         );
  OAI211_X1 U9040 ( .C1(n10204), .C2(n9782), .A(n7401), .B(n7400), .ZN(
        P1_U3289) );
  NOR2_X1 U9041 ( .A1(n9217), .A2(n9330), .ZN(n7404) );
  NAND2_X1 U9042 ( .A1(n9474), .A2(n10222), .ZN(n9224) );
  NAND2_X1 U9043 ( .A1(n7405), .A2(n9224), .ZN(n7619) );
  NAND2_X1 U9044 ( .A1(n9473), .A2(n7526), .ZN(n9339) );
  NAND2_X1 U9045 ( .A1(n9335), .A2(n9339), .ZN(n9264) );
  XNOR2_X1 U9046 ( .A(n7619), .B(n9264), .ZN(n7406) );
  AOI222_X1 U9047 ( .A1(n9772), .A2(n7406), .B1(n9474), .B2(n9938), .C1(n9472), 
        .C2(n9935), .ZN(n7530) );
  NAND2_X1 U9048 ( .A1(n9336), .A2(n9224), .ZN(n9325) );
  INV_X1 U9049 ( .A(n10222), .ZN(n7498) );
  NAND2_X1 U9050 ( .A1(n7410), .A2(n9264), .ZN(n7615) );
  OAI21_X1 U9051 ( .B1(n7410), .B2(n9264), .A(n7615), .ZN(n7528) );
  INV_X1 U9052 ( .A(n9755), .ZN(n7417) );
  OAI211_X1 U9053 ( .C1(n7494), .C2(n7526), .A(n9950), .B(n7627), .ZN(n7525)
         );
  NOR2_X1 U9054 ( .A1(n7411), .A2(n10180), .ZN(n9954) );
  INV_X1 U9055 ( .A(n9954), .ZN(n7911) );
  INV_X1 U9056 ( .A(n7526), .ZN(n7613) );
  OAI22_X1 U9057 ( .A1(n9774), .A2(n7413), .B1(n7412), .B2(n10187), .ZN(n7414)
         );
  AOI21_X1 U9058 ( .B1(n9947), .B2(n7613), .A(n7414), .ZN(n7415) );
  OAI21_X1 U9059 ( .B1(n7525), .B2(n7911), .A(n7415), .ZN(n7416) );
  AOI21_X1 U9060 ( .B1(n7528), .B2(n7417), .A(n7416), .ZN(n7418) );
  OAI21_X1 U9061 ( .B1(n7530), .B2(n10193), .A(n7418), .ZN(P1_U3284) );
  NAND2_X1 U9062 ( .A1(n7420), .A2(n7419), .ZN(n7422) );
  XNOR2_X1 U9063 ( .A(n7422), .B(n7421), .ZN(n7428) );
  INV_X1 U9064 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7423) );
  NOR2_X1 U9065 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7423), .ZN(n10087) );
  INV_X1 U9066 ( .A(n9937), .ZN(n7777) );
  NOR2_X1 U9067 ( .A1(n9117), .A2(n7777), .ZN(n7424) );
  AOI211_X1 U9068 ( .C1(n9134), .C2(n9473), .A(n10087), .B(n7424), .ZN(n7425)
         );
  OAI21_X1 U9069 ( .B1(n9158), .B2(n7625), .A(n7425), .ZN(n7426) );
  AOI21_X1 U9070 ( .B1(n7778), .B2(n9165), .A(n7426), .ZN(n7427) );
  OAI21_X1 U9071 ( .B1(n7428), .B2(n9139), .A(n7427), .ZN(P1_U3219) );
  OAI21_X1 U9072 ( .B1(n7430), .B2(n7329), .A(n7429), .ZN(n7434) );
  XNOR2_X1 U9073 ( .A(n7432), .B(n7431), .ZN(n7433) );
  XNOR2_X1 U9074 ( .A(n7434), .B(n7433), .ZN(n7441) );
  NOR2_X1 U9075 ( .A1(n9151), .A2(n10222), .ZN(n7440) );
  INV_X1 U9076 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7435) );
  NOR2_X1 U9077 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7435), .ZN(n10068) );
  AOI21_X1 U9078 ( .B1(n10469), .B2(n9473), .A(n10068), .ZN(n7438) );
  OR2_X1 U9079 ( .A1(n9161), .A2(n7436), .ZN(n7437) );
  OAI211_X1 U9080 ( .C1(n9158), .C2(n7491), .A(n7438), .B(n7437), .ZN(n7439)
         );
  AOI211_X1 U9081 ( .C1(n7441), .C2(n9152), .A(n7440), .B(n7439), .ZN(n7442)
         );
  INV_X1 U9082 ( .A(n7442), .ZN(P1_U3237) );
  OAI211_X1 U9083 ( .C1(n7445), .C2(n7444), .A(n7443), .B(n8622), .ZN(n7451)
         );
  NAND2_X1 U9084 ( .A1(n8539), .A2(n8643), .ZN(n7446) );
  OAI21_X1 U9085 ( .B1(n8628), .B2(n7577), .A(n7446), .ZN(n7449) );
  OAI21_X1 U9086 ( .B1(n8614), .B2(n7664), .A(n7447), .ZN(n7448) );
  NOR2_X1 U9087 ( .A1(n7449), .A2(n7448), .ZN(n7450) );
  OAI211_X1 U9088 ( .C1(n10359), .C2(n8634), .A(n7451), .B(n7450), .ZN(
        P2_U3223) );
  XOR2_X1 U9089 ( .A(n7458), .B(n7452), .Z(n10269) );
  AOI211_X1 U9090 ( .C1(n10271), .C2(n7454), .A(n4832), .B(n7453), .ZN(n10270)
         );
  NAND2_X1 U9091 ( .A1(n7456), .A2(n7455), .ZN(n7457) );
  XOR2_X1 U9092 ( .A(n7458), .B(n7457), .Z(n7459) );
  OAI222_X1 U9093 ( .A1(n8886), .A2(n6559), .B1(n8884), .B2(n7460), .C1(n9966), 
        .C2(n7459), .ZN(n10276) );
  AOI211_X1 U9094 ( .C1(n10385), .C2(n10271), .A(n10270), .B(n10276), .ZN(
        n7461) );
  OAI21_X1 U9095 ( .B1(n9020), .B2(n10269), .A(n7461), .ZN(n7463) );
  NAND2_X1 U9096 ( .A1(n7463), .A2(n10406), .ZN(n7462) );
  OAI21_X1 U9097 ( .B1(n10406), .B2(n5987), .A(n7462), .ZN(P2_U3525) );
  NAND2_X1 U9098 ( .A1(n7463), .A2(n10395), .ZN(n7464) );
  OAI21_X1 U9099 ( .B1(n10395), .B2(n5983), .A(n7464), .ZN(P2_U3466) );
  INV_X1 U9100 ( .A(n7465), .ZN(n7503) );
  OAI222_X1 U9101 ( .A1(n4480), .A2(n7503), .B1(n7467), .B2(P1_U3084), .C1(
        n7466), .C2(n9896), .ZN(P1_U3333) );
  OR2_X1 U9102 ( .A1(n7468), .A2(n9256), .ZN(n7469) );
  NAND2_X1 U9103 ( .A1(n7470), .A2(n7469), .ZN(n10214) );
  NAND2_X1 U9104 ( .A1(n7471), .A2(n7476), .ZN(n7472) );
  NAND2_X1 U9105 ( .A1(n7473), .A2(n7472), .ZN(n10211) );
  INV_X1 U9106 ( .A(n7474), .ZN(n7475) );
  AOI22_X1 U9107 ( .A1(n9947), .A2(n7476), .B1(n7475), .B2(n9946), .ZN(n7477)
         );
  OAI21_X1 U9108 ( .B1(n9550), .B2(n10211), .A(n7477), .ZN(n7482) );
  XNOR2_X1 U9109 ( .A(n7403), .B(n9256), .ZN(n7480) );
  NAND2_X1 U9110 ( .A1(n10214), .A2(n9943), .ZN(n7479) );
  AOI22_X1 U9111 ( .A1(n9938), .A2(n9477), .B1(n9475), .B2(n9935), .ZN(n7478)
         );
  OAI211_X1 U9112 ( .C1(n7480), .C2(n9940), .A(n7479), .B(n7478), .ZN(n10212)
         );
  MUX2_X1 U9113 ( .A(n10212), .B(P1_REG2_REG_4__SCAN_IN), .S(n10193), .Z(n7481) );
  AOI211_X1 U9114 ( .C1(n9955), .C2(n10214), .A(n7482), .B(n7481), .ZN(n7483)
         );
  INV_X1 U9115 ( .A(n7483), .ZN(P1_U3287) );
  OAI21_X1 U9116 ( .B1(n7485), .B2(n9325), .A(n7484), .ZN(n10226) );
  INV_X1 U9117 ( .A(n10226), .ZN(n7501) );
  NAND2_X1 U9118 ( .A1(n7486), .A2(n9296), .ZN(n7487) );
  XNOR2_X1 U9119 ( .A(n7487), .B(n9325), .ZN(n7490) );
  NAND2_X1 U9120 ( .A1(n10226), .A2(n9943), .ZN(n7489) );
  AOI22_X1 U9121 ( .A1(n9935), .A2(n9473), .B1(n9475), .B2(n9938), .ZN(n7488)
         );
  OAI211_X1 U9122 ( .C1(n7490), .C2(n9940), .A(n7489), .B(n7488), .ZN(n10224)
         );
  NAND2_X1 U9123 ( .A1(n10224), .A2(n9774), .ZN(n7500) );
  OAI22_X1 U9124 ( .A1(n9774), .A2(n7492), .B1(n7491), .B2(n10187), .ZN(n7497)
         );
  AND2_X1 U9125 ( .A1(n7493), .A2(n7498), .ZN(n7495) );
  OR2_X1 U9126 ( .A1(n7495), .A2(n7494), .ZN(n10223) );
  NOR2_X1 U9127 ( .A1(n10223), .A2(n9550), .ZN(n7496) );
  AOI211_X1 U9128 ( .C1(n9947), .C2(n7498), .A(n7497), .B(n7496), .ZN(n7499)
         );
  OAI211_X1 U9129 ( .C1(n7501), .C2(n9782), .A(n7500), .B(n7499), .ZN(P1_U3285) );
  OAI222_X1 U9130 ( .A1(P2_U3152), .A2(n7504), .B1(n4481), .B2(n7503), .C1(
        n7502), .C2(n9050), .ZN(P2_U3338) );
  XNOR2_X1 U9131 ( .A(n10114), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n10110) );
  NOR2_X1 U9132 ( .A1(n10111), .A2(n10110), .ZN(n10109) );
  AOI22_X1 U9133 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7512), .B1(n10127), .B2(
        n7947), .ZN(n10123) );
  NOR2_X1 U9134 ( .A1(n10124), .A2(n10123), .ZN(n10122) );
  XNOR2_X1 U9135 ( .A(n7518), .B(n9506), .ZN(n7507) );
  NAND2_X1 U9136 ( .A1(n7507), .A2(n5453), .ZN(n9507) );
  OAI21_X1 U9137 ( .B1(n7507), .B2(n5453), .A(n9507), .ZN(n7523) );
  INV_X1 U9138 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7521) );
  AOI21_X1 U9139 ( .B1(n10009), .B2(n7509), .A(n7508), .ZN(n10117) );
  MUX2_X1 U9140 ( .A(n7510), .B(P1_REG1_REG_12__SCAN_IN), .S(n10114), .Z(
        n10116) );
  NOR2_X1 U9141 ( .A1(n10117), .A2(n10116), .ZN(n10115) );
  AOI21_X1 U9142 ( .B1(n7510), .B2(n7511), .A(n10115), .ZN(n10130) );
  XNOR2_X1 U9143 ( .A(n10127), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n10129) );
  NOR2_X1 U9144 ( .A1(n10130), .A2(n10129), .ZN(n10128) );
  AOI21_X1 U9145 ( .B1(n7513), .B2(n7512), .A(n10128), .ZN(n7515) );
  AOI22_X1 U9146 ( .A1(n7518), .A2(n9496), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n9505), .ZN(n7514) );
  NOR2_X1 U9147 ( .A1(n7515), .A2(n7514), .ZN(n9495) );
  AOI21_X1 U9148 ( .B1(n7515), .B2(n7514), .A(n9495), .ZN(n7516) );
  OR2_X1 U9149 ( .A1(n7516), .A2(n10131), .ZN(n7520) );
  NAND2_X1 U9150 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9061) );
  INV_X1 U9151 ( .A(n9061), .ZN(n7517) );
  AOI21_X1 U9152 ( .B1(n10168), .B2(n7518), .A(n7517), .ZN(n7519) );
  OAI211_X1 U9153 ( .C1(n7521), .C2(n10175), .A(n7520), .B(n7519), .ZN(n7522)
         );
  AOI21_X1 U9154 ( .B1(n10088), .B2(n7523), .A(n7522), .ZN(n7524) );
  INV_X1 U9155 ( .A(n7524), .ZN(P1_U3255) );
  INV_X1 U9156 ( .A(n9994), .ZN(n10237) );
  OAI21_X1 U9157 ( .B1(n7526), .B2(n10237), .A(n7525), .ZN(n7527) );
  AOI21_X1 U9158 ( .B1(n7528), .B2(n4981), .A(n7527), .ZN(n7529) );
  NAND2_X1 U9159 ( .A1(n7530), .A2(n7529), .ZN(n7558) );
  NAND2_X1 U9160 ( .A1(n7558), .A2(n10255), .ZN(n7531) );
  OAI21_X1 U9161 ( .B1(n10255), .B2(n5257), .A(n7531), .ZN(P1_U3530) );
  XNOR2_X1 U9162 ( .A(n7534), .B(n7533), .ZN(n7535) );
  XNOR2_X1 U9163 ( .A(n7532), .B(n7535), .ZN(n7541) );
  NOR2_X1 U9164 ( .A1(n7777), .A2(n9161), .ZN(n7536) );
  AOI211_X1 U9165 ( .C1(n10469), .C2(n9936), .A(n7537), .B(n7536), .ZN(n7538)
         );
  OAI21_X1 U9166 ( .B1(n9158), .B2(n9944), .A(n7538), .ZN(n7539) );
  AOI21_X1 U9167 ( .B1(n9948), .B2(n9165), .A(n7539), .ZN(n7540) );
  OAI21_X1 U9168 ( .B1(n7541), .B2(n9139), .A(n7540), .ZN(P1_U3215) );
  OAI21_X1 U9169 ( .B1(n6073), .B2(n7543), .A(n7542), .ZN(n7546) );
  MUX2_X1 U9170 ( .A(n7544), .B(P2_REG1_REG_12__SCAN_IN), .S(n7603), .Z(n7545)
         );
  NOR2_X1 U9171 ( .A1(n7546), .A2(n7545), .ZN(n7598) );
  AOI21_X1 U9172 ( .B1(n7546), .B2(n7545), .A(n7598), .ZN(n7549) );
  NOR2_X1 U9173 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7770), .ZN(n7547) );
  AOI21_X1 U9174 ( .B1(n10260), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7547), .ZN(
        n7548) );
  OAI21_X1 U9175 ( .B1(n10262), .B2(n7549), .A(n7548), .ZN(n7556) );
  NAND2_X1 U9176 ( .A1(n7603), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7552) );
  OAI21_X1 U9177 ( .B1(n7603), .B2(P2_REG2_REG_12__SCAN_IN), .A(n7552), .ZN(
        n7553) );
  AOI211_X1 U9178 ( .C1(n7554), .C2(n7553), .A(n7602), .B(n10263), .ZN(n7555)
         );
  AOI211_X1 U9179 ( .C1(n9921), .C2(n7603), .A(n7556), .B(n7555), .ZN(n7557)
         );
  INV_X1 U9180 ( .A(n7557), .ZN(P2_U3257) );
  INV_X1 U9181 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7560) );
  NAND2_X1 U9182 ( .A1(n7558), .A2(n10247), .ZN(n7559) );
  OAI21_X1 U9183 ( .B1(n10247), .B2(n7560), .A(n7559), .ZN(P1_U3475) );
  NOR2_X1 U9184 ( .A1(n5034), .A2(n7562), .ZN(n7563) );
  AND2_X2 U9185 ( .A1(n7564), .A2(n7563), .ZN(n7634) );
  NAND2_X1 U9186 ( .A1(n7573), .A2(n10351), .ZN(n7566) );
  NAND2_X1 U9187 ( .A1(n7567), .A2(n7572), .ZN(n7568) );
  NAND2_X1 U9188 ( .A1(n7676), .A2(n7568), .ZN(n10358) );
  OR2_X1 U9189 ( .A1(n10293), .A2(n7569), .ZN(n8862) );
  OAI21_X1 U9190 ( .B1(n7572), .B2(n7571), .A(n7570), .ZN(n7575) );
  OAI22_X1 U9191 ( .A1(n7664), .A2(n8886), .B1(n7573), .B2(n8884), .ZN(n7574)
         );
  AOI21_X1 U9192 ( .B1(n7575), .B2(n8933), .A(n7574), .ZN(n7576) );
  OAI21_X1 U9193 ( .B1(n10358), .B2(n8845), .A(n7576), .ZN(n10361) );
  NAND2_X1 U9194 ( .A1(n10361), .A2(n8915), .ZN(n7583) );
  OAI22_X1 U9195 ( .A1(n8915), .A2(n7578), .B1(n7577), .B2(n8912), .ZN(n7581)
         );
  NAND2_X1 U9196 ( .A1(n7635), .A2(n7672), .ZN(n7579) );
  NAND2_X1 U9197 ( .A1(n7688), .A2(n7579), .ZN(n10360) );
  NOR2_X1 U9198 ( .A1(n10360), .A2(n7984), .ZN(n7580) );
  AOI211_X1 U9199 ( .C1(n10284), .C2(n7672), .A(n7581), .B(n7580), .ZN(n7582)
         );
  OAI211_X1 U9200 ( .C1(n10358), .C2(n8862), .A(n7583), .B(n7582), .ZN(
        P2_U3288) );
  INV_X1 U9201 ( .A(n7708), .ZN(n10366) );
  NAND2_X1 U9202 ( .A1(n4566), .A2(n7584), .ZN(n7585) );
  XNOR2_X1 U9203 ( .A(n4583), .B(n7585), .ZN(n7587) );
  NAND2_X1 U9204 ( .A1(n7587), .A2(n8622), .ZN(n7593) );
  NAND2_X1 U9205 ( .A1(n8539), .A2(n8642), .ZN(n7588) );
  OAI21_X1 U9206 ( .B1(n8628), .B2(n7686), .A(n7588), .ZN(n7591) );
  OAI21_X1 U9207 ( .B1(n8614), .B2(n7754), .A(n7589), .ZN(n7590) );
  NOR2_X1 U9208 ( .A1(n7591), .A2(n7590), .ZN(n7592) );
  OAI211_X1 U9209 ( .C1(n10366), .C2(n8634), .A(n7593), .B(n7592), .ZN(
        P2_U3233) );
  INV_X1 U9210 ( .A(n7594), .ZN(n7596) );
  OAI222_X1 U9211 ( .A1(n4480), .A2(n7596), .B1(n9290), .B2(P1_U3084), .C1(
        n8162), .C2(n9896), .ZN(P1_U3332) );
  OAI222_X1 U9212 ( .A1(P2_U3152), .A2(n7597), .B1(n4481), .B2(n7596), .C1(
        n7595), .C2(n9050), .ZN(P2_U3337) );
  AOI21_X1 U9213 ( .B1(n7599), .B2(n7544), .A(n7598), .ZN(n7601) );
  AOI22_X1 U9214 ( .A1(n7734), .A2(n7728), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7729), .ZN(n7600) );
  NOR2_X1 U9215 ( .A1(n7601), .A2(n7600), .ZN(n7727) );
  AOI21_X1 U9216 ( .B1(n7601), .B2(n7600), .A(n7727), .ZN(n7612) );
  AOI22_X1 U9217 ( .A1(n7734), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7981), .B2(
        n7729), .ZN(n7604) );
  OAI21_X1 U9218 ( .B1(n7605), .B2(n7604), .A(n7733), .ZN(n7606) );
  NAND2_X1 U9219 ( .A1(n7606), .A2(n10259), .ZN(n7611) );
  INV_X1 U9220 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7608) );
  OAI22_X1 U9221 ( .A1(n8705), .A2(n7608), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7607), .ZN(n7609) );
  AOI21_X1 U9222 ( .B1(n9921), .B2(n7734), .A(n7609), .ZN(n7610) );
  OAI211_X1 U9223 ( .C1(n7612), .C2(n10262), .A(n7611), .B(n7610), .ZN(
        P2_U3258) );
  OR2_X1 U9224 ( .A1(n9473), .A2(n7613), .ZN(n7614) );
  NAND2_X1 U9225 ( .A1(n7615), .A2(n7614), .ZN(n7617) );
  NAND2_X1 U9226 ( .A1(n10229), .A2(n9472), .ZN(n9343) );
  INV_X1 U9227 ( .A(n9472), .ZN(n7781) );
  NAND2_X1 U9228 ( .A1(n7781), .A2(n7778), .ZN(n9349) );
  NAND2_X1 U9229 ( .A1(n7617), .A2(n9266), .ZN(n7618) );
  NAND2_X1 U9230 ( .A1(n7780), .A2(n7618), .ZN(n10228) );
  AOI22_X1 U9231 ( .A1(n9938), .A2(n9473), .B1(n9937), .B2(n9935), .ZN(n7624)
         );
  AND2_X1 U9232 ( .A1(n7621), .A2(n9335), .ZN(n7622) );
  INV_X1 U9233 ( .A(n9335), .ZN(n9328) );
  NOR2_X1 U9234 ( .A1(n7616), .A2(n9328), .ZN(n7620) );
  NAND2_X1 U9235 ( .A1(n7621), .A2(n7620), .ZN(n9932) );
  OAI211_X1 U9236 ( .C1(n7622), .C2(n9266), .A(n9932), .B(n9772), .ZN(n7623)
         );
  OAI211_X1 U9237 ( .C1(n10228), .C2(n9757), .A(n7624), .B(n7623), .ZN(n10231)
         );
  NAND2_X1 U9238 ( .A1(n10231), .A2(n9774), .ZN(n7632) );
  OAI22_X1 U9239 ( .A1(n9774), .A2(n7626), .B1(n7625), .B2(n10187), .ZN(n7630)
         );
  NAND2_X1 U9240 ( .A1(n7627), .A2(n7778), .ZN(n7628) );
  NAND2_X1 U9241 ( .A1(n7787), .A2(n7628), .ZN(n10230) );
  NOR2_X1 U9242 ( .A1(n10230), .A2(n9550), .ZN(n7629) );
  AOI211_X1 U9243 ( .C1(n9947), .C2(n7778), .A(n7630), .B(n7629), .ZN(n7631)
         );
  OAI211_X1 U9244 ( .C1(n10228), .C2(n9782), .A(n7632), .B(n7631), .ZN(
        P1_U3283) );
  OAI21_X1 U9245 ( .B1(n7634), .B2(n7565), .A(n7633), .ZN(n10355) );
  OAI21_X1 U9246 ( .B1(n7636), .B2(n10351), .A(n7635), .ZN(n10352) );
  INV_X1 U9247 ( .A(n7637), .ZN(n7638) );
  AOI22_X1 U9248 ( .A1(n10284), .A2(n7639), .B1(n10283), .B2(n7638), .ZN(n7640) );
  OAI21_X1 U9249 ( .B1(n10352), .B2(n7984), .A(n7640), .ZN(n7646) );
  XOR2_X1 U9250 ( .A(n7642), .B(n7641), .Z(n7643) );
  OAI222_X1 U9251 ( .A1(n8886), .A2(n7644), .B1(n7643), .B2(n9966), .C1(n8884), 
        .C2(n6559), .ZN(n10353) );
  MUX2_X1 U9252 ( .A(n10353), .B(P2_REG2_REG_7__SCAN_IN), .S(n10293), .Z(n7645) );
  AOI211_X1 U9253 ( .C1(n10288), .C2(n10355), .A(n7646), .B(n7645), .ZN(n7647)
         );
  INV_X1 U9254 ( .A(n7647), .ZN(P2_U3289) );
  XNOR2_X1 U9255 ( .A(n7649), .B(n7648), .ZN(n7655) );
  INV_X1 U9256 ( .A(n7899), .ZN(n7940) );
  NOR2_X1 U9257 ( .A1(n7816), .A2(n9161), .ZN(n7650) );
  AOI211_X1 U9258 ( .C1(n10469), .C2(n7940), .A(n7651), .B(n7650), .ZN(n7652)
         );
  OAI21_X1 U9259 ( .B1(n9158), .B2(n7822), .A(n7652), .ZN(n7653) );
  AOI21_X1 U9260 ( .B1(n7895), .B2(n9165), .A(n7653), .ZN(n7654) );
  OAI21_X1 U9261 ( .B1(n7655), .B2(n9139), .A(n7654), .ZN(P1_U3234) );
  INV_X1 U9262 ( .A(n7656), .ZN(n7660) );
  OAI222_X1 U9263 ( .A1(n9901), .A2(n7658), .B1(n4480), .B2(n7660), .C1(
        P1_U3084), .C2(n9452), .ZN(P1_U3331) );
  OAI222_X1 U9264 ( .A1(n7661), .A2(P2_U3152), .B1(n4481), .B2(n7660), .C1(
        n7659), .C2(n9050), .ZN(P2_U3336) );
  XNOR2_X1 U9265 ( .A(n7663), .B(n7662), .ZN(n7671) );
  INV_X1 U9266 ( .A(n7664), .ZN(n8641) );
  NAND2_X1 U9267 ( .A1(n8539), .A2(n8641), .ZN(n7665) );
  OAI21_X1 U9268 ( .B1(n8628), .B2(n7718), .A(n7665), .ZN(n7668) );
  OAI21_X1 U9269 ( .B1(n8614), .B2(n7889), .A(n7666), .ZN(n7667) );
  NOR2_X1 U9270 ( .A1(n7668), .A2(n7667), .ZN(n7670) );
  NAND2_X1 U9271 ( .A1(n7724), .A2(n8618), .ZN(n7669) );
  OAI211_X1 U9272 ( .C1(n7671), .C2(n8620), .A(n7670), .B(n7669), .ZN(P2_U3219) );
  NAND2_X1 U9273 ( .A1(n7672), .A2(n8642), .ZN(n7673) );
  NAND2_X1 U9274 ( .A1(n7676), .A2(n7673), .ZN(n7678) );
  INV_X1 U9275 ( .A(n7680), .ZN(n7674) );
  AND2_X1 U9276 ( .A1(n7674), .A2(n7673), .ZN(n7675) );
  INV_X1 U9277 ( .A(n7710), .ZN(n7677) );
  AOI21_X1 U9278 ( .B1(n7680), .B2(n7678), .A(n7677), .ZN(n10365) );
  INV_X1 U9279 ( .A(n7754), .ZN(n8640) );
  AOI22_X1 U9280 ( .A1(n8928), .A2(n8642), .B1(n8640), .B2(n8930), .ZN(n7685)
         );
  INV_X1 U9281 ( .A(n7570), .ZN(n7681) );
  NOR3_X1 U9282 ( .A1(n7681), .A2(n7680), .A3(n7679), .ZN(n7683) );
  INV_X1 U9283 ( .A(n7682), .ZN(n7712) );
  OAI21_X1 U9284 ( .B1(n7683), .B2(n7712), .A(n8933), .ZN(n7684) );
  OAI211_X1 U9285 ( .C1(n10365), .C2(n8845), .A(n7685), .B(n7684), .ZN(n10368)
         );
  NAND2_X1 U9286 ( .A1(n10368), .A2(n8915), .ZN(n7693) );
  INV_X1 U9287 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7687) );
  OAI22_X1 U9288 ( .A1(n8915), .A2(n7687), .B1(n7686), .B2(n8912), .ZN(n7691)
         );
  AND2_X1 U9289 ( .A1(n7688), .A2(n7708), .ZN(n7689) );
  NOR2_X1 U9290 ( .A1(n7688), .A2(n7708), .ZN(n7720) );
  OR2_X1 U9291 ( .A1(n7689), .A2(n7720), .ZN(n10367) );
  NOR2_X1 U9292 ( .A1(n10367), .A2(n7984), .ZN(n7690) );
  AOI211_X1 U9293 ( .C1(n10284), .C2(n7708), .A(n7691), .B(n7690), .ZN(n7692)
         );
  OAI211_X1 U9294 ( .C1(n10365), .C2(n8862), .A(n7693), .B(n7692), .ZN(
        P2_U3287) );
  INV_X1 U9295 ( .A(n7816), .ZN(n7808) );
  AND2_X1 U9296 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10101) );
  AOI21_X1 U9297 ( .B1(n7808), .B2(n10469), .A(n10101), .ZN(n7695) );
  OR2_X1 U9298 ( .A1(n9161), .A2(n7781), .ZN(n7694) );
  OAI211_X1 U9299 ( .C1(n9158), .C2(n7785), .A(n7695), .B(n7694), .ZN(n7700)
         );
  XOR2_X1 U9300 ( .A(n7696), .B(n7697), .Z(n7698) );
  NOR2_X1 U9301 ( .A1(n7698), .A2(n9139), .ZN(n7699) );
  AOI211_X1 U9302 ( .C1(n10236), .C2(n9165), .A(n7700), .B(n7699), .ZN(n7701)
         );
  INV_X1 U9303 ( .A(n7701), .ZN(P1_U3229) );
  XNOR2_X1 U9304 ( .A(n7703), .B(n7702), .ZN(n7707) );
  OAI22_X1 U9305 ( .A1(n8614), .A2(n7976), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6070), .ZN(n7705) );
  OAI22_X1 U9306 ( .A1(n8615), .A2(n7754), .B1(n7760), .B2(n8628), .ZN(n7704)
         );
  AOI211_X1 U9307 ( .C1(n7877), .C2(n8618), .A(n7705), .B(n7704), .ZN(n7706)
         );
  OAI21_X1 U9308 ( .B1(n7707), .B2(n8620), .A(n7706), .ZN(P2_U3238) );
  OR2_X1 U9309 ( .A1(n7708), .A2(n8641), .ZN(n7709) );
  XNOR2_X1 U9310 ( .A(n7756), .B(n7755), .ZN(n10371) );
  INV_X1 U9311 ( .A(n7889), .ZN(n8639) );
  AOI22_X1 U9312 ( .A1(n8928), .A2(n8641), .B1(n8639), .B2(n8930), .ZN(n7717)
         );
  NOR3_X1 U9313 ( .A1(n7712), .A2(n7755), .A3(n7711), .ZN(n7715) );
  INV_X1 U9314 ( .A(n7713), .ZN(n7714) );
  OAI21_X1 U9315 ( .B1(n7715), .B2(n7714), .A(n8933), .ZN(n7716) );
  OAI211_X1 U9316 ( .C1(n10371), .C2(n8845), .A(n7717), .B(n7716), .ZN(n10374)
         );
  NAND2_X1 U9317 ( .A1(n10374), .A2(n8915), .ZN(n7726) );
  OAI22_X1 U9318 ( .A1(n8915), .A2(n7719), .B1(n7718), .B2(n8912), .ZN(n7723)
         );
  INV_X1 U9319 ( .A(n7724), .ZN(n10372) );
  NOR2_X1 U9320 ( .A1(n7720), .A2(n10372), .ZN(n7721) );
  OR2_X1 U9321 ( .A1(n7762), .A2(n7721), .ZN(n10373) );
  NOR2_X1 U9322 ( .A1(n10373), .A2(n7984), .ZN(n7722) );
  AOI211_X1 U9323 ( .C1(n10284), .C2(n7724), .A(n7723), .B(n7722), .ZN(n7725)
         );
  OAI211_X1 U9324 ( .C1(n10371), .C2(n8862), .A(n7726), .B(n7725), .ZN(
        P2_U3286) );
  AOI21_X1 U9325 ( .B1(n7729), .B2(n7728), .A(n7727), .ZN(n7731) );
  AOI22_X1 U9326 ( .A1(n7866), .A2(n6111), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7873), .ZN(n7730) );
  NOR2_X1 U9327 ( .A1(n7731), .A2(n7730), .ZN(n7872) );
  AOI21_X1 U9328 ( .B1(n7731), .B2(n7730), .A(n7872), .ZN(n7742) );
  NOR2_X1 U9329 ( .A1(n7866), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7732) );
  AOI21_X1 U9330 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7866), .A(n7732), .ZN(
        n7736) );
  NAND2_X1 U9331 ( .A1(n7736), .A2(n7735), .ZN(n7865) );
  OAI21_X1 U9332 ( .B1(n7736), .B2(n7735), .A(n7865), .ZN(n7740) );
  INV_X1 U9333 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U9334 ( .A1(n9921), .A2(n7866), .ZN(n7737) );
  NAND2_X1 U9335 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7929) );
  OAI211_X1 U9336 ( .C1(n7738), .C2(n8705), .A(n7737), .B(n7929), .ZN(n7739)
         );
  AOI21_X1 U9337 ( .B1(n7740), .B2(n10259), .A(n7739), .ZN(n7741) );
  OAI21_X1 U9338 ( .B1(n7742), .B2(n10262), .A(n7741), .ZN(P2_U3259) );
  NAND2_X1 U9339 ( .A1(n7746), .A2(n8014), .ZN(n7744) );
  OR2_X1 U9340 ( .A1(n7743), .A2(P1_U3084), .ZN(n9465) );
  OAI211_X1 U9341 ( .C1(n7745), .C2(n9896), .A(n7744), .B(n9465), .ZN(P1_U3330) );
  NAND2_X1 U9342 ( .A1(n7746), .A2(n8010), .ZN(n7748) );
  OAI211_X1 U9343 ( .C1(n7749), .C2(n9050), .A(n7748), .B(n7747), .ZN(P2_U3335) );
  NAND3_X1 U9344 ( .A1(n7713), .A2(n7757), .A3(n7750), .ZN(n7751) );
  NAND2_X1 U9345 ( .A1(n7752), .A2(n7751), .ZN(n7753) );
  INV_X1 U9346 ( .A(n7976), .ZN(n8638) );
  AOI222_X1 U9347 ( .A1(n8933), .A2(n7753), .B1(n8638), .B2(n8930), .C1(n8640), 
        .C2(n8928), .ZN(n10380) );
  OAI21_X1 U9348 ( .B1(n7758), .B2(n7757), .A(n7879), .ZN(n7759) );
  INV_X1 U9349 ( .A(n7759), .ZN(n10384) );
  NAND2_X1 U9350 ( .A1(n10384), .A2(n10288), .ZN(n7767) );
  INV_X1 U9351 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7761) );
  OAI22_X1 U9352 ( .A1(n8915), .A2(n7761), .B1(n7760), .B2(n8912), .ZN(n7765)
         );
  INV_X1 U9353 ( .A(n7877), .ZN(n10382) );
  NAND2_X1 U9354 ( .A1(n7762), .A2(n10382), .ZN(n7881) );
  OAI211_X1 U9355 ( .C1(n7762), .C2(n10382), .A(n9978), .B(n7881), .ZN(n10379)
         );
  NOR2_X1 U9356 ( .A1(n10379), .A2(n7763), .ZN(n7764) );
  AOI211_X1 U9357 ( .C1(n10284), .C2(n7877), .A(n7765), .B(n7764), .ZN(n7766)
         );
  OAI211_X1 U9358 ( .C1(n10380), .C2(n10293), .A(n7767), .B(n7766), .ZN(
        P2_U3285) );
  XNOR2_X1 U9359 ( .A(n7769), .B(n7768), .ZN(n7774) );
  OAI22_X1 U9360 ( .A1(n8614), .A2(n8115), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7770), .ZN(n7772) );
  OAI22_X1 U9361 ( .A1(n8615), .A2(n7889), .B1(n7883), .B2(n8628), .ZN(n7771)
         );
  AOI211_X1 U9362 ( .C1(n10386), .C2(n8618), .A(n7772), .B(n7771), .ZN(n7773)
         );
  OAI21_X1 U9363 ( .B1(n7774), .B2(n8620), .A(n7773), .ZN(P2_U3226) );
  INV_X1 U9364 ( .A(n7775), .ZN(n7804) );
  OR2_X1 U9365 ( .A1(n10236), .A2(n7777), .ZN(n9182) );
  NAND2_X1 U9366 ( .A1(n10236), .A2(n7777), .ZN(n9929) );
  AND2_X1 U9367 ( .A1(n9182), .A2(n9929), .ZN(n9267) );
  NAND2_X1 U9368 ( .A1(n7778), .A2(n9472), .ZN(n7779) );
  XOR2_X1 U9369 ( .A(n9267), .B(n7807), .Z(n10235) );
  XOR2_X1 U9370 ( .A(n9267), .B(n7811), .Z(n7783) );
  OAI22_X1 U9371 ( .A1(n7781), .A2(n9751), .B1(n7816), .B2(n9769), .ZN(n7782)
         );
  AOI21_X1 U9372 ( .B1(n7783), .B2(n9772), .A(n7782), .ZN(n7784) );
  OAI21_X1 U9373 ( .B1(n10235), .B2(n9757), .A(n7784), .ZN(n10241) );
  NAND2_X1 U9374 ( .A1(n10241), .A2(n9774), .ZN(n7792) );
  OAI22_X1 U9375 ( .A1(n9774), .A2(n7786), .B1(n7785), .B2(n10187), .ZN(n7790)
         );
  AND2_X1 U9376 ( .A1(n7787), .A2(n10236), .ZN(n7788) );
  OR2_X1 U9377 ( .A1(n7788), .A2(n9952), .ZN(n10240) );
  NOR2_X1 U9378 ( .A1(n10240), .A2(n9550), .ZN(n7789) );
  AOI211_X1 U9379 ( .C1(n9947), .C2(n10236), .A(n7790), .B(n7789), .ZN(n7791)
         );
  OAI211_X1 U9380 ( .C1(n10235), .C2(n9782), .A(n7792), .B(n7791), .ZN(
        P1_U3282) );
  INV_X1 U9381 ( .A(n7794), .ZN(n7795) );
  AOI21_X1 U9382 ( .B1(n7796), .B2(n7793), .A(n7795), .ZN(n7802) );
  INV_X1 U9383 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7797) );
  NOR2_X1 U9384 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7797), .ZN(n10113) );
  INV_X1 U9385 ( .A(n9936), .ZN(n7812) );
  NOR2_X1 U9386 ( .A1(n7812), .A2(n9161), .ZN(n7798) );
  AOI211_X1 U9387 ( .C1(n10469), .C2(n9471), .A(n10113), .B(n7798), .ZN(n7799)
         );
  OAI21_X1 U9388 ( .B1(n9158), .B2(n7907), .A(n7799), .ZN(n7800) );
  AOI21_X1 U9389 ( .B1(n9996), .B2(n9165), .A(n7800), .ZN(n7801) );
  OAI21_X1 U9390 ( .B1(n7802), .B2(n9139), .A(n7801), .ZN(P1_U3222) );
  OAI222_X1 U9391 ( .A1(P2_U3152), .A2(n7805), .B1(n4481), .B2(n7804), .C1(
        n7803), .C2(n9050), .ZN(P2_U3334) );
  AND2_X1 U9392 ( .A1(n10236), .A2(n9937), .ZN(n7806) );
  NAND2_X1 U9393 ( .A1(n9948), .A2(n7816), .ZN(n9344) );
  NAND2_X1 U9394 ( .A1(n9351), .A2(n9344), .ZN(n9934) );
  NAND2_X1 U9395 ( .A1(n9928), .A2(n9934), .ZN(n7810) );
  OR2_X1 U9396 ( .A1(n9948), .A2(n7808), .ZN(n7809) );
  XNOR2_X1 U9397 ( .A(n7895), .B(n9936), .ZN(n9356) );
  INV_X1 U9398 ( .A(n9356), .ZN(n9271) );
  XNOR2_X1 U9399 ( .A(n7898), .B(n9271), .ZN(n10006) );
  NAND2_X1 U9400 ( .A1(n9351), .A2(n9182), .ZN(n9346) );
  NAND2_X1 U9401 ( .A1(n9344), .A2(n9929), .ZN(n9352) );
  NAND2_X1 U9402 ( .A1(n9352), .A2(n9351), .ZN(n9181) );
  OR2_X1 U9403 ( .A1(n7895), .A2(n7812), .ZN(n7937) );
  INV_X1 U9404 ( .A(n7937), .ZN(n7815) );
  AOI21_X1 U9405 ( .B1(n7813), .B2(n9271), .A(n9940), .ZN(n7814) );
  OAI21_X1 U9406 ( .B1(n7938), .B2(n7815), .A(n7814), .ZN(n7819) );
  OAI22_X1 U9407 ( .A1(n7816), .A2(n9751), .B1(n7899), .B2(n9769), .ZN(n7817)
         );
  INV_X1 U9408 ( .A(n7817), .ZN(n7818) );
  NAND2_X1 U9409 ( .A1(n7819), .A2(n7818), .ZN(n7820) );
  AOI21_X1 U9410 ( .B1(n10006), .B2(n9943), .A(n7820), .ZN(n10008) );
  INV_X1 U9411 ( .A(n9948), .ZN(n9959) );
  INV_X1 U9412 ( .A(n7895), .ZN(n10003) );
  OR2_X1 U9413 ( .A1(n9949), .A2(n10003), .ZN(n7821) );
  NAND2_X1 U9414 ( .A1(n7905), .A2(n7821), .ZN(n10004) );
  OAI22_X1 U9415 ( .A1(n9774), .A2(n7823), .B1(n7822), .B2(n10187), .ZN(n7824)
         );
  AOI21_X1 U9416 ( .B1(n7895), .B2(n9947), .A(n7824), .ZN(n7825) );
  OAI21_X1 U9417 ( .B1(n10004), .B2(n9550), .A(n7825), .ZN(n7826) );
  AOI21_X1 U9418 ( .B1(n10006), .B2(n9955), .A(n7826), .ZN(n7827) );
  OAI21_X1 U9419 ( .B1(n10008), .B2(n10193), .A(n7827), .ZN(P1_U3280) );
  INV_X1 U9420 ( .A(n7828), .ZN(n7830) );
  NAND2_X1 U9421 ( .A1(n7830), .A2(n7829), .ZN(n7831) );
  XNOR2_X1 U9422 ( .A(n7832), .B(n7831), .ZN(n7837) );
  AND2_X1 U9423 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10126) );
  NOR2_X1 U9424 ( .A1(n7899), .A2(n9161), .ZN(n7833) );
  AOI211_X1 U9425 ( .C1(n10469), .C2(n9767), .A(n10126), .B(n7833), .ZN(n7834)
         );
  OAI21_X1 U9426 ( .B1(n9158), .B2(n7946), .A(n7834), .ZN(n7835) );
  AOI21_X1 U9427 ( .B1(n9869), .B2(n9165), .A(n7835), .ZN(n7836) );
  OAI21_X1 U9428 ( .B1(n7837), .B2(n9139), .A(n7836), .ZN(P1_U3232) );
  XNOR2_X1 U9429 ( .A(n7839), .B(n7838), .ZN(n7843) );
  OAI22_X1 U9430 ( .A1(n8614), .A2(n8018), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7607), .ZN(n7841) );
  OAI22_X1 U9431 ( .A1(n8615), .A2(n7976), .B1(n7980), .B2(n8628), .ZN(n7840)
         );
  AOI211_X1 U9432 ( .C1(n8114), .C2(n8618), .A(n7841), .B(n7840), .ZN(n7842)
         );
  OAI21_X1 U9433 ( .B1(n7843), .B2(n8620), .A(n7842), .ZN(P2_U3236) );
  INV_X1 U9434 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10450) );
  NOR2_X1 U9435 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7844) );
  AOI21_X1 U9436 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7844), .ZN(n10416) );
  NOR2_X1 U9437 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7845) );
  AOI21_X1 U9438 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7845), .ZN(n10419) );
  NOR2_X1 U9439 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n7846) );
  AOI21_X1 U9440 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n7846), .ZN(n10422) );
  NOR2_X1 U9441 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7847) );
  AOI21_X1 U9442 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7847), .ZN(n10425) );
  NOR2_X1 U9443 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7848) );
  AOI21_X1 U9444 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7848), .ZN(n10428) );
  NOR2_X1 U9445 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7849) );
  AOI21_X1 U9446 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7849), .ZN(n10467) );
  NAND2_X1 U9447 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10409) );
  INV_X1 U9448 ( .A(n10409), .ZN(n10411) );
  INV_X1 U9449 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10408) );
  NAND2_X1 U9450 ( .A1(n10409), .A2(n10408), .ZN(n10407) );
  AOI22_X1 U9451 ( .A1(n10411), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(n10407), .ZN(n10443) );
  NAND2_X1 U9452 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7850) );
  OAI21_X1 U9453 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7850), .ZN(n10442) );
  NOR2_X1 U9454 ( .A1(n10443), .A2(n10442), .ZN(n10441) );
  AOI21_X1 U9455 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10441), .ZN(n10464) );
  NAND2_X1 U9456 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7851) );
  OAI21_X1 U9457 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7851), .ZN(n10463) );
  NOR2_X1 U9458 ( .A1(n10464), .A2(n10463), .ZN(n10462) );
  AOI21_X1 U9459 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10462), .ZN(n10466) );
  NAND2_X1 U9460 ( .A1(n10467), .A2(n10466), .ZN(n10465) );
  OAI21_X1 U9461 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10465), .ZN(n7852) );
  INV_X1 U9462 ( .A(n7852), .ZN(n7853) );
  NOR2_X1 U9463 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7853), .ZN(n10445) );
  INV_X1 U9464 ( .A(n10445), .ZN(n10446) );
  INV_X1 U9465 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10448) );
  NAND2_X1 U9466 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7853), .ZN(n10447) );
  NAND2_X1 U9467 ( .A1(n10448), .A2(n10447), .ZN(n10444) );
  NAND2_X1 U9468 ( .A1(n10446), .A2(n10444), .ZN(n7854) );
  INV_X1 U9469 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10080) );
  NOR2_X1 U9470 ( .A1(n7854), .A2(n10080), .ZN(n7855) );
  XNOR2_X1 U9471 ( .A(n7854), .B(n10080), .ZN(n10440) );
  INV_X1 U9472 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10439) );
  INV_X1 U9473 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n8148) );
  AOI22_X1 U9474 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n8148), .B1(
        P2_ADDR_REG_7__SCAN_IN), .B2(n8193), .ZN(n10457) );
  INV_X1 U9475 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n8309) );
  INV_X1 U9476 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10096) );
  AOI22_X1 U9477 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n8309), .B1(
        P2_ADDR_REG_8__SCAN_IN), .B2(n10096), .ZN(n10460) );
  AOI21_X1 U9478 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10459), .ZN(n7856) );
  INV_X1 U9479 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7857) );
  NOR2_X1 U9480 ( .A1(n7856), .A2(n7857), .ZN(n7858) );
  INV_X1 U9481 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10455) );
  XNOR2_X1 U9482 ( .A(n7857), .B(n7856), .ZN(n10454) );
  NAND2_X1 U9483 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7859) );
  OAI21_X1 U9484 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n7859), .ZN(n10436) );
  NAND2_X1 U9485 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7860) );
  OAI21_X1 U9486 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7860), .ZN(n10433) );
  AOI21_X1 U9487 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10432), .ZN(n10431) );
  NOR2_X1 U9488 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7861) );
  AOI21_X1 U9489 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7861), .ZN(n10430) );
  NAND2_X1 U9490 ( .A1(n10431), .A2(n10430), .ZN(n10429) );
  OAI21_X1 U9491 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10429), .ZN(n10427) );
  NAND2_X1 U9492 ( .A1(n10428), .A2(n10427), .ZN(n10426) );
  OAI21_X1 U9493 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10426), .ZN(n10424) );
  NAND2_X1 U9494 ( .A1(n10425), .A2(n10424), .ZN(n10423) );
  OAI21_X1 U9495 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10423), .ZN(n10421) );
  NAND2_X1 U9496 ( .A1(n10422), .A2(n10421), .ZN(n10420) );
  OAI21_X1 U9497 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10420), .ZN(n10418) );
  NAND2_X1 U9498 ( .A1(n10419), .A2(n10418), .ZN(n10417) );
  OAI21_X1 U9499 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10417), .ZN(n10415) );
  NAND2_X1 U9500 ( .A1(n10416), .A2(n10415), .ZN(n10414) );
  OAI21_X1 U9501 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10414), .ZN(n10451) );
  NOR2_X1 U9502 ( .A1(n10450), .A2(n10451), .ZN(n7862) );
  NAND2_X1 U9503 ( .A1(n10450), .A2(n10451), .ZN(n10449) );
  OAI21_X1 U9504 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7862), .A(n10449), .ZN(
        n7864) );
  XNOR2_X1 U9505 ( .A(n4890), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7863) );
  XNOR2_X1 U9506 ( .A(n7864), .B(n7863), .ZN(ADD_1071_U4) );
  OAI21_X1 U9507 ( .B1(n7867), .B2(n6128), .A(n8002), .ZN(n7871) );
  NOR2_X1 U9508 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6143), .ZN(n7868) );
  AOI21_X1 U9509 ( .B1(n10260), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7868), .ZN(
        n7869) );
  OAI21_X1 U9510 ( .B1(n10261), .B2(n8001), .A(n7869), .ZN(n7870) );
  AOI21_X1 U9511 ( .B1(n7871), .B2(n10259), .A(n7870), .ZN(n7876) );
  AOI21_X1 U9512 ( .B1(n7873), .B2(n6111), .A(n7872), .ZN(n7992) );
  XNOR2_X1 U9513 ( .A(n7992), .B(n8001), .ZN(n7874) );
  NAND2_X1 U9514 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7874), .ZN(n7994) );
  OAI211_X1 U9515 ( .C1(n7874), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10258), .B(
        n7994), .ZN(n7875) );
  NAND2_X1 U9516 ( .A1(n7876), .A2(n7875), .ZN(P2_U3260) );
  NAND2_X1 U9517 ( .A1(n7877), .A2(n8639), .ZN(n7878) );
  INV_X1 U9518 ( .A(n7887), .ZN(n7880) );
  OAI21_X1 U9519 ( .B1(n4568), .B2(n7880), .A(n7970), .ZN(n10392) );
  NAND2_X1 U9520 ( .A1(n7881), .A2(n10386), .ZN(n7882) );
  NAND2_X1 U9521 ( .A1(n7982), .A2(n7882), .ZN(n10389) );
  OAI22_X1 U9522 ( .A1(n8915), .A2(n7884), .B1(n7883), .B2(n8912), .ZN(n7885)
         );
  AOI21_X1 U9523 ( .B1(n10386), .B2(n10284), .A(n7885), .ZN(n7886) );
  OAI21_X1 U9524 ( .B1(n10389), .B2(n7984), .A(n7886), .ZN(n7893) );
  XNOR2_X1 U9525 ( .A(n7888), .B(n7887), .ZN(n7891) );
  OAI22_X1 U9526 ( .A1(n8115), .A2(n8886), .B1(n7889), .B2(n8884), .ZN(n7890)
         );
  AOI21_X1 U9527 ( .B1(n7891), .B2(n8933), .A(n7890), .ZN(n10388) );
  NOR2_X1 U9528 ( .A1(n10388), .A2(n10293), .ZN(n7892) );
  AOI211_X1 U9529 ( .C1(n10288), .C2(n10392), .A(n7893), .B(n7892), .ZN(n7894)
         );
  INV_X1 U9530 ( .A(n7894), .ZN(P2_U3284) );
  NOR2_X1 U9531 ( .A1(n7895), .A2(n9936), .ZN(n7897) );
  NAND2_X1 U9532 ( .A1(n7895), .A2(n9936), .ZN(n7896) );
  OR2_X1 U9533 ( .A1(n9996), .A2(n7899), .ZN(n9357) );
  NAND2_X1 U9534 ( .A1(n9996), .A2(n7899), .ZN(n9345) );
  NAND2_X1 U9535 ( .A1(n9357), .A2(n9345), .ZN(n9270) );
  INV_X1 U9536 ( .A(n9270), .ZN(n7900) );
  XNOR2_X1 U9537 ( .A(n7934), .B(n7900), .ZN(n10000) );
  NAND2_X1 U9538 ( .A1(n7938), .A2(n7937), .ZN(n7901) );
  XNOR2_X1 U9539 ( .A(n7901), .B(n7900), .ZN(n7903) );
  AOI22_X1 U9540 ( .A1(n9938), .A2(n9936), .B1(n9471), .B2(n9935), .ZN(n7902)
         );
  OAI21_X1 U9541 ( .B1(n7903), .B2(n9940), .A(n7902), .ZN(n7904) );
  AOI21_X1 U9542 ( .B1(n10000), .B2(n9943), .A(n7904), .ZN(n10002) );
  INV_X1 U9543 ( .A(n9950), .ZN(n10239) );
  AOI21_X1 U9544 ( .B1(n7905), .B2(n9996), .A(n10239), .ZN(n7906) );
  NAND2_X1 U9545 ( .A1(n7906), .A2(n7944), .ZN(n9997) );
  OAI22_X1 U9546 ( .A1(n9774), .A2(n7908), .B1(n7907), .B2(n10187), .ZN(n7909)
         );
  AOI21_X1 U9547 ( .B1(n9996), .B2(n9947), .A(n7909), .ZN(n7910) );
  OAI21_X1 U9548 ( .B1(n9997), .B2(n7911), .A(n7910), .ZN(n7912) );
  AOI21_X1 U9549 ( .B1(n10000), .B2(n9955), .A(n7912), .ZN(n7913) );
  OAI21_X1 U9550 ( .B1(n10002), .B2(n10193), .A(n7913), .ZN(P1_U3279) );
  INV_X1 U9551 ( .A(n7914), .ZN(n7918) );
  OAI222_X1 U9552 ( .A1(n7916), .A2(P2_U3152), .B1(n4481), .B2(n7918), .C1(
        n7915), .C2(n9050), .ZN(P2_U3333) );
  OAI222_X1 U9553 ( .A1(n9901), .A2(n7919), .B1(n4480), .B2(n7918), .C1(n7917), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9554 ( .A(n7920), .ZN(n7952) );
  OAI222_X1 U9555 ( .A1(n4480), .A2(n7952), .B1(P1_U3084), .B2(n7922), .C1(
        n7921), .C2(n9896), .ZN(P1_U3327) );
  INV_X1 U9556 ( .A(n7923), .ZN(n7924) );
  AOI21_X1 U9557 ( .B1(n7926), .B2(n7925), .A(n7924), .ZN(n7933) );
  OR2_X1 U9558 ( .A1(n8115), .A2(n8884), .ZN(n7928) );
  OR2_X1 U9559 ( .A1(n8576), .A2(n8886), .ZN(n7927) );
  NAND2_X1 U9560 ( .A1(n7928), .A2(n7927), .ZN(n9967) );
  NAND2_X1 U9561 ( .A1(n9967), .A2(n8631), .ZN(n7930) );
  OAI211_X1 U9562 ( .C1(n8628), .C2(n9970), .A(n7930), .B(n7929), .ZN(n7931)
         );
  AOI21_X1 U9563 ( .B1(n9972), .B2(n8618), .A(n7931), .ZN(n7932) );
  OAI21_X1 U9564 ( .B1(n7933), .B2(n8620), .A(n7932), .ZN(P2_U3217) );
  NAND2_X1 U9565 ( .A1(n7934), .A2(n9270), .ZN(n7936) );
  NAND2_X1 U9566 ( .A1(n9996), .A2(n7940), .ZN(n7935) );
  NAND2_X1 U9567 ( .A1(n7936), .A2(n7935), .ZN(n7956) );
  XNOR2_X1 U9568 ( .A(n9869), .B(n9471), .ZN(n9273) );
  XNOR2_X1 U9569 ( .A(n7956), .B(n9273), .ZN(n9872) );
  AND2_X1 U9570 ( .A1(n9357), .A2(n7937), .ZN(n9184) );
  NAND2_X1 U9571 ( .A1(n7939), .A2(n9345), .ZN(n7960) );
  XNOR2_X1 U9572 ( .A(n7960), .B(n4767), .ZN(n7942) );
  AOI22_X1 U9573 ( .A1(n7940), .A2(n9938), .B1(n9935), .B2(n9767), .ZN(n7941)
         );
  OAI21_X1 U9574 ( .B1(n7942), .B2(n9940), .A(n7941), .ZN(n7943) );
  AOI21_X1 U9575 ( .B1(n9872), .B2(n9943), .A(n7943), .ZN(n9874) );
  AND2_X1 U9576 ( .A1(n7944), .A2(n9869), .ZN(n7945) );
  OR2_X1 U9577 ( .A1(n7945), .A2(n7957), .ZN(n9870) );
  OAI22_X1 U9578 ( .A1(n9774), .A2(n7947), .B1(n7946), .B2(n10187), .ZN(n7948)
         );
  AOI21_X1 U9579 ( .B1(n9869), .B2(n9947), .A(n7948), .ZN(n7949) );
  OAI21_X1 U9580 ( .B1(n9870), .B2(n9550), .A(n7949), .ZN(n7950) );
  AOI21_X1 U9581 ( .B1(n9872), .B2(n9955), .A(n7950), .ZN(n7951) );
  OAI21_X1 U9582 ( .B1(n9874), .B2(n10193), .A(n7951), .ZN(P1_U3278) );
  OAI222_X1 U9583 ( .A1(P2_U3152), .A2(n7953), .B1(n4481), .B2(n7952), .C1(
        n8321), .C2(n9050), .ZN(P2_U3332) );
  AND2_X1 U9584 ( .A1(n9869), .A2(n9471), .ZN(n7955) );
  OR2_X1 U9585 ( .A1(n9869), .A2(n9471), .ZN(n7954) );
  NAND2_X1 U9586 ( .A1(n9864), .A2(n9162), .ZN(n9190) );
  XNOR2_X1 U9587 ( .A(n8064), .B(n9275), .ZN(n9867) );
  AOI211_X1 U9588 ( .C1(n9864), .C2(n4679), .A(n10239), .B(n9760), .ZN(n9863)
         );
  NOR2_X1 U9589 ( .A1(n9067), .A2(n9742), .ZN(n7959) );
  OAI22_X1 U9590 ( .A1(n9774), .A2(n5453), .B1(n9062), .B2(n10187), .ZN(n7958)
         );
  AOI211_X1 U9591 ( .C1(n9863), .C2(n9954), .A(n7959), .B(n7958), .ZN(n7965)
         );
  INV_X1 U9592 ( .A(n9471), .ZN(n9188) );
  OAI211_X1 U9593 ( .C1(n7961), .C2(n9275), .A(n9762), .B(n9772), .ZN(n7963)
         );
  INV_X1 U9594 ( .A(n9750), .ZN(n9470) );
  AOI22_X1 U9595 ( .A1(n9470), .A2(n9935), .B1(n9938), .B2(n9471), .ZN(n7962)
         );
  NAND2_X1 U9596 ( .A1(n7963), .A2(n7962), .ZN(n9862) );
  NAND2_X1 U9597 ( .A1(n9862), .A2(n9774), .ZN(n7964) );
  OAI211_X1 U9598 ( .C1(n9867), .C2(n9755), .A(n7965), .B(n7964), .ZN(P1_U3277) );
  NAND2_X1 U9599 ( .A1(n7989), .A2(n8014), .ZN(n7967) );
  OAI211_X1 U9600 ( .C1(n9901), .C2(n7968), .A(n7967), .B(n7966), .ZN(P1_U3326) );
  OR2_X1 U9601 ( .A1(n10386), .A2(n8638), .ZN(n7969) );
  NAND2_X1 U9602 ( .A1(n7972), .A2(n7971), .ZN(n7973) );
  NAND2_X1 U9603 ( .A1(n8116), .A2(n7973), .ZN(n9027) );
  XNOR2_X1 U9604 ( .A(n7975), .B(n7974), .ZN(n7979) );
  OAI22_X1 U9605 ( .A1(n8018), .A2(n8886), .B1(n7976), .B2(n8884), .ZN(n7978)
         );
  NOR2_X1 U9606 ( .A1(n9027), .A2(n8845), .ZN(n7977) );
  AOI211_X1 U9607 ( .C1(n8933), .C2(n7979), .A(n7978), .B(n7977), .ZN(n9026)
         );
  OR2_X1 U9608 ( .A1(n9026), .A2(n10293), .ZN(n7988) );
  OAI22_X1 U9609 ( .A1(n8915), .A2(n7981), .B1(n7980), .B2(n8912), .ZN(n7986)
         );
  AND2_X1 U9610 ( .A1(n7982), .A2(n8114), .ZN(n7983) );
  OR2_X1 U9611 ( .A1(n7983), .A2(n4561), .ZN(n9023) );
  NOR2_X1 U9612 ( .A1(n9023), .A2(n7984), .ZN(n7985) );
  AOI211_X1 U9613 ( .C1(n10284), .C2(n8114), .A(n7986), .B(n7985), .ZN(n7987)
         );
  OAI211_X1 U9614 ( .C1(n9027), .C2(n8862), .A(n7988), .B(n7987), .ZN(P2_U3283) );
  INV_X1 U9615 ( .A(n7989), .ZN(n7991) );
  OAI222_X1 U9616 ( .A1(P2_U3152), .A2(n8029), .B1(n4481), .B2(n7991), .C1(
        n7990), .C2(n9050), .ZN(P2_U3331) );
  XNOR2_X1 U9617 ( .A(n8652), .B(n8657), .ZN(n7997) );
  NAND2_X1 U9618 ( .A1(n7993), .A2(n7992), .ZN(n7995) );
  AND2_X1 U9619 ( .A1(n7995), .A2(n7994), .ZN(n7996) );
  NAND2_X1 U9620 ( .A1(n7996), .A2(n7997), .ZN(n8662) );
  OAI21_X1 U9621 ( .B1(n7997), .B2(n7996), .A(n8662), .ZN(n8008) );
  NAND2_X1 U9622 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8575) );
  INV_X1 U9623 ( .A(n8575), .ZN(n7998) );
  AOI21_X1 U9624 ( .B1(n10260), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7998), .ZN(
        n7999) );
  OAI21_X1 U9625 ( .B1(n10261), .B2(n8658), .A(n7999), .ZN(n8007) );
  NAND2_X1 U9626 ( .A1(n8001), .A2(n8000), .ZN(n8003) );
  INV_X1 U9627 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8914) );
  MUX2_X1 U9628 ( .A(n8914), .B(P2_REG2_REG_16__SCAN_IN), .S(n8652), .Z(n8004)
         );
  AOI211_X1 U9629 ( .C1(n8005), .C2(n8004), .A(n10263), .B(n8651), .ZN(n8006)
         );
  AOI211_X1 U9630 ( .C1(n10258), .C2(n8008), .A(n8007), .B(n8006), .ZN(n8009)
         );
  INV_X1 U9631 ( .A(n8009), .ZN(P2_U3261) );
  NAND2_X1 U9632 ( .A1(n8015), .A2(n8010), .ZN(n8012) );
  OAI211_X1 U9633 ( .C1(n9050), .C2(n8013), .A(n8012), .B(n8011), .ZN(P2_U3330) );
  NAND2_X1 U9634 ( .A1(n8015), .A2(n8014), .ZN(n8016) );
  OAI211_X1 U9635 ( .C1(n8017), .C2(n9896), .A(n8016), .B(n9459), .ZN(P1_U3325) );
  XNOR2_X1 U9636 ( .A(n8566), .B(n8567), .ZN(n8570) );
  XNOR2_X1 U9637 ( .A(n8570), .B(n8569), .ZN(n8022) );
  OAI22_X1 U9638 ( .A1(n8614), .A2(n8885), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6143), .ZN(n8020) );
  OAI22_X1 U9639 ( .A1(n8615), .A2(n8018), .B1(n8921), .B2(n8628), .ZN(n8019)
         );
  AOI211_X1 U9640 ( .C1(n9016), .C2(n8618), .A(n8020), .B(n8019), .ZN(n8021)
         );
  OAI21_X1 U9641 ( .B1(n8022), .B2(n8620), .A(n8021), .ZN(P2_U3243) );
  XNOR2_X1 U9642 ( .A(n8024), .B(n8023), .ZN(n8028) );
  OAI22_X1 U9643 ( .A1(n8614), .A2(n8887), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8665), .ZN(n8026) );
  OAI22_X1 U9644 ( .A1(n8615), .A2(n8885), .B1(n8894), .B2(n8628), .ZN(n8025)
         );
  AOI211_X1 U9645 ( .C1(n9005), .C2(n8618), .A(n8026), .B(n8025), .ZN(n8027)
         );
  OAI21_X1 U9646 ( .B1(n8028), .B2(n8620), .A(n8027), .ZN(P2_U3230) );
  INV_X1 U9647 ( .A(n9016), .ZN(n8925) );
  INV_X1 U9648 ( .A(n8994), .ZN(n8847) );
  INV_X1 U9649 ( .A(n8987), .ZN(n8835) );
  NAND2_X1 U9650 ( .A1(n8832), .A2(n8823), .ZN(n8803) );
  INV_X1 U9651 ( .A(n8716), .ZN(n8140) );
  NAND2_X1 U9652 ( .A1(n8939), .A2(n8936), .ZN(n8034) );
  INV_X1 U9653 ( .A(n8029), .ZN(n8030) );
  NAND2_X1 U9654 ( .A1(n8030), .A2(P2_B_REG_SCAN_IN), .ZN(n8031) );
  AND2_X1 U9655 ( .A1(n8930), .A2(n8031), .ZN(n8136) );
  NAND2_X1 U9656 ( .A1(n8032), .A2(n8136), .ZN(n8943) );
  NOR2_X1 U9657 ( .A1(n10293), .A2(n8943), .ZN(n8710) );
  AOI21_X1 U9658 ( .B1(n10293), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8710), .ZN(
        n8033) );
  OAI211_X1 U9659 ( .C1(n8924), .C2(n8941), .A(n8034), .B(n8033), .ZN(P2_U3265) );
  NAND2_X1 U9660 ( .A1(n8035), .A2(n8036), .ZN(n8038) );
  XNOR2_X1 U9661 ( .A(n8038), .B(n8037), .ZN(n8043) );
  AOI22_X1 U9662 ( .A1(n9165), .A2(n8039), .B1(n9134), .B2(n7153), .ZN(n8042)
         );
  AOI22_X1 U9663 ( .A1(n10469), .A2(n9478), .B1(n8040), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n8041) );
  OAI211_X1 U9664 ( .C1(n8043), .C2(n9139), .A(n8042), .B(n8041), .ZN(P1_U3220) );
  NAND2_X1 U9665 ( .A1(n8045), .A2(n8044), .ZN(n8046) );
  XOR2_X1 U9666 ( .A(n8047), .B(n8046), .Z(n8052) );
  INV_X1 U9667 ( .A(n9714), .ZN(n9681) );
  NAND2_X1 U9668 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9517) );
  OAI21_X1 U9669 ( .B1(n9681), .B2(n9117), .A(n9517), .ZN(n8048) );
  AOI21_X1 U9670 ( .B1(n9134), .B2(n9715), .A(n8048), .ZN(n8049) );
  OAI21_X1 U9671 ( .B1(n9158), .B2(n9717), .A(n8049), .ZN(n8050) );
  AOI21_X1 U9672 ( .B1(n9841), .B2(n9165), .A(n8050), .ZN(n8051) );
  OAI21_X1 U9673 ( .B1(n8052), .B2(n9139), .A(n8051), .ZN(P1_U3236) );
  INV_X1 U9674 ( .A(n8053), .ZN(n8055) );
  NOR2_X1 U9675 ( .A1(n8055), .A2(n8054), .ZN(n8056) );
  XNOR2_X1 U9676 ( .A(n8057), .B(n8056), .ZN(n8062) );
  INV_X1 U9677 ( .A(n9106), .ZN(n9731) );
  INV_X1 U9678 ( .A(n9701), .ZN(n9079) );
  NAND2_X1 U9679 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9537) );
  OAI21_X1 U9680 ( .B1(n9079), .B2(n9117), .A(n9537), .ZN(n8058) );
  AOI21_X1 U9681 ( .B1(n9134), .B2(n9731), .A(n8058), .ZN(n8059) );
  OAI21_X1 U9682 ( .B1(n9158), .B2(n9695), .A(n8059), .ZN(n8060) );
  AOI21_X1 U9683 ( .B1(n9836), .B2(n9165), .A(n8060), .ZN(n8061) );
  OAI21_X1 U9684 ( .B1(n8062), .B2(n9139), .A(n8061), .ZN(P1_U3217) );
  INV_X1 U9685 ( .A(n9654), .ZN(n8089) );
  INV_X1 U9686 ( .A(n9770), .ZN(n9730) );
  NOR2_X1 U9687 ( .A1(n9864), .A2(n9767), .ZN(n8063) );
  NOR2_X1 U9688 ( .A1(n9759), .A2(n9750), .ZN(n8065) );
  NAND2_X1 U9689 ( .A1(n9853), .A2(n9770), .ZN(n9377) );
  NOR2_X1 U9690 ( .A1(n9846), .A2(n9715), .ZN(n8066) );
  INV_X1 U9691 ( .A(n9715), .ZN(n9752) );
  INV_X1 U9692 ( .A(n9846), .ZN(n9727) );
  OAI22_X1 U9693 ( .A1(n9722), .A2(n8066), .B1(n9752), .B2(n9727), .ZN(n9707)
         );
  OR2_X1 U9694 ( .A1(n9841), .A2(n9106), .ZN(n9393) );
  NAND2_X1 U9695 ( .A1(n9841), .A2(n9106), .ZN(n9180) );
  NAND2_X1 U9696 ( .A1(n9393), .A2(n9180), .ZN(n9706) );
  INV_X1 U9697 ( .A(n9836), .ZN(n9698) );
  NAND2_X1 U9698 ( .A1(n9827), .A2(n9682), .ZN(n9401) );
  INV_X1 U9699 ( .A(n9682), .ZN(n9653) );
  NAND2_X1 U9700 ( .A1(n9821), .A2(n9666), .ZN(n8068) );
  INV_X1 U9701 ( .A(n9666), .ZN(n8087) );
  AOI22_X1 U9702 ( .A1(n9646), .A2(n8068), .B1(n8087), .B2(n4685), .ZN(n9630)
         );
  NAND2_X1 U9703 ( .A1(n9630), .A2(n8069), .ZN(n8070) );
  NAND2_X1 U9704 ( .A1(n9808), .A2(n9469), .ZN(n9414) );
  NAND2_X1 U9705 ( .A1(n9591), .A2(n9611), .ZN(n8071) );
  INV_X1 U9706 ( .A(n9611), .ZN(n9468) );
  NAND2_X1 U9707 ( .A1(n9796), .A2(n9557), .ZN(n9237) );
  AOI21_X1 U9708 ( .B1(n9570), .B2(n9579), .A(n5025), .ZN(n9553) );
  NAND2_X1 U9709 ( .A1(n9791), .A2(n9580), .ZN(n9238) );
  INV_X1 U9710 ( .A(n9791), .ZN(n9563) );
  NAND2_X1 U9711 ( .A1(n8485), .A2(n5368), .ZN(n8074) );
  OR2_X1 U9712 ( .A1(n9173), .A2(n9902), .ZN(n8073) );
  NAND2_X1 U9713 ( .A1(n9786), .A2(n9556), .ZN(n9432) );
  NAND2_X1 U9714 ( .A1(n9760), .A2(n9759), .ZN(n9758) );
  INV_X1 U9715 ( .A(n9827), .ZN(n8075) );
  INV_X1 U9716 ( .A(n9811), .ZN(n9621) );
  AOI21_X1 U9717 ( .B1(n9786), .B2(n9564), .A(n9544), .ZN(n9787) );
  INV_X1 U9718 ( .A(n8076), .ZN(n8077) );
  AOI22_X1 U9719 ( .A1(n10193), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8077), .B2(
        n9946), .ZN(n8078) );
  OAI21_X1 U9720 ( .B1(n4690), .B2(n9742), .A(n8078), .ZN(n8105) );
  OR2_X1 U9721 ( .A1(n9858), .A2(n9750), .ZN(n9374) );
  NAND2_X1 U9722 ( .A1(n9858), .A2(n9750), .ZN(n9373) );
  NAND2_X1 U9723 ( .A1(n9374), .A2(n9373), .ZN(n9763) );
  INV_X1 U9724 ( .A(n9761), .ZN(n8079) );
  NOR2_X1 U9725 ( .A1(n9763), .A2(n8079), .ZN(n8080) );
  INV_X1 U9726 ( .A(n9748), .ZN(n8081) );
  NOR2_X1 U9727 ( .A1(n9846), .A2(n9752), .ZN(n9255) );
  NAND2_X1 U9728 ( .A1(n9846), .A2(n9752), .ZN(n9253) );
  INV_X1 U9729 ( .A(n9706), .ZN(n9712) );
  OR2_X1 U9730 ( .A1(n9836), .A2(n9681), .ZN(n9392) );
  NAND2_X1 U9731 ( .A1(n9836), .A2(n9681), .ZN(n9396) );
  NAND2_X1 U9732 ( .A1(n9700), .A2(n9699), .ZN(n8083) );
  AND2_X1 U9733 ( .A1(n9833), .A2(n9079), .ZN(n9395) );
  NOR2_X1 U9734 ( .A1(n9660), .A2(n9398), .ZN(n8086) );
  NAND2_X1 U9735 ( .A1(n9662), .A2(n8086), .ZN(n9663) );
  NAND2_X1 U9736 ( .A1(n9663), .A2(n9401), .ZN(n9651) );
  NAND2_X1 U9737 ( .A1(n9651), .A2(n9404), .ZN(n8088) );
  NAND2_X1 U9738 ( .A1(n9821), .A2(n8087), .ZN(n9402) );
  NAND2_X1 U9739 ( .A1(n8088), .A2(n9402), .ZN(n9638) );
  NAND2_X1 U9740 ( .A1(n9816), .A2(n8089), .ZN(n9409) );
  INV_X1 U9741 ( .A(n9642), .ZN(n9612) );
  NAND2_X1 U9742 ( .A1(n9811), .A2(n9612), .ZN(n9410) );
  OR2_X1 U9743 ( .A1(n9811), .A2(n9612), .ZN(n9316) );
  NAND2_X1 U9744 ( .A1(n9316), .A2(n9622), .ZN(n9412) );
  NAND2_X1 U9745 ( .A1(n9412), .A2(n9410), .ZN(n9319) );
  INV_X1 U9746 ( .A(n9415), .ZN(n9235) );
  INV_X1 U9747 ( .A(n9577), .ZN(n9239) );
  NOR2_X1 U9748 ( .A1(n9579), .A2(n9239), .ZN(n8092) );
  INV_X1 U9749 ( .A(n9238), .ZN(n9424) );
  MUX2_X1 U9750 ( .A(n8093), .B(n9426), .S(n9434), .Z(n8096) );
  INV_X1 U9751 ( .A(n9555), .ZN(n8094) );
  NAND3_X1 U9752 ( .A1(n8094), .A2(n9238), .A3(n9434), .ZN(n8095) );
  NAND2_X1 U9753 ( .A1(n8096), .A2(n8095), .ZN(n8097) );
  NAND2_X1 U9754 ( .A1(n8098), .A2(P1_B_REG_SCAN_IN), .ZN(n8099) );
  AND2_X1 U9755 ( .A1(n9935), .A2(n8099), .ZN(n9539) );
  INV_X1 U9756 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9546) );
  NAND2_X1 U9757 ( .A1(n5755), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8103) );
  NAND2_X1 U9758 ( .A1(n8101), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8102) );
  OAI211_X1 U9759 ( .C1(n5806), .C2(n9546), .A(n8103), .B(n8102), .ZN(n9466)
         );
  AOI22_X1 U9760 ( .A1(n8072), .A2(n9938), .B1(n9539), .B2(n9466), .ZN(n8104)
         );
  OAI21_X1 U9761 ( .B1(n9790), .B2(n9755), .A(n8106), .ZN(P1_U3355) );
  AOI22_X1 U9762 ( .A1(n8618), .A2(n8107), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8537), .ZN(n8113) );
  OAI21_X1 U9763 ( .B1(n8109), .B2(n8108), .A(n10334), .ZN(n8110) );
  NAND3_X1 U9764 ( .A1(n8111), .A2(n8622), .A3(n8110), .ZN(n8112) );
  OAI211_X1 U9765 ( .C1(n6530), .C2(n8614), .A(n8113), .B(n8112), .ZN(P2_U3234) );
  INV_X1 U9766 ( .A(n8885), .ZN(n8931) );
  INV_X1 U9767 ( .A(n8114), .ZN(n9022) );
  INV_X1 U9768 ( .A(n8576), .ZN(n8902) );
  INV_X1 U9769 ( .A(n8869), .ZN(n8903) );
  INV_X1 U9770 ( .A(n4584), .ZN(n8875) );
  OR2_X1 U9771 ( .A1(n8994), .A2(n8867), .ZN(n8121) );
  NAND2_X1 U9772 ( .A1(n8844), .A2(n8121), .ZN(n8122) );
  NAND2_X1 U9773 ( .A1(n8122), .A2(n5022), .ZN(n8831) );
  INV_X1 U9774 ( .A(n8548), .ZN(n8853) );
  INV_X1 U9775 ( .A(n8812), .ZN(n8124) );
  NAND2_X1 U9776 ( .A1(n8982), .A2(n8124), .ZN(n8125) );
  NAND2_X1 U9777 ( .A1(n8819), .A2(n8125), .ZN(n8126) );
  INV_X1 U9778 ( .A(n8977), .ZN(n8807) );
  INV_X1 U9779 ( .A(n8972), .ZN(n8797) );
  INV_X1 U9780 ( .A(n8813), .ZN(n8127) );
  NAND2_X1 U9781 ( .A1(n8768), .A2(n8128), .ZN(n8753) );
  INV_X1 U9782 ( .A(n8557), .ZN(n8734) );
  NOR2_X1 U9783 ( .A1(n8946), .A2(n8735), .ZN(n8131) );
  XNOR2_X1 U9784 ( .A(n8132), .B(n8133), .ZN(n8722) );
  NAND2_X1 U9785 ( .A1(n8135), .A2(n8933), .ZN(n8138) );
  AOI22_X1 U9786 ( .A1(n8735), .A2(n8928), .B1(n8136), .B2(n8635), .ZN(n8137)
         );
  XNOR2_X1 U9787 ( .A(n8489), .B(n8716), .ZN(n8717) );
  NAND2_X1 U9788 ( .A1(n8717), .A2(n9978), .ZN(n8139) );
  NAND2_X1 U9789 ( .A1(n10393), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8141) );
  OAI21_X1 U9790 ( .B1(n8143), .B2(n10393), .A(n8141), .ZN(P2_U3517) );
  NOR2_X1 U9791 ( .A1(n10406), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8142) );
  INV_X1 U9792 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U9793 ( .A1(n10378), .A2(keyinput134), .B1(n7510), .B2(keyinput186), 
        .ZN(n8144) );
  OAI221_X1 U9794 ( .B1(n10378), .B2(keyinput134), .C1(n7510), .C2(keyinput186), .A(n8144), .ZN(n8152) );
  AOI22_X1 U9795 ( .A1(n9526), .A2(keyinput191), .B1(keyinput133), .B2(n6813), 
        .ZN(n8145) );
  OAI221_X1 U9796 ( .B1(n9526), .B2(keyinput191), .C1(n6813), .C2(keyinput133), 
        .A(n8145), .ZN(n8151) );
  AOI22_X1 U9797 ( .A1(n9172), .A2(keyinput185), .B1(n6811), .B2(keyinput144), 
        .ZN(n8146) );
  OAI221_X1 U9798 ( .B1(n9172), .B2(keyinput185), .C1(n6811), .C2(keyinput144), 
        .A(n8146), .ZN(n8150) );
  AOI22_X1 U9799 ( .A1(n10195), .A2(keyinput199), .B1(keyinput173), .B2(n8148), 
        .ZN(n8147) );
  OAI221_X1 U9800 ( .B1(n10195), .B2(keyinput199), .C1(n8148), .C2(keyinput173), .A(n8147), .ZN(n8149) );
  NOR4_X1 U9801 ( .A1(n8152), .A2(n8151), .A3(n8150), .A4(n8149), .ZN(n8167)
         );
  INV_X1 U9802 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8154) );
  AOI22_X1 U9803 ( .A1(n8154), .A2(keyinput155), .B1(n5351), .B2(keyinput203), 
        .ZN(n8153) );
  OAI221_X1 U9804 ( .B1(n8154), .B2(keyinput155), .C1(n5351), .C2(keyinput203), 
        .A(n8153), .ZN(n8159) );
  INV_X1 U9805 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8347) );
  AOI22_X1 U9806 ( .A1(n8328), .A2(keyinput204), .B1(keyinput247), .B2(n8347), 
        .ZN(n8155) );
  OAI221_X1 U9807 ( .B1(n8328), .B2(keyinput204), .C1(n8347), .C2(keyinput247), 
        .A(n8155), .ZN(n8158) );
  INV_X1 U9808 ( .A(SI_3_), .ZN(n8319) );
  INV_X1 U9809 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8339) );
  AOI22_X1 U9810 ( .A1(n8319), .A2(keyinput240), .B1(keyinput140), .B2(n8339), 
        .ZN(n8156) );
  OAI221_X1 U9811 ( .B1(n8319), .B2(keyinput240), .C1(n8339), .C2(keyinput140), 
        .A(n8156), .ZN(n8157) );
  NOR3_X1 U9812 ( .A1(n8159), .A2(n8158), .A3(n8157), .ZN(n8166) );
  AOI22_X1 U9813 ( .A1(n10202), .A2(keyinput244), .B1(keyinput213), .B2(n8914), 
        .ZN(n8160) );
  OAI221_X1 U9814 ( .B1(n10202), .B2(keyinput244), .C1(n8914), .C2(keyinput213), .A(n8160), .ZN(n8164) );
  AOI22_X1 U9815 ( .A1(n8162), .A2(keyinput189), .B1(keyinput238), .B2(n7981), 
        .ZN(n8161) );
  OAI221_X1 U9816 ( .B1(n8162), .B2(keyinput189), .C1(n7981), .C2(keyinput238), 
        .A(n8161), .ZN(n8163) );
  NOR2_X1 U9817 ( .A1(n8164), .A2(n8163), .ZN(n8165) );
  NAND3_X1 U9818 ( .A1(n8167), .A2(n8166), .A3(n8165), .ZN(n8285) );
  INV_X1 U9819 ( .A(SI_7_), .ZN(n8311) );
  AOI22_X1 U9820 ( .A1(n8311), .A2(keyinput148), .B1(keyinput223), .B2(n6975), 
        .ZN(n8168) );
  OAI221_X1 U9821 ( .B1(n8311), .B2(keyinput148), .C1(n6975), .C2(keyinput223), 
        .A(n8168), .ZN(n8177) );
  INV_X1 U9822 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8386) );
  AOI22_X1 U9823 ( .A1(n8386), .A2(keyinput222), .B1(n8170), .B2(keyinput241), 
        .ZN(n8169) );
  OAI221_X1 U9824 ( .B1(n8386), .B2(keyinput222), .C1(n8170), .C2(keyinput241), 
        .A(n8169), .ZN(n8176) );
  XNOR2_X1 U9825 ( .A(P1_REG1_REG_25__SCAN_IN), .B(keyinput215), .ZN(n8174) );
  XNOR2_X1 U9826 ( .A(P1_REG3_REG_27__SCAN_IN), .B(keyinput207), .ZN(n8173) );
  XNOR2_X1 U9827 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput254), .ZN(n8172) );
  XNOR2_X1 U9828 ( .A(P2_REG1_REG_16__SCAN_IN), .B(keyinput196), .ZN(n8171) );
  NAND4_X1 U9829 ( .A1(n8174), .A2(n8173), .A3(n8172), .A4(n8171), .ZN(n8175)
         );
  OR3_X1 U9830 ( .A1(n8177), .A2(n8176), .A3(n8175), .ZN(n8190) );
  INV_X1 U9831 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10394) );
  AOI22_X1 U9832 ( .A1(n8337), .A2(keyinput205), .B1(keyinput236), .B2(n10394), 
        .ZN(n8178) );
  OAI221_X1 U9833 ( .B1(n8337), .B2(keyinput205), .C1(n10394), .C2(keyinput236), .A(n8178), .ZN(n8189) );
  XNOR2_X1 U9834 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput201), .ZN(n8182) );
  XNOR2_X1 U9835 ( .A(P2_REG1_REG_13__SCAN_IN), .B(keyinput170), .ZN(n8181) );
  XNOR2_X1 U9836 ( .A(P1_REG1_REG_27__SCAN_IN), .B(keyinput184), .ZN(n8180) );
  XNOR2_X1 U9837 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput202), .ZN(n8179) );
  NAND4_X1 U9838 ( .A1(n8182), .A2(n8181), .A3(n8180), .A4(n8179), .ZN(n8188)
         );
  XNOR2_X1 U9839 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput164), .ZN(n8186) );
  XNOR2_X1 U9840 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput229), .ZN(n8185) );
  XNOR2_X1 U9841 ( .A(P2_REG0_REG_27__SCAN_IN), .B(keyinput129), .ZN(n8184) );
  XNOR2_X1 U9842 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput142), .ZN(n8183) );
  NAND4_X1 U9843 ( .A1(n8186), .A2(n8185), .A3(n8184), .A4(n8183), .ZN(n8187)
         );
  NOR4_X1 U9844 ( .A1(n8190), .A2(n8189), .A3(n8188), .A4(n8187), .ZN(n8209)
         );
  AOI22_X1 U9845 ( .A1(n6009), .A2(keyinput249), .B1(n8352), .B2(keyinput220), 
        .ZN(n8191) );
  OAI221_X1 U9846 ( .B1(n6009), .B2(keyinput249), .C1(n8352), .C2(keyinput220), 
        .A(n8191), .ZN(n8196) );
  AOI22_X1 U9847 ( .A1(n8193), .A2(keyinput153), .B1(keyinput214), .B2(n9546), 
        .ZN(n8192) );
  OAI221_X1 U9848 ( .B1(n8193), .B2(keyinput153), .C1(n9546), .C2(keyinput214), 
        .A(n8192), .ZN(n8195) );
  XNOR2_X1 U9849 ( .A(n10200), .B(keyinput230), .ZN(n8194) );
  NOR3_X1 U9850 ( .A1(n8196), .A2(n8195), .A3(n8194), .ZN(n8208) );
  INV_X1 U9851 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10146) );
  XOR2_X1 U9852 ( .A(keyinput139), .B(n10146), .Z(n8207) );
  AOI22_X1 U9853 ( .A1(n8198), .A2(keyinput135), .B1(n5983), .B2(keyinput180), 
        .ZN(n8197) );
  OAI221_X1 U9854 ( .B1(n8198), .B2(keyinput135), .C1(n5983), .C2(keyinput180), 
        .A(n8197), .ZN(n8205) );
  AOI22_X1 U9855 ( .A1(n8201), .A2(keyinput194), .B1(n8200), .B2(keyinput163), 
        .ZN(n8199) );
  OAI221_X1 U9856 ( .B1(n8201), .B2(keyinput194), .C1(n8200), .C2(keyinput163), 
        .A(n8199), .ZN(n8204) );
  XOR2_X1 U9857 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput245), .Z(n8203) );
  XOR2_X1 U9858 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput248), .Z(n8202) );
  NOR4_X1 U9859 ( .A1(n8205), .A2(n8204), .A3(n8203), .A4(n8202), .ZN(n8206)
         );
  NAND4_X1 U9860 ( .A1(n8209), .A2(n8208), .A3(n8207), .A4(n8206), .ZN(n8284)
         );
  AOI22_X1 U9861 ( .A1(P2_D_REG_25__SCAN_IN), .A2(keyinput179), .B1(
        P1_D_REG_17__SCAN_IN), .B2(keyinput174), .ZN(n8210) );
  OAI221_X1 U9862 ( .B1(P2_D_REG_25__SCAN_IN), .B2(keyinput179), .C1(
        P1_D_REG_17__SCAN_IN), .C2(keyinput174), .A(n8210), .ZN(n8217) );
  AOI22_X1 U9863 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(keyinput239), .B1(
        P1_IR_REG_22__SCAN_IN), .B2(keyinput217), .ZN(n8211) );
  OAI221_X1 U9864 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(keyinput239), .C1(
        P1_IR_REG_22__SCAN_IN), .C2(keyinput217), .A(n8211), .ZN(n8216) );
  AOI22_X1 U9865 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(keyinput167), .B1(
        P1_REG2_REG_26__SCAN_IN), .B2(keyinput145), .ZN(n8212) );
  OAI221_X1 U9866 ( .B1(P2_IR_REG_29__SCAN_IN), .B2(keyinput167), .C1(
        P1_REG2_REG_26__SCAN_IN), .C2(keyinput145), .A(n8212), .ZN(n8215) );
  AOI22_X1 U9867 ( .A1(P2_REG0_REG_26__SCAN_IN), .A2(keyinput165), .B1(
        P1_REG2_REG_23__SCAN_IN), .B2(keyinput210), .ZN(n8213) );
  OAI221_X1 U9868 ( .B1(P2_REG0_REG_26__SCAN_IN), .B2(keyinput165), .C1(
        P1_REG2_REG_23__SCAN_IN), .C2(keyinput210), .A(n8213), .ZN(n8214) );
  NOR4_X1 U9869 ( .A1(n8217), .A2(n8216), .A3(n8215), .A4(n8214), .ZN(n8245)
         );
  AOI22_X1 U9870 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(keyinput156), .B1(
        P1_D_REG_31__SCAN_IN), .B2(keyinput146), .ZN(n8218) );
  OAI221_X1 U9871 ( .B1(P1_DATAO_REG_26__SCAN_IN), .B2(keyinput156), .C1(
        P1_D_REG_31__SCAN_IN), .C2(keyinput146), .A(n8218), .ZN(n8225) );
  AOI22_X1 U9872 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(keyinput211), .B1(
        P1_REG1_REG_19__SCAN_IN), .B2(keyinput171), .ZN(n8219) );
  OAI221_X1 U9873 ( .B1(P2_IR_REG_2__SCAN_IN), .B2(keyinput211), .C1(
        P1_REG1_REG_19__SCAN_IN), .C2(keyinput171), .A(n8219), .ZN(n8224) );
  AOI22_X1 U9874 ( .A1(P2_D_REG_26__SCAN_IN), .A2(keyinput252), .B1(
        P1_REG3_REG_4__SCAN_IN), .B2(keyinput195), .ZN(n8220) );
  OAI221_X1 U9875 ( .B1(P2_D_REG_26__SCAN_IN), .B2(keyinput252), .C1(
        P1_REG3_REG_4__SCAN_IN), .C2(keyinput195), .A(n8220), .ZN(n8223) );
  AOI22_X1 U9876 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(keyinput188), .B1(
        P1_REG0_REG_19__SCAN_IN), .B2(keyinput177), .ZN(n8221) );
  OAI221_X1 U9877 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(keyinput188), .C1(
        P1_REG0_REG_19__SCAN_IN), .C2(keyinput177), .A(n8221), .ZN(n8222) );
  NOR4_X1 U9878 ( .A1(n8225), .A2(n8224), .A3(n8223), .A4(n8222), .ZN(n8244)
         );
  AOI22_X1 U9879 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(keyinput183), .B1(SI_13_), 
        .B2(keyinput228), .ZN(n8226) );
  OAI221_X1 U9880 ( .B1(P1_DATAO_REG_3__SCAN_IN), .B2(keyinput183), .C1(SI_13_), .C2(keyinput228), .A(n8226), .ZN(n8233) );
  AOI22_X1 U9881 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(keyinput209), .B1(
        P2_D_REG_15__SCAN_IN), .B2(keyinput143), .ZN(n8227) );
  OAI221_X1 U9882 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(keyinput209), .C1(
        P2_D_REG_15__SCAN_IN), .C2(keyinput143), .A(n8227), .ZN(n8232) );
  AOI22_X1 U9883 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput242), .B1(
        P2_D_REG_7__SCAN_IN), .B2(keyinput224), .ZN(n8228) );
  OAI221_X1 U9884 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput242), .C1(
        P2_D_REG_7__SCAN_IN), .C2(keyinput224), .A(n8228), .ZN(n8231) );
  AOI22_X1 U9885 ( .A1(P2_REG1_REG_29__SCAN_IN), .A2(keyinput166), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(keyinput161), .ZN(n8229) );
  OAI221_X1 U9886 ( .B1(P2_REG1_REG_29__SCAN_IN), .B2(keyinput166), .C1(
        P1_DATAO_REG_2__SCAN_IN), .C2(keyinput161), .A(n8229), .ZN(n8230) );
  NOR4_X1 U9887 ( .A1(n8233), .A2(n8232), .A3(n8231), .A4(n8230), .ZN(n8243)
         );
  AOI22_X1 U9888 ( .A1(P2_REG0_REG_24__SCAN_IN), .A2(keyinput206), .B1(
        P2_REG0_REG_16__SCAN_IN), .B2(keyinput226), .ZN(n8234) );
  OAI221_X1 U9889 ( .B1(P2_REG0_REG_24__SCAN_IN), .B2(keyinput206), .C1(
        P2_REG0_REG_16__SCAN_IN), .C2(keyinput226), .A(n8234), .ZN(n8241) );
  AOI22_X1 U9890 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(keyinput219), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput227), .ZN(n8235) );
  OAI221_X1 U9891 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(keyinput219), .C1(
        P1_IR_REG_7__SCAN_IN), .C2(keyinput227), .A(n8235), .ZN(n8240) );
  AOI22_X1 U9892 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput152), .B1(
        P2_REG3_REG_25__SCAN_IN), .B2(keyinput225), .ZN(n8236) );
  OAI221_X1 U9893 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput152), .C1(
        P2_REG3_REG_25__SCAN_IN), .C2(keyinput225), .A(n8236), .ZN(n8239) );
  AOI22_X1 U9894 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput147), .B1(
        P2_D_REG_3__SCAN_IN), .B2(keyinput168), .ZN(n8237) );
  OAI221_X1 U9895 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput147), .C1(
        P2_D_REG_3__SCAN_IN), .C2(keyinput168), .A(n8237), .ZN(n8238) );
  NOR4_X1 U9896 ( .A1(n8241), .A2(n8240), .A3(n8239), .A4(n8238), .ZN(n8242)
         );
  NAND4_X1 U9897 ( .A1(n8245), .A2(n8244), .A3(n8243), .A4(n8242), .ZN(n8283)
         );
  AOI22_X1 U9898 ( .A1(P1_REG0_REG_5__SCAN_IN), .A2(keyinput232), .B1(
        P1_REG3_REG_17__SCAN_IN), .B2(keyinput208), .ZN(n8246) );
  OAI221_X1 U9899 ( .B1(P1_REG0_REG_5__SCAN_IN), .B2(keyinput232), .C1(
        P1_REG3_REG_17__SCAN_IN), .C2(keyinput208), .A(n8246), .ZN(n8253) );
  AOI22_X1 U9900 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(keyinput160), .B1(
        P1_REG3_REG_15__SCAN_IN), .B2(keyinput159), .ZN(n8247) );
  OAI221_X1 U9901 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(keyinput160), .C1(
        P1_REG3_REG_15__SCAN_IN), .C2(keyinput159), .A(n8247), .ZN(n8252) );
  AOI22_X1 U9902 ( .A1(P2_REG2_REG_7__SCAN_IN), .A2(keyinput157), .B1(
        P2_D_REG_29__SCAN_IN), .B2(keyinput154), .ZN(n8248) );
  OAI221_X1 U9903 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(keyinput157), .C1(
        P2_D_REG_29__SCAN_IN), .C2(keyinput154), .A(n8248), .ZN(n8251) );
  AOI22_X1 U9904 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(keyinput172), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(keyinput235), .ZN(n8249) );
  OAI221_X1 U9905 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(keyinput172), .C1(
        P2_DATAO_REG_6__SCAN_IN), .C2(keyinput235), .A(n8249), .ZN(n8250) );
  NOR4_X1 U9906 ( .A1(n8253), .A2(n8252), .A3(n8251), .A4(n8250), .ZN(n8281)
         );
  AOI22_X1 U9907 ( .A1(P2_REG0_REG_14__SCAN_IN), .A2(keyinput212), .B1(
        P1_IR_REG_31__SCAN_IN), .B2(keyinput138), .ZN(n8254) );
  OAI221_X1 U9908 ( .B1(P2_REG0_REG_14__SCAN_IN), .B2(keyinput212), .C1(
        P1_IR_REG_31__SCAN_IN), .C2(keyinput138), .A(n8254), .ZN(n8261) );
  AOI22_X1 U9909 ( .A1(P2_REG2_REG_29__SCAN_IN), .A2(keyinput253), .B1(
        P1_REG0_REG_11__SCAN_IN), .B2(keyinput221), .ZN(n8255) );
  OAI221_X1 U9910 ( .B1(P2_REG2_REG_29__SCAN_IN), .B2(keyinput253), .C1(
        P1_REG0_REG_11__SCAN_IN), .C2(keyinput221), .A(n8255), .ZN(n8260) );
  AOI22_X1 U9911 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(keyinput197), .B1(
        P1_REG1_REG_7__SCAN_IN), .B2(keyinput182), .ZN(n8256) );
  OAI221_X1 U9912 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(keyinput197), .C1(
        P1_REG1_REG_7__SCAN_IN), .C2(keyinput182), .A(n8256), .ZN(n8259) );
  AOI22_X1 U9913 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput169), .B1(
        P1_REG2_REG_19__SCAN_IN), .B2(keyinput251), .ZN(n8257) );
  OAI221_X1 U9914 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput169), .C1(
        P1_REG2_REG_19__SCAN_IN), .C2(keyinput251), .A(n8257), .ZN(n8258) );
  NOR4_X1 U9915 ( .A1(n8261), .A2(n8260), .A3(n8259), .A4(n8258), .ZN(n8280)
         );
  AOI22_X1 U9916 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput193), .B1(
        P2_IR_REG_1__SCAN_IN), .B2(keyinput162), .ZN(n8262) );
  OAI221_X1 U9917 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput193), .C1(
        P2_IR_REG_1__SCAN_IN), .C2(keyinput162), .A(n8262), .ZN(n8269) );
  AOI22_X1 U9918 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(keyinput158), .B1(
        P1_D_REG_23__SCAN_IN), .B2(keyinput131), .ZN(n8263) );
  OAI221_X1 U9919 ( .B1(P2_IR_REG_23__SCAN_IN), .B2(keyinput158), .C1(
        P1_D_REG_23__SCAN_IN), .C2(keyinput131), .A(n8263), .ZN(n8268) );
  AOI22_X1 U9920 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(keyinput237), .B1(
        P1_D_REG_28__SCAN_IN), .B2(keyinput200), .ZN(n8264) );
  OAI221_X1 U9921 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(keyinput237), .C1(
        P1_D_REG_28__SCAN_IN), .C2(keyinput200), .A(n8264), .ZN(n8267) );
  AOI22_X1 U9922 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(keyinput218), .B1(
        P1_IR_REG_17__SCAN_IN), .B2(keyinput141), .ZN(n8265) );
  OAI221_X1 U9923 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(keyinput218), .C1(
        P1_IR_REG_17__SCAN_IN), .C2(keyinput141), .A(n8265), .ZN(n8266) );
  NOR4_X1 U9924 ( .A1(n8269), .A2(n8268), .A3(n8267), .A4(n8266), .ZN(n8279)
         );
  AOI22_X1 U9925 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(keyinput255), .B1(
        P1_REG3_REG_24__SCAN_IN), .B2(keyinput151), .ZN(n8270) );
  OAI221_X1 U9926 ( .B1(P2_REG2_REG_28__SCAN_IN), .B2(keyinput255), .C1(
        P1_REG3_REG_24__SCAN_IN), .C2(keyinput151), .A(n8270), .ZN(n8277) );
  AOI22_X1 U9927 ( .A1(P2_D_REG_0__SCAN_IN), .A2(keyinput250), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(keyinput246), .ZN(n8271) );
  OAI221_X1 U9928 ( .B1(P2_D_REG_0__SCAN_IN), .B2(keyinput250), .C1(
        P1_REG2_REG_1__SCAN_IN), .C2(keyinput246), .A(n8271), .ZN(n8276) );
  AOI22_X1 U9929 ( .A1(P2_REG0_REG_13__SCAN_IN), .A2(keyinput178), .B1(
        P2_IR_REG_20__SCAN_IN), .B2(keyinput216), .ZN(n8272) );
  OAI221_X1 U9930 ( .B1(P2_REG0_REG_13__SCAN_IN), .B2(keyinput178), .C1(
        P2_IR_REG_20__SCAN_IN), .C2(keyinput216), .A(n8272), .ZN(n8275) );
  AOI22_X1 U9931 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(keyinput149), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(keyinput137), .ZN(n8273) );
  OAI221_X1 U9932 ( .B1(P1_DATAO_REG_11__SCAN_IN), .B2(keyinput149), .C1(
        P2_DATAO_REG_19__SCAN_IN), .C2(keyinput137), .A(n8273), .ZN(n8274) );
  NOR4_X1 U9933 ( .A1(n8277), .A2(n8276), .A3(n8275), .A4(n8274), .ZN(n8278)
         );
  NAND4_X1 U9934 ( .A1(n8281), .A2(n8280), .A3(n8279), .A4(n8278), .ZN(n8282)
         );
  NOR4_X1 U9935 ( .A1(n8285), .A2(n8284), .A3(n8283), .A4(n8282), .ZN(n8306)
         );
  INV_X1 U9936 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10197) );
  AOI22_X1 U9937 ( .A1(n5376), .A2(keyinput128), .B1(n10197), .B2(keyinput181), 
        .ZN(n8286) );
  OAI221_X1 U9938 ( .B1(n5376), .B2(keyinput128), .C1(n10197), .C2(keyinput181), .A(n8286), .ZN(n8295) );
  AOI22_X1 U9939 ( .A1(n6873), .A2(keyinput234), .B1(n8288), .B2(keyinput243), 
        .ZN(n8287) );
  OAI221_X1 U9940 ( .B1(n6873), .B2(keyinput234), .C1(n8288), .C2(keyinput243), 
        .A(n8287), .ZN(n8294) );
  AOI22_X1 U9941 ( .A1(n8290), .A2(keyinput231), .B1(keyinput175), .B2(n6257), 
        .ZN(n8289) );
  OAI221_X1 U9942 ( .B1(n8290), .B2(keyinput231), .C1(n6257), .C2(keyinput175), 
        .A(n8289), .ZN(n8293) );
  AOI22_X1 U9943 ( .A1(n10299), .A2(keyinput136), .B1(keyinput190), .B2(n8665), 
        .ZN(n8291) );
  OAI221_X1 U9944 ( .B1(n10299), .B2(keyinput136), .C1(n8665), .C2(keyinput190), .A(n8291), .ZN(n8292) );
  NOR4_X1 U9945 ( .A1(n8295), .A2(n8294), .A3(n8293), .A4(n8292), .ZN(n8305)
         );
  AOI22_X1 U9946 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(keyinput192), .B1(
        P1_IR_REG_13__SCAN_IN), .B2(keyinput150), .ZN(n8296) );
  OAI221_X1 U9947 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(keyinput192), .C1(
        P1_IR_REG_13__SCAN_IN), .C2(keyinput150), .A(n8296), .ZN(n8303) );
  AOI22_X1 U9948 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(keyinput132), .B1(
        P1_REG1_REG_5__SCAN_IN), .B2(keyinput187), .ZN(n8297) );
  OAI221_X1 U9949 ( .B1(P2_IR_REG_19__SCAN_IN), .B2(keyinput132), .C1(
        P1_REG1_REG_5__SCAN_IN), .C2(keyinput187), .A(n8297), .ZN(n8302) );
  AOI22_X1 U9950 ( .A1(P2_REG0_REG_18__SCAN_IN), .A2(keyinput233), .B1(
        P1_IR_REG_21__SCAN_IN), .B2(keyinput198), .ZN(n8298) );
  OAI221_X1 U9951 ( .B1(P2_REG0_REG_18__SCAN_IN), .B2(keyinput233), .C1(
        P1_IR_REG_21__SCAN_IN), .C2(keyinput198), .A(n8298), .ZN(n8301) );
  AOI22_X1 U9952 ( .A1(n6122), .A2(keyinput130), .B1(n8388), .B2(keyinput176), 
        .ZN(n8299) );
  OAI221_X1 U9953 ( .B1(n6122), .B2(keyinput130), .C1(n8388), .C2(keyinput176), 
        .A(n8299), .ZN(n8300) );
  NOR4_X1 U9954 ( .A1(n8303), .A2(n8302), .A3(n8301), .A4(n8300), .ZN(n8304)
         );
  NAND3_X1 U9955 ( .A1(n8306), .A2(n8305), .A3(n8304), .ZN(n8482) );
  INV_X1 U9956 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10194) );
  AOI22_X1 U9957 ( .A1(n10194), .A2(keyinput18), .B1(keyinput60), .B2(n6894), 
        .ZN(n8307) );
  OAI221_X1 U9958 ( .B1(n10194), .B2(keyinput18), .C1(n6894), .C2(keyinput60), 
        .A(n8307), .ZN(n8317) );
  AOI22_X1 U9959 ( .A1(n5904), .A2(keyinput4), .B1(keyinput64), .B2(n8309), 
        .ZN(n8308) );
  OAI221_X1 U9960 ( .B1(n5904), .B2(keyinput4), .C1(n8309), .C2(keyinput64), 
        .A(n8308), .ZN(n8316) );
  AOI22_X1 U9961 ( .A1(n8312), .A2(keyinput21), .B1(keyinput20), .B2(n8311), 
        .ZN(n8310) );
  OAI221_X1 U9962 ( .B1(n8312), .B2(keyinput21), .C1(n8311), .C2(keyinput20), 
        .A(n8310), .ZN(n8315) );
  AOI22_X1 U9963 ( .A1(n5097), .A2(keyinput70), .B1(keyinput59), .B2(n5204), 
        .ZN(n8313) );
  OAI221_X1 U9964 ( .B1(n5097), .B2(keyinput70), .C1(n5204), .C2(keyinput59), 
        .A(n8313), .ZN(n8314) );
  NOR4_X1 U9965 ( .A1(n8317), .A2(n8316), .A3(n8315), .A4(n8314), .ZN(n8406)
         );
  AOI22_X1 U9966 ( .A1(n6811), .A2(keyinput16), .B1(n8319), .B2(keyinput112), 
        .ZN(n8318) );
  OAI221_X1 U9967 ( .B1(n6811), .B2(keyinput16), .C1(n8319), .C2(keyinput112), 
        .A(n8318), .ZN(n8325) );
  INV_X1 U9968 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8322) );
  AOI22_X1 U9969 ( .A1(n8322), .A2(keyinput90), .B1(n8321), .B2(keyinput28), 
        .ZN(n8320) );
  OAI221_X1 U9970 ( .B1(n8322), .B2(keyinput90), .C1(n8321), .C2(keyinput28), 
        .A(n8320), .ZN(n8324) );
  INV_X1 U9971 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10325) );
  XNOR2_X1 U9972 ( .A(n10325), .B(keyinput40), .ZN(n8323) );
  NOR3_X1 U9973 ( .A1(n8325), .A2(n8324), .A3(n8323), .ZN(n8344) );
  AOI22_X1 U9974 ( .A1(n10282), .A2(keyinput19), .B1(n7607), .B2(keyinput41), 
        .ZN(n8326) );
  OAI221_X1 U9975 ( .B1(n10282), .B2(keyinput19), .C1(n7607), .C2(keyinput41), 
        .A(n8326), .ZN(n8335) );
  AOI22_X1 U9976 ( .A1(n8329), .A2(keyinput98), .B1(n8328), .B2(keyinput76), 
        .ZN(n8327) );
  OAI221_X1 U9977 ( .B1(n8329), .B2(keyinput98), .C1(n8328), .C2(keyinput76), 
        .A(n8327), .ZN(n8334) );
  AOI22_X1 U9978 ( .A1(n8332), .A2(keyinput55), .B1(n8331), .B2(keyinput100), 
        .ZN(n8330) );
  OAI221_X1 U9979 ( .B1(n8332), .B2(keyinput55), .C1(n8331), .C2(keyinput100), 
        .A(n8330), .ZN(n8333) );
  NOR3_X1 U9980 ( .A1(n8335), .A2(n8334), .A3(n8333), .ZN(n8343) );
  INV_X1 U9981 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U9982 ( .A1(n8337), .A2(keyinput77), .B1(n10196), .B2(keyinput72), 
        .ZN(n8336) );
  OAI221_X1 U9983 ( .B1(n8337), .B2(keyinput77), .C1(n10196), .C2(keyinput72), 
        .A(n8336), .ZN(n8341) );
  INV_X1 U9984 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10198) );
  AOI22_X1 U9985 ( .A1(n8339), .A2(keyinput12), .B1(n10198), .B2(keyinput3), 
        .ZN(n8338) );
  OAI221_X1 U9986 ( .B1(n8339), .B2(keyinput12), .C1(n10198), .C2(keyinput3), 
        .A(n8338), .ZN(n8340) );
  NOR2_X1 U9987 ( .A1(n8341), .A2(n8340), .ZN(n8342) );
  NAND3_X1 U9988 ( .A1(n8344), .A2(n8343), .A3(n8342), .ZN(n8382) );
  AOI22_X1 U9989 ( .A1(n10096), .A2(keyinput69), .B1(n6975), .B2(keyinput95), 
        .ZN(n8345) );
  OAI221_X1 U9990 ( .B1(n10096), .B2(keyinput69), .C1(n6975), .C2(keyinput95), 
        .A(n8345), .ZN(n8349) );
  AOI22_X1 U9991 ( .A1(n8347), .A2(keyinput119), .B1(keyinput108), .B2(n10394), 
        .ZN(n8346) );
  OAI221_X1 U9992 ( .B1(n8347), .B2(keyinput119), .C1(n10394), .C2(keyinput108), .A(n8346), .ZN(n8348) );
  NOR2_X1 U9993 ( .A1(n8349), .A2(n8348), .ZN(n8380) );
  AOI22_X1 U9994 ( .A1(n5937), .A2(keyinput34), .B1(n5351), .B2(keyinput75), 
        .ZN(n8350) );
  OAI221_X1 U9995 ( .B1(n5937), .B2(keyinput34), .C1(n5351), .C2(keyinput75), 
        .A(n8350), .ZN(n8354) );
  AOI22_X1 U9996 ( .A1(n8352), .A2(keyinput92), .B1(keyinput29), .B2(n6912), 
        .ZN(n8351) );
  OAI221_X1 U9997 ( .B1(n8352), .B2(keyinput92), .C1(n6912), .C2(keyinput29), 
        .A(n8351), .ZN(n8353) );
  NOR2_X1 U9998 ( .A1(n8354), .A2(n8353), .ZN(n8379) );
  AOI22_X1 U9999 ( .A1(n8561), .A2(keyinput97), .B1(n10197), .B2(keyinput53), 
        .ZN(n8355) );
  OAI221_X1 U10000 ( .B1(n8561), .B2(keyinput97), .C1(n10197), .C2(keyinput53), 
        .A(n8355), .ZN(n8358) );
  INV_X1 U10001 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U10002 ( .A1(n10413), .A2(keyinput81), .B1(n6128), .B2(keyinput32), 
        .ZN(n8356) );
  OAI221_X1 U10003 ( .B1(n10413), .B2(keyinput81), .C1(n6128), .C2(keyinput32), 
        .A(n8356), .ZN(n8357) );
  NOR2_X1 U10004 ( .A1(n8358), .A2(n8357), .ZN(n8378) );
  AOI22_X1 U10005 ( .A1(n8657), .A2(keyinput68), .B1(keyinput86), .B2(n9546), 
        .ZN(n8359) );
  OAI221_X1 U10006 ( .B1(n8657), .B2(keyinput68), .C1(n9546), .C2(keyinput86), 
        .A(n8359), .ZN(n8360) );
  INV_X1 U10007 ( .A(n8360), .ZN(n8376) );
  XNOR2_X1 U10008 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput14), .ZN(n8363) );
  XNOR2_X1 U10009 ( .A(P1_REG1_REG_18__SCAN_IN), .B(keyinput63), .ZN(n8362) );
  XNOR2_X1 U10010 ( .A(keyinput2), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8361) );
  AND3_X1 U10011 ( .A1(n8363), .A2(n8362), .A3(n8361), .ZN(n8375) );
  XNOR2_X1 U10012 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput36), .ZN(n8367) );
  XNOR2_X1 U10013 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput22), .ZN(n8366) );
  XNOR2_X1 U10014 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput33), .ZN(n8365) );
  XNOR2_X1 U10015 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput109), .ZN(n8364)
         );
  NAND4_X1 U10016 ( .A1(n8367), .A2(n8366), .A3(n8365), .A4(n8364), .ZN(n8373)
         );
  XNOR2_X1 U10017 ( .A(keyinput118), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n8371) );
  XNOR2_X1 U10018 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput126), .ZN(n8370)
         );
  XNOR2_X1 U10019 ( .A(keyinput6), .B(P2_REG0_REG_10__SCAN_IN), .ZN(n8369) );
  XNOR2_X1 U10020 ( .A(keyinput85), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8368) );
  NAND4_X1 U10021 ( .A1(n8371), .A2(n8370), .A3(n8369), .A4(n8368), .ZN(n8372)
         );
  NOR2_X1 U10022 ( .A1(n8373), .A2(n8372), .ZN(n8374) );
  AND3_X1 U10023 ( .A1(n8376), .A2(n8375), .A3(n8374), .ZN(n8377) );
  NAND4_X1 U10024 ( .A1(n8380), .A2(n8379), .A3(n8378), .A4(n8377), .ZN(n8381)
         );
  NOR2_X1 U10025 ( .A1(n8382), .A2(n8381), .ZN(n8405) );
  AOI22_X1 U10026 ( .A1(n5947), .A2(keyinput83), .B1(n5375), .B2(keyinput93), 
        .ZN(n8383) );
  OAI221_X1 U10027 ( .B1(n5947), .B2(keyinput83), .C1(n5375), .C2(keyinput93), 
        .A(n8383), .ZN(n8393) );
  AOI22_X1 U10028 ( .A1(n5584), .A2(keyinput123), .B1(keyinput91), .B2(n5453), 
        .ZN(n8384) );
  OAI221_X1 U10029 ( .B1(n5584), .B2(keyinput123), .C1(n5453), .C2(keyinput91), 
        .A(n8384), .ZN(n8392) );
  AOI22_X1 U10030 ( .A1(n8386), .A2(keyinput94), .B1(n5687), .B2(keyinput82), 
        .ZN(n8385) );
  OAI221_X1 U10031 ( .B1(n8386), .B2(keyinput94), .C1(n5687), .C2(keyinput82), 
        .A(n8385), .ZN(n8391) );
  AOI22_X1 U10032 ( .A1(n8389), .A2(keyinput56), .B1(n8388), .B2(keyinput48), 
        .ZN(n8387) );
  OAI221_X1 U10033 ( .B1(n8389), .B2(keyinput56), .C1(n8388), .C2(keyinput48), 
        .A(n8387), .ZN(n8390) );
  NOR4_X1 U10034 ( .A1(n8393), .A2(n8392), .A3(n8391), .A4(n8390), .ZN(n8404)
         );
  AOI22_X1 U10035 ( .A1(P2_REG2_REG_26__SCAN_IN), .A2(keyinput47), .B1(
        P1_REG3_REG_15__SCAN_IN), .B2(keyinput31), .ZN(n8394) );
  OAI221_X1 U10036 ( .B1(P2_REG2_REG_26__SCAN_IN), .B2(keyinput47), .C1(
        P1_REG3_REG_15__SCAN_IN), .C2(keyinput31), .A(n8394), .ZN(n8402) );
  AOI22_X1 U10037 ( .A1(P2_REG0_REG_18__SCAN_IN), .A2(keyinput105), .B1(
        P2_D_REG_26__SCAN_IN), .B2(keyinput124), .ZN(n8395) );
  OAI221_X1 U10038 ( .B1(P2_REG0_REG_18__SCAN_IN), .B2(keyinput105), .C1(
        P2_D_REG_26__SCAN_IN), .C2(keyinput124), .A(n8395), .ZN(n8401) );
  AOI22_X1 U10039 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(keyinput42), .B1(
        P1_REG2_REG_4__SCAN_IN), .B2(keyinput5), .ZN(n8396) );
  OAI221_X1 U10040 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(keyinput42), .C1(
        P1_REG2_REG_4__SCAN_IN), .C2(keyinput5), .A(n8396), .ZN(n8400) );
  AOI22_X1 U10041 ( .A1(P2_REG0_REG_14__SCAN_IN), .A2(keyinput84), .B1(n8398), 
        .B2(keyinput80), .ZN(n8397) );
  OAI221_X1 U10042 ( .B1(P2_REG0_REG_14__SCAN_IN), .B2(keyinput84), .C1(n8398), 
        .C2(keyinput80), .A(n8397), .ZN(n8399) );
  NOR4_X1 U10043 ( .A1(n8402), .A2(n8401), .A3(n8400), .A4(n8399), .ZN(n8403)
         );
  AND4_X1 U10044 ( .A1(n8406), .A2(n8405), .A3(n8404), .A4(n8403), .ZN(n8481)
         );
  OAI22_X1 U10045 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(keyinput0), .B1(
        keyinput7), .B2(P2_REG1_REG_30__SCAN_IN), .ZN(n8407) );
  AOI221_X1 U10046 ( .B1(P1_REG3_REG_11__SCAN_IN), .B2(keyinput0), .C1(
        P2_REG1_REG_30__SCAN_IN), .C2(keyinput7), .A(n8407), .ZN(n8414) );
  OAI22_X1 U10047 ( .A1(P1_D_REG_10__SCAN_IN), .A2(keyinput102), .B1(
        P2_ADDR_REG_10__SCAN_IN), .B2(keyinput27), .ZN(n8408) );
  AOI221_X1 U10048 ( .B1(P1_D_REG_10__SCAN_IN), .B2(keyinput102), .C1(
        keyinput27), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n8408), .ZN(n8413) );
  OAI22_X1 U10049 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput89), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput115), .ZN(n8409) );
  AOI221_X1 U10050 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput89), .C1(
        keyinput115), .C2(P2_DATAO_REG_13__SCAN_IN), .A(n8409), .ZN(n8412) );
  OAI22_X1 U10051 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput103), .B1(
        P2_REG2_REG_13__SCAN_IN), .B2(keyinput110), .ZN(n8410) );
  AOI221_X1 U10052 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput103), .C1(
        keyinput110), .C2(P2_REG2_REG_13__SCAN_IN), .A(n8410), .ZN(n8411) );
  NAND4_X1 U10053 ( .A1(n8414), .A2(n8413), .A3(n8412), .A4(n8411), .ZN(n8442)
         );
  OAI22_X1 U10054 ( .A1(P1_REG2_REG_26__SCAN_IN), .A2(keyinput17), .B1(
        P2_ADDR_REG_7__SCAN_IN), .B2(keyinput45), .ZN(n8415) );
  AOI221_X1 U10055 ( .B1(P1_REG2_REG_26__SCAN_IN), .B2(keyinput17), .C1(
        keyinput45), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n8415), .ZN(n8422) );
  OAI22_X1 U10056 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput10), .B1(
        P1_ADDR_REG_7__SCAN_IN), .B2(keyinput25), .ZN(n8416) );
  AOI221_X1 U10057 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput10), .C1(
        keyinput25), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n8416), .ZN(n8421) );
  OAI22_X1 U10058 ( .A1(P1_REG1_REG_25__SCAN_IN), .A2(keyinput87), .B1(
        keyinput1), .B2(P2_REG0_REG_27__SCAN_IN), .ZN(n8417) );
  AOI221_X1 U10059 ( .B1(P1_REG1_REG_25__SCAN_IN), .B2(keyinput87), .C1(
        P2_REG0_REG_27__SCAN_IN), .C2(keyinput1), .A(n8417), .ZN(n8420) );
  OAI22_X1 U10060 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(keyinput73), .B1(
        P1_REG1_REG_8__SCAN_IN), .B2(keyinput106), .ZN(n8418) );
  AOI221_X1 U10061 ( .B1(P2_DATAO_REG_2__SCAN_IN), .B2(keyinput73), .C1(
        keyinput106), .C2(P1_REG1_REG_8__SCAN_IN), .A(n8418), .ZN(n8419) );
  NAND4_X1 U10062 ( .A1(n8422), .A2(n8421), .A3(n8420), .A4(n8419), .ZN(n8441)
         );
  OAI22_X1 U10063 ( .A1(P2_D_REG_28__SCAN_IN), .A2(keyinput8), .B1(keyinput38), 
        .B2(P2_REG1_REG_29__SCAN_IN), .ZN(n8423) );
  AOI221_X1 U10064 ( .B1(P2_D_REG_28__SCAN_IN), .B2(keyinput8), .C1(
        P2_REG1_REG_29__SCAN_IN), .C2(keyinput38), .A(n8423), .ZN(n8430) );
  OAI22_X1 U10065 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(keyinput117), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(keyinput24), .ZN(n8424) );
  AOI221_X1 U10066 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(keyinput117), .C1(
        keyinput24), .C2(P2_REG3_REG_12__SCAN_IN), .A(n8424), .ZN(n8429) );
  OAI22_X1 U10067 ( .A1(P1_REG0_REG_19__SCAN_IN), .A2(keyinput49), .B1(
        keyinput37), .B2(P2_REG0_REG_26__SCAN_IN), .ZN(n8425) );
  AOI221_X1 U10068 ( .B1(P1_REG0_REG_19__SCAN_IN), .B2(keyinput49), .C1(
        P2_REG0_REG_26__SCAN_IN), .C2(keyinput37), .A(n8425), .ZN(n8428) );
  OAI22_X1 U10069 ( .A1(P1_REG0_REG_5__SCAN_IN), .A2(keyinput104), .B1(
        keyinput125), .B2(P2_REG2_REG_29__SCAN_IN), .ZN(n8426) );
  AOI221_X1 U10070 ( .B1(P1_REG0_REG_5__SCAN_IN), .B2(keyinput104), .C1(
        P2_REG2_REG_29__SCAN_IN), .C2(keyinput125), .A(n8426), .ZN(n8427) );
  NAND4_X1 U10071 ( .A1(n8430), .A2(n8429), .A3(n8428), .A4(n8427), .ZN(n8440)
         );
  OAI22_X1 U10072 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput13), .B1(
        P2_IR_REG_9__SCAN_IN), .B2(keyinput120), .ZN(n8431) );
  AOI221_X1 U10073 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput13), .C1(
        keyinput120), .C2(P2_IR_REG_9__SCAN_IN), .A(n8431), .ZN(n8438) );
  OAI22_X1 U10074 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput99), .B1(
        P2_REG0_REG_13__SCAN_IN), .B2(keyinput50), .ZN(n8432) );
  AOI221_X1 U10075 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput99), .C1(
        keyinput50), .C2(P2_REG0_REG_13__SCAN_IN), .A(n8432), .ZN(n8437) );
  OAI22_X1 U10076 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(keyinput79), .B1(
        keyinput51), .B2(P2_D_REG_25__SCAN_IN), .ZN(n8433) );
  AOI221_X1 U10077 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(keyinput79), .C1(
        P2_D_REG_25__SCAN_IN), .C2(keyinput51), .A(n8433), .ZN(n8436) );
  OAI22_X1 U10078 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(keyinput30), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(keyinput11), .ZN(n8434) );
  AOI221_X1 U10079 ( .B1(P2_IR_REG_23__SCAN_IN), .B2(keyinput30), .C1(
        keyinput11), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n8434), .ZN(n8435) );
  NAND4_X1 U10080 ( .A1(n8438), .A2(n8437), .A3(n8436), .A4(n8435), .ZN(n8439)
         );
  NOR4_X1 U10081 ( .A1(n8442), .A2(n8441), .A3(n8440), .A4(n8439), .ZN(n8480)
         );
  OAI22_X1 U10082 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput121), .B1(
        keyinput127), .B2(P2_REG2_REG_28__SCAN_IN), .ZN(n8443) );
  AOI221_X1 U10083 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput121), .C1(
        P2_REG2_REG_28__SCAN_IN), .C2(keyinput127), .A(n8443), .ZN(n8450) );
  OAI22_X1 U10084 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(keyinput61), .B1(
        keyinput107), .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8444) );
  AOI221_X1 U10085 ( .B1(P2_DATAO_REG_21__SCAN_IN), .B2(keyinput61), .C1(
        P2_DATAO_REG_6__SCAN_IN), .C2(keyinput107), .A(n8444), .ZN(n8449) );
  OAI22_X1 U10086 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(keyinput88), .B1(
        keyinput96), .B2(P2_D_REG_7__SCAN_IN), .ZN(n8445) );
  AOI221_X1 U10087 ( .B1(P2_IR_REG_20__SCAN_IN), .B2(keyinput88), .C1(
        P2_D_REG_7__SCAN_IN), .C2(keyinput96), .A(n8445), .ZN(n8448) );
  OAI22_X1 U10088 ( .A1(P2_D_REG_15__SCAN_IN), .A2(keyinput15), .B1(
        P2_D_REG_0__SCAN_IN), .B2(keyinput122), .ZN(n8446) );
  AOI221_X1 U10089 ( .B1(P2_D_REG_15__SCAN_IN), .B2(keyinput15), .C1(
        keyinput122), .C2(P2_D_REG_0__SCAN_IN), .A(n8446), .ZN(n8447) );
  NAND4_X1 U10090 ( .A1(n8450), .A2(n8449), .A3(n8448), .A4(n8447), .ZN(n8478)
         );
  OAI22_X1 U10091 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(keyinput101), .B1(
        keyinput52), .B2(P2_REG0_REG_5__SCAN_IN), .ZN(n8451) );
  AOI221_X1 U10092 ( .B1(P2_IR_REG_7__SCAN_IN), .B2(keyinput101), .C1(
        P2_REG0_REG_5__SCAN_IN), .C2(keyinput52), .A(n8451), .ZN(n8458) );
  OAI22_X1 U10093 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(keyinput67), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(keyinput65), .ZN(n8452) );
  AOI221_X1 U10094 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(keyinput67), .C1(
        keyinput65), .C2(P2_DATAO_REG_31__SCAN_IN), .A(n8452), .ZN(n8457) );
  OAI22_X1 U10095 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput74), .B1(
        keyinput23), .B2(P1_REG3_REG_24__SCAN_IN), .ZN(n8453) );
  AOI221_X1 U10096 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput74), .C1(
        P1_REG3_REG_24__SCAN_IN), .C2(keyinput23), .A(n8453), .ZN(n8456) );
  OAI22_X1 U10097 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput116), .B1(
        keyinput114), .B2(P2_REG3_REG_16__SCAN_IN), .ZN(n8454) );
  AOI221_X1 U10098 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput116), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput114), .A(n8454), .ZN(n8455) );
  NAND4_X1 U10099 ( .A1(n8458), .A2(n8457), .A3(n8456), .A4(n8455), .ZN(n8477)
         );
  OAI22_X1 U10100 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(keyinput58), .B1(
        keyinput54), .B2(P1_REG1_REG_7__SCAN_IN), .ZN(n8459) );
  AOI221_X1 U10101 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(keyinput58), .C1(
        P1_REG1_REG_7__SCAN_IN), .C2(keyinput54), .A(n8459), .ZN(n8466) );
  OAI22_X1 U10102 ( .A1(P1_D_REG_30__SCAN_IN), .A2(keyinput71), .B1(
        P2_IR_REG_29__SCAN_IN), .B2(keyinput39), .ZN(n8460) );
  AOI221_X1 U10103 ( .B1(P1_D_REG_30__SCAN_IN), .B2(keyinput71), .C1(
        keyinput39), .C2(P2_IR_REG_29__SCAN_IN), .A(n8460), .ZN(n8465) );
  OAI22_X1 U10104 ( .A1(P1_D_REG_17__SCAN_IN), .A2(keyinput46), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(keyinput57), .ZN(n8461) );
  AOI221_X1 U10105 ( .B1(P1_D_REG_17__SCAN_IN), .B2(keyinput46), .C1(
        keyinput57), .C2(P2_DATAO_REG_30__SCAN_IN), .A(n8461), .ZN(n8464) );
  OAI22_X1 U10106 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput62), .B1(
        P2_REG0_REG_29__SCAN_IN), .B2(keyinput66), .ZN(n8462) );
  AOI221_X1 U10107 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput62), .C1(
        keyinput66), .C2(P2_REG0_REG_29__SCAN_IN), .A(n8462), .ZN(n8463) );
  NAND4_X1 U10108 ( .A1(n8466), .A2(n8465), .A3(n8464), .A4(n8463), .ZN(n8476)
         );
  OAI22_X1 U10109 ( .A1(P1_REG1_REG_19__SCAN_IN), .A2(keyinput43), .B1(
        P2_REG1_REG_17__SCAN_IN), .B2(keyinput111), .ZN(n8467) );
  AOI221_X1 U10110 ( .B1(P1_REG1_REG_19__SCAN_IN), .B2(keyinput43), .C1(
        keyinput111), .C2(P2_REG1_REG_17__SCAN_IN), .A(n8467), .ZN(n8474) );
  OAI22_X1 U10111 ( .A1(P2_REG0_REG_23__SCAN_IN), .A2(keyinput35), .B1(
        keyinput78), .B2(P2_REG0_REG_24__SCAN_IN), .ZN(n8468) );
  AOI221_X1 U10112 ( .B1(P2_REG0_REG_23__SCAN_IN), .B2(keyinput35), .C1(
        P2_REG0_REG_24__SCAN_IN), .C2(keyinput78), .A(n8468), .ZN(n8473) );
  OAI22_X1 U10113 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(keyinput9), .B1(
        keyinput113), .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8469) );
  AOI221_X1 U10114 ( .B1(P2_DATAO_REG_19__SCAN_IN), .B2(keyinput9), .C1(
        P2_DATAO_REG_10__SCAN_IN), .C2(keyinput113), .A(n8469), .ZN(n8472) );
  OAI22_X1 U10115 ( .A1(P2_D_REG_29__SCAN_IN), .A2(keyinput26), .B1(keyinput44), .B2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8470) );
  AOI221_X1 U10116 ( .B1(P2_D_REG_29__SCAN_IN), .B2(keyinput26), .C1(
        P2_ADDR_REG_14__SCAN_IN), .C2(keyinput44), .A(n8470), .ZN(n8471) );
  NAND4_X1 U10117 ( .A1(n8474), .A2(n8473), .A3(n8472), .A4(n8471), .ZN(n8475)
         );
  NOR4_X1 U10118 ( .A1(n8478), .A2(n8477), .A3(n8476), .A4(n8475), .ZN(n8479)
         );
  NAND4_X1 U10119 ( .A1(n8482), .A2(n8481), .A3(n8480), .A4(n8479), .ZN(n8483)
         );
  XNOR2_X1 U10120 ( .A(n8484), .B(n8483), .ZN(P2_U3549) );
  INV_X1 U10121 ( .A(n8485), .ZN(n9904) );
  OAI222_X1 U10122 ( .A1(P2_U3152), .A2(n8487), .B1(n4481), .B2(n9904), .C1(
        n8486), .C2(n9050), .ZN(P2_U3329) );
  XOR2_X1 U10123 ( .A(n8488), .B(n8493), .Z(n8950) );
  AOI21_X1 U10124 ( .B1(n8946), .B2(n8725), .A(n8489), .ZN(n8947) );
  AOI22_X1 U10125 ( .A1(n8490), .A2(n10283), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n10293), .ZN(n8491) );
  OAI21_X1 U10126 ( .B1(n8492), .B2(n8924), .A(n8491), .ZN(n8498) );
  XNOR2_X1 U10127 ( .A(n8494), .B(n8493), .ZN(n8496) );
  INV_X1 U10128 ( .A(n8495), .ZN(n8636) );
  AOI222_X1 U10129 ( .A1(n8933), .A2(n8496), .B1(n8636), .B2(n8930), .C1(n8637), .C2(n8928), .ZN(n8949) );
  NOR2_X1 U10130 ( .A1(n8949), .A2(n10293), .ZN(n8497) );
  AOI211_X1 U10131 ( .C1(n8936), .C2(n8947), .A(n8498), .B(n8497), .ZN(n8499)
         );
  OAI21_X1 U10132 ( .B1(n8950), .B2(n8938), .A(n8499), .ZN(P2_U3268) );
  INV_X1 U10133 ( .A(n9171), .ZN(n9052) );
  OAI222_X1 U10134 ( .A1(n4480), .A2(n9052), .B1(n8500), .B2(P1_U3084), .C1(
        n9172), .C2(n9901), .ZN(P1_U3323) );
  OAI211_X1 U10135 ( .C1(n8503), .C2(n8502), .A(n8501), .B(n8622), .ZN(n8509)
         );
  INV_X1 U10136 ( .A(n8614), .ZN(n8540) );
  INV_X1 U10137 ( .A(n8504), .ZN(n8727) );
  AOI22_X1 U10138 ( .A1(n8727), .A2(n8505), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8506) );
  OAI21_X1 U10139 ( .B1(n8557), .B2(n8615), .A(n8506), .ZN(n8507) );
  AOI21_X1 U10140 ( .B1(n8735), .B2(n8540), .A(n8507), .ZN(n8508) );
  OAI211_X1 U10141 ( .C1(n8729), .C2(n8634), .A(n8509), .B(n8508), .ZN(
        P2_U3216) );
  XNOR2_X1 U10142 ( .A(n8510), .B(n8582), .ZN(n8517) );
  OAI22_X1 U10143 ( .A1(n8512), .A2(n8614), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8511), .ZN(n8515) );
  INV_X1 U10144 ( .A(n8795), .ZN(n8513) );
  OAI22_X1 U10145 ( .A1(n8615), .A2(n8547), .B1(n8513), .B2(n8628), .ZN(n8514)
         );
  AOI211_X1 U10146 ( .C1(n8972), .C2(n8618), .A(n8515), .B(n8514), .ZN(n8516)
         );
  OAI21_X1 U10147 ( .B1(n8517), .B2(n8620), .A(n8516), .ZN(P2_U3218) );
  OAI211_X1 U10148 ( .C1(n8520), .C2(n8519), .A(n8518), .B(n8622), .ZN(n8524)
         );
  AOI22_X1 U10149 ( .A1(n8521), .A2(n8631), .B1(n8618), .B2(n10285), .ZN(n8523) );
  MUX2_X1 U10150 ( .A(n8628), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n8522) );
  NAND3_X1 U10151 ( .A1(n8524), .A2(n8523), .A3(n8522), .ZN(P2_U3220) );
  INV_X1 U10152 ( .A(n8525), .ZN(n8526) );
  AOI21_X1 U10153 ( .B1(n8528), .B2(n8527), .A(n8526), .ZN(n8532) );
  NAND2_X1 U10154 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8704) );
  OAI21_X1 U10155 ( .B1(n8614), .B2(n8548), .A(n8704), .ZN(n8530) );
  OAI22_X1 U10156 ( .A1(n8615), .A2(n8887), .B1(n8857), .B2(n8628), .ZN(n8529)
         );
  AOI211_X1 U10157 ( .C1(n8994), .C2(n8618), .A(n8530), .B(n8529), .ZN(n8531)
         );
  OAI21_X1 U10158 ( .B1(n8532), .B2(n8620), .A(n8531), .ZN(P2_U3221) );
  OAI21_X1 U10159 ( .B1(n8535), .B2(n8534), .A(n8533), .ZN(n8536) );
  NAND2_X1 U10160 ( .A1(n8536), .A2(n8622), .ZN(n8543) );
  AOI22_X1 U10161 ( .A1(n8618), .A2(n8538), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8537), .ZN(n8542) );
  AOI22_X1 U10162 ( .A1(n8540), .A2(n8648), .B1(n8539), .B2(n8650), .ZN(n8541)
         );
  NAND3_X1 U10163 ( .A1(n8543), .A2(n8542), .A3(n8541), .ZN(P2_U3224) );
  XNOR2_X1 U10164 ( .A(n8545), .B(n8544), .ZN(n8552) );
  OAI22_X1 U10165 ( .A1(n8547), .A2(n8614), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8546), .ZN(n8550) );
  OAI22_X1 U10166 ( .A1(n8615), .A2(n8548), .B1(n8820), .B2(n8628), .ZN(n8549)
         );
  AOI211_X1 U10167 ( .C1(n8982), .C2(n8618), .A(n8550), .B(n8549), .ZN(n8551)
         );
  OAI21_X1 U10168 ( .B1(n8552), .B2(n8620), .A(n8551), .ZN(P2_U3225) );
  XNOR2_X1 U10169 ( .A(n8554), .B(n8553), .ZN(n8555) );
  XNOR2_X1 U10170 ( .A(n8556), .B(n8555), .ZN(n8565) );
  OR2_X1 U10171 ( .A1(n8557), .A2(n8886), .ZN(n8559) );
  NAND2_X1 U10172 ( .A1(n8789), .A2(n8928), .ZN(n8558) );
  AND2_X1 U10173 ( .A1(n8559), .A2(n8558), .ZN(n8758) );
  NOR2_X1 U10174 ( .A1(n8758), .A2(n8560), .ZN(n8563) );
  OAI22_X1 U10175 ( .A1(n8761), .A2(n8628), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8561), .ZN(n8562) );
  AOI211_X1 U10176 ( .C1(n8963), .C2(n8618), .A(n8563), .B(n8562), .ZN(n8564)
         );
  OAI21_X1 U10177 ( .B1(n8565), .B2(n8620), .A(n8564), .ZN(P2_U3227) );
  INV_X1 U10178 ( .A(n8566), .ZN(n8568) );
  AOI22_X1 U10179 ( .A1(n8570), .A2(n8569), .B1(n8568), .B2(n8567), .ZN(n8574)
         );
  NAND2_X1 U10180 ( .A1(n8572), .A2(n8571), .ZN(n8573) );
  XNOR2_X1 U10181 ( .A(n8574), .B(n8573), .ZN(n8580) );
  OAI21_X1 U10182 ( .B1(n8614), .B2(n8869), .A(n8575), .ZN(n8578) );
  OAI22_X1 U10183 ( .A1(n8615), .A2(n8576), .B1(n8913), .B2(n8628), .ZN(n8577)
         );
  AOI211_X1 U10184 ( .C1(n9010), .C2(n8618), .A(n8578), .B(n8577), .ZN(n8579)
         );
  OAI21_X1 U10185 ( .B1(n8580), .B2(n8620), .A(n8579), .ZN(P2_U3228) );
  OAI21_X1 U10186 ( .B1(n8510), .B2(n8582), .A(n8581), .ZN(n8586) );
  XNOR2_X1 U10187 ( .A(n8584), .B(n8583), .ZN(n8585) );
  XNOR2_X1 U10188 ( .A(n8586), .B(n8585), .ZN(n8591) );
  OAI22_X1 U10189 ( .A1(n8813), .A2(n8615), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8587), .ZN(n8589) );
  OAI22_X1 U10190 ( .A1(n8777), .A2(n8614), .B1(n8628), .B2(n8781), .ZN(n8588)
         );
  AOI211_X1 U10191 ( .C1(n8966), .C2(n8618), .A(n8589), .B(n8588), .ZN(n8590)
         );
  OAI21_X1 U10192 ( .B1(n8591), .B2(n8620), .A(n8590), .ZN(P2_U3231) );
  XNOR2_X1 U10193 ( .A(n8593), .B(n8592), .ZN(n8599) );
  OAI22_X1 U10194 ( .A1(n8812), .A2(n8614), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8594), .ZN(n8597) );
  INV_X1 U10195 ( .A(n8833), .ZN(n8595) );
  OAI22_X1 U10196 ( .A1(n8615), .A2(n8613), .B1(n8595), .B2(n8628), .ZN(n8596)
         );
  AOI211_X1 U10197 ( .C1(n8987), .C2(n8618), .A(n8597), .B(n8596), .ZN(n8598)
         );
  OAI21_X1 U10198 ( .B1(n8599), .B2(n8620), .A(n8598), .ZN(P2_U3235) );
  OAI21_X1 U10199 ( .B1(n8602), .B2(n8601), .A(n8600), .ZN(n8603) );
  NAND2_X1 U10200 ( .A1(n8603), .A2(n8622), .ZN(n8608) );
  OAI22_X1 U10201 ( .A1(n8813), .A2(n8614), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8604), .ZN(n8606) );
  OAI22_X1 U10202 ( .A1(n8615), .A2(n8812), .B1(n8804), .B2(n8628), .ZN(n8605)
         );
  AOI211_X1 U10203 ( .C1(n8977), .C2(n8618), .A(n8606), .B(n8605), .ZN(n8607)
         );
  NAND2_X1 U10204 ( .A1(n8608), .A2(n8607), .ZN(P2_U3237) );
  NAND2_X1 U10205 ( .A1(n8610), .A2(n8609), .ZN(n8612) );
  XNOR2_X1 U10206 ( .A(n8612), .B(n8611), .ZN(n8621) );
  NAND2_X1 U10207 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8676) );
  OAI21_X1 U10208 ( .B1(n8614), .B2(n8613), .A(n8676), .ZN(n8617) );
  OAI22_X1 U10209 ( .A1(n8615), .A2(n8869), .B1(n8872), .B2(n8628), .ZN(n8616)
         );
  AOI211_X1 U10210 ( .C1(n4584), .C2(n8618), .A(n8617), .B(n8616), .ZN(n8619)
         );
  OAI21_X1 U10211 ( .B1(n8621), .B2(n8620), .A(n8619), .ZN(P2_U3240) );
  OAI211_X1 U10212 ( .C1(n8625), .C2(n8624), .A(n8623), .B(n8622), .ZN(n8633)
         );
  OAI22_X1 U10213 ( .A1(n8626), .A2(n8886), .B1(n8777), .B2(n8884), .ZN(n8748)
         );
  INV_X1 U10214 ( .A(n8743), .ZN(n8629) );
  OAI22_X1 U10215 ( .A1(n8629), .A2(n8628), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8627), .ZN(n8630) );
  AOI21_X1 U10216 ( .B1(n8748), .B2(n8631), .A(n8630), .ZN(n8632) );
  OAI211_X1 U10217 ( .C1(n4597), .C2(n8634), .A(n8633), .B(n8632), .ZN(
        P2_U3242) );
  MUX2_X1 U10218 ( .A(n8635), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8649), .Z(
        P2_U3582) );
  MUX2_X1 U10219 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8636), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U10220 ( .A(n8735), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8649), .Z(
        P2_U3580) );
  MUX2_X1 U10221 ( .A(n8637), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8649), .Z(
        P2_U3579) );
  MUX2_X1 U10222 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8734), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U10223 ( .A(n8789), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8649), .Z(
        P2_U3576) );
  MUX2_X1 U10224 ( .A(n8826), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8649), .Z(
        P2_U3574) );
  MUX2_X1 U10225 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8124), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10226 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8853), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10227 ( .A(n8867), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8649), .Z(
        P2_U3571) );
  MUX2_X1 U10228 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8119), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10229 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8903), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10230 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8931), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10231 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8902), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10232 ( .A(n8929), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8649), .Z(
        P2_U3566) );
  MUX2_X1 U10233 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8638), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U10234 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8639), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10235 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8640), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10236 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8641), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U10237 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8642), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U10238 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8643), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U10239 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8644), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U10240 ( .A(n8645), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8649), .Z(
        P2_U3557) );
  MUX2_X1 U10241 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8646), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U10242 ( .A(n8647), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8649), .Z(
        P2_U3555) );
  MUX2_X1 U10243 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8648), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U10244 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n5941), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U10245 ( .A(n8650), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8649), .Z(
        P2_U3552) );
  NAND2_X1 U10246 ( .A1(n8678), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8653) );
  OAI21_X1 U10247 ( .B1(n8678), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8653), .ZN(
        n8654) );
  AOI211_X1 U10248 ( .C1(n8655), .C2(n8654), .A(n10263), .B(n8672), .ZN(n8671)
         );
  XNOR2_X1 U10249 ( .A(n8678), .B(n8656), .ZN(n8660) );
  NAND2_X1 U10250 ( .A1(n8658), .A2(n8657), .ZN(n8661) );
  AND2_X1 U10251 ( .A1(n8660), .A2(n8661), .ZN(n8659) );
  NAND2_X1 U10252 ( .A1(n8662), .A2(n8659), .ZN(n8684) );
  INV_X1 U10253 ( .A(n8684), .ZN(n8664) );
  AOI21_X1 U10254 ( .B1(n8662), .B2(n8661), .A(n8660), .ZN(n8663) );
  NOR3_X1 U10255 ( .A1(n8664), .A2(n8663), .A3(n10262), .ZN(n8670) );
  NOR2_X1 U10256 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8665), .ZN(n8666) );
  AOI21_X1 U10257 ( .B1(n10260), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8666), .ZN(
        n8667) );
  OAI21_X1 U10258 ( .B1(n10261), .B2(n8668), .A(n8667), .ZN(n8669) );
  OR3_X1 U10259 ( .A1(n8671), .A2(n8670), .A3(n8669), .ZN(P2_U3262) );
  NOR2_X1 U10260 ( .A1(n8674), .A2(n8673), .ZN(n8691) );
  OAI21_X1 U10261 ( .B1(n8675), .B2(P2_REG2_REG_18__SCAN_IN), .A(n10259), .ZN(
        n8689) );
  OAI21_X1 U10262 ( .B1(n8705), .B2(n10450), .A(n8676), .ZN(n8677) );
  AOI21_X1 U10263 ( .B1(n9921), .B2(n8679), .A(n8677), .ZN(n8688) );
  NAND2_X1 U10264 ( .A1(n8678), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8683) );
  OR2_X1 U10265 ( .A1(n8679), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8692) );
  NAND2_X1 U10266 ( .A1(n8679), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8680) );
  AND2_X1 U10267 ( .A1(n8692), .A2(n8680), .ZN(n8682) );
  AND2_X1 U10268 ( .A1(n8683), .A2(n8682), .ZN(n8681) );
  NAND2_X1 U10269 ( .A1(n8684), .A2(n8681), .ZN(n8693) );
  INV_X1 U10270 ( .A(n8693), .ZN(n8686) );
  AOI21_X1 U10271 ( .B1(n8684), .B2(n8683), .A(n8682), .ZN(n8685) );
  OAI21_X1 U10272 ( .B1(n8686), .B2(n8685), .A(n10258), .ZN(n8687) );
  OAI211_X1 U10273 ( .C1(n8690), .C2(n8689), .A(n8688), .B(n8687), .ZN(
        P2_U3263) );
  XNOR2_X1 U10274 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n4508), .ZN(n8700) );
  NAND2_X1 U10275 ( .A1(n8693), .A2(n8692), .ZN(n8695) );
  XNOR2_X1 U10276 ( .A(n8695), .B(n8694), .ZN(n8698) );
  AOI21_X1 U10277 ( .B1(n8698), .B2(n10258), .A(n9921), .ZN(n8696) );
  OAI21_X1 U10278 ( .B1(n8700), .B2(n10263), .A(n8696), .ZN(n8697) );
  INV_X1 U10279 ( .A(n8697), .ZN(n8703) );
  INV_X1 U10280 ( .A(n8698), .ZN(n8699) );
  AOI22_X1 U10281 ( .A1(n8700), .A2(n10259), .B1(n8699), .B2(n10258), .ZN(
        n8702) );
  AOI21_X1 U10282 ( .B1(n8709), .B2(n8708), .A(n8707), .ZN(n8942) );
  NAND2_X1 U10283 ( .A1(n8942), .A2(n8936), .ZN(n8712) );
  AOI21_X1 U10284 ( .B1(n10293), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8710), .ZN(
        n8711) );
  OAI211_X1 U10285 ( .C1(n8945), .C2(n8924), .A(n8712), .B(n8711), .ZN(
        P2_U3266) );
  OAI22_X1 U10286 ( .A1(n8714), .A2(n8912), .B1(n8713), .B2(n8915), .ZN(n8715)
         );
  AOI21_X1 U10287 ( .B1(n8716), .B2(n10284), .A(n8715), .ZN(n8719) );
  NAND2_X1 U10288 ( .A1(n8717), .A2(n8936), .ZN(n8718) );
  OAI211_X1 U10289 ( .C1(n8720), .C2(n10293), .A(n8719), .B(n8718), .ZN(n8721)
         );
  AOI21_X1 U10290 ( .B1(n8722), .B2(n10288), .A(n8721), .ZN(n8723) );
  INV_X1 U10291 ( .A(n8723), .ZN(P2_U3267) );
  XOR2_X1 U10292 ( .A(n8724), .B(n8733), .Z(n8955) );
  INV_X1 U10293 ( .A(n8725), .ZN(n8726) );
  AOI21_X1 U10294 ( .B1(n8951), .B2(n8741), .A(n8726), .ZN(n8952) );
  AOI22_X1 U10295 ( .A1(n8727), .A2(n10283), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n10293), .ZN(n8728) );
  OAI21_X1 U10296 ( .B1(n8729), .B2(n8924), .A(n8728), .ZN(n8738) );
  NAND2_X1 U10297 ( .A1(n8731), .A2(n8730), .ZN(n8732) );
  XOR2_X1 U10298 ( .A(n8733), .B(n8732), .Z(n8736) );
  AOI222_X1 U10299 ( .A1(n8933), .A2(n8736), .B1(n8735), .B2(n8930), .C1(n8734), .C2(n8928), .ZN(n8954) );
  NOR2_X1 U10300 ( .A1(n8954), .A2(n10293), .ZN(n8737) );
  AOI211_X1 U10301 ( .C1(n8936), .C2(n8952), .A(n8738), .B(n8737), .ZN(n8739)
         );
  OAI21_X1 U10302 ( .B1(n8955), .B2(n8938), .A(n8739), .ZN(P2_U3269) );
  XOR2_X1 U10303 ( .A(n8747), .B(n8740), .Z(n8960) );
  INV_X1 U10304 ( .A(n8741), .ZN(n8742) );
  AOI211_X1 U10305 ( .C1(n8957), .C2(n8760), .A(n4832), .B(n8742), .ZN(n8956)
         );
  AOI22_X1 U10306 ( .A1(n8743), .A2(n10283), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n10293), .ZN(n8744) );
  OAI21_X1 U10307 ( .B1(n4597), .B2(n8924), .A(n8744), .ZN(n8751) );
  NAND2_X1 U10308 ( .A1(n8755), .A2(n8745), .ZN(n8746) );
  XOR2_X1 U10309 ( .A(n8747), .B(n8746), .Z(n8749) );
  AOI21_X1 U10310 ( .B1(n8749), .B2(n8933), .A(n8748), .ZN(n8959) );
  NOR2_X1 U10311 ( .A1(n8959), .A2(n10293), .ZN(n8750) );
  AOI211_X1 U10312 ( .C1(n8956), .C2(n10287), .A(n8751), .B(n8750), .ZN(n8752)
         );
  OAI21_X1 U10313 ( .B1(n8960), .B2(n8938), .A(n8752), .ZN(P2_U3270) );
  XNOR2_X1 U10314 ( .A(n8754), .B(n8756), .ZN(n8965) );
  OAI211_X1 U10315 ( .C1(n8757), .C2(n8756), .A(n8755), .B(n8933), .ZN(n8759)
         );
  NAND2_X1 U10316 ( .A1(n8759), .A2(n8758), .ZN(n8961) );
  AOI211_X1 U10317 ( .C1(n8963), .C2(n4489), .A(n4832), .B(n4598), .ZN(n8962)
         );
  NAND2_X1 U10318 ( .A1(n8962), .A2(n10287), .ZN(n8764) );
  INV_X1 U10319 ( .A(n8761), .ZN(n8762) );
  AOI22_X1 U10320 ( .A1(n8762), .A2(n10283), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n10293), .ZN(n8763) );
  OAI211_X1 U10321 ( .C1(n8765), .C2(n8924), .A(n8764), .B(n8763), .ZN(n8766)
         );
  AOI21_X1 U10322 ( .B1(n8961), .B2(n8915), .A(n8766), .ZN(n8767) );
  OAI21_X1 U10323 ( .B1(n8965), .B2(n8938), .A(n8767), .ZN(P2_U3271) );
  INV_X1 U10324 ( .A(n8768), .ZN(n8769) );
  AOI21_X1 U10325 ( .B1(n8771), .B2(n8770), .A(n8769), .ZN(n8970) );
  XNOR2_X1 U10326 ( .A(n8794), .B(n8966), .ZN(n8967) );
  INV_X1 U10327 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8772) );
  OAI22_X1 U10328 ( .A1(n8773), .A2(n8924), .B1(n8915), .B2(n8772), .ZN(n8774)
         );
  AOI21_X1 U10329 ( .B1(n8967), .B2(n8936), .A(n8774), .ZN(n8784) );
  AOI21_X1 U10330 ( .B1(n8776), .B2(n8775), .A(n9966), .ZN(n8780) );
  OAI22_X1 U10331 ( .A1(n8777), .A2(n8886), .B1(n8813), .B2(n8884), .ZN(n8778)
         );
  AOI21_X1 U10332 ( .B1(n8780), .B2(n8779), .A(n8778), .ZN(n8969) );
  OAI21_X1 U10333 ( .B1(n8781), .B2(n8912), .A(n8969), .ZN(n8782) );
  NAND2_X1 U10334 ( .A1(n8782), .A2(n8915), .ZN(n8783) );
  OAI211_X1 U10335 ( .C1(n8970), .C2(n8938), .A(n8784), .B(n8783), .ZN(
        P2_U3272) );
  INV_X1 U10336 ( .A(n8785), .ZN(n8809) );
  OAI21_X1 U10337 ( .B1(n8809), .B2(n8786), .A(n8791), .ZN(n8788) );
  NAND2_X1 U10338 ( .A1(n8788), .A2(n8787), .ZN(n8790) );
  AOI222_X1 U10339 ( .A1(n8933), .A2(n8790), .B1(n8789), .B2(n8930), .C1(n8826), .C2(n8928), .ZN(n8975) );
  OR2_X1 U10340 ( .A1(n8792), .A2(n8791), .ZN(n8971) );
  NAND3_X1 U10341 ( .A1(n8971), .A2(n8793), .A3(n10288), .ZN(n8800) );
  AOI21_X1 U10342 ( .B1(n8972), .B2(n8802), .A(n8794), .ZN(n8973) );
  AOI22_X1 U10343 ( .A1(n8795), .A2(n10283), .B1(n10293), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n8796) );
  OAI21_X1 U10344 ( .B1(n8797), .B2(n8924), .A(n8796), .ZN(n8798) );
  AOI21_X1 U10345 ( .B1(n8973), .B2(n8936), .A(n8798), .ZN(n8799) );
  OAI211_X1 U10346 ( .C1(n10293), .C2(n8975), .A(n8800), .B(n8799), .ZN(
        P2_U3273) );
  XOR2_X1 U10347 ( .A(n8801), .B(n8811), .Z(n8981) );
  AOI21_X1 U10348 ( .B1(n8977), .B2(n8803), .A(n4750), .ZN(n8978) );
  INV_X1 U10349 ( .A(n8804), .ZN(n8805) );
  AOI22_X1 U10350 ( .A1(P2_REG2_REG_22__SCAN_IN), .A2(n10293), .B1(n8805), 
        .B2(n10283), .ZN(n8806) );
  OAI21_X1 U10351 ( .B1(n8807), .B2(n8924), .A(n8806), .ZN(n8817) );
  NAND2_X1 U10352 ( .A1(n8825), .A2(n8808), .ZN(n8810) );
  AOI211_X1 U10353 ( .C1(n8811), .C2(n8810), .A(n9966), .B(n8809), .ZN(n8815)
         );
  OAI22_X1 U10354 ( .A1(n8813), .A2(n8886), .B1(n8812), .B2(n8884), .ZN(n8814)
         );
  NOR2_X1 U10355 ( .A1(n8815), .A2(n8814), .ZN(n8980) );
  NOR2_X1 U10356 ( .A1(n8980), .A2(n10293), .ZN(n8816) );
  AOI211_X1 U10357 ( .C1(n8978), .C2(n8936), .A(n8817), .B(n8816), .ZN(n8818)
         );
  OAI21_X1 U10358 ( .B1(n8981), .B2(n8938), .A(n8818), .ZN(P2_U3274) );
  XOR2_X1 U10359 ( .A(n8819), .B(n8824), .Z(n8986) );
  XNOR2_X1 U10360 ( .A(n8832), .B(n8982), .ZN(n8983) );
  INV_X1 U10361 ( .A(n8820), .ZN(n8821) );
  AOI22_X1 U10362 ( .A1(n10293), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8821), 
        .B2(n10283), .ZN(n8822) );
  OAI21_X1 U10363 ( .B1(n8823), .B2(n8924), .A(n8822), .ZN(n8829) );
  OAI21_X1 U10364 ( .B1(n5032), .B2(n6206), .A(n8825), .ZN(n8827) );
  AOI222_X1 U10365 ( .A1(n8933), .A2(n8827), .B1(n8826), .B2(n8930), .C1(n8853), .C2(n8928), .ZN(n8985) );
  NOR2_X1 U10366 ( .A1(n8985), .A2(n10293), .ZN(n8828) );
  AOI211_X1 U10367 ( .C1(n8983), .C2(n8936), .A(n8829), .B(n8828), .ZN(n8830)
         );
  OAI21_X1 U10368 ( .B1(n8986), .B2(n8938), .A(n8830), .ZN(P2_U3275) );
  XNOR2_X1 U10369 ( .A(n8831), .B(n8839), .ZN(n8991) );
  AOI21_X1 U10370 ( .B1(n8987), .B2(n4551), .A(n8832), .ZN(n8988) );
  AOI22_X1 U10371 ( .A1(n10293), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8833), 
        .B2(n10283), .ZN(n8834) );
  OAI21_X1 U10372 ( .B1(n8835), .B2(n8924), .A(n8834), .ZN(n8842) );
  NAND2_X1 U10373 ( .A1(n8836), .A2(n8837), .ZN(n8838) );
  XOR2_X1 U10374 ( .A(n8839), .B(n8838), .Z(n8840) );
  AOI222_X1 U10375 ( .A1(n8867), .A2(n8928), .B1(n8124), .B2(n8930), .C1(n8933), .C2(n8840), .ZN(n8990) );
  NOR2_X1 U10376 ( .A1(n8990), .A2(n10293), .ZN(n8841) );
  AOI211_X1 U10377 ( .C1(n8988), .C2(n8936), .A(n8842), .B(n8841), .ZN(n8843)
         );
  OAI21_X1 U10378 ( .B1(n8991), .B2(n8938), .A(n8843), .ZN(P2_U3276) );
  XOR2_X1 U10379 ( .A(n8844), .B(n8848), .Z(n8997) );
  NOR2_X1 U10380 ( .A1(n8997), .A2(n8845), .ZN(n8856) );
  OAI211_X1 U10381 ( .C1(n8847), .C2(n8846), .A(n4551), .B(n9978), .ZN(n8992)
         );
  INV_X1 U10382 ( .A(n8848), .ZN(n8850) );
  NAND3_X1 U10383 ( .A1(n8851), .A2(n8850), .A3(n8849), .ZN(n8852) );
  NAND2_X1 U10384 ( .A1(n8836), .A2(n8852), .ZN(n8854) );
  AOI222_X1 U10385 ( .A1(n8933), .A2(n8854), .B1(n8853), .B2(n8930), .C1(n8119), .C2(n8928), .ZN(n8996) );
  OAI21_X1 U10386 ( .B1(n4831), .B2(n8992), .A(n8996), .ZN(n8855) );
  OAI21_X1 U10387 ( .B1(n8856), .B2(n8855), .A(n8915), .ZN(n8861) );
  OAI22_X1 U10388 ( .A1(n8915), .A2(n8858), .B1(n8857), .B2(n8912), .ZN(n8859)
         );
  AOI21_X1 U10389 ( .B1(n8994), .B2(n10284), .A(n8859), .ZN(n8860) );
  OAI211_X1 U10390 ( .C1(n8997), .C2(n8862), .A(n8861), .B(n8860), .ZN(
        P2_U3277) );
  XOR2_X1 U10391 ( .A(n8863), .B(n8865), .Z(n9002) );
  NAND2_X1 U10392 ( .A1(n8881), .A2(n8864), .ZN(n8866) );
  XNOR2_X1 U10393 ( .A(n8866), .B(n8865), .ZN(n8871) );
  NAND2_X1 U10394 ( .A1(n8867), .A2(n8930), .ZN(n8868) );
  OAI21_X1 U10395 ( .B1(n8869), .B2(n8884), .A(n8868), .ZN(n8870) );
  AOI21_X1 U10396 ( .B1(n8871), .B2(n8933), .A(n8870), .ZN(n9001) );
  OAI22_X1 U10397 ( .A1(n8915), .A2(n8873), .B1(n8872), .B2(n8912), .ZN(n8874)
         );
  AOI21_X1 U10398 ( .B1(n4584), .B2(n10284), .A(n8874), .ZN(n8877) );
  XNOR2_X1 U10399 ( .A(n4554), .B(n8875), .ZN(n8999) );
  NAND2_X1 U10400 ( .A1(n8999), .A2(n8936), .ZN(n8876) );
  OAI211_X1 U10401 ( .C1(n9001), .C2(n10293), .A(n8877), .B(n8876), .ZN(n8878)
         );
  INV_X1 U10402 ( .A(n8878), .ZN(n8879) );
  OAI21_X1 U10403 ( .B1(n9002), .B2(n8938), .A(n8879), .ZN(P2_U3278) );
  NAND2_X1 U10404 ( .A1(n8900), .A2(n8880), .ZN(n8883) );
  INV_X1 U10405 ( .A(n8881), .ZN(n8882) );
  AOI211_X1 U10406 ( .C1(n8891), .C2(n8883), .A(n9966), .B(n8882), .ZN(n8889)
         );
  OAI22_X1 U10407 ( .A1(n8887), .A2(n8886), .B1(n8885), .B2(n8884), .ZN(n8888)
         );
  NOR2_X1 U10408 ( .A1(n8889), .A2(n8888), .ZN(n9007) );
  OAI21_X1 U10409 ( .B1(n4564), .B2(n8891), .A(n8890), .ZN(n9003) );
  NAND2_X1 U10410 ( .A1(n9003), .A2(n10288), .ZN(n8899) );
  INV_X1 U10411 ( .A(n4554), .ZN(n8892) );
  AOI211_X1 U10412 ( .C1(n9005), .C2(n8908), .A(n4832), .B(n8892), .ZN(n9004)
         );
  INV_X1 U10413 ( .A(n9005), .ZN(n8893) );
  NOR2_X1 U10414 ( .A1(n8893), .A2(n8924), .ZN(n8897) );
  INV_X1 U10415 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8895) );
  OAI22_X1 U10416 ( .A1(n8915), .A2(n8895), .B1(n8894), .B2(n8912), .ZN(n8896)
         );
  AOI211_X1 U10417 ( .C1(n9004), .C2(n10287), .A(n8897), .B(n8896), .ZN(n8898)
         );
  OAI211_X1 U10418 ( .C1(n10293), .C2(n9007), .A(n8899), .B(n8898), .ZN(
        P2_U3279) );
  OAI21_X1 U10419 ( .B1(n8905), .B2(n8901), .A(n8900), .ZN(n8904) );
  AOI222_X1 U10420 ( .A1(n8933), .A2(n8904), .B1(n8903), .B2(n8930), .C1(n8902), .C2(n8928), .ZN(n9013) );
  INV_X1 U10421 ( .A(n9015), .ZN(n8907) );
  NAND2_X1 U10422 ( .A1(n8906), .A2(n8905), .ZN(n9009) );
  NAND3_X1 U10423 ( .A1(n8907), .A2(n10288), .A3(n9009), .ZN(n8919) );
  INV_X1 U10424 ( .A(n8908), .ZN(n8909) );
  AOI21_X1 U10425 ( .B1(n9010), .B2(n8910), .A(n8909), .ZN(n9011) );
  INV_X1 U10426 ( .A(n9010), .ZN(n8911) );
  NOR2_X1 U10427 ( .A1(n8911), .A2(n8924), .ZN(n8917) );
  OAI22_X1 U10428 ( .A1(n8915), .A2(n8914), .B1(n8913), .B2(n8912), .ZN(n8916)
         );
  AOI211_X1 U10429 ( .C1(n9011), .C2(n8936), .A(n8917), .B(n8916), .ZN(n8918)
         );
  OAI211_X1 U10430 ( .C1(n10293), .C2(n9013), .A(n8919), .B(n8918), .ZN(
        P2_U3280) );
  XOR2_X1 U10431 ( .A(n8927), .B(n8920), .Z(n9021) );
  XNOR2_X1 U10432 ( .A(n9977), .B(n9016), .ZN(n9017) );
  INV_X1 U10433 ( .A(n8921), .ZN(n8922) );
  AOI22_X1 U10434 ( .A1(n10293), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8922), 
        .B2(n10283), .ZN(n8923) );
  OAI21_X1 U10435 ( .B1(n8925), .B2(n8924), .A(n8923), .ZN(n8935) );
  XOR2_X1 U10436 ( .A(n8927), .B(n8926), .Z(n8932) );
  AOI222_X1 U10437 ( .A1(n8933), .A2(n8932), .B1(n8931), .B2(n8930), .C1(n8929), .C2(n8928), .ZN(n9019) );
  NOR2_X1 U10438 ( .A1(n9019), .A2(n10293), .ZN(n8934) );
  AOI211_X1 U10439 ( .C1(n9017), .C2(n8936), .A(n8935), .B(n8934), .ZN(n8937)
         );
  OAI21_X1 U10440 ( .B1(n9021), .B2(n8938), .A(n8937), .ZN(P2_U3281) );
  NAND2_X1 U10441 ( .A1(n8939), .A2(n9978), .ZN(n8940) );
  OAI211_X1 U10442 ( .C1(n10381), .C2(n8941), .A(n8940), .B(n8943), .ZN(n9028)
         );
  MUX2_X1 U10443 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9028), .S(n10406), .Z(
        P2_U3551) );
  NAND2_X1 U10444 ( .A1(n8942), .A2(n9978), .ZN(n8944) );
  OAI211_X1 U10445 ( .C1(n8945), .C2(n10381), .A(n8944), .B(n8943), .ZN(n9029)
         );
  MUX2_X1 U10446 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9029), .S(n10406), .Z(
        P2_U3550) );
  AOI22_X1 U10447 ( .A1(n8947), .A2(n9978), .B1(n10385), .B2(n8946), .ZN(n8948) );
  OAI211_X1 U10448 ( .C1(n8950), .C2(n9020), .A(n8949), .B(n8948), .ZN(n9030)
         );
  MUX2_X1 U10449 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9030), .S(n10406), .Z(
        P2_U3548) );
  AOI22_X1 U10450 ( .A1(n8952), .A2(n9978), .B1(n10385), .B2(n8951), .ZN(n8953) );
  OAI211_X1 U10451 ( .C1(n8955), .C2(n9020), .A(n8954), .B(n8953), .ZN(n9031)
         );
  MUX2_X1 U10452 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9031), .S(n10406), .Z(
        P2_U3547) );
  AOI21_X1 U10453 ( .B1(n10385), .B2(n8957), .A(n8956), .ZN(n8958) );
  OAI211_X1 U10454 ( .C1(n8960), .C2(n9020), .A(n8959), .B(n8958), .ZN(n9032)
         );
  MUX2_X1 U10455 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9032), .S(n10406), .Z(
        P2_U3546) );
  AOI211_X1 U10456 ( .C1(n10385), .C2(n8963), .A(n8962), .B(n8961), .ZN(n8964)
         );
  OAI21_X1 U10457 ( .B1(n8965), .B2(n9020), .A(n8964), .ZN(n9033) );
  MUX2_X1 U10458 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9033), .S(n10406), .Z(
        P2_U3545) );
  AOI22_X1 U10459 ( .A1(n8967), .A2(n9978), .B1(n10385), .B2(n8966), .ZN(n8968) );
  OAI211_X1 U10460 ( .C1(n8970), .C2(n9020), .A(n8969), .B(n8968), .ZN(n9034)
         );
  MUX2_X1 U10461 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9034), .S(n10406), .Z(
        P2_U3544) );
  NAND3_X1 U10462 ( .A1(n8971), .A2(n8793), .A3(n10391), .ZN(n8976) );
  AOI22_X1 U10463 ( .A1(n8973), .A2(n9978), .B1(n10385), .B2(n8972), .ZN(n8974) );
  NAND3_X1 U10464 ( .A1(n8976), .A2(n8975), .A3(n8974), .ZN(n9035) );
  MUX2_X1 U10465 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9035), .S(n10406), .Z(
        P2_U3543) );
  AOI22_X1 U10466 ( .A1(n8978), .A2(n9978), .B1(n10385), .B2(n8977), .ZN(n8979) );
  OAI211_X1 U10467 ( .C1(n8981), .C2(n9020), .A(n8980), .B(n8979), .ZN(n9036)
         );
  MUX2_X1 U10468 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9036), .S(n10406), .Z(
        P2_U3542) );
  AOI22_X1 U10469 ( .A1(n8983), .A2(n9978), .B1(n10385), .B2(n8982), .ZN(n8984) );
  OAI211_X1 U10470 ( .C1(n8986), .C2(n9020), .A(n8985), .B(n8984), .ZN(n9037)
         );
  MUX2_X1 U10471 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9037), .S(n10406), .Z(
        P2_U3541) );
  AOI22_X1 U10472 ( .A1(n8988), .A2(n9978), .B1(n10385), .B2(n8987), .ZN(n8989) );
  OAI211_X1 U10473 ( .C1(n8991), .C2(n9020), .A(n8990), .B(n8989), .ZN(n9038)
         );
  MUX2_X1 U10474 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9038), .S(n10406), .Z(
        P2_U3540) );
  INV_X1 U10475 ( .A(n8992), .ZN(n8993) );
  AOI21_X1 U10476 ( .B1(n10385), .B2(n8994), .A(n8993), .ZN(n8995) );
  OAI211_X1 U10477 ( .C1(n8997), .C2(n9020), .A(n8996), .B(n8995), .ZN(n9039)
         );
  MUX2_X1 U10478 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9039), .S(n10406), .Z(
        P2_U3539) );
  AOI22_X1 U10479 ( .A1(n8999), .A2(n9978), .B1(n10385), .B2(n4584), .ZN(n9000) );
  OAI211_X1 U10480 ( .C1(n9002), .C2(n9020), .A(n9001), .B(n9000), .ZN(n9040)
         );
  MUX2_X1 U10481 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9040), .S(n10406), .Z(
        P2_U3538) );
  INV_X1 U10482 ( .A(n9003), .ZN(n9008) );
  AOI21_X1 U10483 ( .B1(n10385), .B2(n9005), .A(n9004), .ZN(n9006) );
  OAI211_X1 U10484 ( .C1(n9008), .C2(n9020), .A(n9007), .B(n9006), .ZN(n9041)
         );
  MUX2_X1 U10485 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9041), .S(n10406), .Z(
        P2_U3537) );
  NAND2_X1 U10486 ( .A1(n9009), .A2(n10391), .ZN(n9014) );
  AOI22_X1 U10487 ( .A1(n9011), .A2(n9978), .B1(n10385), .B2(n9010), .ZN(n9012) );
  OAI211_X1 U10488 ( .C1(n9015), .C2(n9014), .A(n9013), .B(n9012), .ZN(n9042)
         );
  MUX2_X1 U10489 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9042), .S(n10406), .Z(
        P2_U3536) );
  AOI22_X1 U10490 ( .A1(n9017), .A2(n9978), .B1(n10385), .B2(n9016), .ZN(n9018) );
  OAI211_X1 U10491 ( .C1(n9021), .C2(n9020), .A(n9019), .B(n9018), .ZN(n9043)
         );
  MUX2_X1 U10492 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9043), .S(n10406), .Z(
        P2_U3535) );
  OAI22_X1 U10493 ( .A1(n9023), .A2(n4832), .B1(n9022), .B2(n10381), .ZN(n9024) );
  INV_X1 U10494 ( .A(n9024), .ZN(n9025) );
  OAI211_X1 U10495 ( .C1(n10357), .C2(n9027), .A(n9026), .B(n9025), .ZN(n9044)
         );
  MUX2_X1 U10496 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9044), .S(n10406), .Z(
        P2_U3533) );
  MUX2_X1 U10497 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9028), .S(n10395), .Z(
        P2_U3519) );
  MUX2_X1 U10498 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9029), .S(n10395), .Z(
        P2_U3518) );
  MUX2_X1 U10499 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9030), .S(n10395), .Z(
        P2_U3516) );
  MUX2_X1 U10500 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9031), .S(n10395), .Z(
        P2_U3515) );
  MUX2_X1 U10501 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9032), .S(n10395), .Z(
        P2_U3514) );
  MUX2_X1 U10502 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9033), .S(n10395), .Z(
        P2_U3513) );
  MUX2_X1 U10503 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9034), .S(n10395), .Z(
        P2_U3512) );
  MUX2_X1 U10504 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9035), .S(n10395), .Z(
        P2_U3511) );
  MUX2_X1 U10505 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9036), .S(n10395), .Z(
        P2_U3510) );
  MUX2_X1 U10506 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9037), .S(n10395), .Z(
        P2_U3509) );
  MUX2_X1 U10507 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9038), .S(n10395), .Z(
        P2_U3508) );
  MUX2_X1 U10508 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9039), .S(n10395), .Z(
        P2_U3507) );
  MUX2_X1 U10509 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9040), .S(n10395), .Z(
        P2_U3505) );
  MUX2_X1 U10510 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9041), .S(n10395), .Z(
        P2_U3502) );
  MUX2_X1 U10511 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9042), .S(n10395), .Z(
        P2_U3499) );
  MUX2_X1 U10512 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9043), .S(n10395), .Z(
        P2_U3496) );
  MUX2_X1 U10513 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9044), .S(n10395), .Z(
        P2_U3490) );
  INV_X1 U10514 ( .A(n9169), .ZN(n9900) );
  NOR4_X1 U10515 ( .A1(n9045), .A2(P2_IR_REG_30__SCAN_IN), .A3(n6083), .A4(
        P2_U3152), .ZN(n9046) );
  AOI21_X1 U10516 ( .B1(n9047), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9046), .ZN(
        n9048) );
  OAI21_X1 U10517 ( .B1(n9900), .B2(n4481), .A(n9048), .ZN(P2_U3327) );
  OAI222_X1 U10518 ( .A1(P2_U3152), .A2(n9049), .B1(n4481), .B2(n9052), .C1(
        n9051), .C2(n9050), .ZN(P2_U3328) );
  MUX2_X1 U10519 ( .A(n9053), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10520 ( .A(n9055), .ZN(n9060) );
  AOI21_X1 U10521 ( .B1(n9056), .B2(n9055), .A(n9054), .ZN(n9057) );
  NOR2_X1 U10522 ( .A1(n9057), .A2(n9139), .ZN(n9058) );
  OAI21_X1 U10523 ( .B1(n9060), .B2(n9059), .A(n9058), .ZN(n9066) );
  OAI21_X1 U10524 ( .B1(n9188), .B2(n9161), .A(n9061), .ZN(n9064) );
  NOR2_X1 U10525 ( .A1(n9158), .A2(n9062), .ZN(n9063) );
  AOI211_X1 U10526 ( .C1(n10469), .C2(n9470), .A(n9064), .B(n9063), .ZN(n9065)
         );
  OAI211_X1 U10527 ( .C1(n9067), .C2(n9151), .A(n9066), .B(n9065), .ZN(
        P1_U3213) );
  NOR2_X1 U10528 ( .A1(n9113), .A2(n9068), .ZN(n9069) );
  XOR2_X1 U10529 ( .A(n9070), .B(n9069), .Z(n9075) );
  AOI22_X1 U10530 ( .A1(n10469), .A2(n9642), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9072) );
  NAND2_X1 U10531 ( .A1(n9134), .A2(n9666), .ZN(n9071) );
  OAI211_X1 U10532 ( .C1(n9158), .C2(n9632), .A(n9072), .B(n9071), .ZN(n9073)
         );
  AOI21_X1 U10533 ( .B1(n9816), .B2(n9165), .A(n9073), .ZN(n9074) );
  OAI21_X1 U10534 ( .B1(n9075), .B2(n9139), .A(n9074), .ZN(P1_U3214) );
  XOR2_X1 U10535 ( .A(n9076), .B(n9077), .Z(n9084) );
  OAI22_X1 U10536 ( .A1(n9079), .A2(n9161), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9078), .ZN(n9080) );
  AOI21_X1 U10537 ( .B1(n10469), .B2(n9666), .A(n9080), .ZN(n9081) );
  OAI21_X1 U10538 ( .B1(n9158), .B2(n9673), .A(n9081), .ZN(n9082) );
  AOI21_X1 U10539 ( .B1(n9827), .B2(n9165), .A(n9082), .ZN(n9083) );
  OAI21_X1 U10540 ( .B1(n9084), .B2(n9139), .A(n9083), .ZN(P1_U3221) );
  AOI21_X1 U10541 ( .B1(n9087), .B2(n9086), .A(n9085), .ZN(n9092) );
  AOI22_X1 U10542 ( .A1(n9468), .A2(n10469), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9089) );
  NAND2_X1 U10543 ( .A1(n9134), .A2(n9642), .ZN(n9088) );
  OAI211_X1 U10544 ( .C1(n9158), .C2(n9604), .A(n9089), .B(n9088), .ZN(n9090)
         );
  AOI21_X1 U10545 ( .B1(n9808), .B2(n9165), .A(n9090), .ZN(n9091) );
  OAI21_X1 U10546 ( .B1(n9092), .B2(n9139), .A(n9091), .ZN(P1_U3223) );
  XOR2_X1 U10547 ( .A(n9095), .B(n9094), .Z(n9096) );
  XNOR2_X1 U10548 ( .A(n9093), .B(n9096), .ZN(n9101) );
  NAND2_X1 U10549 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10147)
         );
  OAI21_X1 U10550 ( .B1(n9117), .B2(n9752), .A(n10147), .ZN(n9097) );
  AOI21_X1 U10551 ( .B1(n9134), .B2(n9470), .A(n9097), .ZN(n9098) );
  OAI21_X1 U10552 ( .B1(n9158), .B2(n9744), .A(n9098), .ZN(n9099) );
  AOI21_X1 U10553 ( .B1(n9853), .B2(n9165), .A(n9099), .ZN(n9100) );
  OAI21_X1 U10554 ( .B1(n9101), .B2(n9139), .A(n9100), .ZN(P1_U3224) );
  INV_X1 U10555 ( .A(n9103), .ZN(n9104) );
  AOI21_X1 U10556 ( .B1(n9105), .B2(n9102), .A(n9104), .ZN(n9111) );
  NAND2_X1 U10557 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10160)
         );
  OAI21_X1 U10558 ( .B1(n9117), .B2(n9106), .A(n10160), .ZN(n9108) );
  NOR2_X1 U10559 ( .A1(n9158), .A2(n9724), .ZN(n9107) );
  AOI211_X1 U10560 ( .C1(n9134), .C2(n9730), .A(n9108), .B(n9107), .ZN(n9110)
         );
  NAND2_X1 U10561 ( .A1(n9846), .A2(n9165), .ZN(n9109) );
  OAI211_X1 U10562 ( .C1(n9111), .C2(n9139), .A(n9110), .B(n9109), .ZN(
        P1_U3226) );
  OAI21_X1 U10563 ( .B1(n4518), .B2(n9113), .A(n9112), .ZN(n9114) );
  INV_X1 U10564 ( .A(n9114), .ZN(n9115) );
  OAI21_X1 U10565 ( .B1(n4501), .B2(n9115), .A(n9152), .ZN(n9121) );
  NOR2_X1 U10566 ( .A1(n9158), .A2(n9618), .ZN(n9119) );
  OAI22_X1 U10567 ( .A1(n9117), .A2(n9469), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9116), .ZN(n9118) );
  AOI211_X1 U10568 ( .C1(n9134), .C2(n9654), .A(n9119), .B(n9118), .ZN(n9120)
         );
  OAI211_X1 U10569 ( .C1(n9621), .C2(n9151), .A(n9121), .B(n9120), .ZN(
        P1_U3227) );
  NAND2_X1 U10570 ( .A1(n9124), .A2(n9123), .ZN(n9125) );
  XNOR2_X1 U10571 ( .A(n9122), .B(n9125), .ZN(n9130) );
  AOI22_X1 U10572 ( .A1(n9653), .A2(n10469), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9127) );
  NAND2_X1 U10573 ( .A1(n9714), .A2(n9134), .ZN(n9126) );
  OAI211_X1 U10574 ( .C1(n9158), .C2(n9685), .A(n9127), .B(n9126), .ZN(n9128)
         );
  AOI21_X1 U10575 ( .B1(n9833), .B2(n9165), .A(n9128), .ZN(n9129) );
  OAI21_X1 U10576 ( .B1(n9130), .B2(n9139), .A(n9129), .ZN(P1_U3231) );
  NAND2_X1 U10577 ( .A1(n9131), .A2(n4484), .ZN(n9132) );
  XOR2_X1 U10578 ( .A(n9133), .B(n9132), .Z(n9140) );
  AOI22_X1 U10579 ( .A1(n9653), .A2(n9134), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9136) );
  NAND2_X1 U10580 ( .A1(n10469), .A2(n9654), .ZN(n9135) );
  OAI211_X1 U10581 ( .C1(n9158), .C2(n9648), .A(n9136), .B(n9135), .ZN(n9137)
         );
  AOI21_X1 U10582 ( .B1(n9821), .B2(n9165), .A(n9137), .ZN(n9138) );
  OAI21_X1 U10583 ( .B1(n9140), .B2(n9139), .A(n9138), .ZN(P1_U3233) );
  OAI21_X1 U10584 ( .B1(n9085), .B2(n9143), .A(n9142), .ZN(n9144) );
  NAND3_X1 U10585 ( .A1(n9145), .A2(n9152), .A3(n9144), .ZN(n9150) );
  INV_X1 U10586 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9146) );
  OAI22_X1 U10587 ( .A1(n9469), .A2(n9161), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9146), .ZN(n9148) );
  NOR2_X1 U10588 ( .A1(n9158), .A2(n9588), .ZN(n9147) );
  AOI211_X1 U10589 ( .C1(n10469), .C2(n9595), .A(n9148), .B(n9147), .ZN(n9149)
         );
  OAI211_X1 U10590 ( .C1(n9591), .C2(n9151), .A(n9150), .B(n9149), .ZN(
        P1_U3238) );
  INV_X1 U10591 ( .A(n9157), .ZN(n9154) );
  OAI21_X1 U10592 ( .B1(n9154), .B2(n9153), .A(n9152), .ZN(n9168) );
  AOI21_X1 U10593 ( .B1(n9157), .B2(n9156), .A(n9155), .ZN(n9167) );
  NOR2_X1 U10594 ( .A1(n9158), .A2(n9777), .ZN(n9164) );
  NAND2_X1 U10595 ( .A1(n9730), .A2(n10469), .ZN(n9160) );
  NAND2_X1 U10596 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10136)
         );
  OAI211_X1 U10597 ( .C1(n9162), .C2(n9161), .A(n9160), .B(n10136), .ZN(n9163)
         );
  AOI211_X1 U10598 ( .C1(n9858), .C2(n9165), .A(n9164), .B(n9163), .ZN(n9166)
         );
  OAI21_X1 U10599 ( .B1(n9168), .B2(n9167), .A(n9166), .ZN(P1_U3239) );
  OR2_X1 U10600 ( .A1(n9173), .A2(n6768), .ZN(n9170) );
  INV_X1 U10601 ( .A(n9540), .ZN(n9247) );
  NAND2_X1 U10602 ( .A1(n9783), .A2(n9247), .ZN(n9442) );
  NAND2_X1 U10603 ( .A1(n9171), .A2(n5368), .ZN(n9175) );
  OR2_X1 U10604 ( .A1(n9173), .A2(n9172), .ZN(n9174) );
  INV_X1 U10605 ( .A(n9466), .ZN(n9236) );
  OR2_X1 U10606 ( .A1(n9993), .A2(n9236), .ZN(n9292) );
  NAND2_X1 U10607 ( .A1(n9442), .A2(n9292), .ZN(n9288) );
  NAND2_X1 U10608 ( .A1(n9414), .A2(n9410), .ZN(n9318) );
  INV_X1 U10609 ( .A(n9255), .ZN(n9176) );
  NAND2_X1 U10610 ( .A1(n9176), .A2(n9393), .ZN(n9382) );
  INV_X1 U10611 ( .A(n9382), .ZN(n9179) );
  AND2_X1 U10612 ( .A1(n9396), .A2(n9180), .ZN(n9386) );
  INV_X1 U10613 ( .A(n9386), .ZN(n9178) );
  INV_X1 U10614 ( .A(n9392), .ZN(n9177) );
  NOR2_X1 U10615 ( .A1(n9398), .A2(n9177), .ZN(n9387) );
  OAI211_X1 U10616 ( .C1(n9179), .C2(n9178), .A(n9387), .B(n9399), .ZN(n9223)
         );
  NAND2_X1 U10617 ( .A1(n9180), .A2(n9253), .ZN(n9381) );
  INV_X1 U10618 ( .A(n9377), .ZN(n9200) );
  NAND2_X1 U10619 ( .A1(n9190), .A2(n4530), .ZN(n9367) );
  INV_X1 U10620 ( .A(n9367), .ZN(n9197) );
  NAND2_X1 U10621 ( .A1(n9345), .A2(n4516), .ZN(n9358) );
  OR2_X1 U10622 ( .A1(n9358), .A2(n4797), .ZN(n9195) );
  NAND2_X1 U10623 ( .A1(n9182), .A2(n9343), .ZN(n9348) );
  INV_X1 U10624 ( .A(n9348), .ZN(n9931) );
  AND2_X1 U10625 ( .A1(n9351), .A2(n9931), .ZN(n9186) );
  INV_X1 U10626 ( .A(n9345), .ZN(n9183) );
  NOR2_X1 U10627 ( .A1(n9184), .A2(n9183), .ZN(n9360) );
  INV_X1 U10628 ( .A(n9360), .ZN(n9185) );
  OAI21_X1 U10629 ( .B1(n9195), .B2(n9186), .A(n9185), .ZN(n9187) );
  NAND2_X1 U10630 ( .A1(n9197), .A2(n9187), .ZN(n9191) );
  OR2_X1 U10631 ( .A1(n9869), .A2(n9188), .ZN(n9189) );
  NAND2_X1 U10632 ( .A1(n9761), .A2(n9189), .ZN(n9361) );
  NAND2_X1 U10633 ( .A1(n9361), .A2(n9190), .ZN(n9369) );
  NAND2_X1 U10634 ( .A1(n9191), .A2(n9369), .ZN(n9192) );
  NAND2_X1 U10635 ( .A1(n9192), .A2(n9373), .ZN(n9193) );
  AND3_X1 U10636 ( .A1(n9378), .A2(n9193), .A3(n9374), .ZN(n9194) );
  OR3_X1 U10637 ( .A1(n9381), .A2(n9200), .A3(n9194), .ZN(n9226) );
  INV_X1 U10638 ( .A(n9195), .ZN(n9198) );
  AND2_X1 U10639 ( .A1(n9349), .A2(n9335), .ZN(n9196) );
  NAND4_X1 U10640 ( .A1(n9373), .A2(n9198), .A3(n9197), .A4(n9196), .ZN(n9199)
         );
  OR3_X1 U10641 ( .A1(n9381), .A2(n9200), .A3(n9199), .ZN(n9201) );
  NAND2_X1 U10642 ( .A1(n9226), .A2(n9201), .ZN(n9202) );
  AND2_X1 U10643 ( .A1(n9202), .A2(n9396), .ZN(n9205) );
  NAND2_X1 U10644 ( .A1(n9399), .A2(n9395), .ZN(n9203) );
  AND2_X1 U10645 ( .A1(n9203), .A2(n9401), .ZN(n9204) );
  AND2_X1 U10646 ( .A1(n9402), .A2(n9204), .ZN(n9390) );
  OAI21_X1 U10647 ( .B1(n9223), .B2(n9205), .A(n9390), .ZN(n9206) );
  NAND2_X1 U10648 ( .A1(n9206), .A2(n9404), .ZN(n9207) );
  AND2_X1 U10649 ( .A1(n9207), .A2(n9409), .ZN(n9208) );
  NOR2_X1 U10650 ( .A1(n9412), .A2(n9208), .ZN(n9209) );
  NOR2_X1 U10651 ( .A1(n9318), .A2(n9209), .ZN(n9303) );
  INV_X1 U10652 ( .A(n9210), .ZN(n9212) );
  NAND2_X1 U10653 ( .A1(n9480), .A2(n10185), .ZN(n9211) );
  NAND3_X1 U10654 ( .A1(n9212), .A2(n9453), .A3(n9211), .ZN(n9213) );
  NAND2_X1 U10655 ( .A1(n9213), .A2(n7218), .ZN(n9215) );
  OAI21_X1 U10656 ( .B1(n9216), .B2(n9215), .A(n9214), .ZN(n9222) );
  INV_X1 U10657 ( .A(n9217), .ZN(n9331) );
  NAND2_X1 U10658 ( .A1(n9331), .A2(n9218), .ZN(n9298) );
  INV_X1 U10659 ( .A(n9298), .ZN(n9221) );
  AND2_X1 U10660 ( .A1(n9330), .A2(n9219), .ZN(n9301) );
  INV_X1 U10661 ( .A(n9301), .ZN(n9220) );
  AOI22_X1 U10662 ( .A1(n9222), .A2(n9221), .B1(n9331), .B2(n9220), .ZN(n9231)
         );
  INV_X1 U10663 ( .A(n9223), .ZN(n9228) );
  AND2_X1 U10664 ( .A1(n9339), .A2(n9224), .ZN(n9329) );
  INV_X1 U10665 ( .A(n9329), .ZN(n9225) );
  AOI21_X1 U10666 ( .B1(n4783), .B2(n9336), .A(n9225), .ZN(n9227) );
  NAND4_X1 U10667 ( .A1(n9228), .A2(n9227), .A3(n9404), .A4(n9226), .ZN(n9229)
         );
  OR2_X1 U10668 ( .A1(n9412), .A2(n9229), .ZN(n9304) );
  INV_X1 U10669 ( .A(n9304), .ZN(n9230) );
  OAI21_X1 U10670 ( .B1(n4781), .B2(n9231), .A(n9230), .ZN(n9232) );
  AND2_X1 U10671 ( .A1(n9303), .A2(n9232), .ZN(n9245) );
  NAND2_X1 U10672 ( .A1(n9313), .A2(n9426), .ZN(n9243) );
  INV_X1 U10673 ( .A(n9423), .ZN(n9234) );
  INV_X1 U10674 ( .A(n9419), .ZN(n9233) );
  OR4_X1 U10675 ( .A1(n9243), .A2(n9235), .A3(n9234), .A4(n9233), .ZN(n9295)
         );
  NAND2_X1 U10676 ( .A1(n9993), .A2(n9236), .ZN(n9286) );
  AND2_X1 U10677 ( .A1(n9238), .A2(n9237), .ZN(n9428) );
  INV_X1 U10678 ( .A(n9428), .ZN(n9241) );
  AND2_X1 U10679 ( .A1(n9423), .A2(n9239), .ZN(n9240) );
  NOR2_X1 U10680 ( .A1(n9241), .A2(n9240), .ZN(n9242) );
  OR2_X1 U10681 ( .A1(n9243), .A2(n9242), .ZN(n9244) );
  AND2_X1 U10682 ( .A1(n9244), .A2(n9432), .ZN(n9309) );
  OAI211_X1 U10683 ( .C1(n9245), .C2(n9295), .A(n9286), .B(n9309), .ZN(n9246)
         );
  INV_X1 U10684 ( .A(n9246), .ZN(n9248) );
  OAI21_X1 U10685 ( .B1(n9288), .B2(n9248), .A(n9451), .ZN(n9249) );
  XNOR2_X1 U10686 ( .A(n9249), .B(n10180), .ZN(n9457) );
  INV_X1 U10687 ( .A(n9451), .ZN(n9289) );
  INV_X1 U10688 ( .A(n9434), .ZN(n9285) );
  INV_X1 U10689 ( .A(n9552), .ZN(n9554) );
  INV_X1 U10690 ( .A(n9250), .ZN(n9252) );
  NAND2_X1 U10691 ( .A1(n9404), .A2(n9402), .ZN(n9652) );
  INV_X1 U10692 ( .A(n9660), .ZN(n9664) );
  NOR2_X1 U10693 ( .A1(n9398), .A2(n9395), .ZN(n9679) );
  INV_X1 U10694 ( .A(n9253), .ZN(n9254) );
  OR2_X1 U10695 ( .A1(n9255), .A2(n9254), .ZN(n9728) );
  INV_X1 U10696 ( .A(n9763), .ZN(n9371) );
  INV_X1 U10697 ( .A(n9256), .ZN(n9257) );
  NAND4_X1 U10698 ( .A1(n9260), .A2(n9259), .A3(n9258), .A4(n9257), .ZN(n9263)
         );
  NOR4_X1 U10699 ( .A1(n9263), .A2(n9262), .A3(n9261), .A4(n9325), .ZN(n9268)
         );
  INV_X1 U10700 ( .A(n9264), .ZN(n9265) );
  NAND4_X1 U10701 ( .A1(n9268), .A2(n9267), .A3(n9266), .A4(n9265), .ZN(n9269)
         );
  OR3_X1 U10702 ( .A1(n9270), .A2(n9934), .A3(n9269), .ZN(n9272) );
  NOR2_X1 U10703 ( .A1(n9272), .A2(n9271), .ZN(n9274) );
  NAND4_X1 U10704 ( .A1(n9371), .A2(n9275), .A3(n9274), .A4(n9273), .ZN(n9276)
         );
  OR3_X1 U10705 ( .A1(n9728), .A2(n5009), .A3(n9276), .ZN(n9277) );
  NOR2_X1 U10706 ( .A1(n9706), .A2(n9277), .ZN(n9278) );
  NAND4_X1 U10707 ( .A1(n9664), .A2(n9679), .A3(n9699), .A4(n9278), .ZN(n9279)
         );
  NOR2_X1 U10708 ( .A1(n9652), .A2(n9279), .ZN(n9280) );
  NAND3_X1 U10709 ( .A1(n9624), .A2(n8090), .A3(n9280), .ZN(n9281) );
  NOR2_X1 U10710 ( .A1(n9281), .A2(n9609), .ZN(n9282) );
  NAND2_X1 U10711 ( .A1(n9594), .A2(n9282), .ZN(n9283) );
  NOR2_X1 U10712 ( .A1(n9579), .A2(n9283), .ZN(n9284) );
  NAND4_X1 U10713 ( .A1(n9286), .A2(n9285), .A3(n9554), .A4(n9284), .ZN(n9287)
         );
  OR3_X1 U10714 ( .A1(n9289), .A2(n9288), .A3(n9287), .ZN(n9291) );
  NAND2_X1 U10715 ( .A1(n9291), .A2(n9290), .ZN(n9447) );
  NAND2_X1 U10716 ( .A1(n9292), .A2(n9540), .ZN(n9293) );
  NAND2_X1 U10717 ( .A1(n9293), .A2(n9783), .ZN(n9437) );
  NAND2_X1 U10718 ( .A1(n9540), .A2(n9466), .ZN(n9294) );
  NAND2_X1 U10719 ( .A1(n9993), .A2(n9294), .ZN(n9439) );
  INV_X1 U10720 ( .A(n9295), .ZN(n9307) );
  NAND2_X1 U10721 ( .A1(n9297), .A2(n9296), .ZN(n9322) );
  NAND2_X1 U10722 ( .A1(n9298), .A2(n9322), .ZN(n9299) );
  NAND2_X1 U10723 ( .A1(n9299), .A2(n9336), .ZN(n9300) );
  AOI21_X1 U10724 ( .B1(n9302), .B2(n9301), .A(n9300), .ZN(n9305) );
  OAI21_X1 U10725 ( .B1(n9305), .B2(n9304), .A(n9303), .ZN(n9306) );
  NAND2_X1 U10726 ( .A1(n9307), .A2(n9306), .ZN(n9308) );
  NAND3_X1 U10727 ( .A1(n9439), .A2(n9309), .A3(n9308), .ZN(n9310) );
  NAND2_X1 U10728 ( .A1(n9437), .A2(n9310), .ZN(n9311) );
  NAND3_X1 U10729 ( .A1(n9311), .A2(n9453), .A3(n9451), .ZN(n9312) );
  AND2_X1 U10730 ( .A1(n9447), .A2(n9312), .ZN(n9450) );
  NAND2_X1 U10731 ( .A1(n9437), .A2(n9313), .ZN(n9314) );
  NAND2_X1 U10732 ( .A1(n9314), .A2(n9440), .ZN(n9438) );
  INV_X1 U10733 ( .A(n9579), .ZN(n9422) );
  INV_X1 U10734 ( .A(n9409), .ZN(n9315) );
  AND2_X1 U10735 ( .A1(n9316), .A2(n9315), .ZN(n9317) );
  OR2_X1 U10736 ( .A1(n9318), .A2(n9317), .ZN(n9321) );
  NAND2_X1 U10737 ( .A1(n9319), .A2(n9415), .ZN(n9320) );
  MUX2_X1 U10738 ( .A(n9321), .B(n9320), .S(n9440), .Z(n9418) );
  INV_X1 U10739 ( .A(n9440), .ZN(n9406) );
  NAND2_X1 U10740 ( .A1(n9322), .A2(n9406), .ZN(n9323) );
  INV_X1 U10741 ( .A(n9325), .ZN(n9326) );
  NAND2_X1 U10742 ( .A1(n9327), .A2(n9326), .ZN(n9338) );
  AOI21_X1 U10743 ( .B1(n9338), .B2(n9329), .A(n9328), .ZN(n9341) );
  NAND2_X1 U10744 ( .A1(n7403), .A2(n9330), .ZN(n9332) );
  NAND2_X1 U10745 ( .A1(n9332), .A2(n9331), .ZN(n9334) );
  NAND2_X1 U10746 ( .A1(n9334), .A2(n9333), .ZN(n9337) );
  OAI211_X1 U10747 ( .C1(n9338), .C2(n9337), .A(n9336), .B(n9335), .ZN(n9340)
         );
  NAND2_X1 U10748 ( .A1(n9929), .A2(n9349), .ZN(n9342) );
  AOI21_X1 U10749 ( .B1(n9350), .B2(n9343), .A(n9342), .ZN(n9347) );
  OAI211_X1 U10750 ( .C1(n9347), .C2(n9346), .A(n9345), .B(n9344), .ZN(n9355)
         );
  AOI21_X1 U10751 ( .B1(n9350), .B2(n9349), .A(n9348), .ZN(n9353) );
  OAI21_X1 U10752 ( .B1(n9353), .B2(n9352), .A(n9351), .ZN(n9354) );
  NAND2_X1 U10753 ( .A1(n9357), .A2(n9356), .ZN(n9365) );
  AND2_X1 U10754 ( .A1(n9358), .A2(n9357), .ZN(n9359) );
  NOR2_X1 U10755 ( .A1(n9367), .A2(n9359), .ZN(n9363) );
  NOR2_X1 U10756 ( .A1(n9361), .A2(n9360), .ZN(n9362) );
  MUX2_X1 U10757 ( .A(n9363), .B(n9362), .S(n9440), .Z(n9364) );
  NAND2_X1 U10758 ( .A1(n9367), .A2(n9761), .ZN(n9368) );
  MUX2_X1 U10759 ( .A(n9369), .B(n9368), .S(n9440), .Z(n9370) );
  NAND3_X1 U10760 ( .A1(n9372), .A2(n9371), .A3(n9370), .ZN(n9376) );
  MUX2_X1 U10761 ( .A(n9374), .B(n9373), .S(n9406), .Z(n9375) );
  NAND3_X1 U10762 ( .A1(n9376), .A2(n9738), .A3(n9375), .ZN(n9380) );
  INV_X1 U10763 ( .A(n9728), .ZN(n9721) );
  MUX2_X1 U10764 ( .A(n9378), .B(n9377), .S(n9440), .Z(n9379) );
  NAND3_X1 U10765 ( .A1(n9380), .A2(n9721), .A3(n9379), .ZN(n9385) );
  MUX2_X1 U10766 ( .A(n9382), .B(n9381), .S(n9406), .Z(n9383) );
  INV_X1 U10767 ( .A(n9383), .ZN(n9384) );
  NAND2_X1 U10768 ( .A1(n9385), .A2(n9384), .ZN(n9394) );
  NAND2_X1 U10769 ( .A1(n9394), .A2(n9386), .ZN(n9388) );
  NAND3_X1 U10770 ( .A1(n9388), .A2(n9387), .A3(n9399), .ZN(n9391) );
  INV_X1 U10771 ( .A(n9404), .ZN(n9389) );
  AOI21_X1 U10772 ( .B1(n9391), .B2(n9390), .A(n9389), .ZN(n9408) );
  NAND3_X1 U10773 ( .A1(n9394), .A2(n9393), .A3(n9392), .ZN(n9397) );
  NAND3_X1 U10774 ( .A1(n9397), .A2(n9396), .A3(n8084), .ZN(n9400) );
  INV_X1 U10775 ( .A(n9398), .ZN(n9661) );
  INV_X1 U10776 ( .A(n9402), .ZN(n9403) );
  AOI21_X1 U10777 ( .B1(n9405), .B2(n9404), .A(n9403), .ZN(n9407) );
  NAND2_X1 U10778 ( .A1(n9410), .A2(n9409), .ZN(n9411) );
  OR2_X1 U10779 ( .A1(n9412), .A2(n9411), .ZN(n9413) );
  MUX2_X1 U10780 ( .A(n9415), .B(n9414), .S(n9440), .Z(n9416) );
  OAI211_X1 U10781 ( .C1(n9418), .C2(n9417), .A(n9594), .B(n9416), .ZN(n9421)
         );
  MUX2_X1 U10782 ( .A(n9577), .B(n9419), .S(n9440), .Z(n9420) );
  NAND3_X1 U10783 ( .A1(n9422), .A2(n9421), .A3(n9420), .ZN(n9429) );
  AND2_X1 U10784 ( .A1(n9426), .A2(n9423), .ZN(n9425) );
  AOI21_X1 U10785 ( .B1(n9429), .B2(n9425), .A(n9424), .ZN(n9431) );
  INV_X1 U10786 ( .A(n9426), .ZN(n9427) );
  AOI21_X1 U10787 ( .B1(n9429), .B2(n9428), .A(n9427), .ZN(n9430) );
  OR2_X1 U10788 ( .A1(n9432), .A2(n9440), .ZN(n9433) );
  OAI211_X1 U10789 ( .C1(n9435), .C2(n9434), .A(n9439), .B(n9433), .ZN(n9436)
         );
  INV_X1 U10790 ( .A(n9439), .ZN(n9441) );
  NAND3_X1 U10791 ( .A1(n9442), .A2(n9441), .A3(n9440), .ZN(n9443) );
  AND2_X1 U10792 ( .A1(n9443), .A2(n9451), .ZN(n9444) );
  NAND2_X1 U10793 ( .A1(n9445), .A2(n9444), .ZN(n9454) );
  INV_X1 U10794 ( .A(n9446), .ZN(n9448) );
  OAI21_X1 U10795 ( .B1(n9454), .B2(n9448), .A(n9447), .ZN(n9449) );
  OR2_X1 U10796 ( .A1(n9459), .A2(n9458), .ZN(n9460) );
  NOR2_X1 U10797 ( .A1(n9461), .A2(n9460), .ZN(n9464) );
  OAI21_X1 U10798 ( .B1(n9465), .B2(n9462), .A(P1_B_REG_SCAN_IN), .ZN(n9463)
         );
  MUX2_X1 U10799 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9466), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10800 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9467), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10801 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n8072), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10802 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9595), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10803 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9468), .S(P1_U4006), .Z(
        P1_U3581) );
  INV_X1 U10804 ( .A(n9469), .ZN(n9625) );
  MUX2_X1 U10805 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9625), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10806 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9642), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10807 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9654), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10808 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9666), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10809 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9653), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10810 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9701), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10811 ( .A(n9714), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9479), .Z(
        P1_U3574) );
  MUX2_X1 U10812 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9731), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10813 ( .A(n9715), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9479), .Z(
        P1_U3572) );
  MUX2_X1 U10814 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9730), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10815 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9470), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10816 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9767), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10817 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9471), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10818 ( .A(n9936), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9479), .Z(
        P1_U3566) );
  MUX2_X1 U10819 ( .A(n9937), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9479), .Z(
        P1_U3564) );
  MUX2_X1 U10820 ( .A(n9472), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9479), .Z(
        P1_U3563) );
  MUX2_X1 U10821 ( .A(n9473), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9479), .Z(
        P1_U3562) );
  MUX2_X1 U10822 ( .A(n9474), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9479), .Z(
        P1_U3561) );
  MUX2_X1 U10823 ( .A(n9475), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9479), .Z(
        P1_U3560) );
  MUX2_X1 U10824 ( .A(n9476), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9479), .Z(
        P1_U3559) );
  MUX2_X1 U10825 ( .A(n9477), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9479), .Z(
        P1_U3558) );
  MUX2_X1 U10826 ( .A(n9478), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9479), .Z(
        P1_U3557) );
  MUX2_X1 U10827 ( .A(n9480), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9479), .Z(
        P1_U3556) );
  OAI21_X1 U10828 ( .B1(n10085), .B2(n9483), .A(n9481), .ZN(n9482) );
  AOI21_X1 U10829 ( .B1(n10041), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n9482), .ZN(
        n9494) );
  INV_X1 U10830 ( .A(n10131), .ZN(n10170) );
  MUX2_X1 U10831 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6797), .S(n9483), .Z(n9486)
         );
  NAND3_X1 U10832 ( .A1(n9486), .A2(n9485), .A3(n9484), .ZN(n9487) );
  NAND3_X1 U10833 ( .A1(n10170), .A2(n9488), .A3(n9487), .ZN(n9493) );
  OAI211_X1 U10834 ( .C1(n9491), .C2(n9490), .A(n10088), .B(n9489), .ZN(n9492)
         );
  NAND3_X1 U10835 ( .A1(n9494), .A2(n9493), .A3(n9492), .ZN(P1_U3244) );
  AOI22_X1 U10836 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n9527), .B1(n9523), .B2(
        n9526), .ZN(n9504) );
  XNOR2_X1 U10837 ( .A(n9502), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10172) );
  INV_X1 U10838 ( .A(n10153), .ZN(n9500) );
  XOR2_X1 U10839 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10153), .Z(n10155) );
  AOI21_X1 U10840 ( .B1(n9505), .B2(n9496), .A(n9495), .ZN(n9497) );
  NAND2_X1 U10841 ( .A1(n10141), .A2(n9497), .ZN(n9498) );
  XNOR2_X1 U10842 ( .A(n9497), .B(n9510), .ZN(n10143) );
  NAND2_X1 U10843 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n10143), .ZN(n10142) );
  NAND2_X1 U10844 ( .A1(n9498), .A2(n10142), .ZN(n10156) );
  NAND2_X1 U10845 ( .A1(n10155), .A2(n10156), .ZN(n10154) );
  OAI21_X1 U10846 ( .B1(n9500), .B2(n9499), .A(n10154), .ZN(n10171) );
  NAND2_X1 U10847 ( .A1(n10172), .A2(n10171), .ZN(n10169) );
  OAI21_X1 U10848 ( .B1(n9502), .B2(n9501), .A(n10169), .ZN(n9503) );
  NOR2_X1 U10849 ( .A1(n9504), .A2(n9503), .ZN(n9525) );
  AOI21_X1 U10850 ( .B1(n9504), .B2(n9503), .A(n9525), .ZN(n9521) );
  NAND2_X1 U10851 ( .A1(n9506), .A2(n9505), .ZN(n9508) );
  NAND2_X1 U10852 ( .A1(n9508), .A2(n9507), .ZN(n9509) );
  NOR2_X1 U10853 ( .A1(n9510), .A2(n9509), .ZN(n9511) );
  XNOR2_X1 U10854 ( .A(n9510), .B(n9509), .ZN(n10138) );
  NOR2_X1 U10855 ( .A1(n9778), .A2(n10138), .ZN(n10137) );
  NAND2_X1 U10856 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n10153), .ZN(n9512) );
  OAI21_X1 U10857 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n10153), .A(n9512), .ZN(
        n10149) );
  NOR2_X1 U10858 ( .A1(n10150), .A2(n10149), .ZN(n10148) );
  NAND2_X1 U10859 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n10167), .ZN(n9513) );
  OAI21_X1 U10860 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n10167), .A(n9513), .ZN(
        n10163) );
  NOR2_X1 U10861 ( .A1(n10164), .A2(n10163), .ZN(n10162) );
  AOI22_X1 U10862 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n9527), .B1(n9523), .B2(
        n9709), .ZN(n9514) );
  NOR2_X1 U10863 ( .A1(n9515), .A2(n9514), .ZN(n9522) );
  AOI211_X1 U10864 ( .C1(n9515), .C2(n9514), .A(n9522), .B(n10161), .ZN(n9516)
         );
  INV_X1 U10865 ( .A(n9516), .ZN(n9520) );
  OAI21_X1 U10866 ( .B1(n10085), .B2(n9527), .A(n9517), .ZN(n9518) );
  AOI21_X1 U10867 ( .B1(n10041), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9518), .ZN(
        n9519) );
  OAI211_X1 U10868 ( .C1(n9521), .C2(n10131), .A(n9520), .B(n9519), .ZN(
        P1_U3259) );
  XNOR2_X1 U10869 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9524), .ZN(n9534) );
  INV_X1 U10870 ( .A(n9534), .ZN(n9530) );
  AOI21_X1 U10871 ( .B1(n9527), .B2(n9526), .A(n9525), .ZN(n9529) );
  INV_X1 U10872 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9528) );
  XOR2_X1 U10873 ( .A(n9529), .B(n9528), .Z(n9531) );
  OAI22_X1 U10874 ( .A1(n9530), .A2(n10161), .B1(n9531), .B2(n10131), .ZN(
        n9536) );
  AOI21_X1 U10875 ( .B1(n9531), .B2(n10170), .A(n10168), .ZN(n9532) );
  OAI21_X1 U10876 ( .B1(n9534), .B2(n9533), .A(n9532), .ZN(n9535) );
  INV_X1 U10877 ( .A(n9993), .ZN(n9545) );
  XNOR2_X1 U10878 ( .A(n9543), .B(n9783), .ZN(n9785) );
  NOR2_X1 U10879 ( .A1(n9774), .A2(n9538), .ZN(n9541) );
  NAND2_X1 U10880 ( .A1(n9540), .A2(n9539), .ZN(n9989) );
  NOR2_X1 U10881 ( .A1(n10193), .A2(n9989), .ZN(n9547) );
  AOI211_X1 U10882 ( .C1(n9783), .C2(n9947), .A(n9541), .B(n9547), .ZN(n9542)
         );
  OAI21_X1 U10883 ( .B1(n9785), .B2(n9550), .A(n9542), .ZN(P1_U3261) );
  OAI21_X1 U10884 ( .B1(n9545), .B2(n9544), .A(n9543), .ZN(n9990) );
  NOR2_X1 U10885 ( .A1(n9774), .A2(n9546), .ZN(n9548) );
  AOI211_X1 U10886 ( .C1(n9993), .C2(n9947), .A(n9548), .B(n9547), .ZN(n9549)
         );
  OAI21_X1 U10887 ( .B1(n9990), .B2(n9550), .A(n9549), .ZN(P1_U3262) );
  OAI21_X1 U10888 ( .B1(n9553), .B2(n9552), .A(n9551), .ZN(n9795) );
  XNOR2_X1 U10889 ( .A(n9555), .B(n9554), .ZN(n9559) );
  OAI22_X1 U10890 ( .A1(n9557), .A2(n9751), .B1(n9556), .B2(n9769), .ZN(n9558)
         );
  AOI21_X1 U10891 ( .B1(n9559), .B2(n9772), .A(n9558), .ZN(n9794) );
  OAI22_X1 U10892 ( .A1(n9774), .A2(n9561), .B1(n9560), .B2(n10187), .ZN(n9562) );
  AOI21_X1 U10893 ( .B1(n9791), .B2(n9947), .A(n9562), .ZN(n9567) );
  OR2_X1 U10894 ( .A1(n9563), .A2(n9571), .ZN(n9565) );
  NAND2_X1 U10895 ( .A1(n9792), .A2(n9735), .ZN(n9566) );
  OAI211_X1 U10896 ( .C1(n9794), .C2(n10193), .A(n9567), .B(n9566), .ZN(n9568)
         );
  INV_X1 U10897 ( .A(n9568), .ZN(n9569) );
  OAI21_X1 U10898 ( .B1(n9795), .B2(n9755), .A(n9569), .ZN(P1_U3263) );
  XOR2_X1 U10899 ( .A(n9579), .B(n9570), .Z(n9800) );
  INV_X1 U10900 ( .A(n9587), .ZN(n9572) );
  AOI21_X1 U10901 ( .B1(n9796), .B2(n9572), .A(n9571), .ZN(n9797) );
  INV_X1 U10902 ( .A(n9573), .ZN(n9574) );
  AOI22_X1 U10903 ( .A1(n10193), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9574), 
        .B2(n9946), .ZN(n9575) );
  OAI21_X1 U10904 ( .B1(n9576), .B2(n9742), .A(n9575), .ZN(n9584) );
  NAND2_X1 U10905 ( .A1(n9592), .A2(n9577), .ZN(n9578) );
  AOI211_X1 U10906 ( .C1(n9579), .C2(n9578), .A(n9940), .B(n4514), .ZN(n9582)
         );
  OAI22_X1 U10907 ( .A1(n9611), .A2(n9751), .B1(n9580), .B2(n9769), .ZN(n9581)
         );
  NOR2_X1 U10908 ( .A1(n9582), .A2(n9581), .ZN(n9799) );
  NOR2_X1 U10909 ( .A1(n9799), .A2(n10193), .ZN(n9583) );
  AOI211_X1 U10910 ( .C1(n9735), .C2(n9797), .A(n9584), .B(n9583), .ZN(n9585)
         );
  OAI21_X1 U10911 ( .B1(n9800), .B2(n9755), .A(n9585), .ZN(P1_U3264) );
  XOR2_X1 U10912 ( .A(n9594), .B(n9586), .Z(n9805) );
  AOI211_X1 U10913 ( .C1(n9802), .C2(n9601), .A(n10239), .B(n9587), .ZN(n9801)
         );
  INV_X1 U10914 ( .A(n9588), .ZN(n9589) );
  AOI22_X1 U10915 ( .A1(n10193), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9589), 
        .B2(n9946), .ZN(n9590) );
  OAI21_X1 U10916 ( .B1(n9591), .B2(n9742), .A(n9590), .ZN(n9598) );
  OAI21_X1 U10917 ( .B1(n9594), .B2(n9593), .A(n9592), .ZN(n9596) );
  AOI222_X1 U10918 ( .A1(n9772), .A2(n9596), .B1(n9625), .B2(n9938), .C1(n9595), .C2(n9935), .ZN(n9804) );
  NOR2_X1 U10919 ( .A1(n9804), .A2(n10193), .ZN(n9597) );
  AOI211_X1 U10920 ( .C1(n9801), .C2(n9954), .A(n9598), .B(n9597), .ZN(n9599)
         );
  OAI21_X1 U10921 ( .B1(n9805), .B2(n9755), .A(n9599), .ZN(P1_U3265) );
  XOR2_X1 U10922 ( .A(n9600), .B(n9609), .Z(n9810) );
  INV_X1 U10923 ( .A(n9616), .ZN(n9602) );
  AOI211_X1 U10924 ( .C1(n9808), .C2(n9602), .A(n10239), .B(n4681), .ZN(n9807)
         );
  NOR2_X1 U10925 ( .A1(n9603), .A2(n9742), .ZN(n9607) );
  OAI22_X1 U10926 ( .A1(n9774), .A2(n9605), .B1(n9604), .B2(n10187), .ZN(n9606) );
  AOI211_X1 U10927 ( .C1(n9807), .C2(n9954), .A(n9607), .B(n9606), .ZN(n9614)
         );
  XOR2_X1 U10928 ( .A(n9609), .B(n9608), .Z(n9610) );
  OAI222_X1 U10929 ( .A1(n9751), .A2(n9612), .B1(n9769), .B2(n9611), .C1(n9940), .C2(n9610), .ZN(n9806) );
  NAND2_X1 U10930 ( .A1(n9806), .A2(n9774), .ZN(n9613) );
  OAI211_X1 U10931 ( .C1(n9810), .C2(n9755), .A(n9614), .B(n9613), .ZN(
        P1_U3266) );
  XOR2_X1 U10932 ( .A(n9615), .B(n9624), .Z(n9815) );
  INV_X1 U10933 ( .A(n9631), .ZN(n9617) );
  AOI21_X1 U10934 ( .B1(n9811), .B2(n9617), .A(n9616), .ZN(n9812) );
  INV_X1 U10935 ( .A(n9618), .ZN(n9619) );
  AOI22_X1 U10936 ( .A1(n10193), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9619), 
        .B2(n9946), .ZN(n9620) );
  OAI21_X1 U10937 ( .B1(n9621), .B2(n9742), .A(n9620), .ZN(n9628) );
  NAND2_X1 U10938 ( .A1(n9636), .A2(n9622), .ZN(n9623) );
  XOR2_X1 U10939 ( .A(n9624), .B(n9623), .Z(n9626) );
  AOI222_X1 U10940 ( .A1(n9772), .A2(n9626), .B1(n9654), .B2(n9938), .C1(n9625), .C2(n9935), .ZN(n9814) );
  NOR2_X1 U10941 ( .A1(n9814), .A2(n10193), .ZN(n9627) );
  AOI211_X1 U10942 ( .C1(n9812), .C2(n9735), .A(n9628), .B(n9627), .ZN(n9629)
         );
  OAI21_X1 U10943 ( .B1(n9815), .B2(n9755), .A(n9629), .ZN(P1_U3267) );
  XNOR2_X1 U10944 ( .A(n9630), .B(n9639), .ZN(n9820) );
  AOI21_X1 U10945 ( .B1(n9816), .B2(n9647), .A(n9631), .ZN(n9817) );
  INV_X1 U10946 ( .A(n9632), .ZN(n9633) );
  AOI22_X1 U10947 ( .A1(n10193), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9633), 
        .B2(n9946), .ZN(n9634) );
  OAI21_X1 U10948 ( .B1(n9635), .B2(n9742), .A(n9634), .ZN(n9644) );
  AND2_X1 U10949 ( .A1(n9666), .A2(n9938), .ZN(n9641) );
  INV_X1 U10950 ( .A(n9636), .ZN(n9637) );
  AOI211_X1 U10951 ( .C1(n9639), .C2(n9638), .A(n9940), .B(n9637), .ZN(n9640)
         );
  AOI211_X1 U10952 ( .C1(n9935), .C2(n9642), .A(n9641), .B(n9640), .ZN(n9819)
         );
  NOR2_X1 U10953 ( .A1(n9819), .A2(n10193), .ZN(n9643) );
  AOI211_X1 U10954 ( .C1(n9817), .C2(n9735), .A(n9644), .B(n9643), .ZN(n9645)
         );
  OAI21_X1 U10955 ( .B1(n9820), .B2(n9755), .A(n9645), .ZN(P1_U3268) );
  XOR2_X1 U10956 ( .A(n9646), .B(n9652), .Z(n9825) );
  AOI21_X1 U10957 ( .B1(n9821), .B2(n9668), .A(n4686), .ZN(n9822) );
  INV_X1 U10958 ( .A(n9648), .ZN(n9649) );
  AOI22_X1 U10959 ( .A1(n10193), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9649), 
        .B2(n9946), .ZN(n9650) );
  OAI21_X1 U10960 ( .B1(n4685), .B2(n9742), .A(n9650), .ZN(n9657) );
  XOR2_X1 U10961 ( .A(n9652), .B(n9651), .Z(n9655) );
  AOI222_X1 U10962 ( .A1(n9772), .A2(n9655), .B1(n9654), .B2(n9935), .C1(n9653), .C2(n9938), .ZN(n9824) );
  NOR2_X1 U10963 ( .A1(n9824), .A2(n10193), .ZN(n9656) );
  AOI211_X1 U10964 ( .C1(n9822), .C2(n9735), .A(n9657), .B(n9656), .ZN(n9658)
         );
  OAI21_X1 U10965 ( .B1(n9825), .B2(n9755), .A(n9658), .ZN(P1_U3269) );
  XNOR2_X1 U10966 ( .A(n9659), .B(n9660), .ZN(n9830) );
  AOI22_X1 U10967 ( .A1(n9827), .A2(n9947), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n10193), .ZN(n9676) );
  AND2_X1 U10968 ( .A1(n9662), .A2(n9661), .ZN(n9665) );
  OAI21_X1 U10969 ( .B1(n9665), .B2(n9664), .A(n9663), .ZN(n9667) );
  AOI222_X1 U10970 ( .A1(n9772), .A2(n9667), .B1(n9666), .B2(n9935), .C1(n9701), .C2(n9938), .ZN(n9829) );
  INV_X1 U10971 ( .A(n9683), .ZN(n9670) );
  INV_X1 U10972 ( .A(n9668), .ZN(n9669) );
  AOI211_X1 U10973 ( .C1(n9827), .C2(n9670), .A(n10239), .B(n9669), .ZN(n9826)
         );
  NAND2_X1 U10974 ( .A1(n9826), .A2(n9671), .ZN(n9672) );
  OAI211_X1 U10975 ( .C1(n10187), .C2(n9673), .A(n9829), .B(n9672), .ZN(n9674)
         );
  NAND2_X1 U10976 ( .A1(n9674), .A2(n9774), .ZN(n9675) );
  OAI211_X1 U10977 ( .C1(n9830), .C2(n9755), .A(n9676), .B(n9675), .ZN(
        P1_U3270) );
  XOR2_X1 U10978 ( .A(n9677), .B(n9679), .Z(n9835) );
  XOR2_X1 U10979 ( .A(n9679), .B(n9678), .Z(n9680) );
  OAI222_X1 U10980 ( .A1(n9769), .A2(n9682), .B1(n9751), .B2(n9681), .C1(n9680), .C2(n9940), .ZN(n9831) );
  INV_X1 U10981 ( .A(n9693), .ZN(n9684) );
  AOI211_X1 U10982 ( .C1(n9833), .C2(n9684), .A(n10239), .B(n9683), .ZN(n9832)
         );
  NAND2_X1 U10983 ( .A1(n9832), .A2(n9954), .ZN(n9688) );
  INV_X1 U10984 ( .A(n9685), .ZN(n9686) );
  AOI22_X1 U10985 ( .A1(n10193), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9686), 
        .B2(n9946), .ZN(n9687) );
  OAI211_X1 U10986 ( .C1(n9689), .C2(n9742), .A(n9688), .B(n9687), .ZN(n9690)
         );
  AOI21_X1 U10987 ( .B1(n9831), .B2(n9774), .A(n9690), .ZN(n9691) );
  OAI21_X1 U10988 ( .B1(n9835), .B2(n9755), .A(n9691), .ZN(P1_U3271) );
  XNOR2_X1 U10989 ( .A(n9692), .B(n9699), .ZN(n9840) );
  INV_X1 U10990 ( .A(n9708), .ZN(n9694) );
  AOI21_X1 U10991 ( .B1(n9836), .B2(n9694), .A(n9693), .ZN(n9837) );
  INV_X1 U10992 ( .A(n9695), .ZN(n9696) );
  AOI22_X1 U10993 ( .A1(n10193), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9696), 
        .B2(n9946), .ZN(n9697) );
  OAI21_X1 U10994 ( .B1(n9698), .B2(n9742), .A(n9697), .ZN(n9704) );
  XNOR2_X1 U10995 ( .A(n9700), .B(n9699), .ZN(n9702) );
  AOI222_X1 U10996 ( .A1(n9772), .A2(n9702), .B1(n9731), .B2(n9938), .C1(n9701), .C2(n9935), .ZN(n9839) );
  NOR2_X1 U10997 ( .A1(n9839), .A2(n10193), .ZN(n9703) );
  AOI211_X1 U10998 ( .C1(n9837), .C2(n9735), .A(n9704), .B(n9703), .ZN(n9705)
         );
  OAI21_X1 U10999 ( .B1(n9840), .B2(n9755), .A(n9705), .ZN(P1_U3272) );
  XNOR2_X1 U11000 ( .A(n9707), .B(n9706), .ZN(n9845) );
  AOI21_X1 U11001 ( .B1(n9841), .B2(n9723), .A(n9708), .ZN(n9842) );
  INV_X1 U11002 ( .A(n9841), .ZN(n9710) );
  OAI22_X1 U11003 ( .A1(n9710), .A2(n9742), .B1(n9709), .B2(n9774), .ZN(n9711)
         );
  AOI21_X1 U11004 ( .B1(n9842), .B2(n9735), .A(n9711), .ZN(n9720) );
  XNOR2_X1 U11005 ( .A(n9713), .B(n9712), .ZN(n9716) );
  AOI222_X1 U11006 ( .A1(n9772), .A2(n9716), .B1(n9715), .B2(n9938), .C1(n9714), .C2(n9935), .ZN(n9844) );
  OAI21_X1 U11007 ( .B1(n9717), .B2(n10187), .A(n9844), .ZN(n9718) );
  NAND2_X1 U11008 ( .A1(n9718), .A2(n9774), .ZN(n9719) );
  OAI211_X1 U11009 ( .C1(n9845), .C2(n9755), .A(n9720), .B(n9719), .ZN(
        P1_U3273) );
  XNOR2_X1 U11010 ( .A(n9722), .B(n9721), .ZN(n9850) );
  AOI21_X1 U11011 ( .B1(n9846), .B2(n9740), .A(n4693), .ZN(n9847) );
  INV_X1 U11012 ( .A(n9724), .ZN(n9725) );
  AOI22_X1 U11013 ( .A1(n10193), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9725), 
        .B2(n9946), .ZN(n9726) );
  OAI21_X1 U11014 ( .B1(n9727), .B2(n9742), .A(n9726), .ZN(n9734) );
  XNOR2_X1 U11015 ( .A(n9729), .B(n9728), .ZN(n9732) );
  AOI222_X1 U11016 ( .A1(n9772), .A2(n9732), .B1(n9731), .B2(n9935), .C1(n9730), .C2(n9938), .ZN(n9849) );
  NOR2_X1 U11017 ( .A1(n9849), .A2(n10193), .ZN(n9733) );
  AOI211_X1 U11018 ( .C1(n9847), .C2(n9735), .A(n9734), .B(n9733), .ZN(n9736)
         );
  OAI21_X1 U11019 ( .B1(n9850), .B2(n9755), .A(n9736), .ZN(P1_U3274) );
  AOI21_X1 U11020 ( .B1(n9738), .B2(n9737), .A(n4558), .ZN(n9739) );
  INV_X1 U11021 ( .A(n9739), .ZN(n9855) );
  INV_X1 U11022 ( .A(n9740), .ZN(n9741) );
  AOI211_X1 U11023 ( .C1(n9853), .C2(n9758), .A(n10239), .B(n9741), .ZN(n9852)
         );
  INV_X1 U11024 ( .A(n9853), .ZN(n9743) );
  NOR2_X1 U11025 ( .A1(n9743), .A2(n9742), .ZN(n9747) );
  OAI22_X1 U11026 ( .A1(n9774), .A2(n9745), .B1(n9744), .B2(n10187), .ZN(n9746) );
  AOI211_X1 U11027 ( .C1(n9852), .C2(n9954), .A(n9747), .B(n9746), .ZN(n9754)
         );
  XNOR2_X1 U11028 ( .A(n9748), .B(n5009), .ZN(n9749) );
  OAI222_X1 U11029 ( .A1(n9769), .A2(n9752), .B1(n9751), .B2(n9750), .C1(n9749), .C2(n9940), .ZN(n9851) );
  NAND2_X1 U11030 ( .A1(n9851), .A2(n9774), .ZN(n9753) );
  OAI211_X1 U11031 ( .C1(n9855), .C2(n9755), .A(n9754), .B(n9753), .ZN(
        P1_U3275) );
  XNOR2_X1 U11032 ( .A(n9756), .B(n9763), .ZN(n9861) );
  NOR2_X1 U11033 ( .A1(n9861), .A2(n9757), .ZN(n9776) );
  OAI211_X1 U11034 ( .C1(n9760), .C2(n9759), .A(n9950), .B(n9758), .ZN(n9856)
         );
  NAND2_X1 U11035 ( .A1(n9762), .A2(n9761), .ZN(n9764) );
  NAND2_X1 U11036 ( .A1(n9764), .A2(n9763), .ZN(n9766) );
  NAND2_X1 U11037 ( .A1(n9766), .A2(n9765), .ZN(n9773) );
  NAND2_X1 U11038 ( .A1(n9767), .A2(n9938), .ZN(n9768) );
  OAI21_X1 U11039 ( .B1(n9770), .B2(n9769), .A(n9768), .ZN(n9771) );
  AOI21_X1 U11040 ( .B1(n9773), .B2(n9772), .A(n9771), .ZN(n9860) );
  OAI21_X1 U11041 ( .B1(n10180), .B2(n9856), .A(n9860), .ZN(n9775) );
  OAI21_X1 U11042 ( .B1(n9776), .B2(n9775), .A(n9774), .ZN(n9781) );
  OAI22_X1 U11043 ( .A1(n9774), .A2(n9778), .B1(n9777), .B2(n10187), .ZN(n9779) );
  AOI21_X1 U11044 ( .B1(n9858), .B2(n9947), .A(n9779), .ZN(n9780) );
  OAI211_X1 U11045 ( .C1(n9861), .C2(n9782), .A(n9781), .B(n9780), .ZN(
        P1_U3276) );
  NAND2_X1 U11046 ( .A1(n9783), .A2(n9994), .ZN(n9784) );
  OAI211_X1 U11047 ( .C1(n9785), .C2(n10239), .A(n9989), .B(n9784), .ZN(n9876)
         );
  MUX2_X1 U11048 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9876), .S(n10255), .Z(
        P1_U3554) );
  AOI22_X1 U11049 ( .A1(n9787), .A2(n9950), .B1(n9994), .B2(n9786), .ZN(n9788)
         );
  MUX2_X1 U11050 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9877), .S(n10255), .Z(
        P1_U3552) );
  AOI22_X1 U11051 ( .A1(n9792), .A2(n9950), .B1(n9994), .B2(n9791), .ZN(n9793)
         );
  OAI211_X1 U11052 ( .C1(n9795), .C2(n9866), .A(n9794), .B(n9793), .ZN(n9878)
         );
  MUX2_X1 U11053 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9878), .S(n10255), .Z(
        P1_U3551) );
  AOI22_X1 U11054 ( .A1(n9797), .A2(n9950), .B1(n9994), .B2(n9796), .ZN(n9798)
         );
  OAI211_X1 U11055 ( .C1(n9800), .C2(n9866), .A(n9799), .B(n9798), .ZN(n9879)
         );
  MUX2_X1 U11056 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9879), .S(n10255), .Z(
        P1_U3550) );
  AOI21_X1 U11057 ( .B1(n9994), .B2(n9802), .A(n9801), .ZN(n9803) );
  OAI211_X1 U11058 ( .C1(n9805), .C2(n9866), .A(n9804), .B(n9803), .ZN(n9880)
         );
  MUX2_X1 U11059 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9880), .S(n10255), .Z(
        P1_U3549) );
  AOI211_X1 U11060 ( .C1(n9994), .C2(n9808), .A(n9807), .B(n9806), .ZN(n9809)
         );
  OAI21_X1 U11061 ( .B1(n9810), .B2(n9866), .A(n9809), .ZN(n9881) );
  MUX2_X1 U11062 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9881), .S(n10255), .Z(
        P1_U3548) );
  AOI22_X1 U11063 ( .A1(n9812), .A2(n9950), .B1(n9994), .B2(n9811), .ZN(n9813)
         );
  OAI211_X1 U11064 ( .C1(n9815), .C2(n9866), .A(n9814), .B(n9813), .ZN(n9882)
         );
  MUX2_X1 U11065 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9882), .S(n10255), .Z(
        P1_U3547) );
  AOI22_X1 U11066 ( .A1(n9817), .A2(n9950), .B1(n9994), .B2(n9816), .ZN(n9818)
         );
  OAI211_X1 U11067 ( .C1(n9820), .C2(n9866), .A(n9819), .B(n9818), .ZN(n9883)
         );
  MUX2_X1 U11068 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9883), .S(n10255), .Z(
        P1_U3546) );
  AOI22_X1 U11069 ( .A1(n9822), .A2(n9950), .B1(n9994), .B2(n9821), .ZN(n9823)
         );
  OAI211_X1 U11070 ( .C1(n9825), .C2(n9866), .A(n9824), .B(n9823), .ZN(n9884)
         );
  MUX2_X1 U11071 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9884), .S(n10255), .Z(
        P1_U3545) );
  AOI21_X1 U11072 ( .B1(n9994), .B2(n9827), .A(n9826), .ZN(n9828) );
  OAI211_X1 U11073 ( .C1(n9830), .C2(n9866), .A(n9829), .B(n9828), .ZN(n9885)
         );
  MUX2_X1 U11074 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9885), .S(n10255), .Z(
        P1_U3544) );
  AOI211_X1 U11075 ( .C1(n9994), .C2(n9833), .A(n9832), .B(n9831), .ZN(n9834)
         );
  OAI21_X1 U11076 ( .B1(n9835), .B2(n9866), .A(n9834), .ZN(n9886) );
  MUX2_X1 U11077 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9886), .S(n10255), .Z(
        P1_U3543) );
  AOI22_X1 U11078 ( .A1(n9837), .A2(n9950), .B1(n9994), .B2(n9836), .ZN(n9838)
         );
  OAI211_X1 U11079 ( .C1(n9840), .C2(n9866), .A(n9839), .B(n9838), .ZN(n9887)
         );
  MUX2_X1 U11080 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9887), .S(n10255), .Z(
        P1_U3542) );
  AOI22_X1 U11081 ( .A1(n9842), .A2(n9950), .B1(n9994), .B2(n9841), .ZN(n9843)
         );
  OAI211_X1 U11082 ( .C1(n9845), .C2(n9866), .A(n9844), .B(n9843), .ZN(n9888)
         );
  MUX2_X1 U11083 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9888), .S(n10255), .Z(
        P1_U3541) );
  AOI22_X1 U11084 ( .A1(n9847), .A2(n9950), .B1(n9994), .B2(n9846), .ZN(n9848)
         );
  OAI211_X1 U11085 ( .C1(n9850), .C2(n9866), .A(n9849), .B(n9848), .ZN(n9889)
         );
  MUX2_X1 U11086 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9889), .S(n10255), .Z(
        P1_U3540) );
  AOI211_X1 U11087 ( .C1(n9994), .C2(n9853), .A(n9852), .B(n9851), .ZN(n9854)
         );
  OAI21_X1 U11088 ( .B1(n9855), .B2(n9866), .A(n9854), .ZN(n9890) );
  MUX2_X1 U11089 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9890), .S(n10255), .Z(
        P1_U3539) );
  INV_X1 U11090 ( .A(n9856), .ZN(n9857) );
  AOI21_X1 U11091 ( .B1(n9994), .B2(n9858), .A(n9857), .ZN(n9859) );
  OAI211_X1 U11092 ( .C1(n9861), .C2(n9866), .A(n9860), .B(n9859), .ZN(n9891)
         );
  MUX2_X1 U11093 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9891), .S(n10255), .Z(
        P1_U3538) );
  AOI211_X1 U11094 ( .C1(n9994), .C2(n9864), .A(n9863), .B(n9862), .ZN(n9865)
         );
  OAI21_X1 U11095 ( .B1(n9867), .B2(n9866), .A(n9865), .ZN(n9892) );
  MUX2_X1 U11096 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9892), .S(n10255), .Z(
        P1_U3537) );
  INV_X1 U11097 ( .A(n9868), .ZN(n10244) );
  OAI22_X1 U11098 ( .A1(n9870), .A2(n10239), .B1(n4677), .B2(n10237), .ZN(
        n9871) );
  AOI21_X1 U11099 ( .B1(n9872), .B2(n10244), .A(n9871), .ZN(n9873) );
  NAND2_X1 U11100 ( .A1(n9874), .A2(n9873), .ZN(n9893) );
  MUX2_X1 U11101 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9893), .S(n10255), .Z(
        P1_U3536) );
  MUX2_X1 U11102 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9875), .S(n10255), .Z(
        P1_U3523) );
  MUX2_X1 U11103 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9876), .S(n10247), .Z(
        P1_U3522) );
  MUX2_X1 U11104 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9877), .S(n10247), .Z(
        P1_U3520) );
  MUX2_X1 U11105 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9878), .S(n10247), .Z(
        P1_U3519) );
  MUX2_X1 U11106 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9879), .S(n10247), .Z(
        P1_U3518) );
  MUX2_X1 U11107 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9880), .S(n10247), .Z(
        P1_U3517) );
  MUX2_X1 U11108 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9881), .S(n10247), .Z(
        P1_U3516) );
  MUX2_X1 U11109 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9882), .S(n10247), .Z(
        P1_U3515) );
  MUX2_X1 U11110 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9883), .S(n10247), .Z(
        P1_U3514) );
  MUX2_X1 U11111 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9884), .S(n10247), .Z(
        P1_U3513) );
  MUX2_X1 U11112 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9885), .S(n10247), .Z(
        P1_U3512) );
  MUX2_X1 U11113 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9886), .S(n10247), .Z(
        P1_U3511) );
  MUX2_X1 U11114 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9887), .S(n10247), .Z(
        P1_U3510) );
  MUX2_X1 U11115 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9888), .S(n10247), .Z(
        P1_U3508) );
  MUX2_X1 U11116 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9889), .S(n10247), .Z(
        P1_U3505) );
  MUX2_X1 U11117 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9890), .S(n10247), .Z(
        P1_U3502) );
  MUX2_X1 U11118 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9891), .S(n10247), .Z(
        P1_U3499) );
  MUX2_X1 U11119 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9892), .S(n10247), .Z(
        P1_U3496) );
  MUX2_X1 U11120 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9893), .S(n10247), .Z(
        P1_U3493) );
  NAND3_X1 U11121 ( .A1(n9895), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9897) );
  OAI22_X1 U11122 ( .A1(n9894), .A2(n9897), .B1(n6768), .B2(n9896), .ZN(n9898)
         );
  INV_X1 U11123 ( .A(n9898), .ZN(n9899) );
  OAI21_X1 U11124 ( .B1(n9900), .B2(n4480), .A(n9899), .ZN(P1_U3322) );
  OAI222_X1 U11125 ( .A1(n4480), .A2(n9904), .B1(n9903), .B2(P1_U3084), .C1(
        n9902), .C2(n9901), .ZN(P1_U3324) );
  AOI22_X1 U11126 ( .A1(n10260), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9916) );
  AOI211_X1 U11127 ( .C1(n9907), .C2(n9906), .A(n9905), .B(n10263), .ZN(n9908)
         );
  AOI21_X1 U11128 ( .B1(n9921), .B2(n9909), .A(n9908), .ZN(n9915) );
  INV_X1 U11129 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9910) );
  NOR2_X1 U11130 ( .A1(n9910), .A2(n5916), .ZN(n9913) );
  OAI211_X1 U11131 ( .C1(n9913), .C2(n9912), .A(n10258), .B(n9911), .ZN(n9914)
         );
  NAND3_X1 U11132 ( .A1(n9916), .A2(n9915), .A3(n9914), .ZN(P2_U3246) );
  AOI22_X1 U11133 ( .A1(n10260), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9927) );
  AOI211_X1 U11134 ( .C1(n9919), .C2(n9918), .A(n9917), .B(n10263), .ZN(n9920)
         );
  AOI21_X1 U11135 ( .B1(n9921), .B2(n4697), .A(n9920), .ZN(n9926) );
  OAI211_X1 U11136 ( .C1(n9924), .C2(n9923), .A(n10258), .B(n9922), .ZN(n9925)
         );
  NAND3_X1 U11137 ( .A1(n9927), .A2(n9926), .A3(n9925), .ZN(P2_U3247) );
  XNOR2_X1 U11138 ( .A(n9928), .B(n9934), .ZN(n9963) );
  INV_X1 U11139 ( .A(n9929), .ZN(n9930) );
  AOI21_X1 U11140 ( .B1(n9932), .B2(n9931), .A(n9930), .ZN(n9933) );
  XOR2_X1 U11141 ( .A(n9934), .B(n9933), .Z(n9941) );
  AOI22_X1 U11142 ( .A1(n9938), .A2(n9937), .B1(n9936), .B2(n9935), .ZN(n9939)
         );
  OAI21_X1 U11143 ( .B1(n9941), .B2(n9940), .A(n9939), .ZN(n9942) );
  AOI21_X1 U11144 ( .B1(n9963), .B2(n9943), .A(n9942), .ZN(n9960) );
  INV_X1 U11145 ( .A(n9944), .ZN(n9945) );
  AOI222_X1 U11146 ( .A1(n9948), .A2(n9947), .B1(P1_REG2_REG_10__SCAN_IN), 
        .B2(n10193), .C1(n9946), .C2(n9945), .ZN(n9957) );
  INV_X1 U11147 ( .A(n9949), .ZN(n9951) );
  OAI211_X1 U11148 ( .C1(n9959), .C2(n9952), .A(n9951), .B(n9950), .ZN(n9958)
         );
  INV_X1 U11149 ( .A(n9958), .ZN(n9953) );
  AOI22_X1 U11150 ( .A1(n9963), .A2(n9955), .B1(n9954), .B2(n9953), .ZN(n9956)
         );
  OAI211_X1 U11151 ( .C1(n10193), .C2(n9960), .A(n9957), .B(n9956), .ZN(
        P1_U3281) );
  OAI21_X1 U11152 ( .B1(n9959), .B2(n10237), .A(n9958), .ZN(n9962) );
  INV_X1 U11153 ( .A(n9960), .ZN(n9961) );
  AOI211_X1 U11154 ( .C1(n10244), .C2(n9963), .A(n9962), .B(n9961), .ZN(n9965)
         );
  INV_X1 U11155 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9964) );
  AOI22_X1 U11156 ( .A1(n10247), .A2(n9965), .B1(n9964), .B2(n10245), .ZN(
        P1_U3484) );
  AOI22_X1 U11157 ( .A1(n10255), .A2(n9965), .B1(n6876), .B2(n10256), .ZN(
        P1_U3533) );
  AOI21_X1 U11158 ( .B1(n4557), .B2(n4935), .A(n9966), .ZN(n9969) );
  AOI21_X1 U11159 ( .B1(n9969), .B2(n9968), .A(n9967), .ZN(n9984) );
  INV_X1 U11160 ( .A(n9970), .ZN(n9971) );
  AOI222_X1 U11161 ( .A1(n9972), .A2(n10284), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n10293), .C1(n10283), .C2(n9971), .ZN(n9982) );
  AOI21_X1 U11162 ( .B1(n9975), .B2(n9974), .A(n9973), .ZN(n9976) );
  INV_X1 U11163 ( .A(n9976), .ZN(n9987) );
  INV_X1 U11164 ( .A(n9977), .ZN(n9979) );
  OAI211_X1 U11165 ( .C1(n9985), .C2(n4561), .A(n9979), .B(n9978), .ZN(n9983)
         );
  INV_X1 U11166 ( .A(n9983), .ZN(n9980) );
  AOI22_X1 U11167 ( .A1(n9987), .A2(n10288), .B1(n10287), .B2(n9980), .ZN(
        n9981) );
  OAI211_X1 U11168 ( .C1(n10293), .C2(n9984), .A(n9982), .B(n9981), .ZN(
        P2_U3282) );
  OAI211_X1 U11169 ( .C1(n9985), .C2(n10381), .A(n9984), .B(n9983), .ZN(n9986)
         );
  AOI21_X1 U11170 ( .B1(n9987), .B2(n10391), .A(n9986), .ZN(n9988) );
  AOI22_X1 U11171 ( .A1(n10406), .A2(n9988), .B1(n6111), .B2(n10404), .ZN(
        P2_U3534) );
  AOI22_X1 U11172 ( .A1(n10395), .A2(n9988), .B1(n6115), .B2(n10393), .ZN(
        P2_U3493) );
  INV_X1 U11173 ( .A(n9989), .ZN(n9992) );
  NOR2_X1 U11174 ( .A1(n9990), .A2(n10239), .ZN(n9991) );
  INV_X1 U11175 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9995) );
  AOI22_X1 U11176 ( .A1(n10255), .A2(n10011), .B1(n9995), .B2(n10256), .ZN(
        P1_U3553) );
  INV_X1 U11177 ( .A(n9996), .ZN(n9998) );
  OAI21_X1 U11178 ( .B1(n9998), .B2(n10237), .A(n9997), .ZN(n9999) );
  AOI21_X1 U11179 ( .B1(n10000), .B2(n10244), .A(n9999), .ZN(n10001) );
  AND2_X1 U11180 ( .A1(n10002), .A2(n10001), .ZN(n10013) );
  AOI22_X1 U11181 ( .A1(n10255), .A2(n10013), .B1(n7510), .B2(n10256), .ZN(
        P1_U3535) );
  OAI22_X1 U11182 ( .A1(n10004), .A2(n10239), .B1(n10003), .B2(n10237), .ZN(
        n10005) );
  AOI21_X1 U11183 ( .B1(n10006), .B2(n10244), .A(n10005), .ZN(n10007) );
  AND2_X1 U11184 ( .A1(n10008), .A2(n10007), .ZN(n10014) );
  AOI22_X1 U11185 ( .A1(n10255), .A2(n10014), .B1(n10009), .B2(n10256), .ZN(
        P1_U3534) );
  INV_X1 U11186 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10010) );
  AOI22_X1 U11187 ( .A1(n10247), .A2(n10011), .B1(n10010), .B2(n10245), .ZN(
        P1_U3521) );
  INV_X1 U11188 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10012) );
  AOI22_X1 U11189 ( .A1(n10247), .A2(n10013), .B1(n10012), .B2(n10245), .ZN(
        P1_U3490) );
  AOI22_X1 U11190 ( .A1(n10247), .A2(n10014), .B1(n5375), .B2(n10245), .ZN(
        P1_U3487) );
  XNOR2_X1 U11191 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11192 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U11193 ( .B1(n10017), .B2(n10016), .A(n10015), .ZN(n10022) );
  NAND2_X1 U11194 ( .A1(n10041), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n10021) );
  INV_X1 U11195 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10186) );
  NOR2_X1 U11196 ( .A1(n10186), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10018) );
  AOI21_X1 U11197 ( .B1(n10168), .B2(n10019), .A(n10018), .ZN(n10020) );
  OAI211_X1 U11198 ( .C1(n10161), .C2(n10022), .A(n10021), .B(n10020), .ZN(
        n10023) );
  INV_X1 U11199 ( .A(n10023), .ZN(n10028) );
  OAI211_X1 U11200 ( .C1(n10026), .C2(n10025), .A(n10170), .B(n10024), .ZN(
        n10027) );
  NAND2_X1 U11201 ( .A1(n10028), .A2(n10027), .ZN(P1_U3242) );
  OAI21_X1 U11202 ( .B1(n10031), .B2(n10030), .A(n10029), .ZN(n10034) );
  INV_X1 U11203 ( .A(n10032), .ZN(n10033) );
  AOI22_X1 U11204 ( .A1(n10088), .A2(n10034), .B1(n10033), .B2(n10168), .ZN(
        n10045) );
  OAI21_X1 U11205 ( .B1(n10037), .B2(n10036), .A(n10035), .ZN(n10038) );
  AND2_X1 U11206 ( .A1(n10170), .A2(n10038), .ZN(n10039) );
  AOI211_X1 U11207 ( .C1(P1_ADDR_REG_4__SCAN_IN), .C2(n10041), .A(n10040), .B(
        n10039), .ZN(n10044) );
  INV_X1 U11208 ( .A(n10042), .ZN(n10043) );
  NAND3_X1 U11209 ( .A1(n10045), .A2(n10044), .A3(n10043), .ZN(P1_U3245) );
  OAI21_X1 U11210 ( .B1(n10048), .B2(n10047), .A(n10046), .ZN(n10049) );
  INV_X1 U11211 ( .A(n10049), .ZN(n10054) );
  INV_X1 U11212 ( .A(n10050), .ZN(n10053) );
  NAND2_X1 U11213 ( .A1(n10168), .A2(n10051), .ZN(n10052) );
  OAI211_X1 U11214 ( .C1(n10161), .C2(n10054), .A(n10053), .B(n10052), .ZN(
        n10055) );
  INV_X1 U11215 ( .A(n10055), .ZN(n10062) );
  INV_X1 U11216 ( .A(n10056), .ZN(n10060) );
  INV_X1 U11217 ( .A(n10057), .ZN(n10059) );
  OAI211_X1 U11218 ( .C1(n10060), .C2(n10059), .A(n10170), .B(n10058), .ZN(
        n10061) );
  OAI211_X1 U11219 ( .C1(n10448), .C2(n10175), .A(n10062), .B(n10061), .ZN(
        P1_U3246) );
  INV_X1 U11220 ( .A(n10063), .ZN(n10065) );
  NAND2_X1 U11221 ( .A1(n10065), .A2(n10064), .ZN(n10066) );
  NAND2_X1 U11222 ( .A1(n10067), .A2(n10066), .ZN(n10072) );
  INV_X1 U11223 ( .A(n10068), .ZN(n10071) );
  NAND2_X1 U11224 ( .A1(n10168), .A2(n10069), .ZN(n10070) );
  OAI211_X1 U11225 ( .C1(n10161), .C2(n10072), .A(n10071), .B(n10070), .ZN(
        n10073) );
  INV_X1 U11226 ( .A(n10073), .ZN(n10079) );
  AOI21_X1 U11227 ( .B1(n10076), .B2(n10075), .A(n10074), .ZN(n10077) );
  OR2_X1 U11228 ( .A1(n10131), .A2(n10077), .ZN(n10078) );
  OAI211_X1 U11229 ( .C1(n10080), .C2(n10175), .A(n10079), .B(n10078), .ZN(
        P1_U3247) );
  OAI21_X1 U11230 ( .B1(n10083), .B2(n10082), .A(n10081), .ZN(n10089) );
  NOR2_X1 U11231 ( .A1(n10085), .A2(n10084), .ZN(n10086) );
  AOI211_X1 U11232 ( .C1(n10089), .C2(n10088), .A(n10087), .B(n10086), .ZN(
        n10095) );
  AOI21_X1 U11233 ( .B1(n10092), .B2(n10091), .A(n10090), .ZN(n10093) );
  OR2_X1 U11234 ( .A1(n10093), .A2(n10131), .ZN(n10094) );
  OAI211_X1 U11235 ( .C1(n10175), .C2(n10096), .A(n10095), .B(n10094), .ZN(
        P1_U3249) );
  AOI211_X1 U11236 ( .C1(n10099), .C2(n10098), .A(n10097), .B(n10161), .ZN(
        n10100) );
  AOI211_X1 U11237 ( .C1(n10168), .C2(n10102), .A(n10101), .B(n10100), .ZN(
        n10108) );
  AOI21_X1 U11238 ( .B1(n10105), .B2(n10104), .A(n10103), .ZN(n10106) );
  OR2_X1 U11239 ( .A1(n10106), .A2(n10131), .ZN(n10107) );
  OAI211_X1 U11240 ( .C1(n10455), .C2(n10175), .A(n10108), .B(n10107), .ZN(
        P1_U3250) );
  INV_X1 U11241 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10121) );
  AOI211_X1 U11242 ( .C1(n10111), .C2(n10110), .A(n10161), .B(n10109), .ZN(
        n10112) );
  AOI211_X1 U11243 ( .C1(n10168), .C2(n10114), .A(n10113), .B(n10112), .ZN(
        n10120) );
  AOI21_X1 U11244 ( .B1(n10117), .B2(n10116), .A(n10115), .ZN(n10118) );
  OR2_X1 U11245 ( .A1(n10118), .A2(n10131), .ZN(n10119) );
  OAI211_X1 U11246 ( .C1(n10121), .C2(n10175), .A(n10120), .B(n10119), .ZN(
        P1_U3253) );
  INV_X1 U11247 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10135) );
  AOI211_X1 U11248 ( .C1(n10124), .C2(n10123), .A(n10122), .B(n10161), .ZN(
        n10125) );
  AOI211_X1 U11249 ( .C1(n10168), .C2(n10127), .A(n10126), .B(n10125), .ZN(
        n10134) );
  AOI21_X1 U11250 ( .B1(n10130), .B2(n10129), .A(n10128), .ZN(n10132) );
  OR2_X1 U11251 ( .A1(n10132), .A2(n10131), .ZN(n10133) );
  OAI211_X1 U11252 ( .C1(n10135), .C2(n10175), .A(n10134), .B(n10133), .ZN(
        P1_U3254) );
  INV_X1 U11253 ( .A(n10136), .ZN(n10140) );
  AOI211_X1 U11254 ( .C1(n10138), .C2(n9778), .A(n10137), .B(n10161), .ZN(
        n10139) );
  AOI211_X1 U11255 ( .C1(n10168), .C2(n10141), .A(n10140), .B(n10139), .ZN(
        n10145) );
  OAI211_X1 U11256 ( .C1(n10143), .C2(P1_REG1_REG_15__SCAN_IN), .A(n10170), 
        .B(n10142), .ZN(n10144) );
  OAI211_X1 U11257 ( .C1(n10175), .C2(n10146), .A(n10145), .B(n10144), .ZN(
        P1_U3256) );
  INV_X1 U11258 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10159) );
  INV_X1 U11259 ( .A(n10147), .ZN(n10152) );
  AOI211_X1 U11260 ( .C1(n10150), .C2(n10149), .A(n10148), .B(n10161), .ZN(
        n10151) );
  AOI211_X1 U11261 ( .C1(n10168), .C2(n10153), .A(n10152), .B(n10151), .ZN(
        n10158) );
  OAI211_X1 U11262 ( .C1(n10156), .C2(n10155), .A(n10170), .B(n10154), .ZN(
        n10157) );
  OAI211_X1 U11263 ( .C1(n10159), .C2(n10175), .A(n10158), .B(n10157), .ZN(
        P1_U3257) );
  INV_X1 U11264 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10176) );
  INV_X1 U11265 ( .A(n10160), .ZN(n10166) );
  AOI211_X1 U11266 ( .C1(n10164), .C2(n10163), .A(n10162), .B(n10161), .ZN(
        n10165) );
  AOI211_X1 U11267 ( .C1(n10168), .C2(n10167), .A(n10166), .B(n10165), .ZN(
        n10174) );
  OAI211_X1 U11268 ( .C1(n10172), .C2(n10171), .A(n10170), .B(n10169), .ZN(
        n10173) );
  OAI211_X1 U11269 ( .C1(n10176), .C2(n10175), .A(n10174), .B(n10173), .ZN(
        P1_U3258) );
  INV_X1 U11270 ( .A(n10177), .ZN(n10190) );
  NOR2_X1 U11271 ( .A1(n10179), .A2(n10178), .ZN(n10181) );
  MUX2_X1 U11272 ( .A(n10182), .B(n10181), .S(n10180), .Z(n10189) );
  INV_X1 U11273 ( .A(n10183), .ZN(n10184) );
  OAI22_X1 U11274 ( .A1(n10187), .A2(n10186), .B1(n10185), .B2(n10184), .ZN(
        n10188) );
  NOR3_X1 U11275 ( .A1(n10190), .A2(n10189), .A3(n10188), .ZN(n10191) );
  AOI22_X1 U11276 ( .A1(n10193), .A2(n10192), .B1(n10191), .B2(n9774), .ZN(
        P1_U3290) );
  NOR2_X1 U11277 ( .A1(n10203), .A2(n10194), .ZN(P1_U3292) );
  NOR2_X1 U11278 ( .A1(n10203), .A2(n10195), .ZN(P1_U3293) );
  AND2_X1 U11279 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10201), .ZN(P1_U3294) );
  NOR2_X1 U11280 ( .A1(n10203), .A2(n10196), .ZN(P1_U3295) );
  AND2_X1 U11281 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10201), .ZN(P1_U3296) );
  AND2_X1 U11282 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10201), .ZN(P1_U3297) );
  AND2_X1 U11283 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10201), .ZN(P1_U3298) );
  NOR2_X1 U11284 ( .A1(n10203), .A2(n10197), .ZN(P1_U3299) );
  NOR2_X1 U11285 ( .A1(n10203), .A2(n10198), .ZN(P1_U3300) );
  AND2_X1 U11286 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10201), .ZN(P1_U3301) );
  AND2_X1 U11287 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10201), .ZN(P1_U3302) );
  AND2_X1 U11288 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10201), .ZN(P1_U3303) );
  AND2_X1 U11289 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10201), .ZN(P1_U3304) );
  AND2_X1 U11290 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10201), .ZN(P1_U3305) );
  NOR2_X1 U11291 ( .A1(n10203), .A2(n10199), .ZN(P1_U3306) );
  AND2_X1 U11292 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10201), .ZN(P1_U3307) );
  AND2_X1 U11293 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10201), .ZN(P1_U3308) );
  AND2_X1 U11294 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10201), .ZN(P1_U3309) );
  AND2_X1 U11295 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10201), .ZN(P1_U3310) );
  AND2_X1 U11296 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10201), .ZN(P1_U3311) );
  AND2_X1 U11297 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10201), .ZN(P1_U3312) );
  NOR2_X1 U11298 ( .A1(n10203), .A2(n10200), .ZN(P1_U3313) );
  AND2_X1 U11299 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10201), .ZN(P1_U3314) );
  AND2_X1 U11300 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10201), .ZN(P1_U3315) );
  AND2_X1 U11301 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10201), .ZN(P1_U3316) );
  AND2_X1 U11302 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10201), .ZN(P1_U3317) );
  AND2_X1 U11303 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10201), .ZN(P1_U3318) );
  AND2_X1 U11304 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10201), .ZN(P1_U3319) );
  AND2_X1 U11305 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10201), .ZN(P1_U3320) );
  NOR2_X1 U11306 ( .A1(n10203), .A2(n10202), .ZN(P1_U3321) );
  INV_X1 U11307 ( .A(n10204), .ZN(n10209) );
  OAI22_X1 U11308 ( .A1(n10206), .A2(n10239), .B1(n10205), .B2(n10237), .ZN(
        n10208) );
  AOI211_X1 U11309 ( .C1(n10244), .C2(n10209), .A(n10208), .B(n10207), .ZN(
        n10249) );
  AOI22_X1 U11310 ( .A1(n10247), .A2(n10249), .B1(n5127), .B2(n10245), .ZN(
        P1_U3460) );
  OAI22_X1 U11311 ( .A1(n10211), .A2(n10239), .B1(n10210), .B2(n10237), .ZN(
        n10213) );
  AOI211_X1 U11312 ( .C1(n10244), .C2(n10214), .A(n10213), .B(n10212), .ZN(
        n10251) );
  AOI22_X1 U11313 ( .A1(n10247), .A2(n10251), .B1(n5176), .B2(n10245), .ZN(
        P1_U3466) );
  OAI211_X1 U11314 ( .C1(n10217), .C2(n10237), .A(n10216), .B(n10215), .ZN(
        n10220) );
  INV_X1 U11315 ( .A(n10218), .ZN(n10219) );
  AOI211_X1 U11316 ( .C1(n4981), .C2(n10221), .A(n10220), .B(n10219), .ZN(
        n10252) );
  AOI22_X1 U11317 ( .A1(n10247), .A2(n10252), .B1(n5205), .B2(n10245), .ZN(
        P1_U3469) );
  OAI22_X1 U11318 ( .A1(n10223), .A2(n10239), .B1(n10222), .B2(n10237), .ZN(
        n10225) );
  AOI211_X1 U11319 ( .C1(n10244), .C2(n10226), .A(n10225), .B(n10224), .ZN(
        n10253) );
  INV_X1 U11320 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10227) );
  AOI22_X1 U11321 ( .A1(n10247), .A2(n10253), .B1(n10227), .B2(n10245), .ZN(
        P1_U3472) );
  INV_X1 U11322 ( .A(n10228), .ZN(n10233) );
  OAI22_X1 U11323 ( .A1(n10230), .A2(n10239), .B1(n10229), .B2(n10237), .ZN(
        n10232) );
  AOI211_X1 U11324 ( .C1(n10244), .C2(n10233), .A(n10232), .B(n10231), .ZN(
        n10254) );
  INV_X1 U11325 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10234) );
  AOI22_X1 U11326 ( .A1(n10247), .A2(n10254), .B1(n10234), .B2(n10245), .ZN(
        P1_U3478) );
  INV_X1 U11327 ( .A(n10235), .ZN(n10243) );
  INV_X1 U11328 ( .A(n10236), .ZN(n10238) );
  OAI22_X1 U11329 ( .A1(n10240), .A2(n10239), .B1(n10238), .B2(n10237), .ZN(
        n10242) );
  AOI211_X1 U11330 ( .C1(n10244), .C2(n10243), .A(n10242), .B(n10241), .ZN(
        n10257) );
  INV_X1 U11331 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U11332 ( .A1(n10247), .A2(n10257), .B1(n10246), .B2(n10245), .ZN(
        P1_U3481) );
  AOI22_X1 U11333 ( .A1(n10255), .A2(n10249), .B1(n10248), .B2(n10256), .ZN(
        P1_U3525) );
  AOI22_X1 U11334 ( .A1(n10255), .A2(n10251), .B1(n10250), .B2(n10256), .ZN(
        P1_U3527) );
  AOI22_X1 U11335 ( .A1(n10255), .A2(n10252), .B1(n5204), .B2(n10256), .ZN(
        P1_U3528) );
  AOI22_X1 U11336 ( .A1(n10255), .A2(n10253), .B1(n6801), .B2(n10256), .ZN(
        P1_U3529) );
  AOI22_X1 U11337 ( .A1(n10255), .A2(n10254), .B1(n6873), .B2(n10256), .ZN(
        P1_U3531) );
  AOI22_X1 U11338 ( .A1(n10255), .A2(n10257), .B1(n6874), .B2(n10256), .ZN(
        P1_U3532) );
  AOI22_X1 U11339 ( .A1(n10259), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10258), .ZN(n10268) );
  AOI22_X1 U11340 ( .A1(n10260), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10267) );
  OAI21_X1 U11341 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n10262), .A(n10261), .ZN(
        n10265) );
  NOR2_X1 U11342 ( .A1(n10263), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10264) );
  OAI21_X1 U11343 ( .B1(n10265), .B2(n10264), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n10266) );
  OAI211_X1 U11344 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n10268), .A(n10267), .B(
        n10266), .ZN(P2_U3245) );
  INV_X1 U11345 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10281) );
  INV_X1 U11346 ( .A(n10269), .ZN(n10278) );
  INV_X1 U11347 ( .A(n10270), .ZN(n10275) );
  AOI22_X1 U11348 ( .A1(n10283), .A2(n10273), .B1(n10272), .B2(n10271), .ZN(
        n10274) );
  OAI21_X1 U11349 ( .B1(n10275), .B2(n4831), .A(n10274), .ZN(n10277) );
  AOI211_X1 U11350 ( .C1(n10279), .C2(n10278), .A(n10277), .B(n10276), .ZN(
        n10280) );
  AOI22_X1 U11351 ( .A1(n10293), .A2(n10281), .B1(n10280), .B2(n8915), .ZN(
        P2_U3291) );
  AOI22_X1 U11352 ( .A1(n10283), .A2(n10282), .B1(P2_REG2_REG_3__SCAN_IN), 
        .B2(n10293), .ZN(n10291) );
  AOI222_X1 U11353 ( .A1(n10289), .A2(n10288), .B1(n10287), .B2(n10286), .C1(
        n10285), .C2(n10284), .ZN(n10290) );
  OAI211_X1 U11354 ( .C1(n10293), .C2(n10292), .A(n10291), .B(n10290), .ZN(
        P2_U3293) );
  NOR2_X1 U11355 ( .A1(n10295), .A2(n10294), .ZN(n10308) );
  INV_X1 U11356 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n10296) );
  NOR2_X1 U11357 ( .A1(n10331), .A2(n10296), .ZN(P2_U3297) );
  INV_X1 U11358 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n10297) );
  NOR2_X1 U11359 ( .A1(n10331), .A2(n10297), .ZN(P2_U3298) );
  INV_X1 U11360 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10298) );
  NOR2_X1 U11361 ( .A1(n10308), .A2(n10298), .ZN(P2_U3299) );
  NOR2_X1 U11362 ( .A1(n10308), .A2(n10299), .ZN(P2_U3300) );
  INV_X1 U11363 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10300) );
  NOR2_X1 U11364 ( .A1(n10308), .A2(n10300), .ZN(P2_U3301) );
  INV_X1 U11365 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10301) );
  NOR2_X1 U11366 ( .A1(n10308), .A2(n10301), .ZN(P2_U3302) );
  NOR2_X1 U11367 ( .A1(n10308), .A2(n10302), .ZN(P2_U3303) );
  INV_X1 U11368 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10303) );
  NOR2_X1 U11369 ( .A1(n10308), .A2(n10303), .ZN(P2_U3304) );
  INV_X1 U11370 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10304) );
  NOR2_X1 U11371 ( .A1(n10308), .A2(n10304), .ZN(P2_U3305) );
  INV_X1 U11372 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10305) );
  NOR2_X1 U11373 ( .A1(n10308), .A2(n10305), .ZN(P2_U3306) );
  INV_X1 U11374 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10306) );
  NOR2_X1 U11375 ( .A1(n10308), .A2(n10306), .ZN(P2_U3307) );
  INV_X1 U11376 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10307) );
  NOR2_X1 U11377 ( .A1(n10308), .A2(n10307), .ZN(P2_U3308) );
  INV_X1 U11378 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n10309) );
  NOR2_X1 U11379 ( .A1(n10331), .A2(n10309), .ZN(P2_U3309) );
  INV_X1 U11380 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n10310) );
  NOR2_X1 U11381 ( .A1(n10331), .A2(n10310), .ZN(P2_U3310) );
  INV_X1 U11382 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10311) );
  NOR2_X1 U11383 ( .A1(n10331), .A2(n10311), .ZN(P2_U3311) );
  INV_X1 U11384 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10312) );
  NOR2_X1 U11385 ( .A1(n10331), .A2(n10312), .ZN(P2_U3312) );
  NOR2_X1 U11386 ( .A1(n10331), .A2(n10313), .ZN(P2_U3313) );
  INV_X1 U11387 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10314) );
  NOR2_X1 U11388 ( .A1(n10331), .A2(n10314), .ZN(P2_U3314) );
  INV_X1 U11389 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10315) );
  NOR2_X1 U11390 ( .A1(n10331), .A2(n10315), .ZN(P2_U3315) );
  INV_X1 U11391 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10316) );
  NOR2_X1 U11392 ( .A1(n10331), .A2(n10316), .ZN(P2_U3316) );
  INV_X1 U11393 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10317) );
  NOR2_X1 U11394 ( .A1(n10331), .A2(n10317), .ZN(P2_U3317) );
  INV_X1 U11395 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10318) );
  NOR2_X1 U11396 ( .A1(n10331), .A2(n10318), .ZN(P2_U3318) );
  INV_X1 U11397 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10319) );
  NOR2_X1 U11398 ( .A1(n10331), .A2(n10319), .ZN(P2_U3319) );
  INV_X1 U11399 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n10320) );
  NOR2_X1 U11400 ( .A1(n10331), .A2(n10320), .ZN(P2_U3320) );
  NOR2_X1 U11401 ( .A1(n10331), .A2(n10321), .ZN(P2_U3321) );
  INV_X1 U11402 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10322) );
  NOR2_X1 U11403 ( .A1(n10331), .A2(n10322), .ZN(P2_U3322) );
  INV_X1 U11404 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10323) );
  NOR2_X1 U11405 ( .A1(n10331), .A2(n10323), .ZN(P2_U3323) );
  INV_X1 U11406 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n10324) );
  NOR2_X1 U11407 ( .A1(n10331), .A2(n10324), .ZN(P2_U3324) );
  NOR2_X1 U11408 ( .A1(n10331), .A2(n10325), .ZN(P2_U3325) );
  INV_X1 U11409 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10326) );
  NOR2_X1 U11410 ( .A1(n10331), .A2(n10326), .ZN(P2_U3326) );
  OAI22_X1 U11411 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n10331), .B1(n10327), .B2(
        n10329), .ZN(n10328) );
  INV_X1 U11412 ( .A(n10328), .ZN(P2_U3437) );
  OAI22_X1 U11413 ( .A1(P2_D_REG_1__SCAN_IN), .A2(n10331), .B1(n10330), .B2(
        n10329), .ZN(n10332) );
  INV_X1 U11414 ( .A(n10332), .ZN(P2_U3438) );
  NOR2_X1 U11415 ( .A1(n10334), .A2(n10333), .ZN(n10336) );
  AOI211_X1 U11416 ( .C1(n10337), .C2(n10391), .A(n10336), .B(n10335), .ZN(
        n10396) );
  AOI22_X1 U11417 ( .A1(n10395), .A2(n10396), .B1(n5920), .B2(n10393), .ZN(
        P2_U3451) );
  OAI22_X1 U11418 ( .A1(n10339), .A2(n4832), .B1(n10338), .B2(n10381), .ZN(
        n10341) );
  AOI211_X1 U11419 ( .C1(n10391), .C2(n10342), .A(n10341), .B(n10340), .ZN(
        n10397) );
  AOI22_X1 U11420 ( .A1(n10395), .A2(n10397), .B1(n5930), .B2(n10393), .ZN(
        P2_U3454) );
  NAND3_X1 U11421 ( .A1(n10344), .A2(n10343), .A3(n10391), .ZN(n10348) );
  AOI21_X1 U11422 ( .B1(n10385), .B2(n10346), .A(n10345), .ZN(n10347) );
  AND3_X1 U11423 ( .A1(n10349), .A2(n10348), .A3(n10347), .ZN(n10398) );
  INV_X1 U11424 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U11425 ( .A1(n10395), .A2(n10398), .B1(n10350), .B2(n10393), .ZN(
        P2_U3469) );
  OAI22_X1 U11426 ( .A1(n10352), .A2(n4832), .B1(n10351), .B2(n10381), .ZN(
        n10354) );
  AOI211_X1 U11427 ( .C1(n10391), .C2(n10355), .A(n10354), .B(n10353), .ZN(
        n10399) );
  INV_X1 U11428 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10356) );
  AOI22_X1 U11429 ( .A1(n10395), .A2(n10399), .B1(n10356), .B2(n10393), .ZN(
        P2_U3472) );
  INV_X1 U11430 ( .A(n10357), .ZN(n10377) );
  INV_X1 U11431 ( .A(n10358), .ZN(n10363) );
  OAI22_X1 U11432 ( .A1(n10360), .A2(n4832), .B1(n10359), .B2(n10381), .ZN(
        n10362) );
  AOI211_X1 U11433 ( .C1(n10377), .C2(n10363), .A(n10362), .B(n10361), .ZN(
        n10400) );
  INV_X1 U11434 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U11435 ( .A1(n10395), .A2(n10400), .B1(n10364), .B2(n10393), .ZN(
        P2_U3475) );
  INV_X1 U11436 ( .A(n10365), .ZN(n10370) );
  OAI22_X1 U11437 ( .A1(n10367), .A2(n4832), .B1(n10366), .B2(n10381), .ZN(
        n10369) );
  AOI211_X1 U11438 ( .C1(n10377), .C2(n10370), .A(n10369), .B(n10368), .ZN(
        n10401) );
  AOI22_X1 U11439 ( .A1(n10395), .A2(n10401), .B1(n6038), .B2(n10393), .ZN(
        P2_U3478) );
  INV_X1 U11440 ( .A(n10371), .ZN(n10376) );
  OAI22_X1 U11441 ( .A1(n10373), .A2(n4832), .B1(n10372), .B2(n10381), .ZN(
        n10375) );
  AOI211_X1 U11442 ( .C1(n10377), .C2(n10376), .A(n10375), .B(n10374), .ZN(
        n10402) );
  AOI22_X1 U11443 ( .A1(n10395), .A2(n10402), .B1(n10378), .B2(n10393), .ZN(
        P2_U3481) );
  OAI211_X1 U11444 ( .C1(n10382), .C2(n10381), .A(n10380), .B(n10379), .ZN(
        n10383) );
  AOI21_X1 U11445 ( .B1(n10384), .B2(n10391), .A(n10383), .ZN(n10403) );
  AOI22_X1 U11446 ( .A1(n10395), .A2(n10403), .B1(n6068), .B2(n10393), .ZN(
        P2_U3484) );
  NAND2_X1 U11447 ( .A1(n10386), .A2(n10385), .ZN(n10387) );
  OAI211_X1 U11448 ( .C1(n4832), .C2(n10389), .A(n10388), .B(n10387), .ZN(
        n10390) );
  AOI21_X1 U11449 ( .B1(n10392), .B2(n10391), .A(n10390), .ZN(n10405) );
  AOI22_X1 U11450 ( .A1(n10395), .A2(n10405), .B1(n10394), .B2(n10393), .ZN(
        P2_U3487) );
  AOI22_X1 U11451 ( .A1(n10406), .A2(n10396), .B1(n5916), .B2(n10404), .ZN(
        P2_U3520) );
  AOI22_X1 U11452 ( .A1(n10406), .A2(n10397), .B1(n6837), .B2(n10404), .ZN(
        P2_U3521) );
  AOI22_X1 U11453 ( .A1(n10406), .A2(n10398), .B1(n6903), .B2(n10404), .ZN(
        P2_U3526) );
  AOI22_X1 U11454 ( .A1(n10406), .A2(n10399), .B1(n6918), .B2(n10404), .ZN(
        P2_U3527) );
  AOI22_X1 U11455 ( .A1(n10406), .A2(n10400), .B1(n6975), .B2(n10404), .ZN(
        P2_U3528) );
  AOI22_X1 U11456 ( .A1(n10406), .A2(n10401), .B1(n7070), .B2(n10404), .ZN(
        P2_U3529) );
  AOI22_X1 U11457 ( .A1(n10406), .A2(n10402), .B1(n6058), .B2(n10404), .ZN(
        P2_U3530) );
  AOI22_X1 U11458 ( .A1(n10406), .A2(n10403), .B1(n6073), .B2(n10404), .ZN(
        P2_U3531) );
  AOI22_X1 U11459 ( .A1(n10406), .A2(n10405), .B1(n7544), .B2(n10404), .ZN(
        P2_U3532) );
  OAI21_X1 U11460 ( .B1(n10409), .B2(n10408), .A(n10407), .ZN(n10410) );
  XNOR2_X1 U11461 ( .A(n10410), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(ADD_1071_U5)
         );
  INV_X1 U11462 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10412) );
  AOI21_X1 U11463 ( .B1(n10413), .B2(n10412), .A(n10411), .ZN(ADD_1071_U46) );
  OAI21_X1 U11464 ( .B1(n10416), .B2(n10415), .A(n10414), .ZN(ADD_1071_U56) );
  OAI21_X1 U11465 ( .B1(n10419), .B2(n10418), .A(n10417), .ZN(ADD_1071_U57) );
  OAI21_X1 U11466 ( .B1(n10422), .B2(n10421), .A(n10420), .ZN(ADD_1071_U58) );
  OAI21_X1 U11467 ( .B1(n10425), .B2(n10424), .A(n10423), .ZN(ADD_1071_U59) );
  OAI21_X1 U11468 ( .B1(n10428), .B2(n10427), .A(n10426), .ZN(ADD_1071_U60) );
  OAI21_X1 U11469 ( .B1(n10431), .B2(n10430), .A(n10429), .ZN(ADD_1071_U61) );
  AOI21_X1 U11470 ( .B1(n10434), .B2(n10433), .A(n10432), .ZN(ADD_1071_U62) );
  AOI21_X1 U11471 ( .B1(n10437), .B2(n10436), .A(n10435), .ZN(ADD_1071_U63) );
  AOI21_X1 U11472 ( .B1(n10440), .B2(n10439), .A(n10438), .ZN(ADD_1071_U50) );
  AOI21_X1 U11473 ( .B1(n10443), .B2(n10442), .A(n10441), .ZN(ADD_1071_U54) );
  OAI222_X1 U11474 ( .A1(n10448), .A2(n10447), .B1(n10448), .B2(n10446), .C1(
        n10445), .C2(n10444), .ZN(ADD_1071_U51) );
  OAI21_X1 U11475 ( .B1(n10451), .B2(n10450), .A(n10449), .ZN(n10452) );
  XNOR2_X1 U11476 ( .A(n10452), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11477 ( .B1(n10455), .B2(n10454), .A(n10453), .ZN(ADD_1071_U47) );
  AOI21_X1 U11478 ( .B1(n10458), .B2(n10457), .A(n10456), .ZN(ADD_1071_U49) );
  AOI21_X1 U11479 ( .B1(n10461), .B2(n10460), .A(n10459), .ZN(ADD_1071_U48) );
  AOI21_X1 U11480 ( .B1(n10464), .B2(n10463), .A(n10462), .ZN(ADD_1071_U53) );
  OAI21_X1 U11481 ( .B1(n10467), .B2(n10466), .A(n10465), .ZN(ADD_1071_U52) );
  NAND2_X1 U6139 ( .A1(n5089), .A2(n4523), .ZN(n7152) );
  AND4_X1 U6141 ( .A1(n9454), .A2(n9453), .A3(n9452), .A4(n9451), .ZN(n9455)
         );
  CLKBUF_X1 U4996 ( .A(n5738), .Z(n4593) );
  CLKBUF_X1 U5047 ( .A(n5953), .Z(n6312) );
  CLKBUF_X1 U5151 ( .A(n5578), .Z(n9671) );
  CLKBUF_X1 U5173 ( .A(n9159), .Z(n10469) );
  NOR2_X1 U6110 ( .A1(n5862), .A2(n7159), .ZN(n9159) );
endmodule

