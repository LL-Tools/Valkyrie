

module b15_C_AntiSAT_k_256_7 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
         keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
         keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
         keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
         keyinput144, keyinput145, keyinput146, keyinput147, keyinput148,
         keyinput149, keyinput150, keyinput151, keyinput152, keyinput153,
         keyinput154, keyinput155, keyinput156, keyinput157, keyinput158,
         keyinput159, keyinput160, keyinput161, keyinput162, keyinput163,
         keyinput164, keyinput165, keyinput166, keyinput167, keyinput168,
         keyinput169, keyinput170, keyinput171, keyinput172, keyinput173,
         keyinput174, keyinput175, keyinput176, keyinput177, keyinput178,
         keyinput179, keyinput180, keyinput181, keyinput182, keyinput183,
         keyinput184, keyinput185, keyinput186, keyinput187, keyinput188,
         keyinput189, keyinput190, keyinput191, keyinput192, keyinput193,
         keyinput194, keyinput195, keyinput196, keyinput197, keyinput198,
         keyinput199, keyinput200, keyinput201, keyinput202, keyinput203,
         keyinput204, keyinput205, keyinput206, keyinput207, keyinput208,
         keyinput209, keyinput210, keyinput211, keyinput212, keyinput213,
         keyinput214, keyinput215, keyinput216, keyinput217, keyinput218,
         keyinput219, keyinput220, keyinput221, keyinput222, keyinput223,
         keyinput224, keyinput225, keyinput226, keyinput227, keyinput228,
         keyinput229, keyinput230, keyinput231, keyinput232, keyinput233,
         keyinput234, keyinput235, keyinput236, keyinput237, keyinput238,
         keyinput239, keyinput240, keyinput241, keyinput242, keyinput243,
         keyinput244, keyinput245, keyinput246, keyinput247, keyinput248,
         keyinput249, keyinput250, keyinput251, keyinput252, keyinput253,
         keyinput254, keyinput255;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018;

  OR2_X1 U3635 ( .A1(n4996), .A2(n6457), .ZN(n3195) );
  CLKBUF_X2 U3636 ( .A(n3426), .Z(n3187) );
  CLKBUF_X2 U3637 ( .A(n3428), .Z(n3404) );
  INV_X1 U3638 ( .A(n3720), .ZN(n5955) );
  INV_X1 U3639 ( .A(n4307), .ZN(n5941) );
  INV_X1 U3640 ( .A(n4449), .ZN(n5987) );
  AND4_X1 U3641 ( .A1(n3288), .A2(n3287), .A3(n3286), .A4(n3285), .ZN(n3299)
         );
  AND4_X1 U3642 ( .A1(n3292), .A2(n3291), .A3(n3290), .A4(n3289), .ZN(n3298)
         );
  AND4_X1 U3643 ( .A1(n3316), .A2(n3315), .A3(n3314), .A4(n3313), .ZN(n3317)
         );
  INV_X1 U3644 ( .A(n3837), .ZN(n5960) );
  INV_X1 U3645 ( .A(n3347), .ZN(n5982) );
  NAND2_X1 U3646 ( .A1(n3197), .A2(n3199), .ZN(n3347) );
  AND2_X1 U3647 ( .A1(n3210), .A2(n4477), .ZN(n3426) );
  AND2_X1 U3648 ( .A1(n5012), .A2(n3211), .ZN(n3280) );
  AND2_X1 U3649 ( .A1(n5012), .A2(n4477), .ZN(n3425) );
  AND2_X1 U3650 ( .A1(n4474), .A2(n4578), .ZN(n3406) );
  AND2_X1 U3651 ( .A1(n4729), .A2(n4458), .ZN(n3427) );
  AND2_X1 U3652 ( .A1(n3211), .A2(n4458), .ZN(n3269) );
  NOR2_X2 U3653 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4458) );
  INV_X1 U3654 ( .A(n6457), .ZN(n5851) );
  AOI22_X1 U3655 ( .A1(n6902), .A2(keyinput251), .B1(n6845), .B2(keyinput164), 
        .ZN(n6844) );
  OR2_X1 U3656 ( .A1(n3453), .A2(n3452), .ZN(n3441) );
  OAI221_X1 U3657 ( .B1(n6902), .B2(keyinput251), .C1(n6845), .C2(keyinput164), 
        .A(n6844), .ZN(n6849) );
  AND2_X1 U3658 ( .A1(n3442), .A2(n3441), .ZN(n3443) );
  NAND4_X1 U3659 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3189)
         );
  NAND2_X1 U3660 ( .A1(n5941), .A2(n4297), .ZN(n5111) );
  NAND2_X1 U3661 ( .A1(n4500), .A2(n3925), .ZN(n4521) );
  BUF_X1 U3662 ( .A(n3720), .Z(n4297) );
  INV_X1 U3663 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6799) );
  INV_X1 U3664 ( .A(n5479), .ZN(n5679) );
  AND2_X1 U3665 ( .A1(n5591), .A2(n4237), .ZN(n5654) );
  INV_X1 U3666 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3885) );
  CLKBUF_X3 U3667 ( .A(n3732), .Z(n3191) );
  INV_X4 U3668 ( .A(n4925), .ZN(n3824) );
  NAND2_X2 U3669 ( .A1(n5286), .A2(n5287), .ZN(n5285) );
  INV_X4 U3670 ( .A(n3620), .ZN(n5304) );
  NAND2_X1 U3671 ( .A1(n3444), .A2(n3443), .ZN(n3514) );
  NOR2_X4 U3672 ( .A1(n3344), .A2(n3846), .ZN(n4286) );
  XNOR2_X2 U3673 ( .A(n3453), .B(n3452), .ZN(n3456) );
  OAI21_X2 U3674 ( .B1(n4488), .B2(n3470), .A(n3451), .ZN(n5847) );
  XNOR2_X1 U3675 ( .A(n4748), .B(n4747), .ZN(n5382) );
  NOR2_X2 U3676 ( .A1(n5191), .A2(n5178), .ZN(n5179) );
  NAND2_X1 U3677 ( .A1(n5076), .A2(n5077), .ZN(n5271) );
  INV_X2 U3678 ( .A(n3620), .ZN(n5806) );
  INV_X2 U3679 ( .A(n5654), .ZN(n5717) );
  AND2_X1 U3680 ( .A1(n3895), .A2(n4797), .ZN(n4435) );
  CLKBUF_X1 U3681 ( .A(n3898), .Z(n6217) );
  XNOR2_X1 U3682 ( .A(n3514), .B(n6087), .ZN(n3898) );
  NAND2_X2 U3683 ( .A1(n5204), .A2(n4447), .ZN(n5489) );
  NAND2_X2 U3684 ( .A1(n5733), .A2(n4449), .ZN(n5203) );
  CLKBUF_X1 U3685 ( .A(n4454), .Z(n6270) );
  AND2_X2 U3686 ( .A1(n5814), .A2(n4397), .ZN(n5829) );
  NAND2_X1 U3687 ( .A1(n5637), .A2(n5636), .ZN(n4635) );
  OR2_X1 U3688 ( .A1(n3365), .A2(n3364), .ZN(n3366) );
  CLKBUF_X1 U3689 ( .A(n3884), .Z(n6244) );
  AND2_X1 U3690 ( .A1(n3416), .A2(n3414), .ZN(n3385) );
  CLKBUF_X1 U3691 ( .A(n3354), .Z(n3485) );
  AND2_X1 U3692 ( .A1(n3328), .A2(n4327), .ZN(n3343) );
  OR2_X1 U3693 ( .A1(n4329), .A2(n5941), .ZN(n4277) );
  AND2_X1 U3694 ( .A1(n4441), .A2(n5976), .ZN(n4326) );
  BUF_X4 U3695 ( .A(n5170), .Z(n3188) );
  CLKBUF_X1 U3696 ( .A(n3346), .Z(n5976) );
  AND4_X1 U3697 ( .A1(n3236), .A2(n3235), .A3(n3234), .A4(n3233), .ZN(n3346)
         );
  NAND2_X1 U3698 ( .A1(n3201), .A2(n3198), .ZN(n3837) );
  INV_X2 U3699 ( .A(n3832), .ZN(n5971) );
  OR2_X2 U3700 ( .A1(n3275), .A2(n3274), .ZN(n4449) );
  NAND2_X1 U3701 ( .A1(n3200), .A2(n3203), .ZN(n3832) );
  AND4_X1 U3702 ( .A1(n3308), .A2(n3307), .A3(n3306), .A4(n3305), .ZN(n3319)
         );
  AND4_X1 U3703 ( .A1(n3312), .A2(n3311), .A3(n3310), .A4(n3309), .ZN(n3318)
         );
  AND4_X1 U3704 ( .A1(n3232), .A2(n3231), .A3(n3230), .A4(n3229), .ZN(n3233)
         );
  AND4_X1 U3705 ( .A1(n3304), .A2(n3303), .A3(n3302), .A4(n3301), .ZN(n3320)
         );
  AND4_X1 U3706 ( .A1(n3284), .A2(n3283), .A3(n3282), .A4(n3281), .ZN(n3300)
         );
  BUF_X2 U3707 ( .A(n4765), .Z(n4893) );
  CLKBUF_X2 U3708 ( .A(n3280), .Z(n4894) );
  OR2_X2 U3709 ( .A1(n6523), .A2(n6454), .ZN(n6457) );
  BUF_X2 U3710 ( .A(n3427), .Z(n4895) );
  BUF_X2 U3711 ( .A(n3399), .Z(n4898) );
  BUF_X2 U3712 ( .A(n3425), .Z(n4869) );
  BUF_X2 U3713 ( .A(n3269), .Z(n4905) );
  INV_X2 U3714 ( .A(n6621), .ZN(n6609) );
  BUF_X2 U3715 ( .A(n3406), .Z(n4812) );
  AND2_X2 U3716 ( .A1(n3635), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4729)
         );
  INV_X1 U3717 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5015) );
  AND2_X2 U3718 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4474) );
  AND2_X2 U3719 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4578) );
  INV_X2 U3720 ( .A(n5181), .ZN(n5170) );
  NAND4_X4 U3721 ( .A1(n3300), .A2(n3299), .A3(n3298), .A4(n3297), .ZN(n3720)
         );
  NAND4_X1 U3722 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3190)
         );
  NAND4_X1 U3723 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n4307)
         );
  AOI211_X2 U3724 ( .C1(REIP_REG_31__SCAN_IN), .C2(n4980), .A(n4979), .B(n4978), .ZN(n4981) );
  NAND2_X1 U3725 ( .A1(n5966), .A2(n3190), .ZN(n3732) );
  NOR2_X1 U3726 ( .A1(n3535), .A2(n3534), .ZN(n3549) );
  NAND2_X1 U3727 ( .A1(n5971), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3492) );
  AND3_X1 U3728 ( .A1(n3832), .A2(STATE2_REG_0__SCAN_IN), .A3(n4307), .ZN(
        n3676) );
  OR2_X1 U3729 ( .A1(n4934), .A2(n3612), .ZN(n4734) );
  OR2_X1 U3730 ( .A1(n3571), .A2(n3570), .ZN(n3594) );
  AND4_X1 U3731 ( .A1(n3220), .A2(n3219), .A3(n3218), .A4(n3217), .ZN(n3236)
         );
  AND4_X1 U3732 ( .A1(n3228), .A2(n3227), .A3(n3226), .A4(n3225), .ZN(n3234)
         );
  AND4_X1 U3733 ( .A1(n3224), .A2(n3223), .A3(n3222), .A4(n3221), .ZN(n3235)
         );
  OR2_X1 U3734 ( .A1(n6610), .A2(n4222), .ZN(n5591) );
  OR2_X2 U3735 ( .A1(n5271), .A2(n5189), .ZN(n5191) );
  OR2_X1 U3736 ( .A1(n3378), .A2(n3377), .ZN(n3379) );
  NAND2_X1 U3737 ( .A1(n4438), .A2(n5971), .ZN(n3326) );
  NOR2_X1 U3738 ( .A1(n5028), .A2(n4889), .ZN(n4920) );
  AND2_X1 U3739 ( .A1(n4527), .A2(n4526), .ZN(n4525) );
  OR2_X1 U3740 ( .A1(n4449), .A2(n6799), .ZN(n4861) );
  OR2_X1 U3741 ( .A1(n4687), .A2(n4691), .ZN(n4249) );
  NAND2_X1 U3742 ( .A1(n3463), .A2(n3465), .ZN(n3464) );
  NAND2_X1 U3743 ( .A1(n4454), .A2(n6517), .ZN(n3505) );
  CLKBUF_X1 U3744 ( .A(n4920), .Z(n4890) );
  AND2_X1 U3745 ( .A1(n4806), .A2(n5077), .ZN(n5149) );
  AND2_X1 U3746 ( .A1(n4102), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4103)
         );
  AND2_X1 U3747 ( .A1(n4501), .A2(n4499), .ZN(n3925) );
  NAND2_X1 U3748 ( .A1(n3920), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3919)
         );
  OR2_X1 U3749 ( .A1(n5806), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3629)
         );
  INV_X1 U3750 ( .A(n5285), .ZN(n4744) );
  NAND2_X1 U3751 ( .A1(n4738), .A2(n4737), .ZN(n5293) );
  NAND2_X1 U3752 ( .A1(n3594), .A2(n3593), .ZN(n3606) );
  NAND2_X1 U3753 ( .A1(n3717), .A2(n6515), .ZN(n3859) );
  NAND2_X1 U3754 ( .A1(n3514), .A2(n3447), .ZN(n4488) );
  XNOR2_X1 U3755 ( .A(n4478), .B(n6340), .ZN(n4454) );
  NAND2_X1 U3756 ( .A1(n3689), .A2(n3688), .ZN(n4317) );
  INV_X1 U3757 ( .A(n6052), .ZN(n6051) );
  AND2_X1 U3758 ( .A1(n6458), .A2(n5945), .ZN(n6299) );
  INV_X1 U3759 ( .A(n4243), .ZN(n4244) );
  NOR2_X1 U3760 ( .A1(n5718), .A2(n6970), .ZN(n4245) );
  AND2_X1 U3761 ( .A1(n4972), .A2(n4236), .ZN(n5687) );
  INV_X1 U3762 ( .A(n5696), .ZN(n5718) );
  AND2_X1 U3763 ( .A1(n5204), .A2(n4448), .ZN(n5737) );
  AND2_X1 U3764 ( .A1(n5204), .A2(n4450), .ZN(n5741) );
  INV_X1 U3765 ( .A(n5204), .ZN(n5740) );
  NAND2_X1 U3766 ( .A1(n4758), .A2(n4215), .ZN(n4220) );
  OR2_X1 U3767 ( .A1(n5829), .A2(n4531), .ZN(n5856) );
  XNOR2_X1 U3768 ( .A(n3831), .B(n4927), .ZN(n5026) );
  AND2_X1 U3769 ( .A1(n3204), .A2(n3634), .ZN(n5007) );
  AND2_X1 U3770 ( .A1(n5380), .A2(n3873), .ZN(n5368) );
  NOR2_X1 U3771 ( .A1(n3705), .A2(n3325), .ZN(n3329) );
  OR2_X1 U3772 ( .A1(n3641), .A2(n3644), .ZN(n3643) );
  AND2_X1 U3773 ( .A1(n3669), .A2(n3668), .ZN(n3671) );
  CLKBUF_X1 U3774 ( .A(n3497), .Z(n4897) );
  OR2_X1 U3775 ( .A1(n3396), .A2(n3395), .ZN(n3448) );
  INV_X1 U3776 ( .A(n3448), .ZN(n3457) );
  NAND2_X1 U3777 ( .A1(n3492), .A2(n3491), .ZN(n3683) );
  BUF_X1 U3778 ( .A(n3324), .Z(n3645) );
  INV_X1 U3779 ( .A(n3346), .ZN(n3324) );
  OR2_X1 U3780 ( .A1(n4027), .A2(n4026), .ZN(n4040) );
  NAND2_X1 U3781 ( .A1(n3971), .A2(n3970), .ZN(n4552) );
  INV_X1 U3782 ( .A(n4861), .ZN(n4965) );
  NAND2_X1 U3783 ( .A1(n3571), .A2(n3550), .ZN(n3913) );
  AND2_X1 U3784 ( .A1(n4331), .A2(n3847), .ZN(n4323) );
  AND2_X1 U3785 ( .A1(n3645), .A2(n4297), .ZN(n3640) );
  OR2_X1 U3786 ( .A1(n3434), .A2(n3433), .ZN(n3471) );
  XNOR2_X1 U3787 ( .A(n3382), .B(n3381), .ZN(n3444) );
  AOI22_X1 U3788 ( .A1(n3380), .A2(n3379), .B1(n3676), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3381) );
  MUX2_X1 U3789 ( .A(n3326), .B(n3253), .S(n3347), .Z(n3279) );
  NAND2_X1 U3790 ( .A1(n3363), .A2(n3362), .ZN(n3364) );
  INV_X1 U3791 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6212) );
  AOI21_X1 U3792 ( .B1(n3439), .B2(n3465), .A(n3592), .ZN(n3454) );
  OAI21_X1 U3793 ( .B1(n6616), .B2(n4485), .A(n5009), .ZN(n5940) );
  INV_X1 U3794 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6213) );
  INV_X1 U3795 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5127) );
  AND2_X1 U3796 ( .A1(n3743), .A2(n3742), .ZN(n4427) );
  NAND2_X1 U3797 ( .A1(n3932), .A2(n4052), .ZN(n3939) );
  AND2_X1 U3798 ( .A1(n4847), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4865)
         );
  NAND2_X1 U3799 ( .A1(n4865), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4886)
         );
  AND2_X1 U3800 ( .A1(n5149), .A2(n4829), .ZN(n4830) );
  NOR2_X1 U3801 ( .A1(n4211), .A2(n6970), .ZN(n4796) );
  AND2_X1 U3802 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n4135), .ZN(n4137)
         );
  NAND2_X1 U3803 ( .A1(n4137), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4211)
         );
  NOR2_X1 U3804 ( .A1(n4134), .A2(n5296), .ZN(n4183) );
  NAND2_X1 U3805 ( .A1(n4183), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4184)
         );
  NAND2_X1 U3806 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n4103), .ZN(n4134)
         );
  NOR2_X1 U3807 ( .A1(n4088), .A2(n4087), .ZN(n4102) );
  NAND2_X1 U3808 ( .A1(n4072), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4088)
         );
  OR2_X2 U3809 ( .A1(n4677), .A2(n4944), .ZN(n5196) );
  BUF_X1 U3810 ( .A(n5076), .Z(n5195) );
  NAND2_X1 U3811 ( .A1(n4672), .A2(n4040), .ZN(n4679) );
  CLKBUF_X1 U3812 ( .A(n4677), .Z(n4943) );
  NAND2_X1 U3813 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n4023), .ZN(n4056)
         );
  NAND2_X1 U3814 ( .A1(n4668), .A2(n4669), .ZN(n4672) );
  NOR2_X1 U3815 ( .A1(n6845), .A2(n3974), .ZN(n4023) );
  NOR2_X1 U3816 ( .A1(n4006), .A2(n3973), .ZN(n3991) );
  NAND2_X1 U3817 ( .A1(n3972), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4006)
         );
  INV_X1 U3819 ( .A(n3933), .ZN(n3934) );
  NOR2_X1 U3820 ( .A1(n3919), .A2(n5685), .ZN(n3926) );
  NAND2_X1 U3821 ( .A1(n3924), .A2(n3923), .ZN(n4499) );
  NOR3_X1 U3822 ( .A1(n5138), .A2(n5127), .A3(n3900), .ZN(n3920) );
  INV_X1 U3823 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3900) );
  NAND2_X1 U3824 ( .A1(n5233), .A2(n3630), .ZN(n3632) );
  NAND2_X1 U3825 ( .A1(n3628), .A2(n3627), .ZN(n5251) );
  NOR2_X1 U3826 ( .A1(n3620), .A2(n6782), .ZN(n3627) );
  INV_X1 U3827 ( .A(n5259), .ZN(n3628) );
  AOI21_X1 U3828 ( .B1(n4251), .B2(n3202), .A(n3194), .ZN(n3622) );
  AOI21_X1 U3829 ( .B1(n5404), .B2(n4743), .A(n4742), .ZN(n5286) );
  AND2_X1 U3830 ( .A1(n5303), .A2(n5302), .ZN(n5307) );
  AND2_X1 U3831 ( .A1(n5304), .A2(n4711), .ZN(n4690) );
  OR2_X1 U3832 ( .A1(n5515), .A2(n3610), .ZN(n4687) );
  AND2_X1 U3833 ( .A1(n5517), .A2(n3614), .ZN(n4688) );
  CLKBUF_X1 U3834 ( .A(n4686), .Z(n5516) );
  AND2_X1 U3835 ( .A1(n3484), .A2(n3483), .ZN(n4535) );
  OR2_X1 U3836 ( .A1(n3859), .A2(n4583), .ZN(n4702) );
  NAND2_X1 U3837 ( .A1(n3464), .A2(n3467), .ZN(n3469) );
  AND2_X1 U3839 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4455) );
  NAND2_X1 U3840 ( .A1(n3490), .A2(n3489), .ZN(n6340) );
  OR2_X1 U3841 ( .A1(n6458), .A2(n3882), .ZN(n6368) );
  INV_X1 U3842 ( .A(n3449), .ZN(n5966) );
  INV_X1 U3843 ( .A(n6087), .ZN(n5424) );
  OR4_X1 U3844 ( .A1(n5581), .A2(n6575), .A3(n6571), .A4(n6572), .ZN(n5455) );
  AND2_X1 U3845 ( .A1(n5591), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5696) );
  INV_X1 U3846 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5685) );
  INV_X1 U3847 ( .A(n5667), .ZN(n5612) );
  CLKBUF_X1 U3848 ( .A(n4996), .Z(n4968) );
  INV_X1 U3849 ( .A(n5811), .ZN(n5097) );
  NAND2_X1 U3850 ( .A1(n4445), .A2(n4444), .ZN(n5204) );
  AND2_X1 U3851 ( .A1(n4306), .A2(n4305), .ZN(n5768) );
  CLKBUF_X1 U3852 ( .A(n5769), .Z(n6613) );
  INV_X1 U3853 ( .A(n5762), .ZN(n5775) );
  INV_X1 U3854 ( .A(n4445), .ZN(n5801) );
  OAI21_X1 U3855 ( .B1(n5040), .B2(n5030), .A(n5029), .ZN(n5238) );
  AND2_X1 U3856 ( .A1(n5273), .A2(n5272), .ZN(n5275) );
  XNOR2_X1 U3857 ( .A(n5176), .B(n5066), .ZN(n5499) );
  INV_X1 U3858 ( .A(n5468), .ZN(n5505) );
  AND2_X1 U3859 ( .A1(n5191), .A2(n5190), .ZN(n5734) );
  INV_X1 U3860 ( .A(n5856), .ZN(n5810) );
  INV_X1 U3861 ( .A(n5293), .ZN(n5294) );
  NAND2_X1 U3862 ( .A1(n4535), .A2(n4534), .ZN(n5914) );
  INV_X1 U3863 ( .A(n4702), .ZN(n4339) );
  CLKBUF_X1 U3864 ( .A(n4493), .Z(n6151) );
  BUF_X1 U3865 ( .A(n4488), .Z(n6216) );
  CLKBUF_X1 U3866 ( .A(n3635), .Z(n4732) );
  INV_X1 U3867 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3205) );
  NAND2_X1 U3868 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4317), .ZN(n5009) );
  OAI21_X1 U3869 ( .B1(n6109), .B2(n6600), .A(n6093), .ZN(n6110) );
  INV_X1 U3870 ( .A(n6266), .ZN(n6623) );
  INV_X1 U3871 ( .A(n6335), .ZN(n6324) );
  INV_X1 U3872 ( .A(n6441), .ZN(n6510) );
  INV_X1 U3873 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6517) );
  AOI211_X1 U3874 ( .C1(n5376), .C2(n5687), .A(n4245), .B(n4244), .ZN(n4246)
         );
  INV_X1 U3875 ( .A(n5026), .ZN(n4922) );
  OAI211_X1 U3876 ( .C1(n5856), .C2(n4998), .A(n4997), .B(n3195), .ZN(n4999)
         );
  AND2_X1 U3877 ( .A1(n3877), .A2(n3876), .ZN(n3878) );
  AND4_X1 U3878 ( .A1(n3343), .A2(n3342), .A3(n3711), .A4(n3341), .ZN(n3192)
         );
  NAND2_X1 U3879 ( .A1(n5081), .A2(n5080), .ZN(n5079) );
  NOR2_X1 U3880 ( .A1(n4021), .A2(n4620), .ZN(n3193) );
  INV_X2 U3881 ( .A(n5912), .ZN(n5931) );
  NOR2_X2 U3882 ( .A1(n6545), .A2(n6609), .ZN(n6585) );
  OR2_X1 U3883 ( .A1(n3196), .A2(n3618), .ZN(n3194) );
  NAND2_X1 U3884 ( .A1(n3615), .A2(n4688), .ZN(n3196) );
  AND4_X1 U3885 ( .A1(n3209), .A2(n3208), .A3(n3207), .A4(n3206), .ZN(n3197)
         );
  AND4_X1 U3886 ( .A1(n3252), .A2(n3251), .A3(n3250), .A4(n3249), .ZN(n3198)
         );
  AND4_X1 U3887 ( .A1(n3216), .A2(n3215), .A3(n3214), .A4(n3213), .ZN(n3199)
         );
  AND4_X1 U3888 ( .A1(n3240), .A2(n3239), .A3(n3238), .A4(n3237), .ZN(n3200)
         );
  AND4_X1 U3889 ( .A1(n3248), .A2(n3247), .A3(n3246), .A4(n3245), .ZN(n3201)
         );
  INV_X2 U3890 ( .A(n3606), .ZN(n3620) );
  NOR2_X1 U3891 ( .A1(n4249), .A2(n4734), .ZN(n3202) );
  AND4_X1 U3892 ( .A1(n3244), .A2(n3243), .A3(n3242), .A4(n3241), .ZN(n3203)
         );
  INV_X1 U3893 ( .A(n4551), .ZN(n3970) );
  NAND3_X1 U3894 ( .A1(n3631), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n3632), .ZN(n3204) );
  INV_X1 U3895 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4747) );
  INV_X1 U3896 ( .A(n3683), .ZN(n3660) );
  AND2_X1 U3897 ( .A1(n3639), .A2(n3638), .ZN(n3658) );
  OR2_X1 U3898 ( .A1(n3549), .A2(n3548), .ZN(n3550) );
  NAND2_X1 U3899 ( .A1(n3515), .A2(n6087), .ZN(n3535) );
  INV_X1 U3900 ( .A(n3379), .ZN(n3506) );
  NAND2_X1 U3901 ( .A1(n3884), .A2(n6517), .ZN(n3463) );
  NOR2_X1 U3902 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3212) );
  INV_X1 U3903 ( .A(n3838), .ZN(n3321) );
  OR2_X1 U3904 ( .A1(n3412), .A2(n3411), .ZN(n3595) );
  INV_X1 U3905 ( .A(n3356), .ZN(n3360) );
  INV_X1 U3906 ( .A(n3465), .ZN(n3466) );
  NAND2_X1 U3907 ( .A1(n5941), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3491) );
  INV_X1 U3908 ( .A(n4277), .ZN(n4282) );
  AND2_X2 U3909 ( .A1(n3211), .A2(n4474), .ZN(n4896) );
  INV_X1 U3910 ( .A(n4184), .ZN(n4135) );
  INV_X1 U3911 ( .A(n4552), .ZN(n4022) );
  OAI21_X1 U3912 ( .B1(n3913), .B2(n4070), .A(n3912), .ZN(n4501) );
  NAND2_X1 U3913 ( .A1(n3322), .A2(n3321), .ZN(n3705) );
  AND2_X1 U3914 ( .A1(n3616), .A2(n4252), .ZN(n5302) );
  NAND2_X1 U3915 ( .A1(n5960), .A2(n3449), .ZN(n3838) );
  NAND2_X1 U3916 ( .A1(n3360), .A2(n3359), .ZN(n3383) );
  OR2_X1 U3917 ( .A1(n3467), .A2(n3466), .ZN(n3468) );
  OR2_X1 U3918 ( .A1(n4917), .A2(n5018), .ZN(n4223) );
  NOR2_X1 U3919 ( .A1(n4297), .A2(n4307), .ZN(n4276) );
  INV_X1 U3920 ( .A(n4233), .ZN(n3805) );
  XNOR2_X1 U3921 ( .A(n3594), .B(n3582), .ZN(n3932) );
  OR2_X1 U3922 ( .A1(n4488), .A2(n4070), .ZN(n3895) );
  OR2_X1 U3923 ( .A1(n4886), .A2(n4885), .ZN(n4917) );
  OR2_X1 U3924 ( .A1(n4218), .A2(n5178), .ZN(n4802) );
  NOR2_X1 U3925 ( .A1(n4056), .A2(n5614), .ZN(n4072) );
  INV_X1 U3926 ( .A(n4539), .ZN(n3971) );
  INV_X1 U3927 ( .A(n4070), .ZN(n4052) );
  NOR2_X1 U3928 ( .A1(n5251), .A2(n5235), .ZN(n4983) );
  AND2_X1 U3929 ( .A1(n5419), .A2(n3855), .ZN(n5355) );
  AND2_X1 U3930 ( .A1(n3617), .A2(n5302), .ZN(n4737) );
  AND2_X1 U3931 ( .A1(n5804), .A2(n3607), .ZN(n3608) );
  AND2_X1 U3932 ( .A1(n3759), .A2(n3758), .ZN(n5636) );
  AND2_X1 U3933 ( .A1(n3739), .A2(n3738), .ZN(n5128) );
  NAND2_X1 U3934 ( .A1(n3334), .A2(n3333), .ZN(n3416) );
  NAND2_X1 U3935 ( .A1(n3365), .A2(n3364), .ZN(n4478) );
  AND2_X1 U3936 ( .A1(n5998), .A2(n6466), .ZN(n6246) );
  NAND2_X1 U3937 ( .A1(n3469), .A2(n3468), .ZN(n3882) );
  NAND2_X1 U3938 ( .A1(n3505), .A2(n3504), .ZN(n6087) );
  OR2_X1 U3939 ( .A1(n4791), .A2(n5269), .ZN(n4825) );
  XNOR2_X1 U3940 ( .A(n4223), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4992)
         );
  NAND2_X1 U3941 ( .A1(n4227), .A2(n4226), .ZN(n5667) );
  NAND2_X1 U3942 ( .A1(n5591), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5112) );
  AND2_X1 U3943 ( .A1(n5357), .A2(n5356), .ZN(n5358) );
  AND2_X1 U3944 ( .A1(n5540), .A2(n5539), .ZN(n5542) );
  XNOR2_X1 U3945 ( .A(n4967), .B(n4966), .ZN(n4996) );
  NOR2_X1 U3946 ( .A1(n5191), .A2(n4802), .ZN(n5158) );
  NAND2_X1 U3947 ( .A1(n4679), .A2(n4678), .ZN(n4677) );
  NOR2_X1 U3948 ( .A1(n3954), .A2(n3950), .ZN(n3972) );
  AOI21_X1 U3949 ( .B1(n3931), .B2(n4052), .A(n3930), .ZN(n4522) );
  OAI21_X1 U3950 ( .B1(n4433), .B2(n4434), .A(n4435), .ZN(n3897) );
  NOR2_X1 U3951 ( .A1(n3632), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4982)
         );
  NOR2_X1 U3952 ( .A1(n5250), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5233)
         );
  OAI21_X1 U3953 ( .B1(n3622), .B2(n3621), .A(n3620), .ZN(n3623) );
  OAI21_X1 U3954 ( .B1(n3620), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5285), 
        .ZN(n5279) );
  AND2_X1 U3955 ( .A1(n4741), .A2(n4740), .ZN(n5404) );
  OR2_X1 U3956 ( .A1(n4933), .A2(n4934), .ZN(n5303) );
  OAI21_X1 U3957 ( .B1(n5805), .B2(n3609), .A(n3608), .ZN(n4686) );
  NOR2_X2 U3958 ( .A1(n4528), .A2(n4529), .ZN(n4543) );
  NOR2_X1 U3959 ( .A1(n4700), .A2(n4339), .ZN(n5868) );
  OR2_X1 U3960 ( .A1(n3859), .A2(n4457), .ZN(n5897) );
  XNOR2_X1 U3961 ( .A(n3416), .B(n3415), .ZN(n3884) );
  OR2_X1 U3962 ( .A1(n6217), .A2(n5944), .ZN(n6052) );
  INV_X1 U3963 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6370) );
  INV_X1 U3964 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4724) );
  NOR2_X1 U3965 ( .A1(n4825), .A2(n4824), .ZN(n4847) );
  INV_X1 U3966 ( .A(n4232), .ZN(n5165) );
  NOR2_X2 U3967 ( .A1(n4935), .A2(n4263), .ZN(n5081) );
  AND2_X1 U3968 ( .A1(n4992), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4224) );
  CLKBUF_X1 U3969 ( .A(n4388), .Z(n5143) );
  INV_X1 U3970 ( .A(n5720), .ZN(n5730) );
  NAND2_X1 U3971 ( .A1(n3939), .A2(n3938), .ZN(n4526) );
  INV_X1 U3972 ( .A(n5803), .ZN(n5797) );
  OR2_X1 U3973 ( .A1(n4395), .A2(n4277), .ZN(n4299) );
  XOR2_X1 U3974 ( .A(n5159), .B(n5158), .Z(n5493) );
  INV_X1 U3975 ( .A(n5158), .ZN(n4219) );
  AND2_X1 U3976 ( .A1(n5179), .A2(n5174), .ZN(n5176) );
  AND2_X1 U3977 ( .A1(n4649), .A2(n4634), .ZN(n5811) );
  NAND2_X1 U3978 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n3934), .ZN(n3954)
         );
  NAND2_X1 U3979 ( .A1(n4317), .A2(n6515), .ZN(n4395) );
  OAI22_X1 U3980 ( .A1(n5280), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5279), .B2(n5278), .ZN(n5281) );
  AND2_X1 U3981 ( .A1(n5535), .A2(n3864), .ZN(n5419) );
  OR2_X1 U3982 ( .A1(n3859), .A2(n3835), .ZN(n5903) );
  INV_X1 U3983 ( .A(n5906), .ZN(n5929) );
  INV_X1 U3984 ( .A(n5903), .ZN(n5927) );
  NAND2_X1 U3985 ( .A1(n3475), .A2(n3474), .ZN(n4336) );
  NAND2_X1 U3986 ( .A1(n6517), .A2(n5940), .ZN(n6221) );
  INV_X1 U3987 ( .A(n6075), .ZN(n6078) );
  NOR2_X1 U3988 ( .A1(n6182), .A2(n6368), .ZN(n6150) );
  OR2_X1 U3989 ( .A1(n6223), .A2(n6222), .ZN(n6240) );
  INV_X1 U3990 ( .A(n6631), .ZN(n6291) );
  OR2_X1 U3991 ( .A1(n6345), .A2(n6344), .ZN(n6364) );
  AND2_X1 U3992 ( .A1(n6459), .A2(n6339), .ZN(n6400) );
  AND2_X1 U3993 ( .A1(n6459), .A2(n6369), .ZN(n6438) );
  INV_X1 U3994 ( .A(n4246), .ZN(n4247) );
  INV_X1 U3995 ( .A(n5687), .ZN(n5711) );
  NAND2_X1 U3996 ( .A1(n5591), .A2(n4224), .ZN(n5479) );
  OR2_X1 U3997 ( .A1(n5176), .A2(n5175), .ZN(n5468) );
  AND2_X1 U3998 ( .A1(n4355), .A2(n6515), .ZN(n5733) );
  INV_X1 U3999 ( .A(n4961), .ZN(n4667) );
  INV_X1 U4000 ( .A(n5229), .ZN(n4685) );
  OR2_X1 U4001 ( .A1(n5768), .A2(n6613), .ZN(n5762) );
  INV_X1 U4002 ( .A(n5768), .ZN(n5777) );
  OR2_X1 U4003 ( .A1(n4299), .A2(n4298), .ZN(n4445) );
  OR2_X1 U4004 ( .A1(n4395), .A2(n4607), .ZN(n5803) );
  NAND2_X1 U4005 ( .A1(n4220), .A2(n4219), .ZN(n5223) );
  OR2_X1 U4006 ( .A1(n4395), .A2(n4596), .ZN(n5814) );
  OR2_X1 U4007 ( .A1(n3859), .A2(n3722), .ZN(n5906) );
  INV_X1 U4008 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4721) );
  NAND2_X1 U4009 ( .A1(n6051), .A2(n6339), .ZN(n6025) );
  NAND2_X1 U4010 ( .A1(n6051), .A2(n6410), .ZN(n6075) );
  NAND2_X1 U4011 ( .A1(n6051), .A2(n6299), .ZN(n6113) );
  INV_X1 U4012 ( .A(n6150), .ZN(n6179) );
  OR2_X1 U4013 ( .A1(n6303), .A2(n6368), .ZN(n6631) );
  INV_X1 U4014 ( .A(n6400), .ZN(n6398) );
  INV_X1 U4015 ( .A(n6438), .ZN(n6448) );
  AND2_X1 U4016 ( .A1(n4609), .A2(n4608), .ZN(n6597) );
  OR2_X1 U4017 ( .A1(n4248), .A2(n4247), .ZN(U2804) );
  NOR2_X4 U4018 ( .A1(n3205), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5012)
         );
  AND2_X2 U4019 ( .A1(n3885), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3211)
         );
  AND2_X2 U4021 ( .A1(n3210), .A2(n4578), .ZN(n3367) );
  AOI22_X1 U4022 ( .A1(n3280), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3209) );
  INV_X2 U4023 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3635) );
  AND2_X2 U4024 ( .A1(n5012), .A2(n4729), .ZN(n4765) );
  AOI22_X1 U4025 ( .A1(n4765), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3427), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3208) );
  AND2_X2 U4026 ( .A1(n5012), .A2(n4578), .ZN(n3399) );
  AND2_X2 U4027 ( .A1(n4458), .A2(n4578), .ZN(n3428) );
  AOI22_X1 U4028 ( .A1(n3399), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3207) );
  AND2_X2 U4029 ( .A1(n3210), .A2(n4729), .ZN(n3419) );
  AOI22_X1 U4030 ( .A1(n3419), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3206) );
  NOR2_X4 U4031 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4477) );
  AOI22_X1 U4032 ( .A1(n3425), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3426), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3216) );
  AND2_X2 U4033 ( .A1(n4458), .A2(n4477), .ZN(n3497) );
  AOI22_X1 U4034 ( .A1(n3269), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3215) );
  AND2_X2 U4035 ( .A1(n4477), .A2(n4474), .ZN(n3418) );
  AOI22_X1 U4036 ( .A1(n4896), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3214) );
  AND2_X2 U4037 ( .A1(n4729), .A2(n4474), .ZN(n3258) );
  AND2_X2 U4038 ( .A1(n4455), .A2(n3212), .ZN(n3372) );
  AOI22_X1 U4039 ( .A1(n3258), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3213) );
  NAND2_X1 U4040 ( .A1(n4765), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3220) );
  NAND2_X1 U4041 ( .A1(n3269), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3219) );
  NAND2_X1 U4042 ( .A1(n4896), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3218)
         );
  NAND2_X1 U4043 ( .A1(n3427), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U4044 ( .A1(n3419), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3224) );
  BUF_X4 U4045 ( .A(n3258), .Z(n4874) );
  NAND2_X1 U4046 ( .A1(n4874), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3223)
         );
  NAND2_X1 U4047 ( .A1(n3428), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3222) );
  NAND2_X1 U4048 ( .A1(n3372), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U4049 ( .A1(n3425), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3228) );
  NAND2_X1 U4050 ( .A1(n3426), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3227) );
  NAND2_X1 U4051 ( .A1(n3418), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3226)
         );
  NAND2_X1 U4052 ( .A1(n3406), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3225)
         );
  NAND2_X1 U4053 ( .A1(n3367), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3232) );
  NAND2_X1 U4054 ( .A1(n3280), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3231)
         );
  NAND2_X1 U4055 ( .A1(n3399), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3230)
         );
  NAND2_X1 U4056 ( .A1(n3497), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3229) );
  NAND2_X2 U4057 ( .A1(n3347), .A2(n3346), .ZN(n4438) );
  AOI22_X1 U4058 ( .A1(n3419), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4896), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3240) );
  AOI22_X1 U4059 ( .A1(n3280), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3427), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3239) );
  AOI22_X1 U4060 ( .A1(n3367), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3238) );
  AOI22_X1 U4061 ( .A1(n4765), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3237) );
  AOI22_X1 U4062 ( .A1(n3399), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3258), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3244) );
  AOI22_X1 U4063 ( .A1(n3426), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3243) );
  AOI22_X1 U4064 ( .A1(n3425), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3242) );
  AOI22_X1 U4065 ( .A1(n3269), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3241) );
  AOI22_X1 U4066 ( .A1(n3425), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4896), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3248) );
  AOI22_X1 U4067 ( .A1(n4765), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3247) );
  AOI22_X1 U4068 ( .A1(n3269), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3246) );
  AOI22_X1 U4069 ( .A1(n3418), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3245) );
  AOI22_X1 U4070 ( .A1(n3399), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4874), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U4071 ( .A1(n3280), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3251) );
  AOI22_X1 U4072 ( .A1(n3419), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3427), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3250) );
  AOI22_X1 U4073 ( .A1(n3426), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3249) );
  NAND2_X1 U4074 ( .A1(n4438), .A2(n5960), .ZN(n3253) );
  NAND2_X2 U4075 ( .A1(n5982), .A2(n3324), .ZN(n4446) );
  AOI22_X1 U4076 ( .A1(n4765), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3419), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4077 ( .A1(n3280), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3256) );
  AOI22_X1 U4078 ( .A1(n4896), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3427), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3255) );
  AOI22_X1 U4079 ( .A1(n3399), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3254) );
  NAND4_X1 U4080 ( .A1(n3257), .A2(n3256), .A3(n3255), .A4(n3254), .ZN(n3264)
         );
  BUF_X8 U4081 ( .A(n3258), .Z(n4904) );
  AOI22_X1 U4082 ( .A1(n4904), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3262) );
  AOI22_X1 U4083 ( .A1(n3425), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3261) );
  AOI22_X1 U4084 ( .A1(n3426), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3260) );
  AOI22_X1 U4085 ( .A1(n3269), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3259) );
  NAND4_X1 U4086 ( .A1(n3262), .A2(n3261), .A3(n3260), .A4(n3259), .ZN(n3263)
         );
  OR2_X2 U4087 ( .A1(n3264), .A2(n3263), .ZN(n3449) );
  AOI22_X1 U4088 ( .A1(n4765), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3419), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4089 ( .A1(n3280), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3267) );
  AOI22_X1 U4090 ( .A1(n3428), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3266) );
  AOI22_X1 U4091 ( .A1(n4904), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3265) );
  NAND4_X1 U4092 ( .A1(n3268), .A2(n3267), .A3(n3266), .A4(n3265), .ZN(n3275)
         );
  AOI22_X1 U4093 ( .A1(n3425), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4094 ( .A1(n4896), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3427), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U4095 ( .A1(n3399), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3271) );
  AOI22_X1 U4096 ( .A1(n3426), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3270) );
  NAND4_X1 U4097 ( .A1(n3273), .A2(n3272), .A3(n3271), .A4(n3270), .ZN(n3274)
         );
  AOI21_X1 U4098 ( .B1(n4446), .B2(n3449), .A(n5987), .ZN(n3277) );
  NAND2_X1 U4099 ( .A1(n3326), .A2(n3837), .ZN(n3276) );
  AND2_X1 U4100 ( .A1(n3277), .A2(n3276), .ZN(n3278) );
  NAND2_X2 U4101 ( .A1(n3279), .A2(n3278), .ZN(n3344) );
  NAND2_X1 U4102 ( .A1(n4765), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3284) );
  NAND2_X1 U4103 ( .A1(n3399), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3283)
         );
  NAND2_X1 U4104 ( .A1(n3280), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3282)
         );
  NAND2_X1 U4105 ( .A1(n3269), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3281) );
  NAND2_X1 U4106 ( .A1(n3425), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3288) );
  NAND2_X1 U4107 ( .A1(n3426), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3287) );
  NAND2_X1 U4108 ( .A1(n3419), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3286) );
  NAND2_X1 U4109 ( .A1(n3372), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3285) );
  NAND2_X1 U4110 ( .A1(n4896), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3292)
         );
  NAND2_X1 U4111 ( .A1(n3427), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3291) );
  NAND2_X1 U4112 ( .A1(n3497), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3290) );
  NAND2_X1 U4113 ( .A1(n3406), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3289)
         );
  NAND2_X1 U4114 ( .A1(n3367), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3296) );
  NAND2_X1 U4115 ( .A1(n4874), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3295)
         );
  NAND2_X1 U4116 ( .A1(n3428), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3294) );
  NAND2_X1 U4117 ( .A1(n3418), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3293)
         );
  NAND2_X1 U4119 ( .A1(n4765), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3304) );
  NAND2_X1 U4120 ( .A1(n3419), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3303) );
  NAND2_X1 U4121 ( .A1(n4896), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3302)
         );
  NAND2_X1 U4122 ( .A1(n3427), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3301) );
  NAND2_X1 U4123 ( .A1(n3280), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3308)
         );
  NAND2_X1 U4124 ( .A1(n3399), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3307)
         );
  NAND2_X1 U4125 ( .A1(n3367), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3306) );
  NAND2_X1 U4126 ( .A1(n3497), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3305) );
  NAND2_X1 U4127 ( .A1(n3425), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3312) );
  NAND2_X1 U4128 ( .A1(n3269), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3311) );
  NAND2_X1 U4129 ( .A1(n3418), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3310)
         );
  NAND2_X1 U4130 ( .A1(n3406), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3309)
         );
  NAND2_X1 U4131 ( .A1(n3426), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3316) );
  NAND2_X1 U4132 ( .A1(n4874), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3315)
         );
  NAND2_X1 U4133 ( .A1(n3372), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3314) );
  NAND2_X1 U4134 ( .A1(n3428), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3313) );
  NAND2_X1 U4135 ( .A1(n3344), .A2(n4276), .ZN(n3336) );
  OAI211_X1 U4136 ( .C1(n4446), .C2(n3832), .A(n4449), .B(n4438), .ZN(n3338)
         );
  INV_X1 U4137 ( .A(n3338), .ZN(n3322) );
  NAND2_X1 U4138 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6543) );
  OAI21_X1 U4139 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6543), .ZN(n3690) );
  INV_X1 U4140 ( .A(n3690), .ZN(n3323) );
  NOR2_X1 U4141 ( .A1(n4297), .A2(n3323), .ZN(n3349) );
  OAI21_X1 U4142 ( .B1(n3349), .B2(n3645), .A(n5111), .ZN(n3325) );
  NOR2_X2 U4143 ( .A1(n3326), .A2(n5987), .ZN(n3710) );
  INV_X1 U4144 ( .A(n3710), .ZN(n3327) );
  AND2_X2 U4145 ( .A1(n5955), .A2(n3190), .ZN(n4296) );
  NAND2_X1 U4146 ( .A1(n3327), .A2(n4296), .ZN(n3328) );
  AND2_X2 U4147 ( .A1(n5971), .A2(n3645), .ZN(n3648) );
  AND2_X4 U4148 ( .A1(n3449), .A2(n3720), .ZN(n5181) );
  NAND2_X1 U4149 ( .A1(n3648), .A2(n5181), .ZN(n4327) );
  NAND3_X1 U4150 ( .A1(n3336), .A2(n3329), .A3(n3343), .ZN(n3330) );
  NAND2_X1 U4151 ( .A1(n3330), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3332) );
  NAND2_X1 U4152 ( .A1(n3676), .A2(n4446), .ZN(n3331) );
  NAND2_X1 U4153 ( .A1(n3332), .A2(n3331), .ZN(n3354) );
  NAND2_X1 U4154 ( .A1(n3354), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3334) );
  AND2_X1 U4155 ( .A1(n4724), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3716) );
  NOR2_X1 U4156 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n4725) );
  NAND2_X1 U4157 ( .A1(n4725), .A2(n6517), .ZN(n4396) );
  MUX2_X1 U4158 ( .A(n3716), .B(n4396), .S(n6370), .Z(n3333) );
  INV_X1 U4159 ( .A(n5111), .ZN(n4270) );
  INV_X1 U4160 ( .A(n3648), .ZN(n3718) );
  AOI22_X1 U4161 ( .A1(n4270), .A2(n3718), .B1(n4307), .B2(n3837), .ZN(n3335)
         );
  AND2_X1 U4162 ( .A1(n3336), .A2(n3335), .ZN(n3845) );
  NAND2_X1 U4163 ( .A1(n5960), .A2(n5966), .ZN(n3345) );
  NAND2_X1 U4164 ( .A1(n4725), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5559) );
  INV_X1 U4165 ( .A(n5559), .ZN(n6516) );
  OAI211_X1 U4166 ( .C1(n3345), .C2(n3347), .A(n6516), .B(n3191), .ZN(n3337)
         );
  INV_X1 U4167 ( .A(n3337), .ZN(n3342) );
  INV_X1 U4168 ( .A(n4446), .ZN(n3709) );
  NAND2_X1 U4169 ( .A1(n4296), .A2(n3709), .ZN(n3711) );
  NAND2_X1 U4170 ( .A1(n4446), .A2(n3832), .ZN(n3339) );
  NAND2_X1 U4171 ( .A1(n3339), .A2(n3449), .ZN(n3340) );
  OAI21_X1 U4172 ( .B1(n3338), .B2(n3340), .A(n4297), .ZN(n3341) );
  NAND2_X1 U4173 ( .A1(n3845), .A2(n3192), .ZN(n3414) );
  NAND2_X1 U4174 ( .A1(n3648), .A2(n5941), .ZN(n3846) );
  NAND2_X2 U4175 ( .A1(n4286), .A2(n5955), .ZN(n5550) );
  INV_X1 U4176 ( .A(n3345), .ZN(n4352) );
  AND2_X1 U4177 ( .A1(n4276), .A2(n4352), .ZN(n4441) );
  AND2_X1 U4178 ( .A1(n4449), .A2(n3347), .ZN(n4448) );
  NAND2_X1 U4179 ( .A1(n4326), .A2(n4448), .ZN(n3833) );
  NOR2_X1 U4180 ( .A1(n3838), .A2(n3645), .ZN(n3348) );
  NAND2_X1 U4181 ( .A1(n3710), .A2(n3348), .ZN(n4329) );
  INV_X1 U4182 ( .A(n3349), .ZN(n3350) );
  NAND2_X1 U4183 ( .A1(n4282), .A2(n3350), .ZN(n3351) );
  NAND3_X1 U4184 ( .A1(n5550), .A2(n3833), .A3(n3351), .ZN(n3352) );
  NAND2_X1 U4185 ( .A1(n3352), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3356) );
  INV_X1 U4186 ( .A(n4396), .ZN(n3488) );
  XNOR2_X1 U4187 ( .A(n6370), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6406)
         );
  INV_X1 U4188 ( .A(n3716), .ZN(n3487) );
  AND2_X1 U4189 ( .A1(n3487), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3353)
         );
  AOI21_X1 U4190 ( .B1(n3488), .B2(n6406), .A(n3353), .ZN(n3357) );
  NAND2_X1 U4191 ( .A1(n3354), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3355) );
  NAND3_X1 U4192 ( .A1(n3356), .A2(n3357), .A3(n3355), .ZN(n3384) );
  NAND2_X1 U4193 ( .A1(n3385), .A2(n3384), .ZN(n3361) );
  INV_X1 U4194 ( .A(n3357), .ZN(n3358) );
  OR2_X1 U4195 ( .A1(n3358), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3359)
         );
  NAND2_X1 U4196 ( .A1(n3361), .A2(n3383), .ZN(n3365) );
  NAND2_X1 U4197 ( .A1(n3485), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3363) );
  NAND2_X1 U4198 ( .A1(n6212), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6378) );
  NOR2_X1 U4199 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6212), .ZN(n6267)
         );
  NAND2_X1 U4200 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6267), .ZN(n6301) );
  OAI211_X1 U4201 ( .C1(n6213), .C2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n6378), .B(n6301), .ZN(n5948) );
  AOI22_X1 U4202 ( .A1(n3488), .A2(n5948), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3487), .ZN(n3362) );
  NAND2_X1 U4203 ( .A1(n4478), .A2(n3366), .ZN(n4464) );
  INV_X1 U4204 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6936) );
  AOI22_X1 U4205 ( .A1(n4893), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3420), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3371) );
  INV_X1 U4206 ( .A(n3367), .ZN(n5008) );
  AOI22_X1 U4207 ( .A1(n4894), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3370) );
  BUF_X1 U4208 ( .A(n4896), .Z(n4868) );
  AOI22_X1 U4209 ( .A1(n4868), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4210 ( .A1(n4898), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3368) );
  NAND4_X1 U4211 ( .A1(n3371), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n3378)
         );
  AOI22_X1 U4212 ( .A1(n3187), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4213 ( .A1(n4869), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3375) );
  BUF_X1 U4214 ( .A(n3372), .Z(n4903) );
  AOI22_X1 U4215 ( .A1(n4904), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4216 ( .A1(n4905), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3373) );
  NAND4_X1 U4217 ( .A1(n3376), .A2(n3375), .A3(n3374), .A4(n3373), .ZN(n3377)
         );
  OAI22_X2 U4218 ( .A1(n4464), .A2(STATE2_REG_0__SCAN_IN), .B1(n3506), .B2(
        n3492), .ZN(n3382) );
  INV_X1 U4219 ( .A(n3491), .ZN(n3380) );
  NAND2_X1 U4220 ( .A1(n3384), .A2(n3383), .ZN(n3386) );
  XNOR2_X1 U4221 ( .A(n3386), .B(n3385), .ZN(n4493) );
  NAND2_X1 U4222 ( .A1(n4493), .A2(n6517), .ZN(n3398) );
  AOI22_X1 U4223 ( .A1(n4765), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3420), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4224 ( .A1(n4894), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4225 ( .A1(n4896), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4226 ( .A1(n4898), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3387) );
  NAND4_X1 U4227 ( .A1(n3390), .A2(n3389), .A3(n3388), .A4(n3387), .ZN(n3396)
         );
  AOI22_X1 U4228 ( .A1(n3187), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4229 ( .A1(n4869), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4230 ( .A1(n4904), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3392) );
  AOI22_X1 U4231 ( .A1(n4905), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3391) );
  NAND4_X1 U4232 ( .A1(n3394), .A2(n3393), .A3(n3392), .A4(n3391), .ZN(n3395)
         );
  OR2_X1 U4233 ( .A1(n3492), .A2(n3457), .ZN(n3397) );
  NAND2_X2 U4234 ( .A1(n3398), .A2(n3397), .ZN(n3453) );
  AOI22_X1 U4235 ( .A1(n4893), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3420), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4236 ( .A1(n4894), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3402) );
  AOI22_X1 U4237 ( .A1(n4896), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3401) );
  AOI22_X1 U4238 ( .A1(n4898), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3400) );
  NAND4_X1 U4239 ( .A1(n3403), .A2(n3402), .A3(n3401), .A4(n3400), .ZN(n3412)
         );
  INV_X1 U4240 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n6954) );
  AOI22_X1 U4241 ( .A1(n3187), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4243 ( .A1(n4869), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4244 ( .A1(n4904), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3408) );
  AOI22_X1 U4245 ( .A1(n4905), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3407) );
  NAND4_X1 U4246 ( .A1(n3410), .A2(n3409), .A3(n3408), .A4(n3407), .ZN(n3411)
         );
  OR2_X1 U4247 ( .A1(n3492), .A2(n3595), .ZN(n3417) );
  NAND2_X1 U4248 ( .A1(n3676), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3413) );
  OAI211_X1 U4249 ( .C1(n3457), .C2(n3491), .A(n3417), .B(n3413), .ZN(n3452)
         );
  NAND2_X1 U4250 ( .A1(n3453), .A2(n3452), .ZN(n3440) );
  INV_X1 U4251 ( .A(n3414), .ZN(n3415) );
  NAND2_X1 U4252 ( .A1(n5971), .A2(n3595), .ZN(n3437) );
  NOR2_X1 U4253 ( .A1(n3437), .A2(n6517), .ZN(n3592) );
  INV_X1 U4254 ( .A(n3417), .ZN(n3435) );
  AOI22_X1 U4255 ( .A1(n4893), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4868), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3424) );
  INV_X1 U4256 ( .A(n5008), .ZN(n4811) );
  AOI22_X1 U4257 ( .A1(n4894), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4258 ( .A1(n4904), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3422) );
  BUF_X1 U4259 ( .A(n3419), .Z(n3420) );
  AOI22_X1 U4260 ( .A1(n3420), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3421) );
  NAND4_X1 U4261 ( .A1(n3424), .A2(n3423), .A3(n3422), .A4(n3421), .ZN(n3434)
         );
  AOI22_X1 U4262 ( .A1(n4869), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3187), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3432) );
  AOI22_X1 U4263 ( .A1(n4905), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4264 ( .A1(n4898), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4265 ( .A1(n3404), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3429) );
  NAND4_X1 U4266 ( .A1(n3432), .A2(n3431), .A3(n3430), .A4(n3429), .ZN(n3433)
         );
  MUX2_X1 U4267 ( .A(n3592), .B(n3435), .S(n3471), .Z(n3436) );
  INV_X1 U4268 ( .A(n3436), .ZN(n3467) );
  NAND2_X1 U4269 ( .A1(n3463), .A2(n3467), .ZN(n3439) );
  INV_X1 U4270 ( .A(n3676), .ZN(n3672) );
  INV_X1 U4271 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n6930) );
  AOI21_X1 U4272 ( .B1(n5941), .B2(n3471), .A(n6517), .ZN(n3438) );
  OAI211_X1 U4273 ( .C1(n3672), .C2(n6930), .A(n3438), .B(n3437), .ZN(n3465)
         );
  NAND2_X1 U4274 ( .A1(n3440), .A2(n3454), .ZN(n3442) );
  INV_X1 U4275 ( .A(n3443), .ZN(n3446) );
  INV_X1 U4276 ( .A(n3444), .ZN(n3445) );
  NAND2_X1 U4277 ( .A1(n3446), .A2(n3445), .ZN(n3447) );
  INV_X1 U4278 ( .A(n3640), .ZN(n3470) );
  NAND2_X1 U4279 ( .A1(n3448), .A2(n3471), .ZN(n3507) );
  XNOR2_X1 U4280 ( .A(n3507), .B(n3506), .ZN(n3450) );
  AND2_X1 U4281 ( .A1(n5941), .A2(n3449), .ZN(n3472) );
  AOI21_X1 U4282 ( .B1(n3450), .B2(n4296), .A(n3472), .ZN(n3451) );
  NAND2_X1 U4283 ( .A1(n5847), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3481)
         );
  INV_X1 U4284 ( .A(n3454), .ZN(n3455) );
  XNOR2_X2 U4285 ( .A(n3456), .B(n3455), .ZN(n6458) );
  NAND2_X1 U4286 ( .A1(n6458), .A2(n3640), .ZN(n3462) );
  XNOR2_X1 U4287 ( .A(n3457), .B(n3471), .ZN(n3458) );
  NAND2_X1 U4288 ( .A1(n3458), .A2(n4296), .ZN(n3460) );
  NOR2_X1 U4289 ( .A1(n3838), .A2(n5976), .ZN(n3459) );
  AND2_X1 U4290 ( .A1(n3460), .A2(n3459), .ZN(n3461) );
  NAND2_X1 U4291 ( .A1(n3462), .A2(n3461), .ZN(n4382) );
  OR2_X1 U4292 ( .A1(n3882), .A2(n3470), .ZN(n3475) );
  INV_X1 U4293 ( .A(n3471), .ZN(n3473) );
  AOI21_X1 U4294 ( .B1(n3473), .B2(n4296), .A(n3472), .ZN(n3474) );
  AND2_X1 U4295 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3476) );
  NAND2_X1 U4296 ( .A1(n4336), .A2(n3476), .ZN(n3479) );
  NAND2_X1 U4297 ( .A1(n4336), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3477)
         );
  INV_X1 U4298 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4714) );
  NAND2_X1 U4299 ( .A1(n3477), .A2(n4714), .ZN(n3478) );
  AND2_X1 U4300 ( .A1(n3479), .A2(n3478), .ZN(n4383) );
  INV_X1 U4301 ( .A(n3479), .ZN(n3480) );
  AOI21_X1 U4302 ( .B1(n4382), .B2(n4383), .A(n3480), .ZN(n5849) );
  NAND2_X1 U4303 ( .A1(n3481), .A2(n5849), .ZN(n3484) );
  INV_X1 U4304 ( .A(n5847), .ZN(n3482) );
  INV_X1 U4305 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n5932) );
  NAND2_X1 U4306 ( .A1(n3482), .A2(n5932), .ZN(n3483) );
  NAND2_X1 U4307 ( .A1(n3485), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3490) );
  INV_X1 U4308 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6415) );
  NAND3_X1 U4309 ( .A1(n6415), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6187) );
  INV_X1 U4310 ( .A(n6187), .ZN(n6186) );
  NAND2_X1 U4311 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6186), .ZN(n6181) );
  NAND2_X1 U4312 ( .A1(n6415), .A2(n6181), .ZN(n3486) );
  NAND3_X1 U4313 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6453) );
  INV_X1 U4314 ( .A(n6453), .ZN(n6467) );
  NAND2_X1 U4315 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6467), .ZN(n6450) );
  AND2_X1 U4316 ( .A1(n3486), .A2(n6450), .ZN(n6214) );
  AOI22_X1 U4317 ( .A1(n3488), .A2(n6214), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3487), .ZN(n3489) );
  AOI22_X1 U4318 ( .A1(n4893), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3420), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3496) );
  AOI22_X1 U4319 ( .A1(n4898), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4868), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4320 ( .A1(n3187), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4321 ( .A1(n4905), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3493) );
  NAND4_X1 U4322 ( .A1(n3496), .A2(n3495), .A3(n3494), .A4(n3493), .ZN(n3503)
         );
  AOI22_X1 U4323 ( .A1(n4811), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3501) );
  AOI22_X1 U4324 ( .A1(n4894), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4325 ( .A1(n4904), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4326 ( .A1(n4869), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3498) );
  NAND4_X1 U4327 ( .A1(n3501), .A2(n3500), .A3(n3499), .A4(n3498), .ZN(n3502)
         );
  OR2_X1 U4328 ( .A1(n3503), .A2(n3502), .ZN(n3527) );
  AOI22_X1 U4329 ( .A1(n3683), .A2(n3527), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n3676), .ZN(n3504) );
  NAND2_X1 U4330 ( .A1(n3898), .A2(n3640), .ZN(n3511) );
  NAND2_X1 U4331 ( .A1(n3507), .A2(n3506), .ZN(n3528) );
  INV_X1 U4332 ( .A(n3527), .ZN(n3508) );
  XNOR2_X1 U4333 ( .A(n3528), .B(n3508), .ZN(n3509) );
  NAND2_X1 U4334 ( .A1(n3509), .A2(n4296), .ZN(n3510) );
  NAND2_X1 U4335 ( .A1(n3511), .A2(n3510), .ZN(n3512) );
  INV_X1 U4336 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5920) );
  XNOR2_X1 U4337 ( .A(n3512), .B(n5920), .ZN(n4534) );
  NAND2_X1 U4338 ( .A1(n3512), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3513)
         );
  NAND2_X1 U4339 ( .A1(n5914), .A2(n3513), .ZN(n5839) );
  INV_X1 U4340 ( .A(n3514), .ZN(n3515) );
  AOI22_X1 U4341 ( .A1(n4893), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3420), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3519) );
  AOI22_X1 U4342 ( .A1(n4894), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3518) );
  AOI22_X1 U4343 ( .A1(n4868), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4344 ( .A1(n4898), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3516) );
  NAND4_X1 U4345 ( .A1(n3519), .A2(n3518), .A3(n3517), .A4(n3516), .ZN(n3525)
         );
  AOI22_X1 U4346 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3187), .B1(n3404), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U4347 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4869), .B1(n3405), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4348 ( .A1(n4904), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3521) );
  AOI22_X1 U4349 ( .A1(n4905), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3520) );
  NAND4_X1 U4350 ( .A1(n3523), .A2(n3522), .A3(n3521), .A4(n3520), .ZN(n3524)
         );
  OR2_X1 U4351 ( .A1(n3525), .A2(n3524), .ZN(n3552) );
  AOI22_X1 U4352 ( .A1(n3683), .A2(n3552), .B1(INSTQUEUE_REG_0__4__SCAN_IN), 
        .B2(n3676), .ZN(n3534) );
  INV_X1 U4353 ( .A(n3534), .ZN(n3526) );
  XNOR2_X1 U4354 ( .A(n3535), .B(n3526), .ZN(n3914) );
  NAND2_X1 U4355 ( .A1(n3914), .A2(n3640), .ZN(n3531) );
  NAND2_X1 U4356 ( .A1(n3528), .A2(n3527), .ZN(n3554) );
  XNOR2_X1 U4357 ( .A(n3554), .B(n3552), .ZN(n3529) );
  NAND2_X1 U4358 ( .A1(n3529), .A2(n4296), .ZN(n3530) );
  NAND2_X1 U4359 ( .A1(n3531), .A2(n3530), .ZN(n3532) );
  INV_X1 U4360 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5911) );
  XNOR2_X1 U4361 ( .A(n3532), .B(n5911), .ZN(n5838) );
  NAND2_X1 U4362 ( .A1(n5839), .A2(n5838), .ZN(n5841) );
  NAND2_X1 U4363 ( .A1(n3532), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3533)
         );
  NAND2_X1 U4364 ( .A1(n5841), .A2(n3533), .ZN(n5832) );
  AOI22_X1 U4365 ( .A1(n4898), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4366 ( .A1(n3420), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4367 ( .A1(n3404), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4368 ( .A1(n4869), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3536) );
  NAND4_X1 U4369 ( .A1(n3539), .A2(n3538), .A3(n3537), .A4(n3536), .ZN(n3545)
         );
  AOI22_X1 U4370 ( .A1(n4893), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4868), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4371 ( .A1(n3187), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4874), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4372 ( .A1(n4894), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4373 ( .A1(n4905), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3540) );
  NAND4_X1 U4374 ( .A1(n3543), .A2(n3542), .A3(n3541), .A4(n3540), .ZN(n3544)
         );
  OR2_X1 U4375 ( .A1(n3545), .A2(n3544), .ZN(n3573) );
  NAND2_X1 U4376 ( .A1(n3683), .A2(n3573), .ZN(n3547) );
  NAND2_X1 U4377 ( .A1(n3676), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3546) );
  NAND2_X1 U4378 ( .A1(n3547), .A2(n3546), .ZN(n3548) );
  NAND2_X1 U4379 ( .A1(n3549), .A2(n3548), .ZN(n3571) );
  INV_X1 U4380 ( .A(n3913), .ZN(n3551) );
  NAND2_X1 U4381 ( .A1(n3551), .A2(n3640), .ZN(n3557) );
  INV_X1 U4382 ( .A(n3552), .ZN(n3553) );
  OR2_X1 U4383 ( .A1(n3554), .A2(n3553), .ZN(n3572) );
  XNOR2_X1 U4384 ( .A(n3572), .B(n3573), .ZN(n3555) );
  NAND2_X1 U4385 ( .A1(n3555), .A2(n4296), .ZN(n3556) );
  NAND2_X1 U4386 ( .A1(n3557), .A2(n3556), .ZN(n3558) );
  INV_X1 U4387 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5887) );
  XNOR2_X1 U4388 ( .A(n3558), .B(n5887), .ZN(n5831) );
  NAND2_X1 U4389 ( .A1(n5832), .A2(n5831), .ZN(n5830) );
  NAND2_X1 U4390 ( .A1(n3558), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3559)
         );
  NAND2_X1 U4391 ( .A1(n5830), .A2(n3559), .ZN(n4510) );
  AOI22_X1 U4392 ( .A1(n4893), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3420), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4393 ( .A1(n4894), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4394 ( .A1(n4868), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4395 ( .A1(n4898), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3560) );
  NAND4_X1 U4396 ( .A1(n3563), .A2(n3562), .A3(n3561), .A4(n3560), .ZN(n3569)
         );
  AOI22_X1 U4397 ( .A1(n3187), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3567) );
  AOI22_X1 U4398 ( .A1(n4869), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4399 ( .A1(n4904), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4400 ( .A1(n4905), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3564) );
  NAND4_X1 U4401 ( .A1(n3567), .A2(n3566), .A3(n3565), .A4(n3564), .ZN(n3568)
         );
  OR2_X1 U4402 ( .A1(n3569), .A2(n3568), .ZN(n3584) );
  AOI22_X1 U4403 ( .A1(n3683), .A2(n3584), .B1(n3676), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3570) );
  NAND2_X1 U4404 ( .A1(n3571), .A2(n3570), .ZN(n3931) );
  NAND3_X1 U4405 ( .A1(n3594), .A2(n3931), .A3(n3640), .ZN(n3577) );
  INV_X1 U4406 ( .A(n3572), .ZN(n3574) );
  NAND2_X1 U4407 ( .A1(n3574), .A2(n3573), .ZN(n3583) );
  XNOR2_X1 U4408 ( .A(n3583), .B(n3584), .ZN(n3575) );
  NAND2_X1 U4409 ( .A1(n3575), .A2(n4296), .ZN(n3576) );
  NAND2_X1 U4410 ( .A1(n3577), .A2(n3576), .ZN(n3578) );
  INV_X1 U4411 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3850) );
  XNOR2_X1 U4412 ( .A(n3578), .B(n3850), .ZN(n4509) );
  NAND2_X1 U4413 ( .A1(n4510), .A2(n4509), .ZN(n4508) );
  NAND2_X1 U4414 ( .A1(n3578), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3579)
         );
  NAND2_X1 U4415 ( .A1(n4508), .A2(n3579), .ZN(n5817) );
  NAND2_X1 U4416 ( .A1(n3683), .A2(n3595), .ZN(n3581) );
  NAND2_X1 U4417 ( .A1(n3676), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3580) );
  NAND2_X1 U4418 ( .A1(n3581), .A2(n3580), .ZN(n3582) );
  NAND2_X1 U4419 ( .A1(n3932), .A2(n3640), .ZN(n3588) );
  INV_X1 U4420 ( .A(n3583), .ZN(n3585) );
  NAND2_X1 U4421 ( .A1(n3585), .A2(n3584), .ZN(n3597) );
  XNOR2_X1 U4422 ( .A(n3597), .B(n3595), .ZN(n3586) );
  NAND2_X1 U4423 ( .A1(n3586), .A2(n4296), .ZN(n3587) );
  NAND2_X1 U4424 ( .A1(n3588), .A2(n3587), .ZN(n3590) );
  INV_X1 U4425 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3589) );
  XNOR2_X1 U4426 ( .A(n3590), .B(n3589), .ZN(n5816) );
  NAND2_X1 U4427 ( .A1(n5817), .A2(n5816), .ZN(n5815) );
  NAND2_X1 U4428 ( .A1(n3590), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3591)
         );
  NAND2_X1 U4429 ( .A1(n5815), .A2(n3591), .ZN(n4557) );
  AND2_X1 U4430 ( .A1(n3592), .A2(n3640), .ZN(n3593) );
  NAND2_X1 U4431 ( .A1(n4296), .A2(n3595), .ZN(n3596) );
  OR2_X1 U4432 ( .A1(n3597), .A2(n3596), .ZN(n3598) );
  NAND2_X1 U4433 ( .A1(n5304), .A2(n3598), .ZN(n3599) );
  INV_X1 U4434 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6931) );
  XNOR2_X1 U4435 ( .A(n3599), .B(n6931), .ZN(n4556) );
  NAND2_X1 U4436 ( .A1(n4557), .A2(n4556), .ZN(n4555) );
  NAND2_X1 U4437 ( .A1(n3599), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3600)
         );
  NAND2_X1 U4438 ( .A1(n4555), .A2(n3600), .ZN(n4625) );
  INV_X1 U4439 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4626) );
  NAND2_X1 U4440 ( .A1(n5304), .A2(n4626), .ZN(n3601) );
  NAND2_X1 U4441 ( .A1(n4625), .A2(n3601), .ZN(n3603) );
  NAND2_X1 U4442 ( .A1(n3620), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3602)
         );
  NAND2_X1 U4443 ( .A1(n3603), .A2(n3602), .ZN(n4642) );
  INV_X1 U4444 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3604) );
  NAND2_X1 U4445 ( .A1(n5304), .A2(n3604), .ZN(n4643) );
  NAND2_X1 U4446 ( .A1(n4642), .A2(n4643), .ZN(n5805) );
  INV_X1 U4447 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3605) );
  AND2_X1 U4448 ( .A1(n5304), .A2(n3605), .ZN(n3609) );
  NAND2_X1 U4449 ( .A1(n3620), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U4450 ( .A1(n3620), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3607) );
  INV_X1 U4451 ( .A(n4686), .ZN(n4251) );
  INV_X1 U4452 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4951) );
  NOR2_X1 U4453 ( .A1(n5806), .A2(n4951), .ZN(n5515) );
  XNOR2_X1 U4454 ( .A(n5806), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5519)
         );
  INV_X1 U4455 ( .A(n5519), .ZN(n3610) );
  AND2_X1 U4456 ( .A1(n3620), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4691)
         );
  INV_X1 U4457 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6888) );
  XNOR2_X1 U4458 ( .A(n5806), .B(n6888), .ZN(n4934) );
  INV_X1 U4459 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5534) );
  INV_X1 U4460 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4262) );
  NAND3_X1 U4461 ( .A1(n5534), .A2(n5527), .A3(n4262), .ZN(n3611) );
  AND2_X1 U4462 ( .A1(n3620), .A2(n3611), .ZN(n3612) );
  INV_X1 U4463 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4711) );
  INV_X1 U4464 ( .A(n4690), .ZN(n3615) );
  NAND2_X1 U4465 ( .A1(n5304), .A2(n4951), .ZN(n5517) );
  INV_X1 U4466 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3613) );
  NAND2_X1 U4467 ( .A1(n5304), .A2(n3613), .ZN(n3614) );
  NAND2_X1 U4468 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3854) );
  NAND2_X1 U4469 ( .A1(n5304), .A2(n3854), .ZN(n3617) );
  NAND2_X1 U4470 ( .A1(n5304), .A2(n4262), .ZN(n3616) );
  NAND2_X1 U4471 ( .A1(n5304), .A2(n6888), .ZN(n4252) );
  INV_X1 U4472 ( .A(n4737), .ZN(n3618) );
  NAND2_X1 U4473 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5408) );
  NAND2_X1 U4474 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3868) );
  NOR2_X1 U4475 ( .A1(n5408), .A2(n3868), .ZN(n5377) );
  AND2_X1 U4476 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3871) );
  AND2_X1 U4477 ( .A1(n5377), .A2(n3871), .ZN(n3855) );
  NAND2_X1 U4478 ( .A1(n3622), .A2(n3855), .ZN(n3624) );
  NOR2_X1 U4479 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5409) );
  NOR2_X1 U4480 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3619) );
  INV_X1 U4481 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5397) );
  INV_X1 U4482 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5385) );
  NAND4_X1 U4483 ( .A1(n5409), .A2(n3619), .A3(n5397), .A4(n5385), .ZN(n3621)
         );
  NAND2_X1 U4484 ( .A1(n3624), .A2(n3623), .ZN(n5266) );
  INV_X1 U4485 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3625) );
  XNOR2_X1 U4486 ( .A(n5806), .B(n3625), .ZN(n5267) );
  OR2_X2 U4487 ( .A1(n5266), .A2(n5267), .ZN(n5264) );
  NAND2_X1 U4488 ( .A1(n5304), .A2(n3625), .ZN(n3626) );
  NAND2_X1 U4489 ( .A1(n5264), .A2(n3626), .ZN(n5259) );
  INV_X1 U4490 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6782) );
  NAND2_X1 U4491 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U4492 ( .A1(n4983), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3631) );
  OR2_X2 U4493 ( .A1(n5264), .A2(n3629), .ZN(n5250) );
  INV_X1 U4494 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3821) );
  INV_X1 U4495 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5236) );
  AND2_X1 U4496 ( .A1(n3821), .A2(n5236), .ZN(n3630) );
  INV_X1 U4497 ( .A(n3631), .ZN(n3633) );
  INV_X1 U4498 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3856) );
  AOI21_X1 U4499 ( .B1(n3633), .B2(n3856), .A(n4982), .ZN(n3634) );
  NAND2_X1 U4500 ( .A1(n6212), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3637) );
  NAND2_X1 U4501 ( .A1(n4732), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3636) );
  NAND2_X1 U4502 ( .A1(n3637), .A2(n3636), .ZN(n3641) );
  NAND2_X1 U4503 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6370), .ZN(n3644) );
  NAND2_X1 U4504 ( .A1(n3643), .A2(n3637), .ZN(n3659) );
  NAND2_X1 U4505 ( .A1(n6213), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3639) );
  NAND2_X1 U4506 ( .A1(n4721), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3638) );
  NAND2_X1 U4507 ( .A1(n3659), .A2(n3658), .ZN(n3657) );
  NAND2_X1 U4508 ( .A1(n3657), .A2(n3639), .ZN(n3669) );
  XNOR2_X1 U4509 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3668) );
  AOI21_X1 U4510 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6415), .A(n3671), 
        .ZN(n3682) );
  INV_X1 U4511 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5553) );
  NAND3_X1 U4512 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3682), .A3(n5553), .ZN(n3695) );
  NAND2_X1 U4513 ( .A1(n3676), .A2(n3640), .ZN(n3686) );
  OAI21_X1 U4514 ( .B1(n3660), .B2(n5955), .A(n3645), .ZN(n3655) );
  NAND2_X1 U4515 ( .A1(n3641), .A2(n3644), .ZN(n3642) );
  NAND2_X1 U4516 ( .A1(n3643), .A2(n3642), .ZN(n3692) );
  INV_X1 U4517 ( .A(n3692), .ZN(n3652) );
  OAI21_X1 U4518 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6370), .A(n3644), 
        .ZN(n3647) );
  NOR2_X1 U4519 ( .A1(n3660), .A2(n3647), .ZN(n3650) );
  AND2_X1 U4520 ( .A1(n5955), .A2(n3645), .ZN(n3646) );
  NOR2_X1 U4521 ( .A1(n4276), .A2(n3646), .ZN(n3665) );
  OAI21_X1 U4522 ( .B1(n3648), .B2(n3647), .A(n3190), .ZN(n3649) );
  NAND2_X1 U4523 ( .A1(n3665), .A2(n3649), .ZN(n3651) );
  OAI211_X1 U4524 ( .C1(n3655), .C2(n3652), .A(n3650), .B(n3651), .ZN(n3654)
         );
  INV_X1 U4525 ( .A(n3651), .ZN(n3653) );
  AOI22_X1 U4526 ( .A1(n3686), .A2(n3654), .B1(n3653), .B2(n3652), .ZN(n3664)
         );
  INV_X1 U4527 ( .A(n3655), .ZN(n3656) );
  NOR3_X1 U4528 ( .A1(n3656), .A2(n6517), .A3(n3692), .ZN(n3663) );
  OAI21_X1 U4529 ( .B1(n3659), .B2(n3658), .A(n3657), .ZN(n3691) );
  NOR2_X1 U4530 ( .A1(n3660), .A2(n3691), .ZN(n3667) );
  INV_X1 U4531 ( .A(n3691), .ZN(n3661) );
  OAI21_X1 U4532 ( .B1(n3661), .B2(n3672), .A(n3665), .ZN(n3662) );
  OAI22_X1 U4533 ( .A1(n3664), .A2(n3663), .B1(n3667), .B2(n3662), .ZN(n3674)
         );
  INV_X1 U4534 ( .A(n3665), .ZN(n3666) );
  NAND2_X1 U4535 ( .A1(n3667), .A2(n3666), .ZN(n3673) );
  NOR2_X1 U4536 ( .A1(n3669), .A2(n3668), .ZN(n3670) );
  OR2_X1 U4537 ( .A1(n3671), .A2(n3670), .ZN(n3693) );
  AOI22_X1 U4538 ( .A1(n3674), .A2(n3673), .B1(n3672), .B2(n3693), .ZN(n3678)
         );
  INV_X1 U4539 ( .A(n3693), .ZN(n3675) );
  NOR2_X1 U4540 ( .A1(n3686), .A2(n3675), .ZN(n3677) );
  OAI22_X1 U4541 ( .A1(n3678), .A2(n3677), .B1(n3676), .B2(n3695), .ZN(n3679)
         );
  OAI21_X1 U4542 ( .B1(n3695), .B2(n3686), .A(n3679), .ZN(n3680) );
  AOI21_X1 U4543 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6517), .A(n3680), 
        .ZN(n3685) );
  INV_X1 U4544 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6972) );
  NOR2_X1 U4545 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6972), .ZN(n3681)
         );
  AOI221_X1 U4546 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n3682), .C1(
        n5553), .C2(n3682), .A(n3681), .ZN(n3694) );
  NAND2_X1 U4547 ( .A1(n3694), .A2(n3683), .ZN(n3684) );
  NAND2_X1 U4548 ( .A1(n3685), .A2(n3684), .ZN(n3689) );
  INV_X1 U4549 ( .A(n3686), .ZN(n3687) );
  NAND2_X1 U4550 ( .A1(n3694), .A2(n3687), .ZN(n3688) );
  AND2_X1 U4551 ( .A1(n3709), .A2(n3832), .ZN(n4580) );
  NAND2_X1 U4552 ( .A1(n4580), .A2(n4297), .ZN(n3848) );
  NOR2_X1 U4553 ( .A1(n4317), .A2(n3848), .ZN(n4324) );
  INV_X1 U4554 ( .A(n4324), .ZN(n3715) );
  OR2_X1 U4555 ( .A1(n3690), .A2(STATE_REG_0__SCAN_IN), .ZN(n6533) );
  NAND2_X1 U4556 ( .A1(n4297), .A2(n6533), .ZN(n3698) );
  NOR3_X1 U4557 ( .A1(n3693), .A2(n3692), .A3(n3691), .ZN(n3696) );
  AOI21_X1 U4558 ( .B1(n3696), .B2(n3695), .A(n3694), .ZN(n4288) );
  INV_X1 U4559 ( .A(n4288), .ZN(n3697) );
  NOR2_X1 U4560 ( .A1(n3697), .A2(READY_N), .ZN(n4318) );
  NAND2_X1 U4561 ( .A1(n3698), .A2(n4318), .ZN(n3704) );
  INV_X1 U4562 ( .A(n6533), .ZN(n4305) );
  INV_X1 U4563 ( .A(n4296), .ZN(n6615) );
  OAI21_X1 U4564 ( .B1(n4329), .B2(READY_N), .A(n4307), .ZN(n3699) );
  OAI21_X1 U4565 ( .B1(n4305), .B2(n6615), .A(n3699), .ZN(n3701) );
  INV_X1 U4566 ( .A(n4448), .ZN(n3700) );
  NAND2_X1 U4567 ( .A1(n3701), .A2(n3700), .ZN(n3702) );
  NAND2_X1 U4568 ( .A1(n4317), .A2(n3702), .ZN(n3703) );
  MUX2_X1 U4569 ( .A(n3704), .B(n3703), .S(n5960), .Z(n3714) );
  INV_X1 U4570 ( .A(n3705), .ZN(n3708) );
  INV_X1 U4571 ( .A(n4580), .ZN(n3706) );
  NAND2_X1 U4572 ( .A1(n3706), .A2(n5941), .ZN(n3707) );
  NAND2_X1 U4573 ( .A1(n3708), .A2(n3707), .ZN(n3719) );
  OR3_X1 U4574 ( .A1(n3710), .A2(n5941), .A3(n3709), .ZN(n3712) );
  NAND2_X1 U4575 ( .A1(n3712), .A2(n3711), .ZN(n3843) );
  NOR2_X1 U4576 ( .A1(n3719), .A2(n3843), .ZN(n3713) );
  OR2_X1 U4577 ( .A1(n3713), .A2(n4286), .ZN(n4314) );
  NAND3_X1 U4578 ( .A1(n3715), .A2(n3714), .A3(n4314), .ZN(n3717) );
  AND2_X1 U4579 ( .A1(n3716), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6515) );
  INV_X1 U4580 ( .A(n4276), .ZN(n5108) );
  NOR2_X1 U4581 ( .A1(n3719), .A2(n5108), .ZN(n4316) );
  INV_X1 U4582 ( .A(n4316), .ZN(n4456) );
  OR2_X1 U4583 ( .A1(n3719), .A2(n3718), .ZN(n4596) );
  NAND2_X1 U4584 ( .A1(n4456), .A2(n4596), .ZN(n4283) );
  INV_X1 U4585 ( .A(n5550), .ZN(n4319) );
  NAND2_X4 U4586 ( .A1(n3189), .A2(n3720), .ZN(n3734) );
  OR2_X1 U4587 ( .A1(n4329), .A2(n3734), .ZN(n4310) );
  OAI21_X1 U4588 ( .B1(n5971), .B2(n3833), .A(n4310), .ZN(n3721) );
  NOR3_X1 U4589 ( .A1(n4283), .A2(n4319), .A3(n3721), .ZN(n3722) );
  INV_X1 U4590 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3724) );
  AND2_X1 U4591 ( .A1(n5181), .A2(n3724), .ZN(n3723) );
  INV_X4 U4592 ( .A(n3734), .ZN(n4390) );
  NAND2_X1 U4593 ( .A1(n3723), .A2(n4390), .ZN(n3728) );
  NAND2_X1 U4594 ( .A1(n3732), .A2(n4714), .ZN(n3726) );
  NAND2_X1 U4595 ( .A1(n4390), .A2(n3724), .ZN(n3725) );
  NAND3_X1 U4596 ( .A1(n3726), .A2(n5170), .A3(n3725), .ZN(n3727) );
  NAND2_X1 U4597 ( .A1(n3728), .A2(n3727), .ZN(n3731) );
  NAND2_X1 U4598 ( .A1(n3732), .A2(EBX_REG_0__SCAN_IN), .ZN(n3730) );
  INV_X1 U4599 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4356) );
  NAND2_X1 U4600 ( .A1(n5170), .A2(n4356), .ZN(n3729) );
  NAND2_X1 U4601 ( .A1(n3730), .A2(n3729), .ZN(n4340) );
  XNOR2_X1 U4602 ( .A(n3731), .B(n4340), .ZN(n4388) );
  NAND2_X1 U4603 ( .A1(n4388), .A2(n4390), .ZN(n4389) );
  NAND2_X1 U4604 ( .A1(n4389), .A2(n3731), .ZN(n4422) );
  NAND2_X2 U4605 ( .A1(n3191), .A2(n3188), .ZN(n4930) );
  NAND2_X1 U4606 ( .A1(n4390), .A2(n5170), .ZN(n3819) );
  MUX2_X1 U4607 ( .A(n3819), .B(n3188), .S(EBX_REG_3__SCAN_IN), .Z(n3733) );
  OAI21_X1 U4608 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n4930), .A(n3733), 
        .ZN(n4423) );
  INV_X1 U4609 ( .A(n5181), .ZN(n3735) );
  OR2_X2 U4610 ( .A1(n3735), .A2(n3734), .ZN(n4925) );
  INV_X1 U4611 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6933) );
  NAND2_X1 U4612 ( .A1(n3824), .A2(n6933), .ZN(n3739) );
  NAND2_X1 U4613 ( .A1(n3191), .A2(n5932), .ZN(n3737) );
  NAND2_X1 U4614 ( .A1(n4390), .A2(n6933), .ZN(n3736) );
  NAND3_X1 U4615 ( .A1(n3737), .A2(n3188), .A3(n3736), .ZN(n3738) );
  OR3_X2 U4616 ( .A1(n4422), .A2(n4423), .A3(n5128), .ZN(n4428) );
  INV_X1 U4617 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6834) );
  NAND2_X1 U4618 ( .A1(n3824), .A2(n6834), .ZN(n3743) );
  NAND2_X1 U4619 ( .A1(n3191), .A2(n5911), .ZN(n3741) );
  NAND2_X1 U4620 ( .A1(n4390), .A2(n6834), .ZN(n3740) );
  NAND3_X1 U4621 ( .A1(n3741), .A2(n3188), .A3(n3740), .ZN(n3742) );
  NOR2_X2 U4622 ( .A1(n4428), .A2(n4427), .ZN(n5682) );
  MUX2_X1 U4623 ( .A(n3819), .B(n3188), .S(EBX_REG_5__SCAN_IN), .Z(n3744) );
  OAI21_X1 U4624 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4930), .A(n3744), 
        .ZN(n3745) );
  INV_X1 U4625 ( .A(n3745), .ZN(n5681) );
  NAND2_X1 U4626 ( .A1(n5682), .A2(n5681), .ZN(n5683) );
  INV_X1 U4627 ( .A(EBX_REG_6__SCAN_IN), .ZN(n3746) );
  NAND2_X1 U4628 ( .A1(n3824), .A2(n3746), .ZN(n3750) );
  NAND2_X1 U4629 ( .A1(n3191), .A2(n3850), .ZN(n3748) );
  NAND2_X1 U4630 ( .A1(n4390), .A2(n3746), .ZN(n3747) );
  NAND3_X1 U4631 ( .A1(n3748), .A2(n3188), .A3(n3747), .ZN(n3749) );
  AND2_X1 U4632 ( .A1(n3750), .A2(n3749), .ZN(n4518) );
  OR2_X2 U4633 ( .A1(n5683), .A2(n4518), .ZN(n4528) );
  INV_X1 U4634 ( .A(n4930), .ZN(n3772) );
  NAND2_X1 U4635 ( .A1(n3589), .A2(n3772), .ZN(n3752) );
  MUX2_X1 U4636 ( .A(n3819), .B(n3188), .S(EBX_REG_7__SCAN_IN), .Z(n3751) );
  NAND2_X1 U4637 ( .A1(n3752), .A2(n3751), .ZN(n4529) );
  INV_X1 U4638 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U4639 ( .A1(n3824), .A2(n5650), .ZN(n3756) );
  NAND2_X1 U4640 ( .A1(n3191), .A2(n6931), .ZN(n3754) );
  NAND2_X1 U4641 ( .A1(n4390), .A2(n5650), .ZN(n3753) );
  NAND3_X1 U4642 ( .A1(n3754), .A2(n3188), .A3(n3753), .ZN(n3755) );
  NAND2_X1 U4643 ( .A1(n3756), .A2(n3755), .ZN(n4542) );
  AND2_X2 U4644 ( .A1(n4543), .A2(n4542), .ZN(n5637) );
  INV_X1 U4645 ( .A(n3819), .ZN(n3810) );
  INV_X1 U4646 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U4647 ( .A1(n3810), .A2(n5726), .ZN(n3759) );
  NAND2_X1 U4648 ( .A1(n4390), .A2(n5726), .ZN(n3757) );
  OAI211_X1 U4649 ( .C1(n5181), .C2(n4626), .A(n3757), .B(n3191), .ZN(n3758)
         );
  MUX2_X1 U4650 ( .A(n3819), .B(n3188), .S(EBX_REG_11__SCAN_IN), .Z(n3761) );
  NAND2_X1 U4651 ( .A1(n3605), .A2(n3772), .ZN(n3760) );
  AND2_X1 U4652 ( .A1(n3761), .A2(n3760), .ZN(n4636) );
  INV_X1 U4653 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4624) );
  NAND2_X1 U4654 ( .A1(n3824), .A2(n4624), .ZN(n3766) );
  NAND2_X1 U4655 ( .A1(n3188), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3762) );
  NAND2_X1 U4656 ( .A1(n3191), .A2(n3762), .ZN(n3764) );
  NAND2_X1 U4657 ( .A1(n4390), .A2(n4624), .ZN(n3763) );
  NAND2_X1 U4658 ( .A1(n3764), .A2(n3763), .ZN(n3765) );
  NAND2_X1 U4659 ( .A1(n3766), .A2(n3765), .ZN(n4637) );
  NAND2_X1 U4660 ( .A1(n4636), .A2(n4637), .ZN(n3767) );
  OR2_X2 U4661 ( .A1(n4635), .A2(n3767), .ZN(n4656) );
  OAI21_X1 U4662 ( .B1(n5181), .B2(n4951), .A(n3191), .ZN(n3768) );
  OAI21_X1 U4663 ( .B1(EBX_REG_12__SCAN_IN), .B2(n3734), .A(n3768), .ZN(n3771)
         );
  INV_X1 U4664 ( .A(EBX_REG_12__SCAN_IN), .ZN(n3769) );
  NAND2_X1 U4665 ( .A1(n3824), .A2(n3769), .ZN(n3770) );
  AND2_X1 U4666 ( .A1(n3771), .A2(n3770), .ZN(n4655) );
  NOR2_X2 U4667 ( .A1(n4656), .A2(n4655), .ZN(n5540) );
  MUX2_X1 U4668 ( .A(n3819), .B(n3188), .S(EBX_REG_13__SCAN_IN), .Z(n3774) );
  NAND2_X1 U4669 ( .A1(n3613), .A2(n3772), .ZN(n3773) );
  AND2_X1 U4670 ( .A1(n3774), .A2(n3773), .ZN(n5539) );
  NAND2_X1 U4671 ( .A1(n3188), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3775) );
  NAND2_X1 U4672 ( .A1(n3191), .A2(n3775), .ZN(n3776) );
  OAI21_X1 U4673 ( .B1(EBX_REG_14__SCAN_IN), .B2(n3734), .A(n3776), .ZN(n3777)
         );
  OAI21_X1 U4674 ( .B1(n4925), .B2(EBX_REG_14__SCAN_IN), .A(n3777), .ZN(n4681)
         );
  NAND2_X1 U4675 ( .A1(n5542), .A2(n4681), .ZN(n4680) );
  MUX2_X1 U4676 ( .A(n3819), .B(n3188), .S(EBX_REG_15__SCAN_IN), .Z(n3778) );
  OAI21_X1 U4677 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n4930), .A(n3778), 
        .ZN(n4937) );
  OR2_X2 U4678 ( .A1(n4680), .A2(n4937), .ZN(n4935) );
  INV_X1 U4679 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U4680 ( .A1(n3824), .A2(n5595), .ZN(n3782) );
  NAND2_X1 U4681 ( .A1(n3191), .A2(n4262), .ZN(n3780) );
  NAND2_X1 U4682 ( .A1(n4390), .A2(n5595), .ZN(n3779) );
  NAND3_X1 U4683 ( .A1(n3780), .A2(n3188), .A3(n3779), .ZN(n3781) );
  AND2_X1 U4684 ( .A1(n3782), .A2(n3781), .ZN(n4263) );
  INV_X1 U4685 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6953) );
  NAND2_X1 U4686 ( .A1(n3810), .A2(n6953), .ZN(n3785) );
  NAND2_X1 U4687 ( .A1(n4390), .A2(n6953), .ZN(n3783) );
  OAI211_X1 U4688 ( .C1(n5181), .C2(n5534), .A(n3783), .B(n3191), .ZN(n3784)
         );
  AND2_X1 U4689 ( .A1(n3785), .A2(n3784), .ZN(n5080) );
  INV_X1 U4690 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U4691 ( .A1(n3824), .A2(n5485), .ZN(n3789) );
  INV_X1 U4692 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5418) );
  NAND2_X1 U4693 ( .A1(n3191), .A2(n5418), .ZN(n3787) );
  NAND2_X1 U4694 ( .A1(n4390), .A2(n5485), .ZN(n3786) );
  NAND3_X1 U4695 ( .A1(n3787), .A2(n3188), .A3(n3786), .ZN(n3788) );
  AND2_X1 U4696 ( .A1(n3789), .A2(n3788), .ZN(n5183) );
  OR2_X2 U4697 ( .A1(n5079), .A2(n5183), .ZN(n5169) );
  NAND2_X1 U4698 ( .A1(n4930), .A2(EBX_REG_18__SCAN_IN), .ZN(n3791) );
  NAND2_X1 U4699 ( .A1(n3734), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3790) );
  NAND2_X1 U4700 ( .A1(n3791), .A2(n3790), .ZN(n5182) );
  OR2_X1 U4701 ( .A1(n4930), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3793)
         );
  INV_X1 U4702 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U4703 ( .A1(n4390), .A2(n5177), .ZN(n3792) );
  NAND2_X1 U4704 ( .A1(n3793), .A2(n3792), .ZN(n5172) );
  NAND2_X1 U4705 ( .A1(n5172), .A2(n5182), .ZN(n3795) );
  NAND2_X1 U4706 ( .A1(n5181), .A2(EBX_REG_20__SCAN_IN), .ZN(n3794) );
  OAI211_X1 U4707 ( .C1(n5182), .C2(n5181), .A(n3795), .B(n3794), .ZN(n3796)
         );
  NOR2_X2 U4708 ( .A1(n5169), .A2(n3796), .ZN(n5072) );
  INV_X1 U4709 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5067) );
  NAND2_X1 U4710 ( .A1(n3810), .A2(n5067), .ZN(n3799) );
  NAND2_X1 U4711 ( .A1(n3188), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3797) );
  OAI211_X1 U4712 ( .C1(n3734), .C2(EBX_REG_21__SCAN_IN), .A(n3191), .B(n3797), 
        .ZN(n3798) );
  AND2_X1 U4713 ( .A1(n3799), .A2(n3798), .ZN(n5071) );
  NAND2_X1 U4714 ( .A1(n5072), .A2(n5071), .ZN(n5070) );
  INV_X1 U4715 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6796) );
  NAND2_X1 U4716 ( .A1(n3824), .A2(n6796), .ZN(n3803) );
  NAND2_X1 U4717 ( .A1(n3191), .A2(n5385), .ZN(n3801) );
  NAND2_X1 U4718 ( .A1(n4390), .A2(n6796), .ZN(n3800) );
  NAND3_X1 U4719 ( .A1(n3801), .A2(n3188), .A3(n3800), .ZN(n3802) );
  AND2_X1 U4720 ( .A1(n3803), .A2(n3802), .ZN(n5163) );
  NOR2_X2 U4721 ( .A1(n5070), .A2(n5163), .ZN(n4232) );
  MUX2_X1 U4722 ( .A(n3819), .B(n3188), .S(EBX_REG_23__SCAN_IN), .Z(n3804) );
  OAI21_X1 U4723 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n4930), .A(n3804), 
        .ZN(n4233) );
  NAND2_X1 U4724 ( .A1(n4232), .A2(n3805), .ZN(n5156) );
  INV_X1 U4725 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6924) );
  OAI21_X1 U4726 ( .B1(n5181), .B2(n6924), .A(n3191), .ZN(n3806) );
  OAI21_X1 U4727 ( .B1(EBX_REG_24__SCAN_IN), .B2(n3734), .A(n3806), .ZN(n3809)
         );
  INV_X1 U4728 ( .A(EBX_REG_24__SCAN_IN), .ZN(n3807) );
  NAND2_X1 U4729 ( .A1(n3824), .A2(n3807), .ZN(n3808) );
  AND2_X1 U4730 ( .A1(n3809), .A2(n3808), .ZN(n5155) );
  NOR2_X2 U4731 ( .A1(n5156), .A2(n5155), .ZN(n5357) );
  INV_X1 U4732 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U4733 ( .A1(n3810), .A2(n5488), .ZN(n3813) );
  NAND2_X1 U4734 ( .A1(n3188), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3811) );
  OAI211_X1 U4735 ( .C1(n3734), .C2(EBX_REG_25__SCAN_IN), .A(n3191), .B(n3811), 
        .ZN(n3812) );
  AND2_X1 U4736 ( .A1(n3813), .A2(n3812), .ZN(n5356) );
  NAND2_X1 U4737 ( .A1(n3188), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3814) );
  NAND2_X1 U4738 ( .A1(n3191), .A2(n3814), .ZN(n3817) );
  INV_X1 U4739 ( .A(EBX_REG_26__SCAN_IN), .ZN(n3815) );
  NAND2_X1 U4740 ( .A1(n4390), .A2(n3815), .ZN(n3816) );
  NAND2_X1 U4741 ( .A1(n3817), .A2(n3816), .ZN(n3818) );
  OAI21_X1 U4742 ( .B1(n4925), .B2(EBX_REG_26__SCAN_IN), .A(n3818), .ZN(n5153)
         );
  NAND2_X1 U4743 ( .A1(n5358), .A2(n5153), .ZN(n5057) );
  MUX2_X1 U4744 ( .A(n3819), .B(n3188), .S(EBX_REG_27__SCAN_IN), .Z(n3820) );
  OAI21_X1 U4745 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4930), .A(n3820), 
        .ZN(n5058) );
  OR2_X2 U4746 ( .A1(n5057), .A2(n5058), .ZN(n5060) );
  NAND2_X1 U4747 ( .A1(n3732), .A2(n3821), .ZN(n3822) );
  OAI211_X1 U4748 ( .C1(EBX_REG_28__SCAN_IN), .C2(n3734), .A(n3822), .B(n3188), 
        .ZN(n3826) );
  INV_X1 U4749 ( .A(EBX_REG_28__SCAN_IN), .ZN(n3823) );
  NAND2_X1 U4750 ( .A1(n3824), .A2(n3823), .ZN(n3825) );
  AND2_X1 U4751 ( .A1(n3826), .A2(n3825), .ZN(n5043) );
  NOR2_X4 U4752 ( .A1(n5060), .A2(n5043), .ZN(n5045) );
  OR2_X1 U4753 ( .A1(n4930), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3829)
         );
  INV_X1 U4754 ( .A(EBX_REG_29__SCAN_IN), .ZN(n3827) );
  NAND2_X1 U4755 ( .A1(n4390), .A2(n3827), .ZN(n3828) );
  AND2_X1 U4756 ( .A1(n3829), .A2(n3828), .ZN(n4924) );
  NAND2_X1 U4757 ( .A1(n5045), .A2(n4924), .ZN(n4923) );
  OAI21_X1 U4758 ( .B1(n5045), .B2(n3188), .A(n4923), .ZN(n3831) );
  AND2_X1 U4759 ( .A1(n3734), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3830)
         );
  AOI21_X1 U4760 ( .B1(n4930), .B2(EBX_REG_30__SCAN_IN), .A(n3830), .ZN(n4927)
         );
  OR2_X1 U4761 ( .A1(n4329), .A2(n6615), .ZN(n4607) );
  OR2_X1 U4762 ( .A1(n3833), .A2(n3832), .ZN(n3834) );
  AND2_X1 U4763 ( .A1(n4607), .A2(n3834), .ZN(n3835) );
  OR2_X1 U4764 ( .A1(n4396), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5912) );
  INV_X1 U4765 ( .A(REIP_REG_30__SCAN_IN), .ZN(n3836) );
  NOR2_X1 U4766 ( .A1(n5912), .A2(n3836), .ZN(n5002) );
  NAND2_X1 U4767 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4260) );
  NAND2_X1 U4768 ( .A1(n4286), .A2(n4297), .ZN(n4583) );
  NOR2_X1 U4769 ( .A1(n5932), .A2(n4714), .ZN(n5922) );
  NOR2_X1 U4770 ( .A1(n5911), .A2(n5920), .ZN(n5901) );
  AND2_X1 U4771 ( .A1(n5922), .A2(n5901), .ZN(n5890) );
  NAND3_X1 U4772 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n5890), .ZN(n4566) );
  NOR2_X1 U4773 ( .A1(n6931), .A2(n3589), .ZN(n5867) );
  NAND3_X1 U4774 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n5867), .ZN(n3851) );
  NOR2_X1 U4775 ( .A1(n4566), .A2(n3851), .ZN(n3860) );
  OR2_X1 U4776 ( .A1(n5111), .A2(n3837), .ZN(n4313) );
  NAND2_X1 U4777 ( .A1(n4313), .A2(n4448), .ZN(n3839) );
  OAI21_X1 U4778 ( .B1(n3839), .B2(n4930), .A(n3838), .ZN(n3841) );
  NAND2_X1 U4779 ( .A1(n3338), .A2(n5181), .ZN(n3840) );
  NAND2_X1 U4780 ( .A1(n3841), .A2(n3840), .ZN(n3842) );
  NOR2_X1 U4781 ( .A1(n3843), .A2(n3842), .ZN(n3844) );
  AND2_X1 U4782 ( .A1(n3845), .A2(n3844), .ZN(n4331) );
  OR2_X1 U4783 ( .A1(n3846), .A2(n3188), .ZN(n3847) );
  INV_X1 U4784 ( .A(n3848), .ZN(n3849) );
  NAND2_X1 U4785 ( .A1(n4323), .A2(n3849), .ZN(n4457) );
  INV_X1 U4786 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4723) );
  OAI21_X1 U4787 ( .B1(n4723), .B2(n4714), .A(n5932), .ZN(n5899) );
  NAND2_X1 U4788 ( .A1(n5901), .A2(n5899), .ZN(n5888) );
  OR2_X1 U4789 ( .A1(n5887), .A2(n5888), .ZN(n4512) );
  NOR2_X1 U4790 ( .A1(n3850), .A2(n4512), .ZN(n4564) );
  INV_X1 U4791 ( .A(n4564), .ZN(n4562) );
  NOR2_X1 U4792 ( .A1(n3851), .A2(n4562), .ZN(n3862) );
  INV_X1 U4793 ( .A(n3862), .ZN(n4256) );
  OR2_X1 U4794 ( .A1(n3859), .A2(n4323), .ZN(n3858) );
  NAND2_X1 U4795 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n3860), .ZN(n3852)
         );
  OAI22_X1 U4796 ( .A1(n5897), .A2(n4256), .B1(n3858), .B2(n3852), .ZN(n4704)
         );
  AOI21_X1 U4797 ( .B1(n4339), .B2(n3860), .A(n4704), .ZN(n5548) );
  NAND2_X1 U4798 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4699) );
  NOR2_X1 U4799 ( .A1(n3613), .A2(n4699), .ZN(n4703) );
  INV_X1 U4800 ( .A(n4703), .ZN(n3853) );
  NOR2_X1 U4801 ( .A1(n5548), .A2(n3853), .ZN(n4708) );
  NAND2_X1 U4802 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4708), .ZN(n4940) );
  NOR2_X1 U4803 ( .A1(n4260), .A2(n4940), .ZN(n5535) );
  INV_X1 U4804 ( .A(n3854), .ZN(n3864) );
  AND2_X1 U4805 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U4806 ( .A1(n5355), .A2(n5347), .ZN(n5342) );
  NOR2_X1 U4807 ( .A1(n5342), .A2(n5235), .ZN(n5327) );
  AND3_X1 U4808 ( .A1(n5327), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n3856), 
        .ZN(n3857) );
  AOI211_X1 U4809 ( .C1(n5026), .C2(n5927), .A(n5002), .B(n3857), .ZN(n3877)
         );
  NAND2_X1 U4810 ( .A1(n5897), .A2(n3858), .ZN(n4700) );
  INV_X1 U4811 ( .A(n5868), .ZN(n4513) );
  NAND2_X1 U4812 ( .A1(n3858), .A2(n4702), .ZN(n4567) );
  NAND2_X1 U4813 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4703), .ZN(n4257) );
  NOR2_X1 U4814 ( .A1(n4257), .A2(n4260), .ZN(n3863) );
  INV_X1 U4815 ( .A(n3863), .ZN(n3861) );
  INV_X1 U4816 ( .A(n4567), .ZN(n4511) );
  NAND2_X1 U4817 ( .A1(n5912), .A2(n3859), .ZN(n4337) );
  NAND2_X1 U4818 ( .A1(n4723), .A2(n4700), .ZN(n4341) );
  NAND2_X1 U4819 ( .A1(n4337), .A2(n4341), .ZN(n4385) );
  NAND2_X1 U4820 ( .A1(n5897), .A2(n4385), .ZN(n4563) );
  OAI21_X1 U4821 ( .B1(n4511), .B2(n3860), .A(n4563), .ZN(n4255) );
  AOI21_X1 U4822 ( .B1(n4567), .B2(n3861), .A(n4255), .ZN(n5406) );
  NAND2_X1 U4823 ( .A1(n3863), .A2(n3862), .ZN(n5405) );
  INV_X1 U4824 ( .A(n5408), .ZN(n5386) );
  NAND2_X1 U4825 ( .A1(n5386), .A2(n3864), .ZN(n3865) );
  NOR2_X1 U4826 ( .A1(n5405), .A2(n3865), .ZN(n3866) );
  OR2_X1 U4827 ( .A1(n5868), .A2(n3866), .ZN(n3867) );
  AND2_X1 U4828 ( .A1(n5406), .A2(n3867), .ZN(n5398) );
  INV_X1 U4829 ( .A(n3868), .ZN(n3869) );
  OR2_X1 U4830 ( .A1(n5868), .A2(n3869), .ZN(n3870) );
  AND2_X1 U4831 ( .A1(n5398), .A2(n3870), .ZN(n5380) );
  NOR2_X1 U4832 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n4339), .ZN(n4384)
         );
  NOR2_X1 U4833 ( .A1(n4511), .A2(n4384), .ZN(n5933) );
  INV_X1 U4834 ( .A(n5897), .ZN(n5923) );
  INV_X1 U4835 ( .A(n3871), .ZN(n3872) );
  OAI21_X1 U4836 ( .B1(n5933), .B2(n5923), .A(n3872), .ZN(n3873) );
  NAND2_X1 U4837 ( .A1(n5368), .A2(n5868), .ZN(n3875) );
  NAND2_X1 U4838 ( .A1(n5368), .A2(n5347), .ZN(n3874) );
  AND2_X1 U4839 ( .A1(n3875), .A2(n3874), .ZN(n5344) );
  AOI21_X1 U4840 ( .B1(n5235), .B2(n4513), .A(n5344), .ZN(n4986) );
  NAND2_X1 U4841 ( .A1(n4986), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5326) );
  NAND3_X1 U4842 ( .A1(n5326), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n3875), .ZN(n3876) );
  OAI21_X1 U4843 ( .B1(n5007), .B2(n5906), .A(n3878), .ZN(U2988) );
  NAND2_X1 U4844 ( .A1(n5982), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4070) );
  NAND2_X1 U4845 ( .A1(n6458), .A2(n4052), .ZN(n3881) );
  AND2_X1 U4846 ( .A1(n4448), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3918) );
  INV_X1 U4847 ( .A(EAX_REG_1__SCAN_IN), .ZN(n4301) );
  INV_X1 U4848 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5138) );
  OAI22_X1 U4849 ( .A1(n4861), .A2(n4301), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5138), .ZN(n3879) );
  AOI21_X1 U4850 ( .B1(n3918), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3879), 
        .ZN(n3880) );
  NAND2_X1 U4851 ( .A1(n3881), .A2(n3880), .ZN(n4406) );
  NAND2_X1 U4852 ( .A1(n3882), .A2(n5982), .ZN(n3883) );
  NAND2_X1 U4853 ( .A1(n3883), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4347) );
  INV_X1 U4854 ( .A(n3918), .ZN(n3888) );
  NAND2_X1 U4855 ( .A1(n6799), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3887)
         );
  NAND2_X1 U4856 ( .A1(n4965), .A2(EAX_REG_0__SCAN_IN), .ZN(n3886) );
  OAI211_X1 U4857 ( .C1(n3888), .C2(n3885), .A(n3887), .B(n3886), .ZN(n3889)
         );
  AOI21_X1 U4858 ( .B1(n6244), .B2(n4052), .A(n3889), .ZN(n4346) );
  OR2_X1 U4859 ( .A1(n4347), .A2(n4346), .ZN(n4349) );
  INV_X1 U4860 ( .A(n4346), .ZN(n3890) );
  OR2_X1 U4861 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4798) );
  OR2_X1 U4862 ( .A1(n3890), .A2(n4798), .ZN(n3891) );
  NAND2_X1 U4863 ( .A1(n4349), .A2(n3891), .ZN(n4405) );
  NAND2_X1 U4864 ( .A1(n4406), .A2(n4405), .ZN(n4433) );
  INV_X1 U4865 ( .A(EAX_REG_2__SCAN_IN), .ZN(n3893) );
  NAND2_X1 U4866 ( .A1(n6799), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4797) );
  INV_X1 U4867 ( .A(n4797), .ZN(n4964) );
  INV_X1 U4868 ( .A(n4798), .ZN(n4918) );
  NAND2_X1 U4869 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3899) );
  OAI21_X1 U4870 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3899), .ZN(n5855) );
  AOI22_X1 U4871 ( .A1(n4964), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n4918), 
        .B2(n5855), .ZN(n3892) );
  OAI21_X1 U4872 ( .B1(n4861), .B2(n3893), .A(n3892), .ZN(n3894) );
  AOI21_X1 U4873 ( .B1(n3918), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3894), 
        .ZN(n4434) );
  NAND2_X1 U4874 ( .A1(n4433), .A2(n4434), .ZN(n3896) );
  AND2_X2 U4875 ( .A1(n3897), .A2(n3896), .ZN(n4432) );
  NAND2_X1 U4876 ( .A1(n6217), .A2(n4052), .ZN(n3907) );
  INV_X1 U4877 ( .A(EAX_REG_3__SCAN_IN), .ZN(n3904) );
  INV_X1 U4878 ( .A(n3899), .ZN(n3902) );
  INV_X1 U4879 ( .A(n3920), .ZN(n3901) );
  OAI21_X1 U4880 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3902), .A(n3901), 
        .ZN(n5109) );
  AOI22_X1 U4881 ( .A1(n4918), .A2(n5109), .B1(n4964), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3903) );
  OAI21_X1 U4882 ( .B1(n4861), .B2(n3904), .A(n3903), .ZN(n3905) );
  AOI21_X1 U4883 ( .B1(n3918), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3905), 
        .ZN(n3906) );
  NAND2_X1 U4884 ( .A1(n3907), .A2(n3906), .ZN(n4421) );
  AND2_X2 U4885 ( .A1(n4432), .A2(n4421), .ZN(n4500) );
  INV_X1 U4886 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4505) );
  INV_X1 U4887 ( .A(n3919), .ZN(n3909) );
  INV_X1 U4888 ( .A(n3926), .ZN(n3908) );
  OAI21_X1 U4889 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3909), .A(n3908), 
        .ZN(n5837) );
  AOI22_X1 U4890 ( .A1(n4918), .A2(n5837), .B1(n4964), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3910) );
  OAI21_X1 U4891 ( .B1(n4861), .B2(n4505), .A(n3910), .ZN(n3911) );
  INV_X1 U4892 ( .A(n3911), .ZN(n3912) );
  NAND2_X1 U4893 ( .A1(n3914), .A2(n4052), .ZN(n3924) );
  INV_X1 U4894 ( .A(EAX_REG_4__SCAN_IN), .ZN(n3916) );
  INV_X1 U4895 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3915) );
  OAI22_X1 U4896 ( .A1(n4861), .A2(n3916), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3915), .ZN(n3917) );
  AOI21_X1 U4897 ( .B1(n3918), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n3917), 
        .ZN(n3922) );
  OAI21_X1 U4898 ( .B1(n3920), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3919), 
        .ZN(n5846) );
  INV_X1 U4899 ( .A(n5846), .ZN(n3921) );
  MUX2_X1 U4900 ( .A(n3922), .B(n3921), .S(n4918), .Z(n3923) );
  INV_X1 U4901 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3929) );
  NAND2_X1 U4902 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n3926), .ZN(n3933)
         );
  OAI21_X1 U4903 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n3926), .A(n3933), 
        .ZN(n5828) );
  NAND2_X1 U4904 ( .A1(n5828), .A2(n4918), .ZN(n3928) );
  NAND2_X1 U4905 ( .A1(n4965), .A2(EAX_REG_6__SCAN_IN), .ZN(n3927) );
  OAI211_X1 U4906 ( .C1(n4797), .C2(n3929), .A(n3928), .B(n3927), .ZN(n3930)
         );
  NOR2_X2 U4907 ( .A1(n4521), .A2(n4522), .ZN(n4527) );
  OAI21_X1 U4908 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n3934), .A(n3954), 
        .ZN(n5822) );
  INV_X1 U4909 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3936) );
  INV_X1 U4910 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3935) );
  OAI22_X1 U4911 ( .A1(n4861), .A2(n3936), .B1(n4797), .B2(n3935), .ZN(n3937)
         );
  AOI21_X1 U4912 ( .B1(n5822), .B2(n4918), .A(n3937), .ZN(n3938) );
  AOI22_X1 U4913 ( .A1(n3187), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4874), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4914 ( .A1(n3420), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4905), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4915 ( .A1(n4811), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4916 ( .A1(n4869), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3940) );
  NAND4_X1 U4917 ( .A1(n3943), .A2(n3942), .A3(n3941), .A4(n3940), .ZN(n3949)
         );
  AOI22_X1 U4918 ( .A1(n4894), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4868), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4919 ( .A1(n4898), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4920 ( .A1(n3405), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4921 ( .A1(n4893), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3944) );
  NAND4_X1 U4922 ( .A1(n3947), .A2(n3946), .A3(n3945), .A4(n3944), .ZN(n3948)
         );
  NOR2_X1 U4923 ( .A1(n3949), .A2(n3948), .ZN(n3953) );
  INV_X1 U4924 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3950) );
  XNOR2_X1 U4925 ( .A(n3954), .B(n3950), .ZN(n5652) );
  NAND2_X1 U4926 ( .A1(n5652), .A2(n4918), .ZN(n3952) );
  AOI22_X1 U4927 ( .A1(n4965), .A2(EAX_REG_8__SCAN_IN), .B1(n4964), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3951) );
  OAI211_X1 U4928 ( .C1(n3953), .C2(n4070), .A(n3952), .B(n3951), .ZN(n4538)
         );
  NAND2_X1 U4929 ( .A1(n4525), .A2(n4538), .ZN(n4539) );
  XOR2_X1 U4930 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3972), .Z(n5644) );
  INV_X1 U4931 ( .A(n5644), .ZN(n3969) );
  AOI22_X1 U4932 ( .A1(n4894), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4898), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4933 ( .A1(n3367), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4905), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4934 ( .A1(n3187), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4935 ( .A1(n4869), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3955) );
  NAND4_X1 U4936 ( .A1(n3958), .A2(n3957), .A3(n3956), .A4(n3955), .ZN(n3964)
         );
  AOI22_X1 U4937 ( .A1(n4893), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4938 ( .A1(n4868), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4939 ( .A1(n4904), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4940 ( .A1(n3420), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3959) );
  NAND4_X1 U4941 ( .A1(n3962), .A2(n3961), .A3(n3960), .A4(n3959), .ZN(n3963)
         );
  NOR2_X1 U4942 ( .A1(n3964), .A2(n3963), .ZN(n3967) );
  NAND2_X1 U4943 ( .A1(n4965), .A2(EAX_REG_9__SCAN_IN), .ZN(n3966) );
  NAND2_X1 U4944 ( .A1(n4964), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3965)
         );
  OAI211_X1 U4945 ( .C1(n4070), .C2(n3967), .A(n3966), .B(n3965), .ZN(n3968)
         );
  AOI21_X1 U4946 ( .B1(n3969), .B2(n4918), .A(n3968), .ZN(n4551) );
  INV_X1 U4947 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3973) );
  NAND2_X1 U4948 ( .A1(n3991), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3974)
         );
  INV_X1 U4949 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6845) );
  NAND2_X1 U4950 ( .A1(n3974), .A2(n6845), .ZN(n3976) );
  INV_X1 U4951 ( .A(n4023), .ZN(n3975) );
  NAND2_X1 U4952 ( .A1(n3976), .A2(n3975), .ZN(n4959) );
  AOI22_X1 U4953 ( .A1(n4898), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4868), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4954 ( .A1(n4894), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4874), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4955 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3187), .B1(n3405), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4956 ( .A1(n4893), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3977) );
  NAND4_X1 U4957 ( .A1(n3980), .A2(n3979), .A3(n3978), .A4(n3977), .ZN(n3986)
         );
  AOI22_X1 U4958 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n3367), .B1(n4905), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4959 ( .A1(n4895), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4960 ( .A1(n3420), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4961 ( .A1(n4869), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3981) );
  NAND4_X1 U4962 ( .A1(n3984), .A2(n3983), .A3(n3982), .A4(n3981), .ZN(n3985)
         );
  NOR2_X1 U4963 ( .A1(n3986), .A2(n3985), .ZN(n3989) );
  NAND2_X1 U4964 ( .A1(n4965), .A2(EAX_REG_12__SCAN_IN), .ZN(n3988) );
  NAND2_X1 U4965 ( .A1(n4964), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3987)
         );
  OAI211_X1 U4966 ( .C1(n4070), .C2(n3989), .A(n3988), .B(n3987), .ZN(n3990)
         );
  AOI21_X1 U4967 ( .B1(n4959), .B2(n4918), .A(n3990), .ZN(n4650) );
  INV_X1 U4968 ( .A(n4650), .ZN(n4005) );
  XOR2_X1 U4969 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3991), .Z(n5809) );
  AOI22_X1 U4970 ( .A1(n3420), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4971 ( .A1(n4898), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4868), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4972 ( .A1(n3187), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U4973 ( .A1(n3404), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3992) );
  NAND4_X1 U4974 ( .A1(n3995), .A2(n3994), .A3(n3993), .A4(n3992), .ZN(n4001)
         );
  AOI22_X1 U4975 ( .A1(n4894), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4874), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4976 ( .A1(n4893), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4977 ( .A1(n4869), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4978 ( .A1(n4905), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3996) );
  NAND4_X1 U4979 ( .A1(n3999), .A2(n3998), .A3(n3997), .A4(n3996), .ZN(n4000)
         );
  OR2_X1 U4980 ( .A1(n4001), .A2(n4000), .ZN(n4002) );
  AOI22_X1 U4981 ( .A1(n4052), .A2(n4002), .B1(n4964), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4004) );
  NAND2_X1 U4982 ( .A1(n4965), .A2(EAX_REG_11__SCAN_IN), .ZN(n4003) );
  OAI211_X1 U4983 ( .C1(n5809), .C2(n4798), .A(n4004), .B(n4003), .ZN(n4632)
         );
  NAND2_X1 U4984 ( .A1(n4005), .A2(n4632), .ZN(n4021) );
  XNOR2_X1 U4985 ( .A(n4006), .B(n3973), .ZN(n5099) );
  AOI22_X1 U4986 ( .A1(n4905), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4874), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4987 ( .A1(n4894), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4898), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4988 ( .A1(n4868), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4989 ( .A1(n4811), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4007) );
  NAND4_X1 U4990 ( .A1(n4010), .A2(n4009), .A3(n4008), .A4(n4007), .ZN(n4016)
         );
  AOI22_X1 U4991 ( .A1(n4893), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4869), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U4992 ( .A1(n3405), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4993 ( .A1(n3420), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4994 ( .A1(n3187), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4011) );
  NAND4_X1 U4995 ( .A1(n4014), .A2(n4013), .A3(n4012), .A4(n4011), .ZN(n4015)
         );
  NOR2_X1 U4996 ( .A1(n4016), .A2(n4015), .ZN(n4019) );
  NAND2_X1 U4997 ( .A1(n4965), .A2(EAX_REG_10__SCAN_IN), .ZN(n4018) );
  NAND2_X1 U4998 ( .A1(n4964), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4017)
         );
  OAI211_X1 U4999 ( .C1(n4070), .C2(n4019), .A(n4018), .B(n4017), .ZN(n4020)
         );
  AOI21_X1 U5000 ( .B1(n5099), .B2(n4918), .A(n4020), .ZN(n4620) );
  NAND2_X1 U5001 ( .A1(n4022), .A2(n3193), .ZN(n4027) );
  INV_X1 U5002 ( .A(EAX_REG_13__SCAN_IN), .ZN(n4674) );
  OAI21_X1 U5003 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n4023), .A(n4056), 
        .ZN(n5635) );
  AOI22_X1 U5004 ( .A1(n4918), .A2(n5635), .B1(n4964), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4024) );
  OAI21_X1 U5005 ( .B1(n4861), .B2(n4674), .A(n4024), .ZN(n4025) );
  INV_X1 U5006 ( .A(n4025), .ZN(n4026) );
  NAND2_X1 U5007 ( .A1(n4027), .A2(n4026), .ZN(n4028) );
  AND2_X2 U5008 ( .A1(n4028), .A2(n4040), .ZN(n4668) );
  AOI22_X1 U5009 ( .A1(n4894), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U5010 ( .A1(n4868), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U5011 ( .A1(n3187), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U5012 ( .A1(n4893), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4029) );
  NAND4_X1 U5013 ( .A1(n4032), .A2(n4031), .A3(n4030), .A4(n4029), .ZN(n4038)
         );
  AOI22_X1 U5014 ( .A1(n3420), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4905), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U5015 ( .A1(n3399), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U5016 ( .A1(n4904), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U5017 ( .A1(n4869), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4033) );
  NAND4_X1 U5018 ( .A1(n4036), .A2(n4035), .A3(n4034), .A4(n4033), .ZN(n4037)
         );
  OR2_X1 U5019 ( .A1(n4038), .A2(n4037), .ZN(n4039) );
  AND2_X1 U5020 ( .A1(n4052), .A2(n4039), .ZN(n4669) );
  INV_X1 U5021 ( .A(EAX_REG_14__SCAN_IN), .ZN(n4684) );
  AOI22_X1 U5022 ( .A1(n4893), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4905), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U5023 ( .A1(n4868), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5024 ( .A1(n3418), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U5025 ( .A1(n4894), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4041) );
  NAND4_X1 U5026 ( .A1(n4044), .A2(n4043), .A3(n4042), .A4(n4041), .ZN(n4050)
         );
  AOI22_X1 U5027 ( .A1(n4869), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3419), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U5028 ( .A1(n4898), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U5029 ( .A1(n4904), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U5030 ( .A1(n3187), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4045) );
  NAND4_X1 U5031 ( .A1(n4048), .A2(n4047), .A3(n4046), .A4(n4045), .ZN(n4049)
         );
  OR2_X1 U5032 ( .A1(n4050), .A2(n4049), .ZN(n4051) );
  NAND2_X1 U5033 ( .A1(n4052), .A2(n4051), .ZN(n4055) );
  XNOR2_X1 U5034 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4056), .ZN(n5617)
         );
  INV_X1 U5035 ( .A(n5617), .ZN(n4053) );
  AOI22_X1 U5036 ( .A1(n4964), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n4918), 
        .B2(n4053), .ZN(n4054) );
  OAI211_X1 U5037 ( .C1(n4684), .C2(n4861), .A(n4055), .B(n4054), .ZN(n4678)
         );
  INV_X1 U5038 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5614) );
  XNOR2_X1 U5039 ( .A(n4072), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5602)
         );
  AOI22_X1 U5040 ( .A1(n4893), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5041 ( .A1(n4869), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3187), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U5042 ( .A1(n3428), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U5043 ( .A1(n4868), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4057) );
  NAND4_X1 U5044 ( .A1(n4060), .A2(n4059), .A3(n4058), .A4(n4057), .ZN(n4066)
         );
  AOI22_X1 U5045 ( .A1(n4811), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4904), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5046 ( .A1(n3419), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U5047 ( .A1(n4894), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U5048 ( .A1(n4905), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4061) );
  NAND4_X1 U5049 ( .A1(n4064), .A2(n4063), .A3(n4062), .A4(n4061), .ZN(n4065)
         );
  NOR2_X1 U5050 ( .A1(n4066), .A2(n4065), .ZN(n4069) );
  NAND2_X1 U5051 ( .A1(n4965), .A2(EAX_REG_15__SCAN_IN), .ZN(n4068) );
  NAND2_X1 U5052 ( .A1(n4964), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4067)
         );
  OAI211_X1 U5053 ( .C1(n4070), .C2(n4069), .A(n4068), .B(n4067), .ZN(n4071)
         );
  AOI21_X1 U5054 ( .B1(n5602), .B2(n4918), .A(n4071), .ZN(n4944) );
  XNOR2_X1 U5055 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n4088), .ZN(n5597)
         );
  INV_X1 U5056 ( .A(n5597), .ZN(n4086) );
  NAND2_X1 U5057 ( .A1(n4580), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4915) );
  AOI22_X1 U5058 ( .A1(n3419), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4905), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5059 ( .A1(n4893), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4075) );
  AOI22_X1 U5060 ( .A1(n4898), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4074) );
  AOI22_X1 U5061 ( .A1(n4904), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4073) );
  NAND4_X1 U5062 ( .A1(n4076), .A2(n4075), .A3(n4074), .A4(n4073), .ZN(n4082)
         );
  AOI22_X1 U5063 ( .A1(n4868), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3187), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U5064 ( .A1(n4811), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4079) );
  AOI22_X1 U5065 ( .A1(n4869), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U5066 ( .A1(n4894), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4077) );
  NAND4_X1 U5067 ( .A1(n4080), .A2(n4079), .A3(n4078), .A4(n4077), .ZN(n4081)
         );
  NOR2_X1 U5068 ( .A1(n4082), .A2(n4081), .ZN(n4084) );
  AOI22_X1 U5069 ( .A1(n4965), .A2(EAX_REG_16__SCAN_IN), .B1(n4964), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4083) );
  OAI21_X1 U5070 ( .B1(n4915), .B2(n4084), .A(n4083), .ZN(n4085) );
  AOI21_X1 U5071 ( .B1(n4086), .B2(n4918), .A(n4085), .ZN(n5197) );
  NOR2_X4 U5072 ( .A1(n5196), .A2(n5197), .ZN(n5076) );
  INV_X1 U5073 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4087) );
  XNOR2_X1 U5074 ( .A(n4102), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5313)
         );
  AOI22_X1 U5075 ( .A1(n4869), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3187), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4092) );
  AOI22_X1 U5076 ( .A1(n4893), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U5077 ( .A1(n4904), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U5078 ( .A1(n3419), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4089) );
  NAND4_X1 U5079 ( .A1(n4092), .A2(n4091), .A3(n4090), .A4(n4089), .ZN(n4098)
         );
  AOI22_X1 U5080 ( .A1(n4894), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4868), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4096) );
  AOI22_X1 U5081 ( .A1(n4905), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U5082 ( .A1(n3399), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U5083 ( .A1(n3404), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4093) );
  NAND4_X1 U5084 ( .A1(n4096), .A2(n4095), .A3(n4094), .A4(n4093), .ZN(n4097)
         );
  NOR2_X1 U5085 ( .A1(n4098), .A2(n4097), .ZN(n4100) );
  AOI22_X1 U5086 ( .A1(n4965), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6799), .ZN(n4099) );
  OAI21_X1 U5087 ( .B1(n4915), .B2(n4100), .A(n4099), .ZN(n4101) );
  MUX2_X1 U5088 ( .A(n5313), .B(n4101), .S(n4798), .Z(n5077) );
  OAI21_X1 U5089 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n4103), .A(n4134), 
        .ZN(n5585) );
  INV_X1 U5090 ( .A(n5585), .ZN(n4119) );
  INV_X1 U5091 ( .A(n4915), .ZN(n4844) );
  AOI22_X1 U5092 ( .A1(n4893), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U5093 ( .A1(n4894), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5094 ( .A1(n3187), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4904), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5095 ( .A1(n3420), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4104) );
  NAND4_X1 U5096 ( .A1(n4107), .A2(n4106), .A3(n4105), .A4(n4104), .ZN(n4113)
         );
  AOI22_X1 U5097 ( .A1(n4905), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U5098 ( .A1(n4868), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U5099 ( .A1(n3405), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5100 ( .A1(n4869), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4108) );
  NAND4_X1 U5101 ( .A1(n4111), .A2(n4110), .A3(n4109), .A4(n4108), .ZN(n4112)
         );
  OR2_X1 U5102 ( .A1(n4113), .A2(n4112), .ZN(n4117) );
  INV_X1 U5103 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4115) );
  INV_X1 U5104 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4114) );
  OAI22_X1 U5105 ( .A1(n4861), .A2(n4115), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4114), .ZN(n4116) );
  AOI21_X1 U5106 ( .B1(n4844), .B2(n4117), .A(n4116), .ZN(n4118) );
  MUX2_X1 U5107 ( .A(n4119), .B(n4118), .S(n4798), .Z(n5189) );
  XNOR2_X1 U5108 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n4134), .ZN(n5482)
         );
  AOI22_X1 U5109 ( .A1(n3420), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4868), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5110 ( .A1(n4894), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U5111 ( .A1(n3399), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4904), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U5112 ( .A1(n4905), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4120) );
  NAND4_X1 U5113 ( .A1(n4123), .A2(n4122), .A3(n4121), .A4(n4120), .ZN(n4129)
         );
  AOI22_X1 U5114 ( .A1(n4869), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U5115 ( .A1(n4893), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5116 ( .A1(n3404), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5117 ( .A1(n3187), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4124) );
  NAND4_X1 U5118 ( .A1(n4127), .A2(n4126), .A3(n4125), .A4(n4124), .ZN(n4128)
         );
  OR2_X1 U5119 ( .A1(n4129), .A2(n4128), .ZN(n4132) );
  INV_X1 U5120 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4130) );
  INV_X1 U5121 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5296) );
  OAI22_X1 U5122 ( .A1(n4861), .A2(n4130), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5296), .ZN(n4131) );
  AOI21_X1 U5123 ( .B1(n4844), .B2(n4132), .A(n4131), .ZN(n4133) );
  MUX2_X1 U5124 ( .A(n5482), .B(n4133), .S(n4798), .Z(n5178) );
  INV_X1 U5125 ( .A(n4137), .ZN(n4136) );
  NAND2_X1 U5126 ( .A1(n4136), .A2(n5457), .ZN(n4138) );
  AND2_X1 U5127 ( .A1(n4138), .A2(n4211), .ZN(n5461) );
  AOI22_X1 U5128 ( .A1(n4898), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4868), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U5129 ( .A1(n4893), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4141) );
  AOI22_X1 U5130 ( .A1(n4904), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U5131 ( .A1(n3420), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4139) );
  NAND4_X1 U5132 ( .A1(n4142), .A2(n4141), .A3(n4140), .A4(n4139), .ZN(n4148)
         );
  AOI22_X1 U5133 ( .A1(n4811), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4905), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4146) );
  AOI22_X1 U5134 ( .A1(n4894), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4145) );
  AOI22_X1 U5135 ( .A1(n4869), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U5136 ( .A1(n3187), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4143) );
  NAND4_X1 U5137 ( .A1(n4146), .A2(n4145), .A3(n4144), .A4(n4143), .ZN(n4147)
         );
  OR2_X1 U5138 ( .A1(n4148), .A2(n4147), .ZN(n4151) );
  INV_X1 U5139 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4149) );
  OAI22_X1 U5140 ( .A1(n4861), .A2(n4149), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5457), .ZN(n4150) );
  AOI21_X1 U5141 ( .B1(n4844), .B2(n4151), .A(n4150), .ZN(n4152) );
  MUX2_X1 U5142 ( .A(n5461), .B(n4152), .S(n4798), .Z(n4755) );
  INV_X1 U5143 ( .A(n4755), .ZN(n4187) );
  AOI22_X1 U5144 ( .A1(n4868), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4156) );
  AOI22_X1 U5145 ( .A1(n3420), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U5146 ( .A1(n4898), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5147 ( .A1(n4893), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4153) );
  NAND4_X1 U5148 ( .A1(n4156), .A2(n4155), .A3(n4154), .A4(n4153), .ZN(n4162)
         );
  AOI22_X1 U5149 ( .A1(n4869), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3187), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4160) );
  AOI22_X1 U5150 ( .A1(n4904), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U5151 ( .A1(n4905), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4158) );
  AOI22_X1 U5152 ( .A1(n4894), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4157) );
  NAND4_X1 U5153 ( .A1(n4160), .A2(n4159), .A3(n4158), .A4(n4157), .ZN(n4161)
         );
  NOR2_X1 U5154 ( .A1(n4162), .A2(n4161), .ZN(n4165) );
  INV_X1 U5155 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5288) );
  AOI21_X1 U5156 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5288), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4163) );
  AOI21_X1 U5157 ( .B1(n4965), .B2(EAX_REG_21__SCAN_IN), .A(n4163), .ZN(n4164)
         );
  OAI21_X1 U5158 ( .B1(n4915), .B2(n4165), .A(n4164), .ZN(n4167) );
  XNOR2_X1 U5159 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n4184), .ZN(n5290)
         );
  NAND2_X1 U5160 ( .A1(n4918), .A2(n5290), .ZN(n4166) );
  AND2_X1 U5161 ( .A1(n4167), .A2(n4166), .ZN(n5066) );
  AOI22_X1 U5162 ( .A1(n4894), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4171) );
  AOI22_X1 U5163 ( .A1(n4868), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U5164 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4898), .B1(n4897), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U5165 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3187), .B1(n3404), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4168) );
  NAND4_X1 U5166 ( .A1(n4171), .A2(n4170), .A3(n4169), .A4(n4168), .ZN(n4177)
         );
  AOI22_X1 U5167 ( .A1(n4893), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3420), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U5168 ( .A1(n4904), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U5169 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4869), .B1(n3405), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4173) );
  AOI22_X1 U5170 ( .A1(n4905), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4172) );
  NAND4_X1 U5171 ( .A1(n4175), .A2(n4174), .A3(n4173), .A4(n4172), .ZN(n4176)
         );
  NOR2_X1 U5172 ( .A1(n4177), .A2(n4176), .ZN(n4182) );
  INV_X1 U5173 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4179) );
  INV_X1 U5174 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4178) );
  OAI22_X1 U5175 ( .A1(n4861), .A2(n4179), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4178), .ZN(n4180) );
  INV_X1 U5176 ( .A(n4180), .ZN(n4181) );
  OAI21_X1 U5177 ( .B1(n4915), .B2(n4182), .A(n4181), .ZN(n4186) );
  OR2_X1 U5178 ( .A1(n4183), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4185)
         );
  NAND2_X1 U5179 ( .A1(n4185), .A2(n4184), .ZN(n5509) );
  MUX2_X1 U5180 ( .A(n4186), .B(n5509), .S(n4918), .Z(n5174) );
  AND2_X1 U5181 ( .A1(n5066), .A2(n5174), .ZN(n4754) );
  AND2_X1 U5182 ( .A1(n4187), .A2(n4754), .ZN(n4216) );
  NAND2_X1 U5183 ( .A1(n5179), .A2(n4216), .ZN(n4758) );
  AOI22_X1 U5184 ( .A1(n4765), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3420), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4191) );
  AOI22_X1 U5185 ( .A1(n4894), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4190) );
  AOI22_X1 U5186 ( .A1(n4896), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U5187 ( .A1(n4898), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4188) );
  NAND4_X1 U5188 ( .A1(n4191), .A2(n4190), .A3(n4189), .A4(n4188), .ZN(n4197)
         );
  AOI22_X1 U5189 ( .A1(n3187), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4195) );
  AOI22_X1 U5190 ( .A1(n4869), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4194) );
  AOI22_X1 U5191 ( .A1(n4904), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4193) );
  AOI22_X1 U5192 ( .A1(n4905), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4192) );
  NAND4_X1 U5193 ( .A1(n4195), .A2(n4194), .A3(n4193), .A4(n4192), .ZN(n4196)
         );
  OR2_X1 U5194 ( .A1(n4197), .A2(n4196), .ZN(n4777) );
  AOI22_X1 U5195 ( .A1(n4765), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3420), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4201) );
  AOI22_X1 U5196 ( .A1(n4894), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4200) );
  AOI22_X1 U5197 ( .A1(n4896), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4199) );
  AOI22_X1 U5198 ( .A1(n4898), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4198) );
  NAND4_X1 U5199 ( .A1(n4201), .A2(n4200), .A3(n4199), .A4(n4198), .ZN(n4207)
         );
  AOI22_X1 U5200 ( .A1(n3187), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4205) );
  AOI22_X1 U5201 ( .A1(n4869), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4204) );
  AOI22_X1 U5202 ( .A1(n4904), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4203) );
  AOI22_X1 U5203 ( .A1(n4905), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4202) );
  NAND4_X1 U5204 ( .A1(n4205), .A2(n4204), .A3(n4203), .A4(n4202), .ZN(n4206)
         );
  OR2_X1 U5205 ( .A1(n4207), .A2(n4206), .ZN(n4776) );
  XNOR2_X1 U5206 ( .A(n4777), .B(n4776), .ZN(n4210) );
  NAND2_X1 U5207 ( .A1(n4965), .A2(EAX_REG_23__SCAN_IN), .ZN(n4209) );
  INV_X1 U5208 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6411) );
  OAI21_X1 U5209 ( .B1(n6411), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n6799), 
        .ZN(n4208) );
  OAI211_X1 U5210 ( .C1(n4915), .C2(n4210), .A(n4209), .B(n4208), .ZN(n4214)
         );
  INV_X1 U5211 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6970) );
  AND2_X1 U5212 ( .A1(n4211), .A2(n6970), .ZN(n4212) );
  NOR2_X1 U5213 ( .A1(n4796), .A2(n4212), .ZN(n4751) );
  NAND2_X1 U5214 ( .A1(n4751), .A2(n4918), .ZN(n4213) );
  NAND2_X1 U5215 ( .A1(n4214), .A2(n4213), .ZN(n4215) );
  INV_X1 U5216 ( .A(n4215), .ZN(n4217) );
  NAND2_X1 U5217 ( .A1(n4217), .A2(n4216), .ZN(n4218) );
  NAND2_X1 U5218 ( .A1(n4288), .A2(n4286), .ZN(n4278) );
  INV_X1 U5219 ( .A(n6515), .ZN(n5556) );
  OR2_X1 U5220 ( .A1(n4278), .A2(n5556), .ZN(n4274) );
  NAND2_X1 U5221 ( .A1(n4299), .A2(n4274), .ZN(n6610) );
  INV_X1 U5222 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6600) );
  NAND2_X1 U5223 ( .A1(n4724), .A2(n6799), .ZN(n6521) );
  NOR3_X1 U5224 ( .A1(n6517), .A2(n6600), .A3(n6521), .ZN(n4613) );
  AND2_X1 U5225 ( .A1(n6517), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4401) );
  NAND2_X1 U5226 ( .A1(n4401), .A2(n4918), .ZN(n6519) );
  NAND2_X1 U5227 ( .A1(n6519), .A2(n5912), .ZN(n4221) );
  OR2_X1 U5228 ( .A1(n4613), .A2(n4221), .ZN(n4222) );
  NAND2_X1 U5229 ( .A1(n4796), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4791)
         );
  INV_X1 U5230 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5269) );
  INV_X1 U5231 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4824) );
  INV_X1 U5232 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4885) );
  INV_X1 U5233 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5018) );
  INV_X1 U5234 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6576) );
  INV_X1 U5235 ( .A(n5112), .ZN(n4227) );
  NOR2_X1 U5236 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4239) );
  OAI211_X1 U5237 ( .C1(n4297), .C2(n4305), .A(n4239), .B(n3190), .ZN(n4225)
         );
  INV_X1 U5238 ( .A(n4225), .ZN(n4226) );
  INV_X1 U5239 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6570) );
  INV_X1 U5240 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6566) );
  INV_X1 U5241 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6563) );
  INV_X1 U5242 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6906) );
  INV_X1 U5243 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6601) );
  NAND2_X1 U5244 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n4228) );
  NOR2_X1 U5245 ( .A1(n6601), .A2(n4228), .ZN(n5117) );
  INV_X1 U5246 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6557) );
  INV_X1 U5247 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U5248 ( .A1(REIP_REG_5__SCAN_IN), .A2(REIP_REG_4__SCAN_IN), .ZN(
        n5663) );
  NOR3_X1 U5249 ( .A1(n6557), .A2(n6554), .A3(n5663), .ZN(n5648) );
  NAND3_X1 U5250 ( .A1(REIP_REG_8__SCAN_IN), .A2(n5117), .A3(n5648), .ZN(n5100) );
  NAND2_X1 U5251 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5104) );
  NOR3_X1 U5252 ( .A1(n6906), .A2(n5100), .A3(n5104), .ZN(n4663) );
  NAND2_X1 U5253 ( .A1(REIP_REG_12__SCAN_IN), .A2(n4663), .ZN(n5623) );
  NOR2_X1 U5254 ( .A1(n6563), .A2(n5623), .ZN(n5611) );
  NAND2_X1 U5255 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5611), .ZN(n5589) );
  NOR2_X1 U5256 ( .A1(n6566), .A2(n5589), .ZN(n5592) );
  NAND2_X1 U5257 ( .A1(REIP_REG_16__SCAN_IN), .A2(n5592), .ZN(n5083) );
  NOR2_X1 U5258 ( .A1(n6570), .A2(n5083), .ZN(n4229) );
  NAND2_X1 U5259 ( .A1(n5612), .A2(n4229), .ZN(n5581) );
  INV_X1 U5260 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6575) );
  INV_X1 U5261 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6571) );
  INV_X1 U5262 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6572) );
  NOR2_X1 U5263 ( .A1(n6576), .A2(n5455), .ZN(n5460) );
  AOI21_X1 U5264 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5460), .A(
        REIP_REG_23__SCAN_IN), .ZN(n4231) );
  NAND3_X1 U5265 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n4230) );
  NAND2_X1 U5266 ( .A1(n4229), .A2(n5591), .ZN(n5474) );
  NOR2_X1 U5267 ( .A1(n4230), .A2(n5474), .ZN(n5456) );
  NAND4_X1 U5268 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5456), .ZN(n4969) );
  NAND2_X1 U5269 ( .A1(n5667), .A2(n5591), .ZN(n5473) );
  NAND2_X1 U5270 ( .A1(n4969), .A2(n5473), .ZN(n5447) );
  OAI22_X1 U5271 ( .A1(n5223), .A2(n5479), .B1(n4231), .B2(n5447), .ZN(n4248)
         );
  NAND2_X1 U5272 ( .A1(n5165), .A2(n4233), .ZN(n4234) );
  AND2_X1 U5273 ( .A1(n5156), .A2(n4234), .ZN(n5376) );
  INV_X1 U5274 ( .A(EBX_REG_31__SCAN_IN), .ZN(n4235) );
  NOR2_X1 U5275 ( .A1(n5112), .A2(n4235), .ZN(n4972) );
  NOR2_X1 U5276 ( .A1(n3734), .A2(n4239), .ZN(n4236) );
  NOR2_X1 U5277 ( .A1(n4992), .A2(n4724), .ZN(n4237) );
  INV_X1 U5278 ( .A(n4239), .ZN(n4238) );
  NOR2_X1 U5279 ( .A1(n6533), .A2(n4238), .ZN(n4605) );
  NOR2_X1 U5280 ( .A1(n6615), .A2(n4605), .ZN(n4971) );
  NOR2_X1 U5281 ( .A1(n4239), .A2(EBX_REG_31__SCAN_IN), .ZN(n4240) );
  AND2_X1 U5282 ( .A1(n4307), .A2(n4240), .ZN(n4241) );
  NOR2_X1 U5283 ( .A1(n4971), .A2(n4241), .ZN(n4242) );
  NOR2_X2 U5284 ( .A1(n5112), .A2(n4242), .ZN(n5699) );
  AOI22_X1 U5285 ( .A1(n4751), .A2(n5654), .B1(EBX_REG_23__SCAN_IN), .B2(n5699), .ZN(n4243) );
  INV_X1 U5286 ( .A(n4249), .ZN(n4250) );
  AOI21_X2 U5287 ( .B1(n4251), .B2(n4250), .A(n3196), .ZN(n4933) );
  AND2_X1 U5288 ( .A1(n5303), .A2(n4252), .ZN(n4254) );
  NOR2_X1 U5289 ( .A1(n5806), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5308)
         );
  INV_X1 U5290 ( .A(n5308), .ZN(n5305) );
  OAI21_X1 U5291 ( .B1(n3620), .B2(n4262), .A(n5305), .ZN(n4253) );
  XNOR2_X1 U5292 ( .A(n4254), .B(n4253), .ZN(n5322) );
  NOR2_X1 U5293 ( .A1(n5322), .A2(n5906), .ZN(n4269) );
  AOI21_X1 U5294 ( .B1(n4256), .B2(n5923), .A(n4255), .ZN(n5860) );
  INV_X1 U5295 ( .A(n4257), .ZN(n4258) );
  OR2_X1 U5296 ( .A1(n5868), .A2(n4258), .ZN(n4259) );
  AND2_X1 U5297 ( .A1(n5860), .A2(n4259), .ZN(n4939) );
  NOR2_X1 U5298 ( .A1(n4939), .A2(n4262), .ZN(n4268) );
  INV_X1 U5299 ( .A(n4260), .ZN(n4261) );
  AOI211_X1 U5300 ( .C1(n4262), .C2(n6888), .A(n4261), .B(n4940), .ZN(n4267)
         );
  AND2_X1 U5301 ( .A1(n4935), .A2(n4263), .ZN(n4264) );
  OR2_X1 U5302 ( .A1(n4264), .A2(n5081), .ZN(n5600) );
  NOR2_X1 U5303 ( .A1(n5912), .A2(n6568), .ZN(n5319) );
  INV_X1 U5304 ( .A(n5319), .ZN(n4265) );
  OAI21_X1 U5305 ( .B1(n5600), .B2(n5903), .A(n4265), .ZN(n4266) );
  OR4_X1 U5306 ( .A1(n4269), .A2(n4268), .A3(n4267), .A4(n4266), .ZN(U3002) );
  INV_X1 U5307 ( .A(n6610), .ZN(n4272) );
  OR2_X1 U5308 ( .A1(n4296), .A2(n4270), .ZN(n4281) );
  NOR2_X2 U5309 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6466) );
  NAND2_X1 U5310 ( .A1(n6466), .A2(n4724), .ZN(n4654) );
  INV_X1 U5311 ( .A(n4654), .ZN(n4273) );
  OAI21_X1 U5312 ( .B1(n4273), .B2(READREQUEST_REG_SCAN_IN), .A(n4272), .ZN(
        n4271) );
  OAI21_X1 U5313 ( .B1(n4272), .B2(n4281), .A(n4271), .ZN(U3474) );
  INV_X1 U5314 ( .A(n4299), .ZN(n4295) );
  AOI211_X1 U5315 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4274), .A(n4273), .B(
        n4295), .ZN(n4275) );
  INV_X1 U5316 ( .A(n4275), .ZN(U2788) );
  OR2_X1 U5317 ( .A1(n4317), .A2(n4276), .ZN(n4280) );
  NAND2_X1 U5318 ( .A1(n4278), .A2(n4277), .ZN(n4279) );
  NAND2_X1 U5319 ( .A1(n4280), .A2(n4279), .ZN(n5557) );
  AOI21_X1 U5320 ( .B1(n4281), .B2(n6533), .A(READY_N), .ZN(n6614) );
  NOR2_X1 U5321 ( .A1(n5557), .A2(n6614), .ZN(n4594) );
  OR2_X1 U5322 ( .A1(n4594), .A2(n5556), .ZN(n4292) );
  INV_X1 U5323 ( .A(n4292), .ZN(n5564) );
  INV_X1 U5324 ( .A(MORE_REG_SCAN_IN), .ZN(n4294) );
  NOR2_X1 U5325 ( .A1(n4283), .A2(n4282), .ZN(n4284) );
  OR2_X1 U5326 ( .A1(n4317), .A2(n4284), .ZN(n4291) );
  INV_X1 U5327 ( .A(n4457), .ZN(n4285) );
  NAND2_X1 U5328 ( .A1(n4317), .A2(n4285), .ZN(n4290) );
  INV_X1 U5329 ( .A(n4286), .ZN(n4287) );
  OR2_X1 U5330 ( .A1(n4288), .A2(n4287), .ZN(n4289) );
  AND3_X1 U5331 ( .A1(n4291), .A2(n4290), .A3(n4289), .ZN(n4597) );
  OR2_X1 U5332 ( .A1(n4292), .A2(n4597), .ZN(n4293) );
  OAI21_X1 U5333 ( .B1(n5564), .B2(n4294), .A(n4293), .ZN(U3471) );
  INV_X1 U5334 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n4300) );
  INV_X1 U5335 ( .A(READY_N), .ZN(n6612) );
  OAI21_X1 U5336 ( .B1(n4296), .B2(n6612), .A(n4295), .ZN(n5798) );
  INV_X1 U5337 ( .A(n5798), .ZN(n4410) );
  NAND2_X1 U5338 ( .A1(n4297), .A2(n6612), .ZN(n4298) );
  INV_X1 U5339 ( .A(DATAI_1_), .ZN(n5956) );
  OAI222_X1 U5340 ( .A1(n5803), .A2(n4301), .B1(n4300), .B2(n4410), .C1(n4445), 
        .C2(n5956), .ZN(U2940) );
  INV_X1 U5341 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n4303) );
  INV_X1 U5342 ( .A(DATAI_14_), .ZN(n4302) );
  OAI222_X1 U5343 ( .A1(n5803), .A2(n4684), .B1(n4303), .B2(n4410), .C1(n4445), 
        .C2(n4302), .ZN(U2953) );
  OR2_X1 U5344 ( .A1(n4395), .A2(n4583), .ZN(n4304) );
  NAND2_X1 U5345 ( .A1(n5803), .A2(n4304), .ZN(n4306) );
  NOR2_X1 U5346 ( .A1(n4724), .A2(n6799), .ZN(n4485) );
  NAND2_X1 U5347 ( .A1(n6517), .A2(n4485), .ZN(n5749) );
  INV_X1 U5348 ( .A(n5749), .ZN(n5769) );
  INV_X1 U5349 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n6903) );
  NAND2_X1 U5350 ( .A1(n5768), .A2(n3190), .ZN(n5744) );
  INV_X1 U5351 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n6905) );
  OAI222_X1 U5352 ( .A1(n5762), .A2(n6903), .B1(n5744), .B2(n4179), .C1(n6905), 
        .C2(n5749), .ZN(U2903) );
  INV_X1 U5353 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n6899) );
  INV_X1 U5354 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4308) );
  INV_X1 U5355 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n6919) );
  OAI222_X1 U5356 ( .A1(n5762), .A2(n6899), .B1(n5744), .B2(n4308), .C1(n6919), 
        .C2(n5749), .ZN(U2899) );
  INV_X1 U5357 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n6785) );
  NAND2_X1 U5358 ( .A1(n5801), .A2(DATAI_13_), .ZN(n5799) );
  NAND2_X1 U5359 ( .A1(n5797), .A2(EAX_REG_29__SCAN_IN), .ZN(n4309) );
  OAI211_X1 U5360 ( .C1(n4410), .C2(n6785), .A(n5799), .B(n4309), .ZN(U2937)
         );
  OR2_X1 U5361 ( .A1(n4583), .A2(n3885), .ZN(n4574) );
  INV_X1 U5362 ( .A(n4725), .ZN(n5549) );
  INV_X1 U5363 ( .A(n4310), .ZN(n4312) );
  AOI21_X1 U5364 ( .B1(n4583), .B2(n4329), .A(n6533), .ZN(n4311) );
  OAI211_X1 U5365 ( .C1(n4312), .C2(n4311), .A(n4317), .B(n6612), .ZN(n4315)
         );
  NAND3_X1 U5366 ( .A1(n4315), .A2(n4314), .A3(n4313), .ZN(n4322) );
  NAND2_X1 U5367 ( .A1(n4317), .A2(n4316), .ZN(n4321) );
  NAND2_X1 U5368 ( .A1(n4319), .A2(n4318), .ZN(n4320) );
  NAND2_X1 U5369 ( .A1(n4321), .A2(n4320), .ZN(n4443) );
  NOR2_X1 U5370 ( .A1(n4322), .A2(n4443), .ZN(n4325) );
  NAND2_X1 U5371 ( .A1(n4324), .A2(n4323), .ZN(n4354) );
  NAND2_X1 U5372 ( .A1(n4325), .A2(n4354), .ZN(n4584) );
  NAND2_X1 U5373 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4485), .ZN(n6598) );
  INV_X1 U5374 ( .A(n6598), .ZN(n4614) );
  AOI22_X1 U5375 ( .A1(n4584), .A2(n6515), .B1(n4614), .B2(FLUSH_REG_SCAN_IN), 
        .ZN(n5551) );
  OAI21_X1 U5376 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6600), .A(n5551), .ZN(
        n5554) );
  OAI21_X1 U5377 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5009), .A(n5554), 
        .ZN(n4722) );
  INV_X1 U5378 ( .A(n4326), .ZN(n4328) );
  AND3_X1 U5379 ( .A1(n4329), .A2(n4328), .A3(n4327), .ZN(n4330) );
  AND2_X1 U5380 ( .A1(n5550), .A2(n4330), .ZN(n4332) );
  NAND2_X1 U5381 ( .A1(n4332), .A2(n4331), .ZN(n4577) );
  AND2_X1 U5382 ( .A1(n4580), .A2(n3885), .ZN(n4333) );
  AOI21_X1 U5383 ( .B1(n6244), .B2(n4577), .A(n4333), .ZN(n4576) );
  OAI22_X1 U5384 ( .A1(n4576), .A2(n5549), .B1(n4724), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4334) );
  OAI22_X1 U5385 ( .A1(n4722), .A2(n4334), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5554), .ZN(n4335) );
  OAI21_X1 U5386 ( .B1(n4574), .B2(n5549), .A(n4335), .ZN(U3461) );
  XNOR2_X1 U5387 ( .A(n4336), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4404)
         );
  INV_X1 U5388 ( .A(n4337), .ZN(n4338) );
  OAI21_X1 U5389 ( .B1(n4339), .B2(n4338), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4345) );
  OAI21_X1 U5390 ( .B1(n4930), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4340), 
        .ZN(n5710) );
  INV_X1 U5391 ( .A(n5710), .ZN(n4343) );
  INV_X1 U5392 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6606) );
  OAI21_X1 U5393 ( .B1(n5912), .B2(n6606), .A(n4341), .ZN(n4342) );
  AOI21_X1 U5394 ( .B1(n5927), .B2(n4343), .A(n4342), .ZN(n4344) );
  OAI211_X1 U5395 ( .C1(n4404), .C2(n5906), .A(n4345), .B(n4344), .ZN(U3018)
         );
  NAND2_X1 U5396 ( .A1(n4347), .A2(n4346), .ZN(n4348) );
  AND2_X1 U5397 ( .A1(n4349), .A2(n4348), .ZN(n5715) );
  INV_X1 U5398 ( .A(n5715), .ZN(n4507) );
  INV_X1 U5399 ( .A(n4438), .ZN(n4351) );
  NAND2_X1 U5400 ( .A1(n5987), .A2(n5971), .ZN(n4439) );
  INV_X1 U5401 ( .A(n4439), .ZN(n4350) );
  NAND4_X1 U5402 ( .A1(n4352), .A2(n4351), .A3(n4350), .A4(n4390), .ZN(n4353)
         );
  NAND2_X1 U5403 ( .A1(n4354), .A2(n4353), .ZN(n4355) );
  NAND2_X1 U5404 ( .A1(n5733), .A2(n5987), .ZN(n5720) );
  OAI222_X1 U5405 ( .A1(n4507), .A2(n5203), .B1(n4356), .B2(n5733), .C1(n5710), 
        .C2(n5720), .ZN(U2859) );
  INV_X1 U5406 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6867) );
  AOI22_X1 U5407 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n5769), .B1(n5775), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4357) );
  OAI21_X1 U5408 ( .B1(n6867), .B2(n5744), .A(n4357), .ZN(U2895) );
  INV_X1 U5409 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6887) );
  AOI22_X1 U5410 ( .A1(n5769), .A2(UWORD_REG_0__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4358) );
  OAI21_X1 U5411 ( .B1(n6887), .B2(n5744), .A(n4358), .ZN(U2907) );
  INV_X1 U5412 ( .A(EAX_REG_17__SCAN_IN), .ZN(n5781) );
  AOI22_X1 U5413 ( .A1(n6613), .A2(UWORD_REG_1__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4359) );
  OAI21_X1 U5414 ( .B1(n5781), .B2(n5744), .A(n4359), .ZN(U2906) );
  INV_X1 U5415 ( .A(EAX_REG_30__SCAN_IN), .ZN(n5790) );
  AOI22_X1 U5416 ( .A1(n6613), .A2(UWORD_REG_14__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4360) );
  OAI21_X1 U5417 ( .B1(n5790), .B2(n5744), .A(n4360), .ZN(U2893) );
  INV_X1 U5418 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4362) );
  AOI22_X1 U5419 ( .A1(n5769), .A2(UWORD_REG_7__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4361) );
  OAI21_X1 U5420 ( .B1(n4362), .B2(n5744), .A(n4361), .ZN(U2900) );
  INV_X1 U5421 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4364) );
  AOI22_X1 U5422 ( .A1(n5769), .A2(UWORD_REG_9__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4363) );
  OAI21_X1 U5423 ( .B1(n4364), .B2(n5744), .A(n4363), .ZN(U2898) );
  AOI22_X1 U5424 ( .A1(n5769), .A2(UWORD_REG_10__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4365) );
  OAI21_X1 U5425 ( .B1(n4821), .B2(n5744), .A(n4365), .ZN(U2897) );
  INV_X1 U5426 ( .A(EAX_REG_27__SCAN_IN), .ZN(n5786) );
  AOI22_X1 U5427 ( .A1(n5769), .A2(UWORD_REG_11__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4366) );
  OAI21_X1 U5428 ( .B1(n5786), .B2(n5744), .A(n4366), .ZN(U2896) );
  INV_X1 U5429 ( .A(n4410), .ZN(n4393) );
  AOI22_X1 U5430 ( .A1(n4393), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n5797), .ZN(n4367) );
  NAND2_X1 U5431 ( .A1(n5801), .A2(DATAI_8_), .ZN(n4370) );
  NAND2_X1 U5432 ( .A1(n4367), .A2(n4370), .ZN(U2947) );
  AOI22_X1 U5433 ( .A1(n4393), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n5797), .ZN(n4368) );
  NAND2_X1 U5434 ( .A1(n5801), .A2(DATAI_6_), .ZN(n4373) );
  NAND2_X1 U5435 ( .A1(n4368), .A2(n4373), .ZN(U2930) );
  AOI22_X1 U5436 ( .A1(n4393), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n5797), .ZN(n4369) );
  NAND2_X1 U5437 ( .A1(n5801), .A2(DATAI_3_), .ZN(n4418) );
  NAND2_X1 U5438 ( .A1(n4369), .A2(n4418), .ZN(U2942) );
  AOI22_X1 U5439 ( .A1(n4393), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n5797), .ZN(n4371) );
  NAND2_X1 U5440 ( .A1(n4371), .A2(n4370), .ZN(U2932) );
  AOI22_X1 U5441 ( .A1(n4393), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n5797), .ZN(n4372) );
  NAND2_X1 U5442 ( .A1(n5801), .A2(DATAI_9_), .ZN(n4378) );
  NAND2_X1 U5443 ( .A1(n4372), .A2(n4378), .ZN(U2933) );
  AOI22_X1 U5444 ( .A1(n4393), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n5797), .ZN(n4374) );
  NAND2_X1 U5445 ( .A1(n4374), .A2(n4373), .ZN(U2945) );
  AOI22_X1 U5446 ( .A1(n4393), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n5797), .ZN(n4375) );
  NAND2_X1 U5447 ( .A1(n5801), .A2(DATAI_4_), .ZN(n4376) );
  NAND2_X1 U5448 ( .A1(n4375), .A2(n4376), .ZN(U2943) );
  AOI22_X1 U5449 ( .A1(n4393), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n5797), .ZN(n4377) );
  NAND2_X1 U5450 ( .A1(n4377), .A2(n4376), .ZN(U2928) );
  AOI22_X1 U5451 ( .A1(n4393), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n5797), .ZN(n4379) );
  NAND2_X1 U5452 ( .A1(n4379), .A2(n4378), .ZN(U2948) );
  AOI22_X1 U5453 ( .A1(n4393), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n5797), .ZN(n4380) );
  NAND2_X1 U5454 ( .A1(n5801), .A2(DATAI_2_), .ZN(n4414) );
  NAND2_X1 U5455 ( .A1(n4380), .A2(n4414), .ZN(U2941) );
  AOI22_X1 U5456 ( .A1(n4393), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n5797), .ZN(n4381) );
  INV_X1 U5457 ( .A(DATAI_5_), .ZN(n5977) );
  OR2_X1 U5458 ( .A1(n4445), .A2(n5977), .ZN(n4412) );
  NAND2_X1 U5459 ( .A1(n4381), .A2(n4412), .ZN(U2944) );
  XNOR2_X1 U5460 ( .A(n4383), .B(n4382), .ZN(n4550) );
  NOR2_X1 U5461 ( .A1(n5868), .A2(n4384), .ZN(n4386) );
  MUX2_X1 U5462 ( .A(n4386), .B(n4385), .S(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .Z(n4387) );
  INV_X1 U5463 ( .A(n4387), .ZN(n4392) );
  OAI21_X1 U5464 ( .B1(n5143), .B2(n4390), .A(n4389), .ZN(n4408) );
  AOI22_X1 U5465 ( .A1(n5927), .A2(n4408), .B1(n5931), .B2(REIP_REG_1__SCAN_IN), .ZN(n4391) );
  OAI211_X1 U5466 ( .C1(n4550), .C2(n5906), .A(n4392), .B(n4391), .ZN(U3017)
         );
  INV_X1 U5467 ( .A(DATAI_0_), .ZN(n5942) );
  AOI22_X1 U5468 ( .A1(n4393), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n5797), .ZN(n4394) );
  OAI21_X1 U5469 ( .B1(n5942), .B2(n4445), .A(n4394), .ZN(U2939) );
  INV_X1 U5470 ( .A(n6466), .ZN(n6454) );
  NAND2_X1 U5471 ( .A1(n6454), .A2(n4396), .ZN(n6611) );
  NAND2_X1 U5472 ( .A1(n6611), .A2(n6517), .ZN(n4397) );
  NAND2_X1 U5473 ( .A1(n6517), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4399) );
  NAND2_X1 U5474 ( .A1(n6411), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4398) );
  AND2_X1 U5475 ( .A1(n4399), .A2(n4398), .ZN(n4531) );
  INV_X1 U5476 ( .A(n4531), .ZN(n4400) );
  OAI21_X1 U5477 ( .B1(n5829), .B2(n4400), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4403) );
  NAND2_X1 U5478 ( .A1(n4401), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6523) );
  AOI22_X1 U5479 ( .A1(n5715), .A2(n5851), .B1(n5931), .B2(REIP_REG_0__SCAN_IN), .ZN(n4402) );
  OAI211_X1 U5480 ( .C1(n4404), .C2(n5814), .A(n4403), .B(n4402), .ZN(U2986)
         );
  OR2_X1 U5481 ( .A1(n4406), .A2(n4405), .ZN(n4407) );
  AND2_X1 U5482 ( .A1(n4433), .A2(n4407), .ZN(n5142) );
  INV_X1 U5483 ( .A(n5142), .ZN(n4453) );
  INV_X1 U5484 ( .A(n5733), .ZN(n5201) );
  AOI22_X1 U5485 ( .A1(n5730), .A2(n4408), .B1(EBX_REG_1__SCAN_IN), .B2(n5201), 
        .ZN(n4409) );
  OAI21_X1 U5486 ( .B1(n5203), .B2(n4453), .A(n4409), .ZN(U2858) );
  AOI22_X1 U5487 ( .A1(n4393), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n5797), .ZN(n4411) );
  NAND2_X1 U5488 ( .A1(n5801), .A2(DATAI_7_), .ZN(n4416) );
  NAND2_X1 U5489 ( .A1(n4411), .A2(n4416), .ZN(U2946) );
  AOI22_X1 U5490 ( .A1(n4393), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n5797), .ZN(n4413) );
  NAND2_X1 U5491 ( .A1(n4413), .A2(n4412), .ZN(U2929) );
  AOI22_X1 U5492 ( .A1(n4393), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n5797), .ZN(n4415) );
  NAND2_X1 U5493 ( .A1(n4415), .A2(n4414), .ZN(U2926) );
  AOI22_X1 U5494 ( .A1(n4393), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n5797), .ZN(n4417) );
  NAND2_X1 U5495 ( .A1(n4417), .A2(n4416), .ZN(U2931) );
  AOI22_X1 U5496 ( .A1(n4393), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n5797), .ZN(n4419) );
  NAND2_X1 U5497 ( .A1(n4419), .A2(n4418), .ZN(U2927) );
  INV_X1 U5498 ( .A(n4500), .ZN(n4420) );
  OAI21_X1 U5499 ( .B1(n4432), .B2(n4421), .A(n4420), .ZN(n5123) );
  CLKBUF_X1 U5500 ( .A(n4422), .Z(n5129) );
  OAI21_X1 U5501 ( .B1(n5129), .B2(n5128), .A(n4423), .ZN(n4424) );
  AND2_X1 U5502 ( .A1(n4424), .A2(n4428), .ZN(n5917) );
  AOI22_X1 U5503 ( .A1(n5730), .A2(n5917), .B1(EBX_REG_3__SCAN_IN), .B2(n5201), 
        .ZN(n4425) );
  OAI21_X1 U5504 ( .B1(n5123), .B2(n5203), .A(n4425), .ZN(U2856) );
  INV_X1 U5505 ( .A(n4499), .ZN(n4426) );
  XNOR2_X1 U5506 ( .A(n4500), .B(n4426), .ZN(n5842) );
  INV_X1 U5507 ( .A(n5842), .ZN(n4498) );
  AND2_X1 U5508 ( .A1(n4428), .A2(n4427), .ZN(n4429) );
  OR2_X1 U5509 ( .A1(n4429), .A2(n5682), .ZN(n5902) );
  INV_X1 U5510 ( .A(n5902), .ZN(n4430) );
  AOI22_X1 U5511 ( .A1(n5730), .A2(n4430), .B1(EBX_REG_4__SCAN_IN), .B2(n5201), 
        .ZN(n4431) );
  OAI21_X1 U5512 ( .B1(n4498), .B2(n5203), .A(n4431), .ZN(U2855) );
  INV_X1 U5513 ( .A(n4432), .ZN(n4437) );
  NAND3_X1 U5514 ( .A1(n4435), .A2(n4434), .A3(n4433), .ZN(n4436) );
  NAND2_X1 U5515 ( .A1(n4437), .A2(n4436), .ZN(n5728) );
  NOR2_X1 U5516 ( .A1(n4439), .A2(n4438), .ZN(n4440) );
  AND2_X1 U5517 ( .A1(n4441), .A2(n4440), .ZN(n4442) );
  OAI21_X1 U5518 ( .B1(n4443), .B2(n4442), .A(n6515), .ZN(n4444) );
  NAND2_X1 U5519 ( .A1(n4446), .A2(n4449), .ZN(n4447) );
  INV_X1 U5520 ( .A(n5737), .ZN(n4452) );
  AND2_X1 U5521 ( .A1(n5976), .A2(n4449), .ZN(n4450) );
  INV_X1 U5522 ( .A(n5741), .ZN(n4451) );
  NAND2_X1 U5523 ( .A1(n4452), .A2(n4451), .ZN(n5229) );
  INV_X1 U5524 ( .A(DATAI_2_), .ZN(n5961) );
  OAI222_X1 U5525 ( .A1(n5728), .A2(n5489), .B1(n4685), .B2(n5961), .C1(n5204), 
        .C2(n3893), .ZN(U2889) );
  OAI222_X1 U5526 ( .A1(n4453), .A2(n5489), .B1(n4685), .B2(n5956), .C1(n5204), 
        .C2(n4301), .ZN(U2890) );
  XNOR2_X1 U5527 ( .A(n4455), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4462)
         );
  NAND2_X1 U5528 ( .A1(n4457), .A2(n4456), .ZN(n4466) );
  MUX2_X1 U5529 ( .A(n4458), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4578), 
        .Z(n4459) );
  NOR2_X1 U5530 ( .A1(n4459), .A2(n4474), .ZN(n4460) );
  NAND2_X1 U5531 ( .A1(n4466), .A2(n4460), .ZN(n4461) );
  OAI21_X1 U5532 ( .B1(n4583), .B2(n4462), .A(n4461), .ZN(n4463) );
  AOI21_X1 U5533 ( .B1(n6270), .B2(n4577), .A(n4463), .ZN(n5010) );
  MUX2_X1 U5534 ( .A(n5015), .B(n5010), .S(n4584), .Z(n4591) );
  INV_X1 U5535 ( .A(n4591), .ZN(n4472) );
  OR2_X1 U5536 ( .A1(n4584), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4471)
         );
  INV_X1 U5537 ( .A(n6085), .ZN(n6152) );
  XNOR2_X1 U5538 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4468) );
  XNOR2_X1 U5539 ( .A(n4578), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4465)
         );
  NAND2_X1 U5540 ( .A1(n4466), .A2(n4465), .ZN(n4467) );
  OAI21_X1 U5541 ( .B1(n4468), .B2(n4583), .A(n4467), .ZN(n4469) );
  AOI21_X1 U5542 ( .B1(n6152), .B2(n4577), .A(n4469), .ZN(n4713) );
  NAND2_X1 U5543 ( .A1(n4584), .A2(n4713), .ZN(n4470) );
  AND2_X1 U5544 ( .A1(n4471), .A2(n4470), .ZN(n4590) );
  NAND3_X1 U5545 ( .A1(n4472), .A2(n4590), .A3(n4724), .ZN(n4476) );
  INV_X1 U5546 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5563) );
  NAND2_X1 U5547 ( .A1(n5563), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4480) );
  INV_X1 U5548 ( .A(n4480), .ZN(n4473) );
  NAND2_X1 U5549 ( .A1(n4474), .A2(n4473), .ZN(n4475) );
  NAND2_X1 U5550 ( .A1(n4476), .A2(n4475), .ZN(n4600) );
  INV_X1 U5551 ( .A(n4477), .ZN(n4579) );
  INV_X1 U5552 ( .A(n6340), .ZN(n6089) );
  OR2_X1 U5553 ( .A1(n4478), .A2(n6089), .ZN(n4479) );
  XNOR2_X1 U5554 ( .A(n4479), .B(n5553), .ZN(n5697) );
  OAI22_X1 U5555 ( .A1(n4584), .A2(n5553), .B1(n5550), .B2(n5697), .ZN(n4482)
         );
  NOR2_X1 U5556 ( .A1(n4480), .A2(n5553), .ZN(n4481) );
  AOI21_X1 U5557 ( .B1(n4482), .B2(n4724), .A(n4481), .ZN(n4598) );
  INV_X1 U5558 ( .A(n4598), .ZN(n4483) );
  AOI21_X1 U5559 ( .B1(n4600), .B2(n4579), .A(n4483), .ZN(n4615) );
  AND2_X1 U5560 ( .A1(n4615), .A2(n5563), .ZN(n4484) );
  INV_X1 U5561 ( .A(n6521), .ZN(n6616) );
  OAI21_X1 U5562 ( .B1(n4484), .B2(n6598), .A(n6221), .ZN(n5938) );
  INV_X1 U5563 ( .A(n5938), .ZN(n4497) );
  NAND2_X1 U5564 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6600), .ZN(n5426) );
  INV_X1 U5565 ( .A(n3882), .ZN(n5945) );
  AOI222_X1 U5566 ( .A1(n4615), .A2(n4485), .B1(n6244), .B2(n5426), .C1(n5945), 
        .C2(n6466), .ZN(n4487) );
  NAND2_X1 U5567 ( .A1(n4497), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4486) );
  OAI21_X1 U5568 ( .B1(n4497), .B2(n4487), .A(n4486), .ZN(U3465) );
  NAND2_X1 U5569 ( .A1(n6458), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6302) );
  OAI21_X1 U5570 ( .B1(n6302), .B2(n6216), .A(n6466), .ZN(n5428) );
  AOI21_X1 U5571 ( .B1(n6216), .B2(n6302), .A(n5428), .ZN(n4489) );
  AOI21_X1 U5572 ( .B1(n5426), .B2(n6152), .A(n4489), .ZN(n4491) );
  NAND2_X1 U5573 ( .A1(n4497), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4490) );
  OAI21_X1 U5574 ( .B1(n4497), .B2(n4491), .A(n4490), .ZN(U3463) );
  INV_X1 U5575 ( .A(n6458), .ZN(n4492) );
  AOI21_X1 U5576 ( .B1(n4492), .B2(n6411), .A(n6454), .ZN(n4494) );
  AOI22_X1 U5577 ( .A1(n4494), .A2(n6302), .B1(n6151), .B2(n5426), .ZN(n4496)
         );
  NAND2_X1 U5578 ( .A1(n4497), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4495) );
  OAI21_X1 U5579 ( .B1(n4497), .B2(n4496), .A(n4495), .ZN(U3464) );
  INV_X1 U5580 ( .A(DATAI_4_), .ZN(n6979) );
  OAI222_X1 U5581 ( .A1(n5489), .A2(n4498), .B1(n5204), .B2(n3916), .C1(n6979), 
        .C2(n4685), .ZN(U2887) );
  NAND2_X1 U5582 ( .A1(n4500), .A2(n4499), .ZN(n4503) );
  INV_X1 U5583 ( .A(n4501), .ZN(n4502) );
  NAND2_X1 U5584 ( .A1(n4503), .A2(n4502), .ZN(n4504) );
  AND2_X1 U5585 ( .A1(n4521), .A2(n4504), .ZN(n5834) );
  INV_X1 U5586 ( .A(n5834), .ZN(n4506) );
  OAI222_X1 U5587 ( .A1(n4506), .A2(n5489), .B1(n5977), .B2(n4685), .C1(n4505), 
        .C2(n5204), .ZN(U2886) );
  INV_X1 U5588 ( .A(DATAI_3_), .ZN(n5967) );
  OAI222_X1 U5589 ( .A1(n5123), .A2(n5489), .B1(n4685), .B2(n5967), .C1(n5204), 
        .C2(n3904), .ZN(U2888) );
  INV_X1 U5590 ( .A(EAX_REG_0__SCAN_IN), .ZN(n5778) );
  OAI222_X1 U5591 ( .A1(n4507), .A2(n5489), .B1(n4685), .B2(n5942), .C1(n5204), 
        .C2(n5778), .ZN(U2891) );
  OAI21_X1 U5592 ( .B1(n4510), .B2(n4509), .A(n4508), .ZN(n5823) );
  AOI21_X1 U5593 ( .B1(n5922), .B2(n5933), .A(n5923), .ZN(n5898) );
  NOR2_X1 U5594 ( .A1(n4512), .A2(n5898), .ZN(n4515) );
  OAI21_X1 U5595 ( .B1(n4511), .B2(n5922), .A(n4563), .ZN(n5930) );
  AOI21_X1 U5596 ( .B1(n4513), .B2(n4512), .A(n5930), .ZN(n5896) );
  INV_X1 U5597 ( .A(n5896), .ZN(n4514) );
  MUX2_X1 U5598 ( .A(n4515), .B(n4514), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4516) );
  INV_X1 U5599 ( .A(n4516), .ZN(n4520) );
  INV_X1 U5600 ( .A(n4528), .ZN(n4517) );
  AOI21_X1 U5601 ( .B1(n4518), .B2(n5683), .A(n4517), .ZN(n5672) );
  AOI22_X1 U5602 ( .A1(n5927), .A2(n5672), .B1(n5931), .B2(REIP_REG_6__SCAN_IN), .ZN(n4519) );
  OAI211_X1 U5603 ( .C1(n5823), .C2(n5906), .A(n4520), .B(n4519), .ZN(U3012)
         );
  XOR2_X1 U5604 ( .A(n4522), .B(n4521), .Z(n5824) );
  INV_X1 U5605 ( .A(n5824), .ZN(n4524) );
  AOI22_X1 U5606 ( .A1(n5730), .A2(n5672), .B1(EBX_REG_6__SCAN_IN), .B2(n5201), 
        .ZN(n4523) );
  OAI21_X1 U5607 ( .B1(n4524), .B2(n5203), .A(n4523), .ZN(U2853) );
  INV_X1 U5608 ( .A(EAX_REG_6__SCAN_IN), .ZN(n5767) );
  INV_X1 U5609 ( .A(DATAI_6_), .ZN(n5983) );
  OAI222_X1 U5610 ( .A1(n5489), .A2(n4524), .B1(n5204), .B2(n5767), .C1(n5983), 
        .C2(n4685), .ZN(U2885) );
  INV_X1 U5611 ( .A(n4525), .ZN(n4540) );
  OAI21_X1 U5612 ( .B1(n4527), .B2(n4526), .A(n4540), .ZN(n5660) );
  AOI21_X1 U5613 ( .B1(n4529), .B2(n4528), .A(n4543), .ZN(n5881) );
  AOI22_X1 U5614 ( .A1(n5730), .A2(n5881), .B1(EBX_REG_7__SCAN_IN), .B2(n5201), 
        .ZN(n4530) );
  OAI21_X1 U5615 ( .B1(n5660), .B2(n5203), .A(n4530), .ZN(U2852) );
  INV_X1 U5616 ( .A(DATAI_7_), .ZN(n5989) );
  OAI222_X1 U5617 ( .A1(n5660), .A2(n5489), .B1(n4685), .B2(n5989), .C1(n5204), 
        .C2(n3936), .ZN(U2884) );
  AOI22_X1 U5618 ( .A1(n5829), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n5931), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n4532) );
  OAI21_X1 U5619 ( .B1(n5856), .B2(n5109), .A(n4532), .ZN(n4533) );
  INV_X1 U5620 ( .A(n4533), .ZN(n4537) );
  OR2_X1 U5621 ( .A1(n4535), .A2(n4534), .ZN(n5913) );
  INV_X1 U5622 ( .A(n5814), .ZN(n5850) );
  NAND3_X1 U5623 ( .A1(n5913), .A2(n5914), .A3(n5850), .ZN(n4536) );
  OAI211_X1 U5624 ( .C1(n5123), .C2(n6457), .A(n4537), .B(n4536), .ZN(U2983)
         );
  INV_X1 U5625 ( .A(n4538), .ZN(n4541) );
  INV_X1 U5626 ( .A(n4539), .ZN(n4553) );
  AOI21_X1 U5627 ( .B1(n4541), .B2(n4540), .A(n4553), .ZN(n5655) );
  INV_X1 U5628 ( .A(n5655), .ZN(n4546) );
  NOR2_X1 U5629 ( .A1(n4543), .A2(n4542), .ZN(n4544) );
  OR2_X1 U5630 ( .A1(n5637), .A2(n4544), .ZN(n5649) );
  INV_X1 U5631 ( .A(n5649), .ZN(n4571) );
  AOI22_X1 U5632 ( .A1(n5730), .A2(n4571), .B1(EBX_REG_8__SCAN_IN), .B2(n5201), 
        .ZN(n4545) );
  OAI21_X1 U5633 ( .B1(n4546), .B2(n5203), .A(n4545), .ZN(U2851) );
  INV_X1 U5634 ( .A(DATAI_8_), .ZN(n6809) );
  INV_X1 U5635 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5764) );
  OAI222_X1 U5636 ( .A1(n4546), .A2(n5489), .B1(n4685), .B2(n6809), .C1(n5204), 
        .C2(n5764), .ZN(U2883) );
  AOI22_X1 U5637 ( .A1(n5829), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5931), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4547) );
  OAI21_X1 U5638 ( .B1(n5856), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4547), 
        .ZN(n4548) );
  AOI21_X1 U5639 ( .B1(n5851), .B2(n5142), .A(n4548), .ZN(n4549) );
  OAI21_X1 U5640 ( .B1(n4550), .B2(n5814), .A(n4549), .ZN(U2985) );
  OAI21_X1 U5641 ( .B1(n4553), .B2(n3970), .A(n4619), .ZN(n5643) );
  AOI22_X1 U5642 ( .A1(n5229), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n5740), .ZN(n4554) );
  OAI21_X1 U5643 ( .B1(n5643), .B2(n5489), .A(n4554), .ZN(U2882) );
  OAI21_X1 U5644 ( .B1(n4557), .B2(n4556), .A(n4555), .ZN(n4573) );
  INV_X1 U5645 ( .A(REIP_REG_8__SCAN_IN), .ZN(n4558) );
  NOR2_X1 U5646 ( .A1(n5912), .A2(n4558), .ZN(n4570) );
  AOI21_X1 U5647 ( .B1(n5829), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n4570), 
        .ZN(n4559) );
  OAI21_X1 U5648 ( .B1(n5856), .B2(n5652), .A(n4559), .ZN(n4560) );
  AOI21_X1 U5649 ( .B1(n5655), .B2(n5851), .A(n4560), .ZN(n4561) );
  OAI21_X1 U5650 ( .B1(n4573), .B2(n5814), .A(n4561), .ZN(U2978) );
  NOR2_X1 U5651 ( .A1(n4562), .A2(n5898), .ZN(n5883) );
  OAI21_X1 U5652 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n5883), .ZN(n4568) );
  OAI21_X1 U5653 ( .B1(n4564), .B2(n5897), .A(n4563), .ZN(n4565) );
  AOI21_X1 U5654 ( .B1(n4567), .B2(n4566), .A(n4565), .ZN(n5886) );
  OAI22_X1 U5655 ( .A1(n5867), .A2(n4568), .B1(n5886), .B2(n6931), .ZN(n4569)
         );
  AOI211_X1 U5656 ( .C1(n5927), .C2(n4571), .A(n4570), .B(n4569), .ZN(n4572)
         );
  OAI21_X1 U5657 ( .B1(n5906), .B2(n4573), .A(n4572), .ZN(U3010) );
  AND2_X1 U5658 ( .A1(n4574), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4575)
         );
  AND2_X1 U5659 ( .A1(n4576), .A2(n4575), .ZN(n4588) );
  NAND2_X1 U5660 ( .A1(n6151), .A2(n4577), .ZN(n4582) );
  INV_X1 U5661 ( .A(n4578), .ZN(n4716) );
  NAND3_X1 U5662 ( .A1(n4580), .A2(n4716), .A3(n4579), .ZN(n4581) );
  OAI211_X1 U5663 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n4583), .A(n4582), .B(n4581), .ZN(n4726) );
  INV_X1 U5664 ( .A(n4584), .ZN(n4585) );
  AOI21_X1 U5665 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n4588), .A(n4585), 
        .ZN(n4586) );
  NAND2_X1 U5666 ( .A1(n4726), .A2(n4586), .ZN(n4587) );
  OAI21_X1 U5667 ( .B1(n4588), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n4587), 
        .ZN(n4589) );
  AOI222_X1 U5668 ( .A1(n6213), .A2(n4590), .B1(n6213), .B2(n4589), .C1(n4590), 
        .C2(n4589), .ZN(n4592) );
  AND2_X1 U5669 ( .A1(n4592), .A2(n4591), .ZN(n4593) );
  OAI22_X1 U5670 ( .A1(n4593), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(n4592), .B2(n4591), .ZN(n4602) );
  OAI21_X1 U5671 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n4594), 
        .ZN(n4595) );
  NAND4_X1 U5672 ( .A1(n4598), .A2(n4597), .A3(n4596), .A4(n4595), .ZN(n4599)
         );
  OR2_X1 U5673 ( .A1(n4600), .A2(n4599), .ZN(n4601) );
  AOI21_X1 U5674 ( .B1(n4602), .B2(n6972), .A(n4601), .ZN(n4618) );
  NOR2_X1 U5675 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6612), .ZN(n6525) );
  NAND2_X1 U5676 ( .A1(n4618), .A2(n6515), .ZN(n4604) );
  NAND2_X1 U5677 ( .A1(READY_N), .A2(n6613), .ZN(n4603) );
  NAND2_X1 U5678 ( .A1(n4604), .A2(n4603), .ZN(n4609) );
  INV_X1 U5679 ( .A(n4605), .ZN(n4606) );
  OR2_X1 U5680 ( .A1(n4607), .A2(n4606), .ZN(n4608) );
  NOR2_X1 U5681 ( .A1(n6525), .A2(n6597), .ZN(n4611) );
  OAI21_X1 U5682 ( .B1(n6521), .B2(n5009), .A(n6517), .ZN(n4610) );
  OAI22_X1 U5683 ( .A1(n6517), .A2(n4611), .B1(n6597), .B2(n4610), .ZN(n4612)
         );
  INV_X1 U5684 ( .A(n4612), .ZN(n4617) );
  AOI21_X1 U5685 ( .B1(n4615), .B2(n4614), .A(n4613), .ZN(n4616) );
  OAI211_X1 U5686 ( .C1(n4618), .C2(n5556), .A(n4617), .B(n4616), .ZN(U3148)
         );
  NOR2_X1 U5687 ( .A1(n4619), .A2(n4620), .ZN(n4633) );
  AOI21_X1 U5688 ( .B1(n4620), .B2(n4619), .A(n4633), .ZN(n4621) );
  INV_X1 U5689 ( .A(n4621), .ZN(n5107) );
  AOI22_X1 U5690 ( .A1(n5229), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n5740), .ZN(n4622) );
  OAI21_X1 U5691 ( .B1(n5107), .B2(n5489), .A(n4622), .ZN(U2881) );
  XNOR2_X1 U5692 ( .A(n4635), .B(n4637), .ZN(n5866) );
  INV_X1 U5693 ( .A(n5866), .ZN(n4623) );
  OAI222_X1 U5694 ( .A1(n5107), .A2(n5203), .B1(n4624), .B2(n5733), .C1(n5720), 
        .C2(n4623), .ZN(U2849) );
  XNOR2_X1 U5695 ( .A(n5806), .B(n4626), .ZN(n4627) );
  XNOR2_X1 U5696 ( .A(n4625), .B(n4627), .ZN(n5877) );
  NAND2_X1 U5697 ( .A1(n5877), .A2(n5850), .ZN(n4631) );
  INV_X1 U5698 ( .A(n5829), .ZN(n5297) );
  INV_X1 U5699 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4628) );
  NAND2_X1 U5700 ( .A1(n5931), .A2(REIP_REG_9__SCAN_IN), .ZN(n5873) );
  OAI21_X1 U5701 ( .B1(n5297), .B2(n4628), .A(n5873), .ZN(n4629) );
  AOI21_X1 U5702 ( .B1(n5810), .B2(n5644), .A(n4629), .ZN(n4630) );
  OAI211_X1 U5703 ( .C1(n6457), .C2(n5643), .A(n4631), .B(n4630), .ZN(U2977)
         );
  NAND2_X1 U5704 ( .A1(n4633), .A2(n4632), .ZN(n4649) );
  OR2_X1 U5705 ( .A1(n4633), .A2(n4632), .ZN(n4634) );
  INV_X1 U5706 ( .A(n4635), .ZN(n5638) );
  AOI21_X1 U5707 ( .B1(n5638), .B2(n4637), .A(n4636), .ZN(n4639) );
  INV_X1 U5708 ( .A(n4656), .ZN(n4638) );
  NOR2_X1 U5709 ( .A1(n4639), .A2(n4638), .ZN(n5858) );
  AOI22_X1 U5710 ( .A1(n5730), .A2(n5858), .B1(EBX_REG_11__SCAN_IN), .B2(n5201), .ZN(n4640) );
  OAI21_X1 U5711 ( .B1(n5097), .B2(n5203), .A(n4640), .ZN(U2848) );
  AOI22_X1 U5712 ( .A1(n5229), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n5740), .ZN(n4641) );
  OAI21_X1 U5713 ( .B1(n5097), .B2(n5489), .A(n4641), .ZN(U2880) );
  NAND2_X1 U5714 ( .A1(n5804), .A2(n4643), .ZN(n4644) );
  XNOR2_X1 U5715 ( .A(n4642), .B(n4644), .ZN(n5869) );
  NAND2_X1 U5716 ( .A1(n5869), .A2(n5850), .ZN(n4648) );
  INV_X1 U5717 ( .A(REIP_REG_10__SCAN_IN), .ZN(n4645) );
  NOR2_X1 U5718 ( .A1(n5912), .A2(n4645), .ZN(n5865) );
  NOR2_X1 U5719 ( .A1(n5856), .A2(n5099), .ZN(n4646) );
  AOI211_X1 U5720 ( .C1(n5829), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5865), 
        .B(n4646), .ZN(n4647) );
  OAI211_X1 U5721 ( .C1(n6457), .C2(n5107), .A(n4648), .B(n4647), .ZN(U2976)
         );
  XOR2_X1 U5722 ( .A(n4650), .B(n4649), .Z(n4961) );
  AOI22_X1 U5723 ( .A1(n5229), .A2(DATAI_12_), .B1(EAX_REG_12__SCAN_IN), .B2(
        n5740), .ZN(n4651) );
  OAI21_X1 U5724 ( .B1(n4667), .B2(n5489), .A(n4651), .ZN(U2879) );
  INV_X1 U5725 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6562) );
  NAND2_X1 U5726 ( .A1(n4663), .A2(n6562), .ZN(n4652) );
  NOR2_X1 U5727 ( .A1(n5667), .A2(n4652), .ZN(n5631) );
  INV_X1 U5728 ( .A(n4959), .ZN(n4653) );
  NAND2_X1 U5729 ( .A1(n5654), .A2(n4653), .ZN(n4661) );
  INV_X1 U5730 ( .A(n5591), .ZN(n5137) );
  NOR2_X2 U5731 ( .A1(n5137), .A2(n4654), .ZN(n5695) );
  AND2_X1 U5732 ( .A1(n4656), .A2(n4655), .ZN(n4657) );
  OR2_X1 U5733 ( .A1(n4657), .A2(n5540), .ZN(n4952) );
  OAI22_X1 U5734 ( .A1(n6845), .A2(n5718), .B1(n5711), .B2(n4952), .ZN(n4659)
         );
  INV_X1 U5735 ( .A(n5699), .ZN(n5708) );
  NOR2_X1 U5736 ( .A1(n3769), .A2(n5708), .ZN(n4658) );
  NOR3_X1 U5737 ( .A1(n5695), .A2(n4659), .A3(n4658), .ZN(n4660) );
  NAND2_X1 U5738 ( .A1(n4661), .A2(n4660), .ZN(n4662) );
  NOR2_X1 U5739 ( .A1(n5631), .A2(n4662), .ZN(n4666) );
  OR2_X1 U5740 ( .A1(n5667), .A2(n4663), .ZN(n4664) );
  NAND2_X1 U5741 ( .A1(n4664), .A2(n5591), .ZN(n5632) );
  NAND2_X1 U5742 ( .A1(n5632), .A2(REIP_REG_12__SCAN_IN), .ZN(n4665) );
  OAI211_X1 U5743 ( .C1(n4667), .C2(n5479), .A(n4666), .B(n4665), .ZN(U2815)
         );
  OAI222_X1 U5744 ( .A1(n4952), .A2(n5720), .B1(n5733), .B2(n3769), .C1(n5203), 
        .C2(n4667), .ZN(U2847) );
  INV_X1 U5745 ( .A(n4668), .ZN(n4671) );
  INV_X1 U5746 ( .A(n4669), .ZN(n4670) );
  NAND2_X1 U5747 ( .A1(n4671), .A2(n4670), .ZN(n4673) );
  AND2_X1 U5748 ( .A1(n4673), .A2(n4672), .ZN(n5722) );
  INV_X1 U5749 ( .A(n5722), .ZN(n4676) );
  INV_X1 U5750 ( .A(DATAI_13_), .ZN(n4675) );
  OAI222_X1 U5751 ( .A1(n4676), .A2(n5489), .B1(n4675), .B2(n4685), .C1(n4674), 
        .C2(n5204), .ZN(U2878) );
  OAI21_X1 U5752 ( .B1(n4679), .B2(n4678), .A(n4943), .ZN(n5616) );
  INV_X1 U5753 ( .A(EBX_REG_14__SCAN_IN), .ZN(n4683) );
  OR2_X1 U5754 ( .A1(n5542), .A2(n4681), .ZN(n4682) );
  NAND2_X1 U5755 ( .A1(n4680), .A2(n4682), .ZN(n5613) );
  OAI222_X1 U5756 ( .A1(n5616), .A2(n5203), .B1(n4683), .B2(n5733), .C1(n5720), 
        .C2(n5613), .ZN(U2845) );
  OAI222_X1 U5757 ( .A1(n5616), .A2(n5489), .B1(n4302), .B2(n4685), .C1(n4684), 
        .C2(n5204), .ZN(U2877) );
  OR2_X1 U5758 ( .A1(n5516), .A2(n4687), .ZN(n4689) );
  NAND2_X1 U5759 ( .A1(n4689), .A2(n4688), .ZN(n4693) );
  NOR2_X1 U5760 ( .A1(n4691), .A2(n4690), .ZN(n4692) );
  XNOR2_X1 U5761 ( .A(n4693), .B(n4692), .ZN(n4705) );
  NAND2_X1 U5762 ( .A1(n4705), .A2(n5850), .ZN(n4697) );
  INV_X1 U5763 ( .A(REIP_REG_14__SCAN_IN), .ZN(n4694) );
  NOR2_X1 U5764 ( .A1(n5912), .A2(n4694), .ZN(n4706) );
  AND2_X1 U5765 ( .A1(n5829), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4695)
         );
  AOI211_X1 U5766 ( .C1(n5810), .C2(n5617), .A(n4706), .B(n4695), .ZN(n4696)
         );
  OAI211_X1 U5767 ( .C1(n6457), .C2(n5616), .A(n4697), .B(n4696), .ZN(U2972)
         );
  NOR2_X1 U5768 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n4699), .ZN(n5538)
         );
  INV_X1 U5769 ( .A(n5860), .ZN(n4698) );
  AOI21_X1 U5770 ( .B1(n4700), .B2(n4699), .A(n4698), .ZN(n4701) );
  OAI21_X1 U5771 ( .B1(n4703), .B2(n4702), .A(n4701), .ZN(n5543) );
  AOI21_X1 U5772 ( .B1(n5538), .B2(n4704), .A(n5543), .ZN(n4712) );
  NAND2_X1 U5773 ( .A1(n4705), .A2(n5929), .ZN(n4710) );
  NOR2_X1 U5774 ( .A1(n5903), .A2(n5613), .ZN(n4707) );
  AOI211_X1 U5775 ( .C1(n4708), .C2(n4711), .A(n4707), .B(n4706), .ZN(n4709)
         );
  OAI211_X1 U5776 ( .C1(n4712), .C2(n4711), .A(n4710), .B(n4709), .ZN(U3004)
         );
  INV_X1 U5777 ( .A(n5009), .ZN(n5011) );
  INV_X1 U5778 ( .A(n5554), .ZN(n4731) );
  AOI21_X1 U5779 ( .B1(n4716), .B2(n5011), .A(n4731), .ZN(n5016) );
  INV_X1 U5780 ( .A(n4713), .ZN(n4719) );
  INV_X1 U5781 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4715) );
  AOI22_X1 U5782 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4715), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4714), .ZN(n4728) );
  NOR3_X1 U5783 ( .A1(n4724), .A2(n4723), .A3(n4728), .ZN(n4718) );
  NOR3_X1 U5784 ( .A1(n4716), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5009), 
        .ZN(n4717) );
  AOI211_X1 U5785 ( .C1(n4719), .C2(n4725), .A(n4718), .B(n4717), .ZN(n4720)
         );
  OAI22_X1 U5786 ( .A1(n5016), .A2(n4721), .B1(n4731), .B2(n4720), .ZN(U3459)
         );
  INV_X1 U5787 ( .A(n4722), .ZN(n4733) );
  NOR2_X1 U5788 ( .A1(n4724), .A2(n4723), .ZN(n4727) );
  AOI222_X1 U5789 ( .A1(n5011), .A2(n4729), .B1(n4728), .B2(n4727), .C1(n4726), 
        .C2(n4725), .ZN(n4730) );
  OAI22_X1 U5790 ( .A1(n4733), .A2(n4732), .B1(n4731), .B2(n4730), .ZN(U3460)
         );
  NAND2_X1 U5791 ( .A1(n5303), .A2(n4737), .ZN(n4746) );
  NAND2_X1 U5792 ( .A1(n5304), .A2(n5377), .ZN(n4745) );
  INV_X1 U5793 ( .A(n4933), .ZN(n4736) );
  INV_X1 U5794 ( .A(n4734), .ZN(n4735) );
  NAND2_X1 U5795 ( .A1(n4736), .A2(n4735), .ZN(n4738) );
  XNOR2_X1 U5796 ( .A(n5806), .B(n5418), .ZN(n5295) );
  INV_X1 U5797 ( .A(n5295), .ZN(n4739) );
  NAND2_X1 U5798 ( .A1(n5293), .A2(n4739), .ZN(n4741) );
  NAND2_X1 U5799 ( .A1(n5304), .A2(n5418), .ZN(n4740) );
  INV_X1 U5800 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U5801 ( .A1(n5304), .A2(n5402), .ZN(n4743) );
  NOR2_X1 U5802 ( .A1(n5806), .A2(n5402), .ZN(n4742) );
  XNOR2_X1 U5803 ( .A(n5806), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5287)
         );
  NOR2_X1 U5804 ( .A1(n5304), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4759)
         );
  NAND2_X1 U5805 ( .A1(n4744), .A2(n4759), .ZN(n5280) );
  OAI21_X1 U5806 ( .B1(n4746), .B2(n4745), .A(n5280), .ZN(n4748) );
  NAND2_X1 U5807 ( .A1(n5382), .A2(n5850), .ZN(n4753) );
  INV_X1 U5808 ( .A(REIP_REG_23__SCAN_IN), .ZN(n4749) );
  NOR2_X1 U5809 ( .A1(n5912), .A2(n4749), .ZN(n5375) );
  NOR2_X1 U5810 ( .A1(n5297), .A2(n6970), .ZN(n4750) );
  AOI211_X1 U5811 ( .C1(n5810), .C2(n4751), .A(n5375), .B(n4750), .ZN(n4752)
         );
  OAI211_X1 U5812 ( .C1(n6457), .C2(n5223), .A(n4753), .B(n4752), .ZN(U2963)
         );
  NAND2_X1 U5813 ( .A1(n5179), .A2(n4754), .ZN(n4756) );
  NAND2_X1 U5814 ( .A1(n4756), .A2(n4755), .ZN(n4757) );
  NAND2_X1 U5815 ( .A1(n4758), .A2(n4757), .ZN(n5162) );
  AOI21_X1 U5816 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5806), .A(n4759), 
        .ZN(n4760) );
  XOR2_X1 U5817 ( .A(n4760), .B(n5279), .Z(n5391) );
  NAND2_X1 U5818 ( .A1(n5391), .A2(n5850), .ZN(n4764) );
  INV_X1 U5819 ( .A(REIP_REG_22__SCAN_IN), .ZN(n4761) );
  OR2_X1 U5820 ( .A1(n5912), .A2(n4761), .ZN(n5387) );
  OAI21_X1 U5821 ( .B1(n5297), .B2(n5457), .A(n5387), .ZN(n4762) );
  AOI21_X1 U5822 ( .B1(n5461), .B2(n5810), .A(n4762), .ZN(n4763) );
  OAI211_X1 U5823 ( .C1(n6457), .C2(n5162), .A(n4764), .B(n4763), .ZN(U2964)
         );
  AOI22_X1 U5824 ( .A1(n4894), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4769) );
  AOI22_X1 U5825 ( .A1(n4765), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4768) );
  AOI22_X1 U5826 ( .A1(n4898), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4767) );
  AOI22_X1 U5827 ( .A1(n4869), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4766) );
  NAND4_X1 U5828 ( .A1(n4769), .A2(n4768), .A3(n4767), .A4(n4766), .ZN(n4775)
         );
  AOI22_X1 U5829 ( .A1(n3420), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4868), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4773) );
  AOI22_X1 U5830 ( .A1(n4874), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4772) );
  AOI22_X1 U5831 ( .A1(n3187), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4771) );
  AOI22_X1 U5832 ( .A1(n4905), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4770) );
  NAND4_X1 U5833 ( .A1(n4773), .A2(n4772), .A3(n4771), .A4(n4770), .ZN(n4774)
         );
  OR2_X1 U5834 ( .A1(n4775), .A2(n4774), .ZN(n4793) );
  INV_X1 U5835 ( .A(n4793), .ZN(n4778) );
  NAND2_X1 U5836 ( .A1(n4777), .A2(n4776), .ZN(n4794) );
  OR2_X1 U5837 ( .A1(n4778), .A2(n4794), .ZN(n4819) );
  AOI22_X1 U5838 ( .A1(n4893), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4869), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4782) );
  AOI22_X1 U5839 ( .A1(n4894), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4868), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4781) );
  AOI22_X1 U5840 ( .A1(n3404), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4780) );
  AOI22_X1 U5841 ( .A1(n3399), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4779) );
  NAND4_X1 U5842 ( .A1(n4782), .A2(n4781), .A3(n4780), .A4(n4779), .ZN(n4788)
         );
  AOI22_X1 U5843 ( .A1(n3187), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4874), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4786) );
  AOI22_X1 U5844 ( .A1(n3420), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4905), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4785) );
  AOI22_X1 U5845 ( .A1(n4811), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4784) );
  AOI22_X1 U5846 ( .A1(n3405), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4783) );
  NAND4_X1 U5847 ( .A1(n4786), .A2(n4785), .A3(n4784), .A4(n4783), .ZN(n4787)
         );
  NOR2_X1 U5848 ( .A1(n4788), .A2(n4787), .ZN(n4820) );
  XOR2_X1 U5849 ( .A(n4819), .B(n4820), .Z(n4790) );
  OAI22_X1 U5850 ( .A1(n4861), .A2(n4364), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5269), .ZN(n4789) );
  AOI21_X1 U5851 ( .B1(n4790), .B2(n4844), .A(n4789), .ZN(n4792) );
  XNOR2_X1 U5852 ( .A(n4791), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5440)
         );
  MUX2_X1 U5853 ( .A(n4792), .B(n5440), .S(n4918), .Z(n5274) );
  INV_X1 U5854 ( .A(n5274), .ZN(n4805) );
  XNOR2_X1 U5855 ( .A(n4794), .B(n4793), .ZN(n4795) );
  NAND2_X1 U5856 ( .A1(n4844), .A2(n4795), .ZN(n4801) );
  INV_X1 U5857 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5448) );
  XNOR2_X1 U5858 ( .A(n4796), .B(n5448), .ZN(n5451) );
  OAI22_X1 U5859 ( .A1(n5451), .A2(n4798), .B1(n5448), .B2(n4797), .ZN(n4799)
         );
  AOI21_X1 U5860 ( .B1(n4965), .B2(EAX_REG_24__SCAN_IN), .A(n4799), .ZN(n4800)
         );
  NAND2_X1 U5861 ( .A1(n4801), .A2(n4800), .ZN(n5159) );
  INV_X1 U5862 ( .A(n5159), .ZN(n4803) );
  OR2_X1 U5863 ( .A1(n4803), .A2(n4802), .ZN(n4804) );
  NOR2_X1 U5864 ( .A1(n4804), .A2(n5189), .ZN(n5272) );
  AND2_X1 U5865 ( .A1(n4805), .A2(n5272), .ZN(n4806) );
  AOI22_X1 U5866 ( .A1(n4869), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4905), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4810) );
  AOI22_X1 U5867 ( .A1(n4894), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3420), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4809) );
  AOI22_X1 U5868 ( .A1(n4904), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3404), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4808) );
  AOI22_X1 U5869 ( .A1(n4898), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4807) );
  NAND4_X1 U5870 ( .A1(n4810), .A2(n4809), .A3(n4808), .A4(n4807), .ZN(n4818)
         );
  AOI22_X1 U5871 ( .A1(n4896), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4816) );
  AOI22_X1 U5872 ( .A1(n4765), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4815) );
  AOI22_X1 U5873 ( .A1(n3187), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4814) );
  AOI22_X1 U5874 ( .A1(n3418), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4813) );
  NAND4_X1 U5875 ( .A1(n4816), .A2(n4815), .A3(n4814), .A4(n4813), .ZN(n4817)
         );
  NOR2_X1 U5876 ( .A1(n4818), .A2(n4817), .ZN(n4832) );
  OR2_X1 U5877 ( .A1(n4820), .A2(n4819), .ZN(n4831) );
  XOR2_X1 U5878 ( .A(n4832), .B(n4831), .Z(n4823) );
  INV_X1 U5879 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4821) );
  OAI22_X1 U5880 ( .A1(n4861), .A2(n4821), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4824), .ZN(n4822) );
  AOI21_X1 U5881 ( .B1(n4823), .B2(n4844), .A(n4822), .ZN(n4828) );
  AND2_X1 U5882 ( .A1(n4825), .A2(n4824), .ZN(n4826) );
  OR2_X1 U5883 ( .A1(n4826), .A2(n4847), .ZN(n5438) );
  INV_X1 U5884 ( .A(n5438), .ZN(n4827) );
  MUX2_X1 U5885 ( .A(n4828), .B(n4827), .S(n4918), .Z(n5150) );
  INV_X1 U5886 ( .A(n5150), .ZN(n4829) );
  NAND2_X1 U5887 ( .A1(n5076), .A2(n4830), .ZN(n5053) );
  OR2_X1 U5888 ( .A1(n4832), .A2(n4831), .ZN(n4859) );
  AOI22_X1 U5889 ( .A1(n4765), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3419), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4836) );
  AOI22_X1 U5890 ( .A1(n4896), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4835) );
  AOI22_X1 U5891 ( .A1(n3399), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4834) );
  AOI22_X1 U5892 ( .A1(n4869), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4833) );
  NAND4_X1 U5893 ( .A1(n4836), .A2(n4835), .A3(n4834), .A4(n4833), .ZN(n4842)
         );
  AOI22_X1 U5894 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4894), .B1(n3367), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4840) );
  AOI22_X1 U5895 ( .A1(n4904), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4839) );
  AOI22_X1 U5896 ( .A1(n3187), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4838) );
  AOI22_X1 U5897 ( .A1(n4905), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4837) );
  NAND4_X1 U5898 ( .A1(n4840), .A2(n4839), .A3(n4838), .A4(n4837), .ZN(n4841)
         );
  NOR2_X1 U5899 ( .A1(n4842), .A2(n4841), .ZN(n4860) );
  XOR2_X1 U5900 ( .A(n4859), .B(n4860), .Z(n4845) );
  INV_X1 U5901 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4846) );
  OAI22_X1 U5902 ( .A1(n4861), .A2(n5786), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4846), .ZN(n4843) );
  AOI21_X1 U5903 ( .B1(n4845), .B2(n4844), .A(n4843), .ZN(n4848) );
  XNOR2_X1 U5904 ( .A(n4847), .B(n4846), .ZN(n5061) );
  MUX2_X1 U5905 ( .A(n4848), .B(n5061), .S(n4918), .Z(n5055) );
  NOR2_X2 U5906 ( .A1(n5053), .A2(n5055), .ZN(n5054) );
  AOI22_X1 U5907 ( .A1(n4894), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4852) );
  AOI22_X1 U5908 ( .A1(n3419), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4851) );
  AOI22_X1 U5909 ( .A1(n4904), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4850) );
  AOI22_X1 U5910 ( .A1(n4905), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4849) );
  NAND4_X1 U5911 ( .A1(n4852), .A2(n4851), .A3(n4850), .A4(n4849), .ZN(n4858)
         );
  AOI22_X1 U5912 ( .A1(n4765), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4856) );
  AOI22_X1 U5913 ( .A1(n4896), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4855) );
  AOI22_X1 U5914 ( .A1(n3187), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4854) );
  AOI22_X1 U5915 ( .A1(n4869), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4853) );
  NAND4_X1 U5916 ( .A1(n4856), .A2(n4855), .A3(n4854), .A4(n4853), .ZN(n4857)
         );
  NOR2_X1 U5917 ( .A1(n4858), .A2(n4857), .ZN(n4882) );
  OR2_X1 U5918 ( .A1(n4860), .A2(n4859), .ZN(n4881) );
  XNOR2_X1 U5919 ( .A(n4882), .B(n4881), .ZN(n4864) );
  INV_X1 U5920 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6916) );
  OAI22_X1 U5921 ( .A1(n4861), .A2(n6867), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6916), .ZN(n4862) );
  INV_X1 U5922 ( .A(n4862), .ZN(n4863) );
  OAI21_X1 U5923 ( .B1(n4864), .B2(n4915), .A(n4863), .ZN(n4867) );
  OR2_X1 U5924 ( .A1(n4865), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4866)
         );
  NAND2_X1 U5925 ( .A1(n4886), .A2(n4866), .ZN(n5246) );
  MUX2_X1 U5926 ( .A(n4867), .B(n5246), .S(n4918), .Z(n5039) );
  NAND2_X1 U5927 ( .A1(n5054), .A2(n5039), .ZN(n5028) );
  AOI22_X1 U5928 ( .A1(n3419), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4905), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4873) );
  AOI22_X1 U5929 ( .A1(n4765), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4868), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4872) );
  AOI22_X1 U5930 ( .A1(n3404), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4871) );
  AOI22_X1 U5931 ( .A1(n4869), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3405), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4870) );
  NAND4_X1 U5932 ( .A1(n4873), .A2(n4872), .A3(n4871), .A4(n4870), .ZN(n4880)
         );
  AOI22_X1 U5933 ( .A1(n4894), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4811), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4878) );
  AOI22_X1 U5934 ( .A1(n3187), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4874), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4877) );
  AOI22_X1 U5935 ( .A1(n4898), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3497), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4876) );
  AOI22_X1 U5936 ( .A1(n4895), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4875) );
  NAND4_X1 U5937 ( .A1(n4878), .A2(n4877), .A3(n4876), .A4(n4875), .ZN(n4879)
         );
  NOR2_X1 U5938 ( .A1(n4880), .A2(n4879), .ZN(n4891) );
  OR2_X1 U5939 ( .A1(n4882), .A2(n4881), .ZN(n4892) );
  XNOR2_X1 U5940 ( .A(n4891), .B(n4892), .ZN(n4884) );
  AOI22_X1 U5941 ( .A1(n4965), .A2(EAX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6799), .ZN(n4883) );
  OAI21_X1 U5942 ( .B1(n4884), .B2(n4915), .A(n4883), .ZN(n4888) );
  NAND2_X1 U5943 ( .A1(n4886), .A2(n4885), .ZN(n4887) );
  NAND2_X1 U5944 ( .A1(n4917), .A2(n4887), .ZN(n5240) );
  MUX2_X1 U5945 ( .A(n4888), .B(n5240), .S(n4918), .Z(n5030) );
  INV_X1 U5946 ( .A(n5030), .ZN(n4889) );
  NOR2_X1 U5947 ( .A1(n4892), .A2(n4891), .ZN(n4913) );
  AOI22_X1 U5948 ( .A1(n4893), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3419), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4902) );
  AOI22_X1 U5949 ( .A1(n4894), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4901) );
  AOI22_X1 U5950 ( .A1(n4896), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4895), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4900) );
  AOI22_X1 U5951 ( .A1(n4898), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4897), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4899) );
  NAND4_X1 U5952 ( .A1(n4902), .A2(n4901), .A3(n4900), .A4(n4899), .ZN(n4911)
         );
  AOI22_X1 U5953 ( .A1(n3187), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4909) );
  AOI22_X1 U5954 ( .A1(n4869), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3418), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4908) );
  AOI22_X1 U5955 ( .A1(n4904), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4903), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4907) );
  AOI22_X1 U5956 ( .A1(n4905), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4812), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4906) );
  NAND4_X1 U5957 ( .A1(n4909), .A2(n4908), .A3(n4907), .A4(n4906), .ZN(n4910)
         );
  NOR2_X1 U5958 ( .A1(n4911), .A2(n4910), .ZN(n4912) );
  XOR2_X1 U5959 ( .A(n4913), .B(n4912), .Z(n4916) );
  AOI22_X1 U5960 ( .A1(n4965), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6799), .ZN(n4914) );
  OAI21_X1 U5961 ( .B1(n4916), .B2(n4915), .A(n4914), .ZN(n4919) );
  XNOR2_X1 U5962 ( .A(n4917), .B(n5018), .ZN(n5017) );
  MUX2_X1 U5963 ( .A(n4919), .B(n5017), .S(n4918), .Z(n4921) );
  NAND2_X1 U5964 ( .A1(n4920), .A2(n4921), .ZN(n4967) );
  OAI21_X1 U5965 ( .B1(n4890), .B2(n4921), .A(n4967), .ZN(n5209) );
  INV_X1 U5966 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5024) );
  OAI222_X1 U5967 ( .A1(n5203), .A2(n5209), .B1(n5024), .B2(n5733), .C1(n4922), 
        .C2(n5720), .ZN(U2829) );
  NAND2_X1 U5968 ( .A1(n4923), .A2(n3188), .ZN(n4929) );
  INV_X1 U5969 ( .A(n4924), .ZN(n4926) );
  OAI22_X1 U5970 ( .A1(n4926), .A2(n5181), .B1(EBX_REG_29__SCAN_IN), .B2(n4925), .ZN(n5035) );
  NAND3_X1 U5971 ( .A1(n5045), .A2(n4927), .A3(n5035), .ZN(n4928) );
  NAND2_X1 U5972 ( .A1(n4929), .A2(n4928), .ZN(n4932) );
  OAI22_X1 U5973 ( .A1(n4930), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n3734), .ZN(n4931) );
  XNOR2_X2 U5974 ( .A(n4932), .B(n4931), .ZN(n4977) );
  OAI22_X1 U5975 ( .A1(n4977), .A2(n5720), .B1(n5733), .B2(n4235), .ZN(U2828)
         );
  INV_X1 U5976 ( .A(n5303), .ZN(n5309) );
  AOI21_X1 U5977 ( .B1(n4934), .B2(n4933), .A(n5309), .ZN(n4948) );
  INV_X1 U5978 ( .A(n4935), .ZN(n4936) );
  AOI21_X1 U5979 ( .B1(n4937), .B2(n4680), .A(n4936), .ZN(n5605) );
  NAND2_X1 U5980 ( .A1(n5931), .A2(REIP_REG_15__SCAN_IN), .ZN(n4938) );
  OAI221_X1 U5981 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n4940), .C1(
        n6888), .C2(n4939), .A(n4938), .ZN(n4941) );
  AOI21_X1 U5982 ( .B1(n5605), .B2(n5927), .A(n4941), .ZN(n4942) );
  OAI21_X1 U5983 ( .B1(n4948), .B2(n5906), .A(n4942), .ZN(U3003) );
  XOR2_X1 U5984 ( .A(n4944), .B(n4943), .Z(n5604) );
  AOI22_X1 U5985 ( .A1(n5829), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n5931), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n4945) );
  OAI21_X1 U5986 ( .B1(n5856), .B2(n5602), .A(n4945), .ZN(n4946) );
  AOI21_X1 U5987 ( .B1(n5604), .B2(n5851), .A(n4946), .ZN(n4947) );
  OAI21_X1 U5988 ( .B1(n4948), .B2(n5814), .A(n4947), .ZN(U2971) );
  INV_X1 U5989 ( .A(n5517), .ZN(n4949) );
  NOR2_X1 U5990 ( .A1(n5515), .A2(n4949), .ZN(n4950) );
  XNOR2_X1 U5991 ( .A(n5516), .B(n4950), .ZN(n4963) );
  OR2_X1 U5992 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5548), .ZN(n5863)
         );
  AOI21_X1 U5993 ( .B1(n5860), .B2(n5863), .A(n4951), .ZN(n4955) );
  NOR3_X1 U5994 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n5548), .A3(n3605), 
        .ZN(n4954) );
  NAND2_X1 U5995 ( .A1(n5931), .A2(REIP_REG_12__SCAN_IN), .ZN(n4958) );
  OAI21_X1 U5996 ( .B1(n5903), .B2(n4952), .A(n4958), .ZN(n4953) );
  NOR3_X1 U5997 ( .A1(n4955), .A2(n4954), .A3(n4953), .ZN(n4956) );
  OAI21_X1 U5998 ( .B1(n4963), .B2(n5906), .A(n4956), .ZN(U3006) );
  NAND2_X1 U5999 ( .A1(n5829), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4957)
         );
  OAI211_X1 U6000 ( .C1(n5856), .C2(n4959), .A(n4958), .B(n4957), .ZN(n4960)
         );
  AOI21_X1 U6001 ( .B1(n4961), .B2(n5851), .A(n4960), .ZN(n4962) );
  OAI21_X1 U6002 ( .B1(n4963), .B2(n5814), .A(n4962), .ZN(U2974) );
  AOI22_X1 U6003 ( .A1(n4965), .A2(EAX_REG_31__SCAN_IN), .B1(n4964), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4966) );
  INV_X1 U6004 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6583) );
  INV_X1 U6005 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6582) );
  INV_X1 U6006 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6584) );
  NOR2_X1 U6007 ( .A1(n6582), .A2(n6584), .ZN(n4970) );
  NAND3_X1 U6008 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4973) );
  OAI21_X1 U6009 ( .B1(n4969), .B2(n4973), .A(n5473), .ZN(n5432) );
  OAI21_X1 U6010 ( .B1(n4970), .B2(n5667), .A(n5432), .ZN(n5046) );
  AOI21_X1 U6011 ( .B1(n5612), .B2(n6583), .A(n5046), .ZN(n5019) );
  OAI21_X1 U6012 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5667), .A(n5019), .ZN(n4980) );
  INV_X1 U6013 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4994) );
  NAND2_X1 U6014 ( .A1(n4972), .A2(n4971), .ZN(n4976) );
  INV_X1 U6015 ( .A(REIP_REG_31__SCAN_IN), .ZN(n4974) );
  NAND3_X1 U6016 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        n5460), .ZN(n5441) );
  NOR2_X1 U6017 ( .A1(n5441), .A2(n4973), .ZN(n5064) );
  NAND3_X1 U6018 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .A3(
        n5064), .ZN(n5031) );
  NOR2_X1 U6019 ( .A1(n6583), .A2(n5031), .ZN(n5022) );
  NAND3_X1 U6020 ( .A1(n4974), .A2(REIP_REG_30__SCAN_IN), .A3(n5022), .ZN(
        n4975) );
  OAI211_X1 U6021 ( .C1(n4994), .C2(n5718), .A(n4976), .B(n4975), .ZN(n4979)
         );
  NOR2_X1 U6022 ( .A1(n4977), .A2(n5711), .ZN(n4978) );
  OAI21_X1 U6023 ( .B1(n4968), .B2(n5479), .A(n4981), .ZN(U2796) );
  AND2_X1 U6024 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4987) );
  AOI21_X1 U6025 ( .B1(n4983), .B2(n4987), .A(n4982), .ZN(n4984) );
  XNOR2_X1 U6026 ( .A(n4984), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4985)
         );
  INV_X1 U6027 ( .A(n4985), .ZN(n5001) );
  OAI21_X1 U6028 ( .B1(n4987), .B2(n5868), .A(n4986), .ZN(n4990) );
  NAND3_X1 U6029 ( .A1(n5327), .A2(n4987), .A3(n4715), .ZN(n4988) );
  NAND2_X1 U6030 ( .A1(n5931), .A2(REIP_REG_31__SCAN_IN), .ZN(n4993) );
  OAI211_X1 U6031 ( .C1(n4977), .C2(n5903), .A(n4988), .B(n4993), .ZN(n4989)
         );
  AOI21_X1 U6032 ( .B1(n4990), .B2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n4989), 
        .ZN(n4991) );
  OAI21_X1 U6033 ( .B1(n5001), .B2(n5906), .A(n4991), .ZN(U2987) );
  INV_X1 U6034 ( .A(n4992), .ZN(n4998) );
  OAI21_X1 U6035 ( .B1(n5297), .B2(n4994), .A(n4993), .ZN(n4995) );
  INV_X1 U6036 ( .A(n4995), .ZN(n4997) );
  INV_X1 U6037 ( .A(n4999), .ZN(n5000) );
  OAI21_X1 U6038 ( .B1(n5001), .B2(n5814), .A(n5000), .ZN(U2955) );
  INV_X1 U6039 ( .A(n5209), .ZN(n5005) );
  AOI21_X1 U6040 ( .B1(n5829), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5002), 
        .ZN(n5003) );
  OAI21_X1 U6041 ( .B1(n5856), .B2(n5017), .A(n5003), .ZN(n5004) );
  AOI21_X1 U6042 ( .B1(n5005), .B2(n5851), .A(n5004), .ZN(n5006) );
  OAI21_X1 U6043 ( .B1(n5007), .B2(n5814), .A(n5006), .ZN(U2956) );
  OAI22_X1 U6044 ( .A1(n5010), .A2(n5549), .B1(n5009), .B2(n5008), .ZN(n5013)
         );
  AOI22_X1 U6045 ( .A1(n5554), .A2(n5013), .B1(n5012), .B2(n5011), .ZN(n5014)
         );
  OAI21_X1 U6046 ( .B1(n5016), .B2(n5015), .A(n5014), .ZN(U3456) );
  NOR2_X1 U6047 ( .A1(n5017), .A2(n5717), .ZN(n5021) );
  OAI22_X1 U6048 ( .A1(n5019), .A2(n3836), .B1(n5018), .B2(n5718), .ZN(n5020)
         );
  AOI211_X1 U6049 ( .C1(n3836), .C2(n5022), .A(n5021), .B(n5020), .ZN(n5023)
         );
  OAI21_X1 U6050 ( .B1(n5708), .B2(n5024), .A(n5023), .ZN(n5025) );
  AOI21_X1 U6051 ( .B1(n5026), .B2(n5687), .A(n5025), .ZN(n5027) );
  OAI21_X1 U6052 ( .B1(n5209), .B2(n5479), .A(n5027), .ZN(U2797) );
  INV_X1 U6053 ( .A(n5028), .ZN(n5040) );
  INV_X1 U6054 ( .A(n4890), .ZN(n5029) );
  INV_X1 U6055 ( .A(n5031), .ZN(n5033) );
  OAI22_X1 U6056 ( .A1(n5240), .A2(n5717), .B1(n3827), .B2(n5708), .ZN(n5032)
         );
  AOI21_X1 U6057 ( .B1(n6583), .B2(n5033), .A(n5032), .ZN(n5034) );
  OAI21_X1 U6058 ( .B1(n5718), .B2(n4885), .A(n5034), .ZN(n5037) );
  XNOR2_X1 U6059 ( .A(n5045), .B(n5035), .ZN(n5323) );
  NOR2_X1 U6060 ( .A1(n5323), .A2(n5711), .ZN(n5036) );
  AOI211_X1 U6061 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5046), .A(n5037), .B(n5036), .ZN(n5038) );
  OAI21_X1 U6062 ( .B1(n5238), .B2(n5479), .A(n5038), .ZN(U2798) );
  INV_X1 U6063 ( .A(n5039), .ZN(n5042) );
  INV_X1 U6064 ( .A(n5054), .ZN(n5041) );
  AOI21_X1 U6065 ( .B1(n5042), .B2(n5041), .A(n5040), .ZN(n5248) );
  INV_X1 U6066 ( .A(n5248), .ZN(n5214) );
  AND2_X1 U6067 ( .A1(n5060), .A2(n5043), .ZN(n5044) );
  NOR2_X1 U6068 ( .A1(n5045), .A2(n5044), .ZN(n5332) );
  INV_X1 U6069 ( .A(n5046), .ZN(n5049) );
  OAI22_X1 U6070 ( .A1(n6916), .A2(n5718), .B1(n5717), .B2(n5246), .ZN(n5047)
         );
  AOI21_X1 U6071 ( .B1(n5699), .B2(EBX_REG_28__SCAN_IN), .A(n5047), .ZN(n5048)
         );
  OAI21_X1 U6072 ( .B1(n5049), .B2(n6584), .A(n5048), .ZN(n5050) );
  AOI21_X1 U6073 ( .B1(n5332), .B2(n5687), .A(n5050), .ZN(n5052) );
  NAND3_X1 U6074 ( .A1(n5064), .A2(REIP_REG_27__SCAN_IN), .A3(n6584), .ZN(
        n5051) );
  OAI211_X1 U6075 ( .C1(n5214), .C2(n5479), .A(n5052), .B(n5051), .ZN(U2799)
         );
  AOI21_X1 U6076 ( .B1(n5055), .B2(n5053), .A(n5054), .ZN(n5256) );
  INV_X1 U6077 ( .A(n5256), .ZN(n5217) );
  AOI22_X1 U6078 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n5696), .B1(
        EBX_REG_27__SCAN_IN), .B2(n5699), .ZN(n5056) );
  OAI21_X1 U6079 ( .B1(n6582), .B2(n5432), .A(n5056), .ZN(n5063) );
  NAND2_X1 U6080 ( .A1(n5057), .A2(n5058), .ZN(n5059) );
  NAND2_X1 U6081 ( .A1(n5060), .A2(n5059), .ZN(n5338) );
  INV_X1 U6082 ( .A(n5061), .ZN(n5254) );
  OAI22_X1 U6083 ( .A1(n5338), .A2(n5711), .B1(n5254), .B2(n5717), .ZN(n5062)
         );
  AOI211_X1 U6084 ( .C1(n5064), .C2(n6582), .A(n5063), .B(n5062), .ZN(n5065)
         );
  OAI21_X1 U6085 ( .B1(n5217), .B2(n5479), .A(n5065), .ZN(U2800) );
  INV_X1 U6086 ( .A(n5473), .ZN(n5709) );
  NOR2_X1 U6087 ( .A1(n5709), .A2(n5456), .ZN(n5467) );
  NOR2_X1 U6088 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5455), .ZN(n5069) );
  OAI22_X1 U6089 ( .A1(n5288), .A2(n5718), .B1(n5067), .B2(n5708), .ZN(n5068)
         );
  AOI211_X1 U6090 ( .C1(n5467), .C2(REIP_REG_21__SCAN_IN), .A(n5069), .B(n5068), .ZN(n5075) );
  OR2_X1 U6091 ( .A1(n5072), .A2(n5071), .ZN(n5073) );
  AND2_X1 U6092 ( .A1(n5070), .A2(n5073), .ZN(n5394) );
  AOI22_X1 U6093 ( .A1(n5394), .A2(n5687), .B1(n5654), .B2(n5290), .ZN(n5074)
         );
  OAI211_X1 U6094 ( .C1(n5499), .C2(n5479), .A(n5075), .B(n5074), .ZN(U2806)
         );
  OAI21_X1 U6095 ( .B1(n5195), .B2(n5077), .A(n5271), .ZN(n5228) );
  INV_X1 U6096 ( .A(n5228), .ZN(n5315) );
  INV_X1 U6097 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5078) );
  OAI22_X1 U6098 ( .A1(n5078), .A2(n5718), .B1(n6953), .B2(n5708), .ZN(n5088)
         );
  OAI21_X1 U6099 ( .B1(n5081), .B2(n5080), .A(n5079), .ZN(n5193) );
  INV_X1 U6100 ( .A(n5313), .ZN(n5082) );
  AOI21_X1 U6101 ( .B1(n5654), .B2(n5082), .A(n5695), .ZN(n5086) );
  OAI21_X1 U6102 ( .B1(n5667), .B2(n5083), .A(n6570), .ZN(n5084) );
  NAND3_X1 U6103 ( .A1(n5084), .A2(n5474), .A3(n5473), .ZN(n5085) );
  OAI211_X1 U6104 ( .C1(n5711), .C2(n5193), .A(n5086), .B(n5085), .ZN(n5087)
         );
  AOI211_X1 U6105 ( .C1(n5315), .C2(n5679), .A(n5088), .B(n5087), .ZN(n5089)
         );
  INV_X1 U6106 ( .A(n5089), .ZN(U2810) );
  INV_X1 U6107 ( .A(n5809), .ZN(n5091) );
  AOI22_X1 U6108 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n5696), .B1(n5687), 
        .B2(n5858), .ZN(n5090) );
  INV_X1 U6109 ( .A(n5695), .ZN(n5661) );
  OAI211_X1 U6110 ( .C1(n5717), .C2(n5091), .A(n5090), .B(n5661), .ZN(n5092)
         );
  AOI21_X1 U6111 ( .B1(n5699), .B2(EBX_REG_11__SCAN_IN), .A(n5092), .ZN(n5096)
         );
  INV_X1 U6112 ( .A(n5117), .ZN(n5093) );
  NOR2_X1 U6113 ( .A1(n5667), .A2(n5093), .ZN(n5688) );
  NAND3_X1 U6114 ( .A1(REIP_REG_8__SCAN_IN), .A2(n5648), .A3(n5688), .ZN(n5647) );
  OAI21_X1 U6115 ( .B1(n5104), .B2(n5647), .A(n6906), .ZN(n5094) );
  NAND2_X1 U6116 ( .A1(n5094), .A2(n5632), .ZN(n5095) );
  OAI211_X1 U6117 ( .C1(n5097), .C2(n5479), .A(n5096), .B(n5095), .ZN(U2816)
         );
  INV_X1 U6118 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6969) );
  AOI21_X1 U6119 ( .B1(n4645), .B2(n6969), .A(n5647), .ZN(n5105) );
  AOI21_X1 U6120 ( .B1(n5696), .B2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5695), 
        .ZN(n5098) );
  OAI21_X1 U6121 ( .B1(n5717), .B2(n5099), .A(n5098), .ZN(n5103) );
  OAI21_X1 U6122 ( .B1(n5137), .B2(n5100), .A(n5473), .ZN(n5658) );
  AOI22_X1 U6123 ( .A1(EBX_REG_10__SCAN_IN), .A2(n5699), .B1(n5687), .B2(n5866), .ZN(n5101) );
  OAI21_X1 U6124 ( .B1(n4645), .B2(n5658), .A(n5101), .ZN(n5102) );
  AOI211_X1 U6125 ( .C1(n5105), .C2(n5104), .A(n5103), .B(n5102), .ZN(n5106)
         );
  OAI21_X1 U6126 ( .B1(n5107), .B2(n5479), .A(n5106), .ZN(U2817) );
  OAI21_X1 U6127 ( .B1(n5112), .B2(n5108), .A(n5479), .ZN(n5714) );
  INV_X1 U6128 ( .A(n5714), .ZN(n5136) );
  NAND2_X1 U6129 ( .A1(n5699), .A2(EBX_REG_3__SCAN_IN), .ZN(n5115) );
  INV_X1 U6130 ( .A(n5109), .ZN(n5110) );
  AOI22_X1 U6131 ( .A1(n5110), .A2(n5654), .B1(n5696), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5114) );
  NOR2_X1 U6132 ( .A1(n5112), .A2(n5111), .ZN(n5706) );
  NAND2_X1 U6133 ( .A1(n5706), .A2(n6270), .ZN(n5113) );
  NAND3_X1 U6134 ( .A1(n5115), .A2(n5114), .A3(n5113), .ZN(n5121) );
  INV_X1 U6135 ( .A(REIP_REG_3__SCAN_IN), .ZN(n5119) );
  OAI21_X1 U6136 ( .B1(n5137), .B2(n6601), .A(n5473), .ZN(n5116) );
  NAND2_X1 U6137 ( .A1(n5116), .A2(REIP_REG_2__SCAN_IN), .ZN(n5132) );
  OR2_X1 U6138 ( .A1(n5667), .A2(n5117), .ZN(n5118) );
  NAND2_X1 U6139 ( .A1(n5118), .A2(n5591), .ZN(n5700) );
  INV_X1 U6140 ( .A(n5700), .ZN(n5666) );
  AOI21_X1 U6141 ( .B1(n5119), .B2(n5132), .A(n5666), .ZN(n5120) );
  AOI211_X1 U6142 ( .C1(n5917), .C2(n5687), .A(n5121), .B(n5120), .ZN(n5122)
         );
  OAI21_X1 U6143 ( .B1(n5136), .B2(n5123), .A(n5122), .ZN(U2824) );
  NAND2_X1 U6144 ( .A1(n5706), .A2(n6152), .ZN(n5126) );
  INV_X1 U6145 ( .A(n5855), .ZN(n5124) );
  NAND2_X1 U6146 ( .A1(n5654), .A2(n5124), .ZN(n5125) );
  OAI211_X1 U6147 ( .C1(n5127), .C2(n5718), .A(n5126), .B(n5125), .ZN(n5131)
         );
  XNOR2_X1 U6148 ( .A(n5129), .B(n5128), .ZN(n5729) );
  NOR2_X1 U6149 ( .A1(n5711), .A2(n5729), .ZN(n5130) );
  AOI211_X1 U6150 ( .C1(n5699), .C2(EBX_REG_2__SCAN_IN), .A(n5131), .B(n5130), 
        .ZN(n5135) );
  AND2_X1 U6151 ( .A1(n5612), .A2(REIP_REG_1__SCAN_IN), .ZN(n5133) );
  OAI21_X1 U6152 ( .B1(n5133), .B2(REIP_REG_2__SCAN_IN), .A(n5132), .ZN(n5134)
         );
  OAI211_X1 U6153 ( .C1(n5136), .C2(n5728), .A(n5135), .B(n5134), .ZN(U2825)
         );
  AOI22_X1 U6154 ( .A1(EBX_REG_1__SCAN_IN), .A2(n5699), .B1(n5137), .B2(
        REIP_REG_1__SCAN_IN), .ZN(n5146) );
  AOI22_X1 U6155 ( .A1(n5696), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5654), 
        .B2(n5138), .ZN(n5140) );
  NAND2_X1 U6156 ( .A1(n5706), .A2(n6151), .ZN(n5139) );
  OAI211_X1 U6157 ( .C1(REIP_REG_1__SCAN_IN), .C2(n5667), .A(n5140), .B(n5139), 
        .ZN(n5141) );
  INV_X1 U6158 ( .A(n5141), .ZN(n5145) );
  AOI22_X1 U6159 ( .A1(n5687), .A2(n5143), .B1(n5142), .B2(n5714), .ZN(n5144)
         );
  NAND3_X1 U6160 ( .A1(n5146), .A2(n5145), .A3(n5144), .ZN(U2826) );
  OAI222_X1 U6161 ( .A1(n5238), .A2(n5203), .B1(n3827), .B2(n5733), .C1(n5720), 
        .C2(n5323), .ZN(U2830) );
  AOI22_X1 U6162 ( .A1(n5332), .A2(n5730), .B1(EBX_REG_28__SCAN_IN), .B2(n5201), .ZN(n5147) );
  OAI21_X1 U6163 ( .B1(n5214), .B2(n5203), .A(n5147), .ZN(U2831) );
  INV_X1 U6164 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5148) );
  OAI222_X1 U6165 ( .A1(n5203), .A2(n5217), .B1(n5148), .B2(n5733), .C1(n5338), 
        .C2(n5720), .ZN(U2832) );
  NAND2_X1 U6166 ( .A1(n5195), .A2(n5149), .ZN(n5151) );
  NAND2_X1 U6167 ( .A1(n5151), .A2(n5150), .ZN(n5152) );
  AND2_X1 U6168 ( .A1(n5053), .A2(n5152), .ZN(n5435) );
  INV_X1 U6169 ( .A(n5435), .ZN(n5220) );
  OR2_X1 U6170 ( .A1(n5358), .A2(n5153), .ZN(n5154) );
  NAND2_X1 U6171 ( .A1(n5057), .A2(n5154), .ZN(n5431) );
  OAI222_X1 U6172 ( .A1(n5203), .A2(n5220), .B1(n5733), .B2(n3815), .C1(n5431), 
        .C2(n5720), .ZN(U2833) );
  AND2_X1 U6173 ( .A1(n5156), .A2(n5155), .ZN(n5157) );
  OR2_X1 U6174 ( .A1(n5157), .A2(n5357), .ZN(n5454) );
  INV_X1 U6175 ( .A(n5493), .ZN(n5160) );
  OAI222_X1 U6176 ( .A1(n5720), .A2(n5454), .B1(n5733), .B2(n3807), .C1(n5203), 
        .C2(n5160), .ZN(U2835) );
  AOI22_X1 U6177 ( .A1(n5376), .A2(n5730), .B1(EBX_REG_23__SCAN_IN), .B2(n5201), .ZN(n5161) );
  OAI21_X1 U6178 ( .B1(n5223), .B2(n5203), .A(n5161), .ZN(U2836) );
  INV_X1 U6179 ( .A(n5162), .ZN(n5496) );
  INV_X1 U6180 ( .A(n5203), .ZN(n5731) );
  NAND2_X1 U6181 ( .A1(n5070), .A2(n5163), .ZN(n5164) );
  NAND2_X1 U6182 ( .A1(n5165), .A2(n5164), .ZN(n5464) );
  OAI22_X1 U6183 ( .A1(n5464), .A2(n5720), .B1(n6796), .B2(n5733), .ZN(n5166)
         );
  AOI21_X1 U6184 ( .B1(n5496), .B2(n5731), .A(n5166), .ZN(n5167) );
  INV_X1 U6185 ( .A(n5167), .ZN(U2837) );
  AOI22_X1 U6186 ( .A1(n5394), .A2(n5730), .B1(EBX_REG_21__SCAN_IN), .B2(n5201), .ZN(n5168) );
  OAI21_X1 U6187 ( .B1(n5499), .B2(n5203), .A(n5168), .ZN(U2838) );
  INV_X1 U6188 ( .A(n5182), .ZN(n5171) );
  MUX2_X1 U6189 ( .A(n5171), .B(n3188), .S(n5169), .Z(n5173) );
  XNOR2_X1 U6190 ( .A(n5173), .B(n5172), .ZN(n5469) );
  NOR2_X1 U6191 ( .A1(n5179), .A2(n5174), .ZN(n5175) );
  OAI222_X1 U6192 ( .A1(n5720), .A2(n5469), .B1(n5177), .B2(n5733), .C1(n5468), 
        .C2(n5203), .ZN(U2839) );
  AND2_X1 U6193 ( .A1(n5191), .A2(n5178), .ZN(n5180) );
  OR2_X1 U6194 ( .A1(n5180), .A2(n5179), .ZN(n5480) );
  INV_X1 U6195 ( .A(n5480), .ZN(n5299) );
  XNOR2_X1 U6196 ( .A(n5182), .B(n5181), .ZN(n5186) );
  OR2_X1 U6197 ( .A1(n5079), .A2(n5186), .ZN(n5188) );
  XNOR2_X1 U6198 ( .A(n5188), .B(n5183), .ZN(n5478) );
  OAI22_X1 U6199 ( .A1(n5478), .A2(n5720), .B1(n5485), .B2(n5733), .ZN(n5184)
         );
  AOI21_X1 U6200 ( .B1(n5299), .B2(n5731), .A(n5184), .ZN(n5185) );
  INV_X1 U6201 ( .A(n5185), .ZN(U2840) );
  NAND2_X1 U6202 ( .A1(n5079), .A2(n5186), .ZN(n5187) );
  AND2_X1 U6203 ( .A1(n5188), .A2(n5187), .ZN(n5583) );
  INV_X1 U6204 ( .A(n5583), .ZN(n5523) );
  INV_X1 U6205 ( .A(EBX_REG_18__SCAN_IN), .ZN(n6812) );
  NAND2_X1 U6206 ( .A1(n5271), .A2(n5189), .ZN(n5190) );
  INV_X1 U6207 ( .A(n5734), .ZN(n5192) );
  OAI222_X1 U6208 ( .A1(n5523), .A2(n5720), .B1(n5733), .B2(n6812), .C1(n5192), 
        .C2(n5203), .ZN(U2841) );
  INV_X1 U6209 ( .A(n5193), .ZN(n5530) );
  AOI22_X1 U6210 ( .A1(n5530), .A2(n5730), .B1(EBX_REG_17__SCAN_IN), .B2(n5201), .ZN(n5194) );
  OAI21_X1 U6211 ( .B1(n5228), .B2(n5203), .A(n5194), .ZN(U2842) );
  AOI21_X1 U6212 ( .B1(n5197), .B2(n5196), .A(n5195), .ZN(n5739) );
  INV_X1 U6213 ( .A(n5739), .ZN(n5200) );
  INV_X1 U6214 ( .A(n5600), .ZN(n5198) );
  AOI22_X1 U6215 ( .A1(n5198), .A2(n5730), .B1(EBX_REG_16__SCAN_IN), .B2(n5201), .ZN(n5199) );
  OAI21_X1 U6216 ( .B1(n5200), .B2(n5203), .A(n5199), .ZN(U2843) );
  INV_X1 U6217 ( .A(n5604), .ZN(n5231) );
  AOI22_X1 U6218 ( .A1(n5605), .A2(n5730), .B1(EBX_REG_15__SCAN_IN), .B2(n5201), .ZN(n5202) );
  OAI21_X1 U6219 ( .B1(n5231), .B2(n5203), .A(n5202), .ZN(U2844) );
  NAND2_X1 U6220 ( .A1(n5204), .A2(n5987), .ZN(n5206) );
  AOI22_X1 U6221 ( .A1(n5737), .A2(DATAI_31_), .B1(n5740), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5205) );
  OAI21_X1 U6222 ( .B1(n4968), .B2(n5206), .A(n5205), .ZN(U2860) );
  AOI22_X1 U6223 ( .A1(n5737), .A2(DATAI_30_), .B1(n5740), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5208) );
  NAND2_X1 U6224 ( .A1(n5741), .A2(DATAI_14_), .ZN(n5207) );
  OAI211_X1 U6225 ( .C1(n5209), .C2(n5489), .A(n5208), .B(n5207), .ZN(U2861)
         );
  AOI22_X1 U6226 ( .A1(n5737), .A2(DATAI_29_), .B1(n5740), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6227 ( .A1(n5741), .A2(DATAI_13_), .ZN(n5210) );
  OAI211_X1 U6228 ( .C1(n5238), .C2(n5489), .A(n5211), .B(n5210), .ZN(U2862)
         );
  AOI22_X1 U6229 ( .A1(n5737), .A2(DATAI_28_), .B1(n5740), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6230 ( .A1(n5741), .A2(DATAI_12_), .ZN(n5212) );
  OAI211_X1 U6231 ( .C1(n5214), .C2(n5489), .A(n5213), .B(n5212), .ZN(U2863)
         );
  AOI22_X1 U6232 ( .A1(n5737), .A2(DATAI_27_), .B1(n5740), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6233 ( .A1(n5741), .A2(DATAI_11_), .ZN(n5215) );
  OAI211_X1 U6234 ( .C1(n5217), .C2(n5489), .A(n5216), .B(n5215), .ZN(U2864)
         );
  AOI22_X1 U6235 ( .A1(n5737), .A2(DATAI_26_), .B1(n5740), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5219) );
  NAND2_X1 U6236 ( .A1(n5741), .A2(DATAI_10_), .ZN(n5218) );
  OAI211_X1 U6237 ( .C1(n5220), .C2(n5489), .A(n5219), .B(n5218), .ZN(U2865)
         );
  AOI22_X1 U6238 ( .A1(n5737), .A2(DATAI_23_), .B1(n5740), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U6239 ( .A1(n5741), .A2(DATAI_7_), .ZN(n5221) );
  OAI211_X1 U6240 ( .C1(n5223), .C2(n5489), .A(n5222), .B(n5221), .ZN(U2868)
         );
  AOI22_X1 U6241 ( .A1(n5737), .A2(DATAI_19_), .B1(n5740), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6242 ( .A1(n5741), .A2(DATAI_3_), .ZN(n5224) );
  OAI211_X1 U6243 ( .C1(n5480), .C2(n5489), .A(n5225), .B(n5224), .ZN(U2872)
         );
  AOI22_X1 U6244 ( .A1(n5737), .A2(DATAI_17_), .B1(n5740), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6245 ( .A1(n5741), .A2(DATAI_1_), .ZN(n5226) );
  OAI211_X1 U6246 ( .C1(n5228), .C2(n5489), .A(n5227), .B(n5226), .ZN(U2874)
         );
  AOI22_X1 U6247 ( .A1(n5229), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n5740), .ZN(n5230) );
  OAI21_X1 U6248 ( .B1(n5231), .B2(n5489), .A(n5230), .ZN(U2876) );
  INV_X1 U6249 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5232) );
  NOR2_X1 U6250 ( .A1(n5251), .A2(n5232), .ZN(n5234) );
  OR2_X1 U6251 ( .A1(n5234), .A2(n5233), .ZN(n5244) );
  OAI21_X1 U6252 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5235), .ZN(n5334) );
  NAND2_X1 U6253 ( .A1(n5244), .A2(n5334), .ZN(n5237) );
  XNOR2_X1 U6254 ( .A(n5237), .B(n5236), .ZN(n5330) );
  INV_X1 U6255 ( .A(n5238), .ZN(n5242) );
  NOR2_X1 U6256 ( .A1(n5912), .A2(n6583), .ZN(n5324) );
  AOI21_X1 U6257 ( .B1(n5829), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5324), 
        .ZN(n5239) );
  OAI21_X1 U6258 ( .B1(n5856), .B2(n5240), .A(n5239), .ZN(n5241) );
  AOI21_X1 U6259 ( .B1(n5242), .B2(n5851), .A(n5241), .ZN(n5243) );
  OAI21_X1 U6260 ( .B1(n5814), .B2(n5330), .A(n5243), .ZN(U2957) );
  XNOR2_X1 U6261 ( .A(n5244), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5337)
         );
  NOR2_X1 U6262 ( .A1(n5912), .A2(n6584), .ZN(n5331) );
  AOI21_X1 U6263 ( .B1(n5829), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5331), 
        .ZN(n5245) );
  OAI21_X1 U6264 ( .B1(n5856), .B2(n5246), .A(n5245), .ZN(n5247) );
  AOI21_X1 U6265 ( .B1(n5248), .B2(n5851), .A(n5247), .ZN(n5249) );
  OAI21_X1 U6266 ( .B1(n5337), .B2(n5814), .A(n5249), .ZN(U2958) );
  NAND2_X1 U6267 ( .A1(n5251), .A2(n5250), .ZN(n5252) );
  XNOR2_X1 U6268 ( .A(n5252), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5346)
         );
  NOR2_X1 U6269 ( .A1(n5912), .A2(n6582), .ZN(n5339) );
  AOI21_X1 U6270 ( .B1(n5829), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5339), 
        .ZN(n5253) );
  OAI21_X1 U6271 ( .B1(n5856), .B2(n5254), .A(n5253), .ZN(n5255) );
  AOI21_X1 U6272 ( .B1(n5256), .B2(n5851), .A(n5255), .ZN(n5257) );
  OAI21_X1 U6273 ( .B1(n5346), .B2(n5814), .A(n5257), .ZN(U2959) );
  XNOR2_X1 U6274 ( .A(n3620), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5258)
         );
  XNOR2_X1 U6275 ( .A(n5259), .B(n5258), .ZN(n5354) );
  INV_X1 U6276 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5260) );
  NOR2_X1 U6277 ( .A1(n5912), .A2(n5260), .ZN(n5349) );
  AOI21_X1 U6278 ( .B1(n5829), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5349), 
        .ZN(n5261) );
  OAI21_X1 U6279 ( .B1(n5856), .B2(n5438), .A(n5261), .ZN(n5262) );
  AOI21_X1 U6280 ( .B1(n5435), .B2(n5851), .A(n5262), .ZN(n5263) );
  OAI21_X1 U6281 ( .B1(n5814), .B2(n5354), .A(n5263), .ZN(U2960) );
  INV_X1 U6282 ( .A(n5264), .ZN(n5265) );
  AOI21_X1 U6283 ( .B1(n5267), .B2(n5266), .A(n5265), .ZN(n5367) );
  INV_X1 U6284 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5268) );
  NOR2_X1 U6285 ( .A1(n5912), .A2(n5268), .ZN(n5361) );
  NOR2_X1 U6286 ( .A1(n5297), .A2(n5269), .ZN(n5270) );
  AOI211_X1 U6287 ( .C1(n5810), .C2(n5440), .A(n5361), .B(n5270), .ZN(n5277)
         );
  INV_X1 U6288 ( .A(n5271), .ZN(n5273) );
  XNOR2_X1 U6289 ( .A(n5275), .B(n5274), .ZN(n5490) );
  NAND2_X1 U6290 ( .A1(n5490), .A2(n5851), .ZN(n5276) );
  OAI211_X1 U6291 ( .C1(n5367), .C2(n5814), .A(n5277), .B(n5276), .ZN(U2961)
         );
  NAND3_X1 U6292 ( .A1(n5304), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5278) );
  XNOR2_X1 U6293 ( .A(n5281), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5374)
         );
  NOR2_X1 U6294 ( .A1(n5912), .A2(n6578), .ZN(n5371) );
  NOR2_X1 U6295 ( .A1(n5297), .A2(n5448), .ZN(n5282) );
  AOI211_X1 U6296 ( .C1(n5810), .C2(n5451), .A(n5371), .B(n5282), .ZN(n5284)
         );
  NAND2_X1 U6297 ( .A1(n5493), .A2(n5851), .ZN(n5283) );
  OAI211_X1 U6298 ( .C1(n5374), .C2(n5814), .A(n5284), .B(n5283), .ZN(U2962)
         );
  OAI21_X1 U6299 ( .B1(n5287), .B2(n5286), .A(n5285), .ZN(n5400) );
  NAND2_X1 U6300 ( .A1(n5400), .A2(n5850), .ZN(n5292) );
  NOR2_X1 U6301 ( .A1(n5912), .A2(n6576), .ZN(n5393) );
  NOR2_X1 U6302 ( .A1(n5297), .A2(n5288), .ZN(n5289) );
  AOI211_X1 U6303 ( .C1(n5810), .C2(n5290), .A(n5393), .B(n5289), .ZN(n5291)
         );
  OAI211_X1 U6304 ( .C1(n6457), .C2(n5499), .A(n5292), .B(n5291), .ZN(U2965)
         );
  XOR2_X1 U6305 ( .A(n5295), .B(n5294), .Z(n5423) );
  NOR2_X1 U6306 ( .A1(n5912), .A2(n6571), .ZN(n5416) );
  NOR2_X1 U6307 ( .A1(n5297), .A2(n5296), .ZN(n5298) );
  AOI211_X1 U6308 ( .C1(n5810), .C2(n5482), .A(n5416), .B(n5298), .ZN(n5301)
         );
  NAND2_X1 U6309 ( .A1(n5299), .A2(n5851), .ZN(n5300) );
  OAI211_X1 U6310 ( .C1(n5423), .C2(n5814), .A(n5301), .B(n5300), .ZN(U2967)
         );
  NAND3_X1 U6311 ( .A1(n5307), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5304), .ZN(n5511) );
  INV_X1 U6312 ( .A(n5511), .ZN(n5311) );
  NAND2_X1 U6313 ( .A1(n3620), .A2(n5534), .ZN(n5306) );
  AOI22_X1 U6314 ( .A1(n5307), .A2(n5306), .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5305), .ZN(n5310) );
  NAND3_X1 U6315 ( .A1(n5309), .A2(n5308), .A3(n5534), .ZN(n5510) );
  OAI21_X1 U6316 ( .B1(n5311), .B2(n5310), .A(n5510), .ZN(n5531) );
  INV_X1 U6317 ( .A(n5531), .ZN(n5317) );
  AOI22_X1 U6318 ( .A1(n5829), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .B1(n5931), 
        .B2(REIP_REG_17__SCAN_IN), .ZN(n5312) );
  OAI21_X1 U6319 ( .B1(n5856), .B2(n5313), .A(n5312), .ZN(n5314) );
  AOI21_X1 U6320 ( .B1(n5315), .B2(n5851), .A(n5314), .ZN(n5316) );
  OAI21_X1 U6321 ( .B1(n5317), .B2(n5814), .A(n5316), .ZN(U2969) );
  AND2_X1 U6322 ( .A1(n5829), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5318)
         );
  AOI211_X1 U6323 ( .C1(n5597), .C2(n5810), .A(n5319), .B(n5318), .ZN(n5321)
         );
  NAND2_X1 U6324 ( .A1(n5739), .A2(n5851), .ZN(n5320) );
  OAI211_X1 U6325 ( .C1(n5322), .C2(n5814), .A(n5321), .B(n5320), .ZN(U2970)
         );
  INV_X1 U6326 ( .A(n5323), .ZN(n5325) );
  AOI21_X1 U6327 ( .B1(n5325), .B2(n5927), .A(n5324), .ZN(n5329) );
  OAI21_X1 U6328 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5327), .A(n5326), 
        .ZN(n5328) );
  OAI211_X1 U6329 ( .C1(n5330), .C2(n5906), .A(n5329), .B(n5328), .ZN(U2989)
         );
  AOI21_X1 U6330 ( .B1(n5332), .B2(n5927), .A(n5331), .ZN(n5333) );
  OAI21_X1 U6331 ( .B1(n5342), .B2(n5334), .A(n5333), .ZN(n5335) );
  AOI21_X1 U6332 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n5344), .A(n5335), 
        .ZN(n5336) );
  OAI21_X1 U6333 ( .B1(n5337), .B2(n5906), .A(n5336), .ZN(U2990) );
  INV_X1 U6334 ( .A(n5338), .ZN(n5340) );
  AOI21_X1 U6335 ( .B1(n5340), .B2(n5927), .A(n5339), .ZN(n5341) );
  OAI21_X1 U6336 ( .B1(n5342), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5341), 
        .ZN(n5343) );
  AOI21_X1 U6337 ( .B1(n5344), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5343), 
        .ZN(n5345) );
  OAI21_X1 U6338 ( .B1(n5346), .B2(n5906), .A(n5345), .ZN(U2991) );
  INV_X1 U6339 ( .A(n5368), .ZN(n5365) );
  INV_X1 U6340 ( .A(n5347), .ZN(n5348) );
  OAI211_X1 U6341 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5355), .B(n5348), .ZN(n5351) );
  INV_X1 U6342 ( .A(n5349), .ZN(n5350) );
  OAI211_X1 U6343 ( .C1(n5903), .C2(n5431), .A(n5351), .B(n5350), .ZN(n5352)
         );
  AOI21_X1 U6344 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5365), .A(n5352), 
        .ZN(n5353) );
  OAI21_X1 U6345 ( .B1(n5354), .B2(n5906), .A(n5353), .ZN(U2992) );
  INV_X1 U6346 ( .A(n5355), .ZN(n5363) );
  INV_X1 U6347 ( .A(n5356), .ZN(n5360) );
  INV_X1 U6348 ( .A(n5357), .ZN(n5359) );
  AOI21_X1 U6349 ( .B1(n5360), .B2(n5359), .A(n5358), .ZN(n5486) );
  AOI21_X1 U6350 ( .B1(n5486), .B2(n5927), .A(n5361), .ZN(n5362) );
  OAI21_X1 U6351 ( .B1(n5363), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5362), 
        .ZN(n5364) );
  AOI21_X1 U6352 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5365), .A(n5364), 
        .ZN(n5366) );
  OAI21_X1 U6353 ( .B1(n5367), .B2(n5906), .A(n5366), .ZN(U2993) );
  INV_X1 U6354 ( .A(n5454), .ZN(n5372) );
  NAND3_X1 U6355 ( .A1(n5419), .A2(n5377), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5369) );
  AOI21_X1 U6356 ( .B1(n6924), .B2(n5369), .A(n5368), .ZN(n5370) );
  AOI211_X1 U6357 ( .C1(n5927), .C2(n5372), .A(n5371), .B(n5370), .ZN(n5373)
         );
  OAI21_X1 U6358 ( .B1(n5374), .B2(n5906), .A(n5373), .ZN(U2994) );
  AOI21_X1 U6359 ( .B1(n5376), .B2(n5927), .A(n5375), .ZN(n5379) );
  NAND3_X1 U6360 ( .A1(n5419), .A2(n5377), .A3(n4747), .ZN(n5378) );
  OAI211_X1 U6361 ( .C1(n5380), .C2(n4747), .A(n5379), .B(n5378), .ZN(n5381)
         );
  AOI21_X1 U6362 ( .B1(n5382), .B2(n5929), .A(n5381), .ZN(n5383) );
  INV_X1 U6363 ( .A(n5383), .ZN(U2995) );
  NOR2_X1 U6364 ( .A1(n5408), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5384)
         );
  NAND2_X1 U6365 ( .A1(n5419), .A2(n5384), .ZN(n5396) );
  AOI21_X1 U6366 ( .B1(n5396), .B2(n5398), .A(n5385), .ZN(n5390) );
  NAND4_X1 U6367 ( .A1(n5419), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n5386), .A4(n5385), .ZN(n5388) );
  OAI211_X1 U6368 ( .C1(n5903), .C2(n5464), .A(n5388), .B(n5387), .ZN(n5389)
         );
  AOI211_X1 U6369 ( .C1(n5391), .C2(n5929), .A(n5390), .B(n5389), .ZN(n5392)
         );
  INV_X1 U6370 ( .A(n5392), .ZN(U2996) );
  AOI21_X1 U6371 ( .B1(n5394), .B2(n5927), .A(n5393), .ZN(n5395) );
  OAI211_X1 U6372 ( .C1(n5398), .C2(n5397), .A(n5396), .B(n5395), .ZN(n5399)
         );
  AOI21_X1 U6373 ( .B1(n5400), .B2(n5929), .A(n5399), .ZN(n5401) );
  INV_X1 U6374 ( .A(n5401), .ZN(U2997) );
  XNOR2_X1 U6375 ( .A(n5806), .B(n5402), .ZN(n5403) );
  XNOR2_X1 U6376 ( .A(n5404), .B(n5403), .ZN(n5506) );
  INV_X1 U6377 ( .A(n5506), .ZN(n5415) );
  NOR2_X1 U6378 ( .A1(n5405), .A2(n5534), .ZN(n5407) );
  OAI21_X1 U6379 ( .B1(n5407), .B2(n5897), .A(n5406), .ZN(n5533) );
  AOI21_X1 U6380 ( .B1(n5933), .B2(n5534), .A(n5533), .ZN(n5524) );
  OAI21_X1 U6381 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5868), .A(n5524), 
        .ZN(n5420) );
  AND2_X1 U6382 ( .A1(n5408), .A2(n5419), .ZN(n5411) );
  INV_X1 U6383 ( .A(n5409), .ZN(n5410) );
  AOI22_X1 U6384 ( .A1(n5931), .A2(REIP_REG_20__SCAN_IN), .B1(n5411), .B2(
        n5410), .ZN(n5412) );
  OAI21_X1 U6385 ( .B1(n5469), .B2(n5903), .A(n5412), .ZN(n5413) );
  AOI21_X1 U6386 ( .B1(n5420), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5413), 
        .ZN(n5414) );
  OAI21_X1 U6387 ( .B1(n5415), .B2(n5906), .A(n5414), .ZN(U2998) );
  NOR2_X1 U6388 ( .A1(n5478), .A2(n5903), .ZN(n5417) );
  AOI211_X1 U6389 ( .C1(n5419), .C2(n5418), .A(n5417), .B(n5416), .ZN(n5422)
         );
  NAND2_X1 U6390 ( .A1(n5420), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5421) );
  OAI211_X1 U6391 ( .C1(n5423), .C2(n5906), .A(n5422), .B(n5421), .ZN(U2999)
         );
  INV_X1 U6392 ( .A(n6217), .ZN(n5429) );
  NOR2_X1 U6393 ( .A1(n6216), .A2(n5424), .ZN(n6459) );
  NOR4_X1 U6394 ( .A1(n6459), .A2(n6302), .A3(n6454), .A4(n6216), .ZN(n5425)
         );
  AOI21_X1 U6395 ( .B1(n5426), .B2(n6270), .A(n5425), .ZN(n5427) );
  OAI21_X1 U6396 ( .B1(n5429), .B2(n5428), .A(n5427), .ZN(n5430) );
  MUX2_X1 U6397 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5430), .S(n5938), 
        .Z(U3462) );
  AND2_X1 U6398 ( .A1(n5775), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6399 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n5696), .B1(
        EBX_REG_26__SCAN_IN), .B2(n5699), .ZN(n5437) );
  INV_X1 U6400 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6578) );
  NOR2_X1 U6401 ( .A1(n6578), .A2(n5441), .ZN(n5439) );
  AOI21_X1 U6402 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5439), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5433) );
  OAI22_X1 U6403 ( .A1(n5433), .A2(n5432), .B1(n5431), .B2(n5711), .ZN(n5434)
         );
  AOI21_X1 U6404 ( .B1(n5435), .B2(n5679), .A(n5434), .ZN(n5436) );
  OAI211_X1 U6405 ( .C1(n5438), .C2(n5717), .A(n5437), .B(n5436), .ZN(U2801)
         );
  AOI22_X1 U6406 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n5696), .B1(
        EBX_REG_25__SCAN_IN), .B2(n5699), .ZN(n5446) );
  AOI22_X1 U6407 ( .A1(n5440), .A2(n5654), .B1(n5439), .B2(n5268), .ZN(n5445)
         );
  AOI22_X1 U6408 ( .A1(n5490), .A2(n5679), .B1(n5687), .B2(n5486), .ZN(n5444)
         );
  INV_X1 U6409 ( .A(n5447), .ZN(n5442) );
  NOR2_X1 U6410 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5441), .ZN(n5450) );
  OAI21_X1 U6411 ( .B1(n5442), .B2(n5450), .A(REIP_REG_25__SCAN_IN), .ZN(n5443) );
  NAND4_X1 U6412 ( .A1(n5446), .A2(n5445), .A3(n5444), .A4(n5443), .ZN(U2802)
         );
  OAI22_X1 U6413 ( .A1(n5448), .A2(n5718), .B1(n6578), .B2(n5447), .ZN(n5449)
         );
  AOI211_X1 U6414 ( .C1(n5699), .C2(EBX_REG_24__SCAN_IN), .A(n5450), .B(n5449), 
        .ZN(n5453) );
  AOI22_X1 U6415 ( .A1(n5493), .A2(n5679), .B1(n5451), .B2(n5654), .ZN(n5452)
         );
  OAI211_X1 U6416 ( .C1(n5454), .C2(n5711), .A(n5453), .B(n5452), .ZN(U2803)
         );
  OAI22_X1 U6417 ( .A1(n5709), .A2(n5456), .B1(REIP_REG_21__SCAN_IN), .B2(
        n5455), .ZN(n5459) );
  INV_X1 U6418 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5457) );
  OAI22_X1 U6419 ( .A1(n5457), .A2(n5718), .B1(n6796), .B2(n5708), .ZN(n5458)
         );
  AOI221_X1 U6420 ( .B1(n5460), .B2(n4761), .C1(n5459), .C2(
        REIP_REG_22__SCAN_IN), .A(n5458), .ZN(n5463) );
  AOI22_X1 U6421 ( .A1(n5496), .A2(n5679), .B1(n5461), .B2(n5654), .ZN(n5462)
         );
  OAI211_X1 U6422 ( .C1(n5464), .C2(n5711), .A(n5463), .B(n5462), .ZN(U2805)
         );
  NAND2_X1 U6423 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5465) );
  OAI21_X1 U6424 ( .B1(n5581), .B2(n5465), .A(n6575), .ZN(n5466) );
  AOI22_X1 U6425 ( .A1(EBX_REG_20__SCAN_IN), .A2(n5699), .B1(n5467), .B2(n5466), .ZN(n5472) );
  OAI22_X1 U6426 ( .A1(n5469), .A2(n5711), .B1(n5509), .B2(n5717), .ZN(n5470)
         );
  AOI21_X1 U6427 ( .B1(n5505), .B2(n5679), .A(n5470), .ZN(n5471) );
  OAI211_X1 U6428 ( .C1(n4178), .C2(n5718), .A(n5472), .B(n5471), .ZN(U2807)
         );
  NOR2_X1 U6429 ( .A1(n5581), .A2(n6572), .ZN(n5476) );
  OAI21_X1 U6430 ( .B1(n6572), .B2(n5474), .A(n5473), .ZN(n5580) );
  INV_X1 U6431 ( .A(n5580), .ZN(n5475) );
  MUX2_X1 U6432 ( .A(n5476), .B(n5475), .S(REIP_REG_19__SCAN_IN), .Z(n5477) );
  AOI211_X1 U6433 ( .C1(n5696), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5695), 
        .B(n5477), .ZN(n5484) );
  OAI22_X1 U6434 ( .A1(n5480), .A2(n5479), .B1(n5478), .B2(n5711), .ZN(n5481)
         );
  AOI21_X1 U6435 ( .B1(n5482), .B2(n5654), .A(n5481), .ZN(n5483) );
  OAI211_X1 U6436 ( .C1(n5485), .C2(n5708), .A(n5484), .B(n5483), .ZN(U2808)
         );
  AOI22_X1 U6437 ( .A1(n5490), .A2(n5731), .B1(n5486), .B2(n5730), .ZN(n5487)
         );
  OAI21_X1 U6438 ( .B1(n5733), .B2(n5488), .A(n5487), .ZN(U2834) );
  INV_X1 U6439 ( .A(n5489), .ZN(n5738) );
  AOI22_X1 U6440 ( .A1(n5490), .A2(n5738), .B1(n5737), .B2(DATAI_25_), .ZN(
        n5492) );
  AOI22_X1 U6441 ( .A1(n5741), .A2(DATAI_9_), .B1(n5740), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U6442 ( .A1(n5492), .A2(n5491), .ZN(U2866) );
  AOI22_X1 U6443 ( .A1(n5493), .A2(n5738), .B1(DATAI_24_), .B2(n5737), .ZN(
        n5495) );
  AOI22_X1 U6444 ( .A1(n5741), .A2(DATAI_8_), .B1(n5740), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U6445 ( .A1(n5495), .A2(n5494), .ZN(U2867) );
  AOI22_X1 U6446 ( .A1(n5496), .A2(n5738), .B1(n5737), .B2(DATAI_22_), .ZN(
        n5498) );
  AOI22_X1 U6447 ( .A1(n5741), .A2(DATAI_6_), .B1(n5740), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U6448 ( .A1(n5498), .A2(n5497), .ZN(U2869) );
  INV_X1 U6449 ( .A(n5499), .ZN(n5500) );
  AOI22_X1 U6450 ( .A1(n5500), .A2(n5738), .B1(n5737), .B2(DATAI_21_), .ZN(
        n5502) );
  AOI22_X1 U6451 ( .A1(n5741), .A2(DATAI_5_), .B1(n5740), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U6452 ( .A1(n5502), .A2(n5501), .ZN(U2870) );
  AOI22_X1 U6453 ( .A1(n5505), .A2(n5738), .B1(n5737), .B2(DATAI_20_), .ZN(
        n5504) );
  AOI22_X1 U6454 ( .A1(n5741), .A2(DATAI_4_), .B1(n5740), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U6455 ( .A1(n5504), .A2(n5503), .ZN(U2871) );
  AOI22_X1 U6456 ( .A1(n5829), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .B1(n5931), 
        .B2(REIP_REG_20__SCAN_IN), .ZN(n5508) );
  AOI22_X1 U6457 ( .A1(n5506), .A2(n5850), .B1(n5851), .B2(n5505), .ZN(n5507)
         );
  OAI211_X1 U6458 ( .C1(n5856), .C2(n5509), .A(n5508), .B(n5507), .ZN(U2966)
         );
  AOI22_X1 U6459 ( .A1(n5829), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .B1(n5931), 
        .B2(REIP_REG_18__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U6460 ( .A1(n5511), .A2(n5510), .ZN(n5512) );
  XNOR2_X1 U6461 ( .A(n5512), .B(n5527), .ZN(n5526) );
  AOI22_X1 U6462 ( .A1(n5526), .A2(n5850), .B1(n5851), .B2(n5734), .ZN(n5513)
         );
  OAI211_X1 U6463 ( .C1(n5856), .C2(n5585), .A(n5514), .B(n5513), .ZN(U2968)
         );
  AOI22_X1 U6464 ( .A1(n5829), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .B1(n5931), 
        .B2(REIP_REG_13__SCAN_IN), .ZN(n5522) );
  OR2_X1 U6465 ( .A1(n5516), .A2(n5515), .ZN(n5518) );
  NAND2_X1 U6466 ( .A1(n5518), .A2(n5517), .ZN(n5520) );
  XNOR2_X1 U6467 ( .A(n5520), .B(n5519), .ZN(n5544) );
  AOI22_X1 U6468 ( .A1(n5544), .A2(n5850), .B1(n5851), .B2(n5722), .ZN(n5521)
         );
  OAI211_X1 U6469 ( .C1(n5856), .C2(n5635), .A(n5522), .B(n5521), .ZN(U2973)
         );
  INV_X1 U6470 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5527) );
  OAI22_X1 U6471 ( .A1(n5524), .A2(n5527), .B1(n5903), .B2(n5523), .ZN(n5525)
         );
  AOI21_X1 U6472 ( .B1(n5929), .B2(n5526), .A(n5525), .ZN(n5529) );
  NAND3_X1 U6473 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5535), .A3(n5527), .ZN(n5528) );
  OAI211_X1 U6474 ( .C1(n6572), .C2(n5912), .A(n5529), .B(n5528), .ZN(U3000)
         );
  AOI22_X1 U6475 ( .A1(n5531), .A2(n5929), .B1(n5927), .B2(n5530), .ZN(n5537)
         );
  NOR2_X1 U6476 ( .A1(n5912), .A2(n6570), .ZN(n5532) );
  AOI221_X1 U6477 ( .B1(n5535), .B2(n5534), .C1(n5533), .C2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5532), .ZN(n5536) );
  NAND2_X1 U6478 ( .A1(n5537), .A2(n5536), .ZN(U3001) );
  INV_X1 U6479 ( .A(n5538), .ZN(n5547) );
  NOR2_X1 U6480 ( .A1(n5540), .A2(n5539), .ZN(n5541) );
  OR2_X1 U6481 ( .A1(n5542), .A2(n5541), .ZN(n5719) );
  INV_X1 U6482 ( .A(n5719), .ZN(n5625) );
  AOI22_X1 U6483 ( .A1(n5927), .A2(n5625), .B1(n5931), .B2(
        REIP_REG_13__SCAN_IN), .ZN(n5546) );
  AOI22_X1 U6484 ( .A1(n5544), .A2(n5929), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5543), .ZN(n5545) );
  OAI211_X1 U6485 ( .C1(n5548), .C2(n5547), .A(n5546), .B(n5545), .ZN(U3005)
         );
  OR4_X1 U6486 ( .A1(n5551), .A2(n5550), .A3(n5549), .A4(n5697), .ZN(n5552) );
  OAI21_X1 U6487 ( .B1(n5554), .B2(n5553), .A(n5552), .ZN(U3455) );
  INV_X1 U6488 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6545) );
  INV_X1 U6489 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6527) );
  AOI21_X1 U6490 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6545), .A(n6527), .ZN(n5561) );
  INV_X1 U6491 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5555) );
  INV_X1 U6492 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6535) );
  NOR2_X2 U6493 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6535), .ZN(n6621) );
  AOI21_X1 U6494 ( .B1(n5561), .B2(n5555), .A(n6621), .ZN(U2789) );
  OAI21_X1 U6495 ( .B1(n5557), .B2(n5556), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5558) );
  OAI21_X1 U6496 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5559), .A(n5558), .ZN(
        U2790) );
  NOR2_X1 U6497 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5562) );
  OAI21_X1 U6498 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5562), .A(n6609), .ZN(n5560)
         );
  OAI21_X1 U6499 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6609), .A(n5560), .ZN(
        U2791) );
  NOR2_X1 U6500 ( .A1(n6621), .A2(n5561), .ZN(n6596) );
  OAI21_X1 U6501 ( .B1(BS16_N), .B2(n5562), .A(n6596), .ZN(n6594) );
  OAI21_X1 U6502 ( .B1(n6596), .B2(n6411), .A(n6594), .ZN(U2792) );
  OAI21_X1 U6503 ( .B1(n5564), .B2(n5563), .A(n5814), .ZN(U2793) );
  NOR4_X1 U6504 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n5568) );
  NOR4_X1 U6505 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(DATAWIDTH_REG_13__SCAN_IN), .ZN(n5567)
         );
  NOR4_X1 U6506 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5566) );
  NOR4_X1 U6507 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_22__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n5565) );
  NAND4_X1 U6508 ( .A1(n5568), .A2(n5567), .A3(n5566), .A4(n5565), .ZN(n5574)
         );
  NOR4_X1 U6509 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_28__SCAN_IN), .ZN(n5572) );
  AOI211_X1 U6510 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_3__SCAN_IN), .B(
        DATAWIDTH_REG_8__SCAN_IN), .ZN(n5571) );
  NOR4_X1 U6511 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n5570) );
  NOR4_X1 U6512 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n5569) );
  NAND4_X1 U6513 ( .A1(n5572), .A2(n5571), .A3(n5570), .A4(n5569), .ZN(n5573)
         );
  NOR2_X1 U6514 ( .A1(n5574), .A2(n5573), .ZN(n6604) );
  INV_X1 U6515 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5576) );
  NOR3_X1 U6516 ( .A1(DATAWIDTH_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5577) );
  OAI21_X1 U6517 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5577), .A(n6604), .ZN(n5575)
         );
  OAI21_X1 U6518 ( .B1(n6604), .B2(n5576), .A(n5575), .ZN(U2794) );
  INV_X1 U6519 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6595) );
  AOI21_X1 U6520 ( .B1(n6601), .B2(n6595), .A(n5577), .ZN(n5579) );
  INV_X1 U6521 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5578) );
  INV_X1 U6522 ( .A(n6604), .ZN(n6607) );
  AOI22_X1 U6523 ( .A1(n6604), .A2(n5579), .B1(n5578), .B2(n6607), .ZN(U2795)
         );
  AOI21_X1 U6524 ( .B1(n5581), .B2(n6572), .A(n5580), .ZN(n5582) );
  AOI211_X1 U6525 ( .C1(n5699), .C2(EBX_REG_18__SCAN_IN), .A(n5695), .B(n5582), 
        .ZN(n5588) );
  NAND2_X1 U6526 ( .A1(n5583), .A2(n5687), .ZN(n5584) );
  OAI21_X1 U6527 ( .B1(n5717), .B2(n5585), .A(n5584), .ZN(n5586) );
  AOI21_X1 U6528 ( .B1(n5734), .B2(n5679), .A(n5586), .ZN(n5587) );
  OAI211_X1 U6529 ( .C1(n4114), .C2(n5718), .A(n5588), .B(n5587), .ZN(U2809)
         );
  NOR3_X1 U6530 ( .A1(n5667), .A2(REIP_REG_15__SCAN_IN), .A3(n5589), .ZN(n5601) );
  NAND2_X1 U6531 ( .A1(n5612), .A2(n5589), .ZN(n5590) );
  NAND2_X1 U6532 ( .A1(n5591), .A2(n5590), .ZN(n5610) );
  OAI21_X1 U6533 ( .B1(n5601), .B2(n5610), .A(REIP_REG_16__SCAN_IN), .ZN(n5594) );
  INV_X1 U6534 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6568) );
  NAND3_X1 U6535 ( .A1(n5612), .A2(n6568), .A3(n5592), .ZN(n5593) );
  OAI211_X1 U6536 ( .C1(n5708), .C2(n5595), .A(n5594), .B(n5593), .ZN(n5596)
         );
  AOI211_X1 U6537 ( .C1(n5696), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5695), 
        .B(n5596), .ZN(n5599) );
  AOI22_X1 U6538 ( .A1(n5739), .A2(n5679), .B1(n5654), .B2(n5597), .ZN(n5598)
         );
  OAI211_X1 U6539 ( .C1(n5711), .C2(n5600), .A(n5599), .B(n5598), .ZN(U2811)
         );
  AOI22_X1 U6540 ( .A1(EBX_REG_15__SCAN_IN), .A2(n5699), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5610), .ZN(n5609) );
  AOI211_X1 U6541 ( .C1(n5696), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5695), 
        .B(n5601), .ZN(n5608) );
  INV_X1 U6542 ( .A(n5602), .ZN(n5603) );
  AOI22_X1 U6543 ( .A1(n5604), .A2(n5679), .B1(n5603), .B2(n5654), .ZN(n5607)
         );
  NAND2_X1 U6544 ( .A1(n5687), .A2(n5605), .ZN(n5606) );
  NAND4_X1 U6545 ( .A1(n5609), .A2(n5608), .A3(n5607), .A4(n5606), .ZN(U2812)
         );
  INV_X1 U6546 ( .A(n5610), .ZN(n5622) );
  AOI21_X1 U6547 ( .B1(n5612), .B2(n5611), .A(REIP_REG_14__SCAN_IN), .ZN(n5621) );
  OAI22_X1 U6548 ( .A1(n5614), .A2(n5718), .B1(n5711), .B2(n5613), .ZN(n5615)
         );
  AOI211_X1 U6549 ( .C1(n5699), .C2(EBX_REG_14__SCAN_IN), .A(n5695), .B(n5615), 
        .ZN(n5620) );
  INV_X1 U6550 ( .A(n5616), .ZN(n5618) );
  AOI22_X1 U6551 ( .A1(n5618), .A2(n5679), .B1(n5654), .B2(n5617), .ZN(n5619)
         );
  OAI211_X1 U6552 ( .C1(n5622), .C2(n5621), .A(n5620), .B(n5619), .ZN(U2813)
         );
  INV_X1 U6553 ( .A(n5623), .ZN(n5624) );
  NAND2_X1 U6554 ( .A1(n6563), .A2(n5624), .ZN(n5629) );
  AOI22_X1 U6555 ( .A1(EBX_REG_13__SCAN_IN), .A2(n5699), .B1(n5687), .B2(n5625), .ZN(n5626) );
  NAND2_X1 U6556 ( .A1(n5661), .A2(n5626), .ZN(n5627) );
  AOI21_X1 U6557 ( .B1(n5696), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5627), 
        .ZN(n5628) );
  OAI21_X1 U6558 ( .B1(n5667), .B2(n5629), .A(n5628), .ZN(n5630) );
  AOI21_X1 U6559 ( .B1(n5722), .B2(n5679), .A(n5630), .ZN(n5634) );
  OAI21_X1 U6560 ( .B1(n5632), .B2(n5631), .A(REIP_REG_13__SCAN_IN), .ZN(n5633) );
  OAI211_X1 U6561 ( .C1(n5717), .C2(n5635), .A(n5634), .B(n5633), .ZN(U2814)
         );
  INV_X1 U6562 ( .A(n5636), .ZN(n5640) );
  INV_X1 U6563 ( .A(n5637), .ZN(n5639) );
  AOI21_X1 U6564 ( .B1(n5640), .B2(n5639), .A(n5638), .ZN(n5875) );
  AOI22_X1 U6565 ( .A1(EBX_REG_9__SCAN_IN), .A2(n5699), .B1(n5687), .B2(n5875), 
        .ZN(n5641) );
  OAI21_X1 U6566 ( .B1(n6969), .B2(n5658), .A(n5641), .ZN(n5642) );
  AOI211_X1 U6567 ( .C1(n5696), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n5695), 
        .B(n5642), .ZN(n5646) );
  INV_X1 U6568 ( .A(n5643), .ZN(n5724) );
  AOI22_X1 U6569 ( .A1(n5724), .A2(n5679), .B1(n5654), .B2(n5644), .ZN(n5645)
         );
  OAI211_X1 U6570 ( .C1(REIP_REG_9__SCAN_IN), .C2(n5647), .A(n5646), .B(n5645), 
        .ZN(U2818) );
  AOI21_X1 U6571 ( .B1(n5648), .B2(n5688), .A(REIP_REG_8__SCAN_IN), .ZN(n5659)
         );
  OAI22_X1 U6572 ( .A1(n5650), .A2(n5708), .B1(n5711), .B2(n5649), .ZN(n5651)
         );
  AOI211_X1 U6573 ( .C1(n5696), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n5695), 
        .B(n5651), .ZN(n5657) );
  INV_X1 U6574 ( .A(n5652), .ZN(n5653) );
  AOI22_X1 U6575 ( .A1(n5655), .A2(n5679), .B1(n5654), .B2(n5653), .ZN(n5656)
         );
  OAI211_X1 U6576 ( .C1(n5659), .C2(n5658), .A(n5657), .B(n5656), .ZN(U2819)
         );
  INV_X1 U6577 ( .A(n5660), .ZN(n5819) );
  AOI22_X1 U6578 ( .A1(EBX_REG_7__SCAN_IN), .A2(n5699), .B1(n5687), .B2(n5881), 
        .ZN(n5662) );
  OAI211_X1 U6579 ( .C1(n5718), .C2(n3935), .A(n5662), .B(n5661), .ZN(n5665)
         );
  INV_X1 U6580 ( .A(n5663), .ZN(n5668) );
  NAND2_X1 U6581 ( .A1(n5688), .A2(n5668), .ZN(n5669) );
  NOR3_X1 U6582 ( .A1(n5669), .A2(REIP_REG_7__SCAN_IN), .A3(n6554), .ZN(n5664)
         );
  AOI211_X1 U6583 ( .C1(n5819), .C2(n5679), .A(n5665), .B(n5664), .ZN(n5671)
         );
  OAI21_X1 U6584 ( .B1(n5668), .B2(n5667), .A(n5666), .ZN(n5689) );
  NOR2_X1 U6585 ( .A1(n5669), .A2(REIP_REG_6__SCAN_IN), .ZN(n5673) );
  OAI21_X1 U6586 ( .B1(n5689), .B2(n5673), .A(REIP_REG_7__SCAN_IN), .ZN(n5670)
         );
  OAI211_X1 U6587 ( .C1(n5717), .C2(n5822), .A(n5671), .B(n5670), .ZN(U2820)
         );
  AOI22_X1 U6588 ( .A1(EBX_REG_6__SCAN_IN), .A2(n5699), .B1(
        REIP_REG_6__SCAN_IN), .B2(n5689), .ZN(n5677) );
  AOI21_X1 U6589 ( .B1(n5696), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5695), 
        .ZN(n5676) );
  NAND2_X1 U6590 ( .A1(n5687), .A2(n5672), .ZN(n5675) );
  INV_X1 U6591 ( .A(n5673), .ZN(n5674) );
  NAND4_X1 U6592 ( .A1(n5677), .A2(n5676), .A3(n5675), .A4(n5674), .ZN(n5678)
         );
  AOI21_X1 U6593 ( .B1(n5679), .B2(n5824), .A(n5678), .ZN(n5680) );
  OAI21_X1 U6594 ( .B1(n5828), .B2(n5717), .A(n5680), .ZN(U2821) );
  OR2_X1 U6595 ( .A1(n5682), .A2(n5681), .ZN(n5684) );
  AND2_X1 U6596 ( .A1(n5684), .A2(n5683), .ZN(n5891) );
  INV_X1 U6597 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6653) );
  OAI22_X1 U6598 ( .A1(n5685), .A2(n5718), .B1(n6653), .B2(n5708), .ZN(n5686)
         );
  AOI211_X1 U6599 ( .C1(n5687), .C2(n5891), .A(n5695), .B(n5686), .ZN(n5692)
         );
  INV_X1 U6600 ( .A(n5688), .ZN(n5693) );
  INV_X1 U6601 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6550) );
  INV_X1 U6602 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6552) );
  OAI21_X1 U6603 ( .B1(n5693), .B2(n6550), .A(n6552), .ZN(n5690) );
  AOI22_X1 U6604 ( .A1(n5690), .A2(n5689), .B1(n5834), .B2(n5714), .ZN(n5691)
         );
  OAI211_X1 U6605 ( .C1(n5837), .C2(n5717), .A(n5692), .B(n5691), .ZN(U2822)
         );
  OAI22_X1 U6606 ( .A1(REIP_REG_4__SCAN_IN), .A2(n5693), .B1(n5711), .B2(n5902), .ZN(n5694) );
  AOI211_X1 U6607 ( .C1(n5696), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5695), 
        .B(n5694), .ZN(n5704) );
  INV_X1 U6608 ( .A(n5697), .ZN(n5698) );
  AOI22_X1 U6609 ( .A1(n5699), .A2(EBX_REG_4__SCAN_IN), .B1(n5706), .B2(n5698), 
        .ZN(n5703) );
  NAND2_X1 U6610 ( .A1(n5700), .A2(REIP_REG_4__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U6611 ( .A1(n5842), .A2(n5714), .ZN(n5701) );
  AND4_X1 U6612 ( .A1(n5704), .A2(n5703), .A3(n5702), .A4(n5701), .ZN(n5705)
         );
  OAI21_X1 U6613 ( .B1(n5846), .B2(n5717), .A(n5705), .ZN(U2823) );
  INV_X1 U6614 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n6994) );
  INV_X1 U6615 ( .A(n5706), .ZN(n5707) );
  INV_X1 U6616 ( .A(n6244), .ZN(n6304) );
  OAI22_X1 U6617 ( .A1(n5708), .A2(n4356), .B1(n5707), .B2(n6304), .ZN(n5713)
         );
  OAI22_X1 U6618 ( .A1(n5711), .A2(n5710), .B1(n5709), .B2(n6606), .ZN(n5712)
         );
  AOI211_X1 U6619 ( .C1(n5715), .C2(n5714), .A(n5713), .B(n5712), .ZN(n5716)
         );
  OAI221_X1 U6620 ( .B1(n6994), .B2(n5718), .C1(n6994), .C2(n5717), .A(n5716), 
        .ZN(U2827) );
  INV_X1 U6621 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6902) );
  NOR2_X1 U6622 ( .A1(n5720), .A2(n5719), .ZN(n5721) );
  AOI21_X1 U6623 ( .B1(n5722), .B2(n5731), .A(n5721), .ZN(n5723) );
  OAI21_X1 U6624 ( .B1(n5733), .B2(n6902), .A(n5723), .ZN(U2846) );
  AOI22_X1 U6625 ( .A1(n5724), .A2(n5731), .B1(n5730), .B2(n5875), .ZN(n5725)
         );
  OAI21_X1 U6626 ( .B1(n5733), .B2(n5726), .A(n5725), .ZN(U2850) );
  AOI22_X1 U6627 ( .A1(n5834), .A2(n5731), .B1(n5730), .B2(n5891), .ZN(n5727)
         );
  OAI21_X1 U6628 ( .B1(n5733), .B2(n6653), .A(n5727), .ZN(U2854) );
  INV_X1 U6629 ( .A(n5728), .ZN(n5852) );
  INV_X1 U6630 ( .A(n5729), .ZN(n5926) );
  AOI22_X1 U6631 ( .A1(n5852), .A2(n5731), .B1(n5730), .B2(n5926), .ZN(n5732)
         );
  OAI21_X1 U6632 ( .B1(n5733), .B2(n6933), .A(n5732), .ZN(U2857) );
  AOI22_X1 U6633 ( .A1(n5734), .A2(n5738), .B1(n5737), .B2(DATAI_18_), .ZN(
        n5736) );
  AOI22_X1 U6634 ( .A1(n5741), .A2(DATAI_2_), .B1(n5740), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U6635 ( .A1(n5736), .A2(n5735), .ZN(U2873) );
  AOI22_X1 U6636 ( .A1(n5739), .A2(n5738), .B1(n5737), .B2(DATAI_16_), .ZN(
        n5743) );
  AOI22_X1 U6637 ( .A1(n5741), .A2(DATAI_0_), .B1(n5740), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U6638 ( .A1(n5743), .A2(n5742), .ZN(U2875) );
  INV_X1 U6639 ( .A(n5744), .ZN(n5750) );
  AOI22_X1 U6640 ( .A1(n5775), .A2(DATAO_REG_29__SCAN_IN), .B1(n5750), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5745) );
  OAI21_X1 U6641 ( .B1(n6785), .B2(n5749), .A(n5745), .ZN(U2894) );
  INV_X1 U6642 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n6934) );
  AOI22_X1 U6643 ( .A1(n5750), .A2(EAX_REG_22__SCAN_IN), .B1(n6613), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n5746) );
  OAI21_X1 U6644 ( .B1(n6934), .B2(n5762), .A(n5746), .ZN(U2901) );
  INV_X1 U6645 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n6893) );
  AOI22_X1 U6646 ( .A1(n5750), .A2(EAX_REG_21__SCAN_IN), .B1(n6613), .B2(
        UWORD_REG_5__SCAN_IN), .ZN(n5747) );
  OAI21_X1 U6647 ( .B1(n6893), .B2(n5762), .A(n5747), .ZN(U2902) );
  INV_X1 U6648 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n6921) );
  AOI22_X1 U6649 ( .A1(n5775), .A2(DATAO_REG_19__SCAN_IN), .B1(n5750), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5748) );
  OAI21_X1 U6650 ( .B1(n6921), .B2(n5749), .A(n5748), .ZN(U2904) );
  INV_X1 U6651 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n6891) );
  AOI22_X1 U6652 ( .A1(n5750), .A2(EAX_REG_18__SCAN_IN), .B1(n6613), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n5751) );
  OAI21_X1 U6653 ( .B1(n6891), .B2(n5762), .A(n5751), .ZN(U2905) );
  INV_X1 U6654 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6964) );
  AOI22_X1 U6655 ( .A1(n5769), .A2(LWORD_REG_15__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5752) );
  OAI21_X1 U6656 ( .B1(n6964), .B2(n5777), .A(n5752), .ZN(U2908) );
  AOI22_X1 U6657 ( .A1(n5769), .A2(LWORD_REG_14__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5753) );
  OAI21_X1 U6658 ( .B1(n4684), .B2(n5777), .A(n5753), .ZN(U2909) );
  INV_X1 U6659 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n6847) );
  AOI22_X1 U6660 ( .A1(EAX_REG_13__SCAN_IN), .A2(n5768), .B1(n5769), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n5754) );
  OAI21_X1 U6661 ( .B1(n6847), .B2(n5762), .A(n5754), .ZN(U2910) );
  INV_X1 U6662 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5756) );
  AOI22_X1 U6663 ( .A1(n6613), .A2(LWORD_REG_12__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5755) );
  OAI21_X1 U6664 ( .B1(n5756), .B2(n5777), .A(n5755), .ZN(U2911) );
  INV_X1 U6665 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5758) );
  AOI22_X1 U6666 ( .A1(n6613), .A2(LWORD_REG_11__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5757) );
  OAI21_X1 U6667 ( .B1(n5758), .B2(n5777), .A(n5757), .ZN(U2912) );
  INV_X1 U6668 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5760) );
  AOI22_X1 U6669 ( .A1(n6613), .A2(LWORD_REG_10__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5759) );
  OAI21_X1 U6670 ( .B1(n5760), .B2(n5777), .A(n5759), .ZN(U2913) );
  INV_X1 U6671 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n6980) );
  AOI22_X1 U6672 ( .A1(EAX_REG_9__SCAN_IN), .A2(n5768), .B1(n5769), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n5761) );
  OAI21_X1 U6673 ( .B1(n6980), .B2(n5762), .A(n5761), .ZN(U2914) );
  AOI22_X1 U6674 ( .A1(n6613), .A2(LWORD_REG_8__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5763) );
  OAI21_X1 U6675 ( .B1(n5764), .B2(n5777), .A(n5763), .ZN(U2915) );
  AOI22_X1 U6676 ( .A1(n6613), .A2(LWORD_REG_7__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5765) );
  OAI21_X1 U6677 ( .B1(n3936), .B2(n5777), .A(n5765), .ZN(U2916) );
  AOI22_X1 U6678 ( .A1(n6613), .A2(LWORD_REG_6__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5766) );
  OAI21_X1 U6679 ( .B1(n5767), .B2(n5777), .A(n5766), .ZN(U2917) );
  AOI222_X1 U6680 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n5769), .B1(n5768), .B2(
        EAX_REG_5__SCAN_IN), .C1(n5775), .C2(DATAO_REG_5__SCAN_IN), .ZN(n5770)
         );
  INV_X1 U6681 ( .A(n5770), .ZN(U2918) );
  AOI22_X1 U6682 ( .A1(n6613), .A2(LWORD_REG_4__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5771) );
  OAI21_X1 U6683 ( .B1(n3916), .B2(n5777), .A(n5771), .ZN(U2919) );
  AOI22_X1 U6684 ( .A1(n6613), .A2(LWORD_REG_3__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5772) );
  OAI21_X1 U6685 ( .B1(n3904), .B2(n5777), .A(n5772), .ZN(U2920) );
  AOI22_X1 U6686 ( .A1(n6613), .A2(LWORD_REG_2__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5773) );
  OAI21_X1 U6687 ( .B1(n3893), .B2(n5777), .A(n5773), .ZN(U2921) );
  AOI22_X1 U6688 ( .A1(n6613), .A2(LWORD_REG_1__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5774) );
  OAI21_X1 U6689 ( .B1(n4301), .B2(n5777), .A(n5774), .ZN(U2922) );
  AOI22_X1 U6690 ( .A1(n6613), .A2(LWORD_REG_0__SCAN_IN), .B1(n5775), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5776) );
  OAI21_X1 U6691 ( .B1(n5778), .B2(n5777), .A(n5776), .ZN(U2923) );
  AOI22_X1 U6692 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n5798), .B1(n5801), .B2(
        DATAI_0_), .ZN(n5779) );
  OAI21_X1 U6693 ( .B1(n6887), .B2(n5803), .A(n5779), .ZN(U2924) );
  AOI22_X1 U6694 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n5798), .B1(n5801), .B2(
        DATAI_1_), .ZN(n5780) );
  OAI21_X1 U6695 ( .B1(n5781), .B2(n5803), .A(n5780), .ZN(U2925) );
  NAND2_X1 U6696 ( .A1(n5801), .A2(DATAI_10_), .ZN(n5791) );
  INV_X1 U6697 ( .A(n5791), .ZN(n5782) );
  AOI21_X1 U6698 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n5798), .A(n5782), .ZN(
        n5783) );
  OAI21_X1 U6699 ( .B1(n4821), .B2(n5803), .A(n5783), .ZN(U2934) );
  NAND2_X1 U6700 ( .A1(n5801), .A2(DATAI_11_), .ZN(n5793) );
  INV_X1 U6701 ( .A(n5793), .ZN(n5784) );
  AOI21_X1 U6702 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n5798), .A(n5784), .ZN(
        n5785) );
  OAI21_X1 U6703 ( .B1(n5786), .B2(n5803), .A(n5785), .ZN(U2935) );
  NAND2_X1 U6704 ( .A1(n5801), .A2(DATAI_12_), .ZN(n5795) );
  INV_X1 U6705 ( .A(n5795), .ZN(n5787) );
  AOI21_X1 U6706 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n5798), .A(n5787), .ZN(
        n5788) );
  OAI21_X1 U6707 ( .B1(n6867), .B2(n5803), .A(n5788), .ZN(U2936) );
  AOI22_X1 U6708 ( .A1(UWORD_REG_14__SCAN_IN), .A2(n5798), .B1(n5801), .B2(
        DATAI_14_), .ZN(n5789) );
  OAI21_X1 U6709 ( .B1(n5790), .B2(n5803), .A(n5789), .ZN(U2938) );
  AOI22_X1 U6710 ( .A1(n4393), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n5797), .ZN(n5792) );
  NAND2_X1 U6711 ( .A1(n5792), .A2(n5791), .ZN(U2949) );
  AOI22_X1 U6712 ( .A1(n5798), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n5797), .ZN(n5794) );
  NAND2_X1 U6713 ( .A1(n5794), .A2(n5793), .ZN(U2950) );
  AOI22_X1 U6714 ( .A1(n5798), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n5797), .ZN(n5796) );
  NAND2_X1 U6715 ( .A1(n5796), .A2(n5795), .ZN(U2951) );
  AOI22_X1 U6716 ( .A1(n5798), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n5797), .ZN(n5800) );
  NAND2_X1 U6717 ( .A1(n5800), .A2(n5799), .ZN(U2952) );
  AOI22_X1 U6718 ( .A1(LWORD_REG_15__SCAN_IN), .A2(n5798), .B1(n5801), .B2(
        DATAI_15_), .ZN(n5802) );
  OAI21_X1 U6719 ( .B1(n6964), .B2(n5803), .A(n5802), .ZN(U2954) );
  NAND2_X1 U6720 ( .A1(n5805), .A2(n5804), .ZN(n5808) );
  XNOR2_X1 U6721 ( .A(n5806), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5807)
         );
  XNOR2_X1 U6722 ( .A(n5808), .B(n5807), .ZN(n5857) );
  AOI22_X1 U6723 ( .A1(n5829), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n5931), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n5813) );
  AOI22_X1 U6724 ( .A1(n5811), .A2(n5851), .B1(n5810), .B2(n5809), .ZN(n5812)
         );
  OAI211_X1 U6725 ( .C1(n5857), .C2(n5814), .A(n5813), .B(n5812), .ZN(U2975)
         );
  AOI22_X1 U6726 ( .A1(n5829), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .B1(n5931), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n5821) );
  OAI21_X1 U6727 ( .B1(n5817), .B2(n5816), .A(n5815), .ZN(n5818) );
  INV_X1 U6728 ( .A(n5818), .ZN(n5882) );
  AOI22_X1 U6729 ( .A1(n5882), .A2(n5850), .B1(n5851), .B2(n5819), .ZN(n5820)
         );
  OAI211_X1 U6730 ( .C1(n5856), .C2(n5822), .A(n5821), .B(n5820), .ZN(U2979)
         );
  AOI22_X1 U6731 ( .A1(n5829), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .B1(n5931), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n5827) );
  INV_X1 U6732 ( .A(n5823), .ZN(n5825) );
  AOI22_X1 U6733 ( .A1(n5825), .A2(n5850), .B1(n5851), .B2(n5824), .ZN(n5826)
         );
  OAI211_X1 U6734 ( .C1(n5856), .C2(n5828), .A(n5827), .B(n5826), .ZN(U2980)
         );
  AOI22_X1 U6735 ( .A1(n5829), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n5931), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n5836) );
  OAI21_X1 U6736 ( .B1(n5832), .B2(n5831), .A(n5830), .ZN(n5833) );
  INV_X1 U6737 ( .A(n5833), .ZN(n5892) );
  AOI22_X1 U6738 ( .A1(n5892), .A2(n5850), .B1(n5851), .B2(n5834), .ZN(n5835)
         );
  OAI211_X1 U6739 ( .C1(n5856), .C2(n5837), .A(n5836), .B(n5835), .ZN(U2981)
         );
  AOI22_X1 U6740 ( .A1(n5829), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n5931), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n5845) );
  OR2_X1 U6741 ( .A1(n5839), .A2(n5838), .ZN(n5840) );
  NAND2_X1 U6742 ( .A1(n5841), .A2(n5840), .ZN(n5907) );
  INV_X1 U6743 ( .A(n5907), .ZN(n5843) );
  AOI22_X1 U6744 ( .A1(n5843), .A2(n5850), .B1(n5851), .B2(n5842), .ZN(n5844)
         );
  OAI211_X1 U6745 ( .C1(n5856), .C2(n5846), .A(n5845), .B(n5844), .ZN(U2982)
         );
  AOI22_X1 U6746 ( .A1(n5829), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n5931), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n5854) );
  XNOR2_X1 U6747 ( .A(n5847), .B(n5932), .ZN(n5848) );
  XNOR2_X1 U6748 ( .A(n5849), .B(n5848), .ZN(n5928) );
  AOI22_X1 U6749 ( .A1(n5852), .A2(n5851), .B1(n5850), .B2(n5928), .ZN(n5853)
         );
  OAI211_X1 U6750 ( .C1(n5856), .C2(n5855), .A(n5854), .B(n5853), .ZN(U2984)
         );
  INV_X1 U6751 ( .A(n5857), .ZN(n5862) );
  AOI22_X1 U6752 ( .A1(n5927), .A2(n5858), .B1(n5931), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n5859) );
  OAI21_X1 U6753 ( .B1(n5860), .B2(n3605), .A(n5859), .ZN(n5861) );
  AOI21_X1 U6754 ( .B1(n5862), .B2(n5929), .A(n5861), .ZN(n5864) );
  NAND2_X1 U6755 ( .A1(n5864), .A2(n5863), .ZN(U3007) );
  NAND2_X1 U6756 ( .A1(n5867), .A2(n5883), .ZN(n5880) );
  AOI22_X1 U6757 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n4626), .B1(
        INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n3604), .ZN(n5872) );
  AOI21_X1 U6758 ( .B1(n5927), .B2(n5866), .A(n5865), .ZN(n5871) );
  OAI21_X1 U6759 ( .B1(n5868), .B2(n5867), .A(n5886), .ZN(n5876) );
  AOI22_X1 U6760 ( .A1(n5869), .A2(n5929), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n5876), .ZN(n5870) );
  OAI211_X1 U6761 ( .C1(n5880), .C2(n5872), .A(n5871), .B(n5870), .ZN(U3008)
         );
  INV_X1 U6762 ( .A(n5873), .ZN(n5874) );
  AOI21_X1 U6763 ( .B1(n5927), .B2(n5875), .A(n5874), .ZN(n5879) );
  AOI22_X1 U6764 ( .A1(n5877), .A2(n5929), .B1(n5876), .B2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5878) );
  OAI211_X1 U6765 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n5880), .A(n5879), 
        .B(n5878), .ZN(U3009) );
  AOI22_X1 U6766 ( .A1(n5927), .A2(n5881), .B1(n5931), .B2(REIP_REG_7__SCAN_IN), .ZN(n5885) );
  AOI22_X1 U6767 ( .A1(n3589), .A2(n5883), .B1(n5882), .B2(n5929), .ZN(n5884)
         );
  OAI211_X1 U6768 ( .C1(n5886), .C2(n3589), .A(n5885), .B(n5884), .ZN(U3011)
         );
  OAI21_X1 U6769 ( .B1(n5897), .B2(n5888), .A(n5887), .ZN(n5889) );
  AOI21_X1 U6770 ( .B1(n5890), .B2(n5933), .A(n5889), .ZN(n5895) );
  AOI22_X1 U6771 ( .A1(n5892), .A2(n5929), .B1(n5927), .B2(n5891), .ZN(n5894)
         );
  NAND2_X1 U6772 ( .A1(n5931), .A2(REIP_REG_5__SCAN_IN), .ZN(n5893) );
  OAI211_X1 U6773 ( .C1(n5896), .C2(n5895), .A(n5894), .B(n5893), .ZN(U3013)
         );
  NOR2_X1 U6774 ( .A1(n5897), .A2(n5899), .ZN(n5925) );
  NOR2_X1 U6775 ( .A1(n5925), .A2(n5930), .ZN(n5919) );
  INV_X1 U6776 ( .A(n5898), .ZN(n5900) );
  NAND2_X1 U6777 ( .A1(n5900), .A2(n5899), .ZN(n5921) );
  AOI211_X1 U6778 ( .C1(n5911), .C2(n5920), .A(n5901), .B(n5921), .ZN(n5909)
         );
  OAI22_X1 U6779 ( .A1(n5903), .A2(n5902), .B1(n6550), .B2(n5912), .ZN(n5904)
         );
  INV_X1 U6780 ( .A(n5904), .ZN(n5905) );
  OAI21_X1 U6781 ( .B1(n5907), .B2(n5906), .A(n5905), .ZN(n5908) );
  NOR2_X1 U6782 ( .A1(n5909), .A2(n5908), .ZN(n5910) );
  OAI21_X1 U6783 ( .B1(n5919), .B2(n5911), .A(n5910), .ZN(U3014) );
  NOR2_X1 U6784 ( .A1(n5912), .A2(n5119), .ZN(n5916) );
  AND3_X1 U6785 ( .A1(n5929), .A2(n5914), .A3(n5913), .ZN(n5915) );
  AOI211_X1 U6786 ( .C1(n5927), .C2(n5917), .A(n5916), .B(n5915), .ZN(n5918)
         );
  OAI221_X1 U6787 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n5921), .C1(n5920), .C2(n5919), .A(n5918), .ZN(U3015) );
  AND3_X1 U6788 ( .A1(n5923), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(n5922), 
        .ZN(n5924) );
  AOI211_X1 U6789 ( .C1(n5927), .C2(n5926), .A(n5925), .B(n5924), .ZN(n5937)
         );
  AOI22_X1 U6790 ( .A1(n5930), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n5929), 
        .B2(n5928), .ZN(n5936) );
  NAND2_X1 U6791 ( .A1(n5931), .A2(REIP_REG_2__SCAN_IN), .ZN(n5935) );
  NAND3_X1 U6792 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5933), .A3(n5932), 
        .ZN(n5934) );
  NAND4_X1 U6793 ( .A1(n5937), .A2(n5936), .A3(n5935), .A4(n5934), .ZN(U3016)
         );
  NOR2_X1 U6794 ( .A1(n6972), .A2(n5938), .ZN(U3019) );
  INV_X1 U6795 ( .A(DATAI_24_), .ZN(n5939) );
  NOR2_X1 U6796 ( .A1(n6457), .A2(n5939), .ZN(n6468) );
  INV_X1 U6797 ( .A(n6468), .ZN(n6421) );
  NAND2_X1 U6798 ( .A1(n6459), .A2(n6299), .ZN(n6514) );
  NAND3_X1 U6799 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6517), .A3(n5940), .ZN(
        n5988) );
  NOR2_X2 U6800 ( .A1(n5988), .A2(n5941), .ZN(n6456) );
  NAND3_X1 U6801 ( .A1(n6415), .A2(n6213), .A3(n6212), .ZN(n6001) );
  NOR2_X1 U6802 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6001), .ZN(n5991)
         );
  NOR2_X2 U6803 ( .A1(n5942), .A2(n6221), .ZN(n6455) );
  OR2_X1 U6804 ( .A1(n6270), .A2(n6454), .ZN(n6154) );
  INV_X1 U6805 ( .A(n6151), .ZN(n5943) );
  NAND2_X1 U6806 ( .A1(n5943), .A2(n6085), .ZN(n6219) );
  OR2_X1 U6807 ( .A1(n5948), .A2(n6799), .ZN(n6342) );
  NOR2_X1 U6808 ( .A1(n6406), .A2(n6214), .ZN(n5947) );
  INV_X1 U6809 ( .A(n5947), .ZN(n6086) );
  OAI22_X1 U6810 ( .A1(n6154), .A2(n6219), .B1(n6342), .B2(n6086), .ZN(n5990)
         );
  AOI22_X1 U6811 ( .A1(n6456), .A2(n5991), .B1(n6455), .B2(n5990), .ZN(n5953)
         );
  INV_X1 U6812 ( .A(n6216), .ZN(n5944) );
  OR2_X1 U6813 ( .A1(n6458), .A2(n5945), .ZN(n6218) );
  INV_X1 U6814 ( .A(n6218), .ZN(n6339) );
  AOI21_X1 U6815 ( .B1(n6025), .B2(n6514), .A(n6411), .ZN(n5946) );
  NOR2_X1 U6816 ( .A1(n6270), .A2(n6219), .ZN(n5997) );
  NOR3_X1 U6817 ( .A1(n5946), .A2(n5997), .A3(n6454), .ZN(n5949) );
  INV_X1 U6818 ( .A(n6221), .ZN(n6029) );
  OAI21_X1 U6819 ( .B1(n5947), .B2(n6799), .A(n6029), .ZN(n6091) );
  NAND2_X1 U6820 ( .A1(n5948), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6337) );
  INV_X1 U6821 ( .A(n6337), .ZN(n6407) );
  NOR3_X1 U6822 ( .A1(n5949), .A2(n6091), .A3(n6407), .ZN(n5950) );
  OAI21_X1 U6823 ( .B1(n5991), .B2(n6600), .A(n5950), .ZN(n5994) );
  INV_X1 U6824 ( .A(DATAI_16_), .ZN(n5951) );
  NOR2_X1 U6825 ( .A1(n6457), .A2(n5951), .ZN(n6418) );
  INV_X1 U6826 ( .A(n6025), .ZN(n6008) );
  AOI22_X1 U6827 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n5994), .B1(n6418), 
        .B2(n6008), .ZN(n5952) );
  OAI211_X1 U6828 ( .C1(n6421), .C2(n6514), .A(n5953), .B(n5952), .ZN(U3020)
         );
  INV_X1 U6829 ( .A(DATAI_17_), .ZN(n5954) );
  NOR2_X1 U6830 ( .A1(n6457), .A2(n5954), .ZN(n6348) );
  INV_X1 U6831 ( .A(n6348), .ZN(n6477) );
  NOR2_X2 U6832 ( .A1(n5988), .A2(n5955), .ZN(n6473) );
  NOR2_X2 U6833 ( .A1(n5956), .A2(n6221), .ZN(n6472) );
  AOI22_X1 U6834 ( .A1(n6473), .A2(n5991), .B1(n6472), .B2(n5990), .ZN(n5959)
         );
  INV_X1 U6835 ( .A(DATAI_25_), .ZN(n5957) );
  NOR2_X1 U6836 ( .A1(n6457), .A2(n5957), .ZN(n6474) );
  INV_X1 U6837 ( .A(n6514), .ZN(n5993) );
  AOI22_X1 U6838 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n5994), .B1(n6474), 
        .B2(n5993), .ZN(n5958) );
  OAI211_X1 U6839 ( .C1(n6477), .C2(n6025), .A(n5959), .B(n5958), .ZN(U3021)
         );
  NOR2_X1 U6840 ( .A1(n6457), .A2(n6650), .ZN(n6424) );
  INV_X1 U6841 ( .A(n6424), .ZN(n6483) );
  NOR2_X2 U6842 ( .A1(n5988), .A2(n5960), .ZN(n6479) );
  NOR2_X2 U6843 ( .A1(n5961), .A2(n6221), .ZN(n6478) );
  AOI22_X1 U6844 ( .A1(n6479), .A2(n5991), .B1(n6478), .B2(n5990), .ZN(n5964)
         );
  INV_X1 U6845 ( .A(DATAI_26_), .ZN(n5962) );
  NOR2_X1 U6846 ( .A1(n6457), .A2(n5962), .ZN(n6480) );
  AOI22_X1 U6847 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(n5994), .B1(n6480), 
        .B2(n5993), .ZN(n5963) );
  OAI211_X1 U6848 ( .C1(n6483), .C2(n6025), .A(n5964), .B(n5963), .ZN(U3022)
         );
  INV_X1 U6849 ( .A(DATAI_19_), .ZN(n5965) );
  NOR2_X1 U6850 ( .A1(n6457), .A2(n5965), .ZN(n6387) );
  INV_X1 U6851 ( .A(n6387), .ZN(n6489) );
  NOR2_X2 U6852 ( .A1(n5988), .A2(n5966), .ZN(n6485) );
  NOR2_X2 U6853 ( .A1(n5967), .A2(n6221), .ZN(n6484) );
  AOI22_X1 U6854 ( .A1(n6485), .A2(n5991), .B1(n6484), .B2(n5990), .ZN(n5969)
         );
  INV_X1 U6855 ( .A(DATAI_27_), .ZN(n6983) );
  NOR2_X1 U6856 ( .A1(n6457), .A2(n6983), .ZN(n6486) );
  AOI22_X1 U6857 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n5994), .B1(n6486), 
        .B2(n5993), .ZN(n5968) );
  OAI211_X1 U6858 ( .C1(n6489), .C2(n6025), .A(n5969), .B(n5968), .ZN(U3023)
         );
  INV_X1 U6859 ( .A(DATAI_20_), .ZN(n5970) );
  NOR2_X1 U6860 ( .A1(n6457), .A2(n5970), .ZN(n6430) );
  INV_X1 U6861 ( .A(n6430), .ZN(n6495) );
  NOR2_X2 U6862 ( .A1(n5988), .A2(n5971), .ZN(n6491) );
  NOR2_X2 U6863 ( .A1(n6979), .A2(n6221), .ZN(n6490) );
  AOI22_X1 U6864 ( .A1(n6491), .A2(n5991), .B1(n6490), .B2(n5990), .ZN(n5974)
         );
  INV_X1 U6865 ( .A(DATAI_28_), .ZN(n5972) );
  NOR2_X1 U6866 ( .A1(n6457), .A2(n5972), .ZN(n6492) );
  AOI22_X1 U6867 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n5994), .B1(n6492), 
        .B2(n5993), .ZN(n5973) );
  OAI211_X1 U6868 ( .C1(n6495), .C2(n6025), .A(n5974), .B(n5973), .ZN(U3024)
         );
  INV_X1 U6869 ( .A(DATAI_21_), .ZN(n5975) );
  NOR2_X1 U6870 ( .A1(n6457), .A2(n5975), .ZN(n6434) );
  INV_X1 U6871 ( .A(n6434), .ZN(n6501) );
  NOR2_X2 U6872 ( .A1(n5988), .A2(n5976), .ZN(n6497) );
  NOR2_X2 U6873 ( .A1(n5977), .A2(n6221), .ZN(n6496) );
  AOI22_X1 U6874 ( .A1(n6497), .A2(n5991), .B1(n6496), .B2(n5990), .ZN(n5980)
         );
  INV_X1 U6875 ( .A(DATAI_29_), .ZN(n5978) );
  NOR2_X1 U6876 ( .A1(n6457), .A2(n5978), .ZN(n6498) );
  AOI22_X1 U6877 ( .A1(INSTQUEUE_REG_0__5__SCAN_IN), .A2(n5994), .B1(n6498), 
        .B2(n5993), .ZN(n5979) );
  OAI211_X1 U6878 ( .C1(n6501), .C2(n6025), .A(n5980), .B(n5979), .ZN(U3025)
         );
  INV_X1 U6879 ( .A(DATAI_22_), .ZN(n5981) );
  NOR2_X1 U6880 ( .A1(n6457), .A2(n5981), .ZN(n6395) );
  INV_X1 U6881 ( .A(n6395), .ZN(n6507) );
  NOR2_X2 U6882 ( .A1(n5988), .A2(n5982), .ZN(n6503) );
  NOR2_X2 U6883 ( .A1(n5983), .A2(n6221), .ZN(n6502) );
  AOI22_X1 U6884 ( .A1(n6503), .A2(n5991), .B1(n6502), .B2(n5990), .ZN(n5985)
         );
  INV_X1 U6885 ( .A(DATAI_30_), .ZN(n6784) );
  NOR2_X1 U6886 ( .A1(n6457), .A2(n6784), .ZN(n6504) );
  AOI22_X1 U6887 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(n5994), .B1(n6504), 
        .B2(n5993), .ZN(n5984) );
  OAI211_X1 U6888 ( .C1(n6507), .C2(n6025), .A(n5985), .B(n5984), .ZN(U3026)
         );
  INV_X1 U6889 ( .A(DATAI_23_), .ZN(n5986) );
  NOR2_X1 U6890 ( .A1(n6457), .A2(n5986), .ZN(n6444) );
  INV_X1 U6891 ( .A(n6444), .ZN(n6632) );
  NOR2_X2 U6892 ( .A1(n5988), .A2(n5987), .ZN(n6625) );
  NOR2_X2 U6893 ( .A1(n5989), .A2(n6221), .ZN(n6627) );
  AOI22_X1 U6894 ( .A1(n6625), .A2(n5991), .B1(n6627), .B2(n5990), .ZN(n5996)
         );
  INV_X1 U6895 ( .A(DATAI_31_), .ZN(n5992) );
  NOR2_X1 U6896 ( .A1(n6457), .A2(n5992), .ZN(n6622) );
  AOI22_X1 U6897 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n5994), .B1(n6622), 
        .B2(n5993), .ZN(n5995) );
  OAI211_X1 U6898 ( .C1(n6632), .C2(n6025), .A(n5996), .B(n5995), .ZN(U3027)
         );
  NOR2_X1 U6899 ( .A1(n6370), .A2(n6001), .ZN(n6020) );
  NOR2_X2 U6900 ( .A1(n6052), .A2(n6368), .ZN(n6047) );
  AOI22_X1 U6901 ( .A1(n6456), .A2(n6020), .B1(n6047), .B2(n6418), .ZN(n6005)
         );
  AOI21_X1 U6902 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6370), .A(n6221), .ZN(
        n6465) );
  AOI21_X1 U6903 ( .B1(n5997), .B2(n6244), .A(n6020), .ZN(n6002) );
  OR2_X1 U6904 ( .A1(n6458), .A2(n6411), .ZN(n5998) );
  AOI21_X1 U6905 ( .B1(n6052), .B2(n6466), .A(n6246), .ZN(n6003) );
  INV_X1 U6906 ( .A(n6003), .ZN(n5999) );
  AOI22_X1 U6907 ( .A1(n6002), .A2(n5999), .B1(n6454), .B2(n6001), .ZN(n6000)
         );
  NAND2_X1 U6908 ( .A1(n6465), .A2(n6000), .ZN(n6022) );
  OAI22_X1 U6909 ( .A1(n6003), .A2(n6002), .B1(n6799), .B2(n6001), .ZN(n6021)
         );
  AOI22_X1 U6910 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n6022), .B1(n6455), 
        .B2(n6021), .ZN(n6004) );
  OAI211_X1 U6911 ( .C1(n6421), .C2(n6025), .A(n6005), .B(n6004), .ZN(U3028)
         );
  INV_X1 U6912 ( .A(n6474), .ZN(n6351) );
  AOI22_X1 U6913 ( .A1(n6473), .A2(n6020), .B1(n6047), .B2(n6348), .ZN(n6007)
         );
  AOI22_X1 U6914 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n6022), .B1(n6472), 
        .B2(n6021), .ZN(n6006) );
  OAI211_X1 U6915 ( .C1(n6351), .C2(n6025), .A(n6007), .B(n6006), .ZN(U3029)
         );
  INV_X1 U6916 ( .A(n6047), .ZN(n6011) );
  AOI22_X1 U6917 ( .A1(n6479), .A2(n6020), .B1(n6008), .B2(n6480), .ZN(n6010)
         );
  AOI22_X1 U6918 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n6022), .B1(n6478), 
        .B2(n6021), .ZN(n6009) );
  OAI211_X1 U6919 ( .C1(n6011), .C2(n6483), .A(n6010), .B(n6009), .ZN(U3030)
         );
  INV_X1 U6920 ( .A(n6486), .ZN(n6390) );
  AOI22_X1 U6921 ( .A1(n6485), .A2(n6020), .B1(n6047), .B2(n6387), .ZN(n6013)
         );
  AOI22_X1 U6922 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n6022), .B1(n6484), 
        .B2(n6021), .ZN(n6012) );
  OAI211_X1 U6923 ( .C1(n6390), .C2(n6025), .A(n6013), .B(n6012), .ZN(U3031)
         );
  INV_X1 U6924 ( .A(n6492), .ZN(n6433) );
  AOI22_X1 U6925 ( .A1(n6491), .A2(n6020), .B1(n6047), .B2(n6430), .ZN(n6015)
         );
  AOI22_X1 U6926 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n6022), .B1(n6490), 
        .B2(n6021), .ZN(n6014) );
  OAI211_X1 U6927 ( .C1(n6433), .C2(n6025), .A(n6015), .B(n6014), .ZN(U3032)
         );
  INV_X1 U6928 ( .A(n6498), .ZN(n6437) );
  AOI22_X1 U6929 ( .A1(n6497), .A2(n6020), .B1(n6047), .B2(n6434), .ZN(n6017)
         );
  AOI22_X1 U6930 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n6022), .B1(n6496), 
        .B2(n6021), .ZN(n6016) );
  OAI211_X1 U6931 ( .C1(n6437), .C2(n6025), .A(n6017), .B(n6016), .ZN(U3033)
         );
  INV_X1 U6932 ( .A(n6504), .ZN(n6399) );
  AOI22_X1 U6933 ( .A1(n6503), .A2(n6020), .B1(n6047), .B2(n6395), .ZN(n6019)
         );
  AOI22_X1 U6934 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n6022), .B1(n6502), 
        .B2(n6021), .ZN(n6018) );
  OAI211_X1 U6935 ( .C1(n6399), .C2(n6025), .A(n6019), .B(n6018), .ZN(U3034)
         );
  INV_X1 U6936 ( .A(n6622), .ZN(n6449) );
  AOI22_X1 U6937 ( .A1(n6625), .A2(n6020), .B1(n6047), .B2(n6444), .ZN(n6024)
         );
  AOI22_X1 U6938 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n6022), .B1(n6627), 
        .B2(n6021), .ZN(n6023) );
  OAI211_X1 U6939 ( .C1(n6449), .C2(n6025), .A(n6024), .B(n6023), .ZN(U3035)
         );
  INV_X1 U6940 ( .A(n6418), .ZN(n6471) );
  NAND2_X1 U6941 ( .A1(n6458), .A2(n3882), .ZN(n6268) );
  INV_X1 U6942 ( .A(n6268), .ZN(n6410) );
  NAND2_X1 U6943 ( .A1(n6267), .A2(n6415), .ZN(n6059) );
  NOR2_X1 U6944 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6059), .ZN(n6046)
         );
  INV_X1 U6945 ( .A(n6270), .ZN(n6026) );
  AND2_X1 U6946 ( .A1(n6085), .A2(n6151), .ZN(n6271) );
  NAND2_X1 U6947 ( .A1(n6026), .A2(n6271), .ZN(n6053) );
  INV_X1 U6948 ( .A(n6342), .ZN(n6276) );
  NAND3_X1 U6949 ( .A1(n6276), .A2(n6406), .A3(n6415), .ZN(n6027) );
  OAI21_X1 U6950 ( .B1(n6053), .B2(n6454), .A(n6027), .ZN(n6045) );
  AOI22_X1 U6951 ( .A1(n6456), .A2(n6046), .B1(n6455), .B2(n6045), .ZN(n6032)
         );
  NAND2_X1 U6952 ( .A1(n6466), .A2(n6411), .ZN(n6460) );
  OAI21_X1 U6953 ( .B1(n6078), .B2(n6047), .A(n6460), .ZN(n6028) );
  NAND2_X1 U6954 ( .A1(n6028), .A2(n6053), .ZN(n6030) );
  OAI21_X1 U6955 ( .B1(n6406), .B2(n6799), .A(n6029), .ZN(n6158) );
  NOR2_X1 U6956 ( .A1(n6407), .A2(n6158), .ZN(n6274) );
  OAI221_X1 U6957 ( .B1(n6046), .B2(n6600), .C1(n6046), .C2(n6030), .A(n6274), 
        .ZN(n6048) );
  AOI22_X1 U6958 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n6048), .B1(n6468), 
        .B2(n6047), .ZN(n6031) );
  OAI211_X1 U6959 ( .C1(n6471), .C2(n6075), .A(n6032), .B(n6031), .ZN(U3036)
         );
  AOI22_X1 U6960 ( .A1(n6473), .A2(n6046), .B1(n6472), .B2(n6045), .ZN(n6034)
         );
  AOI22_X1 U6961 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(n6048), .B1(n6047), 
        .B2(n6474), .ZN(n6033) );
  OAI211_X1 U6962 ( .C1(n6075), .C2(n6477), .A(n6034), .B(n6033), .ZN(U3037)
         );
  AOI22_X1 U6963 ( .A1(n6479), .A2(n6046), .B1(n6478), .B2(n6045), .ZN(n6036)
         );
  AOI22_X1 U6964 ( .A1(INSTQUEUE_REG_2__2__SCAN_IN), .A2(n6048), .B1(n6047), 
        .B2(n6480), .ZN(n6035) );
  OAI211_X1 U6965 ( .C1(n6075), .C2(n6483), .A(n6036), .B(n6035), .ZN(U3038)
         );
  AOI22_X1 U6966 ( .A1(n6485), .A2(n6046), .B1(n6484), .B2(n6045), .ZN(n6038)
         );
  AOI22_X1 U6967 ( .A1(INSTQUEUE_REG_2__3__SCAN_IN), .A2(n6048), .B1(n6047), 
        .B2(n6486), .ZN(n6037) );
  OAI211_X1 U6968 ( .C1(n6075), .C2(n6489), .A(n6038), .B(n6037), .ZN(U3039)
         );
  AOI22_X1 U6969 ( .A1(n6491), .A2(n6046), .B1(n6490), .B2(n6045), .ZN(n6040)
         );
  AOI22_X1 U6970 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n6048), .B1(n6047), 
        .B2(n6492), .ZN(n6039) );
  OAI211_X1 U6971 ( .C1(n6075), .C2(n6495), .A(n6040), .B(n6039), .ZN(U3040)
         );
  AOI22_X1 U6972 ( .A1(n6497), .A2(n6046), .B1(n6496), .B2(n6045), .ZN(n6042)
         );
  AOI22_X1 U6973 ( .A1(INSTQUEUE_REG_2__5__SCAN_IN), .A2(n6048), .B1(n6047), 
        .B2(n6498), .ZN(n6041) );
  OAI211_X1 U6974 ( .C1(n6075), .C2(n6501), .A(n6042), .B(n6041), .ZN(U3041)
         );
  AOI22_X1 U6975 ( .A1(n6503), .A2(n6046), .B1(n6502), .B2(n6045), .ZN(n6044)
         );
  AOI22_X1 U6976 ( .A1(INSTQUEUE_REG_2__6__SCAN_IN), .A2(n6048), .B1(n6047), 
        .B2(n6504), .ZN(n6043) );
  OAI211_X1 U6977 ( .C1(n6075), .C2(n6507), .A(n6044), .B(n6043), .ZN(U3042)
         );
  AOI22_X1 U6978 ( .A1(n6625), .A2(n6046), .B1(n6627), .B2(n6045), .ZN(n6050)
         );
  AOI22_X1 U6979 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(n6048), .B1(n6047), 
        .B2(n6622), .ZN(n6049) );
  OAI211_X1 U6980 ( .C1(n6075), .C2(n6632), .A(n6050), .B(n6049), .ZN(U3043)
         );
  NOR2_X1 U6981 ( .A1(n6301), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6079)
         );
  INV_X1 U6982 ( .A(n6113), .ZN(n6072) );
  AOI22_X1 U6983 ( .A1(n6456), .A2(n6079), .B1(n6072), .B2(n6418), .ZN(n6063)
         );
  INV_X1 U6984 ( .A(n6059), .ZN(n6058) );
  OAI21_X1 U6985 ( .B1(n6052), .B2(n6302), .A(n6466), .ZN(n6061) );
  INV_X1 U6986 ( .A(n6061), .ZN(n6056) );
  OR2_X1 U6987 ( .A1(n6053), .A2(n6304), .ZN(n6055) );
  INV_X1 U6988 ( .A(n6079), .ZN(n6054) );
  AND2_X1 U6989 ( .A1(n6055), .A2(n6054), .ZN(n6060) );
  NAND2_X1 U6990 ( .A1(n6056), .A2(n6060), .ZN(n6057) );
  OAI211_X1 U6991 ( .C1(n6466), .C2(n6058), .A(n6057), .B(n6465), .ZN(n6081)
         );
  OAI22_X1 U6992 ( .A1(n6061), .A2(n6060), .B1(n6059), .B2(n6799), .ZN(n6080)
         );
  AOI22_X1 U6993 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6081), .B1(n6455), 
        .B2(n6080), .ZN(n6062) );
  OAI211_X1 U6994 ( .C1(n6075), .C2(n6421), .A(n6063), .B(n6062), .ZN(U3044)
         );
  AOI22_X1 U6995 ( .A1(n6473), .A2(n6079), .B1(n6078), .B2(n6474), .ZN(n6065)
         );
  AOI22_X1 U6996 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6081), .B1(n6472), 
        .B2(n6080), .ZN(n6064) );
  OAI211_X1 U6997 ( .C1(n6477), .C2(n6113), .A(n6065), .B(n6064), .ZN(U3045)
         );
  INV_X1 U6998 ( .A(n6480), .ZN(n6427) );
  AOI22_X1 U6999 ( .A1(n6479), .A2(n6079), .B1(n6072), .B2(n6424), .ZN(n6067)
         );
  AOI22_X1 U7000 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6081), .B1(n6478), 
        .B2(n6080), .ZN(n6066) );
  OAI211_X1 U7001 ( .C1(n6075), .C2(n6427), .A(n6067), .B(n6066), .ZN(U3046)
         );
  AOI22_X1 U7002 ( .A1(n6485), .A2(n6079), .B1(n6072), .B2(n6387), .ZN(n6069)
         );
  AOI22_X1 U7003 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6081), .B1(n6484), 
        .B2(n6080), .ZN(n6068) );
  OAI211_X1 U7004 ( .C1(n6075), .C2(n6390), .A(n6069), .B(n6068), .ZN(U3047)
         );
  AOI22_X1 U7005 ( .A1(n6491), .A2(n6079), .B1(n6072), .B2(n6430), .ZN(n6071)
         );
  AOI22_X1 U7006 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6081), .B1(n6490), 
        .B2(n6080), .ZN(n6070) );
  OAI211_X1 U7007 ( .C1(n6075), .C2(n6433), .A(n6071), .B(n6070), .ZN(U3048)
         );
  AOI22_X1 U7008 ( .A1(n6497), .A2(n6079), .B1(n6072), .B2(n6434), .ZN(n6074)
         );
  AOI22_X1 U7009 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6081), .B1(n6496), 
        .B2(n6080), .ZN(n6073) );
  OAI211_X1 U7010 ( .C1(n6075), .C2(n6437), .A(n6074), .B(n6073), .ZN(U3049)
         );
  AOI22_X1 U7011 ( .A1(n6503), .A2(n6079), .B1(n6078), .B2(n6504), .ZN(n6077)
         );
  AOI22_X1 U7012 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6081), .B1(n6502), 
        .B2(n6080), .ZN(n6076) );
  OAI211_X1 U7013 ( .C1(n6507), .C2(n6113), .A(n6077), .B(n6076), .ZN(U3050)
         );
  AOI22_X1 U7014 ( .A1(n6625), .A2(n6079), .B1(n6078), .B2(n6622), .ZN(n6083)
         );
  AOI22_X1 U7015 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6081), .B1(n6627), 
        .B2(n6080), .ZN(n6082) );
  OAI211_X1 U7016 ( .C1(n6632), .C2(n6113), .A(n6083), .B(n6082), .ZN(U3051)
         );
  NOR2_X1 U7017 ( .A1(n6378), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6121)
         );
  INV_X1 U7018 ( .A(n6121), .ZN(n6084) );
  NOR2_X1 U7019 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6084), .ZN(n6109)
         );
  NOR2_X1 U7020 ( .A1(n6085), .A2(n6151), .ZN(n6371) );
  INV_X1 U7021 ( .A(n6371), .ZN(n6338) );
  OAI22_X1 U7022 ( .A1(n6338), .A2(n6154), .B1(n6337), .B2(n6086), .ZN(n6108)
         );
  AOI22_X1 U7023 ( .A1(n6456), .A2(n6109), .B1(n6455), .B2(n6108), .ZN(n6095)
         );
  OR2_X1 U7024 ( .A1(n6216), .A2(n6087), .ZN(n6182) );
  NOR2_X2 U7025 ( .A1(n6182), .A2(n6218), .ZN(n6144) );
  INV_X1 U7026 ( .A(n6144), .ZN(n6088) );
  AOI21_X1 U7027 ( .B1(n6088), .B2(n6113), .A(n6411), .ZN(n6090) );
  AND2_X1 U7028 ( .A1(n6371), .A2(n6089), .ZN(n6114) );
  NOR3_X1 U7029 ( .A1(n6090), .A2(n6114), .A3(n6454), .ZN(n6092) );
  NOR3_X1 U7030 ( .A1(n6092), .A2(n6091), .A3(n6276), .ZN(n6093) );
  AOI22_X1 U7031 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n6110), .B1(n6418), 
        .B2(n6144), .ZN(n6094) );
  OAI211_X1 U7032 ( .C1(n6421), .C2(n6113), .A(n6095), .B(n6094), .ZN(U3052)
         );
  AOI22_X1 U7033 ( .A1(n6473), .A2(n6109), .B1(n6472), .B2(n6108), .ZN(n6097)
         );
  AOI22_X1 U7034 ( .A1(INSTQUEUE_REG_4__1__SCAN_IN), .A2(n6110), .B1(n6348), 
        .B2(n6144), .ZN(n6096) );
  OAI211_X1 U7035 ( .C1(n6351), .C2(n6113), .A(n6097), .B(n6096), .ZN(U3053)
         );
  AOI22_X1 U7036 ( .A1(n6479), .A2(n6109), .B1(n6478), .B2(n6108), .ZN(n6099)
         );
  AOI22_X1 U7037 ( .A1(INSTQUEUE_REG_4__2__SCAN_IN), .A2(n6110), .B1(n6424), 
        .B2(n6144), .ZN(n6098) );
  OAI211_X1 U7038 ( .C1(n6427), .C2(n6113), .A(n6099), .B(n6098), .ZN(U3054)
         );
  AOI22_X1 U7039 ( .A1(n6485), .A2(n6109), .B1(n6484), .B2(n6108), .ZN(n6101)
         );
  AOI22_X1 U7040 ( .A1(INSTQUEUE_REG_4__3__SCAN_IN), .A2(n6110), .B1(n6387), 
        .B2(n6144), .ZN(n6100) );
  OAI211_X1 U7041 ( .C1(n6390), .C2(n6113), .A(n6101), .B(n6100), .ZN(U3055)
         );
  AOI22_X1 U7042 ( .A1(n6491), .A2(n6109), .B1(n6490), .B2(n6108), .ZN(n6103)
         );
  AOI22_X1 U7043 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n6110), .B1(n6430), 
        .B2(n6144), .ZN(n6102) );
  OAI211_X1 U7044 ( .C1(n6433), .C2(n6113), .A(n6103), .B(n6102), .ZN(U3056)
         );
  AOI22_X1 U7045 ( .A1(n6497), .A2(n6109), .B1(n6496), .B2(n6108), .ZN(n6105)
         );
  AOI22_X1 U7046 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(n6110), .B1(n6434), 
        .B2(n6144), .ZN(n6104) );
  OAI211_X1 U7047 ( .C1(n6437), .C2(n6113), .A(n6105), .B(n6104), .ZN(U3057)
         );
  AOI22_X1 U7048 ( .A1(n6503), .A2(n6109), .B1(n6502), .B2(n6108), .ZN(n6107)
         );
  AOI22_X1 U7049 ( .A1(INSTQUEUE_REG_4__6__SCAN_IN), .A2(n6110), .B1(n6395), 
        .B2(n6144), .ZN(n6106) );
  OAI211_X1 U7050 ( .C1(n6399), .C2(n6113), .A(n6107), .B(n6106), .ZN(U3058)
         );
  AOI22_X1 U7051 ( .A1(n6625), .A2(n6109), .B1(n6627), .B2(n6108), .ZN(n6112)
         );
  AOI22_X1 U7052 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(n6110), .B1(n6444), 
        .B2(n6144), .ZN(n6111) );
  OAI211_X1 U7053 ( .C1(n6449), .C2(n6113), .A(n6112), .B(n6111), .ZN(U3059)
         );
  INV_X1 U7054 ( .A(n6246), .ZN(n6372) );
  INV_X1 U7055 ( .A(n6182), .ZN(n6180) );
  NAND2_X1 U7056 ( .A1(n6372), .A2(n6180), .ZN(n6119) );
  NAND2_X1 U7057 ( .A1(n6114), .A2(n6244), .ZN(n6115) );
  NAND2_X1 U7058 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6121), .ZN(n6116) );
  NAND2_X1 U7059 ( .A1(n6115), .A2(n6116), .ZN(n6117) );
  AOI22_X1 U7060 ( .A1(n6119), .A2(n6117), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6121), .ZN(n6149) );
  INV_X1 U7061 ( .A(n6455), .ZN(n6124) );
  INV_X1 U7062 ( .A(n6116), .ZN(n6143) );
  AOI22_X1 U7063 ( .A1(n6456), .A2(n6143), .B1(n6150), .B2(n6418), .ZN(n6123)
         );
  INV_X1 U7064 ( .A(n6117), .ZN(n6118) );
  NAND2_X1 U7065 ( .A1(n6119), .A2(n6118), .ZN(n6120) );
  OAI211_X1 U7066 ( .C1(n6466), .C2(n6121), .A(n6120), .B(n6465), .ZN(n6145)
         );
  AOI22_X1 U7067 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n6145), .B1(n6468), 
        .B2(n6144), .ZN(n6122) );
  OAI211_X1 U7068 ( .C1(n6149), .C2(n6124), .A(n6123), .B(n6122), .ZN(U3060)
         );
  INV_X1 U7069 ( .A(n6472), .ZN(n6127) );
  AOI22_X1 U7070 ( .A1(n6473), .A2(n6143), .B1(n6144), .B2(n6474), .ZN(n6126)
         );
  AOI22_X1 U7071 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n6145), .B1(n6348), 
        .B2(n6150), .ZN(n6125) );
  OAI211_X1 U7072 ( .C1(n6149), .C2(n6127), .A(n6126), .B(n6125), .ZN(U3061)
         );
  INV_X1 U7073 ( .A(n6478), .ZN(n6130) );
  AOI22_X1 U7074 ( .A1(n6479), .A2(n6143), .B1(n6144), .B2(n6480), .ZN(n6129)
         );
  AOI22_X1 U7075 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n6145), .B1(n6424), 
        .B2(n6150), .ZN(n6128) );
  OAI211_X1 U7076 ( .C1(n6149), .C2(n6130), .A(n6129), .B(n6128), .ZN(U3062)
         );
  INV_X1 U7077 ( .A(n6484), .ZN(n6133) );
  AOI22_X1 U7078 ( .A1(n6485), .A2(n6143), .B1(n6150), .B2(n6387), .ZN(n6132)
         );
  AOI22_X1 U7079 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n6145), .B1(n6486), 
        .B2(n6144), .ZN(n6131) );
  OAI211_X1 U7080 ( .C1(n6149), .C2(n6133), .A(n6132), .B(n6131), .ZN(U3063)
         );
  INV_X1 U7081 ( .A(n6490), .ZN(n6136) );
  AOI22_X1 U7082 ( .A1(n6491), .A2(n6143), .B1(n6150), .B2(n6430), .ZN(n6135)
         );
  AOI22_X1 U7083 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n6145), .B1(n6492), 
        .B2(n6144), .ZN(n6134) );
  OAI211_X1 U7084 ( .C1(n6149), .C2(n6136), .A(n6135), .B(n6134), .ZN(U3064)
         );
  INV_X1 U7085 ( .A(n6496), .ZN(n6139) );
  AOI22_X1 U7086 ( .A1(n6497), .A2(n6143), .B1(n6150), .B2(n6434), .ZN(n6138)
         );
  AOI22_X1 U7087 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n6145), .B1(n6498), 
        .B2(n6144), .ZN(n6137) );
  OAI211_X1 U7088 ( .C1(n6149), .C2(n6139), .A(n6138), .B(n6137), .ZN(U3065)
         );
  INV_X1 U7089 ( .A(n6502), .ZN(n6142) );
  AOI22_X1 U7090 ( .A1(n6503), .A2(n6143), .B1(n6144), .B2(n6504), .ZN(n6141)
         );
  AOI22_X1 U7091 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n6145), .B1(n6395), 
        .B2(n6150), .ZN(n6140) );
  OAI211_X1 U7092 ( .C1(n6149), .C2(n6142), .A(n6141), .B(n6140), .ZN(U3066)
         );
  INV_X1 U7093 ( .A(n6627), .ZN(n6148) );
  AOI22_X1 U7094 ( .A1(n6625), .A2(n6143), .B1(n6150), .B2(n6444), .ZN(n6147)
         );
  AOI22_X1 U7095 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n6145), .B1(n6622), 
        .B2(n6144), .ZN(n6146) );
  OAI211_X1 U7096 ( .C1(n6149), .C2(n6148), .A(n6147), .B(n6146), .ZN(U3067)
         );
  NOR2_X1 U7097 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6187), .ZN(n6175)
         );
  NAND2_X1 U7098 ( .A1(n6152), .A2(n6151), .ZN(n6412) );
  NAND3_X1 U7099 ( .A1(n6407), .A2(n6406), .A3(n6415), .ZN(n6153) );
  OAI21_X1 U7100 ( .B1(n6154), .B2(n6412), .A(n6153), .ZN(n6174) );
  AOI22_X1 U7101 ( .A1(n6456), .A2(n6175), .B1(n6455), .B2(n6174), .ZN(n6161)
         );
  INV_X1 U7102 ( .A(n6175), .ZN(n6157) );
  NOR2_X2 U7103 ( .A1(n6182), .A2(n6268), .ZN(n6202) );
  INV_X1 U7104 ( .A(n6202), .ZN(n6211) );
  NAND3_X1 U7105 ( .A1(n6211), .A2(n6179), .A3(n6466), .ZN(n6155) );
  NOR2_X1 U7106 ( .A1(n6412), .A2(n6340), .ZN(n6183) );
  AOI21_X1 U7107 ( .B1(n6155), .B2(n6460), .A(n6183), .ZN(n6156) );
  AOI21_X1 U7108 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6157), .A(n6156), .ZN(
        n6159) );
  NOR2_X1 U7109 ( .A1(n6276), .A2(n6158), .ZN(n6417) );
  NAND3_X1 U7110 ( .A1(n6415), .A2(n6159), .A3(n6417), .ZN(n6176) );
  AOI22_X1 U7111 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n6176), .B1(n6418), 
        .B2(n6202), .ZN(n6160) );
  OAI211_X1 U7112 ( .C1(n6421), .C2(n6179), .A(n6161), .B(n6160), .ZN(U3068)
         );
  AOI22_X1 U7113 ( .A1(n6473), .A2(n6175), .B1(n6472), .B2(n6174), .ZN(n6163)
         );
  AOI22_X1 U7114 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n6176), .B1(n6348), 
        .B2(n6202), .ZN(n6162) );
  OAI211_X1 U7115 ( .C1(n6351), .C2(n6179), .A(n6163), .B(n6162), .ZN(U3069)
         );
  AOI22_X1 U7116 ( .A1(n6479), .A2(n6175), .B1(n6478), .B2(n6174), .ZN(n6165)
         );
  AOI22_X1 U7117 ( .A1(INSTQUEUE_REG_6__2__SCAN_IN), .A2(n6176), .B1(n6424), 
        .B2(n6202), .ZN(n6164) );
  OAI211_X1 U7118 ( .C1(n6427), .C2(n6179), .A(n6165), .B(n6164), .ZN(U3070)
         );
  AOI22_X1 U7119 ( .A1(n6485), .A2(n6175), .B1(n6484), .B2(n6174), .ZN(n6167)
         );
  AOI22_X1 U7120 ( .A1(INSTQUEUE_REG_6__3__SCAN_IN), .A2(n6176), .B1(n6387), 
        .B2(n6202), .ZN(n6166) );
  OAI211_X1 U7121 ( .C1(n6390), .C2(n6179), .A(n6167), .B(n6166), .ZN(U3071)
         );
  AOI22_X1 U7122 ( .A1(n6491), .A2(n6175), .B1(n6490), .B2(n6174), .ZN(n6169)
         );
  AOI22_X1 U7123 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n6176), .B1(n6430), 
        .B2(n6202), .ZN(n6168) );
  OAI211_X1 U7124 ( .C1(n6433), .C2(n6179), .A(n6169), .B(n6168), .ZN(U3072)
         );
  AOI22_X1 U7125 ( .A1(n6497), .A2(n6175), .B1(n6496), .B2(n6174), .ZN(n6171)
         );
  AOI22_X1 U7126 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n6176), .B1(n6434), 
        .B2(n6202), .ZN(n6170) );
  OAI211_X1 U7127 ( .C1(n6437), .C2(n6179), .A(n6171), .B(n6170), .ZN(U3073)
         );
  AOI22_X1 U7128 ( .A1(n6503), .A2(n6175), .B1(n6502), .B2(n6174), .ZN(n6173)
         );
  AOI22_X1 U7129 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(n6176), .B1(n6395), 
        .B2(n6202), .ZN(n6172) );
  OAI211_X1 U7130 ( .C1(n6399), .C2(n6179), .A(n6173), .B(n6172), .ZN(U3074)
         );
  AOI22_X1 U7131 ( .A1(n6625), .A2(n6175), .B1(n6627), .B2(n6174), .ZN(n6178)
         );
  AOI22_X1 U7132 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n6176), .B1(n6444), 
        .B2(n6202), .ZN(n6177) );
  OAI211_X1 U7133 ( .C1(n6449), .C2(n6179), .A(n6178), .B(n6177), .ZN(U3075)
         );
  NAND2_X1 U7134 ( .A1(n6180), .A2(n6299), .ZN(n6243) );
  INV_X1 U7135 ( .A(n6181), .ZN(n6206) );
  AOI22_X1 U7136 ( .A1(n6456), .A2(n6206), .B1(n6202), .B2(n6468), .ZN(n6191)
         );
  OAI21_X1 U7137 ( .B1(n6182), .B2(n6302), .A(n6466), .ZN(n6189) );
  INV_X1 U7138 ( .A(n6189), .ZN(n6184) );
  AOI21_X1 U7139 ( .B1(n6183), .B2(n6244), .A(n6206), .ZN(n6188) );
  NAND2_X1 U7140 ( .A1(n6184), .A2(n6188), .ZN(n6185) );
  OAI211_X1 U7141 ( .C1(n6466), .C2(n6186), .A(n6185), .B(n6465), .ZN(n6208)
         );
  OAI22_X1 U7142 ( .A1(n6189), .A2(n6188), .B1(n6187), .B2(n6799), .ZN(n6207)
         );
  AOI22_X1 U7143 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6208), .B1(n6455), 
        .B2(n6207), .ZN(n6190) );
  OAI211_X1 U7144 ( .C1(n6471), .C2(n6243), .A(n6191), .B(n6190), .ZN(U3076)
         );
  AOI22_X1 U7145 ( .A1(n6473), .A2(n6206), .B1(n6202), .B2(n6474), .ZN(n6193)
         );
  AOI22_X1 U7146 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6208), .B1(n6472), 
        .B2(n6207), .ZN(n6192) );
  OAI211_X1 U7147 ( .C1(n6477), .C2(n6243), .A(n6193), .B(n6192), .ZN(U3077)
         );
  AOI22_X1 U7148 ( .A1(n6479), .A2(n6206), .B1(n6202), .B2(n6480), .ZN(n6195)
         );
  AOI22_X1 U7149 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6208), .B1(n6478), 
        .B2(n6207), .ZN(n6194) );
  OAI211_X1 U7150 ( .C1(n6483), .C2(n6243), .A(n6195), .B(n6194), .ZN(U3078)
         );
  AOI22_X1 U7151 ( .A1(n6485), .A2(n6206), .B1(n6202), .B2(n6486), .ZN(n6197)
         );
  AOI22_X1 U7152 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6208), .B1(n6484), 
        .B2(n6207), .ZN(n6196) );
  OAI211_X1 U7153 ( .C1(n6489), .C2(n6243), .A(n6197), .B(n6196), .ZN(U3079)
         );
  INV_X1 U7154 ( .A(n6243), .ZN(n6205) );
  AOI22_X1 U7155 ( .A1(n6491), .A2(n6206), .B1(n6205), .B2(n6430), .ZN(n6199)
         );
  AOI22_X1 U7156 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6208), .B1(n6490), 
        .B2(n6207), .ZN(n6198) );
  OAI211_X1 U7157 ( .C1(n6433), .C2(n6211), .A(n6199), .B(n6198), .ZN(U3080)
         );
  AOI22_X1 U7158 ( .A1(n6497), .A2(n6206), .B1(n6202), .B2(n6498), .ZN(n6201)
         );
  AOI22_X1 U7159 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6208), .B1(n6496), 
        .B2(n6207), .ZN(n6200) );
  OAI211_X1 U7160 ( .C1(n6501), .C2(n6243), .A(n6201), .B(n6200), .ZN(U3081)
         );
  AOI22_X1 U7161 ( .A1(n6503), .A2(n6206), .B1(n6202), .B2(n6504), .ZN(n6204)
         );
  AOI22_X1 U7162 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6208), .B1(n6502), 
        .B2(n6207), .ZN(n6203) );
  OAI211_X1 U7163 ( .C1(n6507), .C2(n6243), .A(n6204), .B(n6203), .ZN(U3082)
         );
  AOI22_X1 U7164 ( .A1(n6625), .A2(n6206), .B1(n6205), .B2(n6444), .ZN(n6210)
         );
  AOI22_X1 U7165 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6208), .B1(n6627), 
        .B2(n6207), .ZN(n6209) );
  OAI211_X1 U7166 ( .C1(n6449), .C2(n6211), .A(n6210), .B(n6209), .ZN(U3083)
         );
  NAND3_X1 U7167 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6213), .A3(n6212), .ZN(n6249) );
  NOR2_X1 U7168 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6249), .ZN(n6239)
         );
  NAND2_X1 U7169 ( .A1(n6270), .A2(n6466), .ZN(n6409) );
  INV_X1 U7170 ( .A(n6214), .ZN(n6215) );
  OR2_X1 U7171 ( .A1(n6215), .A2(n6406), .ZN(n6336) );
  OAI22_X1 U7172 ( .A1(n6409), .A2(n6219), .B1(n6342), .B2(n6336), .ZN(n6238)
         );
  AOI22_X1 U7173 ( .A1(n6456), .A2(n6239), .B1(n6455), .B2(n6238), .ZN(n6225)
         );
  NAND2_X1 U7174 ( .A1(n6217), .A2(n6216), .ZN(n6303) );
  OR2_X1 U7175 ( .A1(n6303), .A2(n6218), .ZN(n6266) );
  NAND3_X1 U7176 ( .A1(n6266), .A2(n6466), .A3(n6243), .ZN(n6220) );
  INV_X1 U7177 ( .A(n6219), .ZN(n6245) );
  AOI22_X1 U7178 ( .A1(n6220), .A2(n6460), .B1(n6245), .B2(n6270), .ZN(n6223)
         );
  AOI21_X1 U7179 ( .B1(n6336), .B2(STATE2_REG_2__SCAN_IN), .A(n6221), .ZN(
        n6343) );
  OAI211_X1 U7180 ( .C1(n6600), .C2(n6239), .A(n6337), .B(n6343), .ZN(n6222)
         );
  AOI22_X1 U7181 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n6240), .B1(n6418), 
        .B2(n6623), .ZN(n6224) );
  OAI211_X1 U7182 ( .C1(n6421), .C2(n6243), .A(n6225), .B(n6224), .ZN(U3084)
         );
  AOI22_X1 U7183 ( .A1(n6473), .A2(n6239), .B1(n6472), .B2(n6238), .ZN(n6227)
         );
  AOI22_X1 U7184 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n6240), .B1(n6348), 
        .B2(n6623), .ZN(n6226) );
  OAI211_X1 U7185 ( .C1(n6351), .C2(n6243), .A(n6227), .B(n6226), .ZN(U3085)
         );
  AOI22_X1 U7186 ( .A1(n6479), .A2(n6239), .B1(n6478), .B2(n6238), .ZN(n6229)
         );
  AOI22_X1 U7187 ( .A1(INSTQUEUE_REG_8__2__SCAN_IN), .A2(n6240), .B1(n6424), 
        .B2(n6623), .ZN(n6228) );
  OAI211_X1 U7188 ( .C1(n6427), .C2(n6243), .A(n6229), .B(n6228), .ZN(U3086)
         );
  AOI22_X1 U7189 ( .A1(n6485), .A2(n6239), .B1(n6484), .B2(n6238), .ZN(n6231)
         );
  AOI22_X1 U7190 ( .A1(INSTQUEUE_REG_8__3__SCAN_IN), .A2(n6240), .B1(n6387), 
        .B2(n6623), .ZN(n6230) );
  OAI211_X1 U7191 ( .C1(n6390), .C2(n6243), .A(n6231), .B(n6230), .ZN(U3087)
         );
  AOI22_X1 U7192 ( .A1(n6491), .A2(n6239), .B1(n6490), .B2(n6238), .ZN(n6233)
         );
  AOI22_X1 U7193 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n6240), .B1(n6430), 
        .B2(n6623), .ZN(n6232) );
  OAI211_X1 U7194 ( .C1(n6433), .C2(n6243), .A(n6233), .B(n6232), .ZN(U3088)
         );
  AOI22_X1 U7195 ( .A1(n6497), .A2(n6239), .B1(n6496), .B2(n6238), .ZN(n6235)
         );
  AOI22_X1 U7196 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n6240), .B1(n6434), 
        .B2(n6623), .ZN(n6234) );
  OAI211_X1 U7197 ( .C1(n6437), .C2(n6243), .A(n6235), .B(n6234), .ZN(U3089)
         );
  AOI22_X1 U7198 ( .A1(n6503), .A2(n6239), .B1(n6502), .B2(n6238), .ZN(n6237)
         );
  AOI22_X1 U7199 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(n6240), .B1(n6395), 
        .B2(n6623), .ZN(n6236) );
  OAI211_X1 U7200 ( .C1(n6399), .C2(n6243), .A(n6237), .B(n6236), .ZN(U3090)
         );
  AOI22_X1 U7201 ( .A1(n6625), .A2(n6239), .B1(n6627), .B2(n6238), .ZN(n6242)
         );
  AOI22_X1 U7202 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n6240), .B1(n6444), 
        .B2(n6623), .ZN(n6241) );
  OAI211_X1 U7203 ( .C1(n6449), .C2(n6243), .A(n6242), .B(n6241), .ZN(U3091)
         );
  NOR2_X1 U7204 ( .A1(n6370), .A2(n6249), .ZN(n6624) );
  AOI22_X1 U7205 ( .A1(n6456), .A2(n6624), .B1(n6291), .B2(n6418), .ZN(n6253)
         );
  AND2_X1 U7206 ( .A1(n6270), .A2(n6244), .ZN(n6451) );
  AOI21_X1 U7207 ( .B1(n6451), .B2(n6245), .A(n6624), .ZN(n6250) );
  AOI21_X1 U7208 ( .B1(n6303), .B2(n6466), .A(n6246), .ZN(n6251) );
  INV_X1 U7209 ( .A(n6251), .ZN(n6247) );
  AOI22_X1 U7210 ( .A1(n6250), .A2(n6247), .B1(n6454), .B2(n6249), .ZN(n6248)
         );
  NAND2_X1 U7211 ( .A1(n6465), .A2(n6248), .ZN(n6628) );
  OAI22_X1 U7212 ( .A1(n6251), .A2(n6250), .B1(n6799), .B2(n6249), .ZN(n6626)
         );
  AOI22_X1 U7213 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n6628), .B1(n6455), 
        .B2(n6626), .ZN(n6252) );
  OAI211_X1 U7214 ( .C1(n6421), .C2(n6266), .A(n6253), .B(n6252), .ZN(U3092)
         );
  AOI22_X1 U7215 ( .A1(n6473), .A2(n6624), .B1(n6291), .B2(n6348), .ZN(n6255)
         );
  AOI22_X1 U7216 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n6628), .B1(n6472), 
        .B2(n6626), .ZN(n6254) );
  OAI211_X1 U7217 ( .C1(n6351), .C2(n6266), .A(n6255), .B(n6254), .ZN(U3093)
         );
  AOI22_X1 U7218 ( .A1(n6479), .A2(n6624), .B1(n6623), .B2(n6480), .ZN(n6257)
         );
  AOI22_X1 U7219 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n6628), .B1(n6478), 
        .B2(n6626), .ZN(n6256) );
  OAI211_X1 U7220 ( .C1(n6483), .C2(n6631), .A(n6257), .B(n6256), .ZN(U3094)
         );
  AOI22_X1 U7221 ( .A1(n6485), .A2(n6624), .B1(n6291), .B2(n6387), .ZN(n6259)
         );
  AOI22_X1 U7222 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n6628), .B1(n6484), 
        .B2(n6626), .ZN(n6258) );
  OAI211_X1 U7223 ( .C1(n6390), .C2(n6266), .A(n6259), .B(n6258), .ZN(U3095)
         );
  AOI22_X1 U7224 ( .A1(n6491), .A2(n6624), .B1(n6623), .B2(n6492), .ZN(n6261)
         );
  AOI22_X1 U7225 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n6628), .B1(n6490), 
        .B2(n6626), .ZN(n6260) );
  OAI211_X1 U7226 ( .C1(n6495), .C2(n6631), .A(n6261), .B(n6260), .ZN(U3096)
         );
  AOI22_X1 U7227 ( .A1(n6497), .A2(n6624), .B1(n6291), .B2(n6434), .ZN(n6263)
         );
  AOI22_X1 U7228 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n6628), .B1(n6496), 
        .B2(n6626), .ZN(n6262) );
  OAI211_X1 U7229 ( .C1(n6437), .C2(n6266), .A(n6263), .B(n6262), .ZN(U3097)
         );
  AOI22_X1 U7230 ( .A1(n6503), .A2(n6624), .B1(n6291), .B2(n6395), .ZN(n6265)
         );
  AOI22_X1 U7231 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n6628), .B1(n6502), 
        .B2(n6626), .ZN(n6264) );
  OAI211_X1 U7232 ( .C1(n6399), .C2(n6266), .A(n6265), .B(n6264), .ZN(U3098)
         );
  NAND2_X1 U7233 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6267), .ZN(n6311) );
  NOR2_X1 U7234 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6311), .ZN(n6294)
         );
  OR2_X1 U7235 ( .A1(n6303), .A2(n6268), .ZN(n6335) );
  AOI22_X1 U7236 ( .A1(n6456), .A2(n6294), .B1(n6324), .B2(n6418), .ZN(n6280)
         );
  NAND2_X1 U7237 ( .A1(n6335), .A2(n6631), .ZN(n6269) );
  AOI21_X1 U7238 ( .B1(n6269), .B2(STATEBS16_REG_SCAN_IN), .A(n6454), .ZN(
        n6275) );
  NAND2_X1 U7239 ( .A1(n6271), .A2(n6270), .ZN(n6305) );
  INV_X1 U7240 ( .A(n6294), .ZN(n6272) );
  AOI22_X1 U7241 ( .A1(n6275), .A2(n6305), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n6272), .ZN(n6273) );
  OAI211_X1 U7242 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6799), .A(n6274), .B(n6273), .ZN(n6296) );
  INV_X1 U7243 ( .A(n6275), .ZN(n6278) );
  NAND3_X1 U7244 ( .A1(n6276), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6406), .ZN(n6277) );
  OAI21_X1 U7245 ( .B1(n6278), .B2(n6305), .A(n6277), .ZN(n6295) );
  AOI22_X1 U7246 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n6296), .B1(n6455), 
        .B2(n6295), .ZN(n6279) );
  OAI211_X1 U7247 ( .C1(n6421), .C2(n6631), .A(n6280), .B(n6279), .ZN(U3100)
         );
  AOI22_X1 U7248 ( .A1(n6473), .A2(n6294), .B1(n6291), .B2(n6474), .ZN(n6282)
         );
  AOI22_X1 U7249 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n6296), .B1(n6472), 
        .B2(n6295), .ZN(n6281) );
  OAI211_X1 U7250 ( .C1(n6477), .C2(n6335), .A(n6282), .B(n6281), .ZN(U3101)
         );
  AOI22_X1 U7251 ( .A1(n6479), .A2(n6294), .B1(n6324), .B2(n6424), .ZN(n6284)
         );
  AOI22_X1 U7252 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(n6296), .B1(n6478), 
        .B2(n6295), .ZN(n6283) );
  OAI211_X1 U7253 ( .C1(n6427), .C2(n6631), .A(n6284), .B(n6283), .ZN(U3102)
         );
  AOI22_X1 U7254 ( .A1(n6485), .A2(n6294), .B1(n6324), .B2(n6387), .ZN(n6286)
         );
  AOI22_X1 U7255 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(n6296), .B1(n6484), 
        .B2(n6295), .ZN(n6285) );
  OAI211_X1 U7256 ( .C1(n6390), .C2(n6631), .A(n6286), .B(n6285), .ZN(U3103)
         );
  AOI22_X1 U7257 ( .A1(n6491), .A2(n6294), .B1(n6291), .B2(n6492), .ZN(n6288)
         );
  AOI22_X1 U7258 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n6296), .B1(n6490), 
        .B2(n6295), .ZN(n6287) );
  OAI211_X1 U7259 ( .C1(n6495), .C2(n6335), .A(n6288), .B(n6287), .ZN(U3104)
         );
  AOI22_X1 U7260 ( .A1(n6497), .A2(n6294), .B1(n6324), .B2(n6434), .ZN(n6290)
         );
  AOI22_X1 U7261 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n6296), .B1(n6496), 
        .B2(n6295), .ZN(n6289) );
  OAI211_X1 U7262 ( .C1(n6437), .C2(n6631), .A(n6290), .B(n6289), .ZN(U3105)
         );
  AOI22_X1 U7263 ( .A1(n6503), .A2(n6294), .B1(n6291), .B2(n6504), .ZN(n6293)
         );
  AOI22_X1 U7264 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n6296), .B1(n6502), 
        .B2(n6295), .ZN(n6292) );
  OAI211_X1 U7265 ( .C1(n6507), .C2(n6335), .A(n6293), .B(n6292), .ZN(U3106)
         );
  AOI22_X1 U7266 ( .A1(n6625), .A2(n6294), .B1(n6324), .B2(n6444), .ZN(n6298)
         );
  AOI22_X1 U7267 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n6296), .B1(n6627), 
        .B2(n6295), .ZN(n6297) );
  OAI211_X1 U7268 ( .C1(n6449), .C2(n6631), .A(n6298), .B(n6297), .ZN(U3107)
         );
  INV_X1 U7269 ( .A(n6303), .ZN(n6300) );
  NAND2_X1 U7270 ( .A1(n6300), .A2(n6299), .ZN(n6367) );
  NOR2_X1 U7271 ( .A1(n6415), .A2(n6301), .ZN(n6330) );
  AOI22_X1 U7272 ( .A1(n6456), .A2(n6330), .B1(n6324), .B2(n6468), .ZN(n6315)
         );
  INV_X1 U7273 ( .A(n6311), .ZN(n6309) );
  OAI21_X1 U7274 ( .B1(n6303), .B2(n6302), .A(n6466), .ZN(n6313) );
  OR2_X1 U7275 ( .A1(n6305), .A2(n6304), .ZN(n6307) );
  INV_X1 U7276 ( .A(n6330), .ZN(n6306) );
  NAND2_X1 U7277 ( .A1(n6307), .A2(n6306), .ZN(n6310) );
  OR2_X1 U7278 ( .A1(n6313), .A2(n6310), .ZN(n6308) );
  OAI211_X1 U7279 ( .C1(n6466), .C2(n6309), .A(n6308), .B(n6465), .ZN(n6332)
         );
  INV_X1 U7280 ( .A(n6310), .ZN(n6312) );
  OAI22_X1 U7281 ( .A1(n6313), .A2(n6312), .B1(n6311), .B2(n6799), .ZN(n6331)
         );
  AOI22_X1 U7282 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6332), .B1(n6455), 
        .B2(n6331), .ZN(n6314) );
  OAI211_X1 U7283 ( .C1(n6471), .C2(n6367), .A(n6315), .B(n6314), .ZN(U3108)
         );
  AOI22_X1 U7284 ( .A1(n6473), .A2(n6330), .B1(n6324), .B2(n6474), .ZN(n6317)
         );
  AOI22_X1 U7285 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6332), .B1(n6472), 
        .B2(n6331), .ZN(n6316) );
  OAI211_X1 U7286 ( .C1(n6477), .C2(n6367), .A(n6317), .B(n6316), .ZN(U3109)
         );
  INV_X1 U7287 ( .A(n6367), .ZN(n6329) );
  AOI22_X1 U7288 ( .A1(n6479), .A2(n6330), .B1(n6329), .B2(n6424), .ZN(n6319)
         );
  AOI22_X1 U7289 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6332), .B1(n6478), 
        .B2(n6331), .ZN(n6318) );
  OAI211_X1 U7290 ( .C1(n6427), .C2(n6335), .A(n6319), .B(n6318), .ZN(U3110)
         );
  AOI22_X1 U7291 ( .A1(n6485), .A2(n6330), .B1(n6324), .B2(n6486), .ZN(n6321)
         );
  AOI22_X1 U7292 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6332), .B1(n6484), 
        .B2(n6331), .ZN(n6320) );
  OAI211_X1 U7293 ( .C1(n6489), .C2(n6367), .A(n6321), .B(n6320), .ZN(U3111)
         );
  AOI22_X1 U7294 ( .A1(n6491), .A2(n6330), .B1(n6324), .B2(n6492), .ZN(n6323)
         );
  AOI22_X1 U7295 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6332), .B1(n6490), 
        .B2(n6331), .ZN(n6322) );
  OAI211_X1 U7296 ( .C1(n6495), .C2(n6367), .A(n6323), .B(n6322), .ZN(U3112)
         );
  AOI22_X1 U7297 ( .A1(n6497), .A2(n6330), .B1(n6324), .B2(n6498), .ZN(n6326)
         );
  AOI22_X1 U7298 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6332), .B1(n6496), 
        .B2(n6331), .ZN(n6325) );
  OAI211_X1 U7299 ( .C1(n6501), .C2(n6367), .A(n6326), .B(n6325), .ZN(U3113)
         );
  AOI22_X1 U7300 ( .A1(n6503), .A2(n6330), .B1(n6329), .B2(n6395), .ZN(n6328)
         );
  AOI22_X1 U7301 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6332), .B1(n6502), 
        .B2(n6331), .ZN(n6327) );
  OAI211_X1 U7302 ( .C1(n6399), .C2(n6335), .A(n6328), .B(n6327), .ZN(U3114)
         );
  AOI22_X1 U7303 ( .A1(n6625), .A2(n6330), .B1(n6329), .B2(n6444), .ZN(n6334)
         );
  AOI22_X1 U7304 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6332), .B1(n6627), 
        .B2(n6331), .ZN(n6333) );
  OAI211_X1 U7305 ( .C1(n6449), .C2(n6335), .A(n6334), .B(n6333), .ZN(U3115)
         );
  OR2_X1 U7306 ( .A1(n6415), .A2(n6378), .ZN(n6374) );
  NOR2_X1 U7307 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6374), .ZN(n6363)
         );
  OAI22_X1 U7308 ( .A1(n6338), .A2(n6409), .B1(n6337), .B2(n6336), .ZN(n6362)
         );
  AOI22_X1 U7309 ( .A1(n6456), .A2(n6363), .B1(n6455), .B2(n6362), .ZN(n6347)
         );
  NAND3_X1 U7310 ( .A1(n6398), .A2(n6367), .A3(n6466), .ZN(n6341) );
  AOI22_X1 U7311 ( .A1(n6341), .A2(n6460), .B1(n6371), .B2(n6340), .ZN(n6345)
         );
  OAI211_X1 U7312 ( .C1(n6363), .C2(n6600), .A(n6343), .B(n6342), .ZN(n6344)
         );
  AOI22_X1 U7313 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n6364), .B1(n6418), 
        .B2(n6400), .ZN(n6346) );
  OAI211_X1 U7314 ( .C1(n6421), .C2(n6367), .A(n6347), .B(n6346), .ZN(U3116)
         );
  AOI22_X1 U7315 ( .A1(n6473), .A2(n6363), .B1(n6472), .B2(n6362), .ZN(n6350)
         );
  AOI22_X1 U7316 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n6364), .B1(n6348), 
        .B2(n6400), .ZN(n6349) );
  OAI211_X1 U7317 ( .C1(n6351), .C2(n6367), .A(n6350), .B(n6349), .ZN(U3117)
         );
  AOI22_X1 U7318 ( .A1(n6479), .A2(n6363), .B1(n6478), .B2(n6362), .ZN(n6353)
         );
  AOI22_X1 U7319 ( .A1(INSTQUEUE_REG_12__2__SCAN_IN), .A2(n6364), .B1(n6424), 
        .B2(n6400), .ZN(n6352) );
  OAI211_X1 U7320 ( .C1(n6427), .C2(n6367), .A(n6353), .B(n6352), .ZN(U3118)
         );
  AOI22_X1 U7321 ( .A1(n6485), .A2(n6363), .B1(n6484), .B2(n6362), .ZN(n6355)
         );
  AOI22_X1 U7322 ( .A1(INSTQUEUE_REG_12__3__SCAN_IN), .A2(n6364), .B1(n6387), 
        .B2(n6400), .ZN(n6354) );
  OAI211_X1 U7323 ( .C1(n6390), .C2(n6367), .A(n6355), .B(n6354), .ZN(U3119)
         );
  AOI22_X1 U7324 ( .A1(n6491), .A2(n6363), .B1(n6490), .B2(n6362), .ZN(n6357)
         );
  AOI22_X1 U7325 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n6364), .B1(n6430), 
        .B2(n6400), .ZN(n6356) );
  OAI211_X1 U7326 ( .C1(n6433), .C2(n6367), .A(n6357), .B(n6356), .ZN(U3120)
         );
  AOI22_X1 U7327 ( .A1(n6497), .A2(n6363), .B1(n6496), .B2(n6362), .ZN(n6359)
         );
  AOI22_X1 U7328 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n6364), .B1(n6434), 
        .B2(n6400), .ZN(n6358) );
  OAI211_X1 U7329 ( .C1(n6437), .C2(n6367), .A(n6359), .B(n6358), .ZN(U3121)
         );
  AOI22_X1 U7330 ( .A1(n6503), .A2(n6363), .B1(n6502), .B2(n6362), .ZN(n6361)
         );
  AOI22_X1 U7331 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(n6364), .B1(n6395), 
        .B2(n6400), .ZN(n6360) );
  OAI211_X1 U7332 ( .C1(n6399), .C2(n6367), .A(n6361), .B(n6360), .ZN(U3122)
         );
  AOI22_X1 U7333 ( .A1(n6625), .A2(n6363), .B1(n6627), .B2(n6362), .ZN(n6366)
         );
  AOI22_X1 U7334 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n6364), .B1(n6444), 
        .B2(n6400), .ZN(n6365) );
  OAI211_X1 U7335 ( .C1(n6449), .C2(n6367), .A(n6366), .B(n6365), .ZN(U3123)
         );
  INV_X1 U7336 ( .A(n6368), .ZN(n6369) );
  NOR2_X1 U7337 ( .A1(n6370), .A2(n6374), .ZN(n6401) );
  AOI22_X1 U7338 ( .A1(n6456), .A2(n6401), .B1(n6400), .B2(n6468), .ZN(n6382)
         );
  AOI21_X1 U7339 ( .B1(n6451), .B2(n6371), .A(n6401), .ZN(n6379) );
  OR2_X1 U7340 ( .A1(n6459), .A2(n6454), .ZN(n6373) );
  AND2_X1 U7341 ( .A1(n6373), .A2(n6372), .ZN(n6380) );
  INV_X1 U7342 ( .A(n6380), .ZN(n6375) );
  AOI22_X1 U7343 ( .A1(n6379), .A2(n6375), .B1(n6454), .B2(n6374), .ZN(n6376)
         );
  NAND2_X1 U7344 ( .A1(n6465), .A2(n6376), .ZN(n6403) );
  NAND2_X1 U7345 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        STATE2_REG_2__SCAN_IN), .ZN(n6377) );
  OAI22_X1 U7346 ( .A1(n6380), .A2(n6379), .B1(n6378), .B2(n6377), .ZN(n6402)
         );
  AOI22_X1 U7347 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n6403), .B1(n6455), 
        .B2(n6402), .ZN(n6381) );
  OAI211_X1 U7348 ( .C1(n6471), .C2(n6448), .A(n6382), .B(n6381), .ZN(U3124)
         );
  AOI22_X1 U7349 ( .A1(n6473), .A2(n6401), .B1(n6400), .B2(n6474), .ZN(n6384)
         );
  AOI22_X1 U7350 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n6403), .B1(n6472), 
        .B2(n6402), .ZN(n6383) );
  OAI211_X1 U7351 ( .C1(n6477), .C2(n6448), .A(n6384), .B(n6383), .ZN(U3125)
         );
  AOI22_X1 U7352 ( .A1(n6479), .A2(n6401), .B1(n6438), .B2(n6424), .ZN(n6386)
         );
  AOI22_X1 U7353 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n6403), .B1(n6478), 
        .B2(n6402), .ZN(n6385) );
  OAI211_X1 U7354 ( .C1(n6427), .C2(n6398), .A(n6386), .B(n6385), .ZN(U3126)
         );
  AOI22_X1 U7355 ( .A1(n6485), .A2(n6401), .B1(n6438), .B2(n6387), .ZN(n6389)
         );
  AOI22_X1 U7356 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n6403), .B1(n6484), 
        .B2(n6402), .ZN(n6388) );
  OAI211_X1 U7357 ( .C1(n6390), .C2(n6398), .A(n6389), .B(n6388), .ZN(U3127)
         );
  AOI22_X1 U7358 ( .A1(n6491), .A2(n6401), .B1(n6400), .B2(n6492), .ZN(n6392)
         );
  AOI22_X1 U7359 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n6403), .B1(n6490), 
        .B2(n6402), .ZN(n6391) );
  OAI211_X1 U7360 ( .C1(n6495), .C2(n6448), .A(n6392), .B(n6391), .ZN(U3128)
         );
  AOI22_X1 U7361 ( .A1(n6497), .A2(n6401), .B1(n6438), .B2(n6434), .ZN(n6394)
         );
  AOI22_X1 U7362 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n6403), .B1(n6496), 
        .B2(n6402), .ZN(n6393) );
  OAI211_X1 U7363 ( .C1(n6437), .C2(n6398), .A(n6394), .B(n6393), .ZN(U3129)
         );
  AOI22_X1 U7364 ( .A1(n6503), .A2(n6401), .B1(n6438), .B2(n6395), .ZN(n6397)
         );
  AOI22_X1 U7365 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n6403), .B1(n6502), 
        .B2(n6402), .ZN(n6396) );
  OAI211_X1 U7366 ( .C1(n6399), .C2(n6398), .A(n6397), .B(n6396), .ZN(U3130)
         );
  AOI22_X1 U7367 ( .A1(n6625), .A2(n6401), .B1(n6400), .B2(n6622), .ZN(n6405)
         );
  AOI22_X1 U7368 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n6403), .B1(n6627), 
        .B2(n6402), .ZN(n6404) );
  OAI211_X1 U7369 ( .C1(n6632), .C2(n6448), .A(n6405), .B(n6404), .ZN(U3131)
         );
  NOR2_X1 U7370 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6453), .ZN(n6443)
         );
  NAND3_X1 U7371 ( .A1(n6407), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6406), .ZN(n6408) );
  OAI21_X1 U7372 ( .B1(n6409), .B2(n6412), .A(n6408), .ZN(n6442) );
  AOI22_X1 U7373 ( .A1(n6456), .A2(n6443), .B1(n6455), .B2(n6442), .ZN(n6420)
         );
  NAND2_X1 U7374 ( .A1(n6459), .A2(n6410), .ZN(n6441) );
  AOI21_X1 U7375 ( .B1(n6448), .B2(n6441), .A(n6411), .ZN(n6413) );
  INV_X1 U7376 ( .A(n6412), .ZN(n6452) );
  NOR3_X1 U7377 ( .A1(n6413), .A2(n6452), .A3(n6454), .ZN(n6414) );
  NOR2_X1 U7378 ( .A1(n6415), .A2(n6414), .ZN(n6416) );
  OAI211_X1 U7379 ( .C1(n6443), .C2(n6600), .A(n6417), .B(n6416), .ZN(n6445)
         );
  AOI22_X1 U7380 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n6445), .B1(n6418), 
        .B2(n6510), .ZN(n6419) );
  OAI211_X1 U7381 ( .C1(n6421), .C2(n6448), .A(n6420), .B(n6419), .ZN(U3132)
         );
  AOI22_X1 U7382 ( .A1(n6473), .A2(n6443), .B1(n6472), .B2(n6442), .ZN(n6423)
         );
  AOI22_X1 U7383 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n6445), .B1(n6474), 
        .B2(n6438), .ZN(n6422) );
  OAI211_X1 U7384 ( .C1(n6477), .C2(n6441), .A(n6423), .B(n6422), .ZN(U3133)
         );
  AOI22_X1 U7385 ( .A1(n6479), .A2(n6443), .B1(n6478), .B2(n6442), .ZN(n6426)
         );
  AOI22_X1 U7386 ( .A1(INSTQUEUE_REG_14__2__SCAN_IN), .A2(n6445), .B1(n6424), 
        .B2(n6510), .ZN(n6425) );
  OAI211_X1 U7387 ( .C1(n6427), .C2(n6448), .A(n6426), .B(n6425), .ZN(U3134)
         );
  AOI22_X1 U7388 ( .A1(n6485), .A2(n6443), .B1(n6484), .B2(n6442), .ZN(n6429)
         );
  AOI22_X1 U7389 ( .A1(INSTQUEUE_REG_14__3__SCAN_IN), .A2(n6445), .B1(n6486), 
        .B2(n6438), .ZN(n6428) );
  OAI211_X1 U7390 ( .C1(n6489), .C2(n6441), .A(n6429), .B(n6428), .ZN(U3135)
         );
  AOI22_X1 U7391 ( .A1(n6491), .A2(n6443), .B1(n6490), .B2(n6442), .ZN(n6432)
         );
  AOI22_X1 U7392 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n6445), .B1(n6430), 
        .B2(n6510), .ZN(n6431) );
  OAI211_X1 U7393 ( .C1(n6433), .C2(n6448), .A(n6432), .B(n6431), .ZN(U3136)
         );
  AOI22_X1 U7394 ( .A1(n6497), .A2(n6443), .B1(n6496), .B2(n6442), .ZN(n6436)
         );
  AOI22_X1 U7395 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n6445), .B1(n6434), 
        .B2(n6510), .ZN(n6435) );
  OAI211_X1 U7396 ( .C1(n6437), .C2(n6448), .A(n6436), .B(n6435), .ZN(U3137)
         );
  AOI22_X1 U7397 ( .A1(n6503), .A2(n6443), .B1(n6502), .B2(n6442), .ZN(n6440)
         );
  AOI22_X1 U7398 ( .A1(INSTQUEUE_REG_14__6__SCAN_IN), .A2(n6445), .B1(n6504), 
        .B2(n6438), .ZN(n6439) );
  OAI211_X1 U7399 ( .C1(n6507), .C2(n6441), .A(n6440), .B(n6439), .ZN(U3138)
         );
  AOI22_X1 U7400 ( .A1(n6625), .A2(n6443), .B1(n6627), .B2(n6442), .ZN(n6447)
         );
  AOI22_X1 U7401 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n6445), .B1(n6444), 
        .B2(n6510), .ZN(n6446) );
  OAI211_X1 U7402 ( .C1(n6449), .C2(n6448), .A(n6447), .B(n6446), .ZN(U3139)
         );
  INV_X1 U7403 ( .A(n6450), .ZN(n6509) );
  AOI21_X1 U7404 ( .B1(n6452), .B2(n6451), .A(n6509), .ZN(n6461) );
  OAI22_X1 U7405 ( .A1(n6461), .A2(n6454), .B1(n6453), .B2(n6799), .ZN(n6508)
         );
  AOI22_X1 U7406 ( .A1(n6456), .A2(n6509), .B1(n6455), .B2(n6508), .ZN(n6470)
         );
  AOI21_X1 U7407 ( .B1(n6459), .B2(n6458), .A(n6457), .ZN(n6463) );
  INV_X1 U7408 ( .A(n6460), .ZN(n6462) );
  OAI21_X1 U7409 ( .B1(n6463), .B2(n6462), .A(n6461), .ZN(n6464) );
  OAI211_X1 U7410 ( .C1(n6467), .C2(n6466), .A(n6465), .B(n6464), .ZN(n6511)
         );
  AOI22_X1 U7411 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6511), .B1(n6468), 
        .B2(n6510), .ZN(n6469) );
  OAI211_X1 U7412 ( .C1(n6471), .C2(n6514), .A(n6470), .B(n6469), .ZN(U3140)
         );
  AOI22_X1 U7413 ( .A1(n6473), .A2(n6509), .B1(n6472), .B2(n6508), .ZN(n6476)
         );
  AOI22_X1 U7414 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6511), .B1(n6474), 
        .B2(n6510), .ZN(n6475) );
  OAI211_X1 U7415 ( .C1(n6477), .C2(n6514), .A(n6476), .B(n6475), .ZN(U3141)
         );
  AOI22_X1 U7416 ( .A1(n6479), .A2(n6509), .B1(n6478), .B2(n6508), .ZN(n6482)
         );
  AOI22_X1 U7417 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6511), .B1(n6480), 
        .B2(n6510), .ZN(n6481) );
  OAI211_X1 U7418 ( .C1(n6483), .C2(n6514), .A(n6482), .B(n6481), .ZN(U3142)
         );
  AOI22_X1 U7419 ( .A1(n6485), .A2(n6509), .B1(n6484), .B2(n6508), .ZN(n6488)
         );
  AOI22_X1 U7420 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6511), .B1(n6486), 
        .B2(n6510), .ZN(n6487) );
  OAI211_X1 U7421 ( .C1(n6489), .C2(n6514), .A(n6488), .B(n6487), .ZN(U3143)
         );
  AOI22_X1 U7422 ( .A1(n6491), .A2(n6509), .B1(n6490), .B2(n6508), .ZN(n6494)
         );
  AOI22_X1 U7423 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6511), .B1(n6492), 
        .B2(n6510), .ZN(n6493) );
  OAI211_X1 U7424 ( .C1(n6495), .C2(n6514), .A(n6494), .B(n6493), .ZN(U3144)
         );
  AOI22_X1 U7425 ( .A1(n6497), .A2(n6509), .B1(n6496), .B2(n6508), .ZN(n6500)
         );
  AOI22_X1 U7426 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6511), .B1(n6498), 
        .B2(n6510), .ZN(n6499) );
  OAI211_X1 U7427 ( .C1(n6501), .C2(n6514), .A(n6500), .B(n6499), .ZN(U3145)
         );
  AOI22_X1 U7428 ( .A1(n6503), .A2(n6509), .B1(n6502), .B2(n6508), .ZN(n6506)
         );
  AOI22_X1 U7429 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6511), .B1(n6504), 
        .B2(n6510), .ZN(n6505) );
  OAI211_X1 U7430 ( .C1(n6507), .C2(n6514), .A(n6506), .B(n6505), .ZN(U3146)
         );
  AOI22_X1 U7431 ( .A1(n6625), .A2(n6509), .B1(n6627), .B2(n6508), .ZN(n6513)
         );
  AOI22_X1 U7432 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6511), .B1(n6622), 
        .B2(n6510), .ZN(n6512) );
  OAI211_X1 U7433 ( .C1(n6632), .C2(n6514), .A(n6513), .B(n6512), .ZN(U3147)
         );
  AOI21_X1 U7434 ( .B1(n6516), .B2(n6612), .A(n6515), .ZN(n6520) );
  NAND2_X1 U7435 ( .A1(n6517), .A2(n6799), .ZN(n6522) );
  OAI211_X1 U7436 ( .C1(n6597), .C2(n6525), .A(STATE2_REG_1__SCAN_IN), .B(
        n6522), .ZN(n6518) );
  OAI211_X1 U7437 ( .C1(n6597), .C2(n6520), .A(n6519), .B(n6518), .ZN(U3149)
         );
  NAND3_X1 U7438 ( .A1(n6522), .A2(n6521), .A3(n6598), .ZN(n6524) );
  OAI21_X1 U7439 ( .B1(n6525), .B2(n6524), .A(n6523), .ZN(U3150) );
  INV_X1 U7440 ( .A(n6596), .ZN(n6592) );
  AND2_X1 U7441 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6592), .ZN(U3151) );
  AND2_X1 U7442 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6592), .ZN(U3152) );
  AND2_X1 U7443 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6592), .ZN(U3153) );
  INV_X1 U7444 ( .A(DATAWIDTH_REG_28__SCAN_IN), .ZN(n6868) );
  NOR2_X1 U7445 ( .A1(n6596), .A2(n6868), .ZN(U3154) );
  INV_X1 U7446 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6909) );
  NOR2_X1 U7447 ( .A1(n6596), .A2(n6909), .ZN(U3155) );
  AND2_X1 U7448 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6592), .ZN(U3156) );
  AND2_X1 U7449 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6592), .ZN(U3157) );
  INV_X1 U7450 ( .A(DATAWIDTH_REG_24__SCAN_IN), .ZN(n6940) );
  NOR2_X1 U7451 ( .A1(n6596), .A2(n6940), .ZN(U3158) );
  AND2_X1 U7452 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6592), .ZN(U3159) );
  AND2_X1 U7453 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6592), .ZN(U3160) );
  AND2_X1 U7454 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6592), .ZN(U3161) );
  AND2_X1 U7455 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6592), .ZN(U3162) );
  AND2_X1 U7456 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6592), .ZN(U3163) );
  INV_X1 U7457 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n6855) );
  NOR2_X1 U7458 ( .A1(n6596), .A2(n6855), .ZN(U3164) );
  AND2_X1 U7459 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6592), .ZN(U3165) );
  AND2_X1 U7460 ( .A1(n6592), .A2(DATAWIDTH_REG_16__SCAN_IN), .ZN(U3166) );
  INV_X1 U7461 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6937) );
  NOR2_X1 U7462 ( .A1(n6596), .A2(n6937), .ZN(U3167) );
  AND2_X1 U7463 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6592), .ZN(U3168) );
  AND2_X1 U7464 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6592), .ZN(U3169) );
  AND2_X1 U7465 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6592), .ZN(U3170) );
  AND2_X1 U7466 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6592), .ZN(U3171) );
  INV_X1 U7467 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6966) );
  NOR2_X1 U7468 ( .A1(n6596), .A2(n6966), .ZN(U3172) );
  AND2_X1 U7469 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6592), .ZN(U3173) );
  AND2_X1 U7470 ( .A1(n6592), .A2(DATAWIDTH_REG_8__SCAN_IN), .ZN(U3174) );
  AND2_X1 U7471 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6592), .ZN(U3175) );
  AND2_X1 U7472 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6592), .ZN(U3176) );
  AND2_X1 U7473 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6592), .ZN(U3177) );
  AND2_X1 U7474 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6592), .ZN(U3178) );
  AND2_X1 U7475 ( .A1(n6592), .A2(DATAWIDTH_REG_3__SCAN_IN), .ZN(U3179) );
  AND2_X1 U7476 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6592), .ZN(U3180) );
  INV_X1 U7477 ( .A(n6543), .ZN(n6529) );
  AOI22_X1 U7478 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6544) );
  AND2_X1 U7479 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6530) );
  INV_X1 U7480 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6526) );
  OAI21_X1 U7481 ( .B1(n6530), .B2(n6526), .A(n6609), .ZN(n6528) );
  OAI221_X1 U7482 ( .B1(n6545), .B2(NA_N), .C1(n6545), .C2(n6535), .A(n6527), 
        .ZN(n6540) );
  OAI211_X1 U7483 ( .C1(n6529), .C2(n6544), .A(n6528), .B(n6540), .ZN(U3181)
         );
  NAND2_X1 U7484 ( .A1(STATE_REG_0__SCAN_IN), .A2(REQUESTPENDING_REG_SCAN_IN), 
        .ZN(n6534) );
  INV_X1 U7485 ( .A(n6534), .ZN(n6531) );
  NAND2_X1 U7486 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6537) );
  OAI21_X1 U7487 ( .B1(n6531), .B2(n6530), .A(n6537), .ZN(n6532) );
  OAI211_X1 U7488 ( .C1(n6612), .C2(n6535), .A(n6533), .B(n6532), .ZN(U3182)
         );
  NOR3_X1 U7489 ( .A1(NA_N), .A2(n6612), .A3(n6534), .ZN(n6541) );
  NOR2_X1 U7490 ( .A1(NA_N), .A2(n6612), .ZN(n6536) );
  OAI21_X1 U7491 ( .B1(n6536), .B2(n6535), .A(HOLD), .ZN(n6538) );
  OAI211_X1 U7492 ( .C1(REQUESTPENDING_REG_SCAN_IN), .C2(n6538), .A(
        STATE_REG_0__SCAN_IN), .B(n6537), .ZN(n6539) );
  AOI22_X1 U7493 ( .A1(STATE_REG_1__SCAN_IN), .A2(n6541), .B1(n6540), .B2(
        n6539), .ZN(n6542) );
  OAI21_X1 U7494 ( .B1(n6544), .B2(n6543), .A(n6542), .ZN(U3183) );
  INV_X1 U7495 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6547) );
  NAND2_X1 U7496 ( .A1(n6621), .A2(n6545), .ZN(n6587) );
  AOI22_X1 U7497 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6585), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6609), .ZN(n6546) );
  OAI21_X1 U7498 ( .B1(n6547), .B2(n6587), .A(n6546), .ZN(U3184) );
  AOI22_X1 U7499 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6585), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6609), .ZN(n6548) );
  OAI21_X1 U7500 ( .B1(n5119), .B2(n6587), .A(n6548), .ZN(U3185) );
  AOI22_X1 U7501 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6585), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6609), .ZN(n6549) );
  OAI21_X1 U7502 ( .B1(n6550), .B2(n6587), .A(n6549), .ZN(U3186) );
  AOI22_X1 U7503 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6585), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6609), .ZN(n6551) );
  OAI21_X1 U7504 ( .B1(n6552), .B2(n6587), .A(n6551), .ZN(U3187) );
  AOI22_X1 U7505 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6585), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6609), .ZN(n6553) );
  OAI21_X1 U7506 ( .B1(n6554), .B2(n6587), .A(n6553), .ZN(U3188) );
  AOI22_X1 U7507 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6585), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6609), .ZN(n6555) );
  OAI21_X1 U7508 ( .B1(n6557), .B2(n6587), .A(n6555), .ZN(U3189) );
  INV_X1 U7509 ( .A(n6585), .ZN(n6590) );
  INV_X1 U7510 ( .A(n6587), .ZN(n6588) );
  AOI22_X1 U7511 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6588), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6609), .ZN(n6556) );
  OAI21_X1 U7512 ( .B1(n6557), .B2(n6590), .A(n6556), .ZN(U3190) );
  AOI22_X1 U7513 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6585), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6609), .ZN(n6558) );
  OAI21_X1 U7514 ( .B1(n6969), .B2(n6587), .A(n6558), .ZN(U3191) );
  AOI22_X1 U7515 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6585), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6609), .ZN(n6559) );
  OAI21_X1 U7516 ( .B1(n4645), .B2(n6587), .A(n6559), .ZN(U3192) );
  AOI22_X1 U7517 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6585), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6609), .ZN(n6560) );
  OAI21_X1 U7518 ( .B1(n6906), .B2(n6587), .A(n6560), .ZN(U3193) );
  AOI22_X1 U7519 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6588), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6609), .ZN(n6561) );
  OAI21_X1 U7520 ( .B1(n6906), .B2(n6590), .A(n6561), .ZN(U3194) );
  INV_X1 U7521 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6890) );
  OAI222_X1 U7522 ( .A1(n6590), .A2(n6562), .B1(n6890), .B2(n6621), .C1(n6563), 
        .C2(n6587), .ZN(U3195) );
  INV_X1 U7523 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6823) );
  OAI222_X1 U7524 ( .A1(n6590), .A2(n6563), .B1(n6823), .B2(n6621), .C1(n4694), 
        .C2(n6587), .ZN(U3196) );
  AOI22_X1 U7525 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6588), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6609), .ZN(n6564) );
  OAI21_X1 U7526 ( .B1(n4694), .B2(n6590), .A(n6564), .ZN(U3197) );
  AOI22_X1 U7527 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6588), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6609), .ZN(n6565) );
  OAI21_X1 U7528 ( .B1(n6566), .B2(n6590), .A(n6565), .ZN(U3198) );
  AOI22_X1 U7529 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6588), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6609), .ZN(n6567) );
  OAI21_X1 U7530 ( .B1(n6568), .B2(n6590), .A(n6567), .ZN(U3199) );
  AOI22_X1 U7531 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6588), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6609), .ZN(n6569) );
  OAI21_X1 U7532 ( .B1(n6570), .B2(n6590), .A(n6569), .ZN(U3200) );
  INV_X1 U7533 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6996) );
  OAI222_X1 U7534 ( .A1(n6590), .A2(n6572), .B1(n6996), .B2(n6621), .C1(n6571), 
        .C2(n6587), .ZN(U3201) );
  AOI22_X1 U7535 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6585), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6609), .ZN(n6573) );
  OAI21_X1 U7536 ( .B1(n6575), .B2(n6587), .A(n6573), .ZN(U3202) );
  AOI22_X1 U7537 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6588), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6609), .ZN(n6574) );
  OAI21_X1 U7538 ( .B1(n6575), .B2(n6590), .A(n6574), .ZN(U3203) );
  INV_X1 U7539 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6999) );
  OAI222_X1 U7540 ( .A1(n6590), .A2(n6576), .B1(n6999), .B2(n6621), .C1(n4761), 
        .C2(n6587), .ZN(U3204) );
  INV_X1 U7541 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6856) );
  OAI222_X1 U7542 ( .A1(n6590), .A2(n4761), .B1(n6856), .B2(n6621), .C1(n4749), 
        .C2(n6587), .ZN(U3205) );
  INV_X1 U7543 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n6793) );
  OAI222_X1 U7544 ( .A1(n6590), .A2(n4749), .B1(n6793), .B2(n6621), .C1(n6578), 
        .C2(n6587), .ZN(U3206) );
  AOI22_X1 U7545 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6588), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6609), .ZN(n6577) );
  OAI21_X1 U7546 ( .B1(n6578), .B2(n6590), .A(n6577), .ZN(U3207) );
  AOI22_X1 U7547 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6588), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6609), .ZN(n6579) );
  OAI21_X1 U7548 ( .B1(n5268), .B2(n6590), .A(n6579), .ZN(U3208) );
  AOI22_X1 U7549 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6585), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6609), .ZN(n6580) );
  OAI21_X1 U7550 ( .B1(n6582), .B2(n6587), .A(n6580), .ZN(U3209) );
  AOI22_X1 U7551 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6588), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6609), .ZN(n6581) );
  OAI21_X1 U7552 ( .B1(n6582), .B2(n6590), .A(n6581), .ZN(U3210) );
  INV_X1 U7553 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6884) );
  OAI222_X1 U7554 ( .A1(n6590), .A2(n6584), .B1(n6884), .B2(n6621), .C1(n6583), 
        .C2(n6587), .ZN(U3211) );
  AOI22_X1 U7555 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6585), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6609), .ZN(n6586) );
  OAI21_X1 U7556 ( .B1(n3836), .B2(n6587), .A(n6586), .ZN(U3212) );
  AOI22_X1 U7557 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6588), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6609), .ZN(n6589) );
  OAI21_X1 U7558 ( .B1(n3836), .B2(n6590), .A(n6589), .ZN(U3213) );
  MUX2_X1 U7559 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6621), .Z(U3445) );
  MUX2_X1 U7560 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6621), .Z(U3446) );
  MUX2_X1 U7561 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6621), .Z(U3447) );
  MUX2_X1 U7562 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6621), .Z(U3448) );
  INV_X1 U7563 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6593) );
  INV_X1 U7564 ( .A(n6594), .ZN(n6591) );
  AOI21_X1 U7565 ( .B1(n6593), .B2(n6592), .A(n6591), .ZN(U3451) );
  OAI21_X1 U7566 ( .B1(n6596), .B2(n6595), .A(n6594), .ZN(U3452) );
  INV_X1 U7567 ( .A(n6597), .ZN(n6599) );
  OAI221_X1 U7568 ( .B1(n6600), .B2(STATE2_REG_0__SCAN_IN), .C1(n6600), .C2(
        n6599), .A(n6598), .ZN(U3453) );
  AOI21_X1 U7569 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6602) );
  AOI22_X1 U7570 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6602), .B2(n6601), .ZN(n6603) );
  INV_X1 U7571 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6923) );
  AOI22_X1 U7572 ( .A1(n6604), .A2(n6603), .B1(n6923), .B2(n6607), .ZN(U3468)
         );
  INV_X1 U7573 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6973) );
  NOR2_X1 U7574 ( .A1(n6607), .A2(REIP_REG_1__SCAN_IN), .ZN(n6605) );
  AOI22_X1 U7575 ( .A1(n6973), .A2(n6607), .B1(n6606), .B2(n6605), .ZN(U3469)
         );
  NAND2_X1 U7576 ( .A1(n6609), .A2(W_R_N_REG_SCAN_IN), .ZN(n6608) );
  OAI21_X1 U7577 ( .B1(n6609), .B2(READREQUEST_REG_SCAN_IN), .A(n6608), .ZN(
        U3470) );
  AOI211_X1 U7578 ( .C1(n6613), .C2(n6612), .A(n6611), .B(n6610), .ZN(n6620)
         );
  OAI211_X1 U7579 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6615), .A(n6614), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6617) );
  AOI21_X1 U7580 ( .B1(n6617), .B2(STATE2_REG_0__SCAN_IN), .A(n6616), .ZN(
        n6619) );
  NAND2_X1 U7581 ( .A1(n6620), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6618) );
  OAI21_X1 U7582 ( .B1(n6620), .B2(n6619), .A(n6618), .ZN(U3472) );
  MUX2_X1 U7583 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6621), .Z(U3473) );
  AOI22_X1 U7584 ( .A1(n6625), .A2(n6624), .B1(n6623), .B2(n6622), .ZN(n6630)
         );
  AOI22_X1 U7585 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n6628), .B1(n6627), 
        .B2(n6626), .ZN(n6629) );
  OAI211_X1 U7586 ( .C1(n6632), .C2(n6631), .A(n6630), .B(n6629), .ZN(n7018)
         );
  OAI22_X1 U7587 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(keyinput57), .B1(
        keyinput36), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6633) );
  AOI221_X1 U7588 ( .B1(INSTQUEUE_REG_12__6__SCAN_IN), .B2(keyinput57), .C1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .C2(keyinput36), .A(n6633), .ZN(n6640) );
  OAI22_X1 U7589 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(keyinput111), .B1(
        keyinput11), .B2(ADDRESS_REG_12__SCAN_IN), .ZN(n6634) );
  AOI221_X1 U7590 ( .B1(INSTQUEUE_REG_3__5__SCAN_IN), .B2(keyinput111), .C1(
        ADDRESS_REG_12__SCAN_IN), .C2(keyinput11), .A(n6634), .ZN(n6639) );
  OAI22_X1 U7591 ( .A1(DATAI_29_), .A2(keyinput120), .B1(keyinput70), .B2(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n6635) );
  AOI221_X1 U7592 ( .B1(DATAI_29_), .B2(keyinput120), .C1(
        DATAWIDTH_REG_16__SCAN_IN), .C2(keyinput70), .A(n6635), .ZN(n6638) );
  OAI22_X1 U7593 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(keyinput52), .B1(
        INSTQUEUE_REG_1__5__SCAN_IN), .B2(keyinput19), .ZN(n6636) );
  AOI221_X1 U7594 ( .B1(INSTQUEUE_REG_10__4__SCAN_IN), .B2(keyinput52), .C1(
        keyinput19), .C2(INSTQUEUE_REG_1__5__SCAN_IN), .A(n6636), .ZN(n6637)
         );
  NAND4_X1 U7595 ( .A1(n6640), .A2(n6639), .A3(n6638), .A4(n6637), .ZN(n6671)
         );
  OAI22_X1 U7596 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(keyinput27), .B1(
        keyinput80), .B2(EAX_REG_27__SCAN_IN), .ZN(n6641) );
  AOI221_X1 U7597 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(keyinput27), .C1(
        EAX_REG_27__SCAN_IN), .C2(keyinput80), .A(n6641), .ZN(n6648) );
  OAI22_X1 U7598 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(keyinput125), .B1(
        keyinput13), .B2(REIP_REG_5__SCAN_IN), .ZN(n6642) );
  AOI221_X1 U7599 ( .B1(INSTQUEUE_REG_4__0__SCAN_IN), .B2(keyinput125), .C1(
        REIP_REG_5__SCAN_IN), .C2(keyinput13), .A(n6642), .ZN(n6647) );
  OAI22_X1 U7600 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(keyinput54), .B1(
        keyinput101), .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n6643) );
  AOI221_X1 U7601 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(keyinput54), 
        .C1(INSTQUEUE_REG_9__7__SCAN_IN), .C2(keyinput101), .A(n6643), .ZN(
        n6646) );
  OAI22_X1 U7602 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput12), .B1(
        keyinput126), .B2(DATAWIDTH_REG_28__SCAN_IN), .ZN(n6644) );
  AOI221_X1 U7603 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput12), .C1(
        DATAWIDTH_REG_28__SCAN_IN), .C2(keyinput126), .A(n6644), .ZN(n6645) );
  NAND4_X1 U7604 ( .A1(n6648), .A2(n6647), .A3(n6646), .A4(n6645), .ZN(n6670)
         );
  INV_X1 U7605 ( .A(DATAI_18_), .ZN(n6650) );
  OAI22_X1 U7606 ( .A1(n6650), .A2(keyinput37), .B1(keyinput86), .B2(
        REIP_REG_3__SCAN_IN), .ZN(n6649) );
  AOI221_X1 U7607 ( .B1(n6650), .B2(keyinput37), .C1(REIP_REG_3__SCAN_IN), 
        .C2(keyinput86), .A(n6649), .ZN(n6659) );
  OAI22_X1 U7608 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(keyinput31), .B1(
        keyinput67), .B2(DATAWIDTH_REG_18__SCAN_IN), .ZN(n6651) );
  AOI221_X1 U7609 ( .B1(INSTQUEUE_REG_13__5__SCAN_IN), .B2(keyinput31), .C1(
        DATAWIDTH_REG_18__SCAN_IN), .C2(keyinput67), .A(n6651), .ZN(n6658) );
  OAI22_X1 U7610 ( .A1(n6867), .A2(keyinput23), .B1(n6653), .B2(keyinput50), 
        .ZN(n6652) );
  AOI221_X1 U7611 ( .B1(n6867), .B2(keyinput23), .C1(keyinput50), .C2(n6653), 
        .A(n6652), .ZN(n6657) );
  INV_X1 U7612 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n6655) );
  OAI22_X1 U7613 ( .A1(n6655), .A2(keyinput62), .B1(n6809), .B2(keyinput45), 
        .ZN(n6654) );
  AOI221_X1 U7614 ( .B1(n6655), .B2(keyinput62), .C1(keyinput45), .C2(n6809), 
        .A(n6654), .ZN(n6656) );
  NAND4_X1 U7615 ( .A1(n6659), .A2(n6658), .A3(n6657), .A4(n6656), .ZN(n6669)
         );
  OAI22_X1 U7616 ( .A1(EBX_REG_29__SCAN_IN), .A2(keyinput4), .B1(
        EBX_REG_4__SCAN_IN), .B2(keyinput44), .ZN(n6660) );
  AOI221_X1 U7617 ( .B1(EBX_REG_29__SCAN_IN), .B2(keyinput4), .C1(keyinput44), 
        .C2(EBX_REG_4__SCAN_IN), .A(n6660), .ZN(n6667) );
  OAI22_X1 U7618 ( .A1(EBX_REG_18__SCAN_IN), .A2(keyinput15), .B1(HOLD), .B2(
        keyinput35), .ZN(n6661) );
  AOI221_X1 U7619 ( .B1(EBX_REG_18__SCAN_IN), .B2(keyinput15), .C1(keyinput35), 
        .C2(HOLD), .A(n6661), .ZN(n6666) );
  OAI22_X1 U7620 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(keyinput64), .B1(
        REIP_REG_26__SCAN_IN), .B2(keyinput41), .ZN(n6662) );
  AOI221_X1 U7621 ( .B1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(keyinput64), 
        .C1(keyinput41), .C2(REIP_REG_26__SCAN_IN), .A(n6662), .ZN(n6665) );
  OAI22_X1 U7622 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(keyinput84), .B1(
        EBX_REG_22__SCAN_IN), .B2(keyinput28), .ZN(n6663) );
  AOI221_X1 U7623 ( .B1(INSTQUEUE_REG_6__5__SCAN_IN), .B2(keyinput84), .C1(
        keyinput28), .C2(EBX_REG_22__SCAN_IN), .A(n6663), .ZN(n6664) );
  NAND4_X1 U7624 ( .A1(n6667), .A2(n6666), .A3(n6665), .A4(n6664), .ZN(n6668)
         );
  NOR4_X1 U7625 ( .A1(n6671), .A2(n6670), .A3(n6669), .A4(n6668), .ZN(n7016)
         );
  OAI22_X1 U7626 ( .A1(INSTQUEUE_REG_4__6__SCAN_IN), .A2(keyinput79), .B1(
        keyinput77), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6672) );
  AOI221_X1 U7627 ( .B1(INSTQUEUE_REG_4__6__SCAN_IN), .B2(keyinput79), .C1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .C2(keyinput77), .A(n6672), .ZN(n6679) );
  OAI22_X1 U7628 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(keyinput103), .B1(
        STATE2_REG_3__SCAN_IN), .B2(keyinput82), .ZN(n6673) );
  AOI221_X1 U7629 ( .B1(INSTQUEUE_REG_5__4__SCAN_IN), .B2(keyinput103), .C1(
        keyinput82), .C2(STATE2_REG_3__SCAN_IN), .A(n6673), .ZN(n6678) );
  OAI22_X1 U7630 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(keyinput40), .B1(
        keyinput78), .B2(ADDRESS_REG_22__SCAN_IN), .ZN(n6674) );
  AOI221_X1 U7631 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(keyinput40), 
        .C1(ADDRESS_REG_22__SCAN_IN), .C2(keyinput78), .A(n6674), .ZN(n6677)
         );
  OAI22_X1 U7632 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(keyinput75), .B1(
        DATAWIDTH_REG_3__SCAN_IN), .B2(keyinput47), .ZN(n6675) );
  AOI221_X1 U7633 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput75), 
        .C1(keyinput47), .C2(DATAWIDTH_REG_3__SCAN_IN), .A(n6675), .ZN(n6676)
         );
  NAND4_X1 U7634 ( .A1(n6679), .A2(n6678), .A3(n6677), .A4(n6676), .ZN(n6707)
         );
  OAI22_X1 U7635 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(keyinput89), .B1(
        keyinput10), .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6680) );
  AOI221_X1 U7636 ( .B1(INSTQUEUE_REG_2__1__SCAN_IN), .B2(keyinput89), .C1(
        INSTQUEUE_REG_12__5__SCAN_IN), .C2(keyinput10), .A(n6680), .ZN(n6687)
         );
  OAI22_X1 U7637 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(keyinput24), .B1(
        keyinput3), .B2(DATAI_31_), .ZN(n6681) );
  AOI221_X1 U7638 ( .B1(INSTQUEUE_REG_14__4__SCAN_IN), .B2(keyinput24), .C1(
        DATAI_31_), .C2(keyinput3), .A(n6681), .ZN(n6686) );
  OAI22_X1 U7639 ( .A1(UWORD_REG_13__SCAN_IN), .A2(keyinput55), .B1(
        keyinput116), .B2(DATAO_REG_13__SCAN_IN), .ZN(n6682) );
  AOI221_X1 U7640 ( .B1(UWORD_REG_13__SCAN_IN), .B2(keyinput55), .C1(
        DATAO_REG_13__SCAN_IN), .C2(keyinput116), .A(n6682), .ZN(n6685) );
  OAI22_X1 U7641 ( .A1(DATAI_30_), .A2(keyinput68), .B1(keyinput72), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n6683) );
  AOI221_X1 U7642 ( .B1(DATAI_30_), .B2(keyinput68), .C1(UWORD_REG_12__SCAN_IN), .C2(keyinput72), .A(n6683), .ZN(n6684) );
  NAND4_X1 U7643 ( .A1(n6687), .A2(n6686), .A3(n6685), .A4(n6684), .ZN(n6706)
         );
  OAI22_X1 U7644 ( .A1(STATE2_REG_2__SCAN_IN), .A2(keyinput91), .B1(keyinput1), 
        .B2(REIP_REG_25__SCAN_IN), .ZN(n6688) );
  AOI221_X1 U7645 ( .B1(STATE2_REG_2__SCAN_IN), .B2(keyinput91), .C1(
        REIP_REG_25__SCAN_IN), .C2(keyinput1), .A(n6688), .ZN(n6695) );
  OAI22_X1 U7646 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(keyinput48), .B1(
        DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput108), .ZN(n6689) );
  AOI221_X1 U7647 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(keyinput48), 
        .C1(keyinput108), .C2(DATAWIDTH_REG_8__SCAN_IN), .A(n6689), .ZN(n6694)
         );
  OAI22_X1 U7648 ( .A1(EAX_REG_25__SCAN_IN), .A2(keyinput110), .B1(keyinput38), 
        .B2(ADDRESS_REG_21__SCAN_IN), .ZN(n6690) );
  AOI221_X1 U7649 ( .B1(EAX_REG_25__SCAN_IN), .B2(keyinput110), .C1(
        ADDRESS_REG_21__SCAN_IN), .C2(keyinput38), .A(n6690), .ZN(n6693) );
  OAI22_X1 U7650 ( .A1(REIP_REG_21__SCAN_IN), .A2(keyinput119), .B1(DATAI_2_), 
        .B2(keyinput74), .ZN(n6691) );
  AOI221_X1 U7651 ( .B1(REIP_REG_21__SCAN_IN), .B2(keyinput119), .C1(
        keyinput74), .C2(DATAI_2_), .A(n6691), .ZN(n6692) );
  NAND4_X1 U7652 ( .A1(n6695), .A2(n6694), .A3(n6693), .A4(n6692), .ZN(n6705)
         );
  OAI22_X1 U7653 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(keyinput18), .B1(
        keyinput30), .B2(EAX_REG_8__SCAN_IN), .ZN(n6696) );
  AOI221_X1 U7654 ( .B1(INSTQUEUE_REG_1__3__SCAN_IN), .B2(keyinput18), .C1(
        EAX_REG_8__SCAN_IN), .C2(keyinput30), .A(n6696), .ZN(n6703) );
  OAI22_X1 U7655 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(keyinput51), .B1(
        DATAWIDTH_REG_1__SCAN_IN), .B2(keyinput46), .ZN(n6697) );
  AOI221_X1 U7656 ( .B1(INSTQUEUE_REG_3__0__SCAN_IN), .B2(keyinput51), .C1(
        keyinput46), .C2(DATAWIDTH_REG_1__SCAN_IN), .A(n6697), .ZN(n6702) );
  OAI22_X1 U7657 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(keyinput90), .B1(
        keyinput8), .B2(REIP_REG_14__SCAN_IN), .ZN(n6698) );
  AOI221_X1 U7658 ( .B1(INSTQUEUE_REG_2__0__SCAN_IN), .B2(keyinput90), .C1(
        REIP_REG_14__SCAN_IN), .C2(keyinput8), .A(n6698), .ZN(n6701) );
  OAI22_X1 U7659 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(keyinput117), .B1(
        DATAI_14_), .B2(keyinput71), .ZN(n6699) );
  AOI221_X1 U7660 ( .B1(INSTQUEUE_REG_7__4__SCAN_IN), .B2(keyinput117), .C1(
        keyinput71), .C2(DATAI_14_), .A(n6699), .ZN(n6700) );
  NAND4_X1 U7661 ( .A1(n6703), .A2(n6702), .A3(n6701), .A4(n6700), .ZN(n6704)
         );
  NOR4_X1 U7662 ( .A1(n6707), .A2(n6706), .A3(n6705), .A4(n6704), .ZN(n7015)
         );
  AOI22_X1 U7663 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(keyinput155), .B1(
        INSTQUEUE_REG_7__1__SCAN_IN), .B2(keyinput190), .ZN(n6708) );
  OAI221_X1 U7664 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(keyinput155), .C1(
        INSTQUEUE_REG_7__1__SCAN_IN), .C2(keyinput190), .A(n6708), .ZN(n6715)
         );
  AOI22_X1 U7665 ( .A1(DATAI_31_), .A2(keyinput131), .B1(
        INSTQUEUE_REG_2__7__SCAN_IN), .B2(keyinput177), .ZN(n6709) );
  OAI221_X1 U7666 ( .B1(DATAI_31_), .B2(keyinput131), .C1(
        INSTQUEUE_REG_2__7__SCAN_IN), .C2(keyinput177), .A(n6709), .ZN(n6714)
         );
  AOI22_X1 U7667 ( .A1(DATAI_22_), .A2(keyinput235), .B1(EAX_REG_3__SCAN_IN), 
        .B2(keyinput157), .ZN(n6710) );
  OAI221_X1 U7668 ( .B1(DATAI_22_), .B2(keyinput235), .C1(EAX_REG_3__SCAN_IN), 
        .C2(keyinput157), .A(n6710), .ZN(n6713) );
  AOI22_X1 U7669 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(keyinput198), .B1(
        INSTADDRPOINTER_REG_8__SCAN_IN), .B2(keyinput181), .ZN(n6711) );
  OAI221_X1 U7670 ( .B1(DATAWIDTH_REG_16__SCAN_IN), .B2(keyinput198), .C1(
        INSTADDRPOINTER_REG_8__SCAN_IN), .C2(keyinput181), .A(n6711), .ZN(
        n6712) );
  NOR4_X1 U7671 ( .A1(n6715), .A2(n6714), .A3(n6713), .A4(n6712), .ZN(n6743)
         );
  AOI22_X1 U7672 ( .A1(DATAI_14_), .A2(keyinput199), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput145), .ZN(n6716) );
  OAI221_X1 U7673 ( .B1(DATAI_14_), .B2(keyinput199), .C1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .C2(keyinput145), .A(n6716), .ZN(
        n6723) );
  AOI22_X1 U7674 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(keyinput144), .B1(
        INSTQUEUE_REG_9__7__SCAN_IN), .B2(keyinput229), .ZN(n6717) );
  OAI221_X1 U7675 ( .B1(INSTQUEUE_REG_1__7__SCAN_IN), .B2(keyinput144), .C1(
        INSTQUEUE_REG_9__7__SCAN_IN), .C2(keyinput229), .A(n6717), .ZN(n6722)
         );
  AOI22_X1 U7676 ( .A1(EBX_REG_17__SCAN_IN), .A2(keyinput171), .B1(
        INSTQUEUE_REG_13__4__SCAN_IN), .B2(keyinput243), .ZN(n6718) );
  OAI221_X1 U7677 ( .B1(EBX_REG_17__SCAN_IN), .B2(keyinput171), .C1(
        INSTQUEUE_REG_13__4__SCAN_IN), .C2(keyinput243), .A(n6718), .ZN(n6721)
         );
  AOI22_X1 U7678 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(keyinput245), .B1(
        INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(keyinput168), .ZN(n6719) );
  OAI221_X1 U7679 ( .B1(INSTQUEUE_REG_7__4__SCAN_IN), .B2(keyinput245), .C1(
        INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(keyinput168), .A(n6719), .ZN(
        n6720) );
  NOR4_X1 U7680 ( .A1(n6723), .A2(n6722), .A3(n6721), .A4(n6720), .ZN(n6742)
         );
  AOI22_X1 U7681 ( .A1(HOLD), .A2(keyinput163), .B1(REIP_REG_11__SCAN_IN), 
        .B2(keyinput227), .ZN(n6724) );
  OAI221_X1 U7682 ( .B1(HOLD), .B2(keyinput163), .C1(REIP_REG_11__SCAN_IN), 
        .C2(keyinput227), .A(n6724), .ZN(n6731) );
  AOI22_X1 U7683 ( .A1(DATAWIDTH_REG_1__SCAN_IN), .A2(keyinput174), .B1(
        INSTQUEUE_REG_6__5__SCAN_IN), .B2(keyinput212), .ZN(n6725) );
  OAI221_X1 U7684 ( .B1(DATAWIDTH_REG_1__SCAN_IN), .B2(keyinput174), .C1(
        INSTQUEUE_REG_6__5__SCAN_IN), .C2(keyinput212), .A(n6725), .ZN(n6730)
         );
  AOI22_X1 U7685 ( .A1(ADDRESS_REG_20__SCAN_IN), .A2(keyinput249), .B1(
        EAX_REG_4__SCAN_IN), .B2(keyinput142), .ZN(n6726) );
  OAI221_X1 U7686 ( .B1(ADDRESS_REG_20__SCAN_IN), .B2(keyinput249), .C1(
        EAX_REG_4__SCAN_IN), .C2(keyinput142), .A(n6726), .ZN(n6729) );
  AOI22_X1 U7687 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput140), .B1(
        INSTQUEUE_REG_0__6__SCAN_IN), .B2(keyinput234), .ZN(n6727) );
  OAI221_X1 U7688 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput140), .C1(
        INSTQUEUE_REG_0__6__SCAN_IN), .C2(keyinput234), .A(n6727), .ZN(n6728)
         );
  NOR4_X1 U7689 ( .A1(n6731), .A2(n6730), .A3(n6729), .A4(n6728), .ZN(n6741)
         );
  AOI22_X1 U7690 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(keyinput236), .B1(
        INSTADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput203), .ZN(n6732) );
  OAI221_X1 U7691 ( .B1(DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput236), .C1(
        INSTADDRPOINTER_REG_28__SCAN_IN), .C2(keyinput203), .A(n6732), .ZN(
        n6739) );
  AOI22_X1 U7692 ( .A1(DATAI_18_), .A2(keyinput165), .B1(EBX_REG_5__SCAN_IN), 
        .B2(keyinput178), .ZN(n6733) );
  OAI221_X1 U7693 ( .B1(DATAI_18_), .B2(keyinput165), .C1(EBX_REG_5__SCAN_IN), 
        .C2(keyinput178), .A(n6733), .ZN(n6738) );
  AOI22_X1 U7694 ( .A1(REIP_REG_5__SCAN_IN), .A2(keyinput141), .B1(
        INSTQUEUE_REG_4__0__SCAN_IN), .B2(keyinput253), .ZN(n6734) );
  OAI221_X1 U7695 ( .B1(REIP_REG_5__SCAN_IN), .B2(keyinput141), .C1(
        INSTQUEUE_REG_4__0__SCAN_IN), .C2(keyinput253), .A(n6734), .ZN(n6737)
         );
  AOI22_X1 U7696 ( .A1(DATAO_REG_21__SCAN_IN), .A2(keyinput148), .B1(
        INSTQUEUE_REG_1__3__SCAN_IN), .B2(keyinput146), .ZN(n6735) );
  OAI221_X1 U7697 ( .B1(DATAO_REG_21__SCAN_IN), .B2(keyinput148), .C1(
        INSTQUEUE_REG_1__3__SCAN_IN), .C2(keyinput146), .A(n6735), .ZN(n6736)
         );
  NOR4_X1 U7698 ( .A1(n6739), .A2(n6738), .A3(n6737), .A4(n6736), .ZN(n6740)
         );
  NAND4_X1 U7699 ( .A1(n6743), .A2(n6742), .A3(n6741), .A4(n6740), .ZN(n6882)
         );
  AOI22_X1 U7700 ( .A1(REIP_REG_9__SCAN_IN), .A2(keyinput228), .B1(
        REIP_REG_21__SCAN_IN), .B2(keyinput247), .ZN(n6744) );
  OAI221_X1 U7701 ( .B1(REIP_REG_9__SCAN_IN), .B2(keyinput228), .C1(
        REIP_REG_21__SCAN_IN), .C2(keyinput247), .A(n6744), .ZN(n6751) );
  AOI22_X1 U7702 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput134), .B1(
        STATE2_REG_3__SCAN_IN), .B2(keyinput210), .ZN(n6745) );
  OAI221_X1 U7703 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput134), .C1(
        STATE2_REG_3__SCAN_IN), .C2(keyinput210), .A(n6745), .ZN(n6750) );
  AOI22_X1 U7704 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(keyinput215), .B1(
        INSTQUEUE_REG_14__4__SCAN_IN), .B2(keyinput152), .ZN(n6746) );
  OAI221_X1 U7705 ( .B1(INSTQUEUE_REG_13__0__SCAN_IN), .B2(keyinput215), .C1(
        INSTQUEUE_REG_14__4__SCAN_IN), .C2(keyinput152), .A(n6746), .ZN(n6749)
         );
  AOI22_X1 U7706 ( .A1(EAX_REG_25__SCAN_IN), .A2(keyinput238), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(keyinput205), .ZN(n6747) );
  OAI221_X1 U7707 ( .B1(EAX_REG_25__SCAN_IN), .B2(keyinput238), .C1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .C2(keyinput205), .A(n6747), .ZN(
        n6748) );
  NOR4_X1 U7708 ( .A1(n6751), .A2(n6750), .A3(n6749), .A4(n6748), .ZN(n6779)
         );
  AOI22_X1 U7709 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(keyinput180), .B1(
        INSTQUEUE_REG_0__4__SCAN_IN), .B2(keyinput250), .ZN(n6752) );
  OAI221_X1 U7710 ( .B1(INSTQUEUE_REG_10__4__SCAN_IN), .B2(keyinput180), .C1(
        INSTQUEUE_REG_0__4__SCAN_IN), .C2(keyinput250), .A(n6752), .ZN(n6759)
         );
  AOI22_X1 U7711 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(keyinput175), .B1(
        EBX_REG_26__SCAN_IN), .B2(keyinput225), .ZN(n6753) );
  OAI221_X1 U7712 ( .B1(DATAWIDTH_REG_3__SCAN_IN), .B2(keyinput175), .C1(
        EBX_REG_26__SCAN_IN), .C2(keyinput225), .A(n6753), .ZN(n6758) );
  AOI22_X1 U7713 ( .A1(DATAO_REG_9__SCAN_IN), .A2(keyinput232), .B1(
        INSTADDRPOINTER_REG_24__SCAN_IN), .B2(keyinput246), .ZN(n6754) );
  OAI221_X1 U7714 ( .B1(DATAO_REG_9__SCAN_IN), .B2(keyinput232), .C1(
        INSTADDRPOINTER_REG_24__SCAN_IN), .C2(keyinput246), .A(n6754), .ZN(
        n6757) );
  AOI22_X1 U7715 ( .A1(REIP_REG_25__SCAN_IN), .A2(keyinput129), .B1(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(keyinput182), .ZN(n6755) );
  OAI221_X1 U7716 ( .B1(REIP_REG_25__SCAN_IN), .B2(keyinput129), .C1(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(keyinput182), .A(n6755), .ZN(
        n6756) );
  NOR4_X1 U7717 ( .A1(n6759), .A2(n6758), .A3(n6757), .A4(n6756), .ZN(n6778)
         );
  AOI22_X1 U7718 ( .A1(DATAI_2_), .A2(keyinput202), .B1(EBX_REG_31__SCAN_IN), 
        .B2(keyinput189), .ZN(n6760) );
  OAI221_X1 U7719 ( .B1(DATAI_2_), .B2(keyinput202), .C1(EBX_REG_31__SCAN_IN), 
        .C2(keyinput189), .A(n6760), .ZN(n6767) );
  AOI22_X1 U7720 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(keyinput185), .B1(
        INSTQUEUE_REG_6__0__SCAN_IN), .B2(keyinput170), .ZN(n6761) );
  OAI221_X1 U7721 ( .B1(INSTQUEUE_REG_12__6__SCAN_IN), .B2(keyinput185), .C1(
        INSTQUEUE_REG_6__0__SCAN_IN), .C2(keyinput170), .A(n6761), .ZN(n6766)
         );
  AOI22_X1 U7722 ( .A1(DATAO_REG_24__SCAN_IN), .A2(keyinput241), .B1(
        REIP_REG_14__SCAN_IN), .B2(keyinput136), .ZN(n6762) );
  OAI221_X1 U7723 ( .B1(DATAO_REG_24__SCAN_IN), .B2(keyinput241), .C1(
        REIP_REG_14__SCAN_IN), .C2(keyinput136), .A(n6762), .ZN(n6765) );
  AOI22_X1 U7724 ( .A1(ADDRESS_REG_11__SCAN_IN), .A2(keyinput213), .B1(
        DATAI_29_), .B2(keyinput248), .ZN(n6763) );
  OAI221_X1 U7725 ( .B1(ADDRESS_REG_11__SCAN_IN), .B2(keyinput213), .C1(
        DATAI_29_), .C2(keyinput248), .A(n6763), .ZN(n6764) );
  NOR4_X1 U7726 ( .A1(n6767), .A2(n6766), .A3(n6765), .A4(n6764), .ZN(n6777)
         );
  AOI22_X1 U7727 ( .A1(DATAO_REG_18__SCAN_IN), .A2(keyinput222), .B1(
        REIP_REG_26__SCAN_IN), .B2(keyinput169), .ZN(n6768) );
  OAI221_X1 U7728 ( .B1(DATAO_REG_18__SCAN_IN), .B2(keyinput222), .C1(
        REIP_REG_26__SCAN_IN), .C2(keyinput169), .A(n6768), .ZN(n6775) );
  AOI22_X1 U7729 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(keyinput187), .B1(
        EAX_REG_8__SCAN_IN), .B2(keyinput158), .ZN(n6769) );
  OAI221_X1 U7730 ( .B1(DATAWIDTH_REG_10__SCAN_IN), .B2(keyinput187), .C1(
        EAX_REG_8__SCAN_IN), .C2(keyinput158), .A(n6769), .ZN(n6774) );
  AOI22_X1 U7731 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(keyinput184), .B1(
        EAX_REG_27__SCAN_IN), .B2(keyinput208), .ZN(n6770) );
  OAI221_X1 U7732 ( .B1(DATAWIDTH_REG_27__SCAN_IN), .B2(keyinput184), .C1(
        EAX_REG_27__SCAN_IN), .C2(keyinput208), .A(n6770), .ZN(n6773) );
  AOI22_X1 U7733 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(keyinput193), .B1(
        EAX_REG_2__SCAN_IN), .B2(keyinput130), .ZN(n6771) );
  OAI221_X1 U7734 ( .B1(PHYADDRPOINTER_REG_0__SCAN_IN), .B2(keyinput193), .C1(
        EAX_REG_2__SCAN_IN), .C2(keyinput130), .A(n6771), .ZN(n6772) );
  NOR4_X1 U7735 ( .A1(n6775), .A2(n6774), .A3(n6773), .A4(n6772), .ZN(n6776)
         );
  NAND4_X1 U7736 ( .A1(n6779), .A2(n6778), .A3(n6777), .A4(n6776), .ZN(n6881)
         );
  AOI22_X1 U7737 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(keyinput162), .B1(
        n5119), .B2(keyinput214), .ZN(n6780) );
  OAI221_X1 U7738 ( .B1(INSTQUEUE_REG_14__0__SCAN_IN), .B2(keyinput162), .C1(
        n5119), .C2(keyinput214), .A(n6780), .ZN(n6791) );
  INV_X1 U7739 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6982) );
  AOI22_X1 U7740 ( .A1(n6982), .A2(keyinput216), .B1(keyinput176), .B2(n6782), 
        .ZN(n6781) );
  OAI221_X1 U7741 ( .B1(n6982), .B2(keyinput216), .C1(n6782), .C2(keyinput176), 
        .A(n6781), .ZN(n6790) );
  AOI22_X1 U7742 ( .A1(n6785), .A2(keyinput183), .B1(n6784), .B2(keyinput196), 
        .ZN(n6783) );
  OAI221_X1 U7743 ( .B1(n6785), .B2(keyinput183), .C1(n6784), .C2(keyinput196), 
        .A(n6783), .ZN(n6789) );
  INV_X1 U7744 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n6787) );
  AOI22_X1 U7745 ( .A1(n6983), .A2(keyinput137), .B1(n6787), .B2(keyinput159), 
        .ZN(n6786) );
  OAI221_X1 U7746 ( .B1(n6983), .B2(keyinput137), .C1(n6787), .C2(keyinput159), 
        .A(n6786), .ZN(n6788) );
  NOR4_X1 U7747 ( .A1(n6791), .A2(n6790), .A3(n6789), .A4(n6788), .ZN(n6831)
         );
  INV_X1 U7748 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n6794) );
  AOI22_X1 U7749 ( .A1(n6794), .A2(keyinput179), .B1(keyinput206), .B2(n6793), 
        .ZN(n6792) );
  OAI221_X1 U7750 ( .B1(n6794), .B2(keyinput179), .C1(n6793), .C2(keyinput206), 
        .A(n6792), .ZN(n6806) );
  AOI22_X1 U7751 ( .A1(n6936), .A2(keyinput133), .B1(keyinput156), .B2(n6796), 
        .ZN(n6795) );
  OAI221_X1 U7752 ( .B1(n6936), .B2(keyinput133), .C1(n6796), .C2(keyinput156), 
        .A(n6795), .ZN(n6805) );
  INV_X1 U7753 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n6798) );
  AOI22_X1 U7754 ( .A1(n6799), .A2(keyinput219), .B1(n6798), .B2(keyinput239), 
        .ZN(n6797) );
  OAI221_X1 U7755 ( .B1(n6799), .B2(keyinput219), .C1(n6798), .C2(keyinput239), 
        .A(n6797), .ZN(n6804) );
  INV_X1 U7756 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n6800) );
  XOR2_X1 U7757 ( .A(n6800), .B(keyinput200), .Z(n6802) );
  XNOR2_X1 U7758 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(keyinput192), .ZN(
        n6801) );
  NAND2_X1 U7759 ( .A1(n6802), .A2(n6801), .ZN(n6803) );
  NOR4_X1 U7760 ( .A1(n6806), .A2(n6805), .A3(n6804), .A4(n6803), .ZN(n6830)
         );
  AOI22_X1 U7761 ( .A1(n3929), .A2(keyinput233), .B1(keyinput211), .B2(n6996), 
        .ZN(n6807) );
  OAI221_X1 U7762 ( .B1(n3929), .B2(keyinput233), .C1(n6996), .C2(keyinput211), 
        .A(n6807), .ZN(n6816) );
  AOI22_X1 U7763 ( .A1(n6979), .A2(keyinput255), .B1(n6809), .B2(keyinput173), 
        .ZN(n6808) );
  OAI221_X1 U7764 ( .B1(n6979), .B2(keyinput255), .C1(n6809), .C2(keyinput173), 
        .A(n6808), .ZN(n6815) );
  INV_X1 U7765 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n7002) );
  AOI22_X1 U7766 ( .A1(n6940), .A2(keyinput160), .B1(n7002), .B2(keyinput194), 
        .ZN(n6810) );
  OAI221_X1 U7767 ( .B1(n6940), .B2(keyinput160), .C1(n7002), .C2(keyinput194), 
        .A(n6810), .ZN(n6814) );
  AOI22_X1 U7768 ( .A1(n4645), .A2(keyinput204), .B1(n6812), .B2(keyinput143), 
        .ZN(n6811) );
  OAI221_X1 U7769 ( .B1(n4645), .B2(keyinput204), .C1(n6812), .C2(keyinput143), 
        .A(n6811), .ZN(n6813) );
  NOR4_X1 U7770 ( .A1(n6816), .A2(n6815), .A3(n6814), .A4(n6813), .ZN(n6829)
         );
  INV_X1 U7771 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6818) );
  INV_X1 U7772 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n6950) );
  AOI22_X1 U7773 ( .A1(n6818), .A2(keyinput218), .B1(keyinput186), .B2(n6950), 
        .ZN(n6817) );
  OAI221_X1 U7774 ( .B1(n6818), .B2(keyinput218), .C1(n6950), .C2(keyinput186), 
        .A(n6817), .ZN(n6827) );
  INV_X1 U7775 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n7001) );
  AOI22_X1 U7776 ( .A1(n7001), .A2(keyinput230), .B1(keyinput201), .B2(n6933), 
        .ZN(n6819) );
  OAI221_X1 U7777 ( .B1(n7001), .B2(keyinput230), .C1(n6933), .C2(keyinput201), 
        .A(n6819), .ZN(n6826) );
  INV_X1 U7778 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6821) );
  AOI22_X1 U7779 ( .A1(n6934), .A2(keyinput224), .B1(n6821), .B2(keyinput138), 
        .ZN(n6820) );
  OAI221_X1 U7780 ( .B1(n6934), .B2(keyinput224), .C1(n6821), .C2(keyinput138), 
        .A(n6820), .ZN(n6825) );
  AOI22_X1 U7781 ( .A1(n6823), .A2(keyinput139), .B1(n6887), .B2(keyinput226), 
        .ZN(n6822) );
  OAI221_X1 U7782 ( .B1(n6823), .B2(keyinput139), .C1(n6887), .C2(keyinput226), 
        .A(n6822), .ZN(n6824) );
  NOR4_X1 U7783 ( .A1(n6827), .A2(n6826), .A3(n6825), .A4(n6824), .ZN(n6828)
         );
  NAND4_X1 U7784 ( .A1(n6831), .A2(n6830), .A3(n6829), .A4(n6828), .ZN(n6880)
         );
  AOI22_X1 U7785 ( .A1(n6921), .A2(keyinput135), .B1(n6888), .B2(keyinput220), 
        .ZN(n6832) );
  OAI221_X1 U7786 ( .B1(n6921), .B2(keyinput135), .C1(n6888), .C2(keyinput220), 
        .A(n6832), .ZN(n6841) );
  INV_X1 U7787 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n6835) );
  AOI22_X1 U7788 ( .A1(n6835), .A2(keyinput217), .B1(keyinput172), .B2(n6834), 
        .ZN(n6833) );
  OAI221_X1 U7789 ( .B1(n6835), .B2(keyinput217), .C1(n6834), .C2(keyinput172), 
        .A(n6833), .ZN(n6840) );
  INV_X1 U7790 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6951) );
  AOI22_X1 U7791 ( .A1(n3827), .A2(keyinput132), .B1(n6951), .B2(keyinput188), 
        .ZN(n6836) );
  OAI221_X1 U7792 ( .B1(n3827), .B2(keyinput132), .C1(n6951), .C2(keyinput188), 
        .A(n6836), .ZN(n6839) );
  INV_X1 U7793 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n6988) );
  INV_X1 U7794 ( .A(DATAI_9_), .ZN(n6958) );
  AOI22_X1 U7795 ( .A1(n6988), .A2(keyinput153), .B1(n6958), .B2(keyinput167), 
        .ZN(n6837) );
  OAI221_X1 U7796 ( .B1(n6988), .B2(keyinput153), .C1(n6958), .C2(keyinput167), 
        .A(n6837), .ZN(n6838) );
  NOR4_X1 U7797 ( .A1(n6841), .A2(n6840), .A3(n6839), .A4(n6838), .ZN(n6878)
         );
  AOI22_X1 U7798 ( .A1(n6884), .A2(keyinput154), .B1(n6970), .B2(keyinput252), 
        .ZN(n6842) );
  OAI221_X1 U7799 ( .B1(n6884), .B2(keyinput154), .C1(n6970), .C2(keyinput252), 
        .A(n6842), .ZN(n6851) );
  AOI22_X1 U7800 ( .A1(n6930), .A2(keyinput240), .B1(keyinput209), .B2(n6905), 
        .ZN(n6843) );
  OAI221_X1 U7801 ( .B1(n6930), .B2(keyinput240), .C1(n6905), .C2(keyinput209), 
        .A(n6843), .ZN(n6850) );
  AOI22_X1 U7802 ( .A1(n6847), .A2(keyinput244), .B1(keyinput223), .B2(n6919), 
        .ZN(n6846) );
  OAI221_X1 U7803 ( .B1(n6847), .B2(keyinput244), .C1(n6919), .C2(keyinput223), 
        .A(n6846), .ZN(n6848) );
  NOR4_X1 U7804 ( .A1(n6851), .A2(n6850), .A3(n6849), .A4(n6848), .ZN(n6877)
         );
  INV_X1 U7805 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n6853) );
  AOI22_X1 U7806 ( .A1(n6853), .A2(keyinput147), .B1(keyinput221), .B2(n6954), 
        .ZN(n6852) );
  OAI221_X1 U7807 ( .B1(n6853), .B2(keyinput147), .C1(n6954), .C2(keyinput221), 
        .A(n6852), .ZN(n6862) );
  AOI22_X1 U7808 ( .A1(n6856), .A2(keyinput166), .B1(keyinput195), .B2(n6855), 
        .ZN(n6854) );
  OAI221_X1 U7809 ( .B1(n6856), .B2(keyinput166), .C1(n6855), .C2(keyinput195), 
        .A(n6854), .ZN(n6861) );
  INV_X1 U7810 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n6998) );
  AOI22_X1 U7811 ( .A1(n6972), .A2(keyinput150), .B1(keyinput242), .B2(n6998), 
        .ZN(n6857) );
  OAI221_X1 U7812 ( .B1(n6972), .B2(keyinput150), .C1(n6998), .C2(keyinput242), 
        .A(n6857), .ZN(n6860) );
  AOI22_X1 U7813 ( .A1(n6964), .A2(keyinput128), .B1(keyinput237), .B2(n6937), 
        .ZN(n6858) );
  OAI221_X1 U7814 ( .B1(n6964), .B2(keyinput128), .C1(n6937), .C2(keyinput237), 
        .A(n6858), .ZN(n6859) );
  NOR4_X1 U7815 ( .A1(n6862), .A2(n6861), .A3(n6860), .A4(n6859), .ZN(n6876)
         );
  INV_X1 U7816 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n6864) );
  AOI22_X1 U7817 ( .A1(n6903), .A2(keyinput197), .B1(n6864), .B2(keyinput207), 
        .ZN(n6863) );
  OAI221_X1 U7818 ( .B1(n6903), .B2(keyinput197), .C1(n6864), .C2(keyinput207), 
        .A(n6863), .ZN(n6874) );
  INV_X1 U7819 ( .A(EAX_REG_31__SCAN_IN), .ZN(n6900) );
  INV_X1 U7820 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6967) );
  AOI22_X1 U7821 ( .A1(n6900), .A2(keyinput149), .B1(n6967), .B2(keyinput161), 
        .ZN(n6865) );
  OAI221_X1 U7822 ( .B1(n6900), .B2(keyinput149), .C1(n6967), .C2(keyinput161), 
        .A(n6865), .ZN(n6873) );
  AOI22_X1 U7823 ( .A1(n6868), .A2(keyinput254), .B1(n6867), .B2(keyinput151), 
        .ZN(n6866) );
  OAI221_X1 U7824 ( .B1(n6868), .B2(keyinput254), .C1(n6867), .C2(keyinput151), 
        .A(n6866), .ZN(n6872) );
  INV_X1 U7825 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6870) );
  AOI22_X1 U7826 ( .A1(n6973), .A2(keyinput191), .B1(n6870), .B2(keyinput231), 
        .ZN(n6869) );
  OAI221_X1 U7827 ( .B1(n6973), .B2(keyinput191), .C1(n6870), .C2(keyinput231), 
        .A(n6869), .ZN(n6871) );
  NOR4_X1 U7828 ( .A1(n6874), .A2(n6873), .A3(n6872), .A4(n6871), .ZN(n6875)
         );
  NAND4_X1 U7829 ( .A1(n6878), .A2(n6877), .A3(n6876), .A4(n6875), .ZN(n6879)
         );
  NOR4_X1 U7830 ( .A1(n6882), .A2(n6881), .A3(n6880), .A4(n6879), .ZN(n7013)
         );
  INV_X1 U7831 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n6885) );
  AOI22_X1 U7832 ( .A1(n6885), .A2(keyinput16), .B1(keyinput26), .B2(n6884), 
        .ZN(n6883) );
  OAI221_X1 U7833 ( .B1(n6885), .B2(keyinput16), .C1(n6884), .C2(keyinput26), 
        .A(n6883), .ZN(n6897) );
  AOI22_X1 U7834 ( .A1(n6888), .A2(keyinput92), .B1(keyinput98), .B2(n6887), 
        .ZN(n6886) );
  OAI221_X1 U7835 ( .B1(n6888), .B2(keyinput92), .C1(n6887), .C2(keyinput98), 
        .A(n6886), .ZN(n6896) );
  AOI22_X1 U7836 ( .A1(n6891), .A2(keyinput94), .B1(n6890), .B2(keyinput85), 
        .ZN(n6889) );
  OAI221_X1 U7837 ( .B1(n6891), .B2(keyinput94), .C1(n6890), .C2(keyinput85), 
        .A(n6889), .ZN(n6895) );
  AOI22_X1 U7838 ( .A1(n3815), .A2(keyinput97), .B1(keyinput20), .B2(n6893), 
        .ZN(n6892) );
  OAI221_X1 U7839 ( .B1(n3815), .B2(keyinput97), .C1(n6893), .C2(keyinput20), 
        .A(n6892), .ZN(n6894) );
  NOR4_X1 U7840 ( .A1(n6897), .A2(n6896), .A3(n6895), .A4(n6894), .ZN(n6948)
         );
  AOI22_X1 U7841 ( .A1(n6900), .A2(keyinput21), .B1(keyinput113), .B2(n6899), 
        .ZN(n6898) );
  OAI221_X1 U7842 ( .B1(n6900), .B2(keyinput21), .C1(n6899), .C2(keyinput113), 
        .A(n6898), .ZN(n6913) );
  AOI22_X1 U7843 ( .A1(n6903), .A2(keyinput69), .B1(n6902), .B2(keyinput123), 
        .ZN(n6901) );
  OAI221_X1 U7844 ( .B1(n6903), .B2(keyinput69), .C1(n6902), .C2(keyinput123), 
        .A(n6901), .ZN(n6912) );
  AOI22_X1 U7845 ( .A1(n6906), .A2(keyinput99), .B1(keyinput81), .B2(n6905), 
        .ZN(n6904) );
  OAI221_X1 U7846 ( .B1(n6906), .B2(keyinput99), .C1(n6905), .C2(keyinput81), 
        .A(n6904), .ZN(n6911) );
  INV_X1 U7847 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n6908) );
  AOI22_X1 U7848 ( .A1(n6909), .A2(keyinput56), .B1(n6908), .B2(keyinput106), 
        .ZN(n6907) );
  OAI221_X1 U7849 ( .B1(n6909), .B2(keyinput56), .C1(n6908), .C2(keyinput106), 
        .A(n6907), .ZN(n6910) );
  NOR4_X1 U7850 ( .A1(n6913), .A2(n6912), .A3(n6911), .A4(n6910), .ZN(n6947)
         );
  INV_X1 U7851 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n6915) );
  AOI22_X1 U7852 ( .A1(n6916), .A2(keyinput17), .B1(n6915), .B2(keyinput122), 
        .ZN(n6914) );
  OAI221_X1 U7853 ( .B1(n6916), .B2(keyinput17), .C1(n6915), .C2(keyinput122), 
        .A(n6914), .ZN(n6928) );
  INV_X1 U7854 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6918) );
  AOI22_X1 U7855 ( .A1(n6919), .A2(keyinput95), .B1(n6918), .B2(keyinput49), 
        .ZN(n6917) );
  OAI221_X1 U7856 ( .B1(n6919), .B2(keyinput95), .C1(n6918), .C2(keyinput49), 
        .A(n6917), .ZN(n6927) );
  AOI22_X1 U7857 ( .A1(n6921), .A2(keyinput7), .B1(n3916), .B2(keyinput14), 
        .ZN(n6920) );
  OAI221_X1 U7858 ( .B1(n6921), .B2(keyinput7), .C1(n3916), .C2(keyinput14), 
        .A(n6920), .ZN(n6926) );
  AOI22_X1 U7859 ( .A1(n6924), .A2(keyinput118), .B1(keyinput6), .B2(n6923), 
        .ZN(n6922) );
  OAI221_X1 U7860 ( .B1(n6924), .B2(keyinput118), .C1(n6923), .C2(keyinput6), 
        .A(n6922), .ZN(n6925) );
  NOR4_X1 U7861 ( .A1(n6928), .A2(n6927), .A3(n6926), .A4(n6925), .ZN(n6946)
         );
  AOI22_X1 U7862 ( .A1(n6931), .A2(keyinput53), .B1(n6930), .B2(keyinput112), 
        .ZN(n6929) );
  OAI221_X1 U7863 ( .B1(n6931), .B2(keyinput53), .C1(n6930), .C2(keyinput112), 
        .A(n6929), .ZN(n6944) );
  AOI22_X1 U7864 ( .A1(n6934), .A2(keyinput96), .B1(n6933), .B2(keyinput73), 
        .ZN(n6932) );
  OAI221_X1 U7865 ( .B1(n6934), .B2(keyinput96), .C1(n6933), .C2(keyinput73), 
        .A(n6932), .ZN(n6943) );
  AOI22_X1 U7866 ( .A1(n6937), .A2(keyinput109), .B1(n6936), .B2(keyinput5), 
        .ZN(n6935) );
  OAI221_X1 U7867 ( .B1(n6937), .B2(keyinput109), .C1(n6936), .C2(keyinput5), 
        .A(n6935), .ZN(n6942) );
  INV_X1 U7868 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6939) );
  AOI22_X1 U7869 ( .A1(n6940), .A2(keyinput32), .B1(n6939), .B2(keyinput87), 
        .ZN(n6938) );
  OAI221_X1 U7870 ( .B1(n6940), .B2(keyinput32), .C1(n6939), .C2(keyinput87), 
        .A(n6938), .ZN(n6941) );
  NOR4_X1 U7871 ( .A1(n6944), .A2(n6943), .A3(n6942), .A4(n6941), .ZN(n6945)
         );
  NAND4_X1 U7872 ( .A1(n6948), .A2(n6947), .A3(n6946), .A4(n6945), .ZN(n7012)
         );
  AOI22_X1 U7873 ( .A1(n6951), .A2(keyinput60), .B1(n6950), .B2(keyinput58), 
        .ZN(n6949) );
  OAI221_X1 U7874 ( .B1(n6951), .B2(keyinput60), .C1(n6950), .C2(keyinput58), 
        .A(n6949), .ZN(n6962) );
  AOI22_X1 U7875 ( .A1(n6954), .A2(keyinput93), .B1(keyinput43), .B2(n6953), 
        .ZN(n6952) );
  OAI221_X1 U7876 ( .B1(n6954), .B2(keyinput93), .C1(n6953), .C2(keyinput43), 
        .A(n6952), .ZN(n6961) );
  AOI22_X1 U7877 ( .A1(n3929), .A2(keyinput105), .B1(keyinput107), .B2(n5981), 
        .ZN(n6955) );
  OAI221_X1 U7878 ( .B1(n3929), .B2(keyinput105), .C1(n5981), .C2(keyinput107), 
        .A(n6955), .ZN(n6960) );
  INV_X1 U7879 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n6957) );
  AOI22_X1 U7880 ( .A1(n6958), .A2(keyinput39), .B1(n6957), .B2(keyinput115), 
        .ZN(n6956) );
  OAI221_X1 U7881 ( .B1(n6958), .B2(keyinput39), .C1(n6957), .C2(keyinput115), 
        .A(n6956), .ZN(n6959) );
  NOR4_X1 U7882 ( .A1(n6962), .A2(n6961), .A3(n6960), .A4(n6959), .ZN(n7010)
         );
  AOI22_X1 U7883 ( .A1(n6964), .A2(keyinput0), .B1(keyinput76), .B2(n4645), 
        .ZN(n6963) );
  OAI221_X1 U7884 ( .B1(n6964), .B2(keyinput0), .C1(n4645), .C2(keyinput76), 
        .A(n6963), .ZN(n6977) );
  AOI22_X1 U7885 ( .A1(n6967), .A2(keyinput33), .B1(keyinput59), .B2(n6966), 
        .ZN(n6965) );
  OAI221_X1 U7886 ( .B1(n6967), .B2(keyinput33), .C1(n6966), .C2(keyinput59), 
        .A(n6965), .ZN(n6976) );
  AOI22_X1 U7887 ( .A1(n6970), .A2(keyinput124), .B1(keyinput100), .B2(n6969), 
        .ZN(n6968) );
  OAI221_X1 U7888 ( .B1(n6970), .B2(keyinput124), .C1(n6969), .C2(keyinput100), 
        .A(n6968), .ZN(n6975) );
  AOI22_X1 U7889 ( .A1(n6973), .A2(keyinput63), .B1(n6972), .B2(keyinput22), 
        .ZN(n6971) );
  OAI221_X1 U7890 ( .B1(n6973), .B2(keyinput63), .C1(n6972), .C2(keyinput22), 
        .A(n6971), .ZN(n6974) );
  NOR4_X1 U7891 ( .A1(n6977), .A2(n6976), .A3(n6975), .A4(n6974), .ZN(n7009)
         );
  AOI22_X1 U7892 ( .A1(n6980), .A2(keyinput104), .B1(n6979), .B2(keyinput127), 
        .ZN(n6978) );
  OAI221_X1 U7893 ( .B1(n6980), .B2(keyinput104), .C1(n6979), .C2(keyinput127), 
        .A(n6978), .ZN(n6992) );
  AOI22_X1 U7894 ( .A1(n6983), .A2(keyinput9), .B1(n6982), .B2(keyinput88), 
        .ZN(n6981) );
  OAI221_X1 U7895 ( .B1(n6983), .B2(keyinput9), .C1(n6982), .C2(keyinput88), 
        .A(n6981), .ZN(n6991) );
  INV_X1 U7896 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6985) );
  AOI22_X1 U7897 ( .A1(n3893), .A2(keyinput2), .B1(n6985), .B2(keyinput42), 
        .ZN(n6984) );
  OAI221_X1 U7898 ( .B1(n3893), .B2(keyinput2), .C1(n6985), .C2(keyinput42), 
        .A(n6984), .ZN(n6990) );
  INV_X1 U7899 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n6987) );
  AOI22_X1 U7900 ( .A1(n6988), .A2(keyinput25), .B1(n6987), .B2(keyinput34), 
        .ZN(n6986) );
  OAI221_X1 U7901 ( .B1(n6988), .B2(keyinput25), .C1(n6987), .C2(keyinput34), 
        .A(n6986), .ZN(n6989) );
  NOR4_X1 U7902 ( .A1(n6992), .A2(n6991), .A3(n6990), .A4(n6989), .ZN(n7008)
         );
  AOI22_X1 U7903 ( .A1(n6994), .A2(keyinput65), .B1(keyinput61), .B2(n4235), 
        .ZN(n6993) );
  OAI221_X1 U7904 ( .B1(n6994), .B2(keyinput65), .C1(n4235), .C2(keyinput61), 
        .A(n6993), .ZN(n7006) );
  AOI22_X1 U7905 ( .A1(n6996), .A2(keyinput83), .B1(n3904), .B2(keyinput29), 
        .ZN(n6995) );
  OAI221_X1 U7906 ( .B1(n6996), .B2(keyinput83), .C1(n3904), .C2(keyinput29), 
        .A(n6995), .ZN(n7005) );
  AOI22_X1 U7907 ( .A1(n6999), .A2(keyinput121), .B1(n6998), .B2(keyinput114), 
        .ZN(n6997) );
  OAI221_X1 U7908 ( .B1(n6999), .B2(keyinput121), .C1(n6998), .C2(keyinput114), 
        .A(n6997), .ZN(n7004) );
  AOI22_X1 U7909 ( .A1(n7002), .A2(keyinput66), .B1(keyinput102), .B2(n7001), 
        .ZN(n7000) );
  OAI221_X1 U7910 ( .B1(n7002), .B2(keyinput66), .C1(n7001), .C2(keyinput102), 
        .A(n7000), .ZN(n7003) );
  NOR4_X1 U7911 ( .A1(n7006), .A2(n7005), .A3(n7004), .A4(n7003), .ZN(n7007)
         );
  NAND4_X1 U7912 ( .A1(n7010), .A2(n7009), .A3(n7008), .A4(n7007), .ZN(n7011)
         );
  NOR3_X1 U7913 ( .A1(n7013), .A2(n7012), .A3(n7011), .ZN(n7014) );
  NAND3_X1 U7914 ( .A1(n7016), .A2(n7015), .A3(n7014), .ZN(n7017) );
  XNOR2_X1 U7915 ( .A(n7018), .B(n7017), .ZN(U3099) );
  CLKBUF_X1 U3818 ( .A(n3418), .Z(n3405) );
  AND2_X1 U3838 ( .A1(n5015), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3210)
         );
  AND4_X1 U4020 ( .A1(n3296), .A2(n3295), .A3(n3294), .A4(n3293), .ZN(n3297)
         );
  CLKBUF_X1 U4118 ( .A(n4464), .Z(n6085) );
  CLKBUF_X1 U4242 ( .A(n4552), .Z(n4619) );
endmodule

