

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, 
        P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN, 
        P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN, 
        P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN, 
        P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN, 
        P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN, 
        P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN, 
        P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN, 
        P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN, 
        P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN, 
        P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN,
         P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN,
         P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN,
         P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN,
         P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN,
         P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN,
         P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN,
         P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN,
         P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN,
         P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN,
         P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN,
         P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN,
         P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN,
         P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN,
         P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN,
         P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN,
         P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN,
         P3_ADDR_REG_3__SCAN_IN, P3_ADDR_REG_4__SCAN_IN,
         P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN,
         P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN,
         P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN,
         P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN,
         P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN,
         P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN,
         P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN,
         P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN,
         P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN,
         P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN,
         P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN,
         P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN,
         P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN,
         P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN,
         P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN,
         P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN,
         P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN,
         P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN,
         P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN,
         P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN,
         P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN,
         P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN,
         P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN,
         P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN,
         P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN,
         P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN,
         P3_REG0_REG_3__SCAN_IN, P3_REG0_REG_4__SCAN_IN,
         P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN,
         P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN,
         P3_REG0_REG_9__SCAN_IN, P3_REG0_REG_10__SCAN_IN,
         P3_REG0_REG_11__SCAN_IN, P3_REG0_REG_12__SCAN_IN,
         P3_REG0_REG_13__SCAN_IN, P3_REG0_REG_14__SCAN_IN,
         P3_REG0_REG_15__SCAN_IN, P3_REG0_REG_16__SCAN_IN,
         P3_REG0_REG_17__SCAN_IN, P3_REG0_REG_18__SCAN_IN,
         P3_REG0_REG_19__SCAN_IN, P3_REG0_REG_20__SCAN_IN,
         P3_REG0_REG_21__SCAN_IN, P3_REG0_REG_22__SCAN_IN,
         P3_REG0_REG_23__SCAN_IN, P3_REG0_REG_24__SCAN_IN,
         P3_REG0_REG_25__SCAN_IN, P3_REG0_REG_26__SCAN_IN,
         P3_REG0_REG_27__SCAN_IN, P3_REG0_REG_28__SCAN_IN,
         P3_REG0_REG_29__SCAN_IN, P3_REG0_REG_30__SCAN_IN,
         P3_REG0_REG_31__SCAN_IN, P3_REG1_REG_0__SCAN_IN,
         P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN,
         P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN,
         P3_REG1_REG_5__SCAN_IN, P3_REG1_REG_6__SCAN_IN,
         P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN,
         P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN,
         P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN,
         P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN,
         P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN,
         P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN,
         P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN,
         P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN,
         P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN,
         P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN,
         P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN,
         P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN,
         P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN,
         P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN,
         P3_REG2_REG_3__SCAN_IN, P3_REG2_REG_4__SCAN_IN,
         P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN,
         P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN,
         P3_REG2_REG_9__SCAN_IN, P3_REG2_REG_10__SCAN_IN,
         P3_REG2_REG_11__SCAN_IN, P3_REG2_REG_12__SCAN_IN,
         P3_REG2_REG_13__SCAN_IN, P3_REG2_REG_14__SCAN_IN,
         P3_REG2_REG_15__SCAN_IN, P3_REG2_REG_16__SCAN_IN,
         P3_REG2_REG_17__SCAN_IN, P3_REG2_REG_18__SCAN_IN,
         P3_REG2_REG_19__SCAN_IN, P3_REG2_REG_20__SCAN_IN,
         P3_REG2_REG_21__SCAN_IN, P3_REG2_REG_22__SCAN_IN,
         P3_REG2_REG_23__SCAN_IN, P3_REG2_REG_24__SCAN_IN,
         P3_REG2_REG_25__SCAN_IN, P3_REG2_REG_26__SCAN_IN,
         P3_REG2_REG_27__SCAN_IN, P3_REG2_REG_28__SCAN_IN,
         P3_REG2_REG_29__SCAN_IN, P3_REG2_REG_30__SCAN_IN,
         P3_REG2_REG_31__SCAN_IN, P3_ADDR_REG_19__SCAN_IN,
         P3_ADDR_REG_18__SCAN_IN, P3_ADDR_REG_17__SCAN_IN,
         P3_ADDR_REG_16__SCAN_IN, P3_ADDR_REG_15__SCAN_IN,
         P3_ADDR_REG_14__SCAN_IN, P3_ADDR_REG_13__SCAN_IN,
         P3_ADDR_REG_12__SCAN_IN, P3_ADDR_REG_11__SCAN_IN,
         P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042;

  INV_X4 U7289 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OAI21_X1 U7290 ( .B1(n13602), .B2(n8804), .A(n12698), .ZN(n8805) );
  NAND2_X1 U7291 ( .A1(n11322), .A2(n15925), .ZN(n11535) );
  CLKBUF_X2 U7292 ( .A(n10445), .Z(n7532) );
  INV_X2 U7293 ( .A(n11286), .ZN(n14208) );
  NOR2_X1 U7294 ( .A1(n15450), .A2(n7731), .ZN(n7728) );
  INV_X2 U7295 ( .A(n12956), .ZN(n12965) );
  CLKBUF_X1 U7296 ( .A(n9721), .Z(n7189) );
  CLKBUF_X1 U7298 ( .A(n8380), .Z(n7220) );
  INV_X1 U7299 ( .A(n10514), .ZN(n15739) );
  CLKBUF_X2 U7300 ( .A(n8994), .Z(n9542) );
  INV_X1 U7301 ( .A(n9546), .ZN(n8952) );
  INV_X1 U7302 ( .A(n9104), .ZN(n9571) );
  NAND2_X1 U7303 ( .A1(n8959), .A2(n10395), .ZN(n9209) );
  NAND2_X1 U7304 ( .A1(n8781), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8783) );
  INV_X1 U7305 ( .A(n10404), .ZN(n10395) );
  BUF_X1 U7307 ( .A(n9721), .Z(n14582) );
  INV_X1 U7308 ( .A(n12738), .ZN(n12727) );
  INV_X1 U7309 ( .A(n10520), .ZN(n12335) );
  NAND2_X1 U7311 ( .A1(n10431), .A2(n10697), .ZN(n10503) );
  NAND2_X1 U7312 ( .A1(n11577), .A2(n11576), .ZN(n11578) );
  AND2_X1 U7313 ( .A1(n8297), .A2(n13812), .ZN(n7250) );
  XNOR2_X1 U7314 ( .A(n7711), .B(P3_IR_REG_21__SCAN_IN), .ZN(n10612) );
  NOR2_X2 U7315 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n10264) );
  BUF_X1 U7316 ( .A(n10529), .Z(n12425) );
  INV_X1 U7317 ( .A(n9582), .ZN(n9301) );
  AND4_X1 U7318 ( .A1(n8393), .A2(n8392), .A3(n8391), .A4(n8390), .ZN(n11172)
         );
  XNOR2_X1 U7319 ( .A(n8286), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8297) );
  INV_X2 U7320 ( .A(n10612), .ZN(n12612) );
  AND3_X1 U7321 ( .A1(n7963), .A2(n7964), .A3(n7399), .ZN(n11454) );
  NAND3_X1 U7322 ( .A1(n7500), .A2(n10448), .A3(n7499), .ZN(n12780) );
  INV_X1 U7323 ( .A(n15903), .ZN(n12844) );
  INV_X1 U7324 ( .A(n8297), .ZN(n13808) );
  XNOR2_X1 U7325 ( .A(n7217), .B(n14475), .ZN(n13119) );
  OAI21_X2 U7326 ( .B1(n8020), .B2(n7446), .A(n13937), .ZN(n7445) );
  OR2_X2 U7327 ( .A1(n10262), .A2(n10251), .ZN(n10289) );
  XNOR2_X2 U7328 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n15269) );
  NAND2_X2 U7329 ( .A1(n8475), .A2(n8474), .ZN(n11993) );
  OAI21_X1 U7330 ( .B1(n14507), .B2(n14078), .A(n12766), .ZN(n7188) );
  OAI21_X1 U7331 ( .B1(n14507), .B2(n14078), .A(n12766), .ZN(n10445) );
  AOI21_X2 U7332 ( .B1(n11701), .B2(P2_REG2_REG_13__SCAN_IN), .A(n11700), .ZN(
        n14039) );
  AND2_X2 U7333 ( .A1(n14482), .A2(n13119), .ZN(n10528) );
  AOI21_X2 U7334 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n10226), .A(n10218), .ZN(
        n15358) );
  NOR2_X2 U7335 ( .A1(n8780), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n7712) );
  OAI222_X1 U7336 ( .A1(P3_U3151), .A2(n12602), .B1(n12036), .B2(n10630), .C1(
        n11729), .C2(n13810), .ZN(P3_U3275) );
  XNOR2_X2 U7337 ( .A(n8819), .B(n8818), .ZN(n11232) );
  OAI21_X2 U7338 ( .B1(n9491), .B2(n9490), .A(n9497), .ZN(n9514) );
  XNOR2_X2 U7339 ( .A(n8882), .B(n8881), .ZN(n8888) );
  OAI21_X2 U7340 ( .B1(n11949), .B2(n12654), .A(n12656), .ZN(n12139) );
  OAI222_X1 U7341 ( .A1(P3_U3151), .A2(n8787), .B1(n12036), .B2(n12035), .C1(
        n12034), .C2(n13810), .ZN(P3_U3267) );
  NAND2_X1 U7342 ( .A1(n9781), .A2(n7541), .ZN(n9721) );
  NAND2_X2 U7343 ( .A1(n8369), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7385) );
  XNOR2_X2 U7344 ( .A(n9879), .B(n9880), .ZN(n10447) );
  AOI21_X2 U7345 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(n15350), .A(n15345), .ZN(
        n10220) );
  NOR2_X2 U7346 ( .A1(n15452), .A2(n15451), .ZN(n15450) );
  OAI211_X1 U7347 ( .C1(n10126), .C2(n10275), .A(n8382), .B(n8381), .ZN(n10620) );
  NAND2_X2 U7348 ( .A1(n7676), .A2(n7675), .ZN(n10275) );
  OAI21_X1 U7349 ( .B1(n13050), .B2(n13048), .A(n8205), .ZN(n8207) );
  NOR2_X1 U7350 ( .A1(n7253), .A2(n7366), .ZN(n8272) );
  AOI211_X1 U7351 ( .C1(n15089), .C2(n14917), .A(n14865), .B(n14864), .ZN(
        n14873) );
  OAI21_X1 U7352 ( .B1(n13443), .B2(n13437), .A(n12728), .ZN(n7199) );
  NAND2_X1 U7353 ( .A1(n7195), .A2(n12705), .ZN(n13531) );
  NAND2_X1 U7354 ( .A1(n8805), .A2(n12701), .ZN(n13545) );
  OAI21_X1 U7355 ( .B1(n8722), .B2(n14499), .A(n8358), .ZN(n8733) );
  NAND2_X1 U7356 ( .A1(n7211), .A2(n7484), .ZN(n11618) );
  NAND2_X1 U7357 ( .A1(n11136), .A2(n11135), .ZN(n11302) );
  OR2_X2 U7358 ( .A1(n11535), .A2(n12857), .ZN(n11623) );
  OAI21_X2 U7359 ( .B1(n12139), .B2(n8799), .A(n8798), .ZN(n12205) );
  NAND2_X1 U7360 ( .A1(n10344), .A2(n10343), .ZN(n13239) );
  INV_X1 U7361 ( .A(n10946), .ZN(n10691) );
  INV_X1 U7362 ( .A(n13958), .ZN(n15782) );
  NAND2_X1 U7363 ( .A1(n11168), .A2(n7194), .ZN(n15713) );
  CLKBUF_X2 U7364 ( .A(n11209), .Z(n14607) );
  OR2_X1 U7365 ( .A1(n12576), .A2(n11170), .ZN(n11168) );
  AND2_X1 U7366 ( .A1(n9016), .A2(n9006), .ZN(n10534) );
  INV_X2 U7367 ( .A(n12781), .ZN(n12848) );
  NAND3_X1 U7368 ( .A1(n8376), .A2(n8375), .A3(n8267), .ZN(n13262) );
  AND3_X1 U7369 ( .A1(n8398), .A2(n8397), .A3(n8396), .ZN(n10714) );
  INV_X1 U7370 ( .A(n12602), .ZN(n12749) );
  OR2_X1 U7371 ( .A1(n8380), .A2(n9855), .ZN(n8382) );
  BUF_X1 U7373 ( .A(n8380), .Z(n7219) );
  NAND2_X1 U7374 ( .A1(n8926), .A2(n9649), .ZN(n12052) );
  NAND2_X1 U7375 ( .A1(n7601), .A2(n8887), .ZN(n8994) );
  NOR2_X1 U7376 ( .A1(n8196), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n10157) );
  AND2_X1 U7377 ( .A1(n11040), .A2(n10169), .ZN(n10171) );
  NOR2_X1 U7378 ( .A1(n9609), .A2(n9608), .ZN(n9613) );
  MUX2_X1 U7379 ( .A(n14435), .B(n14434), .S(n15974), .Z(n14436) );
  NOR2_X1 U7380 ( .A1(n14353), .A2(n14352), .ZN(n14434) );
  AND2_X1 U7381 ( .A1(n7705), .A2(n7320), .ZN(n7494) );
  AOI21_X1 U7382 ( .B1(n14422), .B2(n14363), .A(n14362), .ZN(n14364) );
  MUX2_X1 U7383 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14438), .S(n15970), .Z(
        n14362) );
  AOI21_X1 U7384 ( .B1(n7768), .B2(n7763), .A(n7306), .ZN(n7549) );
  NAND2_X1 U7385 ( .A1(n14117), .A2(n7297), .ZN(n7213) );
  AOI21_X1 U7386 ( .B1(n14137), .B2(n14267), .A(n14136), .ZN(n14360) );
  NAND2_X1 U7387 ( .A1(n13906), .A2(n13905), .ZN(n13860) );
  OAI211_X1 U7388 ( .C1(n12934), .C2(n7227), .A(n7251), .B(n12939), .ZN(n12940) );
  NAND2_X1 U7389 ( .A1(n7214), .A2(n13025), .ZN(n14117) );
  NAND2_X1 U7390 ( .A1(n14131), .A2(n14115), .ZN(n7214) );
  NAND2_X1 U7391 ( .A1(n13946), .A2(n13855), .ZN(n13906) );
  AOI21_X1 U7392 ( .B1(n14886), .B2(n14885), .A(n7784), .ZN(n7367) );
  NAND2_X1 U7393 ( .A1(n14132), .A2(n14133), .ZN(n14131) );
  NAND2_X1 U7394 ( .A1(n7551), .A2(n13870), .ZN(n13946) );
  NAND2_X1 U7395 ( .A1(n7646), .A2(n7303), .ZN(n14839) );
  MUX2_X1 U7396 ( .A(n13685), .B(n13754), .S(n15940), .Z(n13686) );
  NAND2_X1 U7397 ( .A1(n14150), .A2(n12420), .ZN(n14132) );
  MUX2_X1 U7398 ( .A(n13755), .B(n13754), .S(n15944), .Z(n13756) );
  AOI21_X1 U7399 ( .B1(n15891), .B2(n13680), .A(n13679), .ZN(n13681) );
  AND2_X1 U7400 ( .A1(n13851), .A2(n8002), .ZN(n7551) );
  NAND2_X1 U7401 ( .A1(n14924), .A2(n14923), .ZN(n14922) );
  AND2_X1 U7402 ( .A1(n14946), .A2(n12521), .ZN(n14924) );
  NAND2_X1 U7403 ( .A1(n14166), .A2(n14147), .ZN(n7939) );
  NAND2_X1 U7404 ( .A1(n14221), .A2(n7226), .ZN(n7945) );
  NAND2_X1 U7405 ( .A1(n13846), .A2(n13845), .ZN(n13848) );
  AND2_X1 U7406 ( .A1(n13452), .A2(n13451), .ZN(n8260) );
  OR2_X1 U7407 ( .A1(n13202), .A2(n13089), .ZN(n13093) );
  AOI21_X1 U7408 ( .B1(n7239), .B2(n7208), .A(n12400), .ZN(n7207) );
  INV_X1 U7409 ( .A(n7239), .ZN(n7209) );
  NAND2_X1 U7410 ( .A1(n7197), .A2(n12717), .ZN(n13492) );
  NAND2_X1 U7411 ( .A1(n14998), .A2(n14997), .ZN(n14996) );
  OR2_X1 U7412 ( .A1(n13479), .A2(n13449), .ZN(n13452) );
  INV_X1 U7413 ( .A(n7226), .ZN(n7208) );
  NAND2_X1 U7414 ( .A1(n8162), .A2(n8161), .ZN(n13193) );
  NAND2_X1 U7415 ( .A1(n14287), .A2(n12331), .ZN(n12333) );
  NAND2_X1 U7416 ( .A1(n7198), .A2(n8807), .ZN(n13512) );
  NAND2_X1 U7417 ( .A1(n13965), .A2(n13964), .ZN(n13963) );
  NAND2_X1 U7418 ( .A1(n14310), .A2(n12323), .ZN(n14287) );
  OAI22_X1 U7419 ( .A1(n13984), .A2(n8013), .B1(n8015), .B2(n8012), .ZN(n13965) );
  NAND2_X1 U7420 ( .A1(n7212), .A2(n14313), .ZN(n14310) );
  NOR2_X1 U7421 ( .A1(n14193), .A2(n14171), .ZN(n12400) );
  NAND2_X1 U7422 ( .A1(n14307), .A2(n14305), .ZN(n7212) );
  OAI21_X1 U7423 ( .B1(n8021), .B2(n7446), .A(n7444), .ZN(n13935) );
  NAND2_X1 U7424 ( .A1(n13531), .A2(n13532), .ZN(n8806) );
  OR2_X1 U7425 ( .A1(n14531), .A2(n14530), .ZN(n8261) );
  NAND2_X1 U7426 ( .A1(n7382), .A2(n7937), .ZN(n14307) );
  NAND2_X1 U7427 ( .A1(n12363), .A2(n12362), .ZN(n14456) );
  AND2_X1 U7428 ( .A1(n13365), .A2(n13385), .ZN(n13366) );
  NAND2_X1 U7429 ( .A1(n7384), .A2(n7383), .ZN(n12058) );
  NAND2_X1 U7430 ( .A1(n8733), .A2(n8732), .ZN(n8735) );
  NAND2_X1 U7431 ( .A1(n14629), .A2(n14525), .ZN(n14529) );
  NAND2_X1 U7432 ( .A1(n13364), .A2(n13379), .ZN(n13385) );
  NAND2_X1 U7433 ( .A1(n12325), .A2(n12324), .ZN(n14408) );
  NAND2_X1 U7434 ( .A1(n14518), .A2(n7284), .ZN(n14629) );
  NAND2_X1 U7435 ( .A1(n12338), .A2(n12337), .ZN(n14461) );
  NAND2_X1 U7436 ( .A1(n8358), .A2(n8357), .ZN(n8722) );
  OR2_X1 U7437 ( .A1(n8356), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U7438 ( .A1(n11618), .A2(n11617), .ZN(n7926) );
  NAND2_X1 U7439 ( .A1(n12190), .A2(n12191), .ZN(n14321) );
  NAND2_X1 U7440 ( .A1(n13635), .A2(n13638), .ZN(n8801) );
  NOR2_X1 U7441 ( .A1(n12224), .A2(n12223), .ZN(n12285) );
  NAND2_X1 U7442 ( .A1(n12322), .A2(n12321), .ZN(n14320) );
  NOR2_X1 U7443 ( .A1(n12016), .A2(n12230), .ZN(n12224) );
  NAND2_X1 U7444 ( .A1(n11136), .A2(n7210), .ZN(n7211) );
  NAND2_X1 U7445 ( .A1(n12172), .A2(n12171), .ZN(n14471) );
  AND2_X1 U7446 ( .A1(n11135), .A2(n11527), .ZN(n7210) );
  NOR2_X2 U7447 ( .A1(n12865), .A2(n11623), .ZN(n11985) );
  AND2_X1 U7448 ( .A1(n7478), .A2(n7477), .ZN(n14028) );
  NAND2_X1 U7449 ( .A1(n7495), .A2(n9310), .ZN(n9325) );
  NAND2_X1 U7450 ( .A1(n12057), .A2(n12056), .ZN(n12877) );
  NAND2_X1 U7451 ( .A1(n7372), .A2(n7370), .ZN(n11074) );
  NAND2_X1 U7452 ( .A1(n11982), .A2(n11981), .ZN(n12873) );
  OR2_X1 U7453 ( .A1(n11027), .A2(n11007), .ZN(n7372) );
  NAND2_X1 U7454 ( .A1(n11300), .A2(n11299), .ZN(n12851) );
  NAND2_X1 U7455 ( .A1(n7215), .A2(n11006), .ZN(n11027) );
  AND2_X1 U7456 ( .A1(n7707), .A2(n11125), .ZN(n15903) );
  NAND2_X1 U7457 ( .A1(n11991), .A2(n12649), .ZN(n11949) );
  NAND2_X1 U7458 ( .A1(n12137), .A2(n8519), .ZN(n12201) );
  OR2_X1 U7459 ( .A1(n12135), .A2(n12658), .ZN(n12137) );
  NOR2_X1 U7460 ( .A1(n15459), .A2(n15296), .ZN(n15463) );
  NAND2_X1 U7461 ( .A1(n11992), .A2(n12647), .ZN(n11991) );
  AND2_X1 U7462 ( .A1(n14001), .A2(n12771), .ZN(n7205) );
  NAND2_X1 U7463 ( .A1(n11633), .A2(n8797), .ZN(n11992) );
  NAND2_X1 U7464 ( .A1(n10872), .A2(n7242), .ZN(n10876) );
  NAND2_X1 U7465 ( .A1(n11634), .A2(n12642), .ZN(n11633) );
  AOI21_X1 U7466 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n11124), .A(n10896), .ZN(
        n10900) );
  OR2_X1 U7467 ( .A1(n10428), .A2(n10427), .ZN(n9727) );
  AOI21_X1 U7468 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n11124), .A(n10903), .ZN(
        n10906) );
  NAND2_X1 U7469 ( .A1(n11190), .A2(n12629), .ZN(n11240) );
  INV_X1 U7470 ( .A(n7203), .ZN(P2_U3532) );
  NAND2_X1 U7471 ( .A1(n9134), .A2(n9133), .ZN(n9138) );
  AOI21_X1 U7472 ( .B1(n14025), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n7204), .ZN(
        n7203) );
  NAND2_X1 U7473 ( .A1(n11191), .A2(n12626), .ZN(n11190) );
  AND2_X1 U7474 ( .A1(n12666), .A2(n12668), .ZN(n12664) );
  NAND2_X1 U7475 ( .A1(n7369), .A2(n10831), .ZN(n7216) );
  NAND2_X1 U7476 ( .A1(n7196), .A2(n12623), .ZN(n11191) );
  NAND2_X1 U7477 ( .A1(n11055), .A2(n11054), .ZN(n7196) );
  NAND2_X1 U7478 ( .A1(n9051), .A2(n9050), .ZN(n10995) );
  NAND2_X1 U7479 ( .A1(n7262), .A2(n7191), .ZN(n7190) );
  INV_X1 U7480 ( .A(n7262), .ZN(n7192) );
  NOR2_X1 U7481 ( .A1(n10625), .A2(n10624), .ZN(n13223) );
  NAND2_X1 U7482 ( .A1(n15713), .A2(n15715), .ZN(n15712) );
  NOR2_X1 U7483 ( .A1(n10668), .A2(n7202), .ZN(n7201) );
  NAND2_X1 U7484 ( .A1(n12994), .A2(n11098), .ZN(n11097) );
  NAND2_X1 U7485 ( .A1(n10829), .A2(n10828), .ZN(n11098) );
  NAND2_X1 U7486 ( .A1(n10535), .A2(n10536), .ZN(n13958) );
  AND3_X1 U7487 ( .A1(n8518), .A2(n8517), .A3(n8516), .ZN(n15892) );
  OR2_X1 U7488 ( .A1(n12992), .A2(n10417), .ZN(n10829) );
  AND2_X1 U7489 ( .A1(n12649), .A2(n12650), .ZN(n12647) );
  AOI21_X1 U7490 ( .B1(n12619), .B2(n7194), .A(n12738), .ZN(n12620) );
  AND2_X1 U7491 ( .A1(n14262), .A2(n7200), .ZN(n7202) );
  NAND2_X1 U7492 ( .A1(n10524), .A2(n10523), .ZN(n12794) );
  AND2_X1 U7493 ( .A1(n10957), .A2(n10815), .ZN(n12994) );
  INV_X1 U7494 ( .A(n12629), .ZN(n7191) );
  AND2_X1 U7495 ( .A1(n9837), .A2(n9735), .ZN(n11209) );
  INV_X4 U7496 ( .A(n12208), .ZN(n11286) );
  NAND2_X1 U7497 ( .A1(n10399), .A2(n10828), .ZN(n12992) );
  INV_X2 U7498 ( .A(n9741), .ZN(n14661) );
  INV_X1 U7499 ( .A(n9721), .ZN(n14615) );
  NAND2_X1 U7500 ( .A1(n9016), .A2(n9015), .ZN(n9020) );
  NAND2_X1 U7501 ( .A1(n7206), .A2(n10440), .ZN(n10399) );
  INV_X1 U7502 ( .A(n12780), .ZN(n15749) );
  NAND4_X1 U7503 ( .A1(n10465), .A2(n10464), .A3(n10463), .A4(n10462), .ZN(
        n14023) );
  INV_X1 U7504 ( .A(n10812), .ZN(n7206) );
  NAND4_X2 U7505 ( .A1(n8999), .A2(n8998), .A3(n8997), .A4(n8996), .ZN(n14748)
         );
  NAND4_X1 U7506 ( .A1(n10533), .A2(n10532), .A3(n10531), .A4(n7252), .ZN(
        n14022) );
  NAND4_X2 U7507 ( .A1(n9037), .A2(n9036), .A3(n9035), .A4(n9034), .ZN(n14747)
         );
  AND3_X1 U7508 ( .A1(n8424), .A2(n8423), .A3(n8422), .ZN(n15772) );
  AND2_X1 U7509 ( .A1(n9706), .A2(n12052), .ZN(n10060) );
  AND4_X1 U7510 ( .A1(n8893), .A2(n8892), .A3(n8891), .A4(n8890), .ZN(n10146)
         );
  AND3_X1 U7511 ( .A1(n8411), .A2(n8410), .A3(n8409), .ZN(n11186) );
  NAND4_X1 U7512 ( .A1(n8956), .A2(n8955), .A3(n8954), .A4(n8953), .ZN(n14750)
         );
  AND4_X1 U7513 ( .A1(n8403), .A2(n8402), .A3(n8401), .A4(n8400), .ZN(n15722)
         );
  AND3_X1 U7514 ( .A1(n8441), .A2(n8440), .A3(n8439), .ZN(n11242) );
  AND4_X1 U7515 ( .A1(n8433), .A2(n8432), .A3(n8431), .A4(n8430), .ZN(n11226)
         );
  NAND4_X1 U7516 ( .A1(n10403), .A2(n10402), .A3(n10401), .A4(n10400), .ZN(
        n12772) );
  NAND2_X1 U7517 ( .A1(n9702), .A2(n9781), .ZN(n14583) );
  CLKBUF_X1 U7518 ( .A(n10528), .Z(n7508) );
  INV_X2 U7519 ( .A(n12960), .ZN(n12336) );
  OR2_X1 U7520 ( .A1(n8404), .A2(n9854), .ZN(n8381) );
  AND2_X2 U7521 ( .A1(n13808), .A2(n8289), .ZN(n8520) );
  AND2_X1 U7522 ( .A1(n10390), .A2(n10389), .ZN(n10529) );
  CLKBUF_X3 U7523 ( .A(n8543), .Z(n8524) );
  CLKBUF_X3 U7524 ( .A(n8404), .Z(n7221) );
  INV_X2 U7525 ( .A(n9209), .ZN(n9595) );
  AND2_X1 U7526 ( .A1(n13119), .A2(n10390), .ZN(n10459) );
  OR2_X1 U7527 ( .A1(n13119), .A2(n10390), .ZN(n10460) );
  XNOR2_X1 U7528 ( .A(n10376), .B(P2_IR_REG_21__SCAN_IN), .ZN(n13030) );
  NAND2_X1 U7529 ( .A1(n8196), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10376) );
  NAND2_X1 U7530 ( .A1(n8924), .A2(n8922), .ZN(n9649) );
  AOI21_X1 U7531 ( .B1(n7571), .B2(n7578), .A(n7569), .ZN(n7568) );
  XNOR2_X1 U7532 ( .A(n8916), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9348) );
  INV_X2 U7533 ( .A(n13798), .ZN(n12036) );
  XNOR2_X1 U7534 ( .A(n8288), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8289) );
  NAND2_X1 U7535 ( .A1(n13801), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8286) );
  OAI21_X1 U7536 ( .B1(n9288), .B2(n9881), .A(n7540), .ZN(n9043) );
  NAND2_X1 U7537 ( .A1(n14474), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7217) );
  NAND2_X2 U7538 ( .A1(n10395), .A2(P1_U3086), .ZN(n15215) );
  XNOR2_X1 U7539 ( .A(n10383), .B(P2_IR_REG_19__SCAN_IN), .ZN(n14078) );
  NAND2_X1 U7540 ( .A1(n7498), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8819) );
  NAND2_X1 U7541 ( .A1(n10171), .A2(n7944), .ZN(n14474) );
  MUX2_X1 U7543 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8884), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n8886) );
  AND2_X1 U7544 ( .A1(n8645), .A2(n8644), .ZN(n8661) );
  NAND2_X1 U7545 ( .A1(n9288), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7540) );
  XNOR2_X1 U7546 ( .A(n7386), .B(n8371), .ZN(n8788) );
  OR2_X1 U7547 ( .A1(n8287), .A2(n8554), .ZN(n8288) );
  INV_X4 U7548 ( .A(n9311), .ZN(n10404) );
  INV_X2 U7549 ( .A(n9311), .ZN(n9288) );
  NOR2_X1 U7550 ( .A1(n8816), .A2(n7910), .ZN(n8287) );
  INV_X1 U7551 ( .A(n8464), .ZN(n7919) );
  NAND2_X1 U7552 ( .A1(n7808), .A2(n7807), .ZN(n8899) );
  NAND2_X1 U7553 ( .A1(n7266), .A2(n7232), .ZN(n8464) );
  AND3_X1 U7554 ( .A1(n7193), .A2(n8282), .A3(n8281), .ZN(n8283) );
  NAND2_X1 U7555 ( .A1(n15272), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n15271) );
  AND4_X1 U7556 ( .A1(n8278), .A2(n8564), .A3(n8529), .A4(n8566), .ZN(n8279)
         );
  AND2_X1 U7557 ( .A1(n8877), .A2(n8917), .ZN(n7718) );
  AND4_X1 U7558 ( .A1(n7871), .A2(n7392), .A3(n8277), .A4(n8449), .ZN(n7232)
         );
  AND2_X1 U7559 ( .A1(n8280), .A2(n8782), .ZN(n7193) );
  AND2_X1 U7560 ( .A1(n9673), .A2(n9672), .ZN(n7378) );
  AND4_X1 U7561 ( .A1(n8873), .A2(n8874), .A3(n8875), .A4(n9210), .ZN(n7719)
         );
  INV_X1 U7562 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10263) );
  INV_X1 U7563 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8566) );
  INV_X1 U7564 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8564) );
  INV_X1 U7565 ( .A(P2_RD_REG_SCAN_IN), .ZN(n15675) );
  INV_X1 U7566 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8449) );
  INV_X1 U7567 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8529) );
  INV_X1 U7568 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n10164) );
  INV_X1 U7569 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7392) );
  NOR2_X1 U7570 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n8919) );
  INV_X1 U7571 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7871) );
  NOR2_X2 U7572 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n8907) );
  NOR2_X1 U7573 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n8281) );
  INV_X1 U7574 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n15326) );
  NOR2_X1 U7575 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n8282) );
  INV_X1 U7576 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8818) );
  NOR2_X1 U7577 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n10281) );
  INV_X4 U7578 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7579 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n9676) );
  NOR2_X1 U7580 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n9675) );
  NOR2_X1 U7581 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n9674) );
  NOR2_X2 U7582 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n9846) );
  NOR2_X1 U7583 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8278) );
  OAI211_X2 U7584 ( .C1(n11190), .C2(n7192), .A(n7746), .B(n7190), .ZN(n11634)
         );
  NAND4_X2 U7585 ( .A1(n7919), .A2(n8820), .A3(n7238), .A4(n8166), .ZN(n8816)
         );
  AND3_X2 U7586 ( .A1(n8283), .A2(n7917), .A3(n7319), .ZN(n7238) );
  NAND2_X1 U7587 ( .A1(n12618), .A2(n7194), .ZN(n12576) );
  NAND2_X1 U7588 ( .A1(n15720), .A2(n10620), .ZN(n7194) );
  NAND2_X1 U7589 ( .A1(n13545), .A2(n13546), .ZN(n7195) );
  OAI21_X1 U7590 ( .B1(n11055), .B2(n11054), .A(n7196), .ZN(n11062) );
  NAND2_X1 U7591 ( .A1(n13512), .A2(n13505), .ZN(n7197) );
  NAND2_X1 U7592 ( .A1(n13523), .A2(n13524), .ZN(n7198) );
  OR2_X1 U7593 ( .A1(n7199), .A2(n12596), .ZN(n7768) );
  XNOR2_X1 U7594 ( .A(n7199), .B(n12732), .ZN(n13428) );
  OAI21_X2 U7596 ( .B1(n8801), .B2(n7754), .A(n7245), .ZN(n13600) );
  NAND2_X1 U7597 ( .A1(n7397), .A2(n12676), .ZN(n13635) );
  CLKBUF_X1 U7598 ( .A(n7206), .Z(n7200) );
  NAND2_X1 U7599 ( .A1(n7206), .A2(n12208), .ZN(n10441) );
  NAND2_X1 U7600 ( .A1(n14242), .A2(n7200), .ZN(n10466) );
  NAND2_X1 U7601 ( .A1(n12848), .A2(n7200), .ZN(n12765) );
  AOI22_X1 U7602 ( .A1(n12848), .A2(n12776), .B1(n12781), .B2(n7200), .ZN(
        n12777) );
  NOR2_X1 U7603 ( .A1(n14025), .A2(n10812), .ZN(n7204) );
  AOI21_X1 U7604 ( .B1(n10490), .B2(n7200), .A(n7205), .ZN(n10488) );
  OAI21_X2 U7605 ( .B1(n14221), .B2(n7209), .A(n7207), .ZN(n14166) );
  NAND2_X2 U7606 ( .A1(n11076), .A2(n11075), .ZN(n11136) );
  NAND2_X1 U7607 ( .A1(n7213), .A2(n14309), .ZN(n7523) );
  NAND2_X1 U7608 ( .A1(n11005), .A2(n12999), .ZN(n7215) );
  OAI21_X1 U7609 ( .B1(n10939), .B2(n7216), .A(n10932), .ZN(n10934) );
  NAND2_X1 U7610 ( .A1(n7216), .A2(n10939), .ZN(n10932) );
  NAND2_X1 U7611 ( .A1(n11097), .A2(n10957), .ZN(n10830) );
  OR2_X2 U7612 ( .A1(n15089), .A2(n15088), .ZN(n7253) );
  NOR2_X1 U7613 ( .A1(n9856), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n7475) );
  NOR2_X1 U7614 ( .A1(n9856), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n7447) );
  NOR2_X2 U7615 ( .A1(n14206), .A2(n14193), .ZN(n14196) );
  XNOR2_X2 U7616 ( .A(n10173), .B(n10172), .ZN(n10179) );
  AOI21_X2 U7617 ( .B1(n12084), .B2(n12083), .A(n12082), .ZN(n12085) );
  INV_X4 U7618 ( .A(n12066), .ZN(n12468) );
  INV_X1 U7619 ( .A(n13106), .ZN(n7218) );
  AND2_X1 U7620 ( .A1(n8888), .A2(n8887), .ZN(n9056) );
  NAND2_X1 U7621 ( .A1(n10126), .A2(n10395), .ZN(n8380) );
  AND2_X4 U7622 ( .A1(n8297), .A2(n8289), .ZN(n8543) );
  NAND2_X1 U7623 ( .A1(n10126), .A2(n10404), .ZN(n8404) );
  AND2_X1 U7624 ( .A1(n13808), .A2(n8289), .ZN(n7222) );
  AND2_X1 U7625 ( .A1(n13808), .A2(n8289), .ZN(n7223) );
  XNOR2_X2 U7626 ( .A(n7385), .B(n8370), .ZN(n8787) );
  OR2_X1 U7627 ( .A1(n14341), .A2(n13865), .ZN(n12455) );
  INV_X1 U7628 ( .A(n9386), .ZN(n9387) );
  AND4_X1 U7629 ( .A1(n8268), .A2(n10168), .A3(n10167), .A4(n10166), .ZN(
        n10169) );
  NOR2_X1 U7630 ( .A1(n12513), .A2(n8192), .ZN(n8191) );
  INV_X1 U7631 ( .A(n8266), .ZN(n8192) );
  NAND2_X1 U7632 ( .A1(n14892), .A2(n8195), .ZN(n8193) );
  NAND2_X1 U7633 ( .A1(n7789), .A2(n7795), .ZN(n9376) );
  NAND2_X1 U7634 ( .A1(n9329), .A2(n7790), .ZN(n7789) );
  NAND2_X1 U7635 ( .A1(n7797), .A2(n7791), .ZN(n7790) );
  INV_X1 U7636 ( .A(n7342), .ZN(n7791) );
  AOI21_X1 U7637 ( .B1(n9044), .B2(n9078), .A(n7411), .ZN(n8187) );
  AND2_X1 U7638 ( .A1(n13057), .A2(n13030), .ZN(n10456) );
  INV_X1 U7639 ( .A(n7508), .ZN(n12471) );
  AND2_X1 U7640 ( .A1(n12455), .A2(n12453), .ZN(n14094) );
  INV_X2 U7641 ( .A(n10521), .ZN(n12959) );
  NAND2_X1 U7642 ( .A1(n16027), .A2(n16001), .ZN(n7989) );
  OAI21_X1 U7643 ( .B1(n12807), .B2(n12920), .A(n12806), .ZN(n12808) );
  NAND2_X1 U7644 ( .A1(n12805), .A2(n12804), .ZN(n12810) );
  NAND2_X1 U7645 ( .A1(n12813), .A2(n12812), .ZN(n12817) );
  NOR2_X1 U7646 ( .A1(n7602), .A2(n7610), .ZN(n7608) );
  INV_X1 U7647 ( .A(n9172), .ZN(n7610) );
  AND2_X1 U7648 ( .A1(n9173), .A2(n7603), .ZN(n7602) );
  NAND2_X1 U7649 ( .A1(n8209), .A2(n7247), .ZN(n8208) );
  NAND2_X1 U7650 ( .A1(n7619), .A2(n7620), .ZN(n9246) );
  AND2_X1 U7651 ( .A1(n7459), .A2(n7456), .ZN(n7455) );
  INV_X1 U7652 ( .A(n12893), .ZN(n7459) );
  NAND2_X1 U7653 ( .A1(n12894), .A2(n7273), .ZN(n7456) );
  AOI22_X1 U7654 ( .A1(n14408), .A2(n12956), .B1(n14008), .B2(n12965), .ZN(
        n12893) );
  NAND2_X1 U7655 ( .A1(n12917), .A2(n12919), .ZN(n8211) );
  OAI21_X1 U7656 ( .B1(n7863), .B2(n7224), .A(n9818), .ZN(n7858) );
  OAI22_X1 U7657 ( .A1(n14372), .A2(n12956), .B1(n14188), .B2(n12920), .ZN(
        n12929) );
  OAI21_X1 U7658 ( .B1(n7977), .B2(n9800), .A(n10787), .ZN(n7364) );
  NAND2_X1 U7659 ( .A1(n13313), .A2(n13314), .ZN(n13339) );
  OR2_X1 U7660 ( .A1(n13116), .A2(n13456), .ZN(n12728) );
  OR2_X1 U7661 ( .A1(n13217), .A2(n13457), .ZN(n12603) );
  NAND2_X1 U7662 ( .A1(n8721), .A2(n7882), .ZN(n7881) );
  NOR2_X1 U7663 ( .A1(n8731), .A2(n7883), .ZN(n7882) );
  INV_X1 U7664 ( .A(n8720), .ZN(n7883) );
  OR2_X1 U7665 ( .A1(n13688), .A2(n13495), .ZN(n8810) );
  NOR2_X1 U7666 ( .A1(n8709), .A2(n7876), .ZN(n7875) );
  INV_X1 U7667 ( .A(n8698), .ZN(n7876) );
  INV_X1 U7668 ( .A(n8685), .ZN(n7879) );
  INV_X1 U7669 ( .A(n13578), .ZN(n7916) );
  INV_X1 U7670 ( .A(n7891), .ZN(n7887) );
  AND2_X1 U7671 ( .A1(n13623), .A2(n8591), .ZN(n12584) );
  AOI21_X1 U7672 ( .B1(n7760), .B2(n7762), .A(n7758), .ZN(n7757) );
  INV_X1 U7673 ( .A(n12672), .ZN(n7758) );
  INV_X1 U7674 ( .A(n12647), .ZN(n7908) );
  OAI21_X1 U7675 ( .B1(n8816), .B2(P3_IR_REG_26__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7386) );
  INV_X1 U7676 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8280) );
  OAI21_X1 U7677 ( .B1(n8643), .B2(n7567), .A(n7564), .ZN(n8344) );
  INV_X1 U7678 ( .A(n8656), .ZN(n7567) );
  AOI21_X1 U7679 ( .B1(n8656), .B2(n7566), .A(n7565), .ZN(n7564) );
  INV_X1 U7680 ( .A(n8343), .ZN(n7565) );
  AOI21_X1 U7681 ( .B1(n8434), .B2(n7577), .A(n7576), .ZN(n7575) );
  INV_X1 U7682 ( .A(n8314), .ZN(n7576) );
  INV_X1 U7683 ( .A(n8311), .ZN(n7577) );
  AND2_X1 U7684 ( .A1(n8022), .A2(n8025), .ZN(n8020) );
  INV_X1 U7685 ( .A(n13916), .ZN(n8025) );
  NAND2_X1 U7686 ( .A1(n12333), .A2(n7947), .ZN(n14261) );
  NOR2_X1 U7687 ( .A1(n14258), .A2(n7948), .ZN(n7947) );
  INV_X1 U7688 ( .A(n12332), .ZN(n7948) );
  NAND2_X1 U7689 ( .A1(n7926), .A2(n13009), .ZN(n11979) );
  AND2_X1 U7690 ( .A1(n11617), .A2(n11517), .ZN(n13008) );
  NOR2_X2 U7691 ( .A1(n12076), .A2(n12877), .ZN(n12190) );
  NAND2_X1 U7692 ( .A1(n8088), .A2(n9750), .ZN(n8087) );
  NOR2_X1 U7693 ( .A1(n7986), .A2(n7985), .ZN(n7984) );
  INV_X1 U7694 ( .A(n12519), .ZN(n7985) );
  INV_X1 U7695 ( .A(n7852), .ZN(n7851) );
  OAI21_X1 U7696 ( .B1(n7854), .B2(n7853), .A(n11483), .ZN(n7852) );
  NAND2_X1 U7697 ( .A1(n14886), .A2(n7782), .ZN(n7779) );
  AOI21_X1 U7698 ( .B1(n14938), .B2(n14937), .A(n12512), .ZN(n14914) );
  AND2_X1 U7699 ( .A1(n12758), .A2(n14757), .ZN(n7868) );
  INV_X1 U7700 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8879) );
  OAI22_X1 U7701 ( .A1(n9514), .A2(n9513), .B1(n9512), .B2(n11714), .ZN(n9553)
         );
  INV_X1 U7702 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8897) );
  XNOR2_X1 U7703 ( .A(n9553), .B(n9551), .ZN(n9529) );
  NOR2_X1 U7704 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n8001) );
  INV_X1 U7705 ( .A(n8178), .ZN(n8177) );
  OAI21_X1 U7706 ( .B1(n8180), .B2(n8179), .A(n9395), .ZN(n8178) );
  OR2_X1 U7707 ( .A1(n9376), .A2(n9375), .ZN(n8183) );
  INV_X1 U7708 ( .A(n9290), .ZN(n7655) );
  NOR2_X1 U7709 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n7651) );
  NOR2_X1 U7710 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n7652) );
  NOR2_X1 U7711 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n7653) );
  NAND2_X1 U7712 ( .A1(n7804), .A2(n9164), .ZN(n7803) );
  AND2_X1 U7713 ( .A1(n7802), .A2(n9189), .ZN(n7801) );
  OR2_X1 U7714 ( .A1(n9129), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n9166) );
  NAND2_X1 U7715 ( .A1(n7412), .A2(n9098), .ZN(n7411) );
  NAND2_X1 U7716 ( .A1(n7414), .A2(n7413), .ZN(n7412) );
  AND2_X1 U7717 ( .A1(n8907), .A2(n8872), .ZN(n8909) );
  INV_X1 U7718 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8872) );
  NAND2_X1 U7719 ( .A1(n13096), .A2(n13486), .ZN(n13155) );
  AOI21_X1 U7720 ( .B1(n11045), .B2(n10875), .A(n11048), .ZN(n8159) );
  NAND2_X1 U7721 ( .A1(n13172), .A2(n8163), .ZN(n8162) );
  NOR2_X1 U7722 ( .A1(n13071), .A2(n8164), .ZN(n8163) );
  INV_X1 U7723 ( .A(n8165), .ZN(n8164) );
  NAND2_X1 U7724 ( .A1(n13158), .A2(n13103), .ZN(n13219) );
  OAI21_X1 U7725 ( .B1(n13421), .B2(n13423), .A(n12563), .ZN(n12600) );
  AND4_X1 U7726 ( .A1(n8575), .A2(n8574), .A3(n8573), .A4(n8572), .ZN(n12306)
         );
  INV_X1 U7727 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8277) );
  INV_X1 U7728 ( .A(n13407), .ZN(n13419) );
  OR2_X1 U7729 ( .A1(n8585), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8614) );
  OR2_X1 U7730 ( .A1(n13789), .A2(n13641), .ZN(n12684) );
  OR2_X1 U7731 ( .A1(n13793), .A2(n13656), .ZN(n13623) );
  INV_X1 U7732 ( .A(n15719), .ZN(n13640) );
  INV_X1 U7733 ( .A(n7220), .ZN(n12560) );
  AND2_X1 U7734 ( .A1(n10336), .A2(n13796), .ZN(n10355) );
  INV_X1 U7735 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7911) );
  OAI21_X1 U7736 ( .B1(n8676), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n8346), .ZN(
        n8688) );
  AND2_X1 U7737 ( .A1(n8339), .A2(n8338), .ZN(n8623) );
  AOI21_X1 U7738 ( .B1(n8607), .B2(n7562), .A(n7561), .ZN(n7560) );
  INV_X1 U7739 ( .A(n8337), .ZN(n7561) );
  INV_X1 U7740 ( .A(n8335), .ZN(n7562) );
  INV_X1 U7741 ( .A(n8607), .ZN(n7563) );
  OAI21_X1 U7742 ( .B1(n8330), .B2(n7823), .A(n7822), .ZN(n8579) );
  AOI21_X1 U7743 ( .B1(n8331), .B2(n10333), .A(n7824), .ZN(n7822) );
  INV_X1 U7744 ( .A(n8576), .ZN(n7824) );
  NAND2_X1 U7745 ( .A1(n8453), .A2(n8315), .ZN(n7836) );
  XNOR2_X1 U7746 ( .A(n13848), .B(n13849), .ZN(n13872) );
  NAND2_X1 U7747 ( .A1(n8034), .A2(n8032), .ZN(n8031) );
  INV_X1 U7748 ( .A(n11289), .ZN(n8032) );
  OR2_X1 U7749 ( .A1(n11955), .A2(n8033), .ZN(n8030) );
  AND2_X1 U7750 ( .A1(n11956), .A2(n11566), .ZN(n8033) );
  NAND2_X1 U7751 ( .A1(n13850), .A2(n13849), .ZN(n13851) );
  NAND2_X1 U7752 ( .A1(n13872), .A2(n13871), .ZN(n13870) );
  NAND2_X1 U7753 ( .A1(n7437), .A2(n7268), .ZN(n7436) );
  OR2_X1 U7754 ( .A1(n11698), .A2(n11697), .ZN(n7478) );
  NAND2_X1 U7755 ( .A1(n12473), .A2(n12472), .ZN(n12474) );
  INV_X1 U7756 ( .A(n8075), .ZN(n8074) );
  AOI21_X1 U7757 ( .B1(n8075), .B2(n8073), .A(n7294), .ZN(n8072) );
  NOR2_X1 U7758 ( .A1(n13025), .A2(n7280), .ZN(n8075) );
  AOI21_X1 U7759 ( .B1(n12486), .B2(n8063), .A(n8062), .ZN(n8061) );
  NOR2_X1 U7760 ( .A1(n14213), .A2(n8064), .ZN(n8063) );
  OAI22_X1 U7761 ( .A1(n14213), .A2(n12488), .B1(n14223), .B2(n14212), .ZN(
        n8062) );
  NAND2_X1 U7762 ( .A1(n7839), .A2(n7838), .ZN(n14247) );
  AND2_X1 U7763 ( .A1(n13014), .A2(n7938), .ZN(n7937) );
  NAND2_X1 U7764 ( .A1(n12058), .A2(n12175), .ZN(n7382) );
  NAND2_X1 U7765 ( .A1(n12074), .A2(n12175), .ZN(n7938) );
  NAND2_X1 U7766 ( .A1(n11519), .A2(n11518), .ZN(n11607) );
  NAND2_X1 U7767 ( .A1(n11122), .A2(n8077), .ZN(n8076) );
  NOR2_X1 U7768 ( .A1(n11314), .A2(n8078), .ZN(n8077) );
  INV_X1 U7769 ( .A(n11121), .ZN(n8078) );
  CLKBUF_X1 U7770 ( .A(n14267), .Z(n14309) );
  AND2_X1 U7771 ( .A1(n10170), .A2(n10172), .ZN(n8054) );
  NAND2_X1 U7772 ( .A1(n10174), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10173) );
  NAND2_X1 U7773 ( .A1(n9687), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9690) );
  NAND2_X1 U7774 ( .A1(n9695), .A2(n9694), .ZN(n9687) );
  XNOR2_X1 U7775 ( .A(n9697), .B(n10164), .ZN(n13051) );
  NOR2_X1 U7776 ( .A1(n9738), .A2(n9737), .ZN(n9734) );
  NAND2_X1 U7777 ( .A1(n7601), .A2(n15200), .ZN(n9031) );
  NOR3_X1 U7778 ( .A1(n14906), .A2(n7723), .A3(n7724), .ZN(n14849) );
  OR2_X1 U7779 ( .A1(n15081), .A2(n14895), .ZN(n7723) );
  AND2_X1 U7780 ( .A1(n8189), .A2(n14857), .ZN(n7645) );
  OR2_X1 U7781 ( .A1(n15107), .A2(n14925), .ZN(n12523) );
  NAND2_X1 U7782 ( .A1(n7990), .A2(n7277), .ZN(n15011) );
  AOI21_X1 U7783 ( .B1(n15028), .B2(n15031), .A(n12506), .ZN(n15007) );
  NAND2_X1 U7784 ( .A1(n12233), .A2(n7638), .ZN(n7637) );
  NOR2_X1 U7785 ( .A1(n12234), .A2(n7639), .ZN(n7638) );
  INV_X1 U7786 ( .A(n12232), .ZN(n7639) );
  OR2_X1 U7787 ( .A1(n11649), .A2(n7236), .ZN(n7991) );
  NAND2_X1 U7788 ( .A1(n7855), .A2(n7854), .ZN(n11379) );
  XNOR2_X1 U7789 ( .A(n7365), .B(n15795), .ZN(n10787) );
  INV_X1 U7790 ( .A(n14747), .ZN(n7365) );
  INV_X1 U7791 ( .A(n15207), .ZN(n9757) );
  NAND2_X1 U7792 ( .A1(n9046), .A2(n9045), .ZN(n9079) );
  NAND2_X1 U7793 ( .A1(n9020), .A2(n9019), .ZN(n9042) );
  OAI21_X1 U7794 ( .B1(n11110), .B2(n7440), .A(n7439), .ZN(n11290) );
  NAND2_X1 U7795 ( .A1(n11285), .A2(n11108), .ZN(n7440) );
  NAND2_X1 U7796 ( .A1(n11113), .A2(n11285), .ZN(n7439) );
  OAI21_X1 U7797 ( .B1(n7299), .B2(n7422), .A(n8273), .ZN(n13050) );
  OAI21_X1 U7798 ( .B1(n12955), .B2(n12954), .A(n12952), .ZN(n7422) );
  INV_X1 U7799 ( .A(n14507), .ZN(n13057) );
  NAND2_X1 U7800 ( .A1(n12443), .A2(n12442), .ZN(n14341) );
  NAND2_X1 U7801 ( .A1(n14351), .A2(n14350), .ZN(n14352) );
  NAND2_X1 U7802 ( .A1(n14348), .A2(n15950), .ZN(n14351) );
  NAND2_X1 U7803 ( .A1(n9351), .A2(n9350), .ZN(n15145) );
  NOR2_X1 U7804 ( .A1(n15461), .A2(n15460), .ZN(n15459) );
  OR2_X1 U7805 ( .A1(n9040), .A2(n9038), .ZN(n7649) );
  AND2_X1 U7806 ( .A1(n7482), .A2(n12810), .ZN(n8204) );
  INV_X1 U7807 ( .A(n12808), .ZN(n7482) );
  NAND2_X1 U7808 ( .A1(n12808), .A2(n12811), .ZN(n8203) );
  NAND2_X1 U7809 ( .A1(n9112), .A2(n7626), .ZN(n7625) );
  OR2_X1 U7810 ( .A1(n8250), .A2(n9086), .ZN(n8249) );
  NAND2_X1 U7811 ( .A1(n9151), .A2(n9152), .ZN(n8241) );
  INV_X1 U7812 ( .A(n12867), .ZN(n7517) );
  INV_X1 U7813 ( .A(n12868), .ZN(n7518) );
  INV_X1 U7814 ( .A(n8208), .ZN(n7468) );
  AND2_X1 U7815 ( .A1(n8231), .A2(n9270), .ZN(n8230) );
  AOI21_X1 U7816 ( .B1(n7617), .B2(n7229), .A(n7615), .ZN(n7614) );
  AND2_X1 U7817 ( .A1(n7329), .A2(n7432), .ZN(n7454) );
  NAND2_X1 U7818 ( .A1(n7455), .A2(n7457), .ZN(n7432) );
  INV_X1 U7819 ( .A(n12894), .ZN(n7457) );
  NOR2_X1 U7820 ( .A1(n7455), .A2(n7458), .ZN(n7431) );
  NOR2_X1 U7821 ( .A1(n12894), .A2(n7273), .ZN(n7458) );
  OR2_X1 U7822 ( .A1(n9343), .A2(n9345), .ZN(n8244) );
  NAND2_X1 U7823 ( .A1(n9381), .A2(n7629), .ZN(n7628) );
  INV_X1 U7824 ( .A(n9380), .ZN(n7629) );
  AOI21_X1 U7825 ( .B1(n12915), .B2(n12914), .A(n12913), .ZN(n7423) );
  OAI21_X1 U7826 ( .B1(n12915), .B2(n12914), .A(n7301), .ZN(n7424) );
  NOR2_X1 U7827 ( .A1(n7473), .A2(n7474), .ZN(n7472) );
  NAND2_X1 U7828 ( .A1(n9431), .A2(n9428), .ZN(n8238) );
  NOR2_X1 U7829 ( .A1(n9431), .A2(n9428), .ZN(n8237) );
  OR2_X1 U7830 ( .A1(n13554), .A2(n13568), .ZN(n12705) );
  AND2_X1 U7831 ( .A1(n7785), .A2(n14885), .ZN(n7782) );
  NAND2_X1 U7832 ( .A1(n14861), .A2(n14841), .ZN(n7785) );
  INV_X1 U7833 ( .A(n7858), .ZN(n7857) );
  INV_X1 U7834 ( .A(n9330), .ZN(n8168) );
  NOR2_X1 U7835 ( .A1(n9257), .A2(n7419), .ZN(n7418) );
  INV_X1 U7836 ( .A(n9237), .ZN(n7419) );
  NAND2_X1 U7837 ( .A1(n15225), .A2(n7738), .ZN(n15227) );
  NAND2_X1 U7838 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n7739), .ZN(n7738) );
  INV_X1 U7839 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7739) );
  AND2_X1 U7840 ( .A1(n8152), .A2(n8146), .ZN(n8145) );
  NAND2_X1 U7841 ( .A1(n8151), .A2(n8148), .ZN(n8146) );
  AND2_X1 U7842 ( .A1(n12038), .A2(n12245), .ZN(n8152) );
  NAND2_X1 U7843 ( .A1(n8145), .A2(n8147), .ZN(n8143) );
  INV_X1 U7844 ( .A(n8148), .ZN(n8147) );
  OAI21_X1 U7845 ( .B1(n11454), .B2(P3_REG1_REG_2__SCAN_IN), .A(n7554), .ZN(
        n10296) );
  NAND2_X1 U7846 ( .A1(n11454), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7554) );
  NAND2_X1 U7847 ( .A1(n15664), .A2(n11466), .ZN(n11673) );
  OR2_X1 U7848 ( .A1(n13680), .A2(n13467), .ZN(n12607) );
  OR2_X1 U7849 ( .A1(n13181), .A2(n13508), .ZN(n7884) );
  NAND2_X1 U7850 ( .A1(n12583), .A2(n12684), .ZN(n7755) );
  INV_X1 U7851 ( .A(n12688), .ZN(n7752) );
  INV_X1 U7852 ( .A(n12684), .ZN(n7756) );
  INV_X1 U7853 ( .A(n12681), .ZN(n7388) );
  INV_X1 U7854 ( .A(n13637), .ZN(n7886) );
  AND2_X1 U7855 ( .A1(n7395), .A2(n8559), .ZN(n7889) );
  NOR2_X1 U7856 ( .A1(n7892), .A2(n8560), .ZN(n7891) );
  INV_X1 U7857 ( .A(n8541), .ZN(n7892) );
  NAND2_X1 U7858 ( .A1(n7749), .A2(n12634), .ZN(n7748) );
  INV_X1 U7859 ( .A(n12639), .ZN(n7747) );
  INV_X1 U7860 ( .A(n7584), .ZN(n7583) );
  OAI21_X1 U7861 ( .B1(n8366), .B2(n7585), .A(n8770), .ZN(n7584) );
  NAND2_X1 U7862 ( .A1(n8553), .A2(n8328), .ZN(n8329) );
  INV_X1 U7863 ( .A(n7575), .ZN(n7572) );
  INV_X1 U7864 ( .A(n7830), .ZN(n7569) );
  AOI21_X1 U7865 ( .B1(n7833), .B2(n7832), .A(n7831), .ZN(n7830) );
  INV_X1 U7866 ( .A(n8315), .ZN(n7832) );
  INV_X1 U7867 ( .A(n8318), .ZN(n7831) );
  INV_X1 U7868 ( .A(n8468), .ZN(n7835) );
  OR2_X1 U7869 ( .A1(n13985), .A2(n8017), .ZN(n8016) );
  NAND2_X1 U7870 ( .A1(n13832), .A2(n13833), .ZN(n8018) );
  OR2_X1 U7871 ( .A1(n14337), .A2(n14341), .ZN(n7843) );
  INV_X1 U7872 ( .A(n12479), .ZN(n8069) );
  NOR2_X1 U7873 ( .A1(n13009), .A2(n8052), .ZN(n8051) );
  NOR2_X1 U7874 ( .A1(n11606), .A2(n8053), .ZN(n8052) );
  INV_X1 U7875 ( .A(n11608), .ZN(n8053) );
  NOR2_X1 U7876 ( .A1(n11305), .A2(n7950), .ZN(n7949) );
  INV_X1 U7877 ( .A(n11301), .ZN(n7950) );
  NAND2_X1 U7878 ( .A1(n15903), .A2(n14016), .ZN(n11301) );
  NOR2_X1 U7879 ( .A1(n12836), .A2(n12828), .ZN(n7837) );
  OR2_X1 U7880 ( .A1(n10887), .A2(n10823), .ZN(n10825) );
  NAND2_X1 U7881 ( .A1(n13030), .A2(n10408), .ZN(n12766) );
  INV_X1 U7882 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9673) );
  INV_X1 U7883 ( .A(n14623), .ZN(n8123) );
  INV_X1 U7884 ( .A(n11209), .ZN(n14613) );
  NOR2_X1 U7885 ( .A1(n7256), .A2(n7246), .ZN(n7596) );
  NAND2_X1 U7886 ( .A1(n9517), .A2(n9519), .ZN(n8252) );
  INV_X1 U7887 ( .A(n7782), .ZN(n7780) );
  NOR2_X1 U7888 ( .A1(n9808), .A2(n8275), .ZN(n7854) );
  NAND2_X1 U7889 ( .A1(n7783), .A2(n7785), .ZN(n7781) );
  NAND2_X1 U7890 ( .A1(n14868), .A2(n7786), .ZN(n7783) );
  AOI21_X1 U7891 ( .B1(n7781), .B2(n7780), .A(n12525), .ZN(n7773) );
  INV_X1 U7892 ( .A(n12052), .ZN(n9825) );
  NAND2_X1 U7893 ( .A1(n9559), .A2(n9558), .ZN(n9563) );
  INV_X1 U7894 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8222) );
  INV_X1 U7895 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U7896 ( .A1(n9325), .A2(n9324), .ZN(n9329) );
  NAND2_X1 U7897 ( .A1(n9329), .A2(n7342), .ZN(n9346) );
  INV_X1 U7898 ( .A(n7699), .ZN(n7696) );
  NAND2_X1 U7899 ( .A1(n8187), .A2(n7788), .ZN(n7787) );
  INV_X1 U7900 ( .A(n9041), .ZN(n7788) );
  AOI21_X1 U7901 ( .B1(n8187), .B2(n8188), .A(n8186), .ZN(n8185) );
  INV_X1 U7902 ( .A(n9098), .ZN(n8186) );
  NAND2_X1 U7903 ( .A1(n8899), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7362) );
  XNOR2_X1 U7904 ( .A(n15227), .B(n7737), .ZN(n15265) );
  OR2_X1 U7905 ( .A1(n15262), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n15229) );
  AND2_X1 U7906 ( .A1(n13122), .A2(n8140), .ZN(n8139) );
  OR2_X1 U7907 ( .A1(n13220), .A2(n13105), .ZN(n8140) );
  NAND2_X1 U7908 ( .A1(n11575), .A2(n13256), .ZN(n8153) );
  AOI21_X1 U7909 ( .B1(n13182), .B2(n13246), .A(n8134), .ZN(n8133) );
  INV_X1 U7910 ( .A(n13183), .ZN(n8134) );
  NAND2_X1 U7911 ( .A1(n7258), .A2(n8149), .ZN(n8148) );
  INV_X1 U7912 ( .A(n12006), .ZN(n8149) );
  OR2_X1 U7913 ( .A1(n13202), .A2(n13509), .ZN(n13200) );
  NAND2_X1 U7914 ( .A1(n13219), .A2(n13220), .ZN(n13218) );
  OR2_X1 U7915 ( .A1(n12601), .A2(n12599), .ZN(n7764) );
  NAND2_X1 U7916 ( .A1(n7767), .A2(n7766), .ZN(n7765) );
  INV_X1 U7917 ( .A(n12597), .ZN(n7766) );
  INV_X1 U7918 ( .A(n12598), .ZN(n7767) );
  OAI21_X1 U7919 ( .B1(n12739), .B2(n12738), .A(n7827), .ZN(n7826) );
  AOI21_X1 U7920 ( .B1(n7829), .B2(n12738), .A(n7828), .ZN(n7827) );
  INV_X1 U7921 ( .A(n12740), .ZN(n7828) );
  INV_X1 U7922 ( .A(n12600), .ZN(n12743) );
  AND4_X1 U7923 ( .A1(n12556), .A2(n12555), .A3(n12554), .A4(n12553), .ZN(
        n13423) );
  AND4_X1 U7924 ( .A1(n8481), .A2(n8480), .A3(n8479), .A4(n8478), .ZN(n12009)
         );
  NAND2_X1 U7925 ( .A1(n7504), .A2(n7503), .ZN(n10291) );
  OR2_X1 U7926 ( .A1(n11454), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7504) );
  NAND2_X1 U7927 ( .A1(n11454), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7503) );
  OR2_X1 U7928 ( .A1(n7964), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n8436) );
  OR2_X1 U7929 ( .A1(n15529), .A2(n15528), .ZN(n7681) );
  XNOR2_X1 U7930 ( .A(n11462), .B(n15601), .ZN(n15604) );
  NOR2_X1 U7931 ( .A1(n15566), .A2(n7260), .ZN(n11397) );
  NAND2_X1 U7932 ( .A1(n15623), .A2(n15622), .ZN(n15621) );
  XNOR2_X1 U7933 ( .A(n11464), .B(n11438), .ZN(n15642) );
  NAND2_X1 U7934 ( .A1(n15642), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n15641) );
  OR2_X1 U7935 ( .A1(n15649), .A2(n15648), .ZN(n7959) );
  NAND2_X1 U7936 ( .A1(n15666), .A2(n15665), .ZN(n15664) );
  NAND2_X1 U7937 ( .A1(n7959), .A2(n7958), .ZN(n7957) );
  NAND2_X1 U7938 ( .A1(n15658), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7958) );
  NOR3_X1 U7939 ( .A1(n13302), .A2(n13301), .A3(n13304), .ZN(n13320) );
  AND2_X1 U7940 ( .A1(n13321), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7682) );
  NAND2_X1 U7941 ( .A1(n13341), .A2(n13342), .ZN(n13357) );
  AOI21_X1 U7942 ( .B1(n13385), .B2(n7952), .A(n7359), .ZN(n7951) );
  INV_X1 U7943 ( .A(n13385), .ZN(n7953) );
  AND2_X1 U7944 ( .A1(n12607), .A2(n12604), .ZN(n13454) );
  NAND2_X1 U7945 ( .A1(n8811), .A2(n12603), .ZN(n13448) );
  NAND2_X1 U7946 ( .A1(n7881), .A2(n7884), .ZN(n13479) );
  NAND2_X1 U7947 ( .A1(n7881), .A2(n7880), .ZN(n13480) );
  AND2_X1 U7948 ( .A1(n13481), .A2(n7884), .ZN(n7880) );
  AND2_X1 U7949 ( .A1(n12609), .A2(n8808), .ZN(n13493) );
  AND4_X1 U7950 ( .A1(n8743), .A2(n8742), .A3(n8741), .A4(n8740), .ZN(n13495)
         );
  INV_X1 U7951 ( .A(n13247), .ZN(n13548) );
  OAI21_X1 U7952 ( .B1(n13608), .B2(n7915), .A(n7912), .ZN(n13566) );
  AOI21_X1 U7953 ( .B1(n7914), .B2(n7913), .A(n7292), .ZN(n7912) );
  INV_X1 U7954 ( .A(n8638), .ZN(n7913) );
  OR2_X1 U7955 ( .A1(n13717), .A2(n13590), .ZN(n13561) );
  AND2_X1 U7956 ( .A1(n13561), .A2(n12693), .ZN(n13578) );
  NAND2_X1 U7957 ( .A1(n13608), .A2(n8638), .ZN(n13588) );
  AND2_X1 U7958 ( .A1(n12690), .A2(n12688), .ZN(n13611) );
  NAND2_X1 U7959 ( .A1(n8801), .A2(n12681), .ZN(n13621) );
  NAND2_X1 U7960 ( .A1(n13621), .A2(n13624), .ZN(n13620) );
  OAI21_X1 U7961 ( .B1(n12205), .B2(n7396), .A(n7394), .ZN(n7397) );
  AOI21_X1 U7962 ( .B1(n7757), .B2(n7761), .A(n7395), .ZN(n7394) );
  INV_X1 U7963 ( .A(n7757), .ZN(n7396) );
  NAND2_X1 U7964 ( .A1(n8542), .A2(n7891), .ZN(n7890) );
  AND2_X1 U7965 ( .A1(n12672), .A2(n12670), .ZN(n12581) );
  INV_X1 U7966 ( .A(n11674), .ZN(n11682) );
  NAND2_X1 U7967 ( .A1(n7909), .A2(n7908), .ZN(n11995) );
  NAND2_X1 U7968 ( .A1(n7897), .A2(n7895), .ZN(n11234) );
  NAND2_X1 U7969 ( .A1(n11193), .A2(n11192), .ZN(n7897) );
  AND4_X1 U7970 ( .A1(n8418), .A2(n8417), .A3(n8416), .A4(n8415), .ZN(n11238)
         );
  AND4_X1 U7971 ( .A1(n8447), .A2(n8446), .A3(n8445), .A4(n8444), .ZN(n11350)
         );
  NAND2_X1 U7972 ( .A1(n11240), .A2(n12632), .ZN(n11239) );
  NAND2_X1 U7973 ( .A1(n10624), .A2(n12727), .ZN(n15723) );
  OR2_X1 U7974 ( .A1(n10624), .A2(n12738), .ZN(n15721) );
  AND2_X1 U7975 ( .A1(n8786), .A2(n8862), .ZN(n15719) );
  NAND2_X1 U7976 ( .A1(n12551), .A2(n12550), .ZN(n13421) );
  NAND2_X1 U7977 ( .A1(n8737), .A2(n8736), .ZN(n13688) );
  OR2_X1 U7978 ( .A1(n7221), .A2(n11713), .ZN(n8736) );
  OR2_X1 U7979 ( .A1(n11329), .A2(n7219), .ZN(n8737) );
  NAND2_X1 U7980 ( .A1(n10751), .A2(n8850), .ZN(n15935) );
  INV_X1 U7981 ( .A(n10620), .ZN(n15697) );
  INV_X1 U7982 ( .A(n15723), .ZN(n13642) );
  NAND2_X1 U7983 ( .A1(n8829), .A2(n8828), .ZN(n10588) );
  NAND2_X1 U7984 ( .A1(n7811), .A2(n8364), .ZN(n8753) );
  XNOR2_X1 U7985 ( .A(n8817), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8833) );
  NOR2_X1 U7986 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(n7920), .ZN(n7917) );
  INV_X1 U7987 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8820) );
  INV_X1 U7988 ( .A(n7920), .ZN(n7918) );
  AOI21_X1 U7989 ( .B1(n8353), .B2(n7592), .A(n7591), .ZN(n7590) );
  INV_X1 U7990 ( .A(n8354), .ZN(n7591) );
  INV_X1 U7991 ( .A(n8349), .ZN(n7592) );
  NAND2_X1 U7992 ( .A1(n8688), .A2(n8348), .ZN(n8350) );
  NAND2_X1 U7993 ( .A1(n8345), .A2(n8346), .ZN(n8676) );
  OR2_X1 U7994 ( .A1(n8344), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8345) );
  AND2_X1 U7995 ( .A1(n8343), .A2(n8342), .ZN(n8656) );
  NAND2_X1 U7996 ( .A1(n7559), .A2(n7557), .ZN(n8626) );
  AOI21_X1 U7997 ( .B1(n7560), .B2(n7563), .A(n7558), .ZN(n7557) );
  INV_X1 U7998 ( .A(n8623), .ZN(n7558) );
  AND2_X1 U7999 ( .A1(n8335), .A2(n8334), .ZN(n8593) );
  AND2_X1 U8000 ( .A1(n8333), .A2(n8332), .ZN(n8576) );
  NAND2_X1 U8001 ( .A1(n8329), .A2(n10334), .ZN(n8331) );
  NAND2_X1 U8002 ( .A1(n7825), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8563) );
  INV_X1 U8003 ( .A(n8561), .ZN(n7825) );
  NAND2_X1 U8004 ( .A1(n8551), .A2(n8550), .ZN(n8553) );
  NOR2_X2 U8005 ( .A1(n8464), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8497) );
  NAND2_X1 U8006 ( .A1(n7573), .A2(n7575), .ZN(n8453) );
  NAND2_X1 U8007 ( .A1(n7574), .A2(n8434), .ZN(n7573) );
  INV_X1 U8008 ( .A(n8306), .ZN(n7821) );
  NAND2_X1 U8009 ( .A1(n8378), .A2(n8304), .ZN(n8395) );
  XNOR2_X1 U8010 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8303) );
  OAI22_X1 U8011 ( .A1(n10811), .A2(n11286), .B1(n12771), .B2(n7188), .ZN(
        n10493) );
  AND2_X1 U8012 ( .A1(n8028), .A2(n11960), .ZN(n8027) );
  NAND2_X1 U8013 ( .A1(n11290), .A2(n8030), .ZN(n8029) );
  NAND2_X1 U8014 ( .A1(n8030), .A2(n8031), .ZN(n8028) );
  NAND2_X1 U8015 ( .A1(n8021), .A2(n8020), .ZN(n13913) );
  AND2_X1 U8016 ( .A1(n13953), .A2(n7438), .ZN(n7435) );
  NAND2_X1 U8017 ( .A1(n7434), .A2(n7433), .ZN(n7437) );
  INV_X1 U8018 ( .A(n10452), .ZN(n7433) );
  INV_X1 U8019 ( .A(n10453), .ZN(n7434) );
  INV_X1 U8020 ( .A(n7445), .ZN(n7444) );
  INV_X1 U8021 ( .A(n13822), .ZN(n7446) );
  OAI21_X1 U8022 ( .B1(n13946), .B2(n7443), .A(n7302), .ZN(n13990) );
  INV_X1 U8023 ( .A(n13905), .ZN(n7443) );
  INV_X1 U8024 ( .A(n14169), .ZN(n14134) );
  NAND2_X1 U8025 ( .A1(n12214), .A2(n12215), .ZN(n12255) );
  NAND2_X1 U8026 ( .A1(n10408), .A2(n14078), .ZN(n13044) );
  NAND2_X1 U8027 ( .A1(n14027), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7477) );
  AND2_X1 U8028 ( .A1(n14115), .A2(n12432), .ZN(n14133) );
  NAND2_X1 U8029 ( .A1(n14177), .A2(n7240), .ZN(n14157) );
  INV_X1 U8030 ( .A(n7941), .ZN(n7940) );
  OAI21_X1 U8031 ( .B1(n13021), .B2(n7942), .A(n14154), .ZN(n7941) );
  NAND2_X1 U8032 ( .A1(n14175), .A2(n14174), .ZN(n14177) );
  AND2_X1 U8033 ( .A1(n12411), .A2(n12410), .ZN(n14188) );
  NAND2_X1 U8034 ( .A1(n7945), .A2(n7946), .ZN(n14187) );
  NOR2_X1 U8035 ( .A1(n12487), .A2(n8066), .ZN(n8065) );
  INV_X1 U8036 ( .A(n12485), .ZN(n8066) );
  AND2_X1 U8037 ( .A1(n12388), .A2(n12387), .ZN(n14223) );
  OR2_X1 U8038 ( .A1(n14221), .A2(n14220), .ZN(n14225) );
  NAND2_X1 U8039 ( .A1(n8056), .A2(n8059), .ZN(n14238) );
  AOI21_X1 U8040 ( .B1(n14258), .B2(n8060), .A(n7293), .ZN(n8059) );
  NAND2_X1 U8041 ( .A1(n12333), .A2(n12332), .ZN(n14259) );
  NOR2_X1 U8042 ( .A1(n13014), .A2(n7225), .ZN(n8071) );
  OR2_X1 U8043 ( .A1(n12058), .A2(n12074), .ZN(n12176) );
  OR2_X1 U8044 ( .A1(n12071), .A2(n12070), .ZN(n12073) );
  NAND2_X1 U8045 ( .A1(n11516), .A2(n11515), .ZN(n12857) );
  NAND2_X1 U8046 ( .A1(n8076), .A2(n7281), .ZN(n11519) );
  NOR2_X1 U8047 ( .A1(n13003), .A2(n7371), .ZN(n7370) );
  INV_X1 U8048 ( .A(n11009), .ZN(n7371) );
  AND2_X1 U8049 ( .A1(n10456), .A2(n10411), .ZN(n14242) );
  NAND2_X1 U8050 ( .A1(n10825), .A2(n8079), .ZN(n11017) );
  NOR2_X1 U8051 ( .A1(n12999), .A2(n8080), .ZN(n8079) );
  INV_X1 U8052 ( .A(n10824), .ZN(n8080) );
  NAND2_X1 U8053 ( .A1(n10818), .A2(n10817), .ZN(n10953) );
  INV_X1 U8054 ( .A(n12993), .ZN(n10956) );
  NAND2_X1 U8055 ( .A1(n12772), .A2(n12771), .ZN(n10811) );
  NOR2_X2 U8056 ( .A1(n7526), .A2(n13044), .ZN(n12761) );
  NAND2_X1 U8057 ( .A1(n12390), .A2(n12389), .ZN(n14193) );
  NAND2_X1 U8058 ( .A1(n12351), .A2(n12350), .ZN(n14396) );
  NAND2_X1 U8059 ( .A1(n11611), .A2(n11610), .ZN(n12865) );
  AND2_X1 U8060 ( .A1(n15778), .A2(n15807), .ZN(n15847) );
  AND2_X1 U8061 ( .A1(n14490), .A2(n10362), .ZN(n15335) );
  AOI21_X1 U8062 ( .B1(n8055), .B2(n7278), .A(n7373), .ZN(n10390) );
  NAND2_X1 U8063 ( .A1(n14474), .A2(n7374), .ZN(n7373) );
  NAND2_X1 U8064 ( .A1(n9690), .A2(n9688), .ZN(n9692) );
  NAND2_X1 U8065 ( .A1(n9686), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9695) );
  NAND2_X1 U8066 ( .A1(n7447), .A2(n7476), .ZN(n10377) );
  NOR2_X1 U8067 ( .A1(n7927), .A2(n9856), .ZN(n11040) );
  INV_X1 U8068 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n10278) );
  NOR2_X1 U8069 ( .A1(n8085), .A2(n8089), .ZN(n8084) );
  INV_X1 U8070 ( .A(n8087), .ZN(n8085) );
  NOR2_X1 U8071 ( .A1(n9751), .A2(n8090), .ZN(n8089) );
  INV_X1 U8072 ( .A(n16000), .ZN(n15050) );
  NAND2_X1 U8073 ( .A1(n11501), .A2(n11500), .ZN(n8098) );
  AND2_X1 U8074 ( .A1(n14658), .A2(n8122), .ZN(n8121) );
  OR2_X1 U8075 ( .A1(n14726), .A2(n8123), .ZN(n8122) );
  NAND2_X1 U8076 ( .A1(n8125), .A2(n9712), .ZN(n8126) );
  AOI21_X1 U8077 ( .B1(n10061), .B2(n14614), .A(n9711), .ZN(n8125) );
  NAND2_X1 U8078 ( .A1(n14750), .A2(n14615), .ZN(n9712) );
  AND2_X1 U8079 ( .A1(n9713), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9711) );
  OR2_X1 U8080 ( .A1(n14641), .A2(n8105), .ZN(n8104) );
  INV_X1 U8081 ( .A(n14597), .ZN(n8105) );
  AND2_X1 U8082 ( .A1(n9716), .A2(n9715), .ZN(n10043) );
  NAND2_X1 U8083 ( .A1(n11209), .A2(n14750), .ZN(n9716) );
  AND2_X1 U8084 ( .A1(n9713), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n9714) );
  AOI21_X1 U8085 ( .B1(n8109), .B2(n8112), .A(n7286), .ZN(n8107) );
  NAND2_X1 U8086 ( .A1(n11931), .A2(n8100), .ZN(n8099) );
  INV_X1 U8087 ( .A(n10800), .ZN(n8092) );
  NAND2_X1 U8088 ( .A1(n10603), .A2(n7491), .ZN(n7490) );
  INV_X1 U8089 ( .A(n9738), .ZN(n7491) );
  INV_X1 U8090 ( .A(n10945), .ZN(n8094) );
  NOR2_X1 U8091 ( .A1(n15200), .A2(n7600), .ZN(n7599) );
  INV_X1 U8092 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7600) );
  NAND2_X1 U8093 ( .A1(n8952), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8955) );
  AND2_X1 U8094 ( .A1(n11586), .A2(n7668), .ZN(n11589) );
  OR2_X1 U8095 ( .A1(n11588), .A2(n11587), .ZN(n7668) );
  NAND2_X1 U8096 ( .A1(n9598), .A2(n9597), .ZN(n14828) );
  NAND2_X1 U8097 ( .A1(n9573), .A2(n9572), .ZN(n14835) );
  NOR2_X1 U8098 ( .A1(n12525), .A2(n7780), .ZN(n7778) );
  OAI21_X1 U8099 ( .B1(n7781), .B2(n12525), .A(n12526), .ZN(n7776) );
  NAND2_X1 U8100 ( .A1(n7646), .A2(n7644), .ZN(n14843) );
  AND2_X1 U8101 ( .A1(n12525), .A2(n7303), .ZN(n7644) );
  AOI21_X1 U8102 ( .B1(n8191), .B2(n8193), .A(n7296), .ZN(n8189) );
  INV_X1 U8103 ( .A(n14874), .ZN(n14885) );
  AOI21_X1 U8104 ( .B1(n7998), .B2(n14913), .A(n7997), .ZN(n7996) );
  INV_X1 U8105 ( .A(n12524), .ZN(n7997) );
  OR2_X1 U8106 ( .A1(n15100), .A2(n14876), .ZN(n8266) );
  OR2_X1 U8107 ( .A1(n15108), .A2(n8193), .ZN(n14891) );
  NAND2_X1 U8108 ( .A1(n14905), .A2(n14904), .ZN(n14903) );
  OAI21_X1 U8109 ( .B1(n14969), .B2(n7633), .A(n7632), .ZN(n14938) );
  INV_X1 U8110 ( .A(n7634), .ZN(n7633) );
  AOI21_X1 U8111 ( .B1(n7634), .B2(n14957), .A(n7291), .ZN(n7632) );
  NAND2_X1 U8112 ( .A1(n7982), .A2(n7981), .ZN(n7800) );
  NAND2_X1 U8113 ( .A1(n7982), .A2(n7799), .ZN(n7798) );
  NOR2_X1 U8114 ( .A1(n14960), .A2(n14961), .ZN(n14959) );
  NAND2_X1 U8115 ( .A1(n15005), .A2(n7611), .ZN(n14991) );
  NOR2_X1 U8116 ( .A1(n14997), .A2(n7612), .ZN(n7611) );
  INV_X1 U8117 ( .A(n12507), .ZN(n7612) );
  NAND2_X1 U8118 ( .A1(n14991), .A2(n7866), .ZN(n14981) );
  NOR2_X1 U8119 ( .A1(n14984), .A2(n7867), .ZN(n7866) );
  INV_X1 U8120 ( .A(n12508), .ZN(n7867) );
  OR2_X1 U8121 ( .A1(n15145), .A2(n15008), .ZN(n12519) );
  NAND2_X1 U8122 ( .A1(n14996), .A2(n7984), .ZN(n14973) );
  NAND2_X1 U8123 ( .A1(n15011), .A2(n8270), .ZN(n14998) );
  NOR2_X1 U8124 ( .A1(n15031), .A2(n7988), .ZN(n7987) );
  INV_X1 U8125 ( .A(n12518), .ZN(n7988) );
  OAI22_X1 U8126 ( .A1(n12517), .A2(n12236), .B1(n15989), .B2(n16000), .ZN(
        n15047) );
  NAND2_X1 U8127 ( .A1(n12283), .A2(n8265), .ZN(n12517) );
  OR2_X1 U8128 ( .A1(n14521), .A2(n14520), .ZN(n8265) );
  NOR2_X1 U8129 ( .A1(n12020), .A2(n7993), .ZN(n7992) );
  INV_X1 U8130 ( .A(n11644), .ZN(n7993) );
  AOI21_X1 U8131 ( .B1(n11556), .B2(n11555), .A(n8263), .ZN(n11558) );
  NAND2_X1 U8132 ( .A1(n7995), .A2(n7994), .ZN(n11645) );
  INV_X1 U8133 ( .A(n11558), .ZN(n7995) );
  OAI21_X1 U8134 ( .B1(n11160), .B2(n7305), .A(n7851), .ZN(n7613) );
  AND2_X1 U8135 ( .A1(n11152), .A2(n7722), .ZN(n11478) );
  NOR2_X1 U8136 ( .A1(n11486), .A2(n11377), .ZN(n7722) );
  INV_X1 U8137 ( .A(n11160), .ZN(n9823) );
  AND2_X1 U8138 ( .A1(n7308), .A2(n9799), .ZN(n7977) );
  NAND2_X1 U8139 ( .A1(n8985), .A2(n7979), .ZN(n10658) );
  OR2_X1 U8140 ( .A1(n9891), .A2(n8984), .ZN(n8985) );
  INV_X1 U8141 ( .A(n7980), .ZN(n7979) );
  OAI22_X1 U8142 ( .A1(n9104), .A2(n9849), .B1(n9870), .B2(n9209), .ZN(n7980)
         );
  NAND2_X1 U8143 ( .A1(n7643), .A2(n8988), .ZN(n10700) );
  INV_X1 U8144 ( .A(n9812), .ZN(n7643) );
  INV_X1 U8145 ( .A(n15049), .ZN(n15033) );
  AND2_X1 U8146 ( .A1(n14914), .A2(n14913), .ZN(n15108) );
  INV_X1 U8147 ( .A(n16016), .ZN(n15985) );
  NAND2_X1 U8148 ( .A1(n11151), .A2(n9807), .ZN(n9809) );
  OR2_X1 U8149 ( .A1(n9209), .A2(n10397), .ZN(n8949) );
  NOR2_X1 U8150 ( .A1(n9756), .A2(n15203), .ZN(n9872) );
  OR2_X1 U8151 ( .A1(n9569), .A2(n9568), .ZN(n9591) );
  INV_X1 U8152 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7641) );
  AND3_X1 U8153 ( .A1(n9105), .A2(n7231), .A3(n7719), .ZN(n9661) );
  OAI21_X1 U8154 ( .B1(n9376), .B2(n7249), .A(n7345), .ZN(n8174) );
  XNOR2_X1 U8155 ( .A(n9442), .B(n9443), .ZN(n12374) );
  INV_X1 U8156 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8921) );
  NAND2_X1 U8157 ( .A1(n8176), .A2(n9388), .ZN(n9396) );
  NAND2_X1 U8158 ( .A1(n8183), .A2(n8180), .ZN(n8176) );
  NAND2_X1 U8159 ( .A1(n9202), .A2(n7805), .ZN(n9238) );
  NOR2_X1 U8160 ( .A1(n9206), .A2(n7806), .ZN(n7805) );
  INV_X1 U8161 ( .A(n9201), .ZN(n7806) );
  NAND2_X1 U8162 ( .A1(n7425), .A2(n7690), .ZN(n9134) );
  INV_X1 U8163 ( .A(n9124), .ZN(n7690) );
  AND2_X1 U8164 ( .A1(n9130), .A2(n9166), .ZN(n10069) );
  NAND2_X1 U8165 ( .A1(n9079), .A2(n9078), .ZN(n9097) );
  NAND2_X1 U8166 ( .A1(n9042), .A2(n9041), .ZN(n9046) );
  INV_X1 U8167 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7672) );
  NAND2_X1 U8168 ( .A1(n8979), .A2(n8978), .ZN(n9001) );
  OAI21_X1 U8169 ( .B1(n15444), .B2(n15445), .A(n7741), .ZN(n7740) );
  XNOR2_X1 U8170 ( .A(n15263), .B(n7265), .ZN(n15264) );
  NAND2_X1 U8171 ( .A1(n15502), .A2(n15504), .ZN(n15290) );
  OAI21_X1 U8172 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n15237), .A(n15236), .ZN(
        n15298) );
  AOI21_X1 U8173 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n15241), .A(n15240), .ZN(
        n15301) );
  NAND2_X1 U8174 ( .A1(n8713), .A2(n8712), .ZN(n13514) );
  OR2_X1 U8175 ( .A1(n7221), .A2(n11723), .ZN(n8712) );
  NAND2_X1 U8176 ( .A1(n10775), .A2(n7483), .ZN(n10872) );
  AND2_X1 U8177 ( .A1(n10776), .A2(n10774), .ZN(n7483) );
  NAND2_X1 U8178 ( .A1(n8373), .A2(n8372), .ZN(n13116) );
  NAND2_X1 U8179 ( .A1(n8690), .A2(n8689), .ZN(n13539) );
  OR2_X1 U8180 ( .A1(n7221), .A2(n10749), .ZN(n8689) );
  AND4_X1 U8181 ( .A1(n8528), .A2(n8527), .A3(n8526), .A4(n8525), .ZN(n12164)
         );
  NOR2_X1 U8182 ( .A1(n13076), .A2(n7275), .ZN(n8161) );
  INV_X1 U8183 ( .A(n13664), .ZN(n13742) );
  NAND2_X1 U8184 ( .A1(n8702), .A2(n8701), .ZN(n13525) );
  INV_X1 U8185 ( .A(n13249), .ZN(n13580) );
  NAND2_X1 U8186 ( .A1(n10356), .A2(n15727), .ZN(n13206) );
  AND4_X1 U8187 ( .A1(n8590), .A2(n8589), .A3(n8588), .A4(n8587), .ZN(n13656)
         );
  AND4_X1 U8188 ( .A1(n12556), .A2(n8778), .A3(n8777), .A4(n8776), .ZN(n13439)
         );
  AND4_X1 U8189 ( .A1(n8301), .A2(n8300), .A3(n8299), .A4(n8298), .ZN(n13456)
         );
  INV_X1 U8190 ( .A(n12306), .ZN(n13644) );
  INV_X1 U8191 ( .A(n12164), .ZN(n13253) );
  XNOR2_X1 U8192 ( .A(n7957), .B(n11674), .ZN(n11403) );
  NOR2_X1 U8193 ( .A1(n11404), .A2(n11403), .ZN(n11668) );
  NAND2_X1 U8194 ( .A1(n11451), .A2(n11450), .ZN(n11687) );
  AND2_X1 U8195 ( .A1(P3_U3897), .A2(n8787), .ZN(n13412) );
  XNOR2_X1 U8196 ( .A(n13403), .B(n13409), .ZN(n7402) );
  AOI211_X1 U8197 ( .C1(n13419), .C2(n15602), .A(n7348), .B(n7972), .ZN(n7971)
         );
  INV_X1 U8198 ( .A(n13418), .ZN(n7972) );
  NAND2_X1 U8199 ( .A1(n8667), .A2(n8666), .ZN(n13713) );
  NAND2_X1 U8200 ( .A1(n8601), .A2(n8600), .ZN(n13789) );
  NAND2_X1 U8201 ( .A1(n8584), .A2(n8583), .ZN(n13793) );
  XNOR2_X1 U8202 ( .A(n8663), .B(n8662), .ZN(n13407) );
  INV_X1 U8203 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8662) );
  NOR2_X1 U8204 ( .A1(n8005), .A2(n10555), .ZN(n8004) );
  NAND2_X1 U8205 ( .A1(n10520), .A2(n14510), .ZN(n7533) );
  NAND2_X1 U8206 ( .A1(n12380), .A2(n12379), .ZN(n14386) );
  OR2_X1 U8207 ( .A1(n14505), .A2(n10521), .ZN(n12380) );
  OR2_X1 U8208 ( .A1(n12960), .A2(n10446), .ZN(n7500) );
  INV_X1 U8209 ( .A(n8206), .ZN(n8205) );
  OAI21_X1 U8210 ( .B1(n13048), .B2(n13049), .A(n13052), .ZN(n8206) );
  INV_X1 U8211 ( .A(n13036), .ZN(n13049) );
  INV_X1 U8212 ( .A(n13050), .ZN(n7421) );
  INV_X1 U8213 ( .A(n14223), .ZN(n14007) );
  AND2_X1 U8214 ( .A1(n10187), .A2(n14487), .ZN(n15419) );
  OR2_X1 U8215 ( .A1(n10181), .A2(n14487), .ZN(n15406) );
  AOI22_X1 U8216 ( .A1(n14095), .A2(n14097), .B1(n14341), .B2(n14114), .ZN(
        n12494) );
  INV_X1 U8217 ( .A(n7928), .ZN(n14339) );
  AOI21_X1 U8218 ( .B1(n7933), .B2(n14309), .A(n12474), .ZN(n7931) );
  INV_X1 U8219 ( .A(n7494), .ZN(n7368) );
  INV_X1 U8220 ( .A(n7522), .ZN(n7521) );
  OAI21_X1 U8221 ( .B1(n14347), .B2(n15778), .A(n14118), .ZN(n7522) );
  NAND2_X1 U8222 ( .A1(n14255), .A2(n14258), .ZN(n14256) );
  NAND2_X1 U8223 ( .A1(n14281), .A2(n12483), .ZN(n14255) );
  INV_X1 U8224 ( .A(n15829), .ZN(n14275) );
  INV_X1 U8225 ( .A(n14234), .ZN(n15823) );
  NAND2_X1 U8226 ( .A1(n15340), .A2(n10477), .ZN(n14318) );
  NAND2_X1 U8227 ( .A1(n10520), .A2(n7849), .ZN(n7848) );
  OAI22_X1 U8228 ( .A1(n10397), .A2(n10395), .B1(n10396), .B2(n10404), .ZN(
        n7849) );
  NAND2_X1 U8229 ( .A1(n14275), .A2(n14073), .ZN(n14234) );
  NAND2_X1 U8230 ( .A1(n12948), .A2(n12947), .ZN(n14330) );
  INV_X1 U8231 ( .A(n14441), .ZN(n14363) );
  NAND2_X1 U8232 ( .A1(n10567), .A2(n10566), .ZN(n15819) );
  NAND2_X1 U8233 ( .A1(n7494), .A2(n7493), .ZN(n14433) );
  INV_X1 U8234 ( .A(n14346), .ZN(n7493) );
  AND2_X1 U8235 ( .A1(n12434), .A2(n12433), .ZN(n14437) );
  AND2_X1 U8236 ( .A1(n10470), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15340) );
  OR3_X1 U8237 ( .A1(n10157), .A2(n9685), .A3(n11039), .ZN(n10162) );
  NOR2_X1 U8238 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n10159) );
  NAND2_X1 U8239 ( .A1(n9516), .A2(n9515), .ZN(n15087) );
  NAND2_X1 U8240 ( .A1(n9244), .A2(n9243), .ZN(n15165) );
  NAND2_X1 U8241 ( .A1(n8098), .A2(n8097), .ZN(n11932) );
  AND2_X1 U8242 ( .A1(n11506), .A2(n7349), .ZN(n8097) );
  NAND2_X1 U8243 ( .A1(n9537), .A2(n9536), .ZN(n15081) );
  INV_X1 U8244 ( .A(n12127), .ZN(n15170) );
  NAND2_X1 U8245 ( .A1(n7361), .A2(n9595), .ZN(n9026) );
  INV_X1 U8246 ( .A(n10549), .ZN(n7361) );
  NAND2_X1 U8247 ( .A1(n9451), .A2(n9450), .ZN(n15107) );
  OR2_X1 U8248 ( .A1(n12264), .A2(n12263), .ZN(n8256) );
  NAND2_X1 U8249 ( .A1(n9171), .A2(n9170), .ZN(n15917) );
  AOI21_X1 U8250 ( .B1(n9609), .B2(n9608), .A(n9607), .ZN(n9610) );
  NAND4_X1 U8251 ( .A1(n8970), .A2(n8969), .A3(n8968), .A4(n8967), .ZN(n14749)
         );
  OR2_X1 U8252 ( .A1(n9546), .A2(n8938), .ZN(n8940) );
  OAI21_X1 U8253 ( .B1(n9333), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U8254 ( .A1(n9427), .A2(n9426), .ZN(n15117) );
  NAND2_X1 U8255 ( .A1(n15218), .A2(n9891), .ZN(n14954) );
  NAND2_X1 U8256 ( .A1(n9315), .A2(n9314), .ZN(n16027) );
  OR2_X1 U8257 ( .A1(n15204), .A2(n9760), .ZN(n15193) );
  CLKBUF_X1 U8258 ( .A(n9705), .Z(n15217) );
  XNOR2_X1 U8259 ( .A(n15270), .B(n7505), .ZN(n15509) );
  NOR2_X1 U8260 ( .A1(n15509), .A2(n15508), .ZN(n15507) );
  NAND2_X1 U8261 ( .A1(n15463), .A2(n15464), .ZN(n15462) );
  XNOR2_X1 U8262 ( .A(n7744), .B(n15305), .ZN(n15478) );
  NAND2_X1 U8263 ( .A1(n15478), .A2(n15477), .ZN(n15476) );
  NOR2_X1 U8264 ( .A1(n15498), .A2(n15497), .ZN(n15496) );
  INV_X1 U8265 ( .A(n12770), .ZN(n7481) );
  OR2_X1 U8266 ( .A1(n12781), .A2(n12768), .ZN(n7507) );
  NAND2_X1 U8267 ( .A1(n12782), .A2(n12783), .ZN(n12786) );
  NAND2_X1 U8268 ( .A1(n8987), .A2(n8986), .ZN(n9009) );
  NAND2_X1 U8269 ( .A1(n9267), .A2(n14749), .ZN(n8987) );
  NAND2_X1 U8270 ( .A1(n9606), .A2(n10658), .ZN(n8986) );
  AND2_X1 U8271 ( .A1(n9623), .A2(n9267), .ZN(n8965) );
  OR2_X1 U8272 ( .A1(n9009), .A2(n9798), .ZN(n8992) );
  MUX2_X1 U8273 ( .A(n9814), .B(n9623), .S(n9606), .Z(n8990) );
  OAI21_X1 U8274 ( .B1(n7288), .B2(n7648), .A(n7647), .ZN(n9064) );
  OR2_X1 U8275 ( .A1(n7650), .A2(n9039), .ZN(n7647) );
  NAND2_X1 U8276 ( .A1(n9014), .A2(n7649), .ZN(n7648) );
  NAND2_X1 U8277 ( .A1(n7464), .A2(n12819), .ZN(n12825) );
  OAI21_X1 U8278 ( .B1(n12809), .B2(n8204), .A(n7547), .ZN(n12819) );
  AND2_X1 U8279 ( .A1(n12818), .A2(n8203), .ZN(n7547) );
  INV_X1 U8280 ( .A(n12831), .ZN(n8212) );
  INV_X1 U8281 ( .A(n9085), .ZN(n8250) );
  INV_X1 U8282 ( .A(n12838), .ZN(n7519) );
  INV_X1 U8283 ( .A(n12839), .ZN(n7520) );
  INV_X1 U8284 ( .A(n9155), .ZN(n7603) );
  AND2_X1 U8285 ( .A1(n8241), .A2(n7624), .ZN(n7623) );
  NAND2_X1 U8286 ( .A1(n9111), .A2(n9113), .ZN(n7624) );
  AOI21_X1 U8287 ( .B1(n8243), .B2(n8242), .A(n11553), .ZN(n8239) );
  INV_X1 U8288 ( .A(n9152), .ZN(n8242) );
  INV_X1 U8289 ( .A(n9151), .ZN(n8243) );
  NAND2_X1 U8290 ( .A1(n9224), .A2(n9227), .ZN(n7620) );
  NOR2_X1 U8291 ( .A1(n9248), .A2(n9245), .ZN(n8233) );
  NAND2_X1 U8292 ( .A1(n9245), .A2(n9248), .ZN(n8232) );
  NAND2_X1 U8293 ( .A1(n9196), .A2(n8227), .ZN(n8226) );
  NAND2_X1 U8294 ( .A1(n7460), .A2(n7283), .ZN(n12868) );
  INV_X1 U8295 ( .A(n12860), .ZN(n8213) );
  NAND2_X1 U8296 ( .A1(n8233), .A2(n8232), .ZN(n8231) );
  INV_X1 U8297 ( .A(n9224), .ZN(n7621) );
  NOR2_X1 U8298 ( .A1(n8233), .A2(n7618), .ZN(n7617) );
  INV_X1 U8299 ( .A(n7620), .ZN(n7618) );
  INV_X1 U8300 ( .A(n8232), .ZN(n7615) );
  NOR2_X1 U8301 ( .A1(n7289), .A2(n7467), .ZN(n7466) );
  NAND2_X1 U8302 ( .A1(n9294), .A2(n9296), .ZN(n8224) );
  NAND2_X1 U8303 ( .A1(n7454), .A2(n7431), .ZN(n7450) );
  NAND2_X1 U8304 ( .A1(n8246), .A2(n8245), .ZN(n9364) );
  OR2_X1 U8305 ( .A1(n8247), .A2(n9344), .ZN(n8245) );
  INV_X1 U8306 ( .A(n9343), .ZN(n8247) );
  NAND2_X1 U8307 ( .A1(n7631), .A2(n9380), .ZN(n7630) );
  INV_X1 U8308 ( .A(n10787), .ZN(n9818) );
  INV_X1 U8309 ( .A(n8710), .ZN(n7589) );
  NOR2_X1 U8310 ( .A1(n7290), .A2(n7472), .ZN(n7471) );
  NOR2_X1 U8311 ( .A1(n7424), .A2(n7423), .ZN(n7470) );
  NOR2_X1 U8312 ( .A1(n8237), .A2(n8235), .ZN(n8234) );
  NOR2_X1 U8313 ( .A1(n7224), .A2(n7861), .ZN(n7860) );
  INV_X1 U8314 ( .A(n9815), .ZN(n7861) );
  NAND2_X1 U8315 ( .A1(n13454), .A2(n12573), .ZN(n12611) );
  OAI21_X1 U8316 ( .B1(n12611), .B2(n7771), .A(n7813), .ZN(n7812) );
  NOR2_X1 U8317 ( .A1(n7814), .A2(n12727), .ZN(n7813) );
  INV_X1 U8318 ( .A(n12610), .ZN(n7814) );
  INV_X1 U8319 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n11892) );
  INV_X1 U8320 ( .A(n12666), .ZN(n7762) );
  INV_X1 U8321 ( .A(n8341), .ZN(n7566) );
  INV_X1 U8322 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9683) );
  NAND2_X1 U8323 ( .A1(n7312), .A2(n7244), .ZN(n7597) );
  NAND2_X1 U8324 ( .A1(n9477), .A2(n8255), .ZN(n8254) );
  NAND2_X1 U8325 ( .A1(n14959), .A2(n14954), .ZN(n14932) );
  NOR2_X1 U8326 ( .A1(n9817), .A2(n7864), .ZN(n7863) );
  INV_X1 U8327 ( .A(n9816), .ZN(n7864) );
  INV_X1 U8328 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8877) );
  INV_X1 U8329 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8917) );
  INV_X1 U8330 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9210) );
  INV_X1 U8331 ( .A(n9190), .ZN(n7804) );
  NOR2_X1 U8332 ( .A1(n9101), .A2(n7700), .ZN(n7699) );
  NOR2_X1 U8333 ( .A1(n7699), .A2(n9018), .ZN(n7694) );
  NAND2_X1 U8334 ( .A1(n9288), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7509) );
  OAI21_X1 U8335 ( .B1(n9288), .B2(n9852), .A(n7501), .ZN(n9002) );
  NAND2_X1 U8336 ( .A1(n9288), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7501) );
  OAI21_X1 U8337 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n15250), .A(n15249), .ZN(
        n15251) );
  NOR2_X1 U8338 ( .A1(n8668), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8669) );
  BUF_X1 U8339 ( .A(n13106), .Z(n7543) );
  NAND2_X1 U8340 ( .A1(n12737), .A2(n12736), .ZN(n7829) );
  INV_X1 U8341 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7391) );
  NAND2_X1 U8342 ( .A1(n13268), .A2(n7350), .ZN(n13292) );
  INV_X1 U8343 ( .A(n13333), .ZN(n7970) );
  OR2_X1 U8344 ( .A1(n13514), .A2(n13522), .ZN(n12717) );
  OR2_X1 U8345 ( .A1(n13539), .A2(n13548), .ZN(n12709) );
  INV_X1 U8346 ( .A(n7906), .ZN(n7899) );
  INV_X1 U8347 ( .A(n7902), .ZN(n7901) );
  OAI21_X1 U8348 ( .B1(n7908), .B2(n7903), .A(n12163), .ZN(n7902) );
  NAND2_X1 U8349 ( .A1(n15697), .A2(n13262), .ZN(n12618) );
  NAND2_X1 U8350 ( .A1(n15712), .A2(n12614), .ZN(n11055) );
  INV_X1 U8351 ( .A(n13264), .ZN(n11173) );
  INV_X1 U8352 ( .A(n8367), .ZN(n7585) );
  AND2_X1 U8353 ( .A1(n7588), .A2(n8355), .ZN(n7587) );
  NAND2_X1 U8354 ( .A1(n7922), .A2(n7921), .ZN(n7920) );
  INV_X1 U8355 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7922) );
  INV_X1 U8356 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7921) );
  INV_X1 U8357 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9289) );
  OAI21_X1 U8358 ( .B1(n8394), .B2(n7821), .A(n8405), .ZN(n7816) );
  NOR2_X1 U8359 ( .A1(n7819), .A2(n7821), .ZN(n7818) );
  INV_X1 U8360 ( .A(n8304), .ZN(n7819) );
  XNOR2_X1 U8361 ( .A(n10440), .B(n10445), .ZN(n10442) );
  INV_X1 U8362 ( .A(n13993), .ZN(n8043) );
  NAND2_X1 U8363 ( .A1(n13905), .A2(n7442), .ZN(n7441) );
  INV_X1 U8364 ( .A(n13855), .ZN(n7442) );
  NAND2_X1 U8365 ( .A1(n8199), .A2(n12938), .ZN(n8198) );
  NAND2_X1 U8366 ( .A1(n7251), .A2(n7227), .ZN(n8199) );
  INV_X1 U8367 ( .A(n12766), .ZN(n12981) );
  INV_X1 U8368 ( .A(n12493), .ZN(n8073) );
  INV_X1 U8369 ( .A(n8065), .ZN(n8064) );
  AOI21_X1 U8370 ( .B1(n7226), .B2(n14220), .A(n7309), .ZN(n7946) );
  NOR2_X1 U8371 ( .A1(n13016), .A2(n8058), .ZN(n8057) );
  INV_X1 U8372 ( .A(n14288), .ZN(n8058) );
  INV_X1 U8373 ( .A(n12483), .ZN(n8060) );
  NOR2_X1 U8374 ( .A1(n12873), .A2(n7704), .ZN(n7703) );
  INV_X1 U8375 ( .A(n11978), .ZN(n7704) );
  NAND2_X1 U8376 ( .A1(n11302), .A2(n7949), .ZN(n11529) );
  OR2_X1 U8377 ( .A1(n10922), .A2(n10921), .ZN(n11079) );
  AND2_X1 U8378 ( .A1(n10820), .A2(n10817), .ZN(n8044) );
  NAND2_X1 U8379 ( .A1(n12993), .A2(n10820), .ZN(n8047) );
  NAND2_X1 U8380 ( .A1(n10812), .A2(n12776), .ZN(n10828) );
  NAND2_X1 U8381 ( .A1(n7375), .A2(n11039), .ZN(n7374) );
  INV_X1 U8382 ( .A(n9677), .ZN(n7380) );
  INV_X1 U8383 ( .A(n14583), .ZN(n9735) );
  AND2_X1 U8384 ( .A1(n14647), .A2(n8110), .ZN(n8109) );
  NAND2_X1 U8385 ( .A1(n8111), .A2(n14554), .ZN(n8110) );
  INV_X1 U8386 ( .A(n14717), .ZN(n8111) );
  INV_X1 U8387 ( .A(n14554), .ZN(n8112) );
  NOR2_X1 U8388 ( .A1(n9731), .A2(n9730), .ZN(n9738) );
  OR2_X1 U8389 ( .A1(n9546), .A2(n8889), .ZN(n8890) );
  NAND2_X1 U8390 ( .A1(n14861), .A2(n14884), .ZN(n7724) );
  INV_X1 U8391 ( .A(n14894), .ZN(n7725) );
  INV_X1 U8392 ( .A(n9401), .ZN(n9402) );
  INV_X1 U8393 ( .A(n7984), .ZN(n7981) );
  NOR2_X1 U8394 ( .A1(n14968), .A2(n7983), .ZN(n7982) );
  INV_X1 U8395 ( .A(n8264), .ZN(n7983) );
  AND2_X1 U8396 ( .A1(n14942), .A2(n12510), .ZN(n7634) );
  NOR2_X1 U8397 ( .A1(n15017), .A2(n15145), .ZN(n7726) );
  AND2_X1 U8398 ( .A1(n9179), .A2(n9178), .ZN(n9215) );
  INV_X1 U8399 ( .A(n11378), .ZN(n7853) );
  INV_X1 U8400 ( .A(n8276), .ZN(n7850) );
  INV_X1 U8401 ( .A(n7364), .ZN(n7975) );
  AND2_X1 U8402 ( .A1(n9027), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9052) );
  OR2_X1 U8403 ( .A1(n14933), .A2(n15107), .ZN(n14906) );
  OR2_X1 U8404 ( .A1(n15117), .A2(n14932), .ZN(n14933) );
  NOR2_X1 U8405 ( .A1(n15057), .A2(n16027), .ZN(n15014) );
  NOR2_X1 U8406 ( .A1(n12269), .A2(n15165), .ZN(n7716) );
  NAND2_X1 U8407 ( .A1(n11379), .A2(n11378), .ZN(n11484) );
  INV_X1 U8408 ( .A(n7862), .ZN(n10788) );
  AOI21_X1 U8409 ( .B1(n7865), .B2(n7863), .A(n7224), .ZN(n7862) );
  NAND2_X1 U8410 ( .A1(n9449), .A2(n9448), .ZN(n9491) );
  INV_X1 U8411 ( .A(n9398), .ZN(n8175) );
  NOR2_X1 U8412 ( .A1(n9389), .A2(n8182), .ZN(n8180) );
  NAND2_X1 U8413 ( .A1(n7417), .A2(n9261), .ZN(n9284) );
  NAND2_X1 U8414 ( .A1(n9238), .A2(n7418), .ZN(n7417) );
  OAI21_X1 U8415 ( .B1(n8973), .B2(n8903), .A(SI_2_), .ZN(n8974) );
  INV_X1 U8416 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n15262) );
  NAND2_X1 U8417 ( .A1(n7404), .A2(n15228), .ZN(n15263) );
  NAND2_X1 U8418 ( .A1(n15265), .A2(n15266), .ZN(n7404) );
  INV_X1 U8419 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15278) );
  INV_X1 U8420 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n15284) );
  AND2_X1 U8421 ( .A1(n13103), .A2(n13101), .ZN(n13156) );
  NAND2_X1 U8422 ( .A1(n7545), .A2(n7544), .ZN(n13172) );
  INV_X1 U8423 ( .A(n13175), .ZN(n7544) );
  AND2_X1 U8424 ( .A1(n13155), .A2(n13098), .ZN(n13183) );
  INV_X1 U8425 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11787) );
  AND2_X1 U8426 ( .A1(n8143), .A2(n12042), .ZN(n8142) );
  INV_X1 U8427 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n11915) );
  INV_X1 U8428 ( .A(SI_22_), .ZN(n9443) );
  OR3_X1 U8429 ( .A1(n8522), .A2(P3_REG3_REG_10__SCAN_IN), .A3(
        P3_REG3_REG_11__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U8430 ( .A1(n13172), .A2(n8165), .ZN(n13210) );
  NOR2_X1 U8431 ( .A1(n11046), .A2(n8269), .ZN(n8158) );
  INV_X1 U8432 ( .A(n8159), .ZN(n8156) );
  NAND2_X1 U8433 ( .A1(n10289), .A2(n10288), .ZN(n10290) );
  NAND2_X1 U8434 ( .A1(n10290), .A2(n10291), .ZN(n11393) );
  NAND2_X1 U8435 ( .A1(n10297), .A2(n10296), .ZN(n11453) );
  NAND2_X1 U8436 ( .A1(n11393), .A2(n7673), .ZN(n11394) );
  NAND2_X1 U8437 ( .A1(n7674), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7673) );
  NAND2_X1 U8438 ( .A1(n11414), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7680) );
  OAI21_X1 U8439 ( .B1(n15604), .B2(n15603), .A(n7556), .ZN(n15623) );
  NAND2_X1 U8440 ( .A1(n11398), .A2(n11461), .ZN(n7955) );
  OR2_X1 U8441 ( .A1(n15589), .A2(n15590), .ZN(n7956) );
  NAND2_X1 U8442 ( .A1(n11436), .A2(n15613), .ZN(n15635) );
  NOR2_X1 U8443 ( .A1(n15609), .A2(n7954), .ZN(n11400) );
  NOR2_X1 U8444 ( .A1(n11463), .A2(n11399), .ZN(n7954) );
  NAND2_X1 U8445 ( .A1(n15641), .A2(n11465), .ZN(n15666) );
  NAND2_X1 U8446 ( .A1(n11675), .A2(n11676), .ZN(n11679) );
  NAND2_X1 U8447 ( .A1(n11679), .A2(n11678), .ZN(n13268) );
  NOR2_X1 U8448 ( .A1(n13265), .A2(n7683), .ZN(n13286) );
  NOR2_X1 U8449 ( .A1(n13269), .A2(n11670), .ZN(n7683) );
  XNOR2_X1 U8450 ( .A(n13292), .B(n13287), .ZN(n13270) );
  XNOR2_X1 U8451 ( .A(n13339), .B(n13337), .ZN(n13315) );
  NAND2_X1 U8452 ( .A1(n13315), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n13341) );
  OR2_X1 U8453 ( .A1(n13311), .A2(n7967), .ZN(n7965) );
  NAND2_X1 U8454 ( .A1(n7970), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7967) );
  NAND2_X1 U8455 ( .A1(n13330), .A2(n7970), .ZN(n7966) );
  OAI21_X1 U8456 ( .B1(n13370), .B2(n7515), .A(n7514), .ZN(n13374) );
  NOR2_X1 U8457 ( .A1(n7516), .A2(n13348), .ZN(n7515) );
  INV_X1 U8458 ( .A(n13373), .ZN(n7514) );
  INV_X1 U8459 ( .A(n13371), .ZN(n7516) );
  AND2_X1 U8460 ( .A1(n7269), .A2(n7555), .ZN(n13360) );
  NAND2_X1 U8461 ( .A1(n13360), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n13395) );
  OR2_X1 U8462 ( .A1(n8757), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n13424) );
  NOR2_X1 U8463 ( .A1(n7772), .A2(n7771), .ZN(n7770) );
  INV_X1 U8464 ( .A(n8810), .ZN(n7772) );
  OR2_X1 U8465 ( .A1(n8738), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U8466 ( .A1(n13492), .A2(n13493), .ZN(n8809) );
  NAND2_X1 U8467 ( .A1(n8721), .A2(n8720), .ZN(n13494) );
  AOI21_X1 U8468 ( .B1(n7875), .B2(n7878), .A(n7234), .ZN(n7873) );
  INV_X1 U8469 ( .A(n7875), .ZN(n7874) );
  NAND2_X1 U8470 ( .A1(n8686), .A2(n8685), .ZN(n13533) );
  AND2_X1 U8471 ( .A1(n12709), .A2(n12710), .ZN(n13532) );
  INV_X1 U8472 ( .A(n12588), .ZN(n13546) );
  AND4_X1 U8473 ( .A1(n8655), .A2(n8654), .A3(n8653), .A4(n8652), .ZN(n13590)
         );
  NAND2_X1 U8474 ( .A1(n7753), .A2(n7388), .ZN(n7387) );
  AOI21_X1 U8475 ( .B1(n7753), .B2(n7756), .A(n7752), .ZN(n7751) );
  INV_X1 U8476 ( .A(n8802), .ZN(n13599) );
  NOR2_X1 U8477 ( .A1(n8614), .A2(n8290), .ZN(n8632) );
  INV_X1 U8478 ( .A(n12584), .ZN(n13638) );
  AOI21_X1 U8479 ( .B1(n7889), .B2(n7887), .A(n7886), .ZN(n7885) );
  INV_X1 U8480 ( .A(n7889), .ZN(n7888) );
  OAI21_X1 U8481 ( .B1(n11993), .B2(n7900), .A(n7898), .ZN(n12135) );
  NOR2_X1 U8482 ( .A1(n7901), .A2(n7904), .ZN(n7900) );
  AOI22_X1 U8483 ( .A1(n7901), .A2(n7903), .B1(n7904), .B2(n7899), .ZN(n7898)
         );
  AOI21_X1 U8484 ( .B1(n12647), .B2(n7906), .A(n7905), .ZN(n7904) );
  AND2_X1 U8485 ( .A1(n8476), .A2(n11890), .ZN(n8491) );
  INV_X1 U8486 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n11890) );
  INV_X1 U8487 ( .A(n12634), .ZN(n7750) );
  INV_X1 U8488 ( .A(n11631), .ZN(n12642) );
  NAND2_X1 U8489 ( .A1(n12576), .A2(n11171), .ZN(n15716) );
  AND2_X1 U8490 ( .A1(n12602), .A2(n13419), .ZN(n11183) );
  NAND2_X1 U8491 ( .A1(n8747), .A2(n8746), .ZN(n13217) );
  OR2_X1 U8492 ( .A1(n7221), .A2(n11714), .ZN(n8746) );
  NAND2_X1 U8493 ( .A1(n8724), .A2(n8723), .ZN(n13181) );
  INV_X1 U8494 ( .A(n15912), .ZN(n13729) );
  AOI21_X1 U8495 ( .B1(n7583), .B2(n7585), .A(n7581), .ZN(n7580) );
  INV_X1 U8496 ( .A(n8772), .ZN(n7581) );
  NAND2_X1 U8497 ( .A1(n8735), .A2(n8361), .ZN(n8745) );
  XNOR2_X1 U8498 ( .A(n8835), .B(n8284), .ZN(n10335) );
  NAND2_X1 U8499 ( .A1(n8661), .A2(n8660), .ZN(n8780) );
  INV_X1 U8500 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8660) );
  AND2_X1 U8501 ( .A1(n8341), .A2(n8340), .ZN(n8640) );
  NAND2_X1 U8502 ( .A1(n8330), .A2(n8331), .ZN(n8561) );
  AND2_X1 U8503 ( .A1(n8328), .A2(n8327), .ZN(n8550) );
  NOR2_X1 U8504 ( .A1(n7572), .A2(n7834), .ZN(n7571) );
  NOR2_X1 U8505 ( .A1(n10723), .A2(n10722), .ZN(n8008) );
  NAND2_X1 U8506 ( .A1(n8010), .A2(n13923), .ZN(n8009) );
  OAI22_X1 U8507 ( .A1(n13886), .A2(n8038), .B1(n13884), .B2(n13885), .ZN(
        n8037) );
  NAND2_X1 U8508 ( .A1(n8042), .A2(n13863), .ZN(n8038) );
  OR2_X1 U8509 ( .A1(n11127), .A2(n11569), .ZN(n11308) );
  INV_X1 U8510 ( .A(n8023), .ZN(n8022) );
  OR2_X1 U8511 ( .A1(n12215), .A2(n12253), .ZN(n8024) );
  INV_X1 U8512 ( .A(n8018), .ZN(n8012) );
  NAND2_X1 U8513 ( .A1(n8018), .A2(n13830), .ZN(n8013) );
  AND2_X1 U8514 ( .A1(n13878), .A2(n8016), .ZN(n8015) );
  OR2_X1 U8515 ( .A1(n12352), .A2(n13968), .ZN(n12365) );
  OR2_X1 U8516 ( .A1(n11290), .A2(n11289), .ZN(n8035) );
  XNOR2_X1 U8517 ( .A(n14408), .B(n7532), .ZN(n13829) );
  NAND2_X1 U8518 ( .A1(n13862), .A2(n13861), .ZN(n13863) );
  XNOR2_X1 U8519 ( .A(n12877), .B(n7532), .ZN(n13815) );
  OAI21_X1 U8520 ( .B1(n13043), .B2(n13037), .A(n13038), .ZN(n13036) );
  OR2_X1 U8521 ( .A1(n10360), .A2(n9698), .ZN(n10178) );
  AOI21_X1 U8522 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n10912), .A(n10318), .ZN(
        n10321) );
  NOR2_X1 U8523 ( .A1(n14029), .A2(n15388), .ZN(n14031) );
  NOR2_X1 U8524 ( .A1(n7843), .A2(n7841), .ZN(n7840) );
  NAND2_X1 U8525 ( .A1(n7842), .A2(n14437), .ZN(n7841) );
  NAND2_X1 U8526 ( .A1(n7935), .A2(n12465), .ZN(n7934) );
  INV_X1 U8527 ( .A(n12455), .ZN(n7935) );
  NAND2_X1 U8528 ( .A1(n13022), .A2(n12455), .ZN(n7936) );
  AND2_X1 U8529 ( .A1(n7932), .A2(n14309), .ZN(n7930) );
  AND2_X1 U8530 ( .A1(n12454), .A2(n12465), .ZN(n7932) );
  NAND2_X1 U8531 ( .A1(n14140), .A2(n14437), .ZN(n14119) );
  AND2_X1 U8532 ( .A1(n12431), .A2(n12430), .ZN(n14151) );
  NAND2_X1 U8533 ( .A1(n7943), .A2(n13021), .ZN(n14168) );
  INV_X1 U8534 ( .A(n14166), .ZN(n7943) );
  NAND2_X1 U8535 ( .A1(n14228), .A2(n14212), .ZN(n14206) );
  INV_X1 U8536 ( .A(n7839), .ZN(n14271) );
  NOR2_X1 U8537 ( .A1(n14313), .A2(n8069), .ZN(n8068) );
  NAND2_X1 U8538 ( .A1(n14282), .A2(n14288), .ZN(n14281) );
  OR2_X1 U8539 ( .A1(n11972), .A2(n11971), .ZN(n12061) );
  AOI21_X1 U8540 ( .B1(n8051), .B2(n8053), .A(n7274), .ZN(n8049) );
  AND2_X1 U8541 ( .A1(n7691), .A2(n13008), .ZN(n7484) );
  OR2_X1 U8542 ( .A1(n7949), .A2(n7692), .ZN(n7691) );
  INV_X1 U8543 ( .A(n11527), .ZN(n7692) );
  NAND2_X1 U8544 ( .A1(n11302), .A2(n11301), .ZN(n11304) );
  NAND2_X1 U8545 ( .A1(n11074), .A2(n11073), .ZN(n11076) );
  AND2_X1 U8546 ( .A1(n11026), .A2(n11016), .ZN(n8081) );
  NAND2_X1 U8547 ( .A1(n11030), .A2(n15864), .ZN(n11090) );
  NAND2_X1 U8548 ( .A1(n7372), .A2(n11009), .ZN(n11010) );
  NAND2_X1 U8549 ( .A1(n10932), .A2(n10832), .ZN(n10884) );
  INV_X1 U8550 ( .A(n13044), .ZN(n12963) );
  INV_X1 U8551 ( .A(n12190), .ZN(n12192) );
  NAND2_X1 U8552 ( .A1(n10825), .A2(n10824), .ZN(n10827) );
  NAND2_X1 U8553 ( .A1(n8046), .A2(n10820), .ZN(n10940) );
  NAND2_X1 U8554 ( .A1(n10953), .A2(n10956), .ZN(n8046) );
  OR2_X1 U8555 ( .A1(n10456), .A2(n10410), .ZN(n15778) );
  NAND2_X1 U8556 ( .A1(n8259), .A2(n13053), .ZN(n15963) );
  AND2_X1 U8557 ( .A1(n14507), .A2(n12963), .ZN(n15950) );
  AND2_X1 U8558 ( .A1(n10360), .A2(n13051), .ZN(n10470) );
  INV_X1 U8559 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9694) );
  INV_X1 U8560 ( .A(n9445), .ZN(n12375) );
  OR2_X1 U8561 ( .A1(n10781), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n11925) );
  OR2_X1 U8562 ( .A1(n10283), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n9931) );
  INV_X1 U8563 ( .A(n9861), .ZN(n7379) );
  OR2_X1 U8564 ( .A1(n14517), .A2(n14516), .ZN(n8274) );
  INV_X1 U8565 ( .A(n9416), .ZN(n9417) );
  AOI21_X1 U8566 ( .B1(n8121), .B2(n8123), .A(n7310), .ZN(n8119) );
  OAI21_X1 U8567 ( .B1(n8084), .B2(n8083), .A(n7255), .ZN(n8082) );
  INV_X1 U8568 ( .A(n11204), .ZN(n8083) );
  INV_X1 U8569 ( .A(n14748), .ZN(n10607) );
  NOR2_X1 U8570 ( .A1(n9355), .A2(n9352), .ZN(n9370) );
  NAND2_X1 U8571 ( .A1(n14671), .A2(n14579), .ZN(n14707) );
  NAND2_X1 U8572 ( .A1(n14547), .A2(n14546), .ZN(n14716) );
  XNOR2_X1 U8573 ( .A(n9747), .B(n14661), .ZN(n8088) );
  OR2_X1 U8574 ( .A1(n9229), .A2(n9228), .ZN(n9250) );
  OR2_X1 U8575 ( .A1(n9250), .A2(n9249), .ZN(n9276) );
  OAI22_X1 U8576 ( .A1(n9540), .A2(n7593), .B1(n7594), .B2(n9541), .ZN(n9609)
         );
  AND2_X1 U8577 ( .A1(n9541), .A2(n7594), .ZN(n7593) );
  INV_X1 U8578 ( .A(n9539), .ZN(n7594) );
  INV_X1 U8579 ( .A(n8994), .ZN(n9157) );
  OR2_X1 U8580 ( .A1(n9542), .A2(n10949), .ZN(n8999) );
  NAND2_X1 U8581 ( .A1(n9976), .A2(n9975), .ZN(n9974) );
  OR2_X1 U8582 ( .A1(n9994), .A2(n9995), .ZN(n7657) );
  NOR2_X1 U8583 ( .A1(n10094), .A2(n7670), .ZN(n10098) );
  AND2_X1 U8584 ( .A1(n10095), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7670) );
  NAND2_X1 U8585 ( .A1(n10098), .A2(n10097), .ZN(n10237) );
  XNOR2_X1 U8586 ( .A(n11589), .B(n9264), .ZN(n15429) );
  NAND2_X1 U8587 ( .A1(n7655), .A2(n7654), .ZN(n9333) );
  AND2_X1 U8588 ( .A1(n8914), .A2(n8915), .ZN(n7654) );
  INV_X1 U8589 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8915) );
  NOR2_X1 U8590 ( .A1(n14834), .A2(n14835), .ZN(n14833) );
  NAND2_X1 U8591 ( .A1(n9561), .A2(n9560), .ZN(n12529) );
  OR2_X1 U8592 ( .A1(n7725), .A2(n7724), .ZN(n14858) );
  INV_X1 U8593 ( .A(n15087), .ZN(n14861) );
  NOR2_X1 U8594 ( .A1(n7725), .A2(n15092), .ZN(n14880) );
  NAND2_X1 U8595 ( .A1(n14948), .A2(n14947), .ZN(n14946) );
  NAND2_X1 U8596 ( .A1(n14967), .A2(n7634), .ZN(n14941) );
  NAND2_X1 U8597 ( .A1(n14969), .A2(n14968), .ZN(n14967) );
  NAND2_X1 U8598 ( .A1(n7726), .A2(n15137), .ZN(n14960) );
  INV_X1 U8599 ( .A(n7726), .ZN(n15000) );
  OR2_X1 U8600 ( .A1(n9298), .A2(n9297), .ZN(n9355) );
  OR2_X1 U8601 ( .A1(n7717), .A2(n16013), .ZN(n15057) );
  NOR2_X1 U8602 ( .A1(n12269), .A2(n14739), .ZN(n12223) );
  NAND2_X1 U8603 ( .A1(n12017), .A2(n15955), .ZN(n12280) );
  NAND2_X1 U8604 ( .A1(n11478), .A2(n7720), .ZN(n11659) );
  AND2_X1 U8605 ( .A1(n11544), .A2(n7721), .ZN(n7720) );
  OR2_X1 U8606 ( .A1(n9115), .A2(n9114), .ZN(n9144) );
  NAND2_X1 U8607 ( .A1(n11478), .A2(n11544), .ZN(n11559) );
  NAND2_X1 U8608 ( .A1(n11152), .A2(n11339), .ZN(n11386) );
  NAND2_X1 U8609 ( .A1(n11149), .A2(n11159), .ZN(n11151) );
  NOR2_X1 U8610 ( .A1(n10654), .A2(n10658), .ZN(n10689) );
  XNOR2_X1 U8611 ( .A(n14749), .B(n10658), .ZN(n10646) );
  NAND2_X1 U8612 ( .A1(n9812), .A2(n9624), .ZN(n10699) );
  NAND2_X1 U8614 ( .A1(n7779), .A2(n7781), .ZN(n14847) );
  INV_X1 U8615 ( .A(n7781), .ZN(n7774) );
  AND2_X1 U8616 ( .A1(n15087), .A2(n16014), .ZN(n15088) );
  NAND2_X1 U8617 ( .A1(n15005), .A2(n12507), .ZN(n14993) );
  NAND2_X1 U8618 ( .A1(n9336), .A2(n9335), .ZN(n15153) );
  INV_X1 U8619 ( .A(n11283), .ZN(n7430) );
  NAND2_X1 U8620 ( .A1(n9142), .A2(n9141), .ZN(n11550) );
  OR2_X1 U8621 ( .A1(n11123), .A2(n9209), .ZN(n9142) );
  OR2_X1 U8622 ( .A1(n10059), .A2(n15217), .ZN(n10987) );
  INV_X1 U8623 ( .A(n16019), .ZN(n15799) );
  OR2_X1 U8624 ( .A1(n9774), .A2(n9773), .ZN(n15954) );
  INV_X1 U8625 ( .A(n15796), .ZN(n16009) );
  AND2_X1 U8626 ( .A1(n9781), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9665) );
  AND2_X1 U8627 ( .A1(n9591), .A2(n9570), .ZN(n13059) );
  OAI21_X1 U8628 ( .B1(n9656), .B2(P1_IR_REG_26__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8898) );
  XNOR2_X1 U8629 ( .A(n9529), .B(n12031), .ZN(n12498) );
  XNOR2_X1 U8630 ( .A(n9657), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9760) );
  INV_X1 U8631 ( .A(n8931), .ZN(n8924) );
  AND2_X1 U8632 ( .A1(n8932), .A2(n8931), .ZN(n9824) );
  NAND2_X1 U8633 ( .A1(n8183), .A2(n8181), .ZN(n9390) );
  NAND2_X1 U8634 ( .A1(n7415), .A2(n9346), .ZN(n9331) );
  NAND2_X1 U8635 ( .A1(n7416), .A2(n11833), .ZN(n7415) );
  NAND2_X1 U8636 ( .A1(n9329), .A2(n9328), .ZN(n7416) );
  NAND2_X1 U8637 ( .A1(n7793), .A2(n9346), .ZN(n9347) );
  NAND2_X1 U8638 ( .A1(n7655), .A2(n8914), .ZN(n9312) );
  NAND2_X1 U8639 ( .A1(n9105), .A2(n7719), .ZN(n9262) );
  NAND2_X1 U8640 ( .A1(n9238), .A2(n9237), .ZN(n9258) );
  NAND2_X1 U8641 ( .A1(n9165), .A2(n9164), .ZN(n9191) );
  NAND2_X1 U8642 ( .A1(n9138), .A2(n9137), .ZN(n9165) );
  NAND2_X1 U8643 ( .A1(n9133), .A2(n7426), .ZN(n9125) );
  AND2_X1 U8644 ( .A1(n8983), .A2(n9021), .ZN(n14766) );
  NAND2_X1 U8645 ( .A1(n8974), .A2(n8172), .ZN(n8979) );
  INV_X1 U8646 ( .A(n8909), .ZN(n8982) );
  INV_X1 U8647 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15224) );
  XNOR2_X1 U8648 ( .A(n15265), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n15274) );
  NOR2_X1 U8649 ( .A1(n15453), .A2(n15283), .ZN(n15288) );
  NOR2_X1 U8650 ( .A1(n15456), .A2(n15291), .ZN(n15294) );
  OAI21_X1 U8651 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n15244), .A(n15243), .ZN(
        n15308) );
  AND2_X1 U8652 ( .A1(n15487), .A2(n7403), .ZN(n15311) );
  OAI21_X1 U8653 ( .B1(n15489), .B2(n15488), .A(n7742), .ZN(n7403) );
  NAND2_X1 U8654 ( .A1(n7714), .A2(n7713), .ZN(n13123) );
  OAI21_X1 U8655 ( .B1(n13219), .B2(n13105), .A(n8139), .ZN(n7713) );
  NAND2_X1 U8656 ( .A1(n13218), .A2(n7241), .ZN(n7714) );
  NAND2_X1 U8657 ( .A1(n12300), .A2(n12299), .ZN(n12303) );
  AND2_X1 U8658 ( .A1(n8162), .A2(n13075), .ZN(n13136) );
  AOI21_X1 U8659 ( .B1(n8139), .B2(n13105), .A(n13108), .ZN(n8138) );
  NAND2_X1 U8660 ( .A1(n11578), .A2(n8153), .ZN(n12007) );
  INV_X1 U8661 ( .A(n13508), .ZN(n13486) );
  NOR2_X1 U8662 ( .A1(n11047), .A2(n11046), .ZN(n11049) );
  NAND2_X1 U8663 ( .A1(n10876), .A2(n11045), .ZN(n8154) );
  NAND2_X1 U8664 ( .A1(n11045), .A2(n7525), .ZN(n10875) );
  OR2_X1 U8665 ( .A1(n10874), .A2(n11238), .ZN(n7525) );
  NOR2_X1 U8666 ( .A1(n10876), .A2(n10875), .ZN(n11047) );
  NAND2_X1 U8667 ( .A1(n11578), .A2(n8150), .ZN(n8144) );
  NAND2_X1 U8668 ( .A1(n8678), .A2(n8677), .ZN(n13554) );
  NAND2_X1 U8669 ( .A1(n13088), .A2(n13090), .ZN(n13202) );
  NAND2_X1 U8670 ( .A1(n10712), .A2(n10711), .ZN(n10775) );
  INV_X1 U8671 ( .A(n13223), .ZN(n13237) );
  INV_X1 U8672 ( .A(n13230), .ZN(n7709) );
  NOR2_X1 U8673 ( .A1(n12600), .A2(n7764), .ZN(n7763) );
  OAI21_X1 U8674 ( .B1(n12747), .B2(n12746), .A(n12745), .ZN(n12748) );
  NAND2_X1 U8675 ( .A1(n12747), .A2(n12744), .ZN(n12745) );
  AOI21_X1 U8676 ( .B1(n7826), .B2(n12743), .A(n12742), .ZN(n12747) );
  INV_X1 U8677 ( .A(n13467), .ZN(n13244) );
  INV_X1 U8678 ( .A(n13656), .ZN(n13627) );
  OR2_X1 U8679 ( .A1(n10336), .A2(n9843), .ZN(n13263) );
  OR2_X1 U8680 ( .A1(n10257), .A2(n10256), .ZN(n10311) );
  NAND2_X1 U8681 ( .A1(n8554), .A2(n7392), .ZN(n7963) );
  AND2_X1 U8682 ( .A1(n8408), .A2(n8436), .ZN(n15521) );
  XNOR2_X1 U8683 ( .A(n11394), .B(n11456), .ZN(n15511) );
  INV_X1 U8684 ( .A(n7681), .ZN(n15527) );
  XNOR2_X1 U8685 ( .A(n7679), .B(n7678), .ZN(n15550) );
  NOR2_X1 U8686 ( .A1(n15550), .A2(n15551), .ZN(n15549) );
  NOR2_X1 U8687 ( .A1(n15549), .A2(n7502), .ZN(n15568) );
  AND2_X1 U8688 ( .A1(n7679), .A2(n7678), .ZN(n7502) );
  XNOR2_X1 U8689 ( .A(n11397), .B(n15601), .ZN(n15589) );
  INV_X1 U8690 ( .A(n7956), .ZN(n15588) );
  OAI22_X1 U8691 ( .A1(n15589), .A2(n7684), .B1(n15610), .B2(n7955), .ZN(
        n15609) );
  OR2_X1 U8692 ( .A1(n15610), .A2(n15590), .ZN(n7684) );
  INV_X1 U8693 ( .A(n7959), .ZN(n15647) );
  INV_X1 U8694 ( .A(n7957), .ZN(n11667) );
  XNOR2_X1 U8695 ( .A(n13286), .B(n13287), .ZN(n13266) );
  NOR2_X1 U8696 ( .A1(n13266), .A2(n13267), .ZN(n13288) );
  AND2_X1 U8697 ( .A1(n13281), .A2(n13280), .ZN(n13302) );
  OAI21_X1 U8698 ( .B1(n7961), .B2(n13266), .A(n7960), .ZN(n13310) );
  NAND2_X1 U8699 ( .A1(n7962), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7961) );
  NAND2_X1 U8700 ( .A1(n13289), .A2(n7962), .ZN(n7960) );
  INV_X1 U8701 ( .A(n13291), .ZN(n7962) );
  INV_X1 U8702 ( .A(n7969), .ZN(n13329) );
  OR2_X1 U8703 ( .A1(n13311), .A2(n13312), .ZN(n7969) );
  INV_X1 U8704 ( .A(n13330), .ZN(n7968) );
  NAND2_X1 U8705 ( .A1(n7965), .A2(n7966), .ZN(n13362) );
  OAI21_X1 U8706 ( .B1(n15657), .B2(n13379), .A(n13369), .ZN(n7687) );
  AOI21_X1 U8707 ( .B1(n13395), .B2(n7269), .A(n13394), .ZN(n13402) );
  OAI21_X1 U8708 ( .B1(n8795), .B2(n15719), .A(n8794), .ZN(n13429) );
  AND2_X1 U8709 ( .A1(n13442), .A2(n13441), .ZN(n13676) );
  OR2_X1 U8710 ( .A1(n7221), .A2(n12031), .ZN(n8754) );
  NAND2_X1 U8711 ( .A1(n13480), .A2(n13464), .ZN(n13465) );
  NAND2_X1 U8712 ( .A1(n7872), .A2(n8698), .ZN(n13520) );
  NAND2_X1 U8713 ( .A1(n8686), .A2(n7877), .ZN(n7872) );
  NAND2_X1 U8714 ( .A1(n13588), .A2(n8639), .ZN(n13577) );
  NAND2_X1 U8715 ( .A1(n13620), .A2(n12684), .ZN(n13605) );
  INV_X1 U8716 ( .A(n7393), .ZN(n13666) );
  AOI21_X1 U8717 ( .B1(n12205), .B2(n7760), .A(n7396), .ZN(n7393) );
  AND2_X1 U8718 ( .A1(n8569), .A2(n8568), .ZN(n13664) );
  NAND2_X1 U8719 ( .A1(n7890), .A2(n8559), .ZN(n13655) );
  NAND2_X1 U8720 ( .A1(n8542), .A2(n8541), .ZN(n12311) );
  AND3_X1 U8721 ( .A1(n8558), .A2(n8557), .A3(n8556), .ZN(n12316) );
  NAND2_X1 U8722 ( .A1(n7759), .A2(n12666), .ZN(n12317) );
  NAND2_X1 U8723 ( .A1(n12205), .A2(n12664), .ZN(n7759) );
  NAND2_X1 U8724 ( .A1(n10595), .A2(n15695), .ZN(n13650) );
  NAND2_X1 U8725 ( .A1(n11995), .A2(n8490), .ZN(n11944) );
  NAND2_X1 U8726 ( .A1(n11239), .A2(n12634), .ZN(n11267) );
  NAND2_X1 U8727 ( .A1(n7897), .A2(n8426), .ZN(n11236) );
  INV_X1 U8728 ( .A(n10714), .ZN(n15730) );
  NAND2_X1 U8729 ( .A1(n10355), .A2(n10354), .ZN(n15727) );
  AND2_X2 U8730 ( .A1(n10591), .A2(n8856), .ZN(n15940) );
  INV_X1 U8731 ( .A(n13421), .ZN(n13745) );
  INV_X1 U8732 ( .A(n12566), .ZN(n13748) );
  INV_X1 U8733 ( .A(n13116), .ZN(n13752) );
  INV_X1 U8734 ( .A(n13181), .ZN(n13762) );
  NAND2_X1 U8736 ( .A1(n15944), .A2(n15891), .ZN(n13794) );
  INV_X1 U8737 ( .A(n15944), .ZN(n15941) );
  INV_X1 U8738 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8285) );
  INV_X1 U8739 ( .A(n8289), .ZN(n13812) );
  NAND2_X1 U8740 ( .A1(n7582), .A2(n8367), .ZN(n8771) );
  INV_X1 U8741 ( .A(SI_26_), .ZN(n11714) );
  XNOR2_X1 U8742 ( .A(n8821), .B(n8820), .ZN(n11328) );
  INV_X1 U8743 ( .A(SI_24_), .ZN(n11828) );
  NAND2_X1 U8744 ( .A1(n8834), .A2(n8284), .ZN(n7498) );
  OAI21_X1 U8745 ( .B1(n8350), .B2(n8699), .A(n7590), .ZN(n8711) );
  NAND2_X1 U8746 ( .A1(n8350), .A2(n8349), .ZN(n8700) );
  NAND2_X1 U8747 ( .A1(n8497), .A2(n7924), .ZN(n8784) );
  AND2_X1 U8748 ( .A1(n8166), .A2(n7925), .ZN(n7924) );
  NOR2_X1 U8749 ( .A1(n10404), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13798) );
  NAND2_X1 U8750 ( .A1(n8657), .A2(n8656), .ZN(n8659) );
  NAND2_X1 U8751 ( .A1(n8643), .A2(n8341), .ZN(n8657) );
  OAI21_X1 U8752 ( .B1(n8596), .B2(n7563), .A(n7560), .ZN(n8624) );
  NAND2_X1 U8753 ( .A1(n8608), .A2(n8607), .ZN(n8610) );
  NAND2_X1 U8754 ( .A1(n8596), .A2(n8335), .ZN(n8608) );
  INV_X1 U8755 ( .A(SI_16_), .ZN(n11845) );
  INV_X1 U8756 ( .A(SI_15_), .ZN(n11711) );
  NAND2_X1 U8757 ( .A1(n8279), .A2(n8514), .ZN(n8597) );
  INV_X1 U8758 ( .A(SI_14_), .ZN(n11818) );
  NAND2_X1 U8759 ( .A1(n8563), .A2(n8331), .ZN(n8577) );
  XNOR2_X1 U8760 ( .A(n8582), .B(n8581), .ZN(n13321) );
  INV_X1 U8761 ( .A(SI_13_), .ZN(n11848) );
  INV_X1 U8762 ( .A(SI_11_), .ZN(n9920) );
  NAND2_X1 U8763 ( .A1(n7836), .A2(n7833), .ZN(n8471) );
  NAND2_X1 U8764 ( .A1(n7836), .A2(n8316), .ZN(n8469) );
  NAND2_X1 U8765 ( .A1(n8312), .A2(n8311), .ZN(n8435) );
  INV_X1 U8766 ( .A(n7820), .ZN(n8406) );
  AOI21_X1 U8767 ( .B1(n8395), .B2(n8394), .A(n7821), .ZN(n7820) );
  INV_X1 U8768 ( .A(n15521), .ZN(n11456) );
  INV_X1 U8769 ( .A(n8303), .ZN(n8377) );
  NAND2_X1 U8770 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7677) );
  NAND2_X1 U8771 ( .A1(n8011), .A2(n7496), .ZN(n10732) );
  OR2_X1 U8772 ( .A1(n10731), .A2(n10730), .ZN(n7496) );
  NAND2_X1 U8773 ( .A1(n8009), .A2(n8007), .ZN(n10733) );
  INV_X1 U8774 ( .A(n8008), .ZN(n8007) );
  NAND2_X1 U8775 ( .A1(n10729), .A2(n10728), .ZN(n15844) );
  INV_X1 U8776 ( .A(n14437), .ZN(n14122) );
  INV_X1 U8777 ( .A(n12873), .ZN(n15964) );
  NAND2_X1 U8778 ( .A1(n13957), .A2(n14262), .ZN(n13998) );
  NAND2_X1 U8779 ( .A1(n8014), .A2(n13830), .ZN(n13879) );
  NAND2_X1 U8780 ( .A1(n13984), .A2(n13985), .ZN(n8014) );
  OAI21_X1 U8781 ( .B1(n13860), .B2(n8039), .A(n8036), .ZN(n13891) );
  OR2_X1 U8782 ( .A1(n13886), .A2(n8040), .ZN(n8039) );
  INV_X1 U8783 ( .A(n8037), .ZN(n8036) );
  INV_X1 U8784 ( .A(n13863), .ZN(n8040) );
  NAND2_X1 U8785 ( .A1(n8026), .A2(n8030), .ZN(n11961) );
  OR2_X1 U8786 ( .A1(n11290), .A2(n8031), .ZN(n8026) );
  XNOR2_X1 U8787 ( .A(n13858), .B(n13856), .ZN(n13905) );
  NAND2_X1 U8788 ( .A1(n12413), .A2(n12412), .ZN(n14158) );
  OR2_X1 U8789 ( .A1(n10475), .A2(n13053), .ZN(n13939) );
  NAND2_X1 U8790 ( .A1(n8021), .A2(n8022), .ZN(n13915) );
  NAND2_X1 U8791 ( .A1(n10552), .A2(n10551), .ZN(n15804) );
  OR2_X1 U8792 ( .A1(n10549), .A2(n10521), .ZN(n10552) );
  NAND2_X1 U8793 ( .A1(n13913), .A2(n13822), .ZN(n13936) );
  INV_X1 U8794 ( .A(n13944), .ZN(n8002) );
  NAND2_X1 U8795 ( .A1(n13870), .A2(n13851), .ZN(n13945) );
  AND2_X1 U8796 ( .A1(n7436), .A2(n7438), .ZN(n13954) );
  NOR2_X1 U8797 ( .A1(n11110), .A2(n11109), .ZN(n11114) );
  INV_X1 U8798 ( .A(n14003), .ZN(n13966) );
  XNOR2_X1 U8799 ( .A(n13844), .B(n13842), .ZN(n13976) );
  AND2_X1 U8800 ( .A1(n8035), .A2(n11566), .ZN(n11957) );
  INV_X1 U8801 ( .A(n7437), .ZN(n10519) );
  INV_X1 U8802 ( .A(n13939), .ZN(n13957) );
  NAND2_X1 U8803 ( .A1(n10577), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13995) );
  NAND2_X1 U8804 ( .A1(n13860), .A2(n13859), .ZN(n13992) );
  NAND2_X1 U8805 ( .A1(n12255), .A2(n12254), .ZN(n13819) );
  NAND2_X1 U8806 ( .A1(n10478), .A2(n14318), .ZN(n14001) );
  NAND2_X1 U8807 ( .A1(n12452), .A2(n12451), .ZN(n14114) );
  OR2_X1 U8808 ( .A1(n14105), .A2(n12458), .ZN(n12452) );
  INV_X1 U8809 ( .A(n14135), .ZN(n14101) );
  NAND4_X1 U8810 ( .A1(n10548), .A2(n10547), .A3(n10546), .A4(n10545), .ZN(
        n14021) );
  NAND2_X1 U8811 ( .A1(n10529), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n10403) );
  OR2_X2 U8812 ( .A1(n10178), .A2(P2_U3088), .ZN(n14025) );
  AOI21_X1 U8813 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n15350), .A(n15342), .ZN(
        n10223) );
  AOI21_X1 U8814 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n10226), .A(n10221), .ZN(
        n15355) );
  AOI21_X1 U8815 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n15372), .A(n15367), .ZN(
        n10213) );
  AOI21_X1 U8816 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n15372), .A(n15364), .ZN(
        n10210) );
  AOI21_X1 U8817 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n15384), .A(n15376), .ZN(
        n10202) );
  AOI21_X1 U8818 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n15384), .A(n15379), .ZN(
        n10199) );
  AOI21_X1 U8819 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n10727), .A(n10197), .ZN(
        n10183) );
  NOR2_X1 U8820 ( .A1(n11355), .A2(n7479), .ZN(n15418) );
  AND2_X1 U8821 ( .A1(n11361), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7479) );
  NAND2_X1 U8822 ( .A1(n15418), .A2(n15417), .ZN(n15416) );
  INV_X1 U8823 ( .A(n7478), .ZN(n14026) );
  NAND2_X1 U8824 ( .A1(n15395), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n15394) );
  OR2_X1 U8825 ( .A1(n14031), .A2(n14030), .ZN(n14057) );
  AND2_X1 U8826 ( .A1(n14051), .A2(n14050), .ZN(n15407) );
  AND2_X1 U8827 ( .A1(n14062), .A2(n14076), .ZN(n14063) );
  OR2_X1 U8828 ( .A1(n14061), .A2(n14060), .ZN(n14062) );
  NAND2_X1 U8829 ( .A1(n14177), .A2(n12490), .ZN(n14155) );
  AND2_X1 U8830 ( .A1(n12402), .A2(n12401), .ZN(n14372) );
  AND2_X1 U8831 ( .A1(n14192), .A2(n14191), .ZN(n14382) );
  AOI21_X1 U8832 ( .B1(n12486), .B2(n8065), .A(n8067), .ZN(n14214) );
  INV_X1 U8833 ( .A(n14386), .ZN(n14212) );
  NAND2_X1 U8834 ( .A1(n14225), .A2(n12373), .ZN(n14203) );
  AND2_X1 U8835 ( .A1(n14270), .A2(n14269), .ZN(n14403) );
  NAND2_X1 U8836 ( .A1(n12480), .A2(n12479), .ZN(n14314) );
  NAND2_X1 U8837 ( .A1(n12176), .A2(n12175), .ZN(n12177) );
  NOR2_X1 U8838 ( .A1(n8070), .A2(n7225), .ZN(n12198) );
  INV_X1 U8839 ( .A(n12196), .ZN(n8070) );
  NAND2_X1 U8840 ( .A1(n8050), .A2(n11608), .ZN(n11984) );
  NAND2_X1 U8841 ( .A1(n11607), .A2(n11606), .ZN(n8050) );
  NAND2_X1 U8842 ( .A1(n8076), .A2(n11316), .ZN(n11317) );
  NAND2_X1 U8843 ( .A1(n11122), .A2(n11121), .ZN(n11315) );
  NAND2_X1 U8844 ( .A1(n11070), .A2(n11069), .ZN(n12836) );
  INV_X1 U8845 ( .A(n9870), .ZN(n10522) );
  INV_X1 U8846 ( .A(n15818), .ZN(n14301) );
  INV_X1 U8847 ( .A(n14318), .ZN(n15816) );
  INV_X1 U8848 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7846) );
  INV_X1 U8849 ( .A(n14330), .ZN(n14427) );
  NAND2_X1 U8850 ( .A1(n14329), .A2(n14331), .ZN(n14424) );
  AND2_X1 U8851 ( .A1(n12422), .A2(n12421), .ZN(n14441) );
  NAND2_X1 U8852 ( .A1(n14360), .A2(n7485), .ZN(n14438) );
  INV_X1 U8853 ( .A(n7486), .ZN(n7485) );
  OAI21_X1 U8854 ( .B1(n14361), .B2(n15847), .A(n14359), .ZN(n7486) );
  INV_X1 U8855 ( .A(n14158), .ZN(n14445) );
  INV_X1 U8856 ( .A(n14320), .ZN(n14468) );
  NAND2_X1 U8857 ( .A1(n10388), .A2(n10387), .ZN(n15339) );
  OR2_X1 U8858 ( .A1(n14490), .A2(n10386), .ZN(n10387) );
  NAND2_X1 U8859 ( .A1(n15335), .A2(n15338), .ZN(n10388) );
  AND2_X1 U8860 ( .A1(n8054), .A2(n7375), .ZN(n7944) );
  INV_X1 U8861 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n14475) );
  NAND2_X1 U8862 ( .A1(n7538), .A2(n7537), .ZN(n10175) );
  NAND2_X1 U8863 ( .A1(n10170), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7537) );
  XNOR2_X1 U8864 ( .A(n9689), .B(P2_IR_REG_26__SCAN_IN), .ZN(n14490) );
  NAND2_X1 U8865 ( .A1(n9692), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9689) );
  NAND2_X1 U8866 ( .A1(n9693), .A2(n9692), .ZN(n14495) );
  XNOR2_X1 U8867 ( .A(n9695), .B(n9694), .ZN(n14498) );
  INV_X1 U8868 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12349) );
  NAND2_X1 U8869 ( .A1(n10379), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n10380) );
  INV_X1 U8870 ( .A(n14078), .ZN(n14073) );
  INV_X1 U8871 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11284) );
  INV_X1 U8872 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10287) );
  AND2_X1 U8873 ( .A1(n10085), .A2(n10053), .ZN(n11124) );
  INV_X1 U8874 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9933) );
  INV_X1 U8875 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9930) );
  INV_X1 U8876 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9883) );
  INV_X1 U8877 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9859) );
  INV_X1 U8878 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9865) );
  INV_X1 U8879 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9871) );
  INV_X1 U8880 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10446) );
  INV_X1 U8881 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10396) );
  NAND2_X1 U8882 ( .A1(n9848), .A2(n9847), .ZN(n10398) );
  NAND2_X1 U8883 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n9845) );
  XNOR2_X1 U8884 ( .A(n9651), .B(n9650), .ZN(n9889) );
  INV_X1 U8885 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9650) );
  OAI21_X1 U8886 ( .B1(n9649), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9651) );
  AOI21_X1 U8887 ( .B1(n7355), .B2(n8093), .A(n8084), .ZN(n11205) );
  INV_X1 U8888 ( .A(n14658), .ZN(n7552) );
  NAND2_X1 U8889 ( .A1(n14518), .A2(n8274), .ZN(n14631) );
  AND2_X1 U8890 ( .A1(n8098), .A2(n7349), .ZN(n11507) );
  NAND2_X1 U8891 ( .A1(n8108), .A2(n14554), .ZN(n14648) );
  NAND2_X1 U8892 ( .A1(n7542), .A2(n14717), .ZN(n8108) );
  AND2_X1 U8893 ( .A1(n8121), .A2(n8124), .ZN(n8114) );
  OAI22_X1 U8894 ( .A1(n8117), .A2(n8116), .B1(n8124), .B2(n8119), .ZN(n8115)
         );
  NOR2_X1 U8895 ( .A1(n8121), .A2(n8124), .ZN(n8117) );
  INV_X1 U8896 ( .A(n8119), .ZN(n8116) );
  NAND2_X1 U8897 ( .A1(n8119), .A2(n14665), .ZN(n8118) );
  NAND2_X1 U8898 ( .A1(n14698), .A2(n14571), .ZN(n14673) );
  NAND2_X1 U8899 ( .A1(n7810), .A2(n9391), .ZN(n14961) );
  NAND2_X1 U8900 ( .A1(n12361), .A2(n9595), .ZN(n7810) );
  AOI21_X1 U8901 ( .B1(n7228), .B2(n8105), .A(n7285), .ZN(n8101) );
  NAND2_X1 U8902 ( .A1(n9476), .A2(n9475), .ZN(n14895) );
  CLKBUF_X1 U8903 ( .A(n15997), .Z(n15998) );
  NAND2_X1 U8904 ( .A1(n8093), .A2(n10943), .ZN(n10802) );
  NAND2_X1 U8905 ( .A1(n8103), .A2(n14597), .ZN(n14687) );
  NAND2_X1 U8906 ( .A1(n14640), .A2(n14641), .ZN(n8103) );
  NAND2_X1 U8907 ( .A1(n9132), .A2(n9131), .ZN(n11486) );
  INV_X1 U8908 ( .A(n15679), .ZN(n10061) );
  NOR2_X1 U8909 ( .A1(n11935), .A2(n8096), .ZN(n8095) );
  INV_X1 U8910 ( .A(n8099), .ZN(n8096) );
  NAND2_X1 U8911 ( .A1(n11932), .A2(n8099), .ZN(n11934) );
  NAND2_X1 U8912 ( .A1(n14691), .A2(n15034), .ZN(n14728) );
  CLKBUF_X1 U8913 ( .A(n14716), .Z(n7542) );
  NAND2_X1 U8914 ( .A1(n8091), .A2(n10799), .ZN(n10994) );
  NAND2_X1 U8915 ( .A1(n7356), .A2(n8093), .ZN(n8091) );
  XNOR2_X1 U8916 ( .A(n14529), .B(n14530), .ZN(n15976) );
  NAND2_X1 U8917 ( .A1(n10045), .A2(P1_STATE_REG_SCAN_IN), .ZN(n16041) );
  INV_X1 U8918 ( .A(n14733), .ZN(n16036) );
  NAND2_X1 U8919 ( .A1(n7599), .A2(n7601), .ZN(n8953) );
  OR2_X1 U8920 ( .A1(n9031), .A2(n8951), .ZN(n8956) );
  NAND2_X1 U8921 ( .A1(n9974), .A2(n7658), .ZN(n9994) );
  OR2_X1 U8922 ( .A1(n9961), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7658) );
  INV_X1 U8923 ( .A(n7657), .ZN(n9993) );
  AND2_X1 U8924 ( .A1(n7657), .A2(n7656), .ZN(n9947) );
  NAND2_X1 U8925 ( .A1(n9963), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7656) );
  NOR2_X1 U8926 ( .A1(n10002), .A2(n7667), .ZN(n10005) );
  AND2_X1 U8927 ( .A1(n10003), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7667) );
  NAND2_X1 U8928 ( .A1(n10005), .A2(n10004), .ZN(n10021) );
  NAND2_X1 U8929 ( .A1(n10021), .A2(n7664), .ZN(n10022) );
  NAND2_X1 U8930 ( .A1(n7666), .A2(n7665), .ZN(n7664) );
  NAND2_X1 U8931 ( .A1(n10022), .A2(n10023), .ZN(n10068) );
  NAND2_X1 U8932 ( .A1(n10237), .A2(n7669), .ZN(n10238) );
  OR2_X1 U8933 ( .A1(n10241), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7669) );
  NAND2_X1 U8934 ( .A1(n10238), .A2(n10239), .ZN(n10632) );
  OR2_X1 U8935 ( .A1(n10864), .A2(n10863), .ZN(n11586) );
  OAI21_X1 U8936 ( .B1(n14824), .B2(n14823), .A(n7662), .ZN(n7661) );
  OR2_X1 U8937 ( .A1(n14822), .A2(n15434), .ZN(n7662) );
  INV_X1 U8938 ( .A(n12529), .ZN(n15075) );
  INV_X1 U8939 ( .A(n7776), .ZN(n7775) );
  OR2_X1 U8940 ( .A1(n15081), .A2(n14871), .ZN(n12514) );
  XNOR2_X1 U8941 ( .A(n7367), .B(n14857), .ZN(n15086) );
  NAND2_X1 U8942 ( .A1(n8190), .A2(n8189), .ZN(n14867) );
  NAND2_X1 U8943 ( .A1(n14891), .A2(n8266), .ZN(n14875) );
  NOR2_X1 U8944 ( .A1(n15108), .A2(n8194), .ZN(n14893) );
  NAND2_X1 U8945 ( .A1(n14903), .A2(n7998), .ZN(n14890) );
  INV_X1 U8946 ( .A(n14961), .ZN(n15129) );
  NAND2_X1 U8947 ( .A1(n14973), .A2(n8264), .ZN(n14958) );
  NAND2_X1 U8948 ( .A1(n14991), .A2(n12508), .ZN(n14983) );
  AND2_X1 U8949 ( .A1(n14996), .A2(n12519), .ZN(n14974) );
  AND2_X1 U8950 ( .A1(n7990), .A2(n7989), .ZN(n15013) );
  NAND2_X1 U8951 ( .A1(n15045), .A2(n12518), .ZN(n15030) );
  NAND2_X1 U8952 ( .A1(n7637), .A2(n7635), .ZN(n15987) );
  NOR2_X1 U8953 ( .A1(n12237), .A2(n7636), .ZN(n7635) );
  INV_X1 U8954 ( .A(n12235), .ZN(n7636) );
  NAND2_X1 U8955 ( .A1(n7637), .A2(n12235), .ZN(n12238) );
  INV_X1 U8956 ( .A(n15165), .ZN(n14521) );
  NAND2_X1 U8957 ( .A1(n12233), .A2(n12232), .ZN(n12278) );
  NAND2_X1 U8958 ( .A1(n9195), .A2(n9194), .ZN(n12127) );
  NAND2_X1 U8959 ( .A1(n11645), .A2(n11644), .ZN(n11646) );
  INV_X1 U8960 ( .A(n14988), .ZN(n15048) );
  AND2_X1 U8961 ( .A1(n7855), .A2(n7856), .ZN(n9829) );
  NAND2_X1 U8962 ( .A1(n7976), .A2(n9801), .ZN(n10786) );
  NAND2_X1 U8963 ( .A1(n7978), .A2(n7977), .ZN(n7976) );
  NAND2_X1 U8964 ( .A1(n7865), .A2(n9816), .ZN(n10686) );
  NAND2_X1 U8965 ( .A1(n7978), .A2(n9799), .ZN(n10684) );
  INV_X1 U8966 ( .A(n15681), .ZN(n15018) );
  OR2_X1 U8967 ( .A1(n10063), .A2(n9888), .ZN(n15035) );
  OAI211_X1 U8968 ( .C1(n9209), .C2(n10449), .A(n8912), .B(n8911), .ZN(n10514)
         );
  INV_X1 U8969 ( .A(n15055), .ZN(n15036) );
  OR2_X1 U8970 ( .A1(n15020), .A2(n9838), .ZN(n15680) );
  NAND2_X1 U8971 ( .A1(n9624), .A2(n9625), .ZN(n15683) );
  OR2_X1 U8972 ( .A1(n9757), .A2(n9760), .ZN(n9875) );
  XNOR2_X1 U8973 ( .A(n9594), .B(n9593), .ZN(n15194) );
  INV_X1 U8974 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8881) );
  NAND2_X1 U8975 ( .A1(n7642), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8882) );
  MUX2_X1 U8976 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8895), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n8896) );
  XNOR2_X1 U8977 ( .A(n9535), .B(n9534), .ZN(n14483) );
  CLKBUF_X1 U8978 ( .A(n9666), .Z(n12531) );
  INV_X1 U8979 ( .A(n9760), .ZN(n15203) );
  AND2_X1 U8980 ( .A1(n9660), .A2(n9656), .ZN(n15204) );
  MUX2_X1 U8981 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9663), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9664) );
  XNOR2_X1 U8982 ( .A(n9425), .B(n9424), .ZN(n15211) );
  AND2_X1 U8983 ( .A1(n10404), .A2(P1_U3086), .ZN(n15212) );
  XNOR2_X1 U8984 ( .A(n9399), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15218) );
  INV_X1 U8985 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11666) );
  INV_X2 U8986 ( .A(n9824), .ZN(n11665) );
  NAND2_X1 U8987 ( .A1(n9332), .A2(n9347), .ZN(n11283) );
  INV_X1 U8988 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11038) );
  INV_X1 U8989 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10895) );
  INV_X1 U8990 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10785) );
  INV_X1 U8991 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10582) );
  NAND2_X1 U8992 ( .A1(n9202), .A2(n9201), .ZN(n9207) );
  INV_X1 U8993 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10276) );
  INV_X1 U8994 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10084) );
  INV_X1 U8995 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10056) );
  NAND2_X1 U8996 ( .A1(n9139), .A2(n9165), .ZN(n11123) );
  OR2_X1 U8997 ( .A1(n9138), .A2(n9137), .ZN(n9139) );
  INV_X1 U8998 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10040) );
  INV_X1 U8999 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9934) );
  NAND2_X1 U9000 ( .A1(n9102), .A2(n9101), .ZN(n9123) );
  NAND2_X1 U9001 ( .A1(n7701), .A2(n7271), .ZN(n9102) );
  OR2_X1 U9002 ( .A1(n9046), .A2(n9045), .ZN(n9047) );
  XNOR2_X1 U9003 ( .A(n7671), .B(P1_IR_REG_4__SCAN_IN), .ZN(n14782) );
  NAND2_X1 U9004 ( .A1(n9021), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7671) );
  NAND2_X1 U9005 ( .A1(n8942), .A2(n8972), .ZN(n8944) );
  NOR2_X1 U9006 ( .A1(n15507), .A2(n15273), .ZN(n15444) );
  XNOR2_X1 U9007 ( .A(n15275), .B(n7736), .ZN(n15449) );
  INV_X1 U9008 ( .A(n15274), .ZN(n7736) );
  NAND2_X1 U9009 ( .A1(n7732), .A2(n15282), .ZN(n7731) );
  OAI21_X1 U9010 ( .B1(n15450), .B2(n15277), .A(n7730), .ZN(n7729) );
  INV_X1 U9011 ( .A(n15282), .ZN(n7730) );
  AND2_X1 U9012 ( .A1(n7729), .A2(n7407), .ZN(n15453) );
  NOR2_X1 U9013 ( .A1(n7728), .A2(n15454), .ZN(n7407) );
  OR2_X1 U9014 ( .A1(n15288), .A2(n15287), .ZN(n15505) );
  NAND2_X1 U9015 ( .A1(n15505), .A2(n15506), .ZN(n15502) );
  XNOR2_X1 U9016 ( .A(n15290), .B(n7745), .ZN(n15457) );
  NOR2_X1 U9017 ( .A1(n15457), .A2(n15458), .ZN(n15456) );
  NAND2_X1 U9018 ( .A1(n7406), .A2(n15462), .ZN(n15467) );
  NOR2_X1 U9019 ( .A1(n15467), .A2(n15468), .ZN(n15466) );
  NAND2_X1 U9020 ( .A1(n15476), .A2(n15307), .ZN(n15481) );
  INV_X1 U9021 ( .A(n7744), .ZN(n15306) );
  NAND2_X1 U9022 ( .A1(n15481), .A2(n15480), .ZN(n15479) );
  NAND2_X1 U9023 ( .A1(n7405), .A2(n15479), .ZN(n15484) );
  OAI21_X1 U9024 ( .B1(n15481), .B2(n15480), .A(n7506), .ZN(n7405) );
  INV_X1 U9025 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7506) );
  OAI21_X1 U9026 ( .B1(n15310), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n15483), .ZN(
        n15489) );
  NOR2_X1 U9027 ( .A1(n15484), .A2(n15485), .ZN(n15310) );
  NAND2_X1 U9028 ( .A1(n15489), .A2(n15488), .ZN(n15487) );
  NOR2_X1 U9029 ( .A1(n15311), .A2(n15312), .ZN(n15492) );
  NAND2_X1 U9030 ( .A1(n15311), .A2(n15312), .ZN(n15494) );
  NAND2_X1 U9031 ( .A1(n15494), .A2(n15495), .ZN(n15491) );
  NOR2_X1 U9032 ( .A1(n15496), .A2(n15314), .ZN(n15501) );
  INV_X1 U9033 ( .A(n13263), .ZN(P3_U3897) );
  NAND2_X1 U9034 ( .A1(n7688), .A2(n7685), .ZN(P3_U3199) );
  AOI21_X1 U9035 ( .B1(n13377), .B2(n15667), .A(n7686), .ZN(n7685) );
  NAND2_X1 U9036 ( .A1(n13367), .A2(n13368), .ZN(n7688) );
  OR2_X1 U9037 ( .A1(n13376), .A2(n7687), .ZN(n7686) );
  OAI211_X1 U9038 ( .C1(n7973), .C2(n15671), .A(n7401), .B(n7287), .ZN(
        P3_U3201) );
  XNOR2_X1 U9039 ( .A(n13417), .B(n13416), .ZN(n7973) );
  NAND2_X1 U9040 ( .A1(n7402), .A2(n15667), .ZN(n7401) );
  NAND2_X1 U9041 ( .A1(n7421), .A2(n7243), .ZN(n7550) );
  AOI211_X1 U9042 ( .C1(n14336), .C2(n15823), .A(n12496), .B(n12495), .ZN(
        n12497) );
  NAND2_X1 U9043 ( .A1(n7368), .A2(n14275), .ZN(n14110) );
  NAND2_X1 U9044 ( .A1(n7847), .A2(n7844), .ZN(P2_U3530) );
  AOI21_X1 U9045 ( .B1(n14330), .B2(n14422), .A(n7845), .ZN(n7844) );
  NAND2_X1 U9046 ( .A1(n14424), .A2(n15970), .ZN(n7847) );
  NOR2_X1 U9047 ( .A1(n15970), .A2(n7846), .ZN(n7845) );
  NAND2_X1 U9048 ( .A1(n14357), .A2(n14356), .ZN(n14358) );
  NAND2_X1 U9049 ( .A1(n7377), .A2(n7376), .ZN(P2_U3495) );
  NAND2_X1 U9050 ( .A1(n15971), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7376) );
  OAI21_X1 U9051 ( .B1(n9655), .B2(n9654), .A(n9653), .ZN(n9670) );
  NAND2_X1 U9052 ( .A1(n7663), .A2(n7659), .ZN(P1_U3262) );
  AOI21_X1 U9053 ( .B1(n7661), .B2(n14825), .A(n7660), .ZN(n7659) );
  NAND2_X1 U9054 ( .A1(n14826), .A2(n9348), .ZN(n7663) );
  OAI21_X1 U9055 ( .B1(n15440), .B2(n8167), .A(n14827), .ZN(n7660) );
  XNOR2_X1 U9056 ( .A(n7734), .B(n7733), .ZN(SUB_1596_U62) );
  INV_X1 U9057 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n7733) );
  NOR2_X1 U9058 ( .A1(n15499), .A2(n7735), .ZN(n7734) );
  AND2_X1 U9059 ( .A1(n15501), .A2(n15500), .ZN(n7735) );
  INV_X1 U9060 ( .A(n11457), .ZN(n7678) );
  AND2_X1 U9061 ( .A1(n14748), .A2(n10691), .ZN(n7224) );
  XNOR2_X1 U9062 ( .A(n14961), .B(n14976), .ZN(n14968) );
  INV_X1 U9063 ( .A(n14968), .ZN(n14957) );
  XNOR2_X1 U9064 ( .A(n11550), .B(n14742), .ZN(n11542) );
  NAND2_X1 U9065 ( .A1(n15092), .A2(n14896), .ZN(n7786) );
  NOR2_X1 U9066 ( .A1(n12877), .A2(n14011), .ZN(n7225) );
  AND2_X1 U9067 ( .A1(n7307), .A2(n12373), .ZN(n7226) );
  AND2_X1 U9068 ( .A1(n8201), .A2(n8200), .ZN(n7227) );
  AND2_X1 U9069 ( .A1(n8104), .A2(n14688), .ZN(n7228) );
  AND2_X1 U9070 ( .A1(n9226), .A2(n7621), .ZN(n7229) );
  AND2_X1 U9071 ( .A1(n8087), .A2(n8092), .ZN(n7230) );
  AND4_X2 U9072 ( .A1(n7322), .A2(n7718), .A3(n8919), .A4(n8876), .ZN(n7231)
         );
  OAI22_X1 U9073 ( .A1(n14212), .A2(n12956), .B1(n14223), .B2(n12920), .ZN(
        n12918) );
  INV_X1 U9074 ( .A(n14892), .ZN(n8000) );
  INV_X1 U9075 ( .A(n13256), .ZN(n11996) );
  NOR2_X1 U9076 ( .A1(n14750), .A2(n15679), .ZN(n8988) );
  AND2_X1 U9077 ( .A1(n8136), .A2(n13522), .ZN(n7233) );
  AND2_X1 U9078 ( .A1(n13525), .A2(n13509), .ZN(n7234) );
  OR2_X1 U9079 ( .A1(n13039), .A2(n13045), .ZN(n7235) );
  AND2_X1 U9080 ( .A1(n15170), .A2(n12124), .ZN(n7236) );
  AND3_X1 U9081 ( .A1(n12870), .A2(n12869), .A3(n7335), .ZN(n7237) );
  AND2_X1 U9082 ( .A1(n7946), .A2(n7279), .ZN(n7239) );
  AND2_X1 U9083 ( .A1(n14148), .A2(n12490), .ZN(n7240) );
  INV_X1 U9084 ( .A(n7761), .ZN(n7760) );
  OAI21_X1 U9085 ( .B1(n12664), .B2(n7762), .A(n12581), .ZN(n7761) );
  NOR2_X1 U9086 ( .A1(n13122), .A2(n13105), .ZN(n7241) );
  OR2_X1 U9087 ( .A1(n10873), .A2(n15722), .ZN(n7242) );
  NOR2_X1 U9088 ( .A1(n7235), .A2(n14501), .ZN(n7243) );
  OAI21_X1 U9089 ( .B1(n10520), .B2(P2_IR_REG_0__SCAN_IN), .A(n7533), .ZN(
        n12768) );
  INV_X1 U9090 ( .A(n12768), .ZN(n12771) );
  NAND2_X1 U9091 ( .A1(n8254), .A2(n7598), .ZN(n7244) );
  AND2_X1 U9092 ( .A1(n7751), .A2(n7387), .ZN(n7245) );
  AND2_X1 U9093 ( .A1(n9500), .A2(n7598), .ZN(n7246) );
  AND2_X1 U9094 ( .A1(n12872), .A2(n12871), .ZN(n7247) );
  OR2_X1 U9095 ( .A1(n7936), .A2(n14289), .ZN(n7248) );
  NAND2_X2 U9096 ( .A1(n10161), .A2(n10162), .ZN(n14507) );
  NAND2_X1 U9097 ( .A1(n9823), .A2(n8276), .ZN(n7855) );
  NAND3_X1 U9098 ( .A1(n9388), .A2(n8184), .A3(n9398), .ZN(n7249) );
  NAND2_X1 U9099 ( .A1(n9266), .A2(n9265), .ZN(n15989) );
  INV_X1 U9100 ( .A(n15989), .ZN(n7715) );
  INV_X1 U9101 ( .A(n7532), .ZN(n13847) );
  INV_X2 U9103 ( .A(n12848), .ZN(n12795) );
  OR2_X1 U9104 ( .A1(n8201), .A2(n8200), .ZN(n7251) );
  NAND2_X1 U9105 ( .A1(n9661), .A2(n8878), .ZN(n9658) );
  OR2_X1 U9106 ( .A1(n10460), .A2(n10530), .ZN(n7252) );
  INV_X1 U9107 ( .A(n7511), .ZN(n8943) );
  OAI211_X1 U9108 ( .C1(n8899), .C2(P2_DATAO_REG_0__SCAN_IN), .A(n7512), .B(
        SI_0_), .ZN(n7511) );
  INV_X1 U9109 ( .A(n13262), .ZN(n15720) );
  AND2_X1 U9110 ( .A1(n12779), .A2(n12778), .ZN(n7254) );
  NAND2_X1 U9111 ( .A1(n10451), .A2(n10450), .ZN(n10517) );
  NAND2_X1 U9112 ( .A1(n11202), .A2(n11203), .ZN(n7255) );
  NOR2_X1 U9113 ( .A1(n9519), .A2(n9517), .ZN(n7256) );
  INV_X1 U9114 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8498) );
  NAND2_X1 U9115 ( .A1(n9499), .A2(n9498), .ZN(n15092) );
  AND2_X1 U9116 ( .A1(n12888), .A2(n12887), .ZN(n7257) );
  INV_X1 U9117 ( .A(n7834), .ZN(n7833) );
  NAND2_X1 U9118 ( .A1(n7835), .A2(n8316), .ZN(n7834) );
  OR2_X1 U9119 ( .A1(n12009), .A2(n12005), .ZN(n7258) );
  AND2_X1 U9120 ( .A1(n8497), .A2(n8498), .ZN(n8514) );
  OR2_X1 U9121 ( .A1(n10520), .A2(n10398), .ZN(n7259) );
  NAND3_X1 U9122 ( .A1(n9757), .A2(n15204), .A3(n9760), .ZN(n9781) );
  AND2_X1 U9123 ( .A1(n11460), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7260) );
  INV_X1 U9124 ( .A(n12923), .ZN(n7474) );
  NOR2_X1 U9125 ( .A1(n10732), .A2(n8008), .ZN(n7261) );
  NAND2_X1 U9126 ( .A1(n8809), .A2(n12609), .ZN(n13477) );
  AND2_X1 U9127 ( .A1(n12637), .A2(n7748), .ZN(n7262) );
  NOR2_X1 U9128 ( .A1(n13217), .A2(n13483), .ZN(n7263) );
  NOR2_X1 U9129 ( .A1(n13680), .A2(n13244), .ZN(n7264) );
  XNOR2_X1 U9130 ( .A(n15262), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n7265) );
  INV_X1 U9131 ( .A(n8888), .ZN(n7601) );
  INV_X1 U9132 ( .A(n14984), .ZN(n7986) );
  INV_X1 U9133 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15266) );
  NAND2_X1 U9134 ( .A1(n10381), .A2(n10380), .ZN(n10408) );
  AND4_X1 U9135 ( .A1(n10263), .A2(n7391), .A3(n7390), .A4(n7389), .ZN(n7266)
         );
  INV_X1 U9136 ( .A(n11192), .ZN(n12626) );
  OR2_X1 U9137 ( .A1(n14119), .A2(n14341), .ZN(n7267) );
  AND2_X1 U9138 ( .A1(n10753), .A2(n10517), .ZN(n7268) );
  NAND2_X1 U9139 ( .A1(n9379), .A2(n9378), .ZN(n14562) );
  INV_X1 U9140 ( .A(n9478), .ZN(n8255) );
  INV_X1 U9141 ( .A(n9197), .ZN(n8227) );
  OR2_X1 U9142 ( .A1(n13359), .A2(n13358), .ZN(n7269) );
  INV_X1 U9143 ( .A(n9455), .ZN(n8235) );
  INV_X1 U9144 ( .A(n13022), .ZN(n12465) );
  OR2_X1 U9145 ( .A1(n12610), .A2(n12738), .ZN(n7270) );
  INV_X1 U9146 ( .A(n14665), .ZN(n8124) );
  NAND2_X1 U9147 ( .A1(n9293), .A2(n9292), .ZN(n16013) );
  AND2_X1 U9148 ( .A1(n8185), .A2(n7787), .ZN(n7271) );
  NOR2_X1 U9149 ( .A1(n12571), .A2(n12570), .ZN(n7272) );
  NAND2_X1 U9150 ( .A1(n10914), .A2(n10913), .ZN(n12828) );
  AND2_X1 U9151 ( .A1(n7257), .A2(n12890), .ZN(n7273) );
  INV_X1 U9152 ( .A(n12269), .ZN(n15955) );
  NAND2_X1 U9153 ( .A1(n9214), .A2(n9213), .ZN(n12269) );
  AND2_X1 U9154 ( .A1(n12865), .A2(n14013), .ZN(n7274) );
  INV_X1 U9155 ( .A(n11649), .ZN(n7994) );
  OR2_X1 U9156 ( .A1(n13181), .A2(n13486), .ZN(n12609) );
  INV_X1 U9157 ( .A(n12609), .ZN(n7771) );
  AND4_X1 U9158 ( .A1(n8496), .A2(n8495), .A3(n8494), .A4(n8493), .ZN(n12163)
         );
  AND2_X1 U9159 ( .A1(n13078), .A2(n13249), .ZN(n7275) );
  AND2_X1 U9160 ( .A1(n14903), .A2(n12523), .ZN(n7276) );
  INV_X1 U9161 ( .A(n15200), .ZN(n8887) );
  AND2_X1 U9162 ( .A1(n15012), .A2(n7989), .ZN(n7277) );
  INV_X1 U9163 ( .A(n13830), .ZN(n8017) );
  NAND2_X1 U9164 ( .A1(n7681), .A2(n7680), .ZN(n7679) );
  INV_X1 U9165 ( .A(n8195), .ZN(n8194) );
  NAND2_X1 U9166 ( .A1(n14912), .A2(n14925), .ZN(n8195) );
  AND2_X1 U9167 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n7278) );
  NAND2_X1 U9168 ( .A1(n14193), .A2(n14171), .ZN(n7279) );
  AND2_X1 U9169 ( .A1(n12493), .A2(n12492), .ZN(n7280) );
  AND2_X1 U9170 ( .A1(n11305), .A2(n11316), .ZN(n7281) );
  INV_X1 U9171 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7505) );
  INV_X1 U9172 ( .A(n7878), .ZN(n7877) );
  OR2_X1 U9173 ( .A1(n8697), .A2(n7879), .ZN(n7878) );
  INV_X1 U9174 ( .A(n15092), .ZN(n14884) );
  AND2_X1 U9175 ( .A1(n7969), .A2(n7968), .ZN(n7282) );
  INV_X1 U9176 ( .A(n8434), .ZN(n7578) );
  OR2_X1 U9177 ( .A1(n8213), .A2(n12861), .ZN(n7283) );
  INV_X1 U9178 ( .A(n8490), .ZN(n7903) );
  AND2_X1 U9179 ( .A1(n14522), .A2(n8274), .ZN(n7284) );
  AND2_X1 U9180 ( .A1(n14603), .A2(n14602), .ZN(n7285) );
  AND2_X1 U9181 ( .A1(n14560), .A2(n14559), .ZN(n7286) );
  AND2_X1 U9182 ( .A1(n14305), .A2(n12174), .ZN(n13014) );
  AND2_X1 U9183 ( .A1(n13420), .A2(n7971), .ZN(n7287) );
  NOR2_X1 U9184 ( .A1(n9013), .A2(n9012), .ZN(n7288) );
  AND2_X1 U9185 ( .A1(n12880), .A2(n8208), .ZN(n7289) );
  AND2_X1 U9186 ( .A1(n12921), .A2(n8211), .ZN(n7290) );
  INV_X1 U9187 ( .A(n12898), .ZN(n12900) );
  NOR2_X1 U9188 ( .A1(n14954), .A2(n14962), .ZN(n7291) );
  NOR2_X1 U9189 ( .A1(n13717), .A2(n13250), .ZN(n7292) );
  NOR2_X1 U9190 ( .A1(n14461), .A2(n14243), .ZN(n7293) );
  NOR2_X1 U9191 ( .A1(n14437), .A2(n14135), .ZN(n7294) );
  INV_X1 U9192 ( .A(n12488), .ZN(n8067) );
  INV_X1 U9193 ( .A(n12935), .ZN(n8200) );
  AND2_X1 U9194 ( .A1(n8897), .A2(n8222), .ZN(n8221) );
  INV_X1 U9195 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8371) );
  AND2_X1 U9196 ( .A1(n7616), .A2(n7614), .ZN(n7295) );
  NOR2_X1 U9197 ( .A1(n15092), .A2(n14870), .ZN(n7296) );
  NAND2_X1 U9198 ( .A1(n9846), .A2(n9879), .ZN(n9861) );
  NAND3_X1 U9199 ( .A1(n14131), .A2(n14116), .A3(n14115), .ZN(n7297) );
  NAND3_X1 U9200 ( .A1(n7919), .A2(n7238), .A3(n8166), .ZN(n7298) );
  AND2_X1 U9201 ( .A1(n12634), .A2(n12635), .ZN(n12632) );
  INV_X1 U9202 ( .A(n12632), .ZN(n7749) );
  INV_X1 U9203 ( .A(n8269), .ZN(n8160) );
  AND2_X1 U9204 ( .A1(n7449), .A2(n7448), .ZN(n7299) );
  NAND2_X1 U9205 ( .A1(n12728), .A2(n12729), .ZN(n13437) );
  INV_X1 U9206 ( .A(n13437), .ZN(n7769) );
  AND2_X1 U9207 ( .A1(n12843), .A2(n12842), .ZN(n7300) );
  OR2_X1 U9208 ( .A1(n12917), .A2(n12919), .ZN(n7301) );
  INV_X1 U9209 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n10165) );
  AND2_X1 U9210 ( .A1(n8041), .A2(n7441), .ZN(n7302) );
  INV_X1 U9211 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9852) );
  INV_X1 U9212 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9881) );
  INV_X1 U9213 ( .A(n7915), .ZN(n7914) );
  NAND2_X1 U9214 ( .A1(n7916), .A2(n8639), .ZN(n7915) );
  INV_X1 U9215 ( .A(n7999), .ZN(n7998) );
  NAND2_X1 U9216 ( .A1(n8000), .A2(n12523), .ZN(n7999) );
  INV_X1 U9217 ( .A(n7754), .ZN(n7753) );
  NAND2_X1 U9218 ( .A1(n13611), .A2(n7755), .ZN(n7754) );
  NAND2_X1 U9219 ( .A1(n10731), .A2(n10730), .ZN(n8011) );
  INV_X1 U9220 ( .A(n8011), .ZN(n8005) );
  INV_X1 U9221 ( .A(n10264), .ZN(n7675) );
  OAI21_X1 U9222 ( .B1(n12454), .B2(n7936), .A(n7934), .ZN(n7933) );
  NAND2_X1 U9223 ( .A1(n15087), .A2(n14841), .ZN(n7303) );
  AND2_X1 U9224 ( .A1(n8943), .A2(n8972), .ZN(n7304) );
  OR2_X1 U9225 ( .A1(n7853), .A2(n7850), .ZN(n7305) );
  AND2_X1 U9226 ( .A1(n12595), .A2(n7272), .ZN(n7306) );
  INV_X1 U9227 ( .A(n10596), .ZN(n7398) );
  NAND2_X1 U9228 ( .A1(n14212), .A2(n14007), .ZN(n7307) );
  OR2_X1 U9229 ( .A1(n14748), .A2(n10946), .ZN(n7308) );
  NOR2_X1 U9230 ( .A1(n14212), .A2(n14007), .ZN(n7309) );
  AND2_X1 U9231 ( .A1(n14657), .A2(n14656), .ZN(n7310) );
  OR2_X1 U9232 ( .A1(n14119), .A2(n7843), .ZN(n7311) );
  NAND2_X1 U9233 ( .A1(n8254), .A2(n9500), .ZN(n7312) );
  INV_X1 U9234 ( .A(n9111), .ZN(n7626) );
  INV_X1 U9235 ( .A(n8042), .ZN(n8041) );
  NAND2_X1 U9236 ( .A1(n8043), .A2(n13859), .ZN(n8042) );
  INV_X1 U9237 ( .A(n8151), .ZN(n8150) );
  NAND2_X1 U9238 ( .A1(n7258), .A2(n8153), .ZN(n8151) );
  AND2_X1 U9239 ( .A1(n9808), .A2(n9807), .ZN(n7313) );
  INV_X1 U9240 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n15226) );
  INV_X1 U9241 ( .A(n9381), .ZN(n7631) );
  AND2_X1 U9242 ( .A1(n14069), .A2(n14068), .ZN(n7314) );
  AND2_X1 U9243 ( .A1(n12122), .A2(n12123), .ZN(n7315) );
  OR2_X1 U9244 ( .A1(n7257), .A2(n12890), .ZN(n7316) );
  OR2_X1 U9245 ( .A1(n12831), .A2(n12833), .ZN(n7317) );
  OR2_X1 U9246 ( .A1(n12860), .A2(n12862), .ZN(n7318) );
  AND2_X1 U9247 ( .A1(n8284), .A2(n8818), .ZN(n7319) );
  AND2_X1 U9248 ( .A1(n14103), .A2(n14102), .ZN(n7320) );
  AND2_X1 U9249 ( .A1(n7716), .A2(n7715), .ZN(n7321) );
  AND3_X1 U9250 ( .A1(n8918), .A2(n8922), .A3(n8913), .ZN(n7322) );
  NOR2_X1 U9251 ( .A1(n13818), .A2(n12253), .ZN(n7323) );
  NAND2_X1 U9252 ( .A1(n12457), .A2(n12456), .ZN(n14337) );
  AND2_X1 U9253 ( .A1(n8001), .A2(n8221), .ZN(n7324) );
  AND2_X1 U9254 ( .A1(n8810), .A2(n13468), .ZN(n13478) );
  AND2_X1 U9255 ( .A1(n7230), .A2(n7255), .ZN(n7325) );
  NAND2_X1 U9256 ( .A1(n9680), .A2(n7380), .ZN(n7927) );
  INV_X1 U9257 ( .A(n7927), .ZN(n7476) );
  AND2_X1 U9258 ( .A1(n14574), .A2(n14571), .ZN(n7326) );
  AND2_X1 U9259 ( .A1(n12301), .A2(n12299), .ZN(n7327) );
  INV_X1 U9260 ( .A(n11955), .ZN(n8034) );
  OR2_X1 U9261 ( .A1(n8212), .A2(n12832), .ZN(n7328) );
  OR2_X1 U9262 ( .A1(n12898), .A2(n8210), .ZN(n7329) );
  INV_X1 U9263 ( .A(n14147), .ZN(n7942) );
  OR2_X1 U9264 ( .A1(n9087), .A2(n9085), .ZN(n7330) );
  OR2_X1 U9265 ( .A1(n8255), .A2(n9477), .ZN(n7331) );
  OR2_X1 U9266 ( .A1(n12900), .A2(n12899), .ZN(n7332) );
  AND2_X1 U9267 ( .A1(n14967), .A2(n12510), .ZN(n7333) );
  OR2_X1 U9268 ( .A1(n9294), .A2(n9296), .ZN(n7334) );
  OR2_X1 U9269 ( .A1(n8209), .A2(n7247), .ZN(n7335) );
  AND2_X1 U9270 ( .A1(n8219), .A2(n7641), .ZN(n7336) );
  NAND2_X1 U9271 ( .A1(n7706), .A2(SI_3_), .ZN(n9000) );
  AND2_X1 U9272 ( .A1(n8249), .A2(n7625), .ZN(n7337) );
  NOR2_X1 U9273 ( .A1(n8227), .A2(n9196), .ZN(n8228) );
  INV_X1 U9274 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n10172) );
  INV_X1 U9275 ( .A(n9501), .ZN(n7598) );
  INV_X1 U9276 ( .A(n8220), .ZN(n8219) );
  NAND2_X1 U9277 ( .A1(n8221), .A2(n8879), .ZN(n8220) );
  INV_X1 U9278 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7375) );
  NAND2_X1 U9279 ( .A1(n15129), .A2(n14573), .ZN(n7338) );
  INV_X1 U9280 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8913) );
  OR2_X1 U9281 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n7339) );
  INV_X1 U9282 ( .A(n7896), .ZN(n7895) );
  NAND2_X1 U9283 ( .A1(n7749), .A2(n8426), .ZN(n7896) );
  OR2_X1 U9284 ( .A1(n7768), .A2(n7765), .ZN(n7340) );
  INV_X1 U9285 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9925) );
  INV_X1 U9286 ( .A(n9056), .ZN(n9582) );
  AND2_X1 U9287 ( .A1(n13935), .A2(n13826), .ZN(n13984) );
  INV_X2 U9288 ( .A(n10460), .ZN(n12064) );
  INV_X1 U9289 ( .A(n14396), .ZN(n7838) );
  NAND2_X1 U9290 ( .A1(n7890), .A2(n7889), .ZN(n13636) );
  NAND2_X1 U9291 ( .A1(n12962), .A2(n12961), .ZN(n14334) );
  INV_X1 U9292 ( .A(n14334), .ZN(n7842) );
  AND2_X1 U9293 ( .A1(n8144), .A2(n8148), .ZN(n7341) );
  INV_X1 U9294 ( .A(n13030), .ZN(n7526) );
  INV_X1 U9295 ( .A(n11454), .ZN(n7674) );
  AND2_X1 U9296 ( .A1(n12676), .A2(n12677), .ZN(n13665) );
  INV_X1 U9297 ( .A(n13665), .ZN(n7395) );
  AND2_X1 U9298 ( .A1(n9328), .A2(SI_18_), .ZN(n7342) );
  INV_X1 U9299 ( .A(n11463), .ZN(n15617) );
  INV_X1 U9300 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7389) );
  NOR2_X1 U9301 ( .A1(n13288), .A2(n13289), .ZN(n7343) );
  AND2_X1 U9302 ( .A1(n13588), .A2(n7914), .ZN(n7344) );
  INV_X1 U9303 ( .A(n7795), .ZN(n7792) );
  NAND2_X1 U9304 ( .A1(n8168), .A2(SI_18_), .ZN(n7795) );
  INV_X1 U9305 ( .A(n8182), .ZN(n8181) );
  NOR2_X1 U9306 ( .A1(n9374), .A2(SI_19_), .ZN(n8182) );
  OR2_X1 U9307 ( .A1(n8177), .A2(n8175), .ZN(n7345) );
  INV_X1 U9308 ( .A(n7786), .ZN(n7784) );
  INV_X1 U9309 ( .A(n7797), .ZN(n7796) );
  AND2_X1 U9310 ( .A1(n11645), .A2(n7992), .ZN(n7346) );
  OR2_X1 U9311 ( .A1(n13066), .A2(n13613), .ZN(n7347) );
  INV_X1 U9312 ( .A(n9388), .ZN(n8179) );
  INV_X1 U9313 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8782) );
  INV_X1 U9314 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9682) );
  INV_X1 U9315 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7390) );
  NAND2_X1 U9317 ( .A1(n10647), .A2(n9815), .ZN(n7865) );
  AND2_X1 U9318 ( .A1(n15663), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7348) );
  INV_X1 U9319 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7665) );
  INV_X1 U9320 ( .A(n15917), .ZN(n7721) );
  NAND2_X1 U9321 ( .A1(n7613), .A2(n11487), .ZN(n11543) );
  OR2_X1 U9322 ( .A1(n11259), .A2(n11258), .ZN(n7349) );
  NAND2_X1 U9323 ( .A1(n7497), .A2(n8833), .ZN(n8827) );
  OR2_X1 U9324 ( .A1(n13269), .A2(n11677), .ZN(n7350) );
  NOR2_X1 U9325 ( .A1(n11114), .A2(n11113), .ZN(n7351) );
  AND2_X1 U9326 ( .A1(n12017), .A2(n7716), .ZN(n7352) );
  INV_X1 U9327 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7745) );
  AND2_X1 U9328 ( .A1(n8154), .A2(n8159), .ZN(n7353) );
  INV_X1 U9329 ( .A(SI_18_), .ZN(n11833) );
  AND2_X1 U9330 ( .A1(n8009), .A2(n7261), .ZN(n7354) );
  AND2_X1 U9331 ( .A1(n10943), .A2(n7230), .ZN(n7355) );
  AND2_X1 U9332 ( .A1(n10943), .A2(n8092), .ZN(n7356) );
  AND2_X1 U9333 ( .A1(n11017), .A2(n11016), .ZN(n7357) );
  AND2_X1 U9334 ( .A1(n7590), .A2(n7589), .ZN(n7358) );
  NAND2_X1 U9335 ( .A1(n10603), .A2(n9734), .ZN(n8086) );
  INV_X1 U9336 ( .A(n10146), .ZN(n10604) );
  INV_X1 U9337 ( .A(n15870), .ZN(n7905) );
  NAND2_X1 U9338 ( .A1(n10174), .A2(n10175), .ZN(n14487) );
  INV_X1 U9339 ( .A(n10799), .ZN(n8090) );
  NAND2_X1 U9340 ( .A1(n13414), .A2(n13384), .ZN(n7359) );
  AND2_X1 U9341 ( .A1(n7956), .A2(n7955), .ZN(n7360) );
  INV_X1 U9342 ( .A(n10024), .ZN(n7666) );
  INV_X1 U9343 ( .A(n9348), .ZN(n14825) );
  INV_X1 U9344 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7743) );
  INV_X1 U9345 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7742) );
  INV_X1 U9346 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8167) );
  INV_X1 U9347 ( .A(SI_7_), .ZN(n7413) );
  INV_X1 U9348 ( .A(SI_9_), .ZN(n7427) );
  INV_X1 U9349 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n7952) );
  INV_X1 U9350 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7737) );
  INV_X1 U9351 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7741) );
  NAND3_X1 U9352 ( .A1(n15326), .A2(n15675), .A3(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7809) );
  OAI21_X1 U9353 ( .B1(n9020), .B2(n9019), .A(n9042), .ZN(n10549) );
  NAND2_X1 U9354 ( .A1(n12285), .A2(n12284), .ZN(n12283) );
  INV_X1 U9355 ( .A(n14996), .ZN(n7799) );
  OAI21_X1 U9356 ( .B1(n8899), .B2(n7363), .A(n7362), .ZN(n8901) );
  INV_X1 U9357 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7363) );
  NAND2_X1 U9358 ( .A1(n7304), .A2(n8942), .ZN(n8971) );
  INV_X1 U9359 ( .A(n8971), .ZN(n8973) );
  NOR2_X1 U9360 ( .A1(n15086), .A2(n15799), .ZN(n7366) );
  AND2_X2 U9361 ( .A1(n14922), .A2(n12522), .ZN(n14905) );
  AOI21_X1 U9362 ( .B1(n7369), .B2(n10958), .A(n14289), .ZN(n10959) );
  NAND2_X1 U9363 ( .A1(n10830), .A2(n12993), .ZN(n7369) );
  NAND2_X1 U9364 ( .A1(n14433), .A2(n15974), .ZN(n7377) );
  NAND2_X2 U9365 ( .A1(n7379), .A2(n7378), .ZN(n9856) );
  NAND2_X1 U9366 ( .A1(n7381), .A2(n10835), .ZN(n11005) );
  NAND2_X1 U9367 ( .A1(n10884), .A2(n10834), .ZN(n7381) );
  NAND2_X1 U9368 ( .A1(n12054), .A2(n12873), .ZN(n7383) );
  NAND2_X1 U9369 ( .A1(n7702), .A2(n12100), .ZN(n7384) );
  NAND2_X2 U9370 ( .A1(n14239), .A2(n12360), .ZN(n14221) );
  NAND2_X1 U9371 ( .A1(n14241), .A2(n14240), .ZN(n14239) );
  AND4_X2 U9372 ( .A1(n10391), .A2(n10393), .A3(n10392), .A4(n10394), .ZN(
        n10812) );
  NAND2_X4 U9373 ( .A1(n8788), .A2(n8787), .ZN(n10126) );
  NAND3_X1 U9374 ( .A1(n10263), .A2(n7871), .A3(n7392), .ZN(n7964) );
  OR2_X1 U9375 ( .A1(n13264), .A2(n7398), .ZN(n11170) );
  NAND2_X1 U9376 ( .A1(n7675), .A2(n7400), .ZN(n7399) );
  NOR2_X1 U9377 ( .A1(n8554), .A2(n7392), .ZN(n7400) );
  INV_X1 U9378 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n15272) );
  OAI21_X1 U9379 ( .B1(n15463), .B2(n15464), .A(n7743), .ZN(n7406) );
  INV_X1 U9380 ( .A(n7408), .ZN(n15471) );
  NAND2_X1 U9381 ( .A1(n7409), .A2(n7408), .ZN(n7744) );
  OR2_X1 U9382 ( .A1(n15473), .A2(n15472), .ZN(n7408) );
  NAND2_X1 U9383 ( .A1(n7410), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7409) );
  NAND2_X1 U9384 ( .A1(n15473), .A2(n15472), .ZN(n7410) );
  XNOR2_X1 U9385 ( .A(n9097), .B(n7411), .ZN(n10726) );
  INV_X1 U9386 ( .A(n9080), .ZN(n7414) );
  NAND2_X1 U9387 ( .A1(n7420), .A2(n9287), .ZN(n9308) );
  NAND2_X1 U9388 ( .A1(n9284), .A2(n9283), .ZN(n7420) );
  INV_X1 U9389 ( .A(n9125), .ZN(n7425) );
  NAND2_X1 U9390 ( .A1(n7428), .A2(n7427), .ZN(n7426) );
  INV_X1 U9391 ( .A(n7429), .ZN(n7428) );
  NAND2_X1 U9392 ( .A1(n7429), .A2(SI_9_), .ZN(n9133) );
  NAND2_X1 U9393 ( .A1(n7695), .A2(n7693), .ZN(n7429) );
  NAND3_X1 U9394 ( .A1(n9332), .A2(n9347), .A3(n12959), .ZN(n12325) );
  NAND2_X1 U9395 ( .A1(n7430), .A2(n9595), .ZN(n9336) );
  NAND2_X1 U9396 ( .A1(n7436), .A2(n7435), .ZN(n13952) );
  NOR2_X1 U9397 ( .A1(n10519), .A2(n10518), .ZN(n10752) );
  NAND2_X1 U9398 ( .A1(n10527), .A2(n10526), .ZN(n7438) );
  NAND3_X1 U9399 ( .A1(n7447), .A2(n7476), .A3(n9681), .ZN(n10382) );
  OAI21_X2 U9400 ( .B1(n13899), .B2(n13898), .A(n13841), .ZN(n13844) );
  INV_X1 U9401 ( .A(n12953), .ZN(n7448) );
  NAND2_X1 U9402 ( .A1(n12955), .A2(n12954), .ZN(n7449) );
  NAND3_X1 U9403 ( .A1(n7451), .A2(n7450), .A3(n7332), .ZN(n12906) );
  NAND3_X1 U9404 ( .A1(n7454), .A2(n7453), .A3(n7452), .ZN(n7451) );
  INV_X1 U9405 ( .A(n7489), .ZN(n7452) );
  INV_X1 U9406 ( .A(n7487), .ZN(n7453) );
  NAND3_X1 U9407 ( .A1(n7462), .A2(n7318), .A3(n7461), .ZN(n7460) );
  OR2_X1 U9408 ( .A1(n12854), .A2(n12853), .ZN(n7461) );
  NAND2_X1 U9409 ( .A1(n7463), .A2(n7534), .ZN(n7462) );
  NAND2_X1 U9410 ( .A1(n12854), .A2(n12853), .ZN(n7463) );
  AOI21_X1 U9411 ( .B1(n12825), .B2(n12824), .A(n12822), .ZN(n12823) );
  OAI21_X1 U9412 ( .B1(n7546), .B2(n7465), .A(n12816), .ZN(n7464) );
  AND2_X1 U9413 ( .A1(n12809), .A2(n8203), .ZN(n7465) );
  OAI22_X1 U9414 ( .A1(n7237), .A2(n7466), .B1(n12881), .B2(n7469), .ZN(n12886) );
  NOR2_X1 U9415 ( .A1(n7468), .A2(n12881), .ZN(n7467) );
  INV_X1 U9416 ( .A(n12880), .ZN(n7469) );
  OAI22_X1 U9417 ( .A1(n7470), .A2(n7471), .B1(n7474), .B2(n12922), .ZN(n12928) );
  INV_X1 U9418 ( .A(n8211), .ZN(n7473) );
  NAND3_X1 U9419 ( .A1(n10169), .A2(n7476), .A3(n7475), .ZN(n10174) );
  NAND2_X2 U9420 ( .A1(n10520), .A2(n10395), .ZN(n12960) );
  NAND2_X2 U9421 ( .A1(n10179), .A2(n14487), .ZN(n10520) );
  NAND2_X1 U9422 ( .A1(n7510), .A2(n12910), .ZN(n12915) );
  OAI21_X1 U9423 ( .B1(n12803), .B2(n12802), .A(n12801), .ZN(n12809) );
  OAI21_X1 U9424 ( .B1(n12789), .B2(n12788), .A(n12787), .ZN(n12798) );
  OAI211_X1 U9425 ( .C1(n14083), .C2(n15406), .A(n7480), .B(n14082), .ZN(
        P2_U3233) );
  NAND2_X1 U9426 ( .A1(n14081), .A2(n15419), .ZN(n7480) );
  AOI21_X1 U9427 ( .B1(n11701), .B2(P2_REG1_REG_13__SCAN_IN), .A(n11695), .ZN(
        n11698) );
  NAND2_X1 U9428 ( .A1(n8019), .A2(n7323), .ZN(n8021) );
  NAND2_X1 U9429 ( .A1(n10442), .A2(n10441), .ZN(n10443) );
  NOR2_X1 U9430 ( .A1(n10918), .A2(n10917), .ZN(n11110) );
  NOR2_X1 U9431 ( .A1(n10492), .A2(n10493), .ZN(n10491) );
  INV_X2 U9432 ( .A(n12776), .ZN(n10440) );
  NAND2_X1 U9433 ( .A1(n12781), .A2(n12776), .ZN(n12764) );
  NAND2_X2 U9434 ( .A1(n7259), .A2(n7848), .ZN(n12776) );
  NAND2_X1 U9435 ( .A1(n8214), .A2(n8216), .ZN(n12854) );
  NAND2_X1 U9436 ( .A1(n12868), .A2(n12867), .ZN(n7530) );
  OAI21_X1 U9437 ( .B1(n8197), .B2(n12937), .A(n12940), .ZN(n12955) );
  OAI21_X1 U9438 ( .B1(n7527), .B2(n12823), .A(n7328), .ZN(n12839) );
  NAND2_X1 U9439 ( .A1(n7481), .A2(n12771), .ZN(n12773) );
  NAND2_X1 U9440 ( .A1(n10157), .A2(n9685), .ZN(n10158) );
  NOR2_X1 U9441 ( .A1(n10160), .A2(n10159), .ZN(n10161) );
  OAI21_X2 U9442 ( .B1(n11350), .B2(n11349), .A(n11348), .ZN(n11577) );
  INV_X1 U9443 ( .A(n13182), .ZN(n8135) );
  NAND2_X1 U9444 ( .A1(n8158), .A2(n10876), .ZN(n8157) );
  OR2_X1 U9445 ( .A1(n8904), .A2(n7511), .ZN(n7488) );
  OAI22_X1 U9446 ( .A1(n13818), .A2(n8024), .B1(n13816), .B2(n13817), .ZN(
        n8023) );
  NAND2_X1 U9447 ( .A1(n10171), .A2(n8054), .ZN(n8055) );
  NAND2_X1 U9448 ( .A1(n13976), .A2(n13975), .ZN(n13846) );
  XNOR2_X1 U9449 ( .A(n15749), .B(n10445), .ZN(n10451) );
  NAND2_X1 U9450 ( .A1(n7528), .A2(n12932), .ZN(n12934) );
  NAND2_X1 U9451 ( .A1(n13924), .A2(n13925), .ZN(n13923) );
  NAND2_X1 U9452 ( .A1(n12096), .A2(n12097), .ZN(n12213) );
  NOR2_X1 U9453 ( .A1(n10491), .A2(n10444), .ZN(n10453) );
  INV_X1 U9454 ( .A(n8171), .ZN(n8170) );
  OAI21_X1 U9455 ( .B1(n12886), .B2(n12885), .A(n7316), .ZN(n7487) );
  NAND3_X1 U9456 ( .A1(n7488), .A2(n8906), .A3(n8905), .ZN(n8976) );
  NAND3_X1 U9457 ( .A1(n8006), .A2(n13923), .A3(n8004), .ZN(n8003) );
  OAI22_X1 U9458 ( .A1(n12786), .A2(n7254), .B1(n12785), .B2(n12784), .ZN(
        n12788) );
  NAND2_X1 U9459 ( .A1(n12781), .A2(n14024), .ZN(n12779) );
  INV_X1 U9460 ( .A(n12837), .ZN(n7535) );
  INV_X1 U9461 ( .A(n12852), .ZN(n7534) );
  NAND2_X1 U9462 ( .A1(n12906), .A2(n12907), .ZN(n12905) );
  NAND2_X1 U9464 ( .A1(n12095), .A2(n12094), .ZN(n12096) );
  AOI21_X1 U9465 ( .B1(n12886), .B2(n12885), .A(n12884), .ZN(n7489) );
  OR2_X1 U9466 ( .A1(n10451), .A2(n10450), .ZN(n7531) );
  NAND2_X1 U9467 ( .A1(n7531), .A2(n10517), .ZN(n10452) );
  NAND2_X1 U9468 ( .A1(n8127), .A2(n8913), .ZN(n9290) );
  NAND2_X2 U9469 ( .A1(n9727), .A2(n8262), .ZN(n10603) );
  NOR2_X1 U9470 ( .A1(n9710), .A2(n9719), .ZN(n10143) );
  XNOR2_X1 U9471 ( .A(n8923), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9705) );
  NAND2_X1 U9472 ( .A1(n12129), .A2(n12128), .ZN(n12265) );
  NOR2_X1 U9473 ( .A1(n12121), .A2(n7315), .ZN(n12129) );
  NAND2_X1 U9474 ( .A1(n7490), .A2(n9737), .ZN(n10943) );
  NAND3_X1 U9475 ( .A1(n7492), .A2(n14267), .A3(n14099), .ZN(n7705) );
  NAND2_X1 U9476 ( .A1(n14098), .A2(n14097), .ZN(n7492) );
  NAND2_X1 U9477 ( .A1(n7939), .A2(n7940), .ZN(n14150) );
  NAND2_X1 U9478 ( .A1(n7523), .A2(n7521), .ZN(n14353) );
  NAND2_X1 U9479 ( .A1(n14434), .A2(n15970), .ZN(n14357) );
  NAND2_X1 U9480 ( .A1(n9308), .A2(n9307), .ZN(n7495) );
  NAND2_X1 U9481 ( .A1(n7787), .A2(n9122), .ZN(n7697) );
  OAI21_X1 U9482 ( .B1(n9288), .B2(n9925), .A(n7509), .ZN(n9080) );
  INV_X1 U9483 ( .A(n7794), .ZN(n7793) );
  OAI22_X1 U9484 ( .A1(n12798), .A2(n12797), .B1(n12800), .B2(n12799), .ZN(
        n12803) );
  NAND2_X1 U9485 ( .A1(n8822), .A2(n11328), .ZN(n7497) );
  NAND2_X1 U9486 ( .A1(n8826), .A2(n8825), .ZN(n10615) );
  NAND2_X1 U9487 ( .A1(n12300), .A2(n7327), .ZN(n13064) );
  OR2_X1 U9488 ( .A1(n13087), .A2(n13086), .ZN(n13088) );
  NAND4_X1 U9489 ( .A1(n7919), .A2(n8166), .A3(n7918), .A4(n7925), .ZN(n7923)
         );
  NAND2_X1 U9490 ( .A1(n9047), .A2(n9079), .ZN(n10565) );
  AND2_X2 U9491 ( .A1(n11932), .A2(n8095), .ZN(n12121) );
  OR2_X1 U9492 ( .A1(n10521), .A2(n10449), .ZN(n7499) );
  NAND2_X1 U9493 ( .A1(n7254), .A2(n12786), .ZN(n12787) );
  NAND3_X1 U9494 ( .A1(n7507), .A2(n12769), .A3(n12770), .ZN(n12775) );
  OAI21_X1 U9495 ( .B1(n8978), .B2(n8173), .A(n9004), .ZN(n8171) );
  NAND2_X1 U9496 ( .A1(n13366), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n13386) );
  AOI21_X1 U9497 ( .B1(n13428), .B2(n15912), .A(n13429), .ZN(n8869) );
  INV_X2 U9498 ( .A(n8796), .ZN(n15715) );
  NAND2_X1 U9499 ( .A1(n7340), .A2(n7549), .ZN(n12750) );
  OR2_X2 U9500 ( .A1(n8816), .A2(n7339), .ZN(n8369) );
  AOI21_X1 U9501 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(n15299), .A(n15466), .ZN(
        n15473) );
  NAND2_X1 U9502 ( .A1(n15443), .A2(n7740), .ZN(n15275) );
  NOR2_X1 U9503 ( .A1(n15501), .A2(n15500), .ZN(n15499) );
  AOI22_X1 U9504 ( .A1(n12336), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n12335), 
        .B2(n15372), .ZN(n10535) );
  INV_X1 U9505 ( .A(n12847), .ZN(n8218) );
  INV_X1 U9506 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7689) );
  NAND2_X1 U9507 ( .A1(n12981), .A2(n12767), .ZN(n12770) );
  NAND3_X1 U9508 ( .A1(n9020), .A2(n8187), .A3(n9019), .ZN(n7701) );
  NAND2_X1 U9509 ( .A1(n7520), .A2(n7519), .ZN(n12840) );
  NAND2_X1 U9510 ( .A1(n7518), .A2(n7517), .ZN(n12869) );
  NAND2_X1 U9511 ( .A1(n8169), .A2(n8170), .ZN(n9016) );
  NAND2_X1 U9512 ( .A1(n12905), .A2(n12904), .ZN(n7510) );
  NAND2_X1 U9513 ( .A1(n8899), .A2(n10405), .ZN(n7512) );
  NAND2_X1 U9514 ( .A1(n9001), .A2(n9000), .ZN(n9005) );
  NOR2_X1 U9515 ( .A1(n13404), .A2(n7513), .ZN(n13411) );
  AND2_X1 U9516 ( .A1(n13406), .A2(n13405), .ZN(n7513) );
  INV_X4 U9517 ( .A(n10129), .ZN(n13408) );
  NOR2_X1 U9518 ( .A1(n14067), .A2(n7314), .ZN(n14071) );
  NAND2_X1 U9519 ( .A1(n14261), .A2(n12347), .ZN(n14241) );
  INV_X1 U9520 ( .A(n12794), .ZN(n15764) );
  NAND2_X1 U9521 ( .A1(n8883), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8884) );
  NAND2_X1 U9522 ( .A1(n8120), .A2(n14623), .ZN(n7553) );
  NAND2_X1 U9523 ( .A1(n7524), .A2(n8082), .ZN(n11215) );
  NAND3_X1 U9524 ( .A1(n10943), .A2(n8093), .A3(n7325), .ZN(n7524) );
  NAND2_X1 U9525 ( .A1(n13064), .A2(n13063), .ZN(n13231) );
  NAND2_X1 U9526 ( .A1(n10874), .A2(n11238), .ZN(n11045) );
  NAND2_X1 U9527 ( .A1(n8156), .A2(n8160), .ZN(n8155) );
  NAND2_X1 U9528 ( .A1(n12085), .A2(n12297), .ZN(n12300) );
  INV_X1 U9529 ( .A(n13174), .ZN(n7545) );
  NAND2_X1 U9530 ( .A1(n7710), .A2(n7709), .ZN(n13232) );
  AOI21_X1 U9531 ( .B1(n7712), .B2(n8782), .A(n8554), .ZN(n7711) );
  OAI21_X1 U9532 ( .B1(n13193), .B2(n13085), .A(n13084), .ZN(n13087) );
  OAI21_X1 U9533 ( .B1(n12825), .B2(n12824), .A(n7317), .ZN(n7527) );
  NAND3_X1 U9534 ( .A1(n12841), .A2(n12840), .A3(n8215), .ZN(n8214) );
  INV_X1 U9535 ( .A(n12866), .ZN(n7529) );
  NAND2_X1 U9536 ( .A1(n12927), .A2(n12926), .ZN(n7528) );
  NAND2_X1 U9537 ( .A1(n12774), .A2(n12775), .ZN(n12785) );
  NAND2_X1 U9538 ( .A1(n7530), .A2(n7529), .ZN(n12870) );
  NAND2_X1 U9539 ( .A1(n13952), .A2(n10540), .ZN(n13924) );
  NAND2_X1 U9540 ( .A1(n12213), .A2(n12212), .ZN(n12214) );
  OAI21_X1 U9541 ( .B1(n10171), .B2(n11039), .A(P2_IR_REG_27__SCAN_IN), .ZN(
        n7538) );
  AOI21_X1 U9542 ( .B1(n12934), .B2(n7251), .A(n8198), .ZN(n8197) );
  NAND2_X1 U9543 ( .A1(n7536), .A2(n7535), .ZN(n12841) );
  NAND2_X1 U9544 ( .A1(n12839), .A2(n12838), .ZN(n7536) );
  NAND2_X1 U9545 ( .A1(n7539), .A2(n8167), .ZN(n7807) );
  NAND3_X1 U9546 ( .A1(n7689), .A2(n15674), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7539) );
  OAI21_X1 U9547 ( .B1(n14130), .B2(n8074), .A(n8072), .ZN(n14095) );
  OAI21_X1 U9548 ( .B1(n7698), .B2(n7697), .A(n7696), .ZN(n7695) );
  INV_X1 U9549 ( .A(n8174), .ZN(n9442) );
  NAND2_X1 U9550 ( .A1(n8943), .A2(n8942), .ZN(n8902) );
  AND2_X2 U9551 ( .A1(n11015), .A2(n11034), .ZN(n11030) );
  AOI22_X1 U9552 ( .A1(n12336), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n12335), 
        .B2(n15361), .ZN(n10524) );
  NOR2_X4 U9553 ( .A1(n14159), .A2(n14363), .ZN(n14140) );
  NOR2_X1 U9554 ( .A1(n11103), .A2(n12794), .ZN(n10961) );
  NAND2_X1 U9555 ( .A1(n9701), .A2(n8271), .ZN(n9704) );
  XNOR2_X1 U9556 ( .A(n7553), .B(n7552), .ZN(n14628) );
  INV_X1 U9557 ( .A(n9702), .ZN(n7541) );
  NOR2_X1 U9558 ( .A1(n10144), .A2(n9719), .ZN(n10428) );
  NAND2_X2 U9559 ( .A1(n14706), .A2(n14590), .ZN(n14640) );
  OAI21_X2 U9560 ( .B1(n13095), .B2(n13094), .A(n13182), .ZN(n13129) );
  NAND2_X1 U9561 ( .A1(n8157), .A2(n8155), .ZN(n11225) );
  NAND2_X1 U9562 ( .A1(n13232), .A2(n7347), .ZN(n13167) );
  INV_X1 U9563 ( .A(n13231), .ZN(n7710) );
  NAND2_X1 U9564 ( .A1(n12749), .A2(n10612), .ZN(n10614) );
  INV_X1 U9565 ( .A(n7712), .ZN(n8781) );
  NAND2_X1 U9566 ( .A1(n8202), .A2(n12817), .ZN(n7546) );
  NAND2_X1 U9567 ( .A1(n8809), .A2(n7770), .ZN(n13469) );
  NAND3_X1 U9568 ( .A1(n7550), .A2(n8207), .A3(n13058), .ZN(P2_U3328) );
  NAND2_X1 U9569 ( .A1(n7809), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7808) );
  INV_X1 U9570 ( .A(n9078), .ZN(n8188) );
  NAND2_X1 U9571 ( .A1(n8029), .A2(n8027), .ZN(n12095) );
  NAND2_X1 U9572 ( .A1(n13990), .A2(n13863), .ZN(n13887) );
  INV_X1 U9573 ( .A(n11123), .ZN(n7708) );
  NAND2_X1 U9574 ( .A1(n7708), .A2(n12959), .ZN(n7707) );
  NAND2_X1 U9575 ( .A1(n8928), .A2(n8921), .ZN(n8931) );
  NAND2_X1 U9576 ( .A1(n13359), .A2(n13358), .ZN(n7555) );
  OR2_X1 U9577 ( .A1(n11462), .A2(n15601), .ZN(n7556) );
  NAND2_X1 U9578 ( .A1(n8596), .A2(n7560), .ZN(n7559) );
  INV_X1 U9579 ( .A(n8312), .ZN(n7574) );
  NAND2_X1 U9580 ( .A1(n7570), .A2(n7568), .ZN(n8484) );
  NAND2_X1 U9581 ( .A1(n8312), .A2(n7571), .ZN(n7570) );
  NAND2_X1 U9582 ( .A1(n8753), .A2(n7583), .ZN(n7579) );
  NAND2_X1 U9583 ( .A1(n7579), .A2(n7580), .ZN(n12543) );
  NAND2_X1 U9584 ( .A1(n8753), .A2(n8366), .ZN(n7582) );
  NAND2_X1 U9585 ( .A1(n8350), .A2(n7358), .ZN(n7586) );
  NAND2_X1 U9586 ( .A1(n7586), .A2(n7587), .ZN(n8356) );
  NAND3_X1 U9587 ( .A1(n7590), .A2(n8699), .A3(n7589), .ZN(n7588) );
  NAND2_X1 U9588 ( .A1(n7595), .A2(n7596), .ZN(n8251) );
  NAND2_X1 U9589 ( .A1(n8253), .A2(n7597), .ZN(n7595) );
  NAND2_X1 U9590 ( .A1(n7605), .A2(n7604), .ZN(n8225) );
  AOI21_X1 U9591 ( .B1(n7608), .B2(n9174), .A(n8228), .ZN(n7604) );
  NAND2_X1 U9592 ( .A1(n9156), .A2(n7606), .ZN(n7605) );
  NAND2_X1 U9593 ( .A1(n7609), .A2(n7607), .ZN(n7606) );
  INV_X1 U9594 ( .A(n7608), .ZN(n7607) );
  NAND2_X1 U9595 ( .A1(n9174), .A2(n9155), .ZN(n7609) );
  OR2_X1 U9596 ( .A1(n9225), .A2(n7229), .ZN(n7619) );
  NAND2_X1 U9597 ( .A1(n9225), .A2(n7617), .ZN(n7616) );
  NAND2_X1 U9598 ( .A1(n8248), .A2(n7337), .ZN(n7622) );
  NAND2_X1 U9599 ( .A1(n7622), .A2(n7623), .ZN(n8240) );
  NAND2_X1 U9600 ( .A1(n7627), .A2(n7630), .ZN(n9410) );
  NAND3_X1 U9601 ( .A1(n9369), .A2(n7628), .A3(n9368), .ZN(n7627) );
  INV_X1 U9602 ( .A(n9656), .ZN(n7640) );
  NAND2_X1 U9603 ( .A1(n7640), .A2(n7336), .ZN(n7642) );
  OR2_X2 U9604 ( .A1(n9656), .A2(n8220), .ZN(n8883) );
  NAND2_X1 U9605 ( .A1(n8190), .A2(n7645), .ZN(n7646) );
  INV_X1 U9606 ( .A(n7646), .ZN(n14866) );
  INV_X1 U9607 ( .A(n9038), .ZN(n7650) );
  AND4_X2 U9608 ( .A1(n8907), .A2(n7651), .A3(n7652), .A4(n7653), .ZN(n9105)
         );
  NAND2_X1 U9609 ( .A1(n8909), .A2(n7672), .ZN(n9021) );
  MUX2_X1 U9610 ( .A(n7677), .B(P3_IR_REG_31__SCAN_IN), .S(n7871), .Z(n7676)
         );
  NOR2_X2 U9611 ( .A1(n13310), .A2(n7682), .ZN(n13328) );
  NOR2_X1 U9612 ( .A1(n15628), .A2(n11401), .ZN(n15649) );
  NAND3_X1 U9613 ( .A1(n8187), .A2(n7694), .A3(n9020), .ZN(n7693) );
  INV_X1 U9614 ( .A(n8185), .ZN(n7698) );
  INV_X1 U9615 ( .A(n9122), .ZN(n7700) );
  NAND2_X1 U9616 ( .A1(n11979), .A2(n7703), .ZN(n7702) );
  NAND2_X1 U9617 ( .A1(n11979), .A2(n11978), .ZN(n12054) );
  OAI21_X1 U9618 ( .B1(n7706), .B2(SI_3_), .A(n9000), .ZN(n8977) );
  MUX2_X1 U9619 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n9311), .Z(n7706) );
  NAND3_X1 U9620 ( .A1(n8166), .A2(n8497), .A3(n8498), .ZN(n8627) );
  NAND2_X2 U9621 ( .A1(n8883), .A2(n8896), .ZN(n12758) );
  NAND2_X1 U9622 ( .A1(n12017), .A2(n7321), .ZN(n7717) );
  INV_X1 U9623 ( .A(n7717), .ZN(n15058) );
  NAND4_X1 U9624 ( .A1(n7231), .A2(n9105), .A3(n7719), .A4(n8001), .ZN(n9656)
         );
  NOR2_X1 U9625 ( .A1(n14906), .A2(n14895), .ZN(n14894) );
  NAND2_X1 U9626 ( .A1(n7729), .A2(n7727), .ZN(n15455) );
  INV_X1 U9627 ( .A(n7728), .ZN(n7727) );
  NOR2_X1 U9628 ( .A1(n15450), .A2(n15277), .ZN(n15281) );
  INV_X1 U9629 ( .A(n15277), .ZN(n7732) );
  AOI21_X1 U9630 ( .B1(n7262), .B2(n7750), .A(n7747), .ZN(n7746) );
  NAND2_X1 U9631 ( .A1(n13469), .A2(n12606), .ZN(n8811) );
  OAI21_X1 U9632 ( .B1(n14886), .B2(n7774), .A(n7773), .ZN(n14845) );
  NAND2_X1 U9633 ( .A1(n7777), .A2(n7775), .ZN(n12528) );
  NAND2_X1 U9634 ( .A1(n14886), .A2(n7778), .ZN(n7777) );
  AOI21_X1 U9635 ( .B1(n9329), .B2(n7796), .A(n7792), .ZN(n7794) );
  NAND2_X1 U9636 ( .A1(n8168), .A2(n9328), .ZN(n7797) );
  NAND3_X1 U9637 ( .A1(n7800), .A2(n7798), .A3(n7338), .ZN(n14948) );
  OAI21_X2 U9638 ( .B1(n9138), .B2(n7803), .A(n7801), .ZN(n9199) );
  NAND3_X1 U9639 ( .A1(n9136), .A2(n9164), .A3(n7804), .ZN(n7802) );
  INV_X2 U9640 ( .A(n8899), .ZN(n9311) );
  NAND2_X1 U9641 ( .A1(n8745), .A2(n8363), .ZN(n7811) );
  NAND3_X1 U9642 ( .A1(n12726), .A2(n7270), .A3(n7812), .ZN(n12734) );
  NAND2_X1 U9643 ( .A1(n7817), .A2(n7815), .ZN(n8309) );
  INV_X1 U9644 ( .A(n7816), .ZN(n7815) );
  NAND2_X1 U9645 ( .A1(n8378), .A2(n7818), .ZN(n7817) );
  INV_X1 U9646 ( .A(n8331), .ZN(n7823) );
  NOR2_X2 U9647 ( .A1(n14321), .A2(n14320), .ZN(n14324) );
  NOR2_X4 U9648 ( .A1(n11142), .A2(n12844), .ZN(n11322) );
  NAND2_X2 U9649 ( .A1(n11030), .A2(n7837), .ZN(n11142) );
  NOR2_X2 U9650 ( .A1(n14247), .A2(n14456), .ZN(n14228) );
  NOR2_X2 U9651 ( .A1(n14293), .A2(n14461), .ZN(n7839) );
  NAND2_X1 U9652 ( .A1(n14140), .A2(n7840), .ZN(n14089) );
  NAND2_X1 U9653 ( .A1(n10520), .A2(n10404), .ZN(n10521) );
  INV_X1 U9654 ( .A(n8275), .ZN(n7856) );
  NAND2_X1 U9655 ( .A1(n10647), .A2(n7860), .ZN(n7859) );
  NAND2_X1 U9656 ( .A1(n7859), .A2(n7857), .ZN(n9820) );
  NAND2_X1 U9657 ( .A1(n9666), .A2(n7868), .ZN(n7869) );
  INV_X2 U9658 ( .A(n8959), .ZN(n9349) );
  NAND2_X2 U9659 ( .A1(n9666), .A2(n12758), .ZN(n8959) );
  AND3_X2 U9660 ( .A1(n8950), .A2(n8949), .A3(n7869), .ZN(n9699) );
  AND2_X1 U9661 ( .A1(n8374), .A2(n7870), .ZN(n8267) );
  NAND3_X1 U9662 ( .A1(n13812), .A2(n8297), .A3(P3_REG2_REG_1__SCAN_IN), .ZN(
        n7870) );
  OAI21_X2 U9663 ( .B1(n8686), .B2(n7874), .A(n7873), .ZN(n13506) );
  OAI21_X1 U9664 ( .B1(n8542), .B2(n7888), .A(n7885), .ZN(n8592) );
  OAI21_X1 U9665 ( .B1(n11193), .B2(n7896), .A(n7893), .ZN(n11268) );
  AND2_X1 U9666 ( .A1(n8456), .A2(n7894), .ZN(n7893) );
  NAND2_X1 U9667 ( .A1(n7895), .A2(n12626), .ZN(n7894) );
  INV_X1 U9668 ( .A(n11993), .ZN(n7909) );
  AND2_X1 U9669 ( .A1(n8490), .A2(n7907), .ZN(n7906) );
  INV_X1 U9670 ( .A(n12163), .ZN(n7907) );
  NAND3_X1 U9671 ( .A1(n8371), .A2(n7911), .A3(n8370), .ZN(n7910) );
  AND2_X1 U9672 ( .A1(n8283), .A2(n8498), .ZN(n7925) );
  INV_X1 U9673 ( .A(n7923), .ZN(n8834) );
  NOR2_X2 U9674 ( .A1(n11153), .A2(n15836), .ZN(n11152) );
  NOR2_X2 U9675 ( .A1(n12127), .A2(n11659), .ZN(n12017) );
  NOR2_X1 U9676 ( .A1(n9856), .A2(n9677), .ZN(n10331) );
  NAND2_X1 U9677 ( .A1(n14117), .A2(n12454), .ZN(n14099) );
  OAI211_X1 U9678 ( .C1(n14117), .C2(n7248), .A(n7931), .B(n7929), .ZN(n7928)
         );
  NAND2_X1 U9679 ( .A1(n14117), .A2(n7930), .ZN(n7929) );
  OAI21_X2 U9680 ( .B1(n13366), .B2(n7953), .A(n7951), .ZN(n13415) );
  NAND3_X1 U9681 ( .A1(n7966), .A2(n7965), .A3(n13332), .ZN(n13364) );
  NAND2_X1 U9682 ( .A1(n11151), .A2(n7313), .ZN(n11374) );
  NAND2_X1 U9683 ( .A1(n7975), .A2(n7974), .ZN(n9803) );
  NAND3_X1 U9684 ( .A1(n10651), .A2(n10652), .A3(n9801), .ZN(n7974) );
  NAND2_X1 U9685 ( .A1(n10651), .A2(n10652), .ZN(n7978) );
  INV_X2 U9686 ( .A(n9104), .ZN(n9596) );
  NAND2_X1 U9687 ( .A1(n8980), .A2(n9001), .ZN(n9870) );
  NAND2_X1 U9688 ( .A1(n15045), .A2(n7987), .ZN(n7990) );
  INV_X1 U9689 ( .A(n7990), .ZN(n15029) );
  OAI22_X1 U9690 ( .A1(n11558), .A2(n7991), .B1(n7992), .B2(n7236), .ZN(n12016) );
  OAI21_X2 U9691 ( .B1(n14905), .B2(n7999), .A(n7996), .ZN(n14886) );
  NAND2_X1 U9692 ( .A1(n9661), .A2(n7324), .ZN(n8894) );
  NOR2_X1 U9693 ( .A1(n10724), .A2(n10555), .ZN(n8010) );
  OAI21_X1 U9694 ( .B1(n8005), .B2(n7261), .A(n8003), .ZN(n10918) );
  INV_X1 U9695 ( .A(n10724), .ZN(n8006) );
  NAND2_X1 U9696 ( .A1(n13923), .A2(n10556), .ZN(n10725) );
  INV_X1 U9697 ( .A(n12214), .ZN(n8019) );
  INV_X1 U9698 ( .A(n8035), .ZN(n11567) );
  NAND2_X1 U9699 ( .A1(n10818), .A2(n8044), .ZN(n8045) );
  NAND3_X1 U9700 ( .A1(n8045), .A2(n8047), .A3(n12996), .ZN(n10822) );
  NAND4_X2 U9701 ( .A1(n10416), .A2(n10415), .A3(n10414), .A4(n10413), .ZN(
        n14024) );
  NAND2_X1 U9702 ( .A1(n14024), .A2(n12848), .ZN(n12783) );
  NAND2_X1 U9703 ( .A1(n11607), .A2(n8051), .ZN(n8048) );
  NAND2_X1 U9704 ( .A1(n8048), .A2(n8049), .ZN(n12071) );
  NAND2_X1 U9705 ( .A1(n14282), .A2(n8057), .ZN(n8056) );
  INV_X1 U9706 ( .A(n8061), .ZN(n14185) );
  NAND2_X1 U9707 ( .A1(n12486), .A2(n12485), .ZN(n14219) );
  NAND2_X1 U9708 ( .A1(n12196), .A2(n8071), .ZN(n12480) );
  NAND2_X1 U9709 ( .A1(n12480), .A2(n8068), .ZN(n12482) );
  OAI21_X1 U9710 ( .B1(n14130), .B2(n12492), .A(n12493), .ZN(n14112) );
  NAND2_X1 U9711 ( .A1(n11017), .A2(n8081), .ZN(n11018) );
  INV_X1 U9712 ( .A(n9727), .ZN(n10601) );
  AND2_X1 U9713 ( .A1(n10143), .A2(n10142), .ZN(n10144) );
  NAND2_X2 U9714 ( .A1(n8086), .A2(n8094), .ZN(n8093) );
  INV_X1 U9715 ( .A(n11933), .ZN(n8100) );
  NAND2_X1 U9716 ( .A1(n14640), .A2(n7228), .ZN(n8102) );
  NAND2_X2 U9717 ( .A1(n8102), .A2(n8101), .ZN(n14680) );
  NAND2_X1 U9718 ( .A1(n14716), .A2(n8109), .ZN(n8106) );
  NAND2_X1 U9719 ( .A1(n8106), .A2(n8107), .ZN(n14697) );
  NAND2_X1 U9720 ( .A1(n14725), .A2(n8114), .ZN(n8113) );
  OAI211_X1 U9721 ( .C1(n14725), .C2(n8118), .A(n8115), .B(n8113), .ZN(n14670)
         );
  NAND2_X1 U9722 ( .A1(n14725), .A2(n14726), .ZN(n8120) );
  NAND2_X2 U9723 ( .A1(n12271), .A2(n12270), .ZN(n14518) );
  NAND2_X1 U9724 ( .A1(n14698), .A2(n7326), .ZN(n14671) );
  NAND2_X2 U9725 ( .A1(n14567), .A2(n14566), .ZN(n14698) );
  INV_X1 U9726 ( .A(n8126), .ZN(n10044) );
  NAND2_X1 U9727 ( .A1(n10043), .A2(n8126), .ZN(n9718) );
  NOR2_X2 U9728 ( .A1(n9290), .A2(n8920), .ZN(n8928) );
  INV_X1 U9729 ( .A(n9262), .ZN(n8127) );
  NAND2_X2 U9730 ( .A1(n9825), .A2(n11665), .ZN(n9702) );
  NAND2_X1 U9731 ( .A1(n10710), .A2(n8128), .ZN(n10623) );
  OR2_X1 U9732 ( .A1(n10622), .A2(n8129), .ZN(n8128) );
  NAND2_X1 U9733 ( .A1(n10622), .A2(n8129), .ZN(n10710) );
  NOR2_X1 U9734 ( .A1(n10708), .A2(n8130), .ZN(n8129) );
  AND2_X1 U9735 ( .A1(n10621), .A2(n13262), .ZN(n8130) );
  INV_X1 U9736 ( .A(n13129), .ZN(n8136) );
  NAND2_X1 U9737 ( .A1(n8131), .A2(n8133), .ZN(n13154) );
  NAND2_X1 U9738 ( .A1(n13129), .A2(n8132), .ZN(n8131) );
  INV_X1 U9739 ( .A(n8135), .ZN(n8132) );
  NAND2_X1 U9740 ( .A1(n8137), .A2(n8138), .ZN(n13111) );
  NAND2_X1 U9741 ( .A1(n13219), .A2(n8139), .ZN(n8137) );
  NAND2_X1 U9742 ( .A1(n11578), .A2(n8145), .ZN(n8141) );
  NAND2_X1 U9743 ( .A1(n8141), .A2(n8142), .ZN(n12084) );
  OR2_X1 U9744 ( .A1(n13070), .A2(n13251), .ZN(n8165) );
  AND2_X2 U9745 ( .A1(n8279), .A2(n8598), .ZN(n8166) );
  INV_X1 U9746 ( .A(n9000), .ZN(n8173) );
  OR2_X2 U9747 ( .A1(n8976), .A2(n8975), .ZN(n8172) );
  NAND3_X1 U9748 ( .A1(n8172), .A2(n9000), .A3(n8974), .ZN(n8169) );
  INV_X1 U9749 ( .A(n9375), .ZN(n8184) );
  NAND2_X1 U9750 ( .A1(n15108), .A2(n8191), .ZN(n8190) );
  NAND2_X1 U9751 ( .A1(n9684), .A2(n8268), .ZN(n8196) );
  INV_X1 U9752 ( .A(n12933), .ZN(n8201) );
  INV_X1 U9753 ( .A(n8204), .ZN(n8202) );
  INV_X1 U9754 ( .A(n12874), .ZN(n8209) );
  INV_X1 U9755 ( .A(n12899), .ZN(n8210) );
  NAND2_X1 U9756 ( .A1(n8217), .A2(n8218), .ZN(n8215) );
  INV_X1 U9757 ( .A(n7300), .ZN(n8217) );
  NAND2_X1 U9758 ( .A1(n7300), .A2(n12847), .ZN(n8216) );
  NAND2_X1 U9759 ( .A1(n8223), .A2(n8224), .ZN(n9318) );
  NAND3_X1 U9760 ( .A1(n9273), .A2(n7334), .A3(n9272), .ZN(n8223) );
  NAND2_X1 U9761 ( .A1(n8225), .A2(n8226), .ZN(n9225) );
  NAND2_X1 U9762 ( .A1(n8229), .A2(n8230), .ZN(n9269) );
  NAND2_X1 U9763 ( .A1(n9246), .A2(n8232), .ZN(n8229) );
  NAND2_X1 U9764 ( .A1(n9429), .A2(n8238), .ZN(n8236) );
  OAI21_X1 U9765 ( .B1(n9429), .B2(n8237), .A(n8238), .ZN(n9454) );
  NAND2_X1 U9766 ( .A1(n8236), .A2(n8234), .ZN(n9453) );
  NAND2_X1 U9767 ( .A1(n8240), .A2(n8239), .ZN(n9156) );
  NAND3_X1 U9768 ( .A1(n9323), .A2(n9322), .A3(n8244), .ZN(n8246) );
  NAND3_X1 U9769 ( .A1(n9069), .A2(n7330), .A3(n9068), .ZN(n8248) );
  NAND2_X1 U9770 ( .A1(n8251), .A2(n8252), .ZN(n9540) );
  NAND3_X1 U9771 ( .A1(n9458), .A2(n7331), .A3(n9457), .ZN(n8253) );
  NOR2_X1 U9772 ( .A1(n15568), .A2(n15567), .ZN(n15566) );
  MUX2_X1 U9773 ( .A(n14433), .B(P2_REG1_REG_28__SCAN_IN), .S(n14355), .Z(
        P2_U3527) );
  AND2_X1 U9774 ( .A1(n11519), .A2(n11318), .ZN(n15928) );
  NAND2_X1 U9775 ( .A1(n8272), .A2(n15091), .ZN(n15180) );
  INV_X1 U9776 ( .A(n10390), .ZN(n14482) );
  INV_X1 U9777 ( .A(n15090), .ZN(n15091) );
  INV_X1 U9778 ( .A(n14474), .ZN(n14476) );
  NAND2_X2 U9779 ( .A1(n14612), .A2(n14611), .ZN(n14725) );
  INV_X1 U9780 ( .A(n12612), .ZN(n10751) );
  NAND2_X2 U9781 ( .A1(n12612), .A2(n12754), .ZN(n12738) );
  INV_X1 U9782 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9879) );
  AND2_X1 U9783 ( .A1(n9709), .A2(n9708), .ZN(n9710) );
  NAND2_X1 U9784 ( .A1(n10529), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n10413) );
  NAND2_X1 U9785 ( .A1(n10376), .A2(n9682), .ZN(n10381) );
  OR2_X1 U9786 ( .A1(n10158), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n9686) );
  NAND2_X1 U9787 ( .A1(n14275), .A2(n12761), .ZN(n14129) );
  NAND4_X1 U9788 ( .A1(n8386), .A2(n8385), .A3(n8384), .A4(n8383), .ZN(n13264)
         );
  NAND2_X2 U9789 ( .A1(n9822), .A2(n9821), .ZN(n11160) );
  AOI21_X1 U9790 ( .B1(n12750), .B2(n12749), .A(n12748), .ZN(n12757) );
  OR2_X1 U9791 ( .A1(n10685), .A2(n9348), .ZN(n10764) );
  NAND2_X1 U9792 ( .A1(n9613), .A2(n9612), .ZN(n9648) );
  MUX2_X1 U9793 ( .A(n9611), .B(n9612), .S(n9610), .Z(n9655) );
  OAI22_X2 U9794 ( .A1(n13566), .A2(n8675), .B1(n13580), .B2(n13143), .ZN(
        n13547) );
  NAND2_X1 U9795 ( .A1(n9656), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9657) );
  AOI21_X2 U9796 ( .B1(n13448), .B2(n13454), .A(n8812), .ZN(n13443) );
  OR2_X1 U9797 ( .A1(n13430), .A2(n13738), .ZN(n8257) );
  OR2_X1 U9798 ( .A1(n13430), .A2(n13794), .ZN(n8258) );
  INV_X2 U9799 ( .A(n15735), .ZN(n13670) );
  INV_X1 U9800 ( .A(n12503), .ZN(n15046) );
  NOR2_X1 U9801 ( .A1(n10599), .A2(n10600), .ZN(n8262) );
  NOR2_X1 U9802 ( .A1(n11554), .A2(n11553), .ZN(n8263) );
  OR2_X1 U9803 ( .A1(n12520), .A2(n15137), .ZN(n8264) );
  AND2_X2 U9804 ( .A1(n9671), .A2(n9889), .ZN(P1_U4016) );
  AND2_X1 U9805 ( .A1(n12534), .A2(n15035), .ZN(n15020) );
  INV_X1 U9806 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8554) );
  INV_X1 U9807 ( .A(n9808), .ZN(n9828) );
  AND2_X1 U9808 ( .A1(n9683), .A2(n9682), .ZN(n8268) );
  INV_X1 U9809 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9685) );
  AND2_X1 U9810 ( .A1(n11223), .A2(n11226), .ZN(n8269) );
  INV_X1 U9811 ( .A(n12527), .ZN(n12515) );
  OR2_X1 U9812 ( .A1(n15153), .A2(n16030), .ZN(n8270) );
  AND4_X1 U9813 ( .A1(n8719), .A2(n8718), .A3(n8717), .A4(n8716), .ZN(n13522)
         );
  OR2_X1 U9814 ( .A1(n9699), .A2(n14583), .ZN(n8271) );
  AND2_X1 U9815 ( .A1(n12980), .A2(n12979), .ZN(n8273) );
  NAND2_X1 U9816 ( .A1(n13047), .A2(n13046), .ZN(n13048) );
  OR2_X1 U9817 ( .A1(n10763), .A2(n10762), .ZN(n16023) );
  INV_X2 U9818 ( .A(n16023), .ZN(n15961) );
  OR2_X1 U9819 ( .A1(n10065), .A2(n10762), .ZN(n16021) );
  AND2_X1 U9820 ( .A1(n15836), .A2(n10997), .ZN(n8275) );
  OR2_X1 U9821 ( .A1(n15836), .A2(n10997), .ZN(n8276) );
  INV_X1 U9822 ( .A(n9039), .ZN(n9040) );
  INV_X1 U9823 ( .A(n12916), .ZN(n12917) );
  INV_X1 U9824 ( .A(n12925), .ZN(n12926) );
  INV_X1 U9825 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n9672) );
  XNOR2_X1 U9826 ( .A(n9348), .B(n15217), .ZN(n9577) );
  NAND2_X1 U9827 ( .A1(n12602), .A2(n12612), .ZN(n10613) );
  INV_X1 U9828 ( .A(n13009), .ZN(n11616) );
  NAND2_X1 U9829 ( .A1(n9577), .A2(n9824), .ZN(n8933) );
  OAI21_X1 U9830 ( .B1(n10615), .B2(n10614), .A(n10613), .ZN(n10616) );
  INV_X1 U9831 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n11913) );
  OR4_X1 U9832 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n9767) );
  INV_X1 U9833 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8918) );
  AND2_X1 U9834 ( .A1(n13083), .A2(n13146), .ZN(n13084) );
  INV_X1 U9835 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n11814) );
  INV_X1 U9836 ( .A(n13513), .ZN(n13505) );
  NAND2_X1 U9837 ( .A1(n8606), .A2(n12583), .ZN(n13606) );
  NAND2_X1 U9838 ( .A1(n12602), .A2(n13407), .ZN(n10617) );
  INV_X1 U9839 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10921) );
  OR3_X1 U9840 ( .A1(n12423), .A2(n13907), .A3(n13994), .ZN(n12435) );
  OR2_X1 U9841 ( .A1(n12381), .A2(n13977), .ZN(n12393) );
  OR2_X1 U9842 ( .A1(n9031), .A2(n9951), .ZN(n8936) );
  INV_X1 U9843 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8878) );
  INV_X1 U9844 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8914) );
  INV_X1 U9845 ( .A(n12304), .ZN(n12301) );
  OR2_X1 U9846 ( .A1(n8714), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8725) );
  OR2_X1 U9847 ( .A1(n13062), .A2(n13627), .ZN(n13063) );
  AND2_X1 U9848 ( .A1(n8632), .A2(n11901), .ZN(n8650) );
  OAI22_X1 U9849 ( .A1(n13456), .A2(n15721), .B1(n13422), .B2(n12565), .ZN(
        n8793) );
  AND2_X1 U9850 ( .A1(n11954), .A2(n11953), .ZN(n11955) );
  NAND2_X1 U9851 ( .A1(n12403), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n12423) );
  INV_X1 U9852 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n12326) );
  INV_X1 U9853 ( .A(n14148), .ZN(n14154) );
  INV_X1 U9854 ( .A(n13016), .ZN(n14258) );
  NAND2_X1 U9855 ( .A1(n15950), .A2(n7526), .ZN(n10476) );
  INV_X1 U9856 ( .A(n14349), .ZN(n14350) );
  NAND2_X1 U9857 ( .A1(n10408), .A2(n14073), .ZN(n13053) );
  INV_X1 U9858 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n10170) );
  INV_X1 U9859 ( .A(n14632), .ZN(n14522) );
  INV_X1 U9860 ( .A(n9432), .ZN(n9433) );
  NAND2_X1 U9861 ( .A1(n15081), .A2(n14737), .ZN(n12526) );
  NAND2_X1 U9862 ( .A1(n14981), .A2(n12509), .ZN(n14969) );
  OR2_X1 U9863 ( .A1(n16013), .A2(n16028), .ZN(n12518) );
  INV_X1 U9864 ( .A(n10970), .ZN(n9804) );
  INV_X1 U9865 ( .A(n14584), .ZN(n9741) );
  INV_X1 U9866 ( .A(n8988), .ZN(n9624) );
  INV_X1 U9867 ( .A(n9705), .ZN(n9706) );
  OR2_X1 U9868 ( .A1(n9192), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9193) );
  INV_X1 U9869 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n15237) );
  INV_X1 U9870 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15248) );
  OR2_X1 U9871 ( .A1(n12738), .A2(n10124), .ZN(n10125) );
  AOI21_X1 U9872 ( .B1(n7398), .B2(n13109), .A(n10619), .ZN(n10622) );
  NOR2_X1 U9873 ( .A1(n8544), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8570) );
  NAND2_X1 U9874 ( .A1(n10351), .A2(n10624), .ZN(n13225) );
  OR2_X1 U9875 ( .A1(n10353), .A2(n10352), .ZN(n10356) );
  AND2_X1 U9876 ( .A1(n8831), .A2(n8830), .ZN(n8832) );
  INV_X1 U9877 ( .A(n15663), .ZN(n15593) );
  OR2_X1 U9878 ( .A1(n13713), .A2(n13580), .ZN(n12701) );
  INV_X1 U9879 ( .A(n12583), .ZN(n13624) );
  OR2_X1 U9880 ( .A1(n8442), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8458) );
  NOR2_X1 U9881 ( .A1(n12746), .A2(n15935), .ZN(n10354) );
  OR2_X1 U9882 ( .A1(n10615), .A2(n10588), .ZN(n8860) );
  INV_X1 U9883 ( .A(n8858), .ZN(n13430) );
  OR2_X1 U9884 ( .A1(n7221), .A2(n11828), .ZN(n8723) );
  OR2_X1 U9885 ( .A1(n8852), .A2(n8850), .ZN(n8848) );
  INV_X1 U9886 ( .A(n11269), .ZN(n12637) );
  INV_X1 U9887 ( .A(n12754), .ZN(n8850) );
  OR2_X1 U9888 ( .A1(n8865), .A2(n8864), .ZN(n10350) );
  OR2_X1 U9889 ( .A1(n8827), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8829) );
  INV_X1 U9890 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8370) );
  AND2_X1 U9891 ( .A1(n8337), .A2(n8336), .ZN(n8607) );
  NOR2_X1 U9892 ( .A1(n8530), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n8565) );
  INV_X1 U9893 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13968) );
  OR2_X1 U9894 ( .A1(n11521), .A2(n11520), .ZN(n11972) );
  INV_X1 U9895 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11569) );
  OR2_X1 U9896 ( .A1(n12327), .A2(n12326), .ZN(n12340) );
  NAND2_X1 U9897 ( .A1(n10528), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n10400) );
  INV_X1 U9898 ( .A(n10190), .ZN(n10192) );
  AND2_X1 U9899 ( .A1(n10192), .A2(n10180), .ZN(n10187) );
  OAI21_X1 U9900 ( .B1(n14507), .B2(n14073), .A(n10419), .ZN(n14267) );
  INV_X1 U9901 ( .A(n15970), .ZN(n14355) );
  XNOR2_X1 U9902 ( .A(n14386), .B(n14007), .ZN(n14213) );
  INV_X1 U9903 ( .A(n14242), .ZN(n14283) );
  INV_X1 U9904 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9688) );
  INV_X1 U9905 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n13234) );
  INV_X1 U9906 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n11039) );
  INV_X1 U9907 ( .A(n14743), .ZN(n11485) );
  AOI21_X1 U9908 ( .B1(n10061), .B2(n14615), .A(n9714), .ZN(n9715) );
  INV_X1 U9909 ( .A(n15978), .ZN(n14520) );
  OR2_X1 U9910 ( .A1(n14545), .A2(n14544), .ZN(n14546) );
  INV_X1 U9911 ( .A(n9646), .ZN(n9647) );
  AND2_X1 U9912 ( .A1(n9370), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9382) );
  INV_X1 U9913 ( .A(n15153), .ZN(n15023) );
  INV_X1 U9914 ( .A(n12237), .ZN(n12236) );
  INV_X1 U9915 ( .A(n14740), .ZN(n12124) );
  INV_X1 U9916 ( .A(n11542), .ZN(n11553) );
  INV_X1 U9917 ( .A(n9873), .ZN(n9888) );
  XNOR2_X1 U9918 ( .A(n15145), .B(n14719), .ZN(n14997) );
  INV_X1 U9919 ( .A(n15954), .ZN(n16014) );
  NAND2_X1 U9920 ( .A1(n15796), .A2(n9348), .ZN(n10063) );
  NAND2_X1 U9921 ( .A1(n9649), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8923) );
  NOR2_X1 U9922 ( .A1(n15235), .A2(n15234), .ZN(n15292) );
  OAI21_X1 U9923 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n15239), .A(n15238), .ZN(
        n15261) );
  AND2_X1 U9924 ( .A1(n10348), .A2(n10355), .ZN(n13221) );
  AND4_X1 U9925 ( .A1(n8763), .A2(n8762), .A3(n8761), .A4(n8760), .ZN(n13467)
         );
  AND4_X1 U9926 ( .A1(n8684), .A2(n8683), .A3(n8682), .A4(n8681), .ZN(n13568)
         );
  AND4_X1 U9927 ( .A1(n8620), .A2(n8619), .A3(n8618), .A4(n8617), .ZN(n13591)
         );
  NAND2_X1 U9928 ( .A1(n8833), .A2(n8832), .ZN(n10336) );
  NOR2_X1 U9929 ( .A1(n11669), .A2(n11668), .ZN(n11672) );
  INV_X1 U9930 ( .A(n15583), .ZN(n15667) );
  INV_X1 U9931 ( .A(n13653), .ZN(n13667) );
  INV_X1 U9932 ( .A(n15727), .ZN(n13648) );
  AND2_X1 U9933 ( .A1(n8855), .A2(n8854), .ZN(n8856) );
  INV_X1 U9934 ( .A(n15935), .ZN(n15891) );
  NAND2_X1 U9935 ( .A1(n8815), .A2(n8848), .ZN(n15937) );
  AND2_X1 U9936 ( .A1(n11183), .A2(n8850), .ZN(n15931) );
  OR2_X1 U9937 ( .A1(n15937), .A2(n15931), .ZN(n15912) );
  XNOR2_X1 U9938 ( .A(n8785), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12754) );
  INV_X1 U9939 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8644) );
  OR2_X1 U9940 ( .A1(n10666), .A2(n15339), .ZN(n10475) );
  AND2_X1 U9941 ( .A1(n12441), .A2(n12440), .ZN(n14135) );
  INV_X1 U9942 ( .A(n12425), .ZN(n12458) );
  NAND2_X1 U9943 ( .A1(n10192), .A2(n10191), .ZN(n14074) );
  INV_X1 U9944 ( .A(n15406), .ZN(n15423) );
  AND2_X1 U9945 ( .A1(n10456), .A2(n10179), .ZN(n14262) );
  INV_X1 U9946 ( .A(n14254), .ZN(n14315) );
  INV_X1 U9947 ( .A(n14417), .ZN(n14422) );
  INV_X1 U9948 ( .A(n15339), .ZN(n10665) );
  INV_X1 U9949 ( .A(n15963), .ZN(n15845) );
  INV_X1 U9950 ( .A(n15778), .ZN(n15812) );
  AND2_X1 U9951 ( .A1(n15333), .A2(n10385), .ZN(n10840) );
  AND2_X1 U9952 ( .A1(n9868), .A2(n9867), .ZN(n15361) );
  INV_X1 U9953 ( .A(n9699), .ZN(n10697) );
  AND2_X1 U9954 ( .A1(n14691), .A2(n15033), .ZN(n16029) );
  NAND2_X1 U9955 ( .A1(n9779), .A2(n15035), .ZN(n14731) );
  NAND2_X1 U9956 ( .A1(n9648), .A2(n9647), .ZN(n9654) );
  AND4_X1 U9957 ( .A1(n9407), .A2(n9406), .A3(n9405), .A4(n9404), .ZN(n14927)
         );
  AND2_X1 U9958 ( .A1(n9895), .A2(n9893), .ZN(n9949) );
  INV_X1 U9959 ( .A(n14819), .ZN(n15434) );
  AND2_X1 U9960 ( .A1(n9949), .A2(n9948), .ZN(n14819) );
  OR2_X1 U9961 ( .A1(n11647), .A2(n7346), .ZN(n15173) );
  OR2_X1 U9962 ( .A1(n15020), .A2(n9837), .ZN(n15681) );
  INV_X1 U9963 ( .A(n15680), .ZN(n15061) );
  INV_X1 U9964 ( .A(n15020), .ZN(n15055) );
  OR2_X1 U9965 ( .A1(n9832), .A2(n9788), .ZN(n10065) );
  AND2_X1 U9966 ( .A1(n9827), .A2(n9826), .ZN(n16016) );
  NAND2_X1 U9967 ( .A1(n10764), .A2(n10987), .ZN(n16019) );
  AND2_X1 U9968 ( .A1(n9889), .A2(n9665), .ZN(n9873) );
  XNOR2_X1 U9969 ( .A(n8898), .B(n8897), .ZN(n9666) );
  AND2_X1 U9970 ( .A1(n10135), .A2(n10134), .ZN(n15663) );
  INV_X1 U9971 ( .A(n12316), .ZN(n15934) );
  INV_X1 U9972 ( .A(n13221), .ZN(n13229) );
  INV_X1 U9973 ( .A(n13206), .ZN(n13242) );
  INV_X1 U9974 ( .A(n13591), .ZN(n13626) );
  INV_X1 U9975 ( .A(n11172), .ZN(n13261) );
  INV_X1 U9976 ( .A(n15602), .ZN(n15657) );
  OR2_X1 U9977 ( .A1(n10136), .A2(n10128), .ZN(n15671) );
  INV_X1 U9978 ( .A(n13412), .ZN(n15659) );
  AND2_X1 U9979 ( .A1(n13594), .A2(n13593), .ZN(n13721) );
  NAND2_X1 U9980 ( .A1(n15735), .A2(n15734), .ZN(n13653) );
  NAND2_X2 U9981 ( .A1(n10594), .A2(n15727), .ZN(n15735) );
  NAND2_X1 U9982 ( .A1(n15940), .A2(n15891), .ZN(n13738) );
  INV_X1 U9983 ( .A(n13217), .ZN(n13757) );
  AND2_X2 U9984 ( .A1(n8868), .A2(n10355), .ZN(n15944) );
  NAND2_X1 U9985 ( .A1(n8827), .A2(n13796), .ZN(n9938) );
  AND2_X1 U9986 ( .A1(n10335), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13796) );
  INV_X1 U9987 ( .A(SI_23_), .ZN(n11723) );
  INV_X1 U9988 ( .A(SI_17_), .ZN(n11840) );
  INV_X1 U9989 ( .A(SI_12_), .ZN(n11850) );
  INV_X1 U9990 ( .A(n15601), .ZN(n11461) );
  AND2_X1 U9991 ( .A1(n10190), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15341) );
  NAND2_X1 U9992 ( .A1(n13957), .A2(n14242), .ZN(n13997) );
  INV_X1 U9993 ( .A(n14001), .ZN(n13974) );
  OR2_X1 U9994 ( .A1(n10475), .A2(n10458), .ZN(n14003) );
  INV_X1 U9995 ( .A(n12958), .ZN(n14085) );
  INV_X1 U9996 ( .A(n14188), .ZN(n14006) );
  OR2_X1 U9997 ( .A1(n12068), .A2(n12067), .ZN(n14010) );
  INV_X1 U9998 ( .A(n15341), .ZN(n15427) );
  AND2_X1 U9999 ( .A1(n12188), .A2(n13918), .ZN(n14419) );
  INV_X1 U10000 ( .A(n14275), .ZN(n15817) );
  AND2_X1 U10001 ( .A1(n10667), .A2(n14318), .ZN(n15829) );
  AND2_X1 U10002 ( .A1(n14129), .A2(n10886), .ZN(n14254) );
  NAND2_X1 U10003 ( .A1(n15970), .A2(n15845), .ZN(n14417) );
  AND2_X2 U10004 ( .A1(n10840), .A2(n10665), .ZN(n15970) );
  INV_X1 U10005 ( .A(n14193), .ZN(n14452) );
  INV_X1 U10006 ( .A(n12865), .ZN(n12154) );
  INV_X1 U10007 ( .A(n15974), .ZN(n15971) );
  AND2_X2 U10008 ( .A1(n10840), .A2(n15339), .ZN(n15974) );
  OR2_X1 U10009 ( .A1(n15337), .A2(n15335), .ZN(n15336) );
  INV_X1 U10010 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14481) );
  INV_X1 U10011 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n14504) );
  INV_X1 U10012 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10333) );
  INV_X1 U10013 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10039) );
  NAND2_X1 U10014 ( .A1(n10395), .A2(P2_U3088), .ZN(n14503) );
  INV_X1 U10015 ( .A(n11550), .ZN(n11544) );
  INV_X1 U10016 ( .A(n11377), .ZN(n11339) );
  INV_X1 U10017 ( .A(n14562), .ZN(n15137) );
  OR2_X1 U10018 ( .A1(n9778), .A2(n9776), .ZN(n14733) );
  INV_X1 U10019 ( .A(n14927), .ZN(n14962) );
  INV_X1 U10020 ( .A(n14791), .ZN(n15440) );
  INV_X1 U10021 ( .A(n14828), .ZN(n15067) );
  OR2_X1 U10022 ( .A1(n15036), .A2(n16016), .ZN(n15064) );
  AND3_X1 U10023 ( .A1(n11658), .A2(n11657), .A3(n11656), .ZN(n15175) );
  OR2_X1 U10024 ( .A1(n15036), .A2(n10685), .ZN(n14988) );
  INV_X1 U10025 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11281) );
  INV_X1 U10026 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10334) );
  INV_X1 U10027 ( .A(n14025), .ZN(P2_U3947) );
  OR4_X1 U10028 ( .A1(n9842), .A2(n9841), .A3(n9840), .A4(n9839), .ZN(P1_U3285) );
  INV_X1 U10029 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8857) );
  INV_X1 U10030 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8284) );
  NAND2_X1 U10031 ( .A1(n8287), .A2(n8285), .ZN(n13801) );
  AND2_X2 U10032 ( .A1(n13808), .A2(n13812), .ZN(n8521) );
  NAND2_X1 U10033 ( .A1(n12552), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8301) );
  NAND2_X1 U10034 ( .A1(n8520), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8300) );
  NOR2_X1 U10035 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8427) );
  INV_X1 U10036 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U10037 ( .A1(n8427), .A2(n8428), .ZN(n8442) );
  NOR2_X1 U10038 ( .A1(n8458), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8476) );
  NAND2_X1 U10039 ( .A1(n8491), .A2(n11787), .ZN(n8522) );
  NAND2_X1 U10040 ( .A1(n8570), .A2(n11915), .ZN(n8585) );
  INV_X1 U10041 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n11816) );
  NAND2_X1 U10042 ( .A1(n11816), .A2(n13234), .ZN(n8290) );
  INV_X1 U10043 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n11901) );
  INV_X1 U10044 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n11801) );
  NAND2_X1 U10045 ( .A1(n8650), .A2(n11801), .ZN(n8668) );
  NAND2_X1 U10046 ( .A1(n11913), .A2(n8669), .ZN(n8691) );
  INV_X1 U10047 ( .A(n8691), .ZN(n8291) );
  NAND2_X1 U10048 ( .A1(n11892), .A2(n8291), .ZN(n8703) );
  INV_X1 U10049 ( .A(n8703), .ZN(n8292) );
  NAND2_X1 U10050 ( .A1(n8292), .A2(n11814), .ZN(n8714) );
  INV_X1 U10051 ( .A(n8725), .ZN(n8293) );
  INV_X1 U10052 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n13186) );
  NAND2_X1 U10053 ( .A1(n8293), .A2(n13186), .ZN(n8738) );
  INV_X1 U10054 ( .A(n8756), .ZN(n8295) );
  NOR2_X1 U10055 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(P3_REG3_REG_26__SCAN_IN), 
        .ZN(n8294) );
  NAND2_X1 U10056 ( .A1(n8295), .A2(n8294), .ZN(n8757) );
  NAND2_X1 U10057 ( .A1(n8757), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8296) );
  NAND2_X1 U10058 ( .A1(n13424), .A2(n8296), .ZN(n13444) );
  NAND2_X1 U10059 ( .A1(n8543), .A2(n13444), .ZN(n8299) );
  NAND2_X1 U10060 ( .A1(n8759), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8298) );
  INV_X1 U10061 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n10405) );
  NAND2_X1 U10062 ( .A1(n10405), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8388) );
  INV_X1 U10063 ( .A(n8388), .ZN(n8302) );
  NAND2_X1 U10064 ( .A1(n8303), .A2(n8302), .ZN(n8378) );
  NAND2_X1 U10065 ( .A1(n10396), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8304) );
  NAND2_X1 U10066 ( .A1(n10446), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8306) );
  INV_X1 U10067 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9844) );
  NAND2_X1 U10068 ( .A1(n9844), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8305) );
  AND2_X1 U10069 ( .A1(n8306), .A2(n8305), .ZN(n8394) );
  NAND2_X1 U10070 ( .A1(n9871), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8308) );
  INV_X1 U10071 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9849) );
  NAND2_X1 U10072 ( .A1(n9849), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8307) );
  AND2_X1 U10073 ( .A1(n8308), .A2(n8307), .ZN(n8405) );
  NAND2_X1 U10074 ( .A1(n8309), .A2(n8308), .ZN(n8420) );
  NAND2_X1 U10075 ( .A1(n9865), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8311) );
  NAND2_X1 U10076 ( .A1(n9852), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8310) );
  AND2_X1 U10077 ( .A1(n8311), .A2(n8310), .ZN(n8419) );
  NAND2_X1 U10078 ( .A1(n8420), .A2(n8419), .ZN(n8312) );
  NAND2_X1 U10079 ( .A1(n9859), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8314) );
  INV_X1 U10080 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9860) );
  NAND2_X1 U10081 ( .A1(n9860), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8313) );
  AND2_X1 U10082 ( .A1(n8314), .A2(n8313), .ZN(n8434) );
  NAND2_X1 U10083 ( .A1(n9881), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8315) );
  NAND2_X1 U10084 ( .A1(n9883), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8316) );
  NAND2_X1 U10085 ( .A1(n9925), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U10086 ( .A1(n9930), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8317) );
  NAND2_X1 U10087 ( .A1(n8318), .A2(n8317), .ZN(n8468) );
  NAND2_X1 U10088 ( .A1(n9934), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8320) );
  NAND2_X1 U10089 ( .A1(n9933), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8319) );
  AND2_X1 U10090 ( .A1(n8320), .A2(n8319), .ZN(n8483) );
  NAND2_X1 U10091 ( .A1(n8484), .A2(n8483), .ZN(n8486) );
  NAND2_X1 U10092 ( .A1(n8486), .A2(n8320), .ZN(n8501) );
  NAND2_X1 U10093 ( .A1(n10040), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U10094 ( .A1(n10039), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8321) );
  AND2_X1 U10095 ( .A1(n8322), .A2(n8321), .ZN(n8500) );
  NAND2_X1 U10096 ( .A1(n8501), .A2(n8500), .ZN(n8503) );
  NAND2_X1 U10097 ( .A1(n8503), .A2(n8322), .ZN(n8511) );
  NAND2_X1 U10098 ( .A1(n10056), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8324) );
  INV_X1 U10099 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10055) );
  NAND2_X1 U10100 ( .A1(n10055), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8323) );
  AND2_X1 U10101 ( .A1(n8324), .A2(n8323), .ZN(n8510) );
  NAND2_X1 U10102 ( .A1(n8511), .A2(n8510), .ZN(n8513) );
  NAND2_X1 U10103 ( .A1(n8513), .A2(n8324), .ZN(n8535) );
  NAND2_X1 U10104 ( .A1(n10084), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8326) );
  INV_X1 U10105 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10089) );
  NAND2_X1 U10106 ( .A1(n10089), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8325) );
  AND2_X1 U10107 ( .A1(n8326), .A2(n8325), .ZN(n8534) );
  NAND2_X1 U10108 ( .A1(n8535), .A2(n8534), .ZN(n8537) );
  NAND2_X1 U10109 ( .A1(n8537), .A2(n8326), .ZN(n8551) );
  NAND2_X1 U10110 ( .A1(n10276), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8328) );
  NAND2_X1 U10111 ( .A1(n10287), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8327) );
  OR2_X1 U10112 ( .A1(n8329), .A2(n10334), .ZN(n8330) );
  NAND2_X1 U10113 ( .A1(n10582), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8333) );
  INV_X1 U10114 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10586) );
  NAND2_X1 U10115 ( .A1(n10586), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8332) );
  NAND2_X1 U10116 ( .A1(n8579), .A2(n8333), .ZN(n8594) );
  NAND2_X1 U10117 ( .A1(n10785), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8335) );
  INV_X1 U10118 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10783) );
  NAND2_X1 U10119 ( .A1(n10783), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8334) );
  NAND2_X1 U10120 ( .A1(n8594), .A2(n8593), .ZN(n8596) );
  NAND2_X1 U10121 ( .A1(n10895), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8337) );
  NAND2_X1 U10122 ( .A1(n9289), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8336) );
  NAND2_X1 U10123 ( .A1(n11038), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8339) );
  INV_X1 U10124 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11044) );
  NAND2_X1 U10125 ( .A1(n11044), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8338) );
  NAND2_X1 U10126 ( .A1(n8626), .A2(n8339), .ZN(n8641) );
  NAND2_X1 U10127 ( .A1(n11281), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8341) );
  NAND2_X1 U10128 ( .A1(n11284), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8340) );
  NAND2_X1 U10129 ( .A1(n8641), .A2(n8640), .ZN(n8643) );
  INV_X1 U10130 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11583) );
  NAND2_X1 U10131 ( .A1(n11583), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8343) );
  INV_X1 U10132 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11585) );
  NAND2_X1 U10133 ( .A1(n11585), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8342) );
  NAND2_X1 U10134 ( .A1(n8344), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8346) );
  INV_X1 U10135 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12053) );
  NAND2_X1 U10136 ( .A1(n12053), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8349) );
  INV_X1 U10137 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12501) );
  NAND2_X1 U10138 ( .A1(n12501), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8347) );
  NAND2_X1 U10139 ( .A1(n8349), .A2(n8347), .ZN(n8687) );
  INV_X1 U10140 ( .A(n8687), .ZN(n8348) );
  INV_X1 U10141 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8351) );
  NAND2_X1 U10142 ( .A1(n8351), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8354) );
  INV_X1 U10143 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n14508) );
  NAND2_X1 U10144 ( .A1(n14508), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8352) );
  NAND2_X1 U10145 ( .A1(n8354), .A2(n8352), .ZN(n8699) );
  INV_X1 U10146 ( .A(n8699), .ZN(n8353) );
  XNOR2_X1 U10147 ( .A(n14504), .B(P2_DATAO_REG_23__SCAN_IN), .ZN(n8710) );
  NAND2_X1 U10148 ( .A1(n14504), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8355) );
  NAND2_X1 U10149 ( .A1(n8356), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8357) );
  INV_X1 U10150 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n14499) );
  INV_X1 U10151 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8359) );
  NAND2_X1 U10152 ( .A1(n8359), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8361) );
  INV_X1 U10153 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14496) );
  NAND2_X1 U10154 ( .A1(n14496), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8360) );
  AND2_X1 U10155 ( .A1(n8361), .A2(n8360), .ZN(n8732) );
  INV_X1 U10156 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15201) );
  NAND2_X1 U10157 ( .A1(n15201), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8364) );
  INV_X1 U10158 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14492) );
  NAND2_X1 U10159 ( .A1(n14492), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8362) );
  NAND2_X1 U10160 ( .A1(n8364), .A2(n8362), .ZN(n8744) );
  INV_X1 U10161 ( .A(n8744), .ZN(n8363) );
  INV_X1 U10162 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n12499) );
  NAND2_X1 U10163 ( .A1(n12499), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8367) );
  INV_X1 U10164 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14489) );
  NAND2_X1 U10165 ( .A1(n14489), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8365) );
  NAND2_X1 U10166 ( .A1(n8367), .A2(n8365), .ZN(n8752) );
  INV_X1 U10167 ( .A(n8752), .ZN(n8366) );
  INV_X1 U10168 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12760) );
  NAND2_X1 U10169 ( .A1(n12760), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8772) );
  INV_X1 U10170 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14486) );
  NAND2_X1 U10171 ( .A1(n14486), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U10172 ( .A1(n8772), .A2(n8368), .ZN(n8769) );
  XNOR2_X1 U10173 ( .A(n8771), .B(n8769), .ZN(n12033) );
  NAND2_X1 U10174 ( .A1(n12033), .A2(n12560), .ZN(n8373) );
  INV_X1 U10175 ( .A(SI_28_), .ZN(n12034) );
  OR2_X1 U10176 ( .A1(n7221), .A2(n12034), .ZN(n8372) );
  NAND2_X1 U10177 ( .A1(n7222), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8376) );
  NAND2_X1 U10178 ( .A1(n8521), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8375) );
  NAND2_X1 U10179 ( .A1(n8543), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8374) );
  NAND2_X1 U10180 ( .A1(n8377), .A2(n8388), .ZN(n8379) );
  AND2_X1 U10181 ( .A1(n8379), .A2(n8378), .ZN(n9855) );
  INV_X1 U10182 ( .A(SI_1_), .ZN(n9854) );
  NAND2_X1 U10183 ( .A1(n7223), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8386) );
  NAND2_X1 U10184 ( .A1(n8521), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8385) );
  NAND2_X1 U10185 ( .A1(n7250), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8384) );
  NAND2_X1 U10186 ( .A1(n8524), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8383) );
  INV_X1 U10187 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8900) );
  NAND2_X1 U10188 ( .A1(n8900), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U10189 ( .A1(n8388), .A2(n8387), .ZN(n8389) );
  MUX2_X1 U10190 ( .A(n8389), .B(SI_0_), .S(n10404), .Z(n13814) );
  MUX2_X1 U10191 ( .A(P3_IR_REG_0__SCAN_IN), .B(n13814), .S(n10126), .Z(n10596) );
  NAND2_X1 U10192 ( .A1(n13264), .A2(n10596), .ZN(n11171) );
  NAND2_X1 U10193 ( .A1(n15720), .A2(n15697), .ZN(n15714) );
  NAND2_X1 U10194 ( .A1(n15716), .A2(n15714), .ZN(n8399) );
  NAND2_X1 U10195 ( .A1(n8524), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8393) );
  NAND2_X1 U10196 ( .A1(n8520), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8392) );
  NAND2_X1 U10197 ( .A1(n7250), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8391) );
  NAND2_X1 U10198 ( .A1(n8521), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8390) );
  OR2_X1 U10199 ( .A1(n7221), .A2(SI_2_), .ZN(n8398) );
  XNOR2_X1 U10200 ( .A(n8395), .B(n8394), .ZN(n9909) );
  OR2_X1 U10201 ( .A1(n7220), .A2(n9909), .ZN(n8397) );
  OR2_X1 U10202 ( .A1(n10126), .A2(n11454), .ZN(n8396) );
  NAND2_X1 U10203 ( .A1(n11172), .A2(n10714), .ZN(n12614) );
  NAND2_X1 U10204 ( .A1(n13261), .A2(n15730), .ZN(n12622) );
  NAND2_X1 U10205 ( .A1(n12614), .A2(n12622), .ZN(n8796) );
  NAND2_X1 U10206 ( .A1(n8399), .A2(n8796), .ZN(n11056) );
  INV_X1 U10207 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11880) );
  NAND2_X1 U10208 ( .A1(n8524), .A2(n11880), .ZN(n8403) );
  NAND2_X1 U10209 ( .A1(n8520), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U10210 ( .A1(n7250), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8401) );
  NAND2_X1 U10211 ( .A1(n8521), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8400) );
  OR2_X1 U10212 ( .A1(n7221), .A2(SI_3_), .ZN(n8411) );
  XNOR2_X1 U10213 ( .A(n8406), .B(n8405), .ZN(n9912) );
  OR2_X1 U10214 ( .A1(n7219), .A2(n9912), .ZN(n8410) );
  NAND2_X1 U10215 ( .A1(n7964), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8407) );
  MUX2_X1 U10216 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8407), .S(
        P3_IR_REG_3__SCAN_IN), .Z(n8408) );
  OR2_X1 U10217 ( .A1(n10126), .A2(n15521), .ZN(n8409) );
  NAND2_X1 U10218 ( .A1(n15722), .A2(n11186), .ZN(n12623) );
  INV_X1 U10219 ( .A(n15722), .ZN(n13260) );
  INV_X1 U10220 ( .A(n11186), .ZN(n11249) );
  NAND2_X1 U10221 ( .A1(n13260), .A2(n11249), .ZN(n12624) );
  NAND2_X1 U10222 ( .A1(n12623), .A2(n12624), .ZN(n12575) );
  NAND2_X1 U10223 ( .A1(n11172), .A2(n15730), .ZN(n11057) );
  AND2_X1 U10224 ( .A1(n12575), .A2(n11057), .ZN(n8412) );
  NAND2_X1 U10225 ( .A1(n11056), .A2(n8412), .ZN(n11058) );
  NAND2_X1 U10226 ( .A1(n13260), .A2(n11186), .ZN(n8413) );
  NAND2_X1 U10227 ( .A1(n11058), .A2(n8413), .ZN(n11193) );
  NAND2_X1 U10228 ( .A1(n8520), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8418) );
  NAND2_X1 U10229 ( .A1(n12552), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8417) );
  AND2_X1 U10230 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8414) );
  OR2_X1 U10231 ( .A1(n8414), .A2(n8427), .ZN(n11197) );
  NAND2_X1 U10232 ( .A1(n8524), .A2(n11197), .ZN(n8416) );
  NAND2_X1 U10233 ( .A1(n7250), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8415) );
  OR2_X1 U10234 ( .A1(n7221), .A2(SI_4_), .ZN(n8424) );
  XNOR2_X1 U10235 ( .A(n8420), .B(n8419), .ZN(n9902) );
  OR2_X1 U10236 ( .A1(n7219), .A2(n9902), .ZN(n8423) );
  NAND2_X1 U10237 ( .A1(n8436), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8421) );
  XNOR2_X1 U10238 ( .A(n8421), .B(P3_IR_REG_4__SCAN_IN), .ZN(n15540) );
  OR2_X1 U10239 ( .A1(n10126), .A2(n15540), .ZN(n8422) );
  NAND2_X1 U10240 ( .A1(n11238), .A2(n15772), .ZN(n12629) );
  INV_X1 U10241 ( .A(n11238), .ZN(n13259) );
  INV_X1 U10242 ( .A(n15772), .ZN(n8425) );
  NAND2_X1 U10243 ( .A1(n13259), .A2(n8425), .ZN(n12630) );
  NAND2_X1 U10244 ( .A1(n12629), .A2(n12630), .ZN(n11192) );
  NAND2_X1 U10245 ( .A1(n13259), .A2(n15772), .ZN(n8426) );
  NAND2_X1 U10246 ( .A1(n8520), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8433) );
  NAND2_X1 U10247 ( .A1(n8521), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8432) );
  OR2_X1 U10248 ( .A1(n8428), .A2(n8427), .ZN(n8429) );
  NAND2_X1 U10249 ( .A1(n8442), .A2(n8429), .ZN(n11241) );
  NAND2_X1 U10250 ( .A1(n8524), .A2(n11241), .ZN(n8431) );
  NAND2_X1 U10251 ( .A1(n7250), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8430) );
  OR2_X1 U10252 ( .A1(n7221), .A2(SI_5_), .ZN(n8441) );
  XNOR2_X1 U10253 ( .A(n8435), .B(n8434), .ZN(n9915) );
  OR2_X1 U10254 ( .A1(n7220), .A2(n9915), .ZN(n8440) );
  INV_X1 U10255 ( .A(n8436), .ZN(n8437) );
  NAND2_X1 U10256 ( .A1(n8437), .A2(n7390), .ZN(n8448) );
  NAND2_X1 U10257 ( .A1(n8448), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8438) );
  XNOR2_X1 U10258 ( .A(n8438), .B(P3_IR_REG_5__SCAN_IN), .ZN(n11457) );
  OR2_X1 U10259 ( .A1(n10126), .A2(n11457), .ZN(n8439) );
  NAND2_X1 U10260 ( .A1(n11226), .A2(n11242), .ZN(n12634) );
  INV_X1 U10261 ( .A(n11226), .ZN(n13258) );
  INV_X1 U10262 ( .A(n11242), .ZN(n15789) );
  NAND2_X1 U10263 ( .A1(n13258), .A2(n15789), .ZN(n12635) );
  NAND2_X1 U10264 ( .A1(n8520), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8447) );
  NAND2_X1 U10265 ( .A1(n12552), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8446) );
  NAND2_X1 U10266 ( .A1(n8442), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8443) );
  NAND2_X1 U10267 ( .A1(n8458), .A2(n8443), .ZN(n11333) );
  NAND2_X1 U10268 ( .A1(n8524), .A2(n11333), .ZN(n8445) );
  NAND2_X1 U10269 ( .A1(n7250), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8444) );
  INV_X1 U10270 ( .A(n8448), .ZN(n8450) );
  NAND2_X1 U10271 ( .A1(n8450), .A2(n8449), .ZN(n8465) );
  NAND2_X1 U10272 ( .A1(n8465), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8451) );
  XNOR2_X1 U10273 ( .A(n8451), .B(n7389), .ZN(n11460) );
  INV_X1 U10274 ( .A(SI_6_), .ZN(n9923) );
  OR2_X1 U10275 ( .A1(n7221), .A2(n9923), .ZN(n8455) );
  XNOR2_X1 U10276 ( .A(n9883), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8452) );
  XNOR2_X1 U10277 ( .A(n8453), .B(n8452), .ZN(n9924) );
  OR2_X1 U10278 ( .A1(n7219), .A2(n9924), .ZN(n8454) );
  OAI211_X1 U10279 ( .C1(n10126), .C2(n11460), .A(n8455), .B(n8454), .ZN(
        n11334) );
  NAND2_X1 U10280 ( .A1(n11350), .A2(n11334), .ZN(n12639) );
  INV_X1 U10281 ( .A(n11350), .ZN(n13257) );
  INV_X1 U10282 ( .A(n11334), .ZN(n11277) );
  NAND2_X1 U10283 ( .A1(n13257), .A2(n11277), .ZN(n12640) );
  NAND2_X1 U10284 ( .A1(n12639), .A2(n12640), .ZN(n11269) );
  NAND2_X1 U10285 ( .A1(n11226), .A2(n15789), .ZN(n11270) );
  AND2_X1 U10286 ( .A1(n11269), .A2(n11270), .ZN(n8456) );
  NAND2_X1 U10287 ( .A1(n13257), .A2(n11334), .ZN(n8457) );
  NAND2_X1 U10288 ( .A1(n11268), .A2(n8457), .ZN(n11632) );
  NAND2_X1 U10289 ( .A1(n7223), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8463) );
  NAND2_X1 U10290 ( .A1(n12552), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8462) );
  AND2_X1 U10291 ( .A1(n8458), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8459) );
  OR2_X1 U10292 ( .A1(n8459), .A2(n8476), .ZN(n11638) );
  NAND2_X1 U10293 ( .A1(n8524), .A2(n11638), .ZN(n8461) );
  NAND2_X1 U10294 ( .A1(n7250), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8460) );
  NAND4_X1 U10295 ( .A1(n8463), .A2(n8462), .A3(n8461), .A4(n8460), .ZN(n13256) );
  OAI21_X1 U10296 ( .B1(n8465), .B2(P3_IR_REG_6__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8466) );
  MUX2_X1 U10297 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8466), .S(
        P3_IR_REG_7__SCAN_IN), .Z(n8467) );
  AND2_X1 U10298 ( .A1(n8464), .A2(n8467), .ZN(n15601) );
  NAND2_X1 U10299 ( .A1(n8469), .A2(n8468), .ZN(n8470) );
  AND2_X1 U10300 ( .A1(n8471), .A2(n8470), .ZN(n9850) );
  OR2_X1 U10301 ( .A1(n7220), .A2(n9850), .ZN(n8473) );
  OR2_X1 U10302 ( .A1(n7221), .A2(SI_7_), .ZN(n8472) );
  OAI211_X1 U10303 ( .C1(n15601), .C2(n10126), .A(n8473), .B(n8472), .ZN(
        n15830) );
  XNOR2_X1 U10304 ( .A(n13256), .B(n15830), .ZN(n11631) );
  NAND2_X1 U10305 ( .A1(n11632), .A2(n11631), .ZN(n8475) );
  INV_X1 U10306 ( .A(n15830), .ZN(n11639) );
  NAND2_X1 U10307 ( .A1(n13256), .A2(n11639), .ZN(n8474) );
  NAND2_X1 U10308 ( .A1(n8521), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U10309 ( .A1(n8520), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8480) );
  NOR2_X1 U10310 ( .A1(n8476), .A2(n11890), .ZN(n8477) );
  OR2_X1 U10311 ( .A1(n8491), .A2(n8477), .ZN(n11999) );
  NAND2_X1 U10312 ( .A1(n8524), .A2(n11999), .ZN(n8479) );
  NAND2_X1 U10313 ( .A1(n7250), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U10314 ( .A1(n8464), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8482) );
  XNOR2_X1 U10315 ( .A(n8482), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11463) );
  INV_X1 U10316 ( .A(SI_8_), .ZN(n9905) );
  OR2_X1 U10317 ( .A1(n7221), .A2(n9905), .ZN(n8488) );
  OR2_X1 U10318 ( .A1(n8484), .A2(n8483), .ZN(n8485) );
  NAND2_X1 U10319 ( .A1(n8486), .A2(n8485), .ZN(n9906) );
  OR2_X1 U10320 ( .A1(n7220), .A2(n9906), .ZN(n8487) );
  OAI211_X1 U10321 ( .C1(n10126), .C2(n15617), .A(n8488), .B(n8487), .ZN(
        n15854) );
  NAND2_X1 U10322 ( .A1(n12009), .A2(n15854), .ZN(n12649) );
  INV_X1 U10323 ( .A(n12009), .ZN(n13255) );
  INV_X1 U10324 ( .A(n15854), .ZN(n8489) );
  NAND2_X1 U10325 ( .A1(n13255), .A2(n8489), .ZN(n12650) );
  NAND2_X1 U10326 ( .A1(n12009), .A2(n8489), .ZN(n8490) );
  NAND2_X1 U10327 ( .A1(n8521), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8496) );
  NAND2_X1 U10328 ( .A1(n8520), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8495) );
  OR2_X1 U10329 ( .A1(n8491), .A2(n11787), .ZN(n8492) );
  NAND2_X1 U10330 ( .A1(n8522), .A2(n8492), .ZN(n12011) );
  NAND2_X1 U10331 ( .A1(n8524), .A2(n12011), .ZN(n8494) );
  NAND2_X1 U10332 ( .A1(n7250), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8493) );
  OR2_X1 U10333 ( .A1(n8497), .A2(n8554), .ZN(n8499) );
  XNOR2_X1 U10334 ( .A(n8499), .B(n8498), .ZN(n15637) );
  INV_X1 U10335 ( .A(n15637), .ZN(n11438) );
  OR2_X1 U10336 ( .A1(n8501), .A2(n8500), .ZN(n8502) );
  AND2_X1 U10337 ( .A1(n8503), .A2(n8502), .ZN(n9907) );
  OR2_X1 U10338 ( .A1(n7219), .A2(n9907), .ZN(n8505) );
  OR2_X1 U10339 ( .A1(n7221), .A2(SI_9_), .ZN(n8504) );
  OAI211_X1 U10340 ( .C1(n11438), .C2(n10126), .A(n8505), .B(n8504), .ZN(
        n15870) );
  NAND2_X1 U10341 ( .A1(n8521), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8509) );
  NAND2_X1 U10342 ( .A1(n8520), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8508) );
  XNOR2_X1 U10343 ( .A(n8522), .B(P3_REG3_REG_10__SCAN_IN), .ZN(n12140) );
  NAND2_X1 U10344 ( .A1(n8524), .A2(n12140), .ZN(n8507) );
  NAND2_X1 U10345 ( .A1(n7250), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8506) );
  NAND4_X1 U10346 ( .A1(n8509), .A2(n8508), .A3(n8507), .A4(n8506), .ZN(n13254) );
  OR2_X1 U10347 ( .A1(n8511), .A2(n8510), .ZN(n8512) );
  AND2_X1 U10348 ( .A1(n8513), .A2(n8512), .ZN(n9899) );
  OR2_X1 U10349 ( .A1(n7219), .A2(n9899), .ZN(n8518) );
  OR2_X1 U10350 ( .A1(n7221), .A2(SI_10_), .ZN(n8517) );
  OR2_X1 U10351 ( .A1(n8514), .A2(n8554), .ZN(n8515) );
  XNOR2_X1 U10352 ( .A(n8515), .B(n8529), .ZN(n15658) );
  INV_X1 U10353 ( .A(n15658), .ZN(n11452) );
  OR2_X1 U10354 ( .A1(n10126), .A2(n11452), .ZN(n8516) );
  XNOR2_X1 U10355 ( .A(n13254), .B(n15892), .ZN(n12658) );
  NAND2_X1 U10356 ( .A1(n13254), .A2(n15892), .ZN(n8519) );
  NAND2_X1 U10357 ( .A1(n8520), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U10358 ( .A1(n8521), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8527) );
  OAI21_X1 U10359 ( .B1(n8522), .B2(P3_REG3_REG_10__SCAN_IN), .A(
        P3_REG3_REG_11__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U10360 ( .A1(n8523), .A2(n8544), .ZN(n12249) );
  NAND2_X1 U10361 ( .A1(n8524), .A2(n12249), .ZN(n8526) );
  NAND2_X1 U10362 ( .A1(n7250), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8525) );
  NAND2_X1 U10363 ( .A1(n8514), .A2(n8529), .ZN(n8530) );
  INV_X1 U10364 ( .A(n8565), .ZN(n8533) );
  NAND2_X1 U10365 ( .A1(n8530), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8531) );
  MUX2_X1 U10366 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8531), .S(
        P3_IR_REG_11__SCAN_IN), .Z(n8532) );
  NAND2_X1 U10367 ( .A1(n8533), .A2(n8532), .ZN(n11674) );
  OR2_X1 U10368 ( .A1(n7221), .A2(SI_11_), .ZN(n8539) );
  OR2_X1 U10369 ( .A1(n8535), .A2(n8534), .ZN(n8536) );
  AND2_X1 U10370 ( .A1(n8537), .A2(n8536), .ZN(n9918) );
  OR2_X1 U10371 ( .A1(n7220), .A2(n9918), .ZN(n8538) );
  OAI211_X1 U10372 ( .C1(n11682), .C2(n10126), .A(n8539), .B(n8538), .ZN(
        n15910) );
  NAND2_X1 U10373 ( .A1(n12164), .A2(n15910), .ZN(n8540) );
  NAND2_X1 U10374 ( .A1(n12201), .A2(n8540), .ZN(n8542) );
  INV_X1 U10375 ( .A(n15910), .ZN(n8800) );
  NAND2_X1 U10376 ( .A1(n13253), .A2(n8800), .ZN(n8541) );
  NAND2_X1 U10377 ( .A1(n12552), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U10378 ( .A1(n8520), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8548) );
  AND2_X1 U10379 ( .A1(n8544), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8545) );
  OR2_X1 U10380 ( .A1(n8545), .A2(n8570), .ZN(n12313) );
  NAND2_X1 U10381 ( .A1(n8524), .A2(n12313), .ZN(n8547) );
  NAND2_X1 U10382 ( .A1(n8759), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8546) );
  NAND4_X1 U10383 ( .A1(n8549), .A2(n8548), .A3(n8547), .A4(n8546), .ZN(n13252) );
  OR2_X1 U10384 ( .A1(n8551), .A2(n8550), .ZN(n8552) );
  AND2_X1 U10385 ( .A1(n8553), .A2(n8552), .ZN(n9921) );
  OR2_X1 U10386 ( .A1(n7219), .A2(n9921), .ZN(n8558) );
  OR2_X1 U10387 ( .A1(n7221), .A2(SI_12_), .ZN(n8557) );
  OR2_X1 U10388 ( .A1(n8565), .A2(n8554), .ZN(n8555) );
  XNOR2_X1 U10389 ( .A(n8555), .B(n8564), .ZN(n13276) );
  INV_X1 U10390 ( .A(n13276), .ZN(n13269) );
  OR2_X1 U10391 ( .A1(n10126), .A2(n13269), .ZN(n8556) );
  AND2_X1 U10392 ( .A1(n13252), .A2(n12316), .ZN(n8560) );
  INV_X1 U10393 ( .A(n13252), .ZN(n13657) );
  NAND2_X1 U10394 ( .A1(n13657), .A2(n15934), .ZN(n8559) );
  NAND2_X1 U10395 ( .A1(n8561), .A2(n10333), .ZN(n8562) );
  NAND2_X1 U10396 ( .A1(n8563), .A2(n8562), .ZN(n9937) );
  NAND2_X1 U10397 ( .A1(n9937), .A2(n12560), .ZN(n8569) );
  INV_X1 U10398 ( .A(n7221), .ZN(n8665) );
  INV_X1 U10399 ( .A(n10126), .ZN(n8664) );
  NAND2_X1 U10400 ( .A1(n8565), .A2(n8564), .ZN(n8580) );
  NAND2_X1 U10401 ( .A1(n8580), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8567) );
  XNOR2_X1 U10402 ( .A(n8567), .B(n8566), .ZN(n13299) );
  AOI22_X1 U10403 ( .A1(n8665), .A2(n11848), .B1(n8664), .B2(n13299), .ZN(
        n8568) );
  NAND2_X1 U10404 ( .A1(n12552), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U10405 ( .A1(n8520), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8574) );
  OR2_X1 U10406 ( .A1(n8570), .A2(n11915), .ZN(n8571) );
  NAND2_X1 U10407 ( .A1(n8585), .A2(n8571), .ZN(n13660) );
  NAND2_X1 U10408 ( .A1(n8524), .A2(n13660), .ZN(n8573) );
  NAND2_X1 U10409 ( .A1(n8759), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8572) );
  NAND2_X1 U10410 ( .A1(n13664), .A2(n12306), .ZN(n12676) );
  NAND2_X1 U10411 ( .A1(n13742), .A2(n13644), .ZN(n12677) );
  NAND2_X1 U10412 ( .A1(n13664), .A2(n13644), .ZN(n13637) );
  OR2_X1 U10413 ( .A1(n8577), .A2(n8576), .ZN(n8578) );
  NAND2_X1 U10414 ( .A1(n8579), .A2(n8578), .ZN(n9986) );
  NAND2_X1 U10415 ( .A1(n9986), .A2(n12560), .ZN(n8584) );
  OAI21_X1 U10416 ( .B1(n8580), .B2(P3_IR_REG_13__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8582) );
  INV_X1 U10417 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8581) );
  AOI22_X1 U10418 ( .A1(n8665), .A2(n11818), .B1(n8664), .B2(n13321), .ZN(
        n8583) );
  NAND2_X1 U10419 ( .A1(n12552), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8590) );
  NAND2_X1 U10420 ( .A1(n8520), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U10421 ( .A1(n8585), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8586) );
  NAND2_X1 U10422 ( .A1(n8614), .A2(n8586), .ZN(n13647) );
  NAND2_X1 U10423 ( .A1(n8524), .A2(n13647), .ZN(n8588) );
  NAND2_X1 U10424 ( .A1(n8759), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8587) );
  NAND2_X1 U10425 ( .A1(n13793), .A2(n13656), .ZN(n8591) );
  NAND2_X1 U10426 ( .A1(n8592), .A2(n12584), .ZN(n13622) );
  NAND2_X1 U10427 ( .A1(n13622), .A2(n13623), .ZN(n8606) );
  OR2_X1 U10428 ( .A1(n8594), .A2(n8593), .ZN(n8595) );
  NAND2_X1 U10429 ( .A1(n8596), .A2(n8595), .ZN(n10041) );
  NAND2_X1 U10430 ( .A1(n10041), .A2(n12560), .ZN(n8601) );
  NAND2_X1 U10431 ( .A1(n8597), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8599) );
  INV_X1 U10432 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8598) );
  XNOR2_X1 U10433 ( .A(n8599), .B(n8598), .ZN(n13340) );
  AOI22_X1 U10434 ( .A1(n8665), .A2(n11711), .B1(n8664), .B2(n13340), .ZN(
        n8600) );
  NAND2_X1 U10435 ( .A1(n12552), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8605) );
  NAND2_X1 U10436 ( .A1(n7223), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8604) );
  XNOR2_X1 U10437 ( .A(n8614), .B(P3_REG3_REG_15__SCAN_IN), .ZN(n13630) );
  NAND2_X1 U10438 ( .A1(n8524), .A2(n13630), .ZN(n8603) );
  NAND2_X1 U10439 ( .A1(n8759), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8602) );
  NAND4_X1 U10440 ( .A1(n8605), .A2(n8604), .A3(n8603), .A4(n8602), .ZN(n13641) );
  NAND2_X1 U10441 ( .A1(n13789), .A2(n13641), .ZN(n12685) );
  NAND2_X1 U10442 ( .A1(n12684), .A2(n12685), .ZN(n12583) );
  INV_X1 U10443 ( .A(n13641), .ZN(n13613) );
  OR2_X1 U10444 ( .A1(n13789), .A2(n13613), .ZN(n13607) );
  OR2_X1 U10445 ( .A1(n8608), .A2(n8607), .ZN(n8609) );
  NAND2_X1 U10446 ( .A1(n8610), .A2(n8609), .ZN(n10042) );
  OR2_X1 U10447 ( .A1(n10042), .A2(n7220), .ZN(n8613) );
  NAND2_X1 U10448 ( .A1(n8627), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8611) );
  XNOR2_X1 U10449 ( .A(n8611), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13348) );
  AOI22_X1 U10450 ( .A1(n8665), .A2(SI_16_), .B1(n8664), .B2(n13348), .ZN(
        n8612) );
  NAND2_X1 U10451 ( .A1(n8613), .A2(n8612), .ZN(n13726) );
  NAND2_X1 U10452 ( .A1(n12552), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8620) );
  NAND2_X1 U10453 ( .A1(n7223), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8619) );
  OAI21_X1 U10454 ( .B1(n8614), .B2(P3_REG3_REG_15__SCAN_IN), .A(
        P3_REG3_REG_16__SCAN_IN), .ZN(n8615) );
  INV_X1 U10455 ( .A(n8615), .ZN(n8616) );
  OR2_X1 U10456 ( .A1(n8616), .A2(n8632), .ZN(n13615) );
  NAND2_X1 U10457 ( .A1(n8524), .A2(n13615), .ZN(n8618) );
  NAND2_X1 U10458 ( .A1(n8759), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8617) );
  OR2_X1 U10459 ( .A1(n13726), .A2(n13591), .ZN(n12690) );
  NAND2_X1 U10460 ( .A1(n13726), .A2(n13591), .ZN(n12688) );
  INV_X1 U10461 ( .A(n13611), .ZN(n8621) );
  AND2_X1 U10462 ( .A1(n13607), .A2(n8621), .ZN(n8622) );
  NAND2_X2 U10463 ( .A1(n13606), .A2(n8622), .ZN(n13608) );
  OR2_X1 U10464 ( .A1(n8624), .A2(n8623), .ZN(n8625) );
  NAND2_X1 U10465 ( .A1(n8626), .A2(n8625), .ZN(n10083) );
  NAND2_X1 U10466 ( .A1(n10083), .A2(n12560), .ZN(n8631) );
  NOR2_X2 U10467 ( .A1(n8627), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n8645) );
  INV_X1 U10468 ( .A(n8645), .ZN(n8628) );
  NAND2_X1 U10469 ( .A1(n8628), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8629) );
  XNOR2_X1 U10470 ( .A(n8629), .B(n8644), .ZN(n13379) );
  AOI22_X1 U10471 ( .A1(n8665), .A2(n11840), .B1(n8664), .B2(n13379), .ZN(
        n8630) );
  NAND2_X1 U10472 ( .A1(n8631), .A2(n8630), .ZN(n13784) );
  NAND2_X1 U10473 ( .A1(n12552), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8637) );
  NAND2_X1 U10474 ( .A1(n7223), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8636) );
  NOR2_X1 U10475 ( .A1(n8632), .A2(n11901), .ZN(n8633) );
  OR2_X1 U10476 ( .A1(n8650), .A2(n8633), .ZN(n13595) );
  NAND2_X1 U10477 ( .A1(n8524), .A2(n13595), .ZN(n8635) );
  NAND2_X1 U10478 ( .A1(n8759), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8634) );
  NAND4_X1 U10479 ( .A1(n8637), .A2(n8636), .A3(n8635), .A4(n8634), .ZN(n13251) );
  OR2_X1 U10480 ( .A1(n13784), .A2(n13251), .ZN(n13575) );
  NAND2_X1 U10481 ( .A1(n13784), .A2(n13251), .ZN(n12694) );
  NAND2_X1 U10482 ( .A1(n13575), .A2(n12694), .ZN(n8802) );
  OR2_X1 U10483 ( .A1(n13726), .A2(n13626), .ZN(n13586) );
  AND2_X1 U10484 ( .A1(n8802), .A2(n13586), .ZN(n8638) );
  INV_X1 U10485 ( .A(n13251), .ZN(n13614) );
  OR2_X1 U10486 ( .A1(n13784), .A2(n13614), .ZN(n8639) );
  OR2_X1 U10487 ( .A1(n8641), .A2(n8640), .ZN(n8642) );
  NAND2_X1 U10488 ( .A1(n8643), .A2(n8642), .ZN(n10106) );
  OR2_X1 U10489 ( .A1(n10106), .A2(n7219), .ZN(n8649) );
  INV_X1 U10490 ( .A(n8661), .ZN(n8646) );
  NAND2_X1 U10491 ( .A1(n8646), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8647) );
  XNOR2_X1 U10492 ( .A(n8647), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13405) );
  AOI22_X1 U10493 ( .A1(n8665), .A2(SI_18_), .B1(n8664), .B2(n13405), .ZN(
        n8648) );
  NAND2_X1 U10494 ( .A1(n8649), .A2(n8648), .ZN(n13717) );
  NAND2_X1 U10495 ( .A1(n12552), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8655) );
  NAND2_X1 U10496 ( .A1(n8520), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8654) );
  OR2_X1 U10497 ( .A1(n8650), .A2(n11801), .ZN(n8651) );
  NAND2_X1 U10498 ( .A1(n8668), .A2(n8651), .ZN(n13581) );
  NAND2_X1 U10499 ( .A1(n8524), .A2(n13581), .ZN(n8653) );
  NAND2_X1 U10500 ( .A1(n8759), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8652) );
  NAND2_X1 U10501 ( .A1(n13717), .A2(n13590), .ZN(n12693) );
  INV_X1 U10502 ( .A(n13590), .ZN(n13250) );
  OR2_X1 U10503 ( .A1(n8657), .A2(n8656), .ZN(n8658) );
  NAND2_X1 U10504 ( .A1(n8659), .A2(n8658), .ZN(n10229) );
  OR2_X1 U10505 ( .A1(n10229), .A2(n7220), .ZN(n8667) );
  NAND2_X1 U10506 ( .A1(n8780), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8663) );
  AOI22_X1 U10507 ( .A1(n8665), .A2(SI_19_), .B1(n8664), .B2(n13419), .ZN(
        n8666) );
  NAND2_X1 U10508 ( .A1(n8520), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8674) );
  NAND2_X1 U10509 ( .A1(n12552), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8673) );
  NAND2_X1 U10510 ( .A1(n8668), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8670) );
  INV_X1 U10511 ( .A(n8669), .ZN(n8679) );
  NAND2_X1 U10512 ( .A1(n8670), .A2(n8679), .ZN(n13569) );
  NAND2_X1 U10513 ( .A1(n8524), .A2(n13569), .ZN(n8672) );
  NAND2_X1 U10514 ( .A1(n8759), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8671) );
  NAND4_X1 U10515 ( .A1(n8674), .A2(n8673), .A3(n8672), .A4(n8671), .ZN(n13249) );
  NOR2_X1 U10516 ( .A1(n13713), .A2(n13249), .ZN(n8675) );
  INV_X1 U10517 ( .A(n13713), .ZN(n13143) );
  XNOR2_X1 U10518 ( .A(n8676), .B(n11666), .ZN(n10629) );
  NAND2_X1 U10519 ( .A1(n10629), .A2(n12560), .ZN(n8678) );
  OR2_X1 U10520 ( .A1(n7221), .A2(n11729), .ZN(n8677) );
  NAND2_X1 U10521 ( .A1(n7223), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8684) );
  NAND2_X1 U10522 ( .A1(n8759), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8683) );
  NAND2_X1 U10523 ( .A1(P3_REG3_REG_20__SCAN_IN), .A2(n8679), .ZN(n8680) );
  NAND2_X1 U10524 ( .A1(n8680), .A2(n8691), .ZN(n13555) );
  NAND2_X1 U10525 ( .A1(n8543), .A2(n13555), .ZN(n8682) );
  NAND2_X1 U10526 ( .A1(n12552), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8681) );
  NAND2_X1 U10527 ( .A1(n13554), .A2(n13568), .ZN(n12706) );
  NAND2_X1 U10528 ( .A1(n12705), .A2(n12706), .ZN(n12588) );
  NAND2_X1 U10529 ( .A1(n13547), .A2(n12588), .ZN(n8686) );
  INV_X1 U10530 ( .A(n13568), .ZN(n13248) );
  NAND2_X1 U10531 ( .A1(n13554), .A2(n13248), .ZN(n8685) );
  XNOR2_X1 U10532 ( .A(n8688), .B(n8687), .ZN(n10748) );
  NAND2_X1 U10533 ( .A1(n10748), .A2(n12560), .ZN(n8690) );
  INV_X1 U10534 ( .A(SI_21_), .ZN(n10749) );
  NAND2_X1 U10535 ( .A1(n8520), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8696) );
  NAND2_X1 U10536 ( .A1(n12552), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8695) );
  NAND2_X1 U10537 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(n8691), .ZN(n8692) );
  NAND2_X1 U10538 ( .A1(n8703), .A2(n8692), .ZN(n13540) );
  NAND2_X1 U10539 ( .A1(n8543), .A2(n13540), .ZN(n8694) );
  NAND2_X1 U10540 ( .A1(n8759), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8693) );
  NAND4_X1 U10541 ( .A1(n8696), .A2(n8695), .A3(n8694), .A4(n8693), .ZN(n13247) );
  AND2_X1 U10542 ( .A1(n13539), .A2(n13247), .ZN(n8697) );
  OR2_X1 U10543 ( .A1(n13539), .A2(n13247), .ZN(n8698) );
  XNOR2_X1 U10544 ( .A(n8700), .B(n8699), .ZN(n10759) );
  NAND2_X1 U10545 ( .A1(n10759), .A2(n12560), .ZN(n8702) );
  OR2_X1 U10546 ( .A1(n7221), .A2(n9443), .ZN(n8701) );
  NAND2_X1 U10547 ( .A1(n7223), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8708) );
  NAND2_X1 U10548 ( .A1(n12552), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8707) );
  NAND2_X1 U10549 ( .A1(n8703), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U10550 ( .A1(n8714), .A2(n8704), .ZN(n13526) );
  NAND2_X1 U10551 ( .A1(n8543), .A2(n13526), .ZN(n8706) );
  NAND2_X1 U10552 ( .A1(n8759), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8705) );
  NAND4_X1 U10553 ( .A1(n8708), .A2(n8707), .A3(n8706), .A4(n8705), .ZN(n13509) );
  NOR2_X1 U10554 ( .A1(n13525), .A2(n13509), .ZN(n8709) );
  XNOR2_X1 U10555 ( .A(n8711), .B(n8710), .ZN(n10882) );
  NAND2_X1 U10556 ( .A1(n10882), .A2(n12560), .ZN(n8713) );
  NAND2_X1 U10557 ( .A1(n12552), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U10558 ( .A1(n7223), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8718) );
  NAND2_X1 U10559 ( .A1(n8714), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U10560 ( .A1(n8725), .A2(n8715), .ZN(n13515) );
  NAND2_X1 U10561 ( .A1(n8543), .A2(n13515), .ZN(n8717) );
  NAND2_X1 U10562 ( .A1(n8759), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8716) );
  NAND2_X1 U10563 ( .A1(n13514), .A2(n13522), .ZN(n12718) );
  NAND2_X1 U10564 ( .A1(n12717), .A2(n12718), .ZN(n13513) );
  NAND2_X1 U10565 ( .A1(n13506), .A2(n13513), .ZN(n8721) );
  INV_X1 U10566 ( .A(n13522), .ZN(n13246) );
  NAND2_X1 U10567 ( .A1(n13514), .A2(n13246), .ZN(n8720) );
  XNOR2_X1 U10568 ( .A(n8722), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n11231) );
  NAND2_X1 U10569 ( .A1(n11231), .A2(n12560), .ZN(n8724) );
  NAND2_X1 U10570 ( .A1(n12552), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8730) );
  NAND2_X1 U10571 ( .A1(n8520), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8729) );
  NAND2_X1 U10572 ( .A1(n8725), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8726) );
  NAND2_X1 U10573 ( .A1(n8738), .A2(n8726), .ZN(n13500) );
  NAND2_X1 U10574 ( .A1(n8543), .A2(n13500), .ZN(n8728) );
  NAND2_X1 U10575 ( .A1(n8759), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8727) );
  NAND4_X1 U10576 ( .A1(n8730), .A2(n8729), .A3(n8728), .A4(n8727), .ZN(n13508) );
  AND2_X1 U10577 ( .A1(n13181), .A2(n13508), .ZN(n8731) );
  OR2_X1 U10578 ( .A1(n8733), .A2(n8732), .ZN(n8734) );
  NAND2_X1 U10579 ( .A1(n8735), .A2(n8734), .ZN(n11329) );
  INV_X1 U10580 ( .A(SI_25_), .ZN(n11713) );
  NAND2_X1 U10581 ( .A1(n12552), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U10582 ( .A1(n7223), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8742) );
  NAND2_X1 U10583 ( .A1(n8738), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8739) );
  NAND2_X1 U10584 ( .A1(n8756), .A2(n8739), .ZN(n13487) );
  NAND2_X1 U10585 ( .A1(n8543), .A2(n13487), .ZN(n8741) );
  NAND2_X1 U10586 ( .A1(n8759), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8740) );
  NAND2_X1 U10587 ( .A1(n13688), .A2(n13495), .ZN(n13468) );
  XNOR2_X1 U10588 ( .A(n8745), .B(n8744), .ZN(n11628) );
  NAND2_X1 U10589 ( .A1(n11628), .A2(n12560), .ZN(n8747) );
  NAND2_X1 U10590 ( .A1(n7223), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8751) );
  NAND2_X1 U10591 ( .A1(n12552), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8750) );
  XNOR2_X1 U10592 ( .A(n8756), .B(P3_REG3_REG_26__SCAN_IN), .ZN(n13472) );
  NAND2_X1 U10593 ( .A1(n8543), .A2(n13472), .ZN(n8749) );
  NAND2_X1 U10594 ( .A1(n8759), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8748) );
  NAND4_X1 U10595 ( .A1(n8751), .A2(n8750), .A3(n8749), .A4(n8748), .ZN(n13483) );
  OR2_X1 U10596 ( .A1(n13478), .A2(n7263), .ZN(n13449) );
  XNOR2_X1 U10597 ( .A(n8753), .B(n8752), .ZN(n12030) );
  NAND2_X1 U10598 ( .A1(n12030), .A2(n12560), .ZN(n8755) );
  INV_X1 U10599 ( .A(SI_27_), .ZN(n12031) );
  NAND2_X2 U10600 ( .A1(n8755), .A2(n8754), .ZN(n13680) );
  NAND2_X1 U10601 ( .A1(n12552), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8763) );
  NAND2_X1 U10602 ( .A1(n7223), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8762) );
  OAI21_X1 U10603 ( .B1(n8756), .B2(P3_REG3_REG_26__SCAN_IN), .A(
        P3_REG3_REG_27__SCAN_IN), .ZN(n8758) );
  NAND2_X1 U10604 ( .A1(n8758), .A2(n8757), .ZN(n13458) );
  NAND2_X1 U10605 ( .A1(n8543), .A2(n13458), .ZN(n8761) );
  NAND2_X1 U10606 ( .A1(n8759), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8760) );
  OR2_X1 U10607 ( .A1(n13449), .A2(n7264), .ZN(n8768) );
  NAND2_X1 U10608 ( .A1(n13680), .A2(n13467), .ZN(n12604) );
  INV_X1 U10609 ( .A(n13454), .ZN(n8766) );
  INV_X1 U10610 ( .A(n13495), .ZN(n13245) );
  NAND2_X1 U10611 ( .A1(n13688), .A2(n13245), .ZN(n13464) );
  NAND2_X1 U10612 ( .A1(n13217), .A2(n13483), .ZN(n8764) );
  AND2_X1 U10613 ( .A1(n13464), .A2(n8764), .ZN(n8765) );
  OR2_X1 U10614 ( .A1(n7263), .A2(n8765), .ZN(n13450) );
  AND2_X1 U10615 ( .A1(n8766), .A2(n13450), .ZN(n13451) );
  OR2_X1 U10616 ( .A1(n7264), .A2(n13451), .ZN(n8767) );
  OAI21_X1 U10617 ( .B1(n13479), .B2(n8768), .A(n8767), .ZN(n13438) );
  NAND2_X1 U10618 ( .A1(n13116), .A2(n13456), .ZN(n12729) );
  NAND2_X1 U10619 ( .A1(n13438), .A2(n13437), .ZN(n13436) );
  OAI21_X1 U10620 ( .B1(n13456), .B2(n13752), .A(n13436), .ZN(n8779) );
  INV_X1 U10621 ( .A(n8769), .ZN(n8770) );
  INV_X1 U10622 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15198) );
  XNOR2_X1 U10623 ( .A(n15198), .B(P1_DATAO_REG_29__SCAN_IN), .ZN(n12541) );
  XNOR2_X1 U10624 ( .A(n12543), .B(n12541), .ZN(n13809) );
  NAND2_X1 U10625 ( .A1(n13809), .A2(n12560), .ZN(n8774) );
  INV_X1 U10626 ( .A(SI_29_), .ZN(n13811) );
  OR2_X1 U10627 ( .A1(n7221), .A2(n13811), .ZN(n8773) );
  NAND2_X1 U10628 ( .A1(n8774), .A2(n8773), .ZN(n8858) );
  INV_X1 U10629 ( .A(n13424), .ZN(n8775) );
  NAND2_X1 U10630 ( .A1(n8543), .A2(n8775), .ZN(n12556) );
  NAND2_X1 U10631 ( .A1(n12552), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8778) );
  NAND2_X1 U10632 ( .A1(n7223), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U10633 ( .A1(n8759), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8776) );
  OR2_X1 U10634 ( .A1(n8858), .A2(n13439), .ZN(n12736) );
  NAND2_X1 U10635 ( .A1(n8858), .A2(n13439), .ZN(n12735) );
  NAND2_X1 U10636 ( .A1(n12736), .A2(n12735), .ZN(n12732) );
  XNOR2_X1 U10637 ( .A(n8779), .B(n12732), .ZN(n8795) );
  XNOR2_X2 U10638 ( .A(n8783), .B(n8782), .ZN(n12602) );
  NAND2_X1 U10639 ( .A1(n12612), .A2(n12749), .ZN(n8786) );
  NAND2_X1 U10640 ( .A1(n8784), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8785) );
  NAND2_X1 U10641 ( .A1(n13419), .A2(n12754), .ZN(n8862) );
  INV_X1 U10642 ( .A(n8787), .ZN(n12751) );
  INV_X1 U10643 ( .A(n8788), .ZN(n10129) );
  NAND2_X1 U10644 ( .A1(n12751), .A2(n10129), .ZN(n10128) );
  NAND2_X1 U10645 ( .A1(n10126), .A2(n10128), .ZN(n10624) );
  AND2_X1 U10646 ( .A1(n12751), .A2(P3_B_REG_SCAN_IN), .ZN(n8789) );
  OR2_X1 U10647 ( .A1(n15723), .A2(n8789), .ZN(n13422) );
  NAND2_X1 U10648 ( .A1(n12552), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8792) );
  NAND2_X1 U10649 ( .A1(n7223), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8791) );
  NAND2_X1 U10650 ( .A1(n8759), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8790) );
  AND4_X1 U10651 ( .A1(n12556), .A2(n8792), .A3(n8791), .A4(n8790), .ZN(n12565) );
  INV_X1 U10652 ( .A(n8793), .ZN(n8794) );
  INV_X1 U10653 ( .A(n12575), .ZN(n11054) );
  NAND2_X1 U10654 ( .A1(n11996), .A2(n11639), .ZN(n8797) );
  NOR2_X1 U10655 ( .A1(n7907), .A2(n15870), .ZN(n12654) );
  NAND2_X1 U10656 ( .A1(n7907), .A2(n15870), .ZN(n12656) );
  INV_X1 U10657 ( .A(n12658), .ZN(n8799) );
  INV_X1 U10658 ( .A(n13254), .ZN(n12246) );
  NAND2_X1 U10659 ( .A1(n12246), .A2(n15892), .ZN(n8798) );
  NAND2_X1 U10660 ( .A1(n12164), .A2(n8800), .ZN(n12666) );
  NAND2_X1 U10661 ( .A1(n13253), .A2(n15910), .ZN(n12668) );
  NAND2_X1 U10662 ( .A1(n13657), .A2(n12316), .ZN(n12672) );
  NAND2_X1 U10663 ( .A1(n13252), .A2(n15934), .ZN(n12670) );
  OR2_X1 U10664 ( .A1(n13793), .A2(n13627), .ZN(n12681) );
  INV_X1 U10665 ( .A(n13561), .ZN(n8804) );
  NAND2_X1 U10666 ( .A1(n13713), .A2(n13580), .ZN(n12702) );
  NAND2_X1 U10667 ( .A1(n12693), .A2(n13575), .ZN(n13562) );
  NAND2_X1 U10668 ( .A1(n13562), .A2(n13561), .ZN(n8803) );
  AND2_X1 U10669 ( .A1(n12702), .A2(n8803), .ZN(n12698) );
  NAND2_X1 U10670 ( .A1(n13539), .A2(n13548), .ZN(n12710) );
  NAND2_X1 U10671 ( .A1(n8806), .A2(n12709), .ZN(n13523) );
  XNOR2_X1 U10672 ( .A(n13525), .B(n13509), .ZN(n13524) );
  INV_X1 U10673 ( .A(n13509), .ZN(n13534) );
  OR2_X1 U10674 ( .A1(n13525), .A2(n13534), .ZN(n8807) );
  NAND2_X1 U10675 ( .A1(n13181), .A2(n13486), .ZN(n8808) );
  INV_X1 U10676 ( .A(n13483), .ZN(n13457) );
  NAND2_X1 U10677 ( .A1(n13217), .A2(n13457), .ZN(n12572) );
  AND2_X1 U10678 ( .A1(n12572), .A2(n13468), .ZN(n12606) );
  INV_X1 U10679 ( .A(n12607), .ZN(n8812) );
  NAND2_X1 U10680 ( .A1(n10751), .A2(n12602), .ZN(n8851) );
  XNOR2_X1 U10681 ( .A(n8851), .B(n12754), .ZN(n8813) );
  NAND2_X1 U10682 ( .A1(n10751), .A2(n13407), .ZN(n12594) );
  NAND2_X1 U10683 ( .A1(n8813), .A2(n12594), .ZN(n10345) );
  INV_X1 U10684 ( .A(n10617), .ZN(n12744) );
  AND2_X1 U10685 ( .A1(n15935), .A2(n12744), .ZN(n8814) );
  NAND2_X1 U10686 ( .A1(n10345), .A2(n8814), .ZN(n8815) );
  NAND2_X1 U10687 ( .A1(n10617), .A2(n8862), .ZN(n8852) );
  NAND2_X1 U10688 ( .A1(n8816), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8817) );
  XNOR2_X1 U10689 ( .A(n11232), .B(P3_B_REG_SCAN_IN), .ZN(n8822) );
  NAND2_X1 U10690 ( .A1(n7298), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8821) );
  INV_X1 U10691 ( .A(n8827), .ZN(n8824) );
  INV_X1 U10692 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8823) );
  NAND2_X1 U10693 ( .A1(n8824), .A2(n8823), .ZN(n8826) );
  INV_X1 U10694 ( .A(n8833), .ZN(n11630) );
  NAND2_X1 U10695 ( .A1(n11630), .A2(n11232), .ZN(n8825) );
  NAND2_X1 U10696 ( .A1(n11630), .A2(n11328), .ZN(n8828) );
  NAND2_X1 U10697 ( .A1(n10615), .A2(n10588), .ZN(n8865) );
  INV_X1 U10698 ( .A(n11328), .ZN(n8831) );
  INV_X1 U10699 ( .A(n11232), .ZN(n8830) );
  NAND2_X1 U10700 ( .A1(n7923), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8835) );
  NOR2_X1 U10701 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n8839) );
  NOR4_X1 U10702 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n8838) );
  NOR4_X1 U10703 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8837) );
  NOR4_X1 U10704 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8836) );
  NAND4_X1 U10705 ( .A1(n8839), .A2(n8838), .A3(n8837), .A4(n8836), .ZN(n8845)
         );
  NOR4_X1 U10706 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8843) );
  NOR4_X1 U10707 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n8842) );
  NOR4_X1 U10708 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n8841) );
  NOR4_X1 U10709 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n8840) );
  NAND4_X1 U10710 ( .A1(n8843), .A2(n8842), .A3(n8841), .A4(n8840), .ZN(n8844)
         );
  NOR2_X1 U10711 ( .A1(n8845), .A2(n8844), .ZN(n8846) );
  OR2_X1 U10712 ( .A1(n8827), .A2(n8846), .ZN(n8863) );
  AND2_X1 U10713 ( .A1(n10355), .A2(n8863), .ZN(n8847) );
  AND3_X1 U10714 ( .A1(n8860), .A2(n8865), .A3(n8847), .ZN(n10591) );
  INV_X1 U10715 ( .A(n10588), .ZN(n13797) );
  NAND2_X1 U10716 ( .A1(n8848), .A2(n12738), .ZN(n10587) );
  OR2_X1 U10717 ( .A1(n12738), .A2(n12744), .ZN(n10590) );
  NAND2_X1 U10718 ( .A1(n10587), .A2(n10590), .ZN(n8849) );
  NAND2_X1 U10719 ( .A1(n13797), .A2(n8849), .ZN(n8855) );
  AOI22_X1 U10720 ( .A1(n10751), .A2(n8852), .B1(n8851), .B2(n8850), .ZN(n8853) );
  NAND2_X1 U10721 ( .A1(n10588), .A2(n8853), .ZN(n8854) );
  MUX2_X1 U10722 ( .A(n8857), .B(n8869), .S(n15940), .Z(n8859) );
  NAND2_X1 U10723 ( .A1(n8859), .A2(n8257), .ZN(P3_U3488) );
  INV_X1 U10724 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8870) );
  INV_X1 U10725 ( .A(n8860), .ZN(n8861) );
  NAND2_X1 U10726 ( .A1(n8861), .A2(n8863), .ZN(n10353) );
  OR2_X1 U10727 ( .A1(n12738), .A2(n10617), .ZN(n10342) );
  OR3_X1 U10728 ( .A1(n12612), .A2(n12602), .A3(n8862), .ZN(n10346) );
  AND2_X1 U10729 ( .A1(n10342), .A2(n10346), .ZN(n8867) );
  INV_X1 U10730 ( .A(n8863), .ZN(n8864) );
  INV_X1 U10731 ( .A(n10345), .ZN(n8866) );
  OAI22_X1 U10732 ( .A1(n10353), .A2(n8867), .B1(n10350), .B2(n8866), .ZN(
        n8868) );
  MUX2_X1 U10733 ( .A(n8870), .B(n8869), .S(n15944), .Z(n8871) );
  NAND2_X1 U10734 ( .A1(n8871), .A2(n8258), .ZN(P3_U3456) );
  NOR2_X1 U10735 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .ZN(n8875) );
  NOR2_X1 U10736 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8874) );
  NOR2_X1 U10737 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), 
        .ZN(n8873) );
  NOR2_X1 U10738 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n8876) );
  INV_X1 U10739 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8880) );
  NAND2_X2 U10740 ( .A1(n8886), .A2(n8885), .ZN(n15200) );
  NAND2_X1 U10741 ( .A1(n9056), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8893) );
  INV_X1 U10742 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9954) );
  OR2_X1 U10743 ( .A1(n9031), .A2(n9954), .ZN(n8892) );
  INV_X1 U10744 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10511) );
  OR2_X1 U10745 ( .A1(n8994), .A2(n10511), .ZN(n8891) );
  NAND2_X4 U10746 ( .A1(n8888), .A2(n15200), .ZN(n9546) );
  INV_X1 U10747 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n8889) );
  NAND2_X1 U10748 ( .A1(n8894), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8895) );
  OR2_X2 U10749 ( .A1(n8901), .A2(SI_1_), .ZN(n8942) );
  INV_X1 U10750 ( .A(SI_0_), .ZN(n8957) );
  NAND2_X1 U10751 ( .A1(n8901), .A2(SI_1_), .ZN(n8972) );
  INV_X1 U10752 ( .A(SI_2_), .ZN(n9911) );
  NAND3_X1 U10753 ( .A1(n8902), .A2(n8972), .A3(n9911), .ZN(n8906) );
  INV_X1 U10754 ( .A(n8972), .ZN(n8903) );
  NAND2_X1 U10755 ( .A1(n8903), .A2(SI_2_), .ZN(n8905) );
  NAND2_X1 U10756 ( .A1(n8942), .A2(SI_2_), .ZN(n8904) );
  MUX2_X1 U10757 ( .A(n9844), .B(n10446), .S(n9288), .Z(n8975) );
  XNOR2_X1 U10758 ( .A(n8976), .B(n8975), .ZN(n10449) );
  NAND2_X2 U10759 ( .A1(n8959), .A2(n10404), .ZN(n9104) );
  NAND2_X1 U10760 ( .A1(n9571), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8912) );
  INV_X1 U10761 ( .A(n8907), .ZN(n8947) );
  NAND2_X1 U10762 ( .A1(n8947), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8908) );
  MUX2_X1 U10763 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8908), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n8910) );
  NAND2_X1 U10764 ( .A1(n8910), .A2(n8982), .ZN(n9953) );
  INV_X1 U10765 ( .A(n9953), .ZN(n10118) );
  NAND2_X1 U10766 ( .A1(n9349), .A2(n10118), .ZN(n8911) );
  NAND2_X1 U10767 ( .A1(n10604), .A2(n15739), .ZN(n9623) );
  NAND3_X1 U10768 ( .A1(n8919), .A2(n8918), .A3(n8917), .ZN(n8920) );
  INV_X1 U10769 ( .A(n9577), .ZN(n8927) );
  NAND2_X1 U10770 ( .A1(n8931), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8925) );
  MUX2_X1 U10771 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8925), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n8926) );
  NAND2_X1 U10772 ( .A1(n8927), .A2(n12052), .ZN(n8934) );
  INV_X1 U10773 ( .A(n8928), .ZN(n8929) );
  NAND2_X1 U10774 ( .A1(n8929), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8930) );
  MUX2_X1 U10775 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8930), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n8932) );
  AND2_X2 U10776 ( .A1(n8934), .A2(n8933), .ZN(n9267) );
  INV_X1 U10777 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n8935) );
  OR2_X1 U10778 ( .A1(n8994), .A2(n8935), .ZN(n8937) );
  INV_X1 U10779 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9951) );
  AND2_X1 U10780 ( .A1(n8937), .A2(n8936), .ZN(n8941) );
  INV_X1 U10781 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n8938) );
  NAND2_X1 U10782 ( .A1(n9056), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8939) );
  NAND3_X2 U10783 ( .A1(n8941), .A2(n8940), .A3(n8939), .ZN(n9700) );
  INV_X2 U10784 ( .A(n9700), .ZN(n10431) );
  NAND2_X1 U10785 ( .A1(n9571), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8950) );
  NAND2_X1 U10786 ( .A1(n8944), .A2(n7511), .ZN(n8945) );
  NAND2_X1 U10787 ( .A1(n8971), .A2(n8945), .ZN(n10397) );
  NAND2_X1 U10788 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8946) );
  MUX2_X1 U10789 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8946), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n8948) );
  NAND2_X1 U10790 ( .A1(n8948), .A2(n8947), .ZN(n9950) );
  INV_X1 U10791 ( .A(n9950), .ZN(n14757) );
  INV_X1 U10792 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8951) );
  NAND2_X1 U10793 ( .A1(n9056), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8954) );
  INV_X1 U10794 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9886) );
  NOR2_X1 U10795 ( .A1(n10404), .A2(n8957), .ZN(n8958) );
  XNOR2_X1 U10796 ( .A(n8958), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n15219) );
  MUX2_X1 U10797 ( .A(n9886), .B(n15219), .S(n9891), .Z(n15679) );
  NAND3_X1 U10798 ( .A1(n10503), .A2(n9624), .A3(n9702), .ZN(n8964) );
  NAND2_X1 U10799 ( .A1(n14750), .A2(n15679), .ZN(n9625) );
  INV_X1 U10800 ( .A(n9625), .ZN(n8960) );
  NAND2_X1 U10801 ( .A1(n8960), .A2(n9700), .ZN(n8963) );
  NAND2_X1 U10802 ( .A1(n9625), .A2(n10431), .ZN(n8961) );
  NAND2_X1 U10803 ( .A1(n8961), .A2(n9699), .ZN(n8962) );
  NAND4_X1 U10804 ( .A1(n8965), .A2(n8964), .A3(n8963), .A4(n8962), .ZN(n8993)
         );
  INV_X4 U10805 ( .A(n9267), .ZN(n9606) );
  INV_X1 U10806 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n8966) );
  OR2_X1 U10807 ( .A1(n9546), .A2(n8966), .ZN(n8970) );
  NAND2_X1 U10808 ( .A1(n9056), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8969) );
  INV_X1 U10809 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9955) );
  OR2_X1 U10810 ( .A1(n9031), .A2(n9955), .ZN(n8968) );
  OR2_X1 U10811 ( .A1(n8994), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8967) );
  INV_X1 U10812 ( .A(n8977), .ZN(n8978) );
  OR2_X1 U10813 ( .A1(n8979), .A2(n8978), .ZN(n8980) );
  NAND2_X1 U10814 ( .A1(n8982), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8981) );
  MUX2_X1 U10815 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8981), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n8983) );
  INV_X1 U10816 ( .A(n14766), .ZN(n8984) );
  NOR2_X1 U10817 ( .A1(n14749), .A2(n10658), .ZN(n9798) );
  NAND2_X1 U10818 ( .A1(n9700), .A2(n9699), .ZN(n9622) );
  NAND2_X1 U10819 ( .A1(n8988), .A2(n9622), .ZN(n8989) );
  NAND2_X1 U10820 ( .A1(n10146), .A2(n10514), .ZN(n9814) );
  NAND4_X1 U10821 ( .A1(n8989), .A2(n9606), .A3(n9814), .A4(n10503), .ZN(n8991) );
  NAND4_X1 U10822 ( .A1(n8993), .A2(n8992), .A3(n8991), .A4(n8990), .ZN(n9011)
         );
  AND2_X1 U10823 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9027) );
  INV_X1 U10824 ( .A(n9027), .ZN(n9029) );
  OAI21_X1 U10825 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9029), .ZN(n10949) );
  NAND2_X1 U10826 ( .A1(n9056), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8998) );
  INV_X1 U10827 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9958) );
  OR2_X1 U10828 ( .A1(n9031), .A2(n9958), .ZN(n8997) );
  INV_X1 U10829 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n8995) );
  OR2_X1 U10830 ( .A1(n9546), .A2(n8995), .ZN(n8996) );
  NAND2_X1 U10831 ( .A1(n9002), .A2(SI_4_), .ZN(n9015) );
  OAI21_X1 U10832 ( .B1(n9002), .B2(SI_4_), .A(n9015), .ZN(n9003) );
  INV_X1 U10833 ( .A(n9003), .ZN(n9004) );
  OR2_X1 U10834 ( .A1(n9005), .A2(n9004), .ZN(n9006) );
  NAND2_X1 U10835 ( .A1(n9595), .A2(n10534), .ZN(n9008) );
  NAND2_X1 U10836 ( .A1(n9349), .A2(n14782), .ZN(n9007) );
  OAI211_X2 U10837 ( .C1(n9104), .C2(n9852), .A(n9008), .B(n9007), .ZN(n10946)
         );
  XNOR2_X1 U10838 ( .A(n14748), .B(n10946), .ZN(n9621) );
  INV_X1 U10839 ( .A(n14749), .ZN(n10430) );
  INV_X1 U10840 ( .A(n10658), .ZN(n15756) );
  OAI21_X1 U10841 ( .B1(n10430), .B2(n15756), .A(n9009), .ZN(n9010) );
  NAND3_X1 U10842 ( .A1(n9011), .A2(n9621), .A3(n9010), .ZN(n9014) );
  AOI21_X1 U10843 ( .B1(n10607), .B2(n9538), .A(n10691), .ZN(n9013) );
  AOI21_X1 U10844 ( .B1(n14748), .B2(n9606), .A(n10946), .ZN(n9012) );
  MUX2_X1 U10845 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9288), .Z(n9017) );
  NAND2_X1 U10846 ( .A1(n9017), .A2(SI_5_), .ZN(n9041) );
  OAI21_X1 U10847 ( .B1(n9017), .B2(SI_5_), .A(n9041), .ZN(n9018) );
  INV_X1 U10848 ( .A(n9018), .ZN(n9019) );
  INV_X1 U10849 ( .A(n9021), .ZN(n9023) );
  INV_X1 U10850 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9022) );
  NAND2_X1 U10851 ( .A1(n9023), .A2(n9022), .ZN(n9048) );
  NAND2_X1 U10852 ( .A1(n9048), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9024) );
  XNOR2_X1 U10853 ( .A(n9024), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9961) );
  AOI22_X1 U10854 ( .A1(n9596), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9349), .B2(
        n9961), .ZN(n9025) );
  NAND2_X1 U10855 ( .A1(n9026), .A2(n9025), .ZN(n15795) );
  INV_X1 U10856 ( .A(n9052), .ZN(n9054) );
  INV_X1 U10857 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U10858 ( .A1(n9029), .A2(n9028), .ZN(n9030) );
  NAND2_X1 U10859 ( .A1(n9054), .A2(n9030), .ZN(n10803) );
  OR2_X1 U10860 ( .A1(n9542), .A2(n10803), .ZN(n9037) );
  NAND2_X1 U10861 ( .A1(n9056), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9036) );
  INV_X1 U10862 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9032) );
  OR2_X1 U10863 ( .A1(n9544), .A2(n9032), .ZN(n9035) );
  INV_X1 U10864 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9033) );
  OR2_X1 U10865 ( .A1(n9546), .A2(n9033), .ZN(n9034) );
  MUX2_X1 U10866 ( .A(n15795), .B(n14747), .S(n9606), .Z(n9039) );
  MUX2_X1 U10867 ( .A(n14747), .B(n15795), .S(n9606), .Z(n9038) );
  NAND2_X1 U10868 ( .A1(n9043), .A2(SI_6_), .ZN(n9078) );
  OAI21_X1 U10869 ( .B1(SI_6_), .B2(n9043), .A(n9078), .ZN(n9044) );
  INV_X1 U10870 ( .A(n9044), .ZN(n9045) );
  OR2_X1 U10871 ( .A1(n10565), .A2(n9209), .ZN(n9051) );
  OR2_X1 U10872 ( .A1(n9048), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9081) );
  NAND2_X1 U10873 ( .A1(n9081), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9049) );
  XNOR2_X1 U10874 ( .A(n9049), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9963) );
  AOI22_X1 U10875 ( .A1(n9596), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9349), .B2(
        n9963), .ZN(n9050) );
  NAND2_X1 U10876 ( .A1(n9052), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9071) );
  INV_X1 U10877 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9053) );
  NAND2_X1 U10878 ( .A1(n9054), .A2(n9053), .ZN(n9055) );
  NAND2_X1 U10879 ( .A1(n9071), .A2(n9055), .ZN(n10996) );
  OR2_X1 U10880 ( .A1(n9542), .A2(n10996), .ZN(n9061) );
  NAND2_X1 U10881 ( .A1(n9056), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9060) );
  INV_X1 U10882 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9962) );
  OR2_X1 U10883 ( .A1(n9544), .A2(n9962), .ZN(n9059) );
  INV_X1 U10884 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9057) );
  OR2_X1 U10885 ( .A1(n9546), .A2(n9057), .ZN(n9058) );
  NAND4_X1 U10886 ( .A1(n9061), .A2(n9060), .A3(n9059), .A4(n9058), .ZN(n14746) );
  MUX2_X1 U10887 ( .A(n10995), .B(n14746), .S(n9538), .Z(n9065) );
  NAND2_X1 U10888 ( .A1(n9064), .A2(n9065), .ZN(n9063) );
  MUX2_X1 U10889 ( .A(n10995), .B(n14746), .S(n9606), .Z(n9062) );
  NAND2_X1 U10890 ( .A1(n9063), .A2(n9062), .ZN(n9069) );
  INV_X1 U10891 ( .A(n9064), .ZN(n9067) );
  INV_X1 U10892 ( .A(n9065), .ZN(n9066) );
  NAND2_X1 U10893 ( .A1(n9067), .A2(n9066), .ZN(n9068) );
  INV_X1 U10894 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9070) );
  NOR2_X1 U10895 ( .A1(n9071), .A2(n9070), .ZN(n9088) );
  INV_X1 U10896 ( .A(n9088), .ZN(n9090) );
  NAND2_X1 U10897 ( .A1(n9071), .A2(n9070), .ZN(n9072) );
  NAND2_X1 U10898 ( .A1(n9090), .A2(n9072), .ZN(n11156) );
  OR2_X1 U10899 ( .A1(n9542), .A2(n11156), .ZN(n9077) );
  NAND2_X1 U10900 ( .A1(n9056), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9076) );
  INV_X1 U10901 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10006) );
  OR2_X1 U10902 ( .A1(n9544), .A2(n10006), .ZN(n9075) );
  INV_X1 U10903 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9073) );
  OR2_X1 U10904 ( .A1(n9546), .A2(n9073), .ZN(n9074) );
  NAND4_X1 U10905 ( .A1(n9077), .A2(n9076), .A3(n9075), .A4(n9074), .ZN(n14745) );
  NAND2_X1 U10906 ( .A1(n9080), .A2(SI_7_), .ZN(n9098) );
  NAND2_X1 U10907 ( .A1(n10726), .A2(n9595), .ZN(n9084) );
  OAI21_X1 U10908 ( .B1(n9081), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9082) );
  XNOR2_X1 U10909 ( .A(n9082), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10003) );
  AOI22_X1 U10910 ( .A1(n9596), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9349), .B2(
        n10003), .ZN(n9083) );
  NAND2_X2 U10911 ( .A1(n9084), .A2(n9083), .ZN(n15836) );
  MUX2_X1 U10912 ( .A(n14745), .B(n15836), .S(n9267), .Z(n9086) );
  MUX2_X1 U10913 ( .A(n14745), .B(n15836), .S(n9606), .Z(n9085) );
  INV_X1 U10914 ( .A(n9086), .ZN(n9087) );
  NAND2_X1 U10915 ( .A1(n9088), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9115) );
  INV_X1 U10916 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9089) );
  NAND2_X1 U10917 ( .A1(n9090), .A2(n9089), .ZN(n9091) );
  NAND2_X1 U10918 ( .A1(n9115), .A2(n9091), .ZN(n11217) );
  OR2_X1 U10919 ( .A1(n9542), .A2(n11217), .ZN(n9096) );
  NAND2_X1 U10920 ( .A1(n9056), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9095) );
  INV_X1 U10921 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10008) );
  OR2_X1 U10922 ( .A1(n9544), .A2(n10008), .ZN(n9094) );
  INV_X1 U10923 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9092) );
  OR2_X1 U10924 ( .A1(n9546), .A2(n9092), .ZN(n9093) );
  NAND4_X1 U10925 ( .A1(n9096), .A2(n9095), .A3(n9094), .A4(n9093), .ZN(n14744) );
  MUX2_X1 U10926 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9288), .Z(n9099) );
  NAND2_X1 U10927 ( .A1(n9099), .A2(SI_8_), .ZN(n9122) );
  OAI21_X1 U10928 ( .B1(SI_8_), .B2(n9099), .A(n9122), .ZN(n9100) );
  INV_X1 U10929 ( .A(n9100), .ZN(n9101) );
  OR2_X1 U10930 ( .A1(n9102), .A2(n9101), .ZN(n9103) );
  NAND2_X1 U10931 ( .A1(n9123), .A2(n9103), .ZN(n10911) );
  OR2_X1 U10932 ( .A1(n10911), .A2(n9209), .ZN(n9110) );
  INV_X1 U10933 ( .A(n9105), .ZN(n9107) );
  NAND2_X1 U10934 ( .A1(n9107), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9108) );
  XNOR2_X1 U10935 ( .A(n9108), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10024) );
  AOI22_X1 U10936 ( .A1(n9596), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9349), .B2(
        n10024), .ZN(n9109) );
  NAND2_X1 U10937 ( .A1(n9110), .A2(n9109), .ZN(n11377) );
  MUX2_X1 U10938 ( .A(n14744), .B(n11377), .S(n9606), .Z(n9112) );
  MUX2_X1 U10939 ( .A(n14744), .B(n11377), .S(n9267), .Z(n9111) );
  INV_X1 U10940 ( .A(n9112), .ZN(n9113) );
  INV_X1 U10941 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9114) );
  NAND2_X1 U10942 ( .A1(n9115), .A2(n9114), .ZN(n9116) );
  NAND2_X1 U10943 ( .A1(n9144), .A2(n9116), .ZN(n11387) );
  OR2_X1 U10944 ( .A1(n9542), .A2(n11387), .ZN(n9121) );
  NAND2_X1 U10945 ( .A1(n9301), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9120) );
  OR2_X1 U10946 ( .A1(n9544), .A2(n10025), .ZN(n9119) );
  INV_X1 U10947 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9117) );
  OR2_X1 U10948 ( .A1(n9546), .A2(n9117), .ZN(n9118) );
  NAND4_X1 U10949 ( .A1(n9121), .A2(n9120), .A3(n9119), .A4(n9118), .ZN(n14743) );
  MUX2_X1 U10950 ( .A(n10040), .B(n10039), .S(n10404), .Z(n9124) );
  NAND2_X1 U10951 ( .A1(n9125), .A2(n9124), .ZN(n9126) );
  NAND2_X1 U10952 ( .A1(n9134), .A2(n9126), .ZN(n11067) );
  OR2_X1 U10953 ( .A1(n11067), .A2(n9209), .ZN(n9132) );
  INV_X1 U10954 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9127) );
  NAND2_X1 U10955 ( .A1(n9105), .A2(n9127), .ZN(n9129) );
  NAND2_X1 U10956 ( .A1(n9129), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9128) );
  MUX2_X1 U10957 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9128), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n9130) );
  AOI22_X1 U10958 ( .A1(n9596), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9349), .B2(
        n10069), .ZN(n9131) );
  MUX2_X1 U10959 ( .A(n14743), .B(n11486), .S(n9538), .Z(n9152) );
  MUX2_X1 U10960 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10404), .Z(n9135) );
  NAND2_X1 U10961 ( .A1(n9135), .A2(SI_10_), .ZN(n9164) );
  OAI21_X1 U10962 ( .B1(n9135), .B2(SI_10_), .A(n9164), .ZN(n9136) );
  INV_X1 U10963 ( .A(n9136), .ZN(n9137) );
  NAND2_X1 U10964 ( .A1(n9166), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9140) );
  XNOR2_X1 U10965 ( .A(n9140), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10095) );
  AOI22_X1 U10966 ( .A1(n9596), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9349), 
        .B2(n10095), .ZN(n9141) );
  INV_X1 U10967 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9143) );
  NOR2_X1 U10968 ( .A1(n9144), .A2(n9143), .ZN(n9179) );
  INV_X1 U10969 ( .A(n9179), .ZN(n9177) );
  NAND2_X1 U10970 ( .A1(n9144), .A2(n9143), .ZN(n9145) );
  NAND2_X1 U10971 ( .A1(n9177), .A2(n9145), .ZN(n11508) );
  OR2_X1 U10972 ( .A1(n9542), .A2(n11508), .ZN(n9150) );
  NAND2_X1 U10973 ( .A1(n9301), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9149) );
  INV_X1 U10974 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11493) );
  OR2_X1 U10975 ( .A1(n9544), .A2(n11493), .ZN(n9148) );
  INV_X1 U10976 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9146) );
  OR2_X1 U10977 ( .A1(n9546), .A2(n9146), .ZN(n9147) );
  NAND4_X1 U10978 ( .A1(n9150), .A2(n9149), .A3(n9148), .A4(n9147), .ZN(n14742) );
  INV_X1 U10979 ( .A(n11486), .ZN(n15877) );
  MUX2_X1 U10980 ( .A(n11485), .B(n15877), .S(n9606), .Z(n9151) );
  AND2_X1 U10981 ( .A1(n14742), .A2(n9606), .ZN(n9154) );
  OAI21_X1 U10982 ( .B1(n9606), .B2(n14742), .A(n11550), .ZN(n9153) );
  OAI21_X1 U10983 ( .B1(n9154), .B2(n11550), .A(n9153), .ZN(n9155) );
  NAND2_X1 U10984 ( .A1(n9301), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9163) );
  XNOR2_X1 U10985 ( .A(n9177), .B(P1_REG3_REG_11__SCAN_IN), .ZN(n11939) );
  NAND2_X1 U10986 ( .A1(n9157), .A2(n11939), .ZN(n9162) );
  INV_X1 U10987 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9158) );
  OR2_X1 U10988 ( .A1(n9544), .A2(n9158), .ZN(n9161) );
  INV_X1 U10989 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9159) );
  OR2_X1 U10990 ( .A1(n9546), .A2(n9159), .ZN(n9160) );
  NAND4_X1 U10991 ( .A1(n9163), .A2(n9162), .A3(n9161), .A4(n9160), .ZN(n14741) );
  MUX2_X1 U10992 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n10404), .Z(n9187) );
  XNOR2_X1 U10993 ( .A(n9187), .B(SI_11_), .ZN(n9190) );
  XNOR2_X1 U10994 ( .A(n9191), .B(n9190), .ZN(n11298) );
  NAND2_X1 U10995 ( .A1(n11298), .A2(n9595), .ZN(n9171) );
  INV_X1 U10996 ( .A(n9166), .ZN(n9168) );
  INV_X1 U10997 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9167) );
  NAND2_X1 U10998 ( .A1(n9168), .A2(n9167), .ZN(n9192) );
  NAND2_X1 U10999 ( .A1(n9192), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9169) );
  XNOR2_X1 U11000 ( .A(n9169), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10241) );
  AOI22_X1 U11001 ( .A1(n9596), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9349), 
        .B2(n10241), .ZN(n9170) );
  MUX2_X1 U11002 ( .A(n14741), .B(n15917), .S(n9538), .Z(n9173) );
  MUX2_X1 U11003 ( .A(n14741), .B(n15917), .S(n9606), .Z(n9172) );
  INV_X1 U11004 ( .A(n9173), .ZN(n9174) );
  INV_X1 U11005 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9176) );
  INV_X1 U11006 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9175) );
  OAI21_X1 U11007 ( .B1(n9177), .B2(n9176), .A(n9175), .ZN(n9180) );
  AND2_X1 U11008 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n9178) );
  INV_X1 U11009 ( .A(n9215), .ZN(n9216) );
  NAND2_X1 U11010 ( .A1(n9180), .A2(n9216), .ZN(n12130) );
  OR2_X1 U11011 ( .A1(n9542), .A2(n12130), .ZN(n9186) );
  NAND2_X1 U11012 ( .A1(n9301), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9185) );
  INV_X1 U11013 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9181) );
  OR2_X1 U11014 ( .A1(n9544), .A2(n9181), .ZN(n9184) );
  INV_X1 U11015 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9182) );
  OR2_X1 U11016 ( .A1(n9546), .A2(n9182), .ZN(n9183) );
  NAND4_X1 U11017 ( .A1(n9186), .A2(n9185), .A3(n9184), .A4(n9183), .ZN(n14740) );
  INV_X1 U11018 ( .A(n9187), .ZN(n9188) );
  NAND2_X1 U11019 ( .A1(n9188), .A2(n9920), .ZN(n9189) );
  MUX2_X1 U11020 ( .A(n10276), .B(n10287), .S(n10404), .Z(n9200) );
  XNOR2_X1 U11021 ( .A(n9200), .B(SI_12_), .ZN(n9198) );
  XNOR2_X1 U11022 ( .A(n9199), .B(n9198), .ZN(n11514) );
  NAND2_X1 U11023 ( .A1(n11514), .A2(n9595), .ZN(n9195) );
  NAND2_X1 U11024 ( .A1(n9193), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9211) );
  XNOR2_X1 U11025 ( .A(n9211), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10636) );
  AOI22_X1 U11026 ( .A1(n9596), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9349), 
        .B2(n10636), .ZN(n9194) );
  MUX2_X1 U11027 ( .A(n14740), .B(n12127), .S(n9606), .Z(n9197) );
  MUX2_X1 U11028 ( .A(n14740), .B(n12127), .S(n9538), .Z(n9196) );
  NAND2_X1 U11029 ( .A1(n9199), .A2(n9198), .ZN(n9202) );
  NAND2_X1 U11030 ( .A1(n9200), .A2(n11850), .ZN(n9201) );
  MUX2_X1 U11031 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n10404), .Z(n9203) );
  NAND2_X1 U11032 ( .A1(n9203), .A2(SI_13_), .ZN(n9237) );
  INV_X1 U11033 ( .A(n9203), .ZN(n9204) );
  NAND2_X1 U11034 ( .A1(n9204), .A2(n11848), .ZN(n9205) );
  NAND2_X1 U11035 ( .A1(n9237), .A2(n9205), .ZN(n9206) );
  NAND2_X1 U11036 ( .A1(n9207), .A2(n9206), .ZN(n9208) );
  NAND2_X1 U11037 ( .A1(n9238), .A2(n9208), .ZN(n11609) );
  OR2_X1 U11038 ( .A1(n11609), .A2(n9209), .ZN(n9214) );
  NAND2_X1 U11039 ( .A1(n9211), .A2(n9210), .ZN(n9212) );
  NAND2_X1 U11040 ( .A1(n9212), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9240) );
  XNOR2_X1 U11041 ( .A(n9240), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U11042 ( .A1(n9596), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9349), 
        .B2(n10862), .ZN(n9213) );
  NAND2_X1 U11043 ( .A1(n9215), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9229) );
  INV_X1 U11044 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n12273) );
  NAND2_X1 U11045 ( .A1(n9216), .A2(n12273), .ZN(n9217) );
  NAND2_X1 U11046 ( .A1(n9229), .A2(n9217), .ZN(n12272) );
  OR2_X1 U11047 ( .A1(n9542), .A2(n12272), .ZN(n9223) );
  NAND2_X1 U11048 ( .A1(n9301), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9222) );
  INV_X1 U11049 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9218) );
  OR2_X1 U11050 ( .A1(n9544), .A2(n9218), .ZN(n9221) );
  INV_X1 U11051 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9219) );
  OR2_X1 U11052 ( .A1(n9546), .A2(n9219), .ZN(n9220) );
  NAND4_X1 U11053 ( .A1(n9223), .A2(n9222), .A3(n9221), .A4(n9220), .ZN(n14739) );
  MUX2_X1 U11054 ( .A(n12269), .B(n14739), .S(n9606), .Z(n9226) );
  MUX2_X1 U11055 ( .A(n12269), .B(n14739), .S(n9538), .Z(n9224) );
  INV_X1 U11056 ( .A(n9226), .ZN(n9227) );
  INV_X1 U11057 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9228) );
  NAND2_X1 U11058 ( .A1(n9229), .A2(n9228), .ZN(n9230) );
  NAND2_X1 U11059 ( .A1(n9250), .A2(n9230), .ZN(n14636) );
  OR2_X1 U11060 ( .A1(n9542), .A2(n14636), .ZN(n9236) );
  NAND2_X1 U11061 ( .A1(n9301), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9235) );
  INV_X1 U11062 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9231) );
  OR2_X1 U11063 ( .A1(n9544), .A2(n9231), .ZN(n9234) );
  INV_X1 U11064 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9232) );
  OR2_X1 U11065 ( .A1(n9546), .A2(n9232), .ZN(n9233) );
  NAND4_X1 U11066 ( .A1(n9236), .A2(n9235), .A3(n9234), .A4(n9233), .ZN(n15978) );
  MUX2_X1 U11067 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n10404), .Z(n9259) );
  XNOR2_X1 U11068 ( .A(n9259), .B(SI_14_), .ZN(n9257) );
  XNOR2_X1 U11069 ( .A(n9258), .B(n9257), .ZN(n11980) );
  NAND2_X1 U11070 ( .A1(n11980), .A2(n9595), .ZN(n9244) );
  INV_X1 U11071 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9239) );
  NAND2_X1 U11072 ( .A1(n9240), .A2(n9239), .ZN(n9241) );
  NAND2_X1 U11073 ( .A1(n9241), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9242) );
  XNOR2_X1 U11074 ( .A(n9242), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U11075 ( .A1(n9596), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n9349), 
        .B2(n11595), .ZN(n9243) );
  MUX2_X1 U11076 ( .A(n15978), .B(n15165), .S(n9606), .Z(n9247) );
  MUX2_X1 U11077 ( .A(n15978), .B(n15165), .S(n9538), .Z(n9245) );
  INV_X1 U11078 ( .A(n9247), .ZN(n9248) );
  INV_X1 U11079 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9249) );
  NAND2_X1 U11080 ( .A1(n9250), .A2(n9249), .ZN(n9251) );
  NAND2_X1 U11081 ( .A1(n9276), .A2(n9251), .ZN(n15984) );
  OR2_X1 U11082 ( .A1(n9542), .A2(n15984), .ZN(n9256) );
  NAND2_X1 U11083 ( .A1(n9301), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9255) );
  INV_X1 U11084 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n12227) );
  OR2_X1 U11085 ( .A1(n9544), .A2(n12227), .ZN(n9254) );
  INV_X1 U11086 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9252) );
  OR2_X1 U11087 ( .A1(n9546), .A2(n9252), .ZN(n9253) );
  NAND4_X1 U11088 ( .A1(n9256), .A2(n9255), .A3(n9254), .A4(n9253), .ZN(n16000) );
  INV_X1 U11089 ( .A(n9259), .ZN(n9260) );
  NAND2_X1 U11090 ( .A1(n9260), .A2(n11818), .ZN(n9261) );
  MUX2_X1 U11091 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n10404), .Z(n9285) );
  XNOR2_X1 U11092 ( .A(n9285), .B(n11711), .ZN(n9283) );
  XNOR2_X1 U11093 ( .A(n9284), .B(n9283), .ZN(n12055) );
  NAND2_X1 U11094 ( .A1(n12055), .A2(n9595), .ZN(n9266) );
  NAND2_X1 U11095 ( .A1(n9262), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9263) );
  XNOR2_X1 U11096 ( .A(n9263), .B(n8913), .ZN(n15433) );
  INV_X1 U11097 ( .A(n15433), .ZN(n9264) );
  AOI22_X1 U11098 ( .A1(n9596), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9349), 
        .B2(n9264), .ZN(n9265) );
  MUX2_X1 U11099 ( .A(n16000), .B(n15989), .S(n9538), .Z(n9270) );
  MUX2_X1 U11100 ( .A(n16000), .B(n15989), .S(n9606), .Z(n9268) );
  NAND2_X1 U11101 ( .A1(n9269), .A2(n9268), .ZN(n9273) );
  INV_X1 U11102 ( .A(n9270), .ZN(n9271) );
  NAND2_X1 U11103 ( .A1(n7295), .A2(n9271), .ZN(n9272) );
  INV_X1 U11104 ( .A(n9276), .ZN(n9274) );
  NAND2_X1 U11105 ( .A1(n9274), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9298) );
  INV_X1 U11106 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9275) );
  NAND2_X1 U11107 ( .A1(n9276), .A2(n9275), .ZN(n9277) );
  NAND2_X1 U11108 ( .A1(n9298), .A2(n9277), .ZN(n16008) );
  OR2_X1 U11109 ( .A1(n9542), .A2(n16008), .ZN(n9282) );
  NAND2_X1 U11110 ( .A1(n9301), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9281) );
  INV_X1 U11111 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n15056) );
  OR2_X1 U11112 ( .A1(n9544), .A2(n15056), .ZN(n9280) );
  INV_X1 U11113 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9278) );
  OR2_X1 U11114 ( .A1(n9546), .A2(n9278), .ZN(n9279) );
  NAND4_X1 U11115 ( .A1(n9282), .A2(n9281), .A3(n9280), .A4(n9279), .ZN(n16028) );
  INV_X1 U11116 ( .A(n9285), .ZN(n9286) );
  NAND2_X1 U11117 ( .A1(n9286), .A2(n11711), .ZN(n9287) );
  MUX2_X1 U11118 ( .A(n10895), .B(n9289), .S(n10404), .Z(n9309) );
  XNOR2_X1 U11119 ( .A(n9309), .B(SI_16_), .ZN(n9307) );
  XNOR2_X1 U11120 ( .A(n9308), .B(n9307), .ZN(n12170) );
  NAND2_X1 U11121 ( .A1(n12170), .A2(n9595), .ZN(n9293) );
  NAND2_X1 U11122 ( .A1(n9290), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9291) );
  XNOR2_X1 U11123 ( .A(n9291), .B(P1_IR_REG_16__SCAN_IN), .ZN(n12112) );
  AOI22_X1 U11124 ( .A1(n9596), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9349), 
        .B2(n12112), .ZN(n9292) );
  MUX2_X1 U11125 ( .A(n16028), .B(n16013), .S(n9606), .Z(n9295) );
  MUX2_X1 U11126 ( .A(n16028), .B(n16013), .S(n9538), .Z(n9294) );
  INV_X1 U11127 ( .A(n9295), .ZN(n9296) );
  INV_X1 U11128 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9297) );
  NAND2_X1 U11129 ( .A1(n9298), .A2(n9297), .ZN(n9299) );
  NAND2_X1 U11130 ( .A1(n9355), .A2(n9299), .ZN(n16040) );
  INV_X1 U11131 ( .A(n16040), .ZN(n9300) );
  NAND2_X1 U11132 ( .A1(n9300), .A2(n9157), .ZN(n9306) );
  NAND2_X1 U11133 ( .A1(n9301), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9305) );
  INV_X1 U11134 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15032) );
  OR2_X1 U11135 ( .A1(n9544), .A2(n15032), .ZN(n9304) );
  INV_X1 U11136 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9302) );
  OR2_X1 U11137 ( .A1(n9546), .A2(n9302), .ZN(n9303) );
  NAND4_X1 U11138 ( .A1(n9306), .A2(n9305), .A3(n9304), .A4(n9303), .ZN(n16001) );
  NAND2_X1 U11139 ( .A1(n9309), .A2(n11845), .ZN(n9310) );
  MUX2_X1 U11140 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n10404), .Z(n9326) );
  XNOR2_X1 U11141 ( .A(n9326), .B(n11840), .ZN(n9324) );
  XNOR2_X1 U11142 ( .A(n9325), .B(n9324), .ZN(n12320) );
  NAND2_X1 U11143 ( .A1(n12320), .A2(n9595), .ZN(n9315) );
  NAND2_X1 U11144 ( .A1(n9312), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9313) );
  XNOR2_X1 U11145 ( .A(n9313), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14797) );
  AOI22_X1 U11146 ( .A1(n9596), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9349), 
        .B2(n14797), .ZN(n9314) );
  MUX2_X1 U11147 ( .A(n16001), .B(n16027), .S(n9538), .Z(n9319) );
  NAND2_X1 U11148 ( .A1(n9318), .A2(n9319), .ZN(n9317) );
  MUX2_X1 U11149 ( .A(n16001), .B(n16027), .S(n9606), .Z(n9316) );
  NAND2_X1 U11150 ( .A1(n9317), .A2(n9316), .ZN(n9323) );
  INV_X1 U11151 ( .A(n9318), .ZN(n9321) );
  INV_X1 U11152 ( .A(n9319), .ZN(n9320) );
  NAND2_X1 U11153 ( .A1(n9321), .A2(n9320), .ZN(n9322) );
  INV_X1 U11154 ( .A(n9326), .ZN(n9327) );
  NAND2_X1 U11155 ( .A1(n9327), .A2(n11840), .ZN(n9328) );
  MUX2_X1 U11156 ( .A(n11281), .B(n11284), .S(n10404), .Z(n9330) );
  NAND2_X1 U11157 ( .A1(n9331), .A2(n9330), .ZN(n9332) );
  NAND2_X1 U11158 ( .A1(n9333), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9334) );
  XNOR2_X1 U11159 ( .A(n9334), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14814) );
  AOI22_X1 U11160 ( .A1(n9596), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9349), 
        .B2(n14814), .ZN(n9335) );
  INV_X1 U11161 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14799) );
  INV_X1 U11162 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9337) );
  OR2_X1 U11163 ( .A1(n9544), .A2(n9337), .ZN(n9340) );
  INV_X1 U11164 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9338) );
  OR2_X1 U11165 ( .A1(n9546), .A2(n9338), .ZN(n9339) );
  AND2_X1 U11166 ( .A1(n9340), .A2(n9339), .ZN(n9342) );
  XNOR2_X1 U11167 ( .A(n9355), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n15019) );
  NAND2_X1 U11168 ( .A1(n15019), .A2(n9157), .ZN(n9341) );
  OAI211_X1 U11169 ( .C1(n9582), .C2(n14799), .A(n9342), .B(n9341), .ZN(n16030) );
  MUX2_X1 U11170 ( .A(n15153), .B(n16030), .S(n9538), .Z(n9344) );
  MUX2_X1 U11171 ( .A(n15153), .B(n16030), .S(n9606), .Z(n9343) );
  INV_X1 U11172 ( .A(n9344), .ZN(n9345) );
  MUX2_X1 U11173 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10404), .Z(n9374) );
  XNOR2_X1 U11174 ( .A(n9374), .B(SI_19_), .ZN(n9375) );
  XNOR2_X1 U11175 ( .A(n9376), .B(n9375), .ZN(n12334) );
  NAND2_X1 U11176 ( .A1(n12334), .A2(n9595), .ZN(n9351) );
  AOI22_X1 U11177 ( .A1(n9596), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9349), 
        .B2(n9348), .ZN(n9350) );
  NAND2_X1 U11178 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n9352) );
  INV_X1 U11179 ( .A(n9370), .ZN(n9357) );
  INV_X1 U11180 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9354) );
  INV_X1 U11181 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9353) );
  OAI21_X1 U11182 ( .B1(n9355), .B2(n9354), .A(n9353), .ZN(n9356) );
  NAND2_X1 U11183 ( .A1(n9357), .A2(n9356), .ZN(n14989) );
  NAND2_X1 U11184 ( .A1(n9301), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n9359) );
  INV_X1 U11185 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14817) );
  OR2_X1 U11186 ( .A1(n9544), .A2(n14817), .ZN(n9358) );
  AND2_X1 U11187 ( .A1(n9359), .A2(n9358), .ZN(n9361) );
  NAND2_X1 U11188 ( .A1(n8952), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9360) );
  OAI211_X1 U11189 ( .C1(n14989), .C2(n9542), .A(n9361), .B(n9360), .ZN(n15008) );
  MUX2_X1 U11190 ( .A(n15145), .B(n15008), .S(n9606), .Z(n9365) );
  NAND2_X1 U11191 ( .A1(n9364), .A2(n9365), .ZN(n9363) );
  MUX2_X1 U11192 ( .A(n15008), .B(n15145), .S(n9606), .Z(n9362) );
  NAND2_X1 U11193 ( .A1(n9363), .A2(n9362), .ZN(n9369) );
  INV_X1 U11194 ( .A(n9364), .ZN(n9367) );
  INV_X1 U11195 ( .A(n9365), .ZN(n9366) );
  NAND2_X1 U11196 ( .A1(n9367), .A2(n9366), .ZN(n9368) );
  NOR2_X1 U11197 ( .A1(n9370), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9371) );
  OR2_X1 U11198 ( .A1(n9382), .A2(n9371), .ZN(n14977) );
  INV_X1 U11199 ( .A(n9544), .ZN(n9578) );
  AOI22_X1 U11200 ( .A1(n9301), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n9578), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9373) );
  NAND2_X1 U11201 ( .A1(n8952), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9372) );
  OAI211_X1 U11202 ( .C1(n14977), .C2(n9542), .A(n9373), .B(n9372), .ZN(n14963) );
  MUX2_X1 U11203 ( .A(n11666), .B(n12349), .S(n10404), .Z(n9386) );
  XNOR2_X1 U11204 ( .A(n9386), .B(SI_20_), .ZN(n9377) );
  XNOR2_X1 U11205 ( .A(n9390), .B(n9377), .ZN(n12348) );
  NAND2_X1 U11206 ( .A1(n12348), .A2(n9595), .ZN(n9379) );
  NAND2_X1 U11207 ( .A1(n9596), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9378) );
  MUX2_X1 U11208 ( .A(n14963), .B(n14562), .S(n9606), .Z(n9381) );
  MUX2_X1 U11209 ( .A(n14963), .B(n14562), .S(n9538), .Z(n9380) );
  OR2_X1 U11210 ( .A1(n9382), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9383) );
  NAND2_X1 U11211 ( .A1(n9382), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9401) );
  NAND2_X1 U11212 ( .A1(n9383), .A2(n9401), .ZN(n14964) );
  AOI22_X1 U11213 ( .A1(n9578), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n8952), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n9385) );
  NAND2_X1 U11214 ( .A1(n9301), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9384) );
  OAI211_X1 U11215 ( .C1(n14964), .C2(n9542), .A(n9385), .B(n9384), .ZN(n14976) );
  NOR2_X1 U11216 ( .A1(n9387), .A2(SI_20_), .ZN(n9389) );
  NAND2_X1 U11217 ( .A1(n9387), .A2(SI_20_), .ZN(n9388) );
  MUX2_X1 U11218 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10404), .Z(n9397) );
  XNOR2_X1 U11219 ( .A(n9397), .B(SI_21_), .ZN(n9394) );
  XNOR2_X1 U11220 ( .A(n9396), .B(n9394), .ZN(n12361) );
  NAND2_X1 U11221 ( .A1(n9596), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9391) );
  MUX2_X1 U11222 ( .A(n14976), .B(n14961), .S(n9538), .Z(n9409) );
  NAND2_X1 U11223 ( .A1(n9410), .A2(n9409), .ZN(n9393) );
  MUX2_X1 U11224 ( .A(n14976), .B(n14961), .S(n9606), .Z(n9392) );
  NAND2_X1 U11225 ( .A1(n9393), .A2(n9392), .ZN(n9408) );
  INV_X1 U11226 ( .A(n9394), .ZN(n9395) );
  NAND2_X1 U11227 ( .A1(n9397), .A2(SI_21_), .ZN(n9398) );
  NAND2_X1 U11228 ( .A1(n12374), .A2(n10395), .ZN(n9399) );
  NAND2_X1 U11229 ( .A1(n9301), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n9407) );
  INV_X1 U11230 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9400) );
  OR2_X1 U11231 ( .A1(n9544), .A2(n9400), .ZN(n9406) );
  NAND2_X1 U11232 ( .A1(n9402), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9416) );
  OAI21_X1 U11233 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n9402), .A(n9416), .ZN(
        n14710) );
  OR2_X1 U11234 ( .A1(n9542), .A2(n14710), .ZN(n9405) );
  INV_X1 U11235 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9403) );
  OR2_X1 U11236 ( .A1(n9546), .A2(n9403), .ZN(n9404) );
  XNOR2_X1 U11237 ( .A(n14954), .B(n14927), .ZN(n14942) );
  OAI211_X1 U11238 ( .C1(n9410), .C2(n9409), .A(n9408), .B(n14942), .ZN(n9415)
         );
  NOR2_X1 U11239 ( .A1(n14962), .A2(n9606), .ZN(n9413) );
  NAND2_X1 U11240 ( .A1(n14962), .A2(n9606), .ZN(n9411) );
  NAND2_X1 U11241 ( .A1(n14954), .A2(n9411), .ZN(n9412) );
  OAI21_X1 U11242 ( .B1(n14954), .B2(n9413), .A(n9412), .ZN(n9414) );
  NAND2_X1 U11243 ( .A1(n9415), .A2(n9414), .ZN(n9429) );
  NAND2_X1 U11244 ( .A1(n9417), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9432) );
  OAI21_X1 U11245 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n9417), .A(n9432), .ZN(
        n14928) );
  OR2_X1 U11246 ( .A1(n9542), .A2(n14928), .ZN(n9422) );
  NAND2_X1 U11247 ( .A1(n9301), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9421) );
  INV_X1 U11248 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14931) );
  OR2_X1 U11249 ( .A1(n9544), .A2(n14931), .ZN(n9420) );
  INV_X1 U11250 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9418) );
  OR2_X1 U11251 ( .A1(n9546), .A2(n9418), .ZN(n9419) );
  NAND4_X1 U11252 ( .A1(n9422), .A2(n9421), .A3(n9420), .A4(n9419), .ZN(n14738) );
  MUX2_X1 U11253 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10404), .Z(n9445) );
  NAND2_X1 U11254 ( .A1(n12374), .A2(n9445), .ZN(n12378) );
  NAND2_X1 U11255 ( .A1(n9442), .A2(SI_22_), .ZN(n9423) );
  NAND2_X1 U11256 ( .A1(n12378), .A2(n9423), .ZN(n9425) );
  MUX2_X1 U11257 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10404), .Z(n9446) );
  XNOR2_X1 U11258 ( .A(n9446), .B(SI_23_), .ZN(n9424) );
  NAND2_X1 U11259 ( .A1(n15211), .A2(n9595), .ZN(n9427) );
  NAND2_X1 U11260 ( .A1(n9596), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9426) );
  MUX2_X1 U11261 ( .A(n14738), .B(n15117), .S(n9538), .Z(n9430) );
  MUX2_X1 U11262 ( .A(n14738), .B(n15117), .S(n9606), .Z(n9428) );
  INV_X1 U11263 ( .A(n9430), .ZN(n9431) );
  NAND2_X1 U11264 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n9433), .ZN(n9461) );
  OAI21_X1 U11265 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n9433), .A(n9461), .ZN(
        n14908) );
  OR2_X1 U11266 ( .A1(n9542), .A2(n14908), .ZN(n9439) );
  NAND2_X1 U11267 ( .A1(n9301), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9438) );
  INV_X1 U11268 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9434) );
  OR2_X1 U11269 ( .A1(n9544), .A2(n9434), .ZN(n9437) );
  INV_X1 U11270 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9435) );
  OR2_X1 U11271 ( .A1(n9546), .A2(n9435), .ZN(n9436) );
  NAND4_X1 U11272 ( .A1(n9439), .A2(n9438), .A3(n9437), .A4(n9436), .ZN(n14925) );
  INV_X1 U11273 ( .A(n9446), .ZN(n9440) );
  AOI22_X1 U11274 ( .A1(n9443), .A2(n12375), .B1(n9440), .B2(n11723), .ZN(
        n9441) );
  NAND2_X1 U11275 ( .A1(n9442), .A2(n9441), .ZN(n9449) );
  OAI21_X1 U11276 ( .B1(n12375), .B2(n9443), .A(n11723), .ZN(n9447) );
  AND2_X1 U11277 ( .A1(SI_22_), .A2(SI_23_), .ZN(n9444) );
  AOI22_X1 U11278 ( .A1(n9447), .A2(n9446), .B1(n9445), .B2(n9444), .ZN(n9448)
         );
  XNOR2_X1 U11279 ( .A(n9491), .B(SI_24_), .ZN(n9470) );
  MUX2_X1 U11280 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10404), .Z(n9492) );
  XNOR2_X1 U11281 ( .A(n9470), .B(n9492), .ZN(n14497) );
  NAND2_X1 U11282 ( .A1(n14497), .A2(n9595), .ZN(n9451) );
  NAND2_X1 U11283 ( .A1(n9596), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9450) );
  MUX2_X1 U11284 ( .A(n14925), .B(n15107), .S(n9606), .Z(n9455) );
  MUX2_X1 U11285 ( .A(n14925), .B(n15107), .S(n9538), .Z(n9452) );
  NAND2_X1 U11286 ( .A1(n9453), .A2(n9452), .ZN(n9458) );
  INV_X1 U11287 ( .A(n9454), .ZN(n9456) );
  NAND2_X1 U11288 ( .A1(n9456), .A2(n8235), .ZN(n9457) );
  INV_X1 U11289 ( .A(n9461), .ZN(n9459) );
  NAND2_X1 U11290 ( .A1(n9459), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9481) );
  INV_X1 U11291 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9460) );
  NAND2_X1 U11292 ( .A1(n9461), .A2(n9460), .ZN(n9462) );
  NAND2_X1 U11293 ( .A1(n9481), .A2(n9462), .ZN(n14897) );
  OR2_X1 U11294 ( .A1(n9542), .A2(n14897), .ZN(n9468) );
  NAND2_X1 U11295 ( .A1(n9301), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9467) );
  INV_X1 U11296 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9463) );
  OR2_X1 U11297 ( .A1(n9544), .A2(n9463), .ZN(n9466) );
  INV_X1 U11298 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9464) );
  OR2_X1 U11299 ( .A1(n9546), .A2(n9464), .ZN(n9465) );
  NAND4_X1 U11300 ( .A1(n9468), .A2(n9467), .A3(n9466), .A4(n9465), .ZN(n14876) );
  INV_X1 U11301 ( .A(n9492), .ZN(n9489) );
  INV_X1 U11302 ( .A(n9491), .ZN(n9469) );
  OAI22_X1 U11303 ( .A1(n9470), .A2(n9489), .B1(n9469), .B2(n11828), .ZN(n9474) );
  MUX2_X1 U11304 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n10404), .Z(n9471) );
  NAND2_X1 U11305 ( .A1(n9471), .A2(SI_25_), .ZN(n9495) );
  INV_X1 U11306 ( .A(n9471), .ZN(n9472) );
  NAND2_X1 U11307 ( .A1(n9472), .A2(n11713), .ZN(n9493) );
  NAND2_X1 U11308 ( .A1(n9495), .A2(n9493), .ZN(n9473) );
  XNOR2_X1 U11309 ( .A(n9474), .B(n9473), .ZN(n14494) );
  NAND2_X1 U11310 ( .A1(n14494), .A2(n9595), .ZN(n9476) );
  NAND2_X1 U11311 ( .A1(n9596), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9475) );
  MUX2_X1 U11312 ( .A(n14876), .B(n14895), .S(n9538), .Z(n9478) );
  MUX2_X1 U11313 ( .A(n14876), .B(n14895), .S(n9606), .Z(n9477) );
  INV_X1 U11314 ( .A(n9481), .ZN(n9479) );
  NAND2_X1 U11315 ( .A1(n9479), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9504) );
  INV_X1 U11316 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9480) );
  NAND2_X1 U11317 ( .A1(n9481), .A2(n9480), .ZN(n9482) );
  NAND2_X1 U11318 ( .A1(n9504), .A2(n9482), .ZN(n14881) );
  OR2_X1 U11319 ( .A1(n9542), .A2(n14881), .ZN(n9488) );
  NAND2_X1 U11320 ( .A1(n9301), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9487) );
  INV_X1 U11321 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9483) );
  OR2_X1 U11322 ( .A1(n9544), .A2(n9483), .ZN(n9486) );
  INV_X1 U11323 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9484) );
  OR2_X1 U11324 ( .A1(n9546), .A2(n9484), .ZN(n9485) );
  NAND4_X1 U11325 ( .A1(n9488), .A2(n9487), .A3(n9486), .A4(n9485), .ZN(n14896) );
  OAI21_X1 U11326 ( .B1(n11828), .B2(n9489), .A(n9495), .ZN(n9490) );
  NOR2_X1 U11327 ( .A1(n9492), .A2(SI_24_), .ZN(n9496) );
  INV_X1 U11328 ( .A(n9493), .ZN(n9494) );
  AOI21_X1 U11329 ( .B1(n9496), .B2(n9495), .A(n9494), .ZN(n9497) );
  MUX2_X1 U11330 ( .A(n15201), .B(n14492), .S(n10404), .Z(n9512) );
  XNOR2_X1 U11331 ( .A(n9512), .B(SI_26_), .ZN(n9511) );
  XNOR2_X1 U11332 ( .A(n9514), .B(n9511), .ZN(n14491) );
  NAND2_X1 U11333 ( .A1(n14491), .A2(n9595), .ZN(n9499) );
  NAND2_X1 U11334 ( .A1(n9571), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9498) );
  MUX2_X1 U11335 ( .A(n14896), .B(n15092), .S(n9606), .Z(n9501) );
  MUX2_X1 U11336 ( .A(n15092), .B(n14896), .S(n9606), .Z(n9500) );
  INV_X1 U11337 ( .A(n9504), .ZN(n9502) );
  NAND2_X1 U11338 ( .A1(n9502), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9522) );
  INV_X1 U11339 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9503) );
  NAND2_X1 U11340 ( .A1(n9504), .A2(n9503), .ZN(n9505) );
  NAND2_X1 U11341 ( .A1(n9522), .A2(n9505), .ZN(n14862) );
  OR2_X1 U11342 ( .A1(n9542), .A2(n14862), .ZN(n9510) );
  NAND2_X1 U11343 ( .A1(n9301), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9509) );
  INV_X1 U11344 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14863) );
  OR2_X1 U11345 ( .A1(n9544), .A2(n14863), .ZN(n9508) );
  INV_X1 U11346 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9506) );
  OR2_X1 U11347 ( .A1(n9546), .A2(n9506), .ZN(n9507) );
  NAND4_X1 U11348 ( .A1(n9510), .A2(n9509), .A3(n9508), .A4(n9507), .ZN(n14877) );
  INV_X1 U11349 ( .A(n9511), .ZN(n9513) );
  MUX2_X1 U11350 ( .A(n12499), .B(n14489), .S(n10404), .Z(n9551) );
  NAND2_X1 U11351 ( .A1(n12498), .A2(n9595), .ZN(n9516) );
  NAND2_X1 U11352 ( .A1(n9596), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9515) );
  MUX2_X1 U11353 ( .A(n14877), .B(n15087), .S(n9538), .Z(n9518) );
  MUX2_X1 U11354 ( .A(n14877), .B(n15087), .S(n9606), .Z(n9517) );
  INV_X1 U11355 ( .A(n9518), .ZN(n9519) );
  INV_X1 U11356 ( .A(n9522), .ZN(n9520) );
  NAND2_X1 U11357 ( .A1(n9520), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n12533) );
  INV_X1 U11358 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9521) );
  NAND2_X1 U11359 ( .A1(n9522), .A2(n9521), .ZN(n9523) );
  NAND2_X1 U11360 ( .A1(n12533), .A2(n9523), .ZN(n14851) );
  OR2_X1 U11361 ( .A1(n9542), .A2(n14851), .ZN(n9528) );
  NAND2_X1 U11362 ( .A1(n9301), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9527) );
  INV_X1 U11363 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n14852) );
  OR2_X1 U11364 ( .A1(n9544), .A2(n14852), .ZN(n9526) );
  INV_X1 U11365 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9524) );
  OR2_X1 U11366 ( .A1(n9546), .A2(n9524), .ZN(n9525) );
  NAND4_X1 U11367 ( .A1(n9528), .A2(n9527), .A3(n9526), .A4(n9525), .ZN(n14737) );
  NAND2_X1 U11368 ( .A1(n9529), .A2(SI_27_), .ZN(n9531) );
  INV_X1 U11369 ( .A(n9551), .ZN(n9554) );
  NAND2_X1 U11370 ( .A1(n9553), .A2(n9554), .ZN(n9530) );
  NAND2_X1 U11371 ( .A1(n9531), .A2(n9530), .ZN(n9535) );
  MUX2_X1 U11372 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n10404), .Z(n9532) );
  NAND2_X1 U11373 ( .A1(n9532), .A2(SI_28_), .ZN(n9556) );
  NOR2_X1 U11374 ( .A1(n9532), .A2(SI_28_), .ZN(n9555) );
  INV_X1 U11375 ( .A(n9555), .ZN(n9533) );
  NAND2_X1 U11376 ( .A1(n9556), .A2(n9533), .ZN(n9534) );
  NAND2_X1 U11377 ( .A1(n14483), .A2(n9595), .ZN(n9537) );
  NAND2_X1 U11378 ( .A1(n9571), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9536) );
  MUX2_X1 U11379 ( .A(n14737), .B(n15081), .S(n9606), .Z(n9541) );
  MUX2_X1 U11380 ( .A(n14737), .B(n15081), .S(n9538), .Z(n9539) );
  OR2_X1 U11381 ( .A1(n9542), .A2(n12533), .ZN(n9550) );
  NAND2_X1 U11382 ( .A1(n9301), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9549) );
  INV_X1 U11383 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9543) );
  OR2_X1 U11384 ( .A1(n9544), .A2(n9543), .ZN(n9548) );
  INV_X1 U11385 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9545) );
  OR2_X1 U11386 ( .A1(n9546), .A2(n9545), .ZN(n9547) );
  NAND4_X1 U11387 ( .A1(n9550), .A2(n9549), .A3(n9548), .A4(n9547), .ZN(n14736) );
  OAI21_X1 U11388 ( .B1(n9551), .B2(n12031), .A(n9556), .ZN(n9552) );
  OR2_X1 U11389 ( .A1(n9553), .A2(n9552), .ZN(n9559) );
  NOR2_X1 U11390 ( .A1(n9554), .A2(SI_27_), .ZN(n9557) );
  AOI21_X1 U11391 ( .B1(n9557), .B2(n9556), .A(n9555), .ZN(n9558) );
  MUX2_X1 U11392 ( .A(n15198), .B(n14481), .S(n10404), .Z(n9564) );
  XNOR2_X1 U11393 ( .A(n9564), .B(SI_29_), .ZN(n9562) );
  XNOR2_X1 U11394 ( .A(n9563), .B(n9562), .ZN(n14480) );
  NAND2_X1 U11395 ( .A1(n14480), .A2(n9595), .ZN(n9561) );
  NAND2_X1 U11396 ( .A1(n9596), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9560) );
  MUX2_X1 U11397 ( .A(n14736), .B(n12529), .S(n9267), .Z(n9608) );
  NAND2_X1 U11398 ( .A1(n9563), .A2(n9562), .ZN(n9566) );
  NAND2_X1 U11399 ( .A1(n9564), .A2(n13811), .ZN(n9565) );
  NAND2_X1 U11400 ( .A1(n9566), .A2(n9565), .ZN(n9569) );
  MUX2_X1 U11401 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10404), .Z(n9567) );
  NAND2_X1 U11402 ( .A1(n9567), .A2(SI_30_), .ZN(n9590) );
  OAI21_X1 U11403 ( .B1(SI_30_), .B2(n9567), .A(n9590), .ZN(n9568) );
  NAND2_X1 U11404 ( .A1(n9569), .A2(n9568), .ZN(n9570) );
  NAND2_X1 U11405 ( .A1(n13059), .A2(n9595), .ZN(n9573) );
  NAND2_X1 U11406 ( .A1(n9571), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9572) );
  INV_X1 U11407 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9576) );
  NAND2_X1 U11408 ( .A1(n9578), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9575) );
  NAND2_X1 U11409 ( .A1(n8952), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9574) );
  OAI211_X1 U11410 ( .C1(n9582), .C2(n9576), .A(n9575), .B(n9574), .ZN(n14830)
         );
  INV_X1 U11411 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9581) );
  NAND2_X1 U11412 ( .A1(n9578), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9580) );
  NAND2_X1 U11413 ( .A1(n8952), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9579) );
  OAI211_X1 U11414 ( .C1(n9582), .C2(n9581), .A(n9580), .B(n9579), .ZN(n14735)
         );
  OAI21_X1 U11415 ( .B1(n14830), .B2(n8927), .A(n14735), .ZN(n9583) );
  INV_X1 U11416 ( .A(n9583), .ZN(n9584) );
  MUX2_X1 U11417 ( .A(n14835), .B(n9584), .S(n9606), .Z(n9603) );
  INV_X1 U11418 ( .A(n9603), .ZN(n9587) );
  OAI21_X1 U11419 ( .B1(n14830), .B2(n11665), .A(n14735), .ZN(n9585) );
  INV_X1 U11420 ( .A(n9585), .ZN(n9586) );
  MUX2_X1 U11421 ( .A(n14835), .B(n9586), .S(n9538), .Z(n9602) );
  NAND2_X1 U11422 ( .A1(n9587), .A2(n9602), .ZN(n9616) );
  NAND2_X1 U11423 ( .A1(n15217), .A2(n9825), .ZN(n9775) );
  NAND2_X1 U11424 ( .A1(n9706), .A2(n11665), .ZN(n9588) );
  NAND2_X1 U11425 ( .A1(n9775), .A2(n9588), .ZN(n9589) );
  NAND2_X1 U11426 ( .A1(n7541), .A2(n9348), .ZN(n9836) );
  AND2_X1 U11427 ( .A1(n9589), .A2(n9836), .ZN(n9615) );
  NAND2_X1 U11428 ( .A1(n9591), .A2(n9590), .ZN(n9594) );
  MUX2_X1 U11429 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10404), .Z(n9592) );
  XNOR2_X1 U11430 ( .A(n9592), .B(SI_31_), .ZN(n9593) );
  NAND2_X1 U11431 ( .A1(n15194), .A2(n9595), .ZN(n9598) );
  NAND2_X1 U11432 ( .A1(n9596), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n9597) );
  XNOR2_X1 U11433 ( .A(n14828), .B(n14830), .ZN(n9636) );
  NAND3_X1 U11434 ( .A1(n9616), .A2(n9615), .A3(n9636), .ZN(n9644) );
  NOR2_X1 U11435 ( .A1(n9613), .A2(n9644), .ZN(n9611) );
  NAND2_X1 U11436 ( .A1(n15067), .A2(n14830), .ZN(n9601) );
  INV_X1 U11437 ( .A(n14830), .ZN(n9599) );
  NAND2_X1 U11438 ( .A1(n14828), .A2(n9599), .ZN(n9600) );
  MUX2_X1 U11439 ( .A(n9601), .B(n9600), .S(n9606), .Z(n9618) );
  INV_X1 U11440 ( .A(n9602), .ZN(n9604) );
  NAND2_X1 U11441 ( .A1(n9604), .A2(n9603), .ZN(n9645) );
  NAND2_X1 U11442 ( .A1(n12052), .A2(n9824), .ZN(n9639) );
  INV_X1 U11443 ( .A(n9615), .ZN(n9617) );
  AND3_X1 U11444 ( .A1(n9645), .A2(n9639), .A3(n9617), .ZN(n9605) );
  AND2_X1 U11445 ( .A1(n9618), .A2(n9605), .ZN(n9612) );
  INV_X1 U11446 ( .A(n14736), .ZN(n14840) );
  MUX2_X1 U11447 ( .A(n14840), .B(n15075), .S(n9606), .Z(n9607) );
  INV_X1 U11448 ( .A(n9618), .ZN(n9614) );
  AOI211_X1 U11449 ( .C1(n9616), .C2(n9636), .A(n9615), .B(n9614), .ZN(n9642)
         );
  OAI21_X1 U11450 ( .B1(n9618), .B2(n9617), .A(n9639), .ZN(n9641) );
  XOR2_X1 U11451 ( .A(n14736), .B(n12529), .Z(n12527) );
  XNOR2_X1 U11452 ( .A(n14835), .B(n14735), .ZN(n9619) );
  XNOR2_X1 U11453 ( .A(n15107), .B(n14925), .ZN(n14913) );
  NAND2_X1 U11454 ( .A1(n9619), .A2(n14913), .ZN(n9634) );
  INV_X1 U11455 ( .A(n14738), .ZN(n12511) );
  XNOR2_X1 U11456 ( .A(n15117), .B(n12511), .ZN(n14923) );
  NAND2_X1 U11457 ( .A1(n14895), .A2(n14876), .ZN(n12524) );
  OR2_X1 U11458 ( .A1(n14895), .A2(n14876), .ZN(n9620) );
  NAND2_X1 U11459 ( .A1(n12524), .A2(n9620), .ZN(n14892) );
  INV_X1 U11460 ( .A(n14976), .ZN(n14573) );
  INV_X1 U11461 ( .A(n14963), .ZN(n12520) );
  XNOR2_X1 U11462 ( .A(n14562), .B(n12520), .ZN(n14984) );
  INV_X1 U11463 ( .A(n15008), .ZN(n14719) );
  XNOR2_X1 U11464 ( .A(n15153), .B(n16030), .ZN(n15006) );
  XNOR2_X1 U11465 ( .A(n15989), .B(n15050), .ZN(n12237) );
  XNOR2_X1 U11466 ( .A(n15165), .B(n14520), .ZN(n12284) );
  XNOR2_X1 U11467 ( .A(n12127), .B(n12124), .ZN(n11654) );
  XNOR2_X1 U11468 ( .A(n12269), .B(n14739), .ZN(n12230) );
  XNOR2_X1 U11469 ( .A(n11486), .B(n11485), .ZN(n11380) );
  INV_X1 U11470 ( .A(n14744), .ZN(n11376) );
  XNOR2_X1 U11471 ( .A(n11377), .B(n11376), .ZN(n9808) );
  INV_X1 U11472 ( .A(n14745), .ZN(n10997) );
  XNOR2_X1 U11473 ( .A(n15836), .B(n10997), .ZN(n11159) );
  INV_X1 U11474 ( .A(n9621), .ZN(n10687) );
  NAND2_X2 U11475 ( .A1(n9622), .A2(n10503), .ZN(n9812) );
  NAND2_X1 U11476 ( .A1(n9814), .A2(n9623), .ZN(n10504) );
  NOR4_X1 U11477 ( .A1(n10687), .A2(n9812), .A3(n10504), .A4(n15683), .ZN(
        n9626) );
  XNOR2_X1 U11478 ( .A(n10995), .B(n14746), .ZN(n10970) );
  NAND4_X1 U11479 ( .A1(n9626), .A2(n10970), .A3(n9818), .A4(n10646), .ZN(
        n9627) );
  NOR4_X1 U11480 ( .A1(n11380), .A2(n9808), .A3(n11159), .A4(n9627), .ZN(n9628) );
  XNOR2_X1 U11481 ( .A(n15917), .B(n14741), .ZN(n11649) );
  NAND4_X1 U11482 ( .A1(n12230), .A2(n9628), .A3(n11649), .A4(n11542), .ZN(
        n9629) );
  NOR4_X1 U11483 ( .A1(n12237), .A2(n12284), .A3(n11654), .A4(n9629), .ZN(
        n9630) );
  XNOR2_X1 U11484 ( .A(n16027), .B(n16001), .ZN(n15031) );
  XNOR2_X1 U11485 ( .A(n16013), .B(n16028), .ZN(n12503) );
  NAND4_X1 U11486 ( .A1(n15006), .A2(n9630), .A3(n15031), .A4(n12503), .ZN(
        n9631) );
  NOR4_X1 U11487 ( .A1(n14957), .A2(n14984), .A3(n14997), .A4(n9631), .ZN(
        n9632) );
  XNOR2_X1 U11488 ( .A(n15092), .B(n14896), .ZN(n14874) );
  NAND4_X1 U11489 ( .A1(n14892), .A2(n14942), .A3(n9632), .A4(n14874), .ZN(
        n9633) );
  NOR4_X1 U11490 ( .A1(n12527), .A2(n9634), .A3(n14923), .A4(n9633), .ZN(n9637) );
  OR2_X1 U11491 ( .A1(n15081), .A2(n14737), .ZN(n9635) );
  NAND2_X1 U11492 ( .A1(n12526), .A2(n9635), .ZN(n12525) );
  XNOR2_X1 U11493 ( .A(n15087), .B(n14877), .ZN(n14857) );
  NAND4_X1 U11494 ( .A1(n9637), .A2(n12525), .A3(n14857), .A4(n9636), .ZN(
        n9638) );
  XNOR2_X1 U11495 ( .A(n9638), .B(n9348), .ZN(n9640) );
  OAI22_X1 U11496 ( .A1(n9642), .A2(n9641), .B1(n9640), .B2(n9639), .ZN(n9643)
         );
  OAI21_X1 U11497 ( .B1(n9645), .B2(n9644), .A(n9643), .ZN(n9646) );
  INV_X1 U11498 ( .A(n9889), .ZN(n9652) );
  NAND2_X1 U11499 ( .A1(n9652), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15213) );
  INV_X1 U11500 ( .A(n15213), .ZN(n9653) );
  NAND2_X1 U11501 ( .A1(n9658), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9659) );
  MUX2_X1 U11502 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9659), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9660) );
  INV_X1 U11503 ( .A(n9661), .ZN(n9662) );
  NAND2_X1 U11504 ( .A1(n9662), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9663) );
  NAND2_X1 U11505 ( .A1(n9664), .A2(n9658), .ZN(n15207) );
  INV_X1 U11506 ( .A(n9775), .ZN(n9890) );
  NAND2_X1 U11507 ( .A1(n14825), .A2(n11665), .ZN(n9772) );
  NAND2_X1 U11508 ( .A1(n9890), .A2(n9772), .ZN(n9782) );
  NAND2_X1 U11509 ( .A1(n9873), .A2(n9782), .ZN(n9785) );
  INV_X1 U11510 ( .A(n12758), .ZN(n10111) );
  NAND2_X1 U11511 ( .A1(n10111), .A2(n9890), .ZN(n15049) );
  NOR3_X1 U11512 ( .A1(n9785), .A2(n15049), .A3(n12531), .ZN(n9668) );
  OAI21_X1 U11513 ( .B1(n15213), .B2(n15217), .A(P1_B_REG_SCAN_IN), .ZN(n9667)
         );
  OR2_X1 U11514 ( .A1(n9668), .A2(n9667), .ZN(n9669) );
  NAND2_X1 U11515 ( .A1(n9670), .A2(n9669), .ZN(P1_U3242) );
  NOR2_X1 U11516 ( .A1(n9781), .A2(P1_U3086), .ZN(n9671) );
  NAND4_X1 U11517 ( .A1(n10281), .A2(n9676), .A3(n9675), .A4(n9674), .ZN(n9677) );
  NOR2_X1 U11518 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), 
        .ZN(n9679) );
  NOR2_X1 U11519 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), 
        .ZN(n9678) );
  AND2_X1 U11520 ( .A1(n9679), .A2(n9678), .ZN(n9680) );
  INV_X1 U11521 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n9681) );
  INV_X1 U11522 ( .A(n10382), .ZN(n9684) );
  INV_X1 U11523 ( .A(n9690), .ZN(n9691) );
  NAND2_X1 U11524 ( .A1(n9691), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n9693) );
  NOR2_X1 U11525 ( .A1(n14495), .A2(n14498), .ZN(n9696) );
  NAND2_X1 U11526 ( .A1(n14490), .A2(n9696), .ZN(n10360) );
  NAND2_X1 U11527 ( .A1(n10158), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9697) );
  INV_X1 U11528 ( .A(n13051), .ZN(n9698) );
  INV_X1 U11529 ( .A(n9781), .ZN(n9713) );
  NAND2_X1 U11530 ( .A1(n9700), .A2(n14615), .ZN(n9701) );
  NAND2_X1 U11531 ( .A1(n14825), .A2(n9705), .ZN(n9703) );
  NAND2_X2 U11532 ( .A1(n9703), .A2(n9702), .ZN(n14584) );
  XNOR2_X1 U11533 ( .A(n9704), .B(n14584), .ZN(n9709) );
  AND2_X4 U11534 ( .A1(n10060), .A2(n11665), .ZN(n15796) );
  NAND2_X1 U11535 ( .A1(n15796), .A2(n14825), .ZN(n9837) );
  NAND2_X1 U11536 ( .A1(n9700), .A2(n11209), .ZN(n9707) );
  OAI21_X1 U11537 ( .B1(n9699), .B2(n9721), .A(n9707), .ZN(n9708) );
  NOR2_X1 U11538 ( .A1(n9709), .A2(n9708), .ZN(n9719) );
  INV_X2 U11539 ( .A(n14582), .ZN(n14659) );
  NAND2_X1 U11540 ( .A1(n10044), .A2(n14584), .ZN(n9717) );
  NAND2_X1 U11541 ( .A1(n9718), .A2(n9717), .ZN(n10142) );
  OAI22_X1 U11542 ( .A1(n10146), .A2(n9721), .B1(n15739), .B2(n14583), .ZN(
        n9720) );
  XNOR2_X1 U11543 ( .A(n9720), .B(n14661), .ZN(n9726) );
  OAI22_X1 U11544 ( .A1(n10146), .A2(n14613), .B1(n15739), .B2(n7189), .ZN(
        n9725) );
  XNOR2_X1 U11545 ( .A(n9726), .B(n9725), .ZN(n10427) );
  NAND2_X1 U11546 ( .A1(n14749), .A2(n14615), .ZN(n9723) );
  INV_X2 U11547 ( .A(n14583), .ZN(n14614) );
  NAND2_X1 U11548 ( .A1(n10658), .A2(n14614), .ZN(n9722) );
  NAND2_X1 U11549 ( .A1(n9723), .A2(n9722), .ZN(n9724) );
  XNOR2_X1 U11550 ( .A(n9724), .B(n14661), .ZN(n9728) );
  OAI22_X1 U11551 ( .A1(n10430), .A2(n14613), .B1(n15756), .B2(n14582), .ZN(
        n9729) );
  XNOR2_X1 U11552 ( .A(n9728), .B(n9729), .ZN(n10599) );
  NOR2_X1 U11553 ( .A1(n9726), .A2(n9725), .ZN(n10600) );
  INV_X1 U11554 ( .A(n9728), .ZN(n9731) );
  INV_X1 U11555 ( .A(n9729), .ZN(n9730) );
  NAND2_X1 U11556 ( .A1(n14748), .A2(n14607), .ZN(n9733) );
  NAND2_X1 U11557 ( .A1(n10946), .A2(n14659), .ZN(n9732) );
  NAND2_X1 U11558 ( .A1(n9733), .A2(n9732), .ZN(n9737) );
  OAI22_X1 U11559 ( .A1(n10607), .A2(n14582), .B1(n10691), .B2(n14583), .ZN(
        n9736) );
  XOR2_X1 U11560 ( .A(n14584), .B(n9736), .Z(n10945) );
  NAND2_X1 U11561 ( .A1(n14747), .A2(n14659), .ZN(n9740) );
  NAND2_X1 U11562 ( .A1(n15795), .A2(n14614), .ZN(n9739) );
  NAND2_X1 U11563 ( .A1(n9740), .A2(n9739), .ZN(n9742) );
  XNOR2_X1 U11564 ( .A(n9742), .B(n9741), .ZN(n9744) );
  AOI22_X1 U11565 ( .A1(n14747), .A2(n14607), .B1(n15795), .B2(n14659), .ZN(
        n9743) );
  NOR2_X1 U11566 ( .A1(n9744), .A2(n9743), .ZN(n10800) );
  NAND2_X1 U11567 ( .A1(n9744), .A2(n9743), .ZN(n10799) );
  NAND2_X1 U11568 ( .A1(n10995), .A2(n14614), .ZN(n9746) );
  NAND2_X1 U11569 ( .A1(n14746), .A2(n14659), .ZN(n9745) );
  NAND2_X1 U11570 ( .A1(n9746), .A2(n9745), .ZN(n9747) );
  NAND2_X1 U11571 ( .A1(n10995), .A2(n14659), .ZN(n9749) );
  NAND2_X1 U11572 ( .A1(n14746), .A2(n14607), .ZN(n9748) );
  NAND2_X1 U11573 ( .A1(n9749), .A2(n9748), .ZN(n9750) );
  NOR2_X1 U11574 ( .A1(n8088), .A2(n9750), .ZN(n9751) );
  INV_X1 U11575 ( .A(n9750), .ZN(n10992) );
  NAND2_X1 U11576 ( .A1(n15836), .A2(n14614), .ZN(n9753) );
  NAND2_X1 U11577 ( .A1(n14745), .A2(n14659), .ZN(n9752) );
  NAND2_X1 U11578 ( .A1(n9753), .A2(n9752), .ZN(n9754) );
  XNOR2_X1 U11579 ( .A(n9754), .B(n14584), .ZN(n11202) );
  AOI22_X1 U11580 ( .A1(n15836), .A2(n14659), .B1(n14607), .B2(n14745), .ZN(
        n11201) );
  XNOR2_X1 U11581 ( .A(n11202), .B(n11201), .ZN(n11204) );
  XNOR2_X1 U11582 ( .A(n11205), .B(n11204), .ZN(n9777) );
  INV_X1 U11583 ( .A(P1_B_REG_SCAN_IN), .ZN(n12530) );
  NOR2_X1 U11584 ( .A1(n15204), .A2(n12530), .ZN(n9755) );
  MUX2_X1 U11585 ( .A(n9755), .B(n12530), .S(n9757), .Z(n9756) );
  INV_X1 U11586 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9877) );
  NAND2_X1 U11587 ( .A1(n9872), .A2(n9877), .ZN(n9758) );
  NAND2_X1 U11588 ( .A1(n9758), .A2(n9875), .ZN(n9788) );
  INV_X1 U11589 ( .A(n9788), .ZN(n9833) );
  INV_X1 U11590 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9759) );
  NAND2_X1 U11591 ( .A1(n9872), .A2(n9759), .ZN(n9761) );
  NAND2_X1 U11592 ( .A1(n9761), .A2(n15193), .ZN(n10064) );
  INV_X1 U11593 ( .A(n10064), .ZN(n9834) );
  NOR4_X1 U11594 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9770) );
  NOR4_X1 U11595 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9769) );
  NOR4_X1 U11596 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n9765) );
  NOR4_X1 U11597 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n9764) );
  NOR4_X1 U11598 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n9763) );
  NOR4_X1 U11599 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n9762) );
  NAND4_X1 U11600 ( .A1(n9765), .A2(n9764), .A3(n9763), .A4(n9762), .ZN(n9766)
         );
  NOR4_X1 U11601 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n9767), .A4(n9766), .ZN(n9768) );
  NAND3_X1 U11602 ( .A1(n9770), .A2(n9769), .A3(n9768), .ZN(n9771) );
  NAND2_X1 U11603 ( .A1(n9872), .A2(n9771), .ZN(n9786) );
  NAND4_X1 U11604 ( .A1(n9833), .A2(n9834), .A3(n9873), .A4(n9786), .ZN(n9778)
         );
  INV_X1 U11605 ( .A(n10060), .ZN(n9774) );
  INV_X1 U11606 ( .A(n9772), .ZN(n9773) );
  NAND2_X1 U11607 ( .A1(n15954), .A2(n9775), .ZN(n9776) );
  NOR2_X1 U11608 ( .A1(n9777), .A2(n14733), .ZN(n9793) );
  NAND2_X1 U11609 ( .A1(n10060), .A2(n9824), .ZN(n9838) );
  OR2_X1 U11610 ( .A1(n9778), .A2(n9838), .ZN(n9779) );
  AND2_X1 U11611 ( .A1(n15836), .A2(n14731), .ZN(n9792) );
  NAND3_X1 U11612 ( .A1(n9833), .A2(n9834), .A3(n9786), .ZN(n9780) );
  NAND2_X1 U11613 ( .A1(n9780), .A2(n10063), .ZN(n9784) );
  AND3_X1 U11614 ( .A1(n9782), .A2(n9889), .A3(n9781), .ZN(n9783) );
  NAND2_X1 U11615 ( .A1(n9784), .A2(n9783), .ZN(n10045) );
  NOR2_X1 U11616 ( .A1(n16041), .A2(n11156), .ZN(n9791) );
  INV_X1 U11617 ( .A(n9785), .ZN(n9787) );
  NAND2_X1 U11618 ( .A1(n9787), .A2(n9786), .ZN(n9832) );
  NOR2_X1 U11619 ( .A1(n10065), .A2(n10064), .ZN(n14691) );
  NAND2_X1 U11620 ( .A1(n9890), .A2(n12758), .ZN(n15051) );
  INV_X2 U11621 ( .A(n15051), .ZN(n15034) );
  NAND2_X1 U11622 ( .A1(n16029), .A2(n14746), .ZN(n9789) );
  NAND2_X1 U11623 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9968) );
  OAI211_X1 U11624 ( .C1(n11376), .C2(n14728), .A(n9789), .B(n9968), .ZN(n9790) );
  OR4_X1 U11625 ( .A1(n9793), .A2(n9792), .A3(n9791), .A4(n9790), .ZN(P1_U3213) );
  NAND2_X1 U11626 ( .A1(n14750), .A2(n10061), .ZN(n10696) );
  NAND2_X1 U11627 ( .A1(n9812), .A2(n10696), .ZN(n9795) );
  NAND2_X1 U11628 ( .A1(n10431), .A2(n9699), .ZN(n9794) );
  NAND2_X1 U11629 ( .A1(n9795), .A2(n9794), .ZN(n10500) );
  NAND2_X1 U11630 ( .A1(n10500), .A2(n10504), .ZN(n9797) );
  NAND2_X1 U11631 ( .A1(n10146), .A2(n15739), .ZN(n9796) );
  NAND2_X1 U11632 ( .A1(n9797), .A2(n9796), .ZN(n10651) );
  INV_X1 U11633 ( .A(n10646), .ZN(n10652) );
  INV_X1 U11634 ( .A(n9798), .ZN(n9799) );
  AND2_X1 U11635 ( .A1(n14748), .A2(n10946), .ZN(n9800) );
  INV_X1 U11636 ( .A(n9800), .ZN(n9801) );
  NAND2_X1 U11637 ( .A1(n14747), .A2(n15795), .ZN(n9802) );
  NAND2_X1 U11638 ( .A1(n9803), .A2(n9802), .ZN(n10966) );
  INV_X1 U11639 ( .A(n10966), .ZN(n9805) );
  NAND2_X1 U11640 ( .A1(n9805), .A2(n9804), .ZN(n10968) );
  OR2_X1 U11641 ( .A1(n10995), .A2(n14746), .ZN(n9806) );
  NAND2_X1 U11642 ( .A1(n10968), .A2(n9806), .ZN(n11149) );
  OR2_X1 U11643 ( .A1(n15836), .A2(n14745), .ZN(n9807) );
  NAND2_X1 U11644 ( .A1(n9809), .A2(n9828), .ZN(n9810) );
  NAND2_X1 U11645 ( .A1(n11374), .A2(n9810), .ZN(n11338) );
  NAND2_X1 U11646 ( .A1(n7541), .A2(n15217), .ZN(n9811) );
  NAND2_X1 U11647 ( .A1(n9811), .A2(n14584), .ZN(n10685) );
  AOI22_X1 U11648 ( .A1(n15034), .A2(n14743), .B1(n14745), .B2(n15033), .ZN(
        n9831) );
  NAND2_X1 U11649 ( .A1(n10700), .A2(n10503), .ZN(n9813) );
  INV_X1 U11650 ( .A(n10504), .ZN(n10501) );
  NAND2_X1 U11651 ( .A1(n9813), .A2(n10501), .ZN(n10502) );
  NAND2_X1 U11652 ( .A1(n10502), .A2(n9814), .ZN(n10647) );
  NAND2_X1 U11653 ( .A1(n14749), .A2(n15756), .ZN(n9815) );
  NAND2_X1 U11654 ( .A1(n10430), .A2(n10658), .ZN(n9816) );
  NOR2_X1 U11655 ( .A1(n14748), .A2(n10691), .ZN(n9817) );
  INV_X1 U11656 ( .A(n15795), .ZN(n10795) );
  NAND2_X1 U11657 ( .A1(n10795), .A2(n14747), .ZN(n9819) );
  NAND2_X1 U11658 ( .A1(n9820), .A2(n9819), .ZN(n10969) );
  NAND2_X1 U11659 ( .A1(n10969), .A2(n10970), .ZN(n9822) );
  INV_X1 U11660 ( .A(n10995), .ZN(n10979) );
  NAND2_X1 U11661 ( .A1(n10979), .A2(n14746), .ZN(n9821) );
  NAND2_X1 U11662 ( .A1(n15217), .A2(n9348), .ZN(n9827) );
  NAND2_X1 U11663 ( .A1(n9825), .A2(n9824), .ZN(n9826) );
  OAI211_X1 U11664 ( .C1(n9829), .C2(n9828), .A(n11379), .B(n15985), .ZN(n9830) );
  OAI211_X1 U11665 ( .C1(n11338), .C2(n10764), .A(n9831), .B(n9830), .ZN(
        n11341) );
  OR2_X1 U11666 ( .A1(n9833), .A2(n9832), .ZN(n10763) );
  INV_X1 U11667 ( .A(n10763), .ZN(n9835) );
  NAND2_X1 U11668 ( .A1(n9835), .A2(n9834), .ZN(n12534) );
  MUX2_X1 U11669 ( .A(n11341), .B(P1_REG2_REG_8__SCAN_IN), .S(n15036), .Z(
        n9842) );
  OR2_X1 U11670 ( .A1(n15036), .A2(n9836), .ZN(n11391) );
  NOR2_X1 U11671 ( .A1(n11338), .A2(n11391), .ZN(n9841) );
  NAND3_X1 U11672 ( .A1(n15739), .A2(n9699), .A3(n15679), .ZN(n10654) );
  NAND2_X1 U11673 ( .A1(n10689), .A2(n10691), .ZN(n10793) );
  OR2_X1 U11674 ( .A1(n10793), .A2(n15795), .ZN(n10978) );
  OR2_X1 U11675 ( .A1(n10978), .A2(n10995), .ZN(n11153) );
  OAI21_X1 U11676 ( .B1(n11152), .B2(n11339), .A(n11386), .ZN(n11340) );
  NOR2_X1 U11677 ( .A1(n11340), .A2(n15681), .ZN(n9840) );
  OAI22_X1 U11678 ( .A1(n11339), .A2(n15680), .B1(n11217), .B2(n15035), .ZN(
        n9839) );
  INV_X4 U11679 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U11680 ( .A(n13796), .ZN(n9843) );
  INV_X2 U11681 ( .A(n15212), .ZN(n15210) );
  OAI222_X1 U11682 ( .A1(n15210), .A2(n9844), .B1(n15215), .B2(n10449), .C1(
        n9953), .C2(P1_U3086), .ZN(P1_U3353) );
  AND2_X1 U11683 ( .A1(n10404), .A2(P2_U3088), .ZN(n14500) );
  INV_X2 U11684 ( .A(n14500), .ZN(n14506) );
  MUX2_X1 U11685 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9845), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n9848) );
  INV_X1 U11686 ( .A(n9846), .ZN(n9847) );
  OAI222_X1 U11687 ( .A1(n14506), .A2(n10397), .B1(n14503), .B2(n10396), .C1(
        P2_U3088), .C2(n10398), .ZN(P2_U3326) );
  OAI222_X1 U11688 ( .A1(n15210), .A2(n9849), .B1(n15215), .B2(n9870), .C1(
        n8984), .C2(P1_U3086), .ZN(P1_U3352) );
  OAI222_X1 U11689 ( .A1(P1_U3086), .A2(n9950), .B1(n15215), .B2(n10397), .C1(
        n7363), .C2(n15210), .ZN(P1_U3354) );
  NAND2_X2 U11690 ( .A1(n10404), .A2(P3_U3151), .ZN(n13810) );
  INV_X1 U11691 ( .A(n9850), .ZN(n9851) );
  OAI222_X1 U11692 ( .A1(P3_U3151), .A2(n11461), .B1(n13810), .B2(n7413), .C1(
        n12036), .C2(n9851), .ZN(P3_U3288) );
  INV_X1 U11693 ( .A(n14782), .ZN(n9853) );
  INV_X1 U11694 ( .A(n10534), .ZN(n9864) );
  OAI222_X1 U11695 ( .A1(P1_U3086), .A2(n9853), .B1(n15215), .B2(n9864), .C1(
        n9852), .C2(n15210), .ZN(P1_U3351) );
  OAI222_X1 U11696 ( .A1(n10275), .A2(P3_U3151), .B1(n12036), .B2(n9855), .C1(
        n9854), .C2(n13810), .ZN(P3_U3294) );
  NAND2_X1 U11697 ( .A1(n9856), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9857) );
  XNOR2_X1 U11698 ( .A(n9857), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10550) );
  INV_X1 U11699 ( .A(n10550), .ZN(n9858) );
  OAI222_X1 U11700 ( .A1(n14503), .A2(n9859), .B1(n14506), .B2(n10549), .C1(
        n9858), .C2(P2_U3088), .ZN(P2_U3322) );
  INV_X1 U11701 ( .A(n9961), .ZN(n9985) );
  OAI222_X1 U11702 ( .A1(n15210), .A2(n9860), .B1(n15215), .B2(n10549), .C1(
        n9985), .C2(P1_U3086), .ZN(P1_U3350) );
  INV_X1 U11703 ( .A(n14503), .ZN(n11927) );
  INV_X1 U11704 ( .A(n11927), .ZN(n14509) );
  OR2_X1 U11705 ( .A1(n9861), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n9867) );
  NAND2_X1 U11706 ( .A1(n9867), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9862) );
  XNOR2_X1 U11707 ( .A(n9862), .B(P2_IR_REG_4__SCAN_IN), .ZN(n15372) );
  INV_X1 U11708 ( .A(n15372), .ZN(n9863) );
  OAI222_X1 U11709 ( .A1(n14509), .A2(n9865), .B1(n14506), .B2(n9864), .C1(
        n9863), .C2(P2_U3088), .ZN(P2_U3323) );
  NAND2_X1 U11710 ( .A1(n9861), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9866) );
  MUX2_X1 U11711 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9866), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n9868) );
  INV_X1 U11712 ( .A(n15361), .ZN(n9869) );
  OAI222_X1 U11713 ( .A1(n14509), .A2(n9871), .B1(n14506), .B2(n9870), .C1(
        n9869), .C2(P2_U3088), .ZN(P2_U3324) );
  INV_X1 U11714 ( .A(n9872), .ZN(n9874) );
  NAND2_X1 U11715 ( .A1(n9874), .A2(n9873), .ZN(n15332) );
  INV_X1 U11716 ( .A(n15332), .ZN(n9878) );
  NAND2_X1 U11717 ( .A1(n9878), .A2(n9875), .ZN(n9876) );
  OAI21_X1 U11718 ( .B1(n9878), .B2(n9877), .A(n9876), .ZN(P1_U3445) );
  OR2_X1 U11719 ( .A1(n9846), .A2(n11039), .ZN(n9880) );
  OAI222_X1 U11720 ( .A1(P2_U3088), .A2(n10447), .B1(n14506), .B2(n10449), 
        .C1(n10446), .C2(n14509), .ZN(P2_U3325) );
  INV_X1 U11721 ( .A(n9963), .ZN(n9998) );
  OAI222_X1 U11722 ( .A1(P1_U3086), .A2(n9998), .B1(n15215), .B2(n10565), .C1(
        n9881), .C2(n15210), .ZN(P1_U3349) );
  NOR2_X1 U11723 ( .A1(n9856), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n9927) );
  OR2_X1 U11724 ( .A1(n9927), .A2(n11039), .ZN(n9882) );
  XNOR2_X1 U11725 ( .A(n9882), .B(P2_IR_REG_6__SCAN_IN), .ZN(n15384) );
  INV_X1 U11726 ( .A(n15384), .ZN(n9884) );
  OAI222_X1 U11727 ( .A1(P2_U3088), .A2(n9884), .B1(n14506), .B2(n10565), .C1(
        n9883), .C2(n14503), .ZN(P2_U3321) );
  INV_X1 U11728 ( .A(n12531), .ZN(n9885) );
  AOI21_X1 U11729 ( .B1(n9885), .B2(n8951), .A(n12758), .ZN(n10109) );
  OAI21_X1 U11730 ( .B1(n9885), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10109), .ZN(
        n9887) );
  XNOR2_X1 U11731 ( .A(n9887), .B(n9886), .ZN(n9898) );
  NAND2_X1 U11732 ( .A1(n9888), .A2(n15213), .ZN(n9895) );
  NAND2_X1 U11733 ( .A1(n9890), .A2(n9889), .ZN(n9892) );
  NAND2_X1 U11734 ( .A1(n9892), .A2(n9891), .ZN(n9894) );
  INV_X1 U11735 ( .A(n9894), .ZN(n9893) );
  INV_X1 U11736 ( .A(n9949), .ZN(n9897) );
  AND2_X1 U11737 ( .A1(n9895), .A2(n9894), .ZN(n14791) );
  AOI22_X1 U11738 ( .A1(n14791), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9896) );
  OAI21_X1 U11739 ( .B1(n9898), .B2(n9897), .A(n9896), .ZN(P1_U3243) );
  INV_X1 U11740 ( .A(SI_10_), .ZN(n9901) );
  INV_X1 U11741 ( .A(n9899), .ZN(n9900) );
  OAI222_X1 U11742 ( .A1(P3_U3151), .A2(n15658), .B1(n13810), .B2(n9901), .C1(
        n12036), .C2(n9900), .ZN(P3_U3285) );
  INV_X1 U11743 ( .A(n15540), .ZN(n11414) );
  INV_X1 U11744 ( .A(SI_4_), .ZN(n9904) );
  INV_X1 U11745 ( .A(n9902), .ZN(n9903) );
  OAI222_X1 U11746 ( .A1(P3_U3151), .A2(n11414), .B1(n13810), .B2(n9904), .C1(
        n12036), .C2(n9903), .ZN(P3_U3291) );
  OAI222_X1 U11747 ( .A1(n12036), .A2(n9906), .B1(n13810), .B2(n9905), .C1(
        P3_U3151), .C2(n15617), .ZN(P3_U3287) );
  INV_X1 U11748 ( .A(n9907), .ZN(n9908) );
  OAI222_X1 U11749 ( .A1(P3_U3151), .A2(n15637), .B1(n13810), .B2(n7427), .C1(
        n12036), .C2(n9908), .ZN(P3_U3286) );
  INV_X1 U11750 ( .A(n9909), .ZN(n9910) );
  OAI222_X1 U11751 ( .A1(P3_U3151), .A2(n7674), .B1(n13810), .B2(n9911), .C1(
        n12036), .C2(n9910), .ZN(P3_U3293) );
  INV_X1 U11752 ( .A(SI_3_), .ZN(n9914) );
  INV_X1 U11753 ( .A(n9912), .ZN(n9913) );
  OAI222_X1 U11754 ( .A1(P3_U3151), .A2(n11456), .B1(n13810), .B2(n9914), .C1(
        n12036), .C2(n9913), .ZN(P3_U3292) );
  INV_X1 U11755 ( .A(SI_5_), .ZN(n9917) );
  INV_X1 U11756 ( .A(n9915), .ZN(n9916) );
  OAI222_X1 U11757 ( .A1(P3_U3151), .A2(n7678), .B1(n13810), .B2(n9917), .C1(
        n12036), .C2(n9916), .ZN(P3_U3290) );
  INV_X1 U11758 ( .A(n9918), .ZN(n9919) );
  OAI222_X1 U11759 ( .A1(P3_U3151), .A2(n11674), .B1(n13810), .B2(n9920), .C1(
        n12036), .C2(n9919), .ZN(P3_U3284) );
  INV_X1 U11760 ( .A(n9921), .ZN(n9922) );
  OAI222_X1 U11761 ( .A1(n13276), .A2(P3_U3151), .B1(n12036), .B2(n9922), .C1(
        n13810), .C2(n11850), .ZN(P3_U3283) );
  OAI222_X1 U11762 ( .A1(P3_U3151), .A2(n11460), .B1(n12036), .B2(n9924), .C1(
        n9923), .C2(n13810), .ZN(P3_U3289) );
  INV_X1 U11763 ( .A(n10726), .ZN(n9929) );
  INV_X1 U11764 ( .A(n10003), .ZN(n10007) );
  OAI222_X1 U11765 ( .A1(n15210), .A2(n9925), .B1(n15215), .B2(n9929), .C1(
        P1_U3086), .C2(n10007), .ZN(P1_U3348) );
  INV_X1 U11766 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U11767 ( .A1(n9927), .A2(n9926), .ZN(n10283) );
  NAND2_X1 U11768 ( .A1(n10283), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9928) );
  XNOR2_X1 U11769 ( .A(n9928), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10727) );
  INV_X1 U11770 ( .A(n10727), .ZN(n10204) );
  OAI222_X1 U11771 ( .A1(n14509), .A2(n9930), .B1(n14506), .B2(n9929), .C1(
        P2_U3088), .C2(n10204), .ZN(P2_U3320) );
  NAND2_X1 U11772 ( .A1(n9931), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10036) );
  XNOR2_X1 U11773 ( .A(n10036), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10912) );
  INV_X1 U11774 ( .A(n10912), .ZN(n9932) );
  OAI222_X1 U11775 ( .A1(n14509), .A2(n9933), .B1(n14506), .B2(n10911), .C1(
        n9932), .C2(P2_U3088), .ZN(P2_U3319) );
  OAI222_X1 U11776 ( .A1(n15210), .A2(n9934), .B1(n15215), .B2(n10911), .C1(
        n7666), .C2(P1_U3086), .ZN(P1_U3347) );
  INV_X1 U11777 ( .A(n10615), .ZN(n9935) );
  NAND2_X1 U11778 ( .A1(n9935), .A2(n13796), .ZN(n9936) );
  OAI21_X1 U11779 ( .B1(n13796), .B2(n8823), .A(n9936), .ZN(P3_U3376) );
  OAI222_X1 U11780 ( .A1(P3_U3151), .A2(n13299), .B1(n13810), .B2(n11848), 
        .C1(n12036), .C2(n9937), .ZN(P3_U3282) );
  AND2_X1 U11781 ( .A1(n9938), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U11782 ( .A1(n9938), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U11783 ( .A1(n9938), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U11784 ( .A1(n9938), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U11785 ( .A1(n9938), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U11786 ( .A1(n9938), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U11787 ( .A1(n9938), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U11788 ( .A1(n9938), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U11789 ( .A1(n9938), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U11790 ( .A1(n9938), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U11791 ( .A1(n9938), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U11792 ( .A1(n9938), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U11793 ( .A1(n9938), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U11794 ( .A1(n9938), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U11795 ( .A1(n9938), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U11796 ( .A1(n9938), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U11797 ( .A1(n9938), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U11798 ( .A1(n9938), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U11799 ( .A1(n9938), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U11800 ( .A1(n9938), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U11801 ( .A1(n9938), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U11802 ( .A1(n9938), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U11803 ( .A1(n9938), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U11804 ( .A1(n9938), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U11805 ( .A1(n9938), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U11806 ( .A1(n9938), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U11807 ( .A1(n9938), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U11808 ( .A1(n9938), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U11809 ( .A1(n9938), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U11810 ( .A1(n9938), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  NOR2_X1 U11811 ( .A1(n14791), .A2(P1_U4016), .ZN(P1_U3085) );
  XNOR2_X1 U11812 ( .A(n9950), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n14753) );
  AND2_X1 U11813 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14752) );
  NAND2_X1 U11814 ( .A1(n14753), .A2(n14752), .ZN(n14751) );
  NAND2_X1 U11815 ( .A1(n14757), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9939) );
  NAND2_X1 U11816 ( .A1(n14751), .A2(n9939), .ZN(n10116) );
  XNOR2_X1 U11817 ( .A(n9953), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n10117) );
  NAND2_X1 U11818 ( .A1(n10116), .A2(n10117), .ZN(n10115) );
  NAND2_X1 U11819 ( .A1(n10118), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9940) );
  NAND2_X1 U11820 ( .A1(n10115), .A2(n9940), .ZN(n14763) );
  INV_X1 U11821 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9941) );
  XNOR2_X1 U11822 ( .A(n14766), .B(n9941), .ZN(n14764) );
  NAND2_X1 U11823 ( .A1(n14763), .A2(n14764), .ZN(n14762) );
  NAND2_X1 U11824 ( .A1(n14766), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9942) );
  NAND2_X1 U11825 ( .A1(n14762), .A2(n9942), .ZN(n14785) );
  INV_X1 U11826 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10772) );
  MUX2_X1 U11827 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10772), .S(n14782), .Z(
        n14786) );
  AND2_X1 U11828 ( .A1(n14785), .A2(n14786), .ZN(n14783) );
  AOI21_X1 U11829 ( .B1(n14782), .B2(P1_REG1_REG_4__SCAN_IN), .A(n14783), .ZN(
        n9976) );
  INV_X1 U11830 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9943) );
  MUX2_X1 U11831 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9943), .S(n9961), .Z(n9975)
         );
  INV_X1 U11832 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9944) );
  MUX2_X1 U11833 ( .A(n9944), .B(P1_REG1_REG_6__SCAN_IN), .S(n9963), .Z(n9995)
         );
  INV_X1 U11834 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9945) );
  MUX2_X1 U11835 ( .A(n9945), .B(P1_REG1_REG_7__SCAN_IN), .S(n10003), .Z(n9946) );
  NAND2_X1 U11836 ( .A1(n9949), .A2(n12531), .ZN(n14823) );
  NOR2_X1 U11837 ( .A1(n9947), .A2(n9946), .ZN(n10002) );
  AOI211_X1 U11838 ( .C1(n9947), .C2(n9946), .A(n14823), .B(n10002), .ZN(n9973) );
  NAND2_X1 U11839 ( .A1(n9949), .A2(n12758), .ZN(n15432) );
  NOR2_X1 U11840 ( .A1(n12758), .A2(n12531), .ZN(n9948) );
  MUX2_X1 U11841 ( .A(n9951), .B(P1_REG2_REG_1__SCAN_IN), .S(n9950), .Z(n14755) );
  AND2_X1 U11842 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14756) );
  NAND2_X1 U11843 ( .A1(n14755), .A2(n14756), .ZN(n14754) );
  NAND2_X1 U11844 ( .A1(n14757), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U11845 ( .A1(n14754), .A2(n9952), .ZN(n10113) );
  MUX2_X1 U11846 ( .A(n9954), .B(P1_REG2_REG_2__SCAN_IN), .S(n9953), .Z(n10114) );
  NAND2_X1 U11847 ( .A1(n10113), .A2(n10114), .ZN(n14768) );
  NAND2_X1 U11848 ( .A1(n10118), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14767) );
  NAND2_X1 U11849 ( .A1(n14768), .A2(n14767), .ZN(n9957) );
  MUX2_X1 U11850 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9955), .S(n14766), .Z(n9956) );
  NAND2_X1 U11851 ( .A1(n9957), .A2(n9956), .ZN(n14778) );
  NAND2_X1 U11852 ( .A1(n14766), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14777) );
  NAND2_X1 U11853 ( .A1(n14778), .A2(n14777), .ZN(n9960) );
  MUX2_X1 U11854 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9958), .S(n14782), .Z(n9959) );
  NAND2_X1 U11855 ( .A1(n9960), .A2(n9959), .ZN(n14780) );
  NAND2_X1 U11856 ( .A1(n14782), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9978) );
  MUX2_X1 U11857 ( .A(n9032), .B(P1_REG2_REG_5__SCAN_IN), .S(n9961), .Z(n9977)
         );
  AOI21_X1 U11858 ( .B1(n14780), .B2(n9978), .A(n9977), .ZN(n9990) );
  NOR2_X1 U11859 ( .A1(n9985), .A2(n9032), .ZN(n9989) );
  MUX2_X1 U11860 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9962), .S(n9963), .Z(n9988)
         );
  OAI21_X1 U11861 ( .B1(n9990), .B2(n9989), .A(n9988), .ZN(n9987) );
  NAND2_X1 U11862 ( .A1(n9963), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9965) );
  MUX2_X1 U11863 ( .A(n10006), .B(P1_REG2_REG_7__SCAN_IN), .S(n10003), .Z(
        n9964) );
  AOI21_X1 U11864 ( .B1(n9987), .B2(n9965), .A(n9964), .ZN(n10011) );
  INV_X1 U11865 ( .A(n10011), .ZN(n9967) );
  NAND3_X1 U11866 ( .A1(n9987), .A2(n9965), .A3(n9964), .ZN(n9966) );
  NAND3_X1 U11867 ( .A1(n14819), .A2(n9967), .A3(n9966), .ZN(n9971) );
  INV_X1 U11868 ( .A(n9968), .ZN(n9969) );
  AOI21_X1 U11869 ( .B1(n14791), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9969), .ZN(
        n9970) );
  OAI211_X1 U11870 ( .C1(n15432), .C2(n10007), .A(n9971), .B(n9970), .ZN(n9972) );
  OR2_X1 U11871 ( .A1(n9973), .A2(n9972), .ZN(P1_U3250) );
  INV_X1 U11872 ( .A(n14823), .ZN(n15437) );
  OAI21_X1 U11873 ( .B1(n9976), .B2(n9975), .A(n9974), .ZN(n9981) );
  AND3_X1 U11874 ( .A1(n14780), .A2(n9978), .A3(n9977), .ZN(n9979) );
  NOR3_X1 U11875 ( .A1(n15434), .A2(n9990), .A3(n9979), .ZN(n9980) );
  AOI21_X1 U11876 ( .B1(n15437), .B2(n9981), .A(n9980), .ZN(n9984) );
  NAND2_X1 U11877 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n10805) );
  INV_X1 U11878 ( .A(n10805), .ZN(n9982) );
  AOI21_X1 U11879 ( .B1(n14791), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n9982), .ZN(
        n9983) );
  OAI211_X1 U11880 ( .C1(n9985), .C2(n15432), .A(n9984), .B(n9983), .ZN(
        P1_U3248) );
  OAI222_X1 U11881 ( .A1(n13321), .A2(P3_U3151), .B1(n12036), .B2(n9986), .C1(
        n13810), .C2(n11818), .ZN(P3_U3281) );
  INV_X1 U11882 ( .A(n9987), .ZN(n9992) );
  NOR3_X1 U11883 ( .A1(n9990), .A2(n9989), .A3(n9988), .ZN(n9991) );
  NOR3_X1 U11884 ( .A1(n15434), .A2(n9992), .A3(n9991), .ZN(n10001) );
  AOI211_X1 U11885 ( .C1(n9995), .C2(n9994), .A(n9993), .B(n14823), .ZN(n10000) );
  AND2_X1 U11886 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9996) );
  AOI21_X1 U11887 ( .B1(n14791), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n9996), .ZN(
        n9997) );
  OAI21_X1 U11888 ( .B1(n15432), .B2(n9998), .A(n9997), .ZN(n9999) );
  OR3_X1 U11889 ( .A1(n10001), .A2(n10000), .A3(n9999), .ZN(P1_U3249) );
  MUX2_X1 U11890 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n7665), .S(n10024), .Z(
        n10004) );
  OAI21_X1 U11891 ( .B1(n10005), .B2(n10004), .A(n10021), .ZN(n10018) );
  NOR2_X1 U11892 ( .A1(n10007), .A2(n10006), .ZN(n10010) );
  MUX2_X1 U11893 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10008), .S(n10024), .Z(
        n10009) );
  OAI21_X1 U11894 ( .B1(n10011), .B2(n10010), .A(n10009), .ZN(n10028) );
  INV_X1 U11895 ( .A(n10028), .ZN(n10013) );
  NOR3_X1 U11896 ( .A1(n10011), .A2(n10010), .A3(n10009), .ZN(n10012) );
  NOR3_X1 U11897 ( .A1(n15434), .A2(n10013), .A3(n10012), .ZN(n10017) );
  NAND2_X1 U11898 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11218) );
  INV_X1 U11899 ( .A(n11218), .ZN(n10014) );
  AOI21_X1 U11900 ( .B1(n14791), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n10014), .ZN(
        n10015) );
  OAI21_X1 U11901 ( .B1(n15432), .B2(n7666), .A(n10015), .ZN(n10016) );
  AOI211_X1 U11902 ( .C1(n10018), .C2(n15437), .A(n10017), .B(n10016), .ZN(
        n10019) );
  INV_X1 U11903 ( .A(n10019), .ZN(P1_U3251) );
  INV_X1 U11904 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10020) );
  MUX2_X1 U11905 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10020), .S(n10069), .Z(
        n10023) );
  OAI21_X1 U11906 ( .B1(n10023), .B2(n10022), .A(n10068), .ZN(n10033) );
  NAND2_X1 U11907 ( .A1(n10024), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10027) );
  INV_X1 U11908 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10025) );
  MUX2_X1 U11909 ( .A(n10025), .B(P1_REG2_REG_9__SCAN_IN), .S(n10069), .Z(
        n10026) );
  AOI21_X1 U11910 ( .B1(n10028), .B2(n10027), .A(n10026), .ZN(n10075) );
  AND3_X1 U11911 ( .A1(n10028), .A2(n10027), .A3(n10026), .ZN(n10029) );
  NOR3_X1 U11912 ( .A1(n10075), .A2(n15434), .A3(n10029), .ZN(n10032) );
  INV_X1 U11913 ( .A(n10069), .ZN(n10072) );
  NAND2_X1 U11914 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n11261) );
  NAND2_X1 U11915 ( .A1(n14791), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n10030) );
  OAI211_X1 U11916 ( .C1(n15432), .C2(n10072), .A(n11261), .B(n10030), .ZN(
        n10031) );
  AOI211_X1 U11917 ( .C1(n10033), .C2(n15437), .A(n10032), .B(n10031), .ZN(
        n10034) );
  INV_X1 U11918 ( .A(n10034), .ZN(P1_U3252) );
  INV_X1 U11919 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n10035) );
  NAND2_X1 U11920 ( .A1(n10036), .A2(n10035), .ZN(n10037) );
  NAND2_X1 U11921 ( .A1(n10037), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10050) );
  XNOR2_X1 U11922 ( .A(n10050), .B(P2_IR_REG_9__SCAN_IN), .ZN(n11068) );
  INV_X1 U11923 ( .A(n11068), .ZN(n10038) );
  OAI222_X1 U11924 ( .A1(n14503), .A2(n10039), .B1(n14506), .B2(n11067), .C1(
        n10038), .C2(P2_U3088), .ZN(P2_U3318) );
  OAI222_X1 U11925 ( .A1(n15210), .A2(n10040), .B1(n15215), .B2(n11067), .C1(
        n10072), .C2(P1_U3086), .ZN(P1_U3346) );
  OAI222_X1 U11926 ( .A1(n13340), .A2(P3_U3151), .B1(n12036), .B2(n10041), 
        .C1(n13810), .C2(n11711), .ZN(P3_U3280) );
  INV_X1 U11927 ( .A(n13348), .ZN(n13372) );
  OAI222_X1 U11928 ( .A1(n13810), .A2(n11845), .B1(n12036), .B2(n10042), .C1(
        n13372), .C2(P3_U3151), .ZN(P3_U3279) );
  XNOR2_X1 U11929 ( .A(n10044), .B(n10043), .ZN(n10108) );
  AND2_X1 U11930 ( .A1(n9700), .A2(n15034), .ZN(n10057) );
  AOI22_X1 U11931 ( .A1(n14691), .A2(n10057), .B1(n14731), .B2(n10061), .ZN(
        n10048) );
  NOR2_X1 U11932 ( .A1(n10045), .A2(P1_U3086), .ZN(n10429) );
  INV_X1 U11933 ( .A(n10429), .ZN(n10046) );
  NAND2_X1 U11934 ( .A1(n10046), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n10047) );
  OAI211_X1 U11935 ( .C1(n10108), .C2(n14733), .A(n10048), .B(n10047), .ZN(
        P1_U3232) );
  INV_X1 U11936 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n10049) );
  NAND2_X1 U11937 ( .A1(n10050), .A2(n10049), .ZN(n10051) );
  NAND2_X1 U11938 ( .A1(n10051), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10052) );
  NAND2_X1 U11939 ( .A1(n10052), .A2(n10278), .ZN(n10085) );
  OR2_X1 U11940 ( .A1(n10052), .A2(n10278), .ZN(n10053) );
  INV_X1 U11941 ( .A(n11124), .ZN(n10054) );
  OAI222_X1 U11942 ( .A1(n14503), .A2(n10055), .B1(n14506), .B2(n11123), .C1(
        n10054), .C2(P2_U3088), .ZN(P2_U3317) );
  INV_X1 U11943 ( .A(n10095), .ZN(n10079) );
  OAI222_X1 U11944 ( .A1(P1_U3086), .A2(n10079), .B1(n15215), .B2(n11123), 
        .C1(n10056), .C2(n15210), .ZN(P1_U3345) );
  NAND2_X1 U11945 ( .A1(n10764), .A2(n16016), .ZN(n10058) );
  AOI21_X1 U11946 ( .B1(n15683), .B2(n10058), .A(n10057), .ZN(n15687) );
  NAND2_X1 U11947 ( .A1(n9348), .A2(n11665), .ZN(n10059) );
  INV_X1 U11948 ( .A(n10987), .ZN(n15881) );
  AOI22_X1 U11949 ( .A1(n15683), .A2(n15881), .B1(n10061), .B2(n10060), .ZN(
        n10062) );
  AND2_X1 U11950 ( .A1(n15687), .A2(n10062), .ZN(n15677) );
  NAND2_X1 U11951 ( .A1(n10064), .A2(n10063), .ZN(n10762) );
  NAND2_X1 U11952 ( .A1(n16021), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10066) );
  OAI21_X1 U11953 ( .B1(n15677), .B2(n16021), .A(n10066), .ZN(P1_U3528) );
  INV_X1 U11954 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10067) );
  MUX2_X1 U11955 ( .A(n10067), .B(P1_REG1_REG_10__SCAN_IN), .S(n10095), .Z(
        n10071) );
  OAI21_X1 U11956 ( .B1(n10069), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10068), .ZN(
        n10070) );
  NOR2_X1 U11957 ( .A1(n10070), .A2(n10071), .ZN(n10094) );
  AOI211_X1 U11958 ( .C1(n10071), .C2(n10070), .A(n14823), .B(n10094), .ZN(
        n10082) );
  NOR2_X1 U11959 ( .A1(n10072), .A2(n10025), .ZN(n10074) );
  MUX2_X1 U11960 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11493), .S(n10095), .Z(
        n10073) );
  OAI21_X1 U11961 ( .B1(n10075), .B2(n10074), .A(n10073), .ZN(n10092) );
  INV_X1 U11962 ( .A(n10092), .ZN(n10077) );
  NOR3_X1 U11963 ( .A1(n10075), .A2(n10074), .A3(n10073), .ZN(n10076) );
  NOR3_X1 U11964 ( .A1(n10077), .A2(n10076), .A3(n15434), .ZN(n10081) );
  AND2_X1 U11965 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11510) );
  AOI21_X1 U11966 ( .B1(n14791), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n11510), 
        .ZN(n10078) );
  OAI21_X1 U11967 ( .B1(n15432), .B2(n10079), .A(n10078), .ZN(n10080) );
  OR3_X1 U11968 ( .A1(n10082), .A2(n10081), .A3(n10080), .ZN(P1_U3253) );
  OAI222_X1 U11969 ( .A1(n13379), .A2(P3_U3151), .B1(n12036), .B2(n10083), 
        .C1(n13810), .C2(n11840), .ZN(P3_U3278) );
  INV_X1 U11970 ( .A(n11298), .ZN(n10088) );
  INV_X1 U11971 ( .A(n10241), .ZN(n10100) );
  OAI222_X1 U11972 ( .A1(n15210), .A2(n10084), .B1(n15215), .B2(n10088), .C1(
        P1_U3086), .C2(n10100), .ZN(P1_U3344) );
  NAND2_X1 U11973 ( .A1(n10085), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10086) );
  XNOR2_X1 U11974 ( .A(n10086), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11361) );
  INV_X1 U11975 ( .A(n11361), .ZN(n10087) );
  OAI222_X1 U11976 ( .A1(n14503), .A2(n10089), .B1(n14506), .B2(n10088), .C1(
        P2_U3088), .C2(n10087), .ZN(P2_U3316) );
  NAND2_X1 U11977 ( .A1(n10095), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10091) );
  MUX2_X1 U11978 ( .A(n9158), .B(P1_REG2_REG_11__SCAN_IN), .S(n10241), .Z(
        n10090) );
  AOI21_X1 U11979 ( .B1(n10092), .B2(n10091), .A(n10090), .ZN(n10240) );
  NAND3_X1 U11980 ( .A1(n10092), .A2(n10091), .A3(n10090), .ZN(n10093) );
  NAND2_X1 U11981 ( .A1(n10093), .A2(n14819), .ZN(n10105) );
  INV_X1 U11982 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10096) );
  MUX2_X1 U11983 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10096), .S(n10241), .Z(
        n10097) );
  OAI21_X1 U11984 ( .B1(n10098), .B2(n10097), .A(n10237), .ZN(n10099) );
  NAND2_X1 U11985 ( .A1(n10099), .A2(n15437), .ZN(n10104) );
  NAND2_X1 U11986 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n11936)
         );
  INV_X1 U11987 ( .A(n11936), .ZN(n10102) );
  NOR2_X1 U11988 ( .A1(n15432), .A2(n10100), .ZN(n10101) );
  AOI211_X1 U11989 ( .C1(n14791), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10102), 
        .B(n10101), .ZN(n10103) );
  OAI211_X1 U11990 ( .C1(n10240), .C2(n10105), .A(n10104), .B(n10103), .ZN(
        P1_U3254) );
  INV_X1 U11991 ( .A(n13405), .ZN(n10107) );
  OAI222_X1 U11992 ( .A1(P3_U3151), .A2(n10107), .B1(n13810), .B2(n11833), 
        .C1(n12036), .C2(n10106), .ZN(P3_U3277) );
  MUX2_X1 U11993 ( .A(n14756), .B(n10108), .S(n12531), .Z(n10112) );
  OAI21_X1 U11994 ( .B1(n10109), .B2(P1_IR_REG_0__SCAN_IN), .A(P1_U4016), .ZN(
        n10110) );
  AOI21_X1 U11995 ( .B1(n10112), .B2(n10111), .A(n10110), .ZN(n14775) );
  AOI22_X1 U11996 ( .A1(n14791), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10122) );
  OAI211_X1 U11997 ( .C1(n10114), .C2(n10113), .A(n14819), .B(n14768), .ZN(
        n10121) );
  OAI211_X1 U11998 ( .C1(n10117), .C2(n10116), .A(n15437), .B(n10115), .ZN(
        n10120) );
  INV_X1 U11999 ( .A(n15432), .ZN(n14795) );
  NAND2_X1 U12000 ( .A1(n14795), .A2(n10118), .ZN(n10119) );
  NAND4_X1 U12001 ( .A1(n10122), .A2(n10121), .A3(n10120), .A4(n10119), .ZN(
        n10123) );
  OR2_X1 U12002 ( .A1(n14775), .A2(n10123), .ZN(P1_U3245) );
  INV_X1 U12003 ( .A(n10335), .ZN(n10124) );
  NAND2_X1 U12004 ( .A1(n10126), .A2(n10125), .ZN(n10134) );
  OR2_X1 U12005 ( .A1(n10335), .A2(P3_U3151), .ZN(n12756) );
  INV_X1 U12006 ( .A(n12756), .ZN(n10127) );
  NOR2_X1 U12007 ( .A1(n10355), .A2(n10127), .ZN(n10133) );
  OR2_X1 U12008 ( .A1(n10134), .A2(n10133), .ZN(n10136) );
  INV_X1 U12009 ( .A(n15671), .ZN(n13368) );
  OR2_X1 U12010 ( .A1(n10136), .A2(n10129), .ZN(n15583) );
  NOR3_X1 U12011 ( .A1(n13368), .A2(n15667), .A3(n13412), .ZN(n10141) );
  MUX2_X1 U12012 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n13408), .Z(n10132) );
  INV_X1 U12013 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10593) );
  INV_X1 U12014 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10130) );
  MUX2_X1 U12015 ( .A(n10593), .B(n10130), .S(n13408), .Z(n10131) );
  NAND2_X1 U12016 ( .A1(n10131), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10256) );
  INV_X1 U12017 ( .A(n10256), .ZN(n10258) );
  AOI21_X1 U12018 ( .B1(n10263), .B2(n10132), .A(n10258), .ZN(n10140) );
  INV_X1 U12019 ( .A(n10133), .ZN(n10135) );
  AOI22_X1 U12020 ( .A1(n15663), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n10139) );
  INV_X1 U12021 ( .A(n10136), .ZN(n10137) );
  MUX2_X1 U12022 ( .A(P3_U3897), .B(n10137), .S(n8787), .Z(n15602) );
  NAND2_X1 U12023 ( .A1(n15602), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10138) );
  OAI211_X1 U12024 ( .C1(n10141), .C2(n10140), .A(n10139), .B(n10138), .ZN(
        P3_U3182) );
  NOR2_X1 U12025 ( .A1(n10143), .A2(n10142), .ZN(n10145) );
  OAI21_X1 U12026 ( .B1(n10145), .B2(n10144), .A(n16036), .ZN(n10150) );
  INV_X1 U12027 ( .A(n16029), .ZN(n14701) );
  INV_X1 U12028 ( .A(n14750), .ZN(n10147) );
  OAI22_X1 U12029 ( .A1(n14701), .A2(n10147), .B1(n10146), .B2(n14728), .ZN(
        n10148) );
  AOI21_X1 U12030 ( .B1(n10697), .B2(n14731), .A(n10148), .ZN(n10149) );
  OAI211_X1 U12031 ( .C1(n10429), .C2(n8935), .A(n10150), .B(n10149), .ZN(
        P1_U3222) );
  INV_X1 U12032 ( .A(n10447), .ZN(n10226) );
  INV_X1 U12033 ( .A(n10398), .ZN(n15350) );
  INV_X1 U12034 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10151) );
  XNOR2_X1 U12035 ( .A(n10398), .B(n10151), .ZN(n15343) );
  INV_X1 U12036 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10152) );
  INV_X1 U12037 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10407) );
  NOR3_X1 U12038 ( .A1(n15343), .A2(n10152), .A3(n10407), .ZN(n15342) );
  XOR2_X1 U12039 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10447), .Z(n10222) );
  NOR2_X1 U12040 ( .A1(n10223), .A2(n10222), .ZN(n10221) );
  XNOR2_X1 U12041 ( .A(n15361), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n15354) );
  NOR2_X1 U12042 ( .A1(n15355), .A2(n15354), .ZN(n15353) );
  AOI21_X1 U12043 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n15361), .A(n15353), .ZN(
        n15366) );
  XNOR2_X1 U12044 ( .A(n15372), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n15365) );
  NOR2_X1 U12045 ( .A1(n15366), .A2(n15365), .ZN(n15364) );
  INV_X1 U12046 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10153) );
  MUX2_X1 U12047 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10153), .S(n10550), .Z(
        n10154) );
  INV_X1 U12048 ( .A(n10154), .ZN(n10209) );
  NOR2_X1 U12049 ( .A1(n10210), .A2(n10209), .ZN(n10208) );
  AOI21_X1 U12050 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n10550), .A(n10208), .ZN(
        n15381) );
  XNOR2_X1 U12051 ( .A(n15384), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n15380) );
  NOR2_X1 U12052 ( .A1(n15381), .A2(n15380), .ZN(n15379) );
  XNOR2_X1 U12053 ( .A(n10727), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n10198) );
  NOR2_X1 U12054 ( .A1(n10199), .A2(n10198), .ZN(n10197) );
  INV_X1 U12055 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10155) );
  MUX2_X1 U12056 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10155), .S(n10912), .Z(
        n10156) );
  INV_X1 U12057 ( .A(n10156), .ZN(n10182) );
  INV_X1 U12058 ( .A(n10158), .ZN(n10160) );
  NAND2_X1 U12059 ( .A1(n10456), .A2(n13051), .ZN(n10176) );
  INV_X1 U12060 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n10163) );
  AND4_X1 U12061 ( .A1(n9681), .A2(n10165), .A3(n10164), .A4(n10163), .ZN(
        n10168) );
  NOR2_X1 U12062 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n10167) );
  NOR2_X1 U12063 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n10166) );
  NAND2_X1 U12064 ( .A1(n10176), .A2(n10520), .ZN(n10177) );
  AND2_X1 U12065 ( .A1(n10178), .A2(n10177), .ZN(n10190) );
  OR2_X1 U12066 ( .A1(n10179), .A2(P2_U3088), .ZN(n14484) );
  INV_X1 U12067 ( .A(n14484), .ZN(n10180) );
  INV_X1 U12068 ( .A(n10187), .ZN(n10181) );
  NOR2_X1 U12069 ( .A1(n10183), .A2(n10182), .ZN(n10325) );
  AOI211_X1 U12070 ( .C1(n10183), .C2(n10182), .A(n15406), .B(n10325), .ZN(
        n10196) );
  INV_X1 U12071 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10184) );
  XNOR2_X1 U12072 ( .A(n10398), .B(n10184), .ZN(n15346) );
  INV_X1 U12073 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n15691) );
  NOR3_X1 U12074 ( .A1(n15346), .A2(n15691), .A3(n10407), .ZN(n15345) );
  XOR2_X1 U12075 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10447), .Z(n10219) );
  NOR2_X1 U12076 ( .A1(n10220), .A2(n10219), .ZN(n10218) );
  XNOR2_X1 U12077 ( .A(n15361), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n15357) );
  NOR2_X1 U12078 ( .A1(n15358), .A2(n15357), .ZN(n15356) );
  AOI21_X1 U12079 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n15361), .A(n15356), .ZN(
        n15369) );
  XNOR2_X1 U12080 ( .A(n15372), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n15368) );
  NOR2_X1 U12081 ( .A1(n15369), .A2(n15368), .ZN(n15367) );
  INV_X1 U12082 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10185) );
  MUX2_X1 U12083 ( .A(n10185), .B(P2_REG1_REG_5__SCAN_IN), .S(n10550), .Z(
        n10212) );
  NOR2_X1 U12084 ( .A1(n10213), .A2(n10212), .ZN(n10211) );
  AOI21_X1 U12085 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n10550), .A(n10211), .ZN(
        n15378) );
  XNOR2_X1 U12086 ( .A(n15384), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n15377) );
  NOR2_X1 U12087 ( .A1(n15378), .A2(n15377), .ZN(n15376) );
  XNOR2_X1 U12088 ( .A(n10727), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n10201) );
  NOR2_X1 U12089 ( .A1(n10202), .A2(n10201), .ZN(n10200) );
  AOI21_X1 U12090 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n10727), .A(n10200), .ZN(
        n10189) );
  INV_X1 U12091 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10186) );
  MUX2_X1 U12092 ( .A(n10186), .B(P2_REG1_REG_8__SCAN_IN), .S(n10912), .Z(
        n10188) );
  INV_X1 U12093 ( .A(n15419), .ZN(n15387) );
  NOR2_X1 U12094 ( .A1(n10189), .A2(n10188), .ZN(n10318) );
  AOI211_X1 U12095 ( .C1(n10189), .C2(n10188), .A(n15387), .B(n10318), .ZN(
        n10195) );
  INV_X1 U12096 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n15460) );
  AND2_X1 U12097 ( .A1(n10179), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10191) );
  INV_X1 U12098 ( .A(n14074), .ZN(n15421) );
  NAND2_X1 U12099 ( .A1(n15421), .A2(n10912), .ZN(n10193) );
  NAND2_X1 U12100 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n10919) );
  OAI211_X1 U12101 ( .C1(n15427), .C2(n15460), .A(n10193), .B(n10919), .ZN(
        n10194) );
  OR3_X1 U12102 ( .A1(n10196), .A2(n10195), .A3(n10194), .ZN(P2_U3222) );
  AOI211_X1 U12103 ( .C1(n10199), .C2(n10198), .A(n15406), .B(n10197), .ZN(
        n10207) );
  AOI211_X1 U12104 ( .C1(n10202), .C2(n10201), .A(n15387), .B(n10200), .ZN(
        n10206) );
  NAND2_X1 U12105 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10734) );
  NAND2_X1 U12106 ( .A1(n15341), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n10203) );
  OAI211_X1 U12107 ( .C1(n14074), .C2(n10204), .A(n10734), .B(n10203), .ZN(
        n10205) );
  OR3_X1 U12108 ( .A1(n10207), .A2(n10206), .A3(n10205), .ZN(P2_U3221) );
  AOI211_X1 U12109 ( .C1(n10210), .C2(n10209), .A(n15406), .B(n10208), .ZN(
        n10217) );
  AOI211_X1 U12110 ( .C1(n10213), .C2(n10212), .A(n15387), .B(n10211), .ZN(
        n10216) );
  INV_X1 U12111 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15454) );
  NAND2_X1 U12112 ( .A1(n15421), .A2(n10550), .ZN(n10214) );
  NAND2_X1 U12113 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n13928) );
  OAI211_X1 U12114 ( .C1(n15427), .C2(n15454), .A(n10214), .B(n13928), .ZN(
        n10215) );
  OR3_X1 U12115 ( .A1(n10217), .A2(n10216), .A3(n10215), .ZN(P2_U3219) );
  AOI211_X1 U12116 ( .C1(n10220), .C2(n10219), .A(n10218), .B(n15387), .ZN(
        n10225) );
  AOI211_X1 U12117 ( .C1(n10223), .C2(n10222), .A(n10221), .B(n15406), .ZN(
        n10224) );
  NOR2_X1 U12118 ( .A1(n10225), .A2(n10224), .ZN(n10228) );
  AOI22_X1 U12119 ( .A1(n15421), .A2(n10226), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10227) );
  OAI211_X1 U12120 ( .C1(n15427), .C2(n7741), .A(n10228), .B(n10227), .ZN(
        P2_U3216) );
  INV_X1 U12121 ( .A(SI_19_), .ZN(n11728) );
  OAI222_X1 U12122 ( .A1(n13810), .A2(n11728), .B1(P3_U3151), .B2(n13407), 
        .C1(n12036), .C2(n10229), .ZN(P3_U3276) );
  NAND2_X1 U12123 ( .A1(n15419), .A2(n15691), .ZN(n10230) );
  OAI211_X1 U12124 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n15406), .A(n10230), .B(
        n14074), .ZN(n10231) );
  INV_X1 U12125 ( .A(n10231), .ZN(n10233) );
  AOI22_X1 U12126 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15423), .B1(n15419), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n10232) );
  MUX2_X1 U12127 ( .A(n10233), .B(n10232), .S(n10407), .Z(n10235) );
  AOI22_X1 U12128 ( .A1(n15341), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10234) );
  NAND2_X1 U12129 ( .A1(n10235), .A2(n10234), .ZN(P2_U3214) );
  INV_X1 U12130 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10236) );
  MUX2_X1 U12131 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10236), .S(n10636), .Z(
        n10239) );
  OAI21_X1 U12132 ( .B1(n10239), .B2(n10238), .A(n10632), .ZN(n10248) );
  INV_X1 U12133 ( .A(n10636), .ZN(n10277) );
  MUX2_X1 U12134 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n9181), .S(n10636), .Z(
        n10243) );
  AOI21_X1 U12135 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n10241), .A(n10240), 
        .ZN(n10242) );
  NAND2_X1 U12136 ( .A1(n10242), .A2(n10243), .ZN(n10635) );
  OAI21_X1 U12137 ( .B1(n10243), .B2(n10242), .A(n10635), .ZN(n10244) );
  NAND2_X1 U12138 ( .A1(n10244), .A2(n14819), .ZN(n10246) );
  AOI22_X1 U12139 ( .A1(n14791), .A2(P1_ADDR_REG_12__SCAN_IN), .B1(
        P1_REG3_REG_12__SCAN_IN), .B2(P1_U3086), .ZN(n10245) );
  OAI211_X1 U12140 ( .C1(n15432), .C2(n10277), .A(n10246), .B(n10245), .ZN(
        n10247) );
  AOI21_X1 U12141 ( .B1(n10248), .B2(n15437), .A(n10247), .ZN(n10249) );
  INV_X1 U12142 ( .A(n10249), .ZN(P1_U3255) );
  INV_X1 U12143 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10251) );
  INV_X1 U12144 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10250) );
  MUX2_X1 U12145 ( .A(n10251), .B(n10250), .S(n13408), .Z(n10253) );
  INV_X1 U12146 ( .A(n10275), .ZN(n10252) );
  NAND2_X1 U12147 ( .A1(n10253), .A2(n10252), .ZN(n10312) );
  INV_X1 U12148 ( .A(n10253), .ZN(n10254) );
  NAND2_X1 U12149 ( .A1(n10254), .A2(n10275), .ZN(n10255) );
  NAND2_X1 U12150 ( .A1(n10312), .A2(n10255), .ZN(n10257) );
  INV_X1 U12151 ( .A(n10257), .ZN(n10259) );
  OAI21_X1 U12152 ( .B1(n10259), .B2(n10258), .A(n10311), .ZN(n10273) );
  AND2_X1 U12153 ( .A1(n10263), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10260) );
  NAND2_X1 U12154 ( .A1(n10264), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10288) );
  OAI21_X1 U12155 ( .B1(n10275), .B2(n10260), .A(n10288), .ZN(n10262) );
  INV_X1 U12156 ( .A(n10289), .ZN(n10261) );
  AOI21_X1 U12157 ( .B1(n10251), .B2(n10262), .A(n10261), .ZN(n10271) );
  AOI22_X1 U12158 ( .A1(n15663), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10270) );
  NAND2_X1 U12159 ( .A1(n10264), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10294) );
  NAND2_X1 U12160 ( .A1(n10275), .A2(n10294), .ZN(n10267) );
  NAND2_X1 U12161 ( .A1(n10263), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10265) );
  OR2_X1 U12162 ( .A1(n10265), .A2(n10264), .ZN(n10266) );
  NAND2_X1 U12163 ( .A1(n10267), .A2(n10266), .ZN(n10293) );
  XNOR2_X1 U12164 ( .A(n10293), .B(P3_REG1_REG_1__SCAN_IN), .ZN(n10268) );
  NAND2_X1 U12165 ( .A1(n15667), .A2(n10268), .ZN(n10269) );
  OAI211_X1 U12166 ( .C1(n10271), .C2(n15671), .A(n10270), .B(n10269), .ZN(
        n10272) );
  AOI21_X1 U12167 ( .B1(n13412), .B2(n10273), .A(n10272), .ZN(n10274) );
  OAI21_X1 U12168 ( .B1(n10275), .B2(n15657), .A(n10274), .ZN(P3_U3183) );
  INV_X1 U12169 ( .A(n11514), .ZN(n10286) );
  OAI222_X1 U12170 ( .A1(P1_U3086), .A2(n10277), .B1(n15215), .B2(n10286), 
        .C1(n10276), .C2(n15210), .ZN(P1_U3343) );
  INV_X1 U12171 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n10280) );
  INV_X1 U12172 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n10279) );
  NAND4_X1 U12173 ( .A1(n10281), .A2(n10280), .A3(n10279), .A4(n10278), .ZN(
        n10282) );
  OAI21_X1 U12174 ( .B1(n10283), .B2(n10282), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n10284) );
  XNOR2_X1 U12175 ( .A(n10284), .B(P2_IR_REG_12__SCAN_IN), .ZN(n15422) );
  INV_X1 U12176 ( .A(n15422), .ZN(n10285) );
  OAI222_X1 U12177 ( .A1(n14503), .A2(n10287), .B1(n14506), .B2(n10286), .C1(
        n10285), .C2(P2_U3088), .ZN(P2_U3315) );
  AOI22_X1 U12178 ( .A1(n15663), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10304) );
  INV_X1 U12179 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15737) );
  OAI21_X1 U12180 ( .B1(n10291), .B2(n10290), .A(n11393), .ZN(n10292) );
  NAND2_X1 U12181 ( .A1(n13368), .A2(n10292), .ZN(n10303) );
  INV_X1 U12182 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10305) );
  NAND2_X1 U12183 ( .A1(n10293), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10295) );
  NAND2_X1 U12184 ( .A1(n10295), .A2(n10294), .ZN(n10297) );
  INV_X1 U12185 ( .A(n10296), .ZN(n10299) );
  INV_X1 U12186 ( .A(n10297), .ZN(n10298) );
  NAND2_X1 U12187 ( .A1(n10299), .A2(n10298), .ZN(n10300) );
  NAND2_X1 U12188 ( .A1(n11453), .A2(n10300), .ZN(n10301) );
  NAND2_X1 U12189 ( .A1(n15667), .A2(n10301), .ZN(n10302) );
  NAND3_X1 U12190 ( .A1(n10304), .A2(n10303), .A3(n10302), .ZN(n10316) );
  NAND2_X1 U12191 ( .A1(n10311), .A2(n10312), .ZN(n10309) );
  MUX2_X1 U12192 ( .A(n15737), .B(n10305), .S(n13408), .Z(n10306) );
  NAND2_X1 U12193 ( .A1(n10306), .A2(n11454), .ZN(n15516) );
  INV_X1 U12194 ( .A(n10306), .ZN(n10307) );
  NAND2_X1 U12195 ( .A1(n10307), .A2(n7674), .ZN(n10308) );
  AND2_X1 U12196 ( .A1(n15516), .A2(n10308), .ZN(n10310) );
  NAND2_X1 U12197 ( .A1(n10309), .A2(n10310), .ZN(n15517) );
  INV_X1 U12198 ( .A(n10310), .ZN(n10313) );
  NAND3_X1 U12199 ( .A1(n10313), .A2(n10312), .A3(n10311), .ZN(n10314) );
  AOI21_X1 U12200 ( .B1(n15517), .B2(n10314), .A(n15659), .ZN(n10315) );
  AOI211_X1 U12201 ( .C1(n15602), .C2(n11454), .A(n10316), .B(n10315), .ZN(
        n10317) );
  INV_X1 U12202 ( .A(n10317), .ZN(P3_U3184) );
  INV_X1 U12203 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10319) );
  MUX2_X1 U12204 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10319), .S(n11068), .Z(
        n10320) );
  NAND2_X1 U12205 ( .A1(n10321), .A2(n10320), .ZN(n10674) );
  OAI21_X1 U12206 ( .B1(n10321), .B2(n10320), .A(n10674), .ZN(n10324) );
  NAND2_X1 U12207 ( .A1(n15421), .A2(n11068), .ZN(n10322) );
  NAND2_X1 U12208 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n11115) );
  OAI211_X1 U12209 ( .C1(n15427), .C2(n7743), .A(n10322), .B(n11115), .ZN(
        n10323) );
  AOI21_X1 U12210 ( .B1(n10324), .B2(n15419), .A(n10323), .ZN(n10330) );
  INV_X1 U12211 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11089) );
  XNOR2_X1 U12212 ( .A(n11068), .B(n11089), .ZN(n10327) );
  AOI21_X1 U12213 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n10912), .A(n10325), .ZN(
        n10326) );
  NAND2_X1 U12214 ( .A1(n10326), .A2(n10327), .ZN(n10677) );
  OAI21_X1 U12215 ( .B1(n10327), .B2(n10326), .A(n10677), .ZN(n10328) );
  NAND2_X1 U12216 ( .A1(n10328), .A2(n15423), .ZN(n10329) );
  NAND2_X1 U12217 ( .A1(n10330), .A2(n10329), .ZN(P2_U3223) );
  OR2_X1 U12218 ( .A1(n10331), .A2(n11039), .ZN(n10332) );
  XNOR2_X1 U12219 ( .A(n10332), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11701) );
  INV_X1 U12220 ( .A(n11701), .ZN(n11368) );
  OAI222_X1 U12221 ( .A1(n14503), .A2(n10333), .B1(n14506), .B2(n11609), .C1(
        n11368), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U12222 ( .A(n10862), .ZN(n10642) );
  OAI222_X1 U12223 ( .A1(n15210), .A2(n10334), .B1(n15215), .B2(n11609), .C1(
        n10642), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U12224 ( .A(n10346), .ZN(n10338) );
  NAND3_X1 U12225 ( .A1(n10590), .A2(n10336), .A3(n10335), .ZN(n10337) );
  AOI21_X1 U12226 ( .B1(n10350), .B2(n10338), .A(n10337), .ZN(n10340) );
  NAND2_X1 U12227 ( .A1(n10353), .A2(n10345), .ZN(n10339) );
  NAND2_X1 U12228 ( .A1(n10340), .A2(n10339), .ZN(n10341) );
  NAND2_X1 U12229 ( .A1(n10341), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10344) );
  INV_X1 U12230 ( .A(n10342), .ZN(n10436) );
  NAND2_X1 U12231 ( .A1(n10355), .A2(n10436), .ZN(n10349) );
  INV_X1 U12232 ( .A(n10349), .ZN(n12752) );
  NAND2_X1 U12233 ( .A1(n10350), .A2(n12752), .ZN(n10343) );
  NOR2_X1 U12234 ( .A1(n13239), .A2(P3_U3151), .ZN(n10720) );
  INV_X1 U12235 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10359) );
  NAND2_X1 U12236 ( .A1(n10345), .A2(n15935), .ZN(n10347) );
  OAI22_X1 U12237 ( .A1(n10353), .A2(n10347), .B1(n10350), .B2(n10346), .ZN(
        n10348) );
  NAND2_X1 U12238 ( .A1(n13264), .A2(n7398), .ZN(n12617) );
  NAND2_X1 U12239 ( .A1(n11170), .A2(n12617), .ZN(n12574) );
  OR2_X1 U12240 ( .A1(n10350), .A2(n10349), .ZN(n10625) );
  INV_X1 U12241 ( .A(n10625), .ZN(n10351) );
  NAND2_X1 U12242 ( .A1(n10355), .A2(n15891), .ZN(n10352) );
  INV_X1 U12243 ( .A(n11183), .ZN(n12746) );
  OAI22_X1 U12244 ( .A1(n15720), .A2(n13225), .B1(n7398), .B2(n13242), .ZN(
        n10357) );
  AOI21_X1 U12245 ( .B1(n13221), .B2(n12574), .A(n10357), .ZN(n10358) );
  OAI21_X1 U12246 ( .B1(n10720), .B2(n10359), .A(n10358), .ZN(P3_U3172) );
  INV_X1 U12247 ( .A(P2_B_REG_SCAN_IN), .ZN(n12466) );
  XOR2_X1 U12248 ( .A(n14498), .B(n12466), .Z(n10361) );
  NAND2_X1 U12249 ( .A1(n14495), .A2(n10361), .ZN(n10362) );
  INV_X1 U12250 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15334) );
  NAND2_X1 U12251 ( .A1(n15335), .A2(n15334), .ZN(n10365) );
  INV_X1 U12252 ( .A(n14495), .ZN(n10363) );
  OR2_X1 U12253 ( .A1(n14490), .A2(n10363), .ZN(n10364) );
  NAND2_X1 U12254 ( .A1(n10365), .A2(n10364), .ZN(n10455) );
  AND2_X1 U12255 ( .A1(n15340), .A2(n10455), .ZN(n15333) );
  NOR4_X1 U12256 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n10374) );
  OR4_X1 U12257 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n10371) );
  NOR4_X1 U12258 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n10369) );
  NOR4_X1 U12259 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n10368) );
  NOR4_X1 U12260 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n10367) );
  NOR4_X1 U12261 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n10366) );
  NAND4_X1 U12262 ( .A1(n10369), .A2(n10368), .A3(n10367), .A4(n10366), .ZN(
        n10370) );
  NOR4_X1 U12263 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        n10371), .A4(n10370), .ZN(n10373) );
  NOR4_X1 U12264 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n10372) );
  NAND3_X1 U12265 ( .A1(n10374), .A2(n10373), .A3(n10372), .ZN(n10375) );
  AND2_X1 U12266 ( .A1(n10375), .A2(n15335), .ZN(n10454) );
  NAND2_X1 U12267 ( .A1(n10377), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n11282) );
  OAI21_X1 U12268 ( .B1(P2_IR_REG_18__SCAN_IN), .B2(P2_IR_REG_19__SCAN_IN), 
        .A(P2_IR_REG_31__SCAN_IN), .ZN(n10378) );
  NAND2_X1 U12269 ( .A1(n11282), .A2(n10378), .ZN(n10379) );
  NAND2_X1 U12270 ( .A1(n10382), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10383) );
  NAND2_X1 U12271 ( .A1(n10456), .A2(n13053), .ZN(n10663) );
  NAND2_X1 U12272 ( .A1(n10663), .A2(n10476), .ZN(n10384) );
  NOR2_X1 U12273 ( .A1(n10454), .A2(n10384), .ZN(n10385) );
  INV_X1 U12274 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15338) );
  INV_X1 U12275 ( .A(n14498), .ZN(n10386) );
  INV_X1 U12276 ( .A(n13119), .ZN(n10389) );
  NAND2_X1 U12277 ( .A1(n10529), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n10394) );
  NAND2_X1 U12278 ( .A1(n10528), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n10393) );
  NAND2_X1 U12279 ( .A1(n10459), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10392) );
  INV_X1 U12280 ( .A(n10460), .ZN(n10412) );
  NAND2_X1 U12281 ( .A1(n10412), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10391) );
  NAND2_X1 U12282 ( .A1(n10412), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10402) );
  NAND2_X1 U12283 ( .A1(n10459), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10401) );
  NAND2_X1 U12284 ( .A1(n10404), .A2(SI_0_), .ZN(n10406) );
  XNOR2_X1 U12285 ( .A(n10406), .B(n10405), .ZN(n14510) );
  XNOR2_X1 U12286 ( .A(n12992), .B(n10811), .ZN(n10853) );
  NAND2_X1 U12287 ( .A1(n14507), .A2(n12766), .ZN(n10409) );
  NAND2_X1 U12288 ( .A1(n10409), .A2(n14073), .ZN(n10410) );
  NAND2_X1 U12289 ( .A1(n10853), .A2(n15812), .ZN(n10423) );
  INV_X1 U12290 ( .A(n10179), .ZN(n10411) );
  NAND2_X1 U12291 ( .A1(n10412), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10416) );
  NAND2_X1 U12292 ( .A1(n10459), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10415) );
  NAND2_X1 U12293 ( .A1(n10528), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U12294 ( .A1(n14242), .A2(n12772), .B1(n14262), .B2(n14024), .ZN(
        n10422) );
  INV_X1 U12295 ( .A(n12772), .ZN(n10499) );
  NAND2_X1 U12296 ( .A1(n10499), .A2(n12771), .ZN(n10417) );
  NAND2_X1 U12297 ( .A1(n12992), .A2(n10417), .ZN(n10418) );
  NAND2_X1 U12298 ( .A1(n10829), .A2(n10418), .ZN(n10420) );
  INV_X1 U12299 ( .A(n10408), .ZN(n10473) );
  NAND2_X1 U12300 ( .A1(n10473), .A2(n13030), .ZN(n10419) );
  NAND2_X1 U12301 ( .A1(n10420), .A2(n14267), .ZN(n10421) );
  NAND3_X1 U12302 ( .A1(n10423), .A2(n10422), .A3(n10421), .ZN(n10849) );
  NAND2_X1 U12303 ( .A1(n10853), .A2(n15950), .ZN(n10424) );
  NAND2_X2 U12304 ( .A1(n8259), .A2(n10408), .ZN(n12208) );
  NAND2_X1 U12305 ( .A1(n10440), .A2(n12768), .ZN(n11102) );
  OAI211_X1 U12306 ( .C1(n10440), .C2(n12768), .A(n11286), .B(n11102), .ZN(
        n10856) );
  OAI211_X1 U12307 ( .C1(n10440), .C2(n15963), .A(n10424), .B(n10856), .ZN(
        n10425) );
  NOR2_X1 U12308 ( .A1(n10849), .A2(n10425), .ZN(n15711) );
  NAND2_X1 U12309 ( .A1(n14355), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10426) );
  OAI21_X1 U12310 ( .B1(n14355), .B2(n15711), .A(n10426), .ZN(P2_U3500) );
  AOI21_X1 U12311 ( .B1(n10428), .B2(n10427), .A(n10601), .ZN(n10435) );
  NOR2_X1 U12312 ( .A1(n10429), .A2(n10511), .ZN(n10433) );
  OAI22_X1 U12313 ( .A1(n14701), .A2(n10431), .B1(n10430), .B2(n14728), .ZN(
        n10432) );
  AOI211_X1 U12314 ( .C1(n10514), .C2(n14731), .A(n10433), .B(n10432), .ZN(
        n10434) );
  OAI21_X1 U12315 ( .B1(n10435), .B2(n14733), .A(n10434), .ZN(P1_U3237) );
  NOR2_X1 U12316 ( .A1(n10436), .A2(n15891), .ZN(n10437) );
  AOI22_X1 U12317 ( .A1(n12574), .A2(n10437), .B1(n13642), .B2(n13262), .ZN(
        n10592) );
  INV_X1 U12318 ( .A(n15940), .ZN(n15939) );
  OAI22_X1 U12319 ( .A1(n13738), .A2(n7398), .B1(n15940), .B2(n10130), .ZN(
        n10438) );
  INV_X1 U12320 ( .A(n10438), .ZN(n10439) );
  OAI21_X1 U12321 ( .B1(n10592), .B2(n15939), .A(n10439), .ZN(P3_U3459) );
  OAI21_X1 U12322 ( .B1(n10442), .B2(n10441), .A(n10443), .ZN(n10492) );
  INV_X1 U12323 ( .A(n10443), .ZN(n10444) );
  OR2_X1 U12324 ( .A1(n10520), .A2(n10447), .ZN(n10448) );
  NAND2_X1 U12325 ( .A1(n14024), .A2(n12208), .ZN(n10450) );
  AOI21_X1 U12326 ( .B1(n10453), .B2(n10452), .A(n10519), .ZN(n10481) );
  NOR2_X1 U12327 ( .A1(n10455), .A2(n10454), .ZN(n10468) );
  NAND2_X1 U12328 ( .A1(n10468), .A2(n15340), .ZN(n10666) );
  INV_X1 U12329 ( .A(n10456), .ZN(n10457) );
  NAND2_X1 U12330 ( .A1(n10457), .A2(n15963), .ZN(n10458) );
  INV_X1 U12331 ( .A(n10459), .ZN(n12066) );
  NAND2_X1 U12332 ( .A1(n12468), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10465) );
  NAND2_X1 U12333 ( .A1(n12064), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10464) );
  INV_X1 U12334 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10461) );
  NAND2_X1 U12335 ( .A1(n12425), .A2(n10461), .ZN(n10463) );
  NAND2_X1 U12336 ( .A1(n10528), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n10462) );
  NAND2_X1 U12337 ( .A1(n14262), .A2(n14023), .ZN(n10467) );
  NAND2_X1 U12338 ( .A1(n10467), .A2(n10466), .ZN(n11099) );
  INV_X1 U12339 ( .A(n10468), .ZN(n10469) );
  OAI21_X1 U12340 ( .B1(n10469), .B2(n15339), .A(n10476), .ZN(n10472) );
  AND2_X1 U12341 ( .A1(n10470), .A2(n10663), .ZN(n10471) );
  NAND2_X1 U12342 ( .A1(n10472), .A2(n10471), .ZN(n10577) );
  OR2_X1 U12343 ( .A1(n10577), .A2(P2_U3088), .ZN(n10496) );
  AOI22_X1 U12344 ( .A1(n13957), .A2(n11099), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n10496), .ZN(n10480) );
  NAND2_X1 U12345 ( .A1(n10473), .A2(n7526), .ZN(n12983) );
  INV_X1 U12346 ( .A(n12983), .ZN(n10474) );
  NAND2_X1 U12347 ( .A1(n14507), .A2(n10474), .ZN(n10852) );
  OR2_X1 U12348 ( .A1(n10475), .A2(n10852), .ZN(n10478) );
  INV_X1 U12349 ( .A(n10476), .ZN(n10477) );
  NAND2_X1 U12350 ( .A1(n14001), .A2(n12780), .ZN(n10479) );
  OAI211_X1 U12351 ( .C1(n10481), .C2(n14003), .A(n10480), .B(n10479), .ZN(
        P2_U3209) );
  INV_X1 U12352 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10482) );
  OAI22_X1 U12353 ( .A1(n13794), .A2(n7398), .B1(n15944), .B2(n10482), .ZN(
        n10483) );
  INV_X1 U12354 ( .A(n10483), .ZN(n10484) );
  OAI21_X1 U12355 ( .B1(n10592), .B2(n15941), .A(n10484), .ZN(P3_U3390) );
  NAND2_X1 U12356 ( .A1(n13263), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10485) );
  OAI21_X1 U12357 ( .B1(n12565), .B2(n13263), .A(n10485), .ZN(P3_U3521) );
  NAND2_X1 U12358 ( .A1(n13263), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10486) );
  OAI21_X1 U12359 ( .B1(n13439), .B2(n13263), .A(n10486), .ZN(P3_U3520) );
  XNOR2_X1 U12360 ( .A(n12772), .B(n12771), .ZN(n15689) );
  MUX2_X1 U12361 ( .A(n15689), .B(n12768), .S(n11286), .Z(n10489) );
  INV_X1 U12362 ( .A(n13998), .ZN(n10490) );
  NAND2_X1 U12363 ( .A1(n10496), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n10487) );
  OAI211_X1 U12364 ( .C1(n10489), .C2(n14003), .A(n10488), .B(n10487), .ZN(
        P2_U3204) );
  AOI22_X1 U12365 ( .A1(n10490), .A2(n14024), .B1(n12776), .B2(n14001), .ZN(
        n10498) );
  AOI21_X1 U12366 ( .B1(n10493), .B2(n10492), .A(n10491), .ZN(n10494) );
  NOR2_X1 U12367 ( .A1(n14003), .A2(n10494), .ZN(n10495) );
  AOI21_X1 U12368 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n10496), .A(n10495), .ZN(
        n10497) );
  OAI211_X1 U12369 ( .C1(n10499), .C2(n13997), .A(n10498), .B(n10497), .ZN(
        P2_U3194) );
  XNOR2_X1 U12370 ( .A(n10500), .B(n10501), .ZN(n15738) );
  INV_X1 U12371 ( .A(n10502), .ZN(n10506) );
  AND3_X1 U12372 ( .A1(n10700), .A2(n10504), .A3(n10503), .ZN(n10505) );
  OAI21_X1 U12373 ( .B1(n10506), .B2(n10505), .A(n15985), .ZN(n10508) );
  AOI22_X1 U12374 ( .A1(n15034), .A2(n14749), .B1(n9700), .B2(n15033), .ZN(
        n10507) );
  OAI211_X1 U12375 ( .C1(n15738), .C2(n10764), .A(n10508), .B(n10507), .ZN(
        n15741) );
  NAND2_X1 U12376 ( .A1(n15741), .A2(n15055), .ZN(n10516) );
  NAND2_X1 U12377 ( .A1(n9699), .A2(n15679), .ZN(n10509) );
  NAND2_X1 U12378 ( .A1(n10509), .A2(n10514), .ZN(n10510) );
  NAND2_X1 U12379 ( .A1(n10654), .A2(n10510), .ZN(n15740) );
  NOR2_X1 U12380 ( .A1(n15681), .A2(n15740), .ZN(n10513) );
  OAI22_X1 U12381 ( .A1(n15055), .A2(n9954), .B1(n10511), .B2(n15035), .ZN(
        n10512) );
  AOI211_X1 U12382 ( .C1(n15061), .C2(n10514), .A(n10513), .B(n10512), .ZN(
        n10515) );
  OAI211_X1 U12383 ( .C1(n15738), .C2(n11391), .A(n10516), .B(n10515), .ZN(
        P1_U3291) );
  INV_X1 U12384 ( .A(n10517), .ZN(n10518) );
  NAND2_X1 U12385 ( .A1(n10522), .A2(n12959), .ZN(n10523) );
  XNOR2_X1 U12386 ( .A(n7188), .B(n12794), .ZN(n10526) );
  NAND2_X1 U12387 ( .A1(n14023), .A2(n14208), .ZN(n10525) );
  XNOR2_X1 U12388 ( .A(n10526), .B(n10525), .ZN(n10753) );
  INV_X1 U12389 ( .A(n10525), .ZN(n10527) );
  NAND2_X1 U12390 ( .A1(n12468), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10533) );
  NAND2_X1 U12391 ( .A1(n10528), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n10532) );
  NAND2_X1 U12392 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n10543) );
  OAI21_X1 U12393 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n10543), .ZN(n10935) );
  INV_X1 U12394 ( .A(n10935), .ZN(n13959) );
  NAND2_X1 U12395 ( .A1(n10529), .A2(n13959), .ZN(n10531) );
  INV_X1 U12396 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10530) );
  INV_X2 U12397 ( .A(n11286), .ZN(n14295) );
  AND2_X1 U12398 ( .A1(n14022), .A2(n14295), .ZN(n10538) );
  NAND2_X1 U12399 ( .A1(n10534), .A2(n12959), .ZN(n10536) );
  XNOR2_X1 U12400 ( .A(n13958), .B(n7188), .ZN(n10537) );
  NOR2_X1 U12401 ( .A1(n10537), .A2(n10538), .ZN(n10539) );
  AOI21_X1 U12402 ( .B1(n10538), .B2(n10537), .A(n10539), .ZN(n13953) );
  INV_X1 U12403 ( .A(n10539), .ZN(n10540) );
  NAND2_X1 U12404 ( .A1(n12064), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10548) );
  NAND2_X1 U12405 ( .A1(n12468), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10547) );
  INV_X1 U12406 ( .A(n10543), .ZN(n10541) );
  NAND2_X1 U12407 ( .A1(n10541), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10559) );
  INV_X1 U12408 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10542) );
  NAND2_X1 U12409 ( .A1(n10543), .A2(n10542), .ZN(n10544) );
  AND2_X1 U12410 ( .A1(n10559), .A2(n10544), .ZN(n13931) );
  NAND2_X1 U12411 ( .A1(n12425), .A2(n13931), .ZN(n10546) );
  NAND2_X1 U12412 ( .A1(n10528), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n10545) );
  AND2_X1 U12413 ( .A1(n14021), .A2(n14295), .ZN(n10554) );
  AOI22_X1 U12414 ( .A1(n12336), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n12335), 
        .B2(n10550), .ZN(n10551) );
  XNOR2_X1 U12415 ( .A(n15804), .B(n7532), .ZN(n10553) );
  NOR2_X1 U12416 ( .A1(n10553), .A2(n10554), .ZN(n10555) );
  AOI21_X1 U12417 ( .B1(n10554), .B2(n10553), .A(n10555), .ZN(n13925) );
  INV_X1 U12418 ( .A(n10555), .ZN(n10556) );
  NAND2_X1 U12419 ( .A1(n12468), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10564) );
  NAND2_X1 U12420 ( .A1(n10528), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n10563) );
  INV_X1 U12421 ( .A(n10559), .ZN(n10557) );
  NAND2_X1 U12422 ( .A1(n10557), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10570) );
  INV_X1 U12423 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10558) );
  NAND2_X1 U12424 ( .A1(n10559), .A2(n10558), .ZN(n10560) );
  AND2_X1 U12425 ( .A1(n10570), .A2(n10560), .ZN(n15815) );
  NAND2_X1 U12426 ( .A1(n12425), .A2(n15815), .ZN(n10562) );
  NAND2_X1 U12427 ( .A1(n12064), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10561) );
  NAND4_X1 U12428 ( .A1(n10564), .A2(n10563), .A3(n10562), .A4(n10561), .ZN(
        n14020) );
  NAND2_X1 U12429 ( .A1(n14020), .A2(n14208), .ZN(n10722) );
  OR2_X1 U12430 ( .A1(n10565), .A2(n10521), .ZN(n10567) );
  AOI22_X1 U12431 ( .A1(n12336), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n12335), 
        .B2(n15384), .ZN(n10566) );
  XNOR2_X1 U12432 ( .A(n15819), .B(n7532), .ZN(n10721) );
  XOR2_X1 U12433 ( .A(n10722), .B(n10721), .Z(n10724) );
  XNOR2_X1 U12434 ( .A(n10725), .B(n10724), .ZN(n10580) );
  NAND2_X1 U12435 ( .A1(n12064), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10575) );
  NAND2_X1 U12436 ( .A1(n12468), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10574) );
  INV_X1 U12437 ( .A(n10570), .ZN(n10568) );
  NAND2_X1 U12438 ( .A1(n10568), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10737) );
  INV_X1 U12439 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10569) );
  NAND2_X1 U12440 ( .A1(n10570), .A2(n10569), .ZN(n10571) );
  AND2_X1 U12441 ( .A1(n10737), .A2(n10571), .ZN(n11032) );
  NAND2_X1 U12442 ( .A1(n12425), .A2(n11032), .ZN(n10573) );
  NAND2_X1 U12443 ( .A1(n7508), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n10572) );
  NAND4_X1 U12444 ( .A1(n10575), .A2(n10574), .A3(n10573), .A4(n10572), .ZN(
        n14019) );
  AOI22_X1 U12445 ( .A1(n14242), .A2(n14021), .B1(n14262), .B2(n14019), .ZN(
        n10836) );
  INV_X1 U12446 ( .A(n10836), .ZN(n10576) );
  AOI22_X1 U12447 ( .A1(n13957), .A2(n10576), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10579) );
  INV_X1 U12448 ( .A(n13995), .ZN(n13971) );
  AOI22_X1 U12449 ( .A1(n13971), .A2(n15815), .B1(n14001), .B2(n15819), .ZN(
        n10578) );
  OAI211_X1 U12450 ( .C1(n10580), .C2(n14003), .A(n10579), .B(n10578), .ZN(
        P2_U3211) );
  NAND2_X1 U12451 ( .A1(n13263), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n10581) );
  OAI21_X1 U12452 ( .B1(n13456), .B2(n13263), .A(n10581), .ZN(P3_U3519) );
  INV_X1 U12453 ( .A(n11980), .ZN(n10585) );
  INV_X1 U12454 ( .A(n11595), .ZN(n11587) );
  OAI222_X1 U12455 ( .A1(n15210), .A2(n10582), .B1(n15215), .B2(n10585), .C1(
        P1_U3086), .C2(n11587), .ZN(P1_U3341) );
  INV_X1 U12456 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n10583) );
  NAND2_X1 U12457 ( .A1(n10331), .A2(n10583), .ZN(n10781) );
  NAND2_X1 U12458 ( .A1(n10781), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10584) );
  XNOR2_X1 U12459 ( .A(n10584), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14027) );
  INV_X1 U12460 ( .A(n14027), .ZN(n14037) );
  OAI222_X1 U12461 ( .A1(n14509), .A2(n10586), .B1(n14506), .B2(n10585), .C1(
        P2_U3088), .C2(n14037), .ZN(P2_U3313) );
  XNOR2_X1 U12462 ( .A(n10588), .B(n10587), .ZN(n10589) );
  NAND3_X1 U12463 ( .A1(n10591), .A2(n10590), .A3(n10589), .ZN(n10594) );
  MUX2_X1 U12464 ( .A(n10593), .B(n10592), .S(n15735), .Z(n10598) );
  INV_X1 U12465 ( .A(n10594), .ZN(n10595) );
  NOR2_X1 U12466 ( .A1(n15935), .A2(n11183), .ZN(n15695) );
  INV_X1 U12467 ( .A(n13650), .ZN(n13663) );
  AOI22_X1 U12468 ( .A1(n13663), .A2(n10596), .B1(n13648), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10597) );
  NAND2_X1 U12469 ( .A1(n10598), .A2(n10597), .ZN(P3_U3233) );
  OAI21_X1 U12470 ( .B1(n10601), .B2(n10600), .A(n10599), .ZN(n10602) );
  NAND3_X1 U12471 ( .A1(n10603), .A2(n16036), .A3(n10602), .ZN(n10611) );
  INV_X1 U12472 ( .A(n14731), .ZN(n16033) );
  NAND2_X1 U12473 ( .A1(n16029), .A2(n10604), .ZN(n10605) );
  OAI21_X1 U12474 ( .B1(n16033), .B2(n15756), .A(n10605), .ZN(n10609) );
  INV_X1 U12475 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10606) );
  OAI22_X1 U12476 ( .A1(n14728), .A2(n10607), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10606), .ZN(n10608) );
  NOR2_X1 U12477 ( .A1(n10609), .A2(n10608), .ZN(n10610) );
  OAI211_X1 U12478 ( .C1(n16041), .C2(P1_REG3_REG_3__SCAN_IN), .A(n10611), .B(
        n10610), .ZN(P1_U3218) );
  INV_X1 U12479 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15696) );
  INV_X1 U12480 ( .A(n10616), .ZN(n10618) );
  AND2_X4 U12481 ( .A1(n10618), .A2(n10617), .ZN(n13106) );
  INV_X4 U12482 ( .A(n13106), .ZN(n13109) );
  INV_X1 U12483 ( .A(n11171), .ZN(n10619) );
  XNOR2_X1 U12484 ( .A(n10620), .B(n13106), .ZN(n10621) );
  NOR2_X1 U12485 ( .A1(n13262), .A2(n10621), .ZN(n10708) );
  NAND2_X1 U12486 ( .A1(n10623), .A2(n13221), .ZN(n10628) );
  OAI22_X1 U12487 ( .A1(n11172), .A2(n13225), .B1(n15697), .B2(n13242), .ZN(
        n10626) );
  AOI21_X1 U12488 ( .B1(n13223), .B2(n13264), .A(n10626), .ZN(n10627) );
  OAI211_X1 U12489 ( .C1(n10720), .C2(n15696), .A(n10628), .B(n10627), .ZN(
        P3_U3162) );
  INV_X1 U12490 ( .A(n10629), .ZN(n10630) );
  INV_X1 U12491 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10631) );
  MUX2_X1 U12492 ( .A(n10631), .B(P1_REG1_REG_13__SCAN_IN), .S(n10862), .Z(
        n10634) );
  OAI21_X1 U12493 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n10636), .A(n10632), 
        .ZN(n10633) );
  NOR2_X1 U12494 ( .A1(n10633), .A2(n10634), .ZN(n10861) );
  AOI211_X1 U12495 ( .C1(n10634), .C2(n10633), .A(n14823), .B(n10861), .ZN(
        n10645) );
  OAI21_X1 U12496 ( .B1(n10636), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10635), 
        .ZN(n10639) );
  MUX2_X1 U12497 ( .A(n9218), .B(P1_REG2_REG_13__SCAN_IN), .S(n10862), .Z(
        n10638) );
  OR2_X1 U12498 ( .A1(n10639), .A2(n10638), .ZN(n10859) );
  INV_X1 U12499 ( .A(n10859), .ZN(n10637) );
  AOI211_X1 U12500 ( .C1(n10639), .C2(n10638), .A(n15434), .B(n10637), .ZN(
        n10644) );
  NOR2_X1 U12501 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n12273), .ZN(n10640) );
  AOI21_X1 U12502 ( .B1(n14791), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10640), 
        .ZN(n10641) );
  OAI21_X1 U12503 ( .B1(n15432), .B2(n10642), .A(n10641), .ZN(n10643) );
  OR3_X1 U12504 ( .A1(n10645), .A2(n10644), .A3(n10643), .ZN(P1_U3256) );
  XNOR2_X1 U12505 ( .A(n10647), .B(n10646), .ZN(n10648) );
  NAND2_X1 U12506 ( .A1(n10648), .A2(n15985), .ZN(n10650) );
  AOI22_X1 U12507 ( .A1(n10604), .A2(n15033), .B1(n15034), .B2(n14748), .ZN(
        n10649) );
  NAND2_X1 U12508 ( .A1(n10650), .A2(n10649), .ZN(n15758) );
  INV_X1 U12509 ( .A(n15758), .ZN(n10662) );
  XNOR2_X1 U12510 ( .A(n10651), .B(n10652), .ZN(n15760) );
  OR2_X1 U12511 ( .A1(n15036), .A2(n10764), .ZN(n10653) );
  NAND2_X1 U12512 ( .A1(n11391), .A2(n10653), .ZN(n15025) );
  INV_X1 U12513 ( .A(n10654), .ZN(n10656) );
  INV_X1 U12514 ( .A(n10689), .ZN(n10655) );
  OAI21_X1 U12515 ( .B1(n15756), .B2(n10656), .A(n10655), .ZN(n15757) );
  OAI22_X1 U12516 ( .A1(n15055), .A2(n9955), .B1(n15035), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n10657) );
  AOI21_X1 U12517 ( .B1(n15061), .B2(n10658), .A(n10657), .ZN(n10659) );
  OAI21_X1 U12518 ( .B1(n15681), .B2(n15757), .A(n10659), .ZN(n10660) );
  AOI21_X1 U12519 ( .B1(n15760), .B2(n15025), .A(n10660), .ZN(n10661) );
  OAI21_X1 U12520 ( .B1(n10662), .B2(n15020), .A(n10661), .ZN(P1_U3290) );
  INV_X1 U12521 ( .A(n10663), .ZN(n10664) );
  OR3_X1 U12522 ( .A1(n10666), .A2(n10665), .A3(n10664), .ZN(n10667) );
  NAND2_X1 U12523 ( .A1(n8259), .A2(n12771), .ZN(n15688) );
  INV_X1 U12524 ( .A(n14267), .ZN(n14289) );
  AOI21_X1 U12525 ( .B1(n14289), .B2(n15778), .A(n15689), .ZN(n10668) );
  OAI21_X1 U12526 ( .B1(n12963), .B2(n15688), .A(n7201), .ZN(n10669) );
  AOI21_X1 U12527 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n15816), .A(n10669), .ZN(
        n10670) );
  NOR2_X1 U12528 ( .A1(n10670), .A2(n15817), .ZN(n10671) );
  AOI21_X1 U12529 ( .B1(n15817), .B2(P2_REG2_REG_0__SCAN_IN), .A(n10671), .ZN(
        n10672) );
  OAI21_X1 U12530 ( .B1(n15689), .B2(n14129), .A(n10672), .ZN(P2_U3265) );
  INV_X1 U12531 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10673) );
  MUX2_X1 U12532 ( .A(n10673), .B(P2_REG1_REG_10__SCAN_IN), .S(n11124), .Z(
        n10676) );
  OAI21_X1 U12533 ( .B1(n11068), .B2(P2_REG1_REG_9__SCAN_IN), .A(n10674), .ZN(
        n10675) );
  NOR2_X1 U12534 ( .A1(n10675), .A2(n10676), .ZN(n10903) );
  AOI211_X1 U12535 ( .C1(n10676), .C2(n10675), .A(n15387), .B(n10903), .ZN(
        n10683) );
  XNOR2_X1 U12536 ( .A(n11124), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n10679) );
  OAI21_X1 U12537 ( .B1(n11068), .B2(P2_REG2_REG_9__SCAN_IN), .A(n10677), .ZN(
        n10678) );
  NOR2_X1 U12538 ( .A1(n10678), .A2(n10679), .ZN(n10896) );
  AOI211_X1 U12539 ( .C1(n10679), .C2(n10678), .A(n15406), .B(n10896), .ZN(
        n10682) );
  INV_X1 U12540 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15470) );
  NAND2_X1 U12541 ( .A1(n15421), .A2(n11124), .ZN(n10680) );
  NAND2_X1 U12542 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11291)
         );
  OAI211_X1 U12543 ( .C1(n15427), .C2(n15470), .A(n10680), .B(n11291), .ZN(
        n10681) );
  OR3_X1 U12544 ( .A1(n10683), .A2(n10682), .A3(n10681), .ZN(P2_U3224) );
  XOR2_X1 U12545 ( .A(n10687), .B(n10684), .Z(n10768) );
  XOR2_X1 U12546 ( .A(n10687), .B(n10686), .Z(n10688) );
  AOI222_X1 U12547 ( .A1(n10688), .A2(n15985), .B1(n14747), .B2(n15034), .C1(
        n14749), .C2(n15033), .ZN(n10767) );
  OR2_X1 U12548 ( .A1(n10767), .A2(n15036), .ZN(n10695) );
  OR2_X1 U12549 ( .A1(n10689), .A2(n10691), .ZN(n10690) );
  AND2_X1 U12550 ( .A1(n10793), .A2(n10690), .ZN(n10765) );
  NOR2_X1 U12551 ( .A1(n15680), .A2(n10691), .ZN(n10693) );
  OAI22_X1 U12552 ( .A1(n15055), .A2(n9958), .B1(n10949), .B2(n15035), .ZN(
        n10692) );
  AOI211_X1 U12553 ( .C1(n10765), .C2(n15018), .A(n10693), .B(n10692), .ZN(
        n10694) );
  OAI211_X1 U12554 ( .C1(n10768), .C2(n14988), .A(n10695), .B(n10694), .ZN(
        P1_U3289) );
  INV_X1 U12555 ( .A(n11391), .ZN(n15684) );
  XNOR2_X1 U12556 ( .A(n9812), .B(n10696), .ZN(n15707) );
  XNOR2_X1 U12557 ( .A(n9699), .B(n15679), .ZN(n15704) );
  INV_X1 U12558 ( .A(n15035), .ZN(n15678) );
  AOI22_X1 U12559 ( .A1(n15061), .A2(n10697), .B1(n15678), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n10698) );
  OAI21_X1 U12560 ( .B1(n15704), .B2(n15681), .A(n10698), .ZN(n10706) );
  INV_X1 U12561 ( .A(n10764), .ZN(n11648) );
  NAND2_X1 U12562 ( .A1(n15707), .A2(n11648), .ZN(n10704) );
  AOI22_X1 U12563 ( .A1(n10604), .A2(n15034), .B1(n15033), .B2(n14750), .ZN(
        n10703) );
  NAND2_X1 U12564 ( .A1(n10700), .A2(n10699), .ZN(n10701) );
  NAND2_X1 U12565 ( .A1(n10701), .A2(n15985), .ZN(n10702) );
  NAND3_X1 U12566 ( .A1(n10704), .A2(n10703), .A3(n10702), .ZN(n15705) );
  MUX2_X1 U12567 ( .A(n15705), .B(P1_REG2_REG_1__SCAN_IN), .S(n15036), .Z(
        n10705) );
  AOI211_X1 U12568 ( .C1(n15684), .C2(n15707), .A(n10706), .B(n10705), .ZN(
        n10707) );
  INV_X1 U12569 ( .A(n10707), .ZN(P1_U3292) );
  INV_X1 U12570 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15728) );
  XNOR2_X1 U12571 ( .A(n10714), .B(n7218), .ZN(n10773) );
  XNOR2_X1 U12572 ( .A(n13261), .B(n10773), .ZN(n10712) );
  INV_X1 U12573 ( .A(n10708), .ZN(n10709) );
  NAND2_X1 U12574 ( .A1(n10710), .A2(n10709), .ZN(n10711) );
  OAI21_X1 U12575 ( .B1(n10712), .B2(n10711), .A(n10775), .ZN(n10713) );
  NAND2_X1 U12576 ( .A1(n10713), .A2(n13221), .ZN(n10719) );
  OR2_X1 U12577 ( .A1(n15720), .A2(n13237), .ZN(n10716) );
  NAND2_X1 U12578 ( .A1(n13206), .A2(n10714), .ZN(n10715) );
  OAI211_X1 U12579 ( .C1(n15722), .C2(n13225), .A(n10716), .B(n10715), .ZN(
        n10717) );
  INV_X1 U12580 ( .A(n10717), .ZN(n10718) );
  OAI211_X1 U12581 ( .C1(n10720), .C2(n15728), .A(n10719), .B(n10718), .ZN(
        P3_U3177) );
  INV_X1 U12582 ( .A(n10721), .ZN(n10723) );
  NAND2_X1 U12583 ( .A1(n10726), .A2(n12959), .ZN(n10729) );
  AOI22_X1 U12584 ( .A1(n12336), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n12335), 
        .B2(n10727), .ZN(n10728) );
  XNOR2_X1 U12585 ( .A(n15844), .B(n13847), .ZN(n10731) );
  NAND2_X1 U12586 ( .A1(n14019), .A2(n14208), .ZN(n10730) );
  AOI21_X1 U12587 ( .B1(n10733), .B2(n10732), .A(n7354), .ZN(n10747) );
  INV_X1 U12588 ( .A(n10734), .ZN(n10744) );
  NAND2_X1 U12589 ( .A1(n12064), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10742) );
  NAND2_X1 U12590 ( .A1(n12468), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10741) );
  INV_X1 U12591 ( .A(n10737), .ZN(n10735) );
  NAND2_X1 U12592 ( .A1(n10735), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10922) );
  INV_X1 U12593 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10736) );
  NAND2_X1 U12594 ( .A1(n10737), .A2(n10736), .ZN(n10738) );
  AND2_X1 U12595 ( .A1(n10922), .A2(n10738), .ZN(n11020) );
  NAND2_X1 U12596 ( .A1(n12425), .A2(n11020), .ZN(n10740) );
  NAND2_X1 U12597 ( .A1(n7508), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n10739) );
  NAND4_X1 U12598 ( .A1(n10742), .A2(n10741), .A3(n10740), .A4(n10739), .ZN(
        n14018) );
  AOI22_X1 U12599 ( .A1(n14242), .A2(n14020), .B1(n14262), .B2(n14018), .ZN(
        n11028) );
  NOR2_X1 U12600 ( .A1(n13939), .A2(n11028), .ZN(n10743) );
  AOI211_X1 U12601 ( .C1(n13971), .C2(n11032), .A(n10744), .B(n10743), .ZN(
        n10746) );
  NAND2_X1 U12602 ( .A1(n14001), .A2(n15844), .ZN(n10745) );
  OAI211_X1 U12603 ( .C1(n10747), .C2(n14003), .A(n10746), .B(n10745), .ZN(
        P2_U3185) );
  INV_X1 U12604 ( .A(n10748), .ZN(n10750) );
  OAI222_X1 U12605 ( .A1(P3_U3151), .A2(n10751), .B1(n12036), .B2(n10750), 
        .C1(n10749), .C2(n13810), .ZN(P3_U3274) );
  XNOR2_X1 U12606 ( .A(n10752), .B(n10753), .ZN(n10758) );
  INV_X1 U12607 ( .A(n13997), .ZN(n10756) );
  OAI22_X1 U12608 ( .A1(n13995), .A2(P2_REG3_REG_3__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n10461), .ZN(n10755) );
  INV_X1 U12609 ( .A(n14022), .ZN(n10954) );
  OAI22_X1 U12610 ( .A1(n13998), .A2(n10954), .B1(n13974), .B2(n15764), .ZN(
        n10754) );
  AOI211_X1 U12611 ( .C1(n10756), .C2(n14024), .A(n10755), .B(n10754), .ZN(
        n10757) );
  OAI21_X1 U12612 ( .B1(n10758), .B2(n14003), .A(n10757), .ZN(P2_U3190) );
  INV_X1 U12613 ( .A(n10759), .ZN(n10761) );
  OAI22_X1 U12614 ( .A1(n12754), .A2(P3_U3151), .B1(SI_22_), .B2(n13810), .ZN(
        n10760) );
  AOI21_X1 U12615 ( .B1(n10761), .B2(n13798), .A(n10760), .ZN(P3_U3273) );
  AOI22_X1 U12616 ( .A1(n10765), .A2(n15796), .B1(n16014), .B2(n10946), .ZN(
        n10766) );
  OAI211_X1 U12617 ( .C1(n15799), .C2(n10768), .A(n10767), .B(n10766), .ZN(
        n10770) );
  NAND2_X1 U12618 ( .A1(n10770), .A2(n15961), .ZN(n10769) );
  OAI21_X1 U12619 ( .B1(n15961), .B2(n8995), .A(n10769), .ZN(P1_U3471) );
  INV_X2 U12620 ( .A(n16021), .ZN(n15922) );
  NAND2_X1 U12621 ( .A1(n10770), .A2(n15922), .ZN(n10771) );
  OAI21_X1 U12622 ( .B1(n15922), .B2(n10772), .A(n10771), .ZN(P1_U3532) );
  INV_X1 U12623 ( .A(n13239), .ZN(n12169) );
  NAND2_X1 U12624 ( .A1(n10773), .A2(n11172), .ZN(n10774) );
  AND2_X1 U12625 ( .A1(n10775), .A2(n10774), .ZN(n10777) );
  XNOR2_X1 U12626 ( .A(n7543), .B(n11186), .ZN(n10871) );
  XNOR2_X1 U12627 ( .A(n10871), .B(n15722), .ZN(n10776) );
  OAI211_X1 U12628 ( .C1(n10777), .C2(n10776), .A(n13221), .B(n10872), .ZN(
        n10780) );
  NOR2_X1 U12629 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11880), .ZN(n15512) );
  OAI22_X1 U12630 ( .A1(n11172), .A2(n13237), .B1(n11238), .B2(n13225), .ZN(
        n10778) );
  AOI211_X1 U12631 ( .C1(n11186), .C2(n13206), .A(n15512), .B(n10778), .ZN(
        n10779) );
  OAI211_X1 U12632 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12169), .A(n10780), .B(
        n10779), .ZN(P3_U3158) );
  INV_X1 U12633 ( .A(n12055), .ZN(n10784) );
  NAND2_X1 U12634 ( .A1(n11925), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10782) );
  XNOR2_X1 U12635 ( .A(n10782), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15393) );
  INV_X1 U12636 ( .A(n15393), .ZN(n14040) );
  OAI222_X1 U12637 ( .A1(n14509), .A2(n10783), .B1(n14506), .B2(n10784), .C1(
        n14040), .C2(P2_U3088), .ZN(P2_U3312) );
  OAI222_X1 U12638 ( .A1(n15210), .A2(n10785), .B1(n15215), .B2(n10784), .C1(
        n15433), .C2(P1_U3086), .ZN(P1_U3340) );
  XNOR2_X1 U12639 ( .A(n10786), .B(n10787), .ZN(n15800) );
  XNOR2_X1 U12640 ( .A(n10788), .B(n10787), .ZN(n10789) );
  NAND2_X1 U12641 ( .A1(n10789), .A2(n15985), .ZN(n10791) );
  AOI22_X1 U12642 ( .A1(n15033), .A2(n14748), .B1(n14746), .B2(n15034), .ZN(
        n10790) );
  NAND2_X1 U12643 ( .A1(n10791), .A2(n10790), .ZN(n15802) );
  MUX2_X1 U12644 ( .A(n15802), .B(P1_REG2_REG_5__SCAN_IN), .S(n15036), .Z(
        n10792) );
  INV_X1 U12645 ( .A(n10792), .ZN(n10798) );
  NAND2_X1 U12646 ( .A1(n10793), .A2(n15795), .ZN(n10794) );
  AND2_X1 U12647 ( .A1(n10978), .A2(n10794), .ZN(n15797) );
  OAI22_X1 U12648 ( .A1(n15680), .A2(n10795), .B1(n15035), .B2(n10803), .ZN(
        n10796) );
  AOI21_X1 U12649 ( .B1(n15797), .B2(n15018), .A(n10796), .ZN(n10797) );
  OAI211_X1 U12650 ( .C1(n15800), .C2(n14988), .A(n10798), .B(n10797), .ZN(
        P1_U3288) );
  NOR2_X1 U12651 ( .A1(n10800), .A2(n8090), .ZN(n10801) );
  XNOR2_X1 U12652 ( .A(n10802), .B(n10801), .ZN(n10810) );
  AOI22_X1 U12653 ( .A1(n16029), .A2(n14748), .B1(n15795), .B2(n14731), .ZN(
        n10809) );
  INV_X1 U12654 ( .A(n14746), .ZN(n10806) );
  OR2_X1 U12655 ( .A1(n16041), .A2(n10803), .ZN(n10804) );
  OAI211_X1 U12656 ( .C1(n14728), .C2(n10806), .A(n10805), .B(n10804), .ZN(
        n10807) );
  INV_X1 U12657 ( .A(n10807), .ZN(n10808) );
  OAI211_X1 U12658 ( .C1(n10810), .C2(n14733), .A(n10809), .B(n10808), .ZN(
        P1_U3227) );
  XNOR2_X1 U12659 ( .A(n15819), .B(n14020), .ZN(n12999) );
  NAND2_X1 U12660 ( .A1(n12992), .A2(n10811), .ZN(n10814) );
  NAND2_X1 U12661 ( .A1(n10812), .A2(n10440), .ZN(n10813) );
  NAND2_X1 U12662 ( .A1(n10814), .A2(n10813), .ZN(n11096) );
  INV_X1 U12663 ( .A(n14024), .ZN(n10955) );
  NAND2_X1 U12664 ( .A1(n10955), .A2(n12780), .ZN(n10957) );
  NAND2_X1 U12665 ( .A1(n14024), .A2(n15749), .ZN(n10815) );
  INV_X1 U12666 ( .A(n12994), .ZN(n10816) );
  NAND2_X1 U12667 ( .A1(n11096), .A2(n10816), .ZN(n10818) );
  NAND2_X1 U12668 ( .A1(n10955), .A2(n15749), .ZN(n10817) );
  INV_X1 U12669 ( .A(n14023), .ZN(n10933) );
  NAND2_X1 U12670 ( .A1(n10933), .A2(n12794), .ZN(n10831) );
  NAND2_X1 U12671 ( .A1(n14023), .A2(n15764), .ZN(n10819) );
  AND2_X1 U12672 ( .A1(n10831), .A2(n10819), .ZN(n12993) );
  NAND2_X1 U12673 ( .A1(n10933), .A2(n15764), .ZN(n10820) );
  XNOR2_X1 U12674 ( .A(n15782), .B(n14022), .ZN(n12996) );
  NAND2_X1 U12675 ( .A1(n15782), .A2(n10954), .ZN(n10821) );
  NAND2_X1 U12676 ( .A1(n10822), .A2(n10821), .ZN(n10887) );
  NOR2_X1 U12677 ( .A1(n15804), .A2(n14021), .ZN(n10823) );
  NAND2_X1 U12678 ( .A1(n15804), .A2(n14021), .ZN(n10824) );
  INV_X1 U12679 ( .A(n11017), .ZN(n10826) );
  AOI21_X1 U12680 ( .B1(n12999), .B2(n10827), .A(n10826), .ZN(n15820) );
  INV_X1 U12681 ( .A(n15950), .ZN(n15807) );
  INV_X1 U12682 ( .A(n12996), .ZN(n10939) );
  NAND2_X1 U12683 ( .A1(n10954), .A2(n13958), .ZN(n10832) );
  INV_X1 U12684 ( .A(n15804), .ZN(n10833) );
  NAND2_X1 U12685 ( .A1(n10833), .A2(n14021), .ZN(n10834) );
  INV_X1 U12686 ( .A(n14021), .ZN(n12807) );
  NAND2_X1 U12687 ( .A1(n15804), .A2(n12807), .ZN(n10835) );
  XNOR2_X1 U12688 ( .A(n11005), .B(n12999), .ZN(n10838) );
  OAI21_X1 U12689 ( .B1(n15820), .B2(n15778), .A(n10836), .ZN(n10837) );
  AOI21_X1 U12690 ( .B1(n14309), .B2(n10838), .A(n10837), .ZN(n15828) );
  INV_X1 U12691 ( .A(n15819), .ZN(n10842) );
  OR2_X1 U12692 ( .A1(n11102), .A2(n12780), .ZN(n11103) );
  NAND2_X1 U12693 ( .A1(n10961), .A2(n15782), .ZN(n10936) );
  OR2_X1 U12694 ( .A1(n10936), .A2(n15804), .ZN(n10888) );
  INV_X1 U12695 ( .A(n10888), .ZN(n10839) );
  NOR2_X1 U12696 ( .A1(n10888), .A2(n15819), .ZN(n11015) );
  INV_X1 U12697 ( .A(n11015), .ZN(n11031) );
  OAI211_X1 U12698 ( .C1(n10842), .C2(n10839), .A(n11031), .B(n11286), .ZN(
        n15821) );
  OAI211_X1 U12699 ( .C1(n15820), .C2(n15807), .A(n15828), .B(n15821), .ZN(
        n10845) );
  NAND2_X1 U12700 ( .A1(n15974), .A2(n15845), .ZN(n14467) );
  INV_X1 U12701 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10841) );
  OAI22_X1 U12702 ( .A1(n14467), .A2(n10842), .B1(n15974), .B2(n10841), .ZN(
        n10843) );
  AOI21_X1 U12703 ( .B1(n10845), .B2(n15974), .A(n10843), .ZN(n10844) );
  INV_X1 U12704 ( .A(n10844), .ZN(P2_U3448) );
  INV_X1 U12705 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10848) );
  NAND2_X1 U12706 ( .A1(n10845), .A2(n15970), .ZN(n10847) );
  NAND2_X1 U12707 ( .A1(n14422), .A2(n15819), .ZN(n10846) );
  OAI211_X1 U12708 ( .C1(n15970), .C2(n10848), .A(n10847), .B(n10846), .ZN(
        P2_U3505) );
  AOI22_X1 U12709 ( .A1(n14275), .A2(n10849), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n15816), .ZN(n10850) );
  INV_X1 U12710 ( .A(n10850), .ZN(n10851) );
  AOI21_X1 U12711 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n15817), .A(n10851), .ZN(
        n10855) );
  INV_X1 U12712 ( .A(n14129), .ZN(n15824) );
  NOR2_X2 U12713 ( .A1(n15817), .A2(n10852), .ZN(n15818) );
  AOI22_X1 U12714 ( .A1(n15824), .A2(n10853), .B1(n15818), .B2(n12776), .ZN(
        n10854) );
  OAI211_X1 U12715 ( .C1(n14234), .C2(n10856), .A(n10855), .B(n10854), .ZN(
        P2_U3264) );
  NAND2_X1 U12716 ( .A1(n10862), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10858) );
  MUX2_X1 U12717 ( .A(n9231), .B(P1_REG2_REG_14__SCAN_IN), .S(n11595), .Z(
        n10857) );
  AOI21_X1 U12718 ( .B1(n10859), .B2(n10858), .A(n10857), .ZN(n11594) );
  NAND3_X1 U12719 ( .A1(n10859), .A2(n10858), .A3(n10857), .ZN(n10860) );
  NAND2_X1 U12720 ( .A1(n10860), .A2(n14819), .ZN(n10870) );
  AOI21_X1 U12721 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n10862), .A(n10861), 
        .ZN(n11588) );
  XNOR2_X1 U12722 ( .A(n11588), .B(n11587), .ZN(n10864) );
  INV_X1 U12723 ( .A(n10864), .ZN(n10865) );
  INV_X1 U12724 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10863) );
  OAI211_X1 U12725 ( .C1(n10865), .C2(P1_REG1_REG_14__SCAN_IN), .A(n11586), 
        .B(n15437), .ZN(n10869) );
  NAND2_X1 U12726 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14633)
         );
  INV_X1 U12727 ( .A(n14633), .ZN(n10867) );
  NOR2_X1 U12728 ( .A1(n15432), .A2(n11587), .ZN(n10866) );
  AOI211_X1 U12729 ( .C1(n14791), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n10867), 
        .B(n10866), .ZN(n10868) );
  OAI211_X1 U12730 ( .C1(n11594), .C2(n10870), .A(n10869), .B(n10868), .ZN(
        P1_U3257) );
  INV_X1 U12731 ( .A(n10871), .ZN(n10873) );
  XNOR2_X1 U12732 ( .A(n15772), .B(n13109), .ZN(n10874) );
  AOI21_X1 U12733 ( .B1(n10876), .B2(n10875), .A(n11047), .ZN(n10881) );
  INV_X1 U12734 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10877) );
  NOR2_X1 U12735 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10877), .ZN(n15530) );
  OAI22_X1 U12736 ( .A1(n15722), .A2(n13237), .B1(n11226), .B2(n13225), .ZN(
        n10878) );
  AOI211_X1 U12737 ( .C1(n15772), .C2(n13206), .A(n15530), .B(n10878), .ZN(
        n10880) );
  NAND2_X1 U12738 ( .A1(n13239), .A2(n11197), .ZN(n10879) );
  OAI211_X1 U12739 ( .C1(n10881), .C2(n13229), .A(n10880), .B(n10879), .ZN(
        P3_U3170) );
  NAND2_X1 U12740 ( .A1(n10882), .A2(n13798), .ZN(n10883) );
  OAI211_X1 U12741 ( .C1(n11723), .C2(n13810), .A(n10883), .B(n12756), .ZN(
        P3_U3272) );
  XNOR2_X1 U12742 ( .A(n15804), .B(n14021), .ZN(n12998) );
  XOR2_X1 U12743 ( .A(n10884), .B(n12998), .Z(n10885) );
  AOI22_X1 U12744 ( .A1(n14242), .A2(n14022), .B1(n14262), .B2(n14020), .ZN(
        n13927) );
  OAI21_X1 U12745 ( .B1(n10885), .B2(n14289), .A(n13927), .ZN(n15809) );
  MUX2_X1 U12746 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n15809), .S(n14275), .Z(
        n10893) );
  NAND2_X1 U12747 ( .A1(n14275), .A2(n15812), .ZN(n10886) );
  XNOR2_X1 U12748 ( .A(n10887), .B(n12998), .ZN(n15808) );
  AOI22_X1 U12749 ( .A1(n15818), .A2(n15804), .B1(n15816), .B2(n13931), .ZN(
        n10891) );
  AOI21_X1 U12750 ( .B1(n10936), .B2(n15804), .A(n14295), .ZN(n10889) );
  NAND2_X1 U12751 ( .A1(n10889), .A2(n10888), .ZN(n15806) );
  OR2_X1 U12752 ( .A1(n14234), .A2(n15806), .ZN(n10890) );
  OAI211_X1 U12753 ( .C1(n14254), .C2(n15808), .A(n10891), .B(n10890), .ZN(
        n10892) );
  OR2_X1 U12754 ( .A1(n10893), .A2(n10892), .ZN(P2_U3260) );
  INV_X1 U12755 ( .A(n12170), .ZN(n10894) );
  INV_X1 U12756 ( .A(n12112), .ZN(n11603) );
  OAI222_X1 U12757 ( .A1(n15210), .A2(n10895), .B1(n15215), .B2(n10894), .C1(
        n11603), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U12758 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10897) );
  MUX2_X1 U12759 ( .A(n10897), .B(P2_REG2_REG_11__SCAN_IN), .S(n11361), .Z(
        n10898) );
  INV_X1 U12760 ( .A(n10898), .ZN(n10899) );
  NAND2_X1 U12761 ( .A1(n10900), .A2(n10899), .ZN(n11360) );
  OAI21_X1 U12762 ( .B1(n10900), .B2(n10899), .A(n11360), .ZN(n10909) );
  INV_X1 U12763 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n15475) );
  NAND2_X1 U12764 ( .A1(n15421), .A2(n11361), .ZN(n10902) );
  NAND2_X1 U12765 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n10901)
         );
  OAI211_X1 U12766 ( .C1(n15427), .C2(n15475), .A(n10902), .B(n10901), .ZN(
        n10908) );
  INV_X1 U12767 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10904) );
  MUX2_X1 U12768 ( .A(n10904), .B(P2_REG1_REG_11__SCAN_IN), .S(n11361), .Z(
        n10905) );
  NOR2_X1 U12769 ( .A1(n10906), .A2(n10905), .ZN(n11355) );
  AOI211_X1 U12770 ( .C1(n10906), .C2(n10905), .A(n15387), .B(n11355), .ZN(
        n10907) );
  AOI211_X1 U12771 ( .C1(n15423), .C2(n10909), .A(n10908), .B(n10907), .ZN(
        n10910) );
  INV_X1 U12772 ( .A(n10910), .ZN(P2_U3225) );
  OR2_X1 U12773 ( .A1(n10911), .A2(n10521), .ZN(n10914) );
  AOI22_X1 U12774 ( .A1(n12336), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n12335), 
        .B2(n10912), .ZN(n10913) );
  XNOR2_X1 U12775 ( .A(n12828), .B(n13847), .ZN(n10916) );
  NAND2_X1 U12776 ( .A1(n14018), .A2(n14208), .ZN(n10915) );
  NAND2_X1 U12777 ( .A1(n10916), .A2(n10915), .ZN(n11108) );
  OAI21_X1 U12778 ( .B1(n10916), .B2(n10915), .A(n11108), .ZN(n10917) );
  AOI21_X1 U12779 ( .B1(n10918), .B2(n10917), .A(n11110), .ZN(n10931) );
  INV_X1 U12780 ( .A(n11020), .ZN(n10920) );
  OAI21_X1 U12781 ( .B1(n13995), .B2(n10920), .A(n10919), .ZN(n10929) );
  INV_X1 U12782 ( .A(n14019), .ZN(n11008) );
  NAND2_X1 U12783 ( .A1(n12064), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10927) );
  NAND2_X1 U12784 ( .A1(n12468), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10926) );
  NAND2_X1 U12785 ( .A1(n10922), .A2(n10921), .ZN(n10923) );
  AND2_X1 U12786 ( .A1(n11079), .A2(n10923), .ZN(n11088) );
  NAND2_X1 U12787 ( .A1(n12425), .A2(n11088), .ZN(n10925) );
  NAND2_X1 U12788 ( .A1(n7508), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n10924) );
  NAND4_X1 U12789 ( .A1(n10927), .A2(n10926), .A3(n10925), .A4(n10924), .ZN(
        n14017) );
  INV_X1 U12790 ( .A(n14017), .ZN(n11293) );
  OAI22_X1 U12791 ( .A1(n11008), .A2(n13997), .B1(n13998), .B2(n11293), .ZN(
        n10928) );
  AOI211_X1 U12792 ( .C1(n12828), .C2(n14001), .A(n10929), .B(n10928), .ZN(
        n10930) );
  OAI21_X1 U12793 ( .B1(n10931), .B2(n14003), .A(n10930), .ZN(P2_U3193) );
  INV_X1 U12794 ( .A(n14262), .ZN(n14285) );
  OAI22_X1 U12795 ( .A1(n10933), .A2(n14283), .B1(n14285), .B2(n12807), .ZN(
        n13956) );
  AOI21_X1 U12796 ( .B1(n10934), .B2(n14309), .A(n13956), .ZN(n15781) );
  OAI22_X1 U12797 ( .A1(n14275), .A2(n10530), .B1(n10935), .B2(n14318), .ZN(
        n10938) );
  OAI211_X1 U12798 ( .C1(n10961), .C2(n15782), .A(n10936), .B(n11286), .ZN(
        n15780) );
  NOR2_X1 U12799 ( .A1(n14234), .A2(n15780), .ZN(n10937) );
  AOI211_X1 U12800 ( .C1(n15818), .C2(n13958), .A(n10938), .B(n10937), .ZN(
        n10942) );
  XNOR2_X1 U12801 ( .A(n10940), .B(n10939), .ZN(n15779) );
  INV_X1 U12802 ( .A(n15779), .ZN(n15785) );
  NAND2_X1 U12803 ( .A1(n14315), .A2(n15785), .ZN(n10941) );
  OAI211_X1 U12804 ( .C1(n15829), .C2(n15781), .A(n10942), .B(n10941), .ZN(
        P2_U3261) );
  NAND2_X1 U12805 ( .A1(n10943), .A2(n8086), .ZN(n10944) );
  XOR2_X1 U12806 ( .A(n10945), .B(n10944), .Z(n10951) );
  INV_X1 U12807 ( .A(n14728), .ZN(n16031) );
  AOI22_X1 U12808 ( .A1(n16031), .A2(n14747), .B1(n10946), .B2(n14731), .ZN(
        n10948) );
  AOI22_X1 U12809 ( .A1(n16029), .A2(n14749), .B1(P1_REG3_REG_4__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10947) );
  OAI211_X1 U12810 ( .C1(n10949), .C2(n16041), .A(n10948), .B(n10947), .ZN(
        n10950) );
  AOI21_X1 U12811 ( .B1(n10951), .B2(n16036), .A(n10950), .ZN(n10952) );
  INV_X1 U12812 ( .A(n10952), .ZN(P1_U3230) );
  XNOR2_X1 U12813 ( .A(n10953), .B(n10956), .ZN(n15768) );
  OAI22_X1 U12814 ( .A1(n10955), .A2(n14283), .B1(n14285), .B2(n10954), .ZN(
        n10960) );
  NAND3_X1 U12815 ( .A1(n11097), .A2(n10957), .A3(n10956), .ZN(n10958) );
  AOI211_X1 U12816 ( .C1(n15812), .C2(n15768), .A(n10960), .B(n10959), .ZN(
        n15765) );
  AOI211_X1 U12817 ( .C1(n12794), .C2(n11103), .A(n14208), .B(n10961), .ZN(
        n15762) );
  AOI22_X1 U12818 ( .A1(n15824), .A2(n15768), .B1(n15823), .B2(n15762), .ZN(
        n10965) );
  INV_X1 U12819 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10962) );
  OAI22_X1 U12820 ( .A1(n14275), .A2(n10962), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14318), .ZN(n10963) );
  AOI21_X1 U12821 ( .B1(n15818), .B2(n12794), .A(n10963), .ZN(n10964) );
  OAI211_X1 U12822 ( .C1(n15829), .C2(n15765), .A(n10965), .B(n10964), .ZN(
        P2_U3262) );
  NAND2_X1 U12823 ( .A1(n10966), .A2(n10970), .ZN(n10967) );
  NAND2_X1 U12824 ( .A1(n10968), .A2(n10967), .ZN(n10972) );
  INV_X1 U12825 ( .A(n10972), .ZN(n10988) );
  XNOR2_X1 U12826 ( .A(n10969), .B(n9804), .ZN(n10971) );
  NAND2_X1 U12827 ( .A1(n10971), .A2(n15985), .ZN(n10975) );
  AOI22_X1 U12828 ( .A1(n15033), .A2(n14747), .B1(n14745), .B2(n15034), .ZN(
        n10974) );
  NAND2_X1 U12829 ( .A1(n10972), .A2(n11648), .ZN(n10973) );
  NAND3_X1 U12830 ( .A1(n10975), .A2(n10974), .A3(n10973), .ZN(n10983) );
  MUX2_X1 U12831 ( .A(n10983), .B(P1_REG2_REG_6__SCAN_IN), .S(n15036), .Z(
        n10976) );
  INV_X1 U12832 ( .A(n10976), .ZN(n10982) );
  INV_X1 U12833 ( .A(n11153), .ZN(n10977) );
  AOI21_X1 U12834 ( .B1(n10995), .B2(n10978), .A(n10977), .ZN(n10984) );
  OAI22_X1 U12835 ( .A1(n15680), .A2(n10979), .B1(n10996), .B2(n15035), .ZN(
        n10980) );
  AOI21_X1 U12836 ( .B1(n10984), .B2(n15018), .A(n10980), .ZN(n10981) );
  OAI211_X1 U12837 ( .C1(n10988), .C2(n11391), .A(n10982), .B(n10981), .ZN(
        P1_U3287) );
  INV_X1 U12838 ( .A(n10983), .ZN(n10986) );
  AOI22_X1 U12839 ( .A1(n10984), .A2(n15796), .B1(n16014), .B2(n10995), .ZN(
        n10985) );
  OAI211_X1 U12840 ( .C1(n10988), .C2(n10987), .A(n10986), .B(n10985), .ZN(
        n10990) );
  NAND2_X1 U12841 ( .A1(n10990), .A2(n15922), .ZN(n10989) );
  OAI21_X1 U12842 ( .B1(n15922), .B2(n9944), .A(n10989), .ZN(P1_U3534) );
  NAND2_X1 U12843 ( .A1(n10990), .A2(n15961), .ZN(n10991) );
  OAI21_X1 U12844 ( .B1(n15961), .B2(n9057), .A(n10991), .ZN(P1_U3477) );
  XNOR2_X1 U12845 ( .A(n8088), .B(n10992), .ZN(n10993) );
  XNOR2_X1 U12846 ( .A(n10994), .B(n10993), .ZN(n11003) );
  AOI22_X1 U12847 ( .A1(n16029), .A2(n14747), .B1(P1_REG3_REG_6__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11001) );
  NAND2_X1 U12848 ( .A1(n10995), .A2(n14731), .ZN(n11000) );
  OR2_X1 U12849 ( .A1(n16041), .A2(n10996), .ZN(n10999) );
  OR2_X1 U12850 ( .A1(n10997), .A2(n14728), .ZN(n10998) );
  NAND4_X1 U12851 ( .A1(n11001), .A2(n11000), .A3(n10999), .A4(n10998), .ZN(
        n11002) );
  AOI21_X1 U12852 ( .B1(n11003), .B2(n16036), .A(n11002), .ZN(n11004) );
  INV_X1 U12853 ( .A(n11004), .ZN(P1_U3239) );
  INV_X1 U12854 ( .A(n14020), .ZN(n12815) );
  NAND2_X1 U12855 ( .A1(n15819), .A2(n12815), .ZN(n11006) );
  AND2_X1 U12856 ( .A1(n15844), .A2(n11008), .ZN(n11007) );
  OR2_X1 U12857 ( .A1(n15844), .A2(n11008), .ZN(n11009) );
  INV_X1 U12858 ( .A(n14018), .ZN(n12830) );
  XNOR2_X1 U12859 ( .A(n12828), .B(n12830), .ZN(n13003) );
  NAND2_X1 U12860 ( .A1(n11010), .A2(n13003), .ZN(n11011) );
  NAND2_X1 U12861 ( .A1(n11074), .A2(n11011), .ZN(n11012) );
  NAND2_X1 U12862 ( .A1(n11012), .A2(n14309), .ZN(n11014) );
  AOI22_X1 U12863 ( .A1(n14242), .A2(n14019), .B1(n14262), .B2(n14017), .ZN(
        n11013) );
  NAND2_X1 U12864 ( .A1(n11014), .A2(n11013), .ZN(n15866) );
  MUX2_X1 U12865 ( .A(n15866), .B(P2_REG2_REG_8__SCAN_IN), .S(n15829), .Z(
        n11024) );
  INV_X1 U12866 ( .A(n15844), .ZN(n11034) );
  INV_X1 U12867 ( .A(n12828), .ZN(n15864) );
  OAI211_X1 U12868 ( .C1(n11030), .C2(n15864), .A(n11286), .B(n11090), .ZN(
        n15862) );
  OR2_X1 U12869 ( .A1(n15819), .A2(n14020), .ZN(n11016) );
  OR2_X1 U12870 ( .A1(n15844), .A2(n14019), .ZN(n11026) );
  NAND2_X1 U12871 ( .A1(n15844), .A2(n14019), .ZN(n11025) );
  NAND2_X1 U12872 ( .A1(n11018), .A2(n11025), .ZN(n11019) );
  OR2_X1 U12873 ( .A1(n11019), .A2(n13003), .ZN(n15861) );
  NAND2_X1 U12874 ( .A1(n11019), .A2(n13003), .ZN(n15860) );
  NAND3_X1 U12875 ( .A1(n15861), .A2(n15860), .A3(n14315), .ZN(n11022) );
  AOI22_X1 U12876 ( .A1(n15818), .A2(n12828), .B1(n15816), .B2(n11020), .ZN(
        n11021) );
  OAI211_X1 U12877 ( .C1(n14234), .C2(n15862), .A(n11022), .B(n11021), .ZN(
        n11023) );
  OR2_X1 U12878 ( .A1(n11024), .A2(n11023), .ZN(P2_U3257) );
  NAND2_X1 U12879 ( .A1(n11026), .A2(n11025), .ZN(n13001) );
  XOR2_X1 U12880 ( .A(n13001), .B(n7357), .Z(n15848) );
  XOR2_X1 U12881 ( .A(n13001), .B(n11027), .Z(n11029) );
  OAI21_X1 U12882 ( .B1(n11029), .B2(n14289), .A(n11028), .ZN(n15849) );
  NAND2_X1 U12883 ( .A1(n15849), .A2(n14275), .ZN(n11037) );
  AOI211_X1 U12884 ( .C1(n15844), .C2(n11031), .A(n14208), .B(n11030), .ZN(
        n15843) );
  AOI22_X1 U12885 ( .A1(n15829), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n11032), 
        .B2(n15816), .ZN(n11033) );
  OAI21_X1 U12886 ( .B1(n14301), .B2(n11034), .A(n11033), .ZN(n11035) );
  AOI21_X1 U12887 ( .B1(n15823), .B2(n15843), .A(n11035), .ZN(n11036) );
  OAI211_X1 U12888 ( .C1(n14254), .C2(n15848), .A(n11037), .B(n11036), .ZN(
        P2_U3258) );
  INV_X1 U12889 ( .A(n14797), .ZN(n14803) );
  INV_X1 U12890 ( .A(n12320), .ZN(n11043) );
  OAI222_X1 U12891 ( .A1(P1_U3086), .A2(n14803), .B1(n15215), .B2(n11043), 
        .C1(n11038), .C2(n15210), .ZN(P1_U3338) );
  OR2_X1 U12892 ( .A1(n11040), .A2(n11039), .ZN(n11041) );
  XNOR2_X1 U12893 ( .A(n11041), .B(P2_IR_REG_17__SCAN_IN), .ZN(n15404) );
  INV_X1 U12894 ( .A(n15404), .ZN(n11042) );
  OAI222_X1 U12895 ( .A1(n14509), .A2(n11044), .B1(n14506), .B2(n11043), .C1(
        n11042), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U12896 ( .A(n11045), .ZN(n11046) );
  XNOR2_X1 U12897 ( .A(n11242), .B(n13109), .ZN(n11223) );
  XNOR2_X1 U12898 ( .A(n11223), .B(n11226), .ZN(n11048) );
  AOI21_X1 U12899 ( .B1(n11049), .B2(n11048), .A(n7353), .ZN(n11053) );
  NOR2_X1 U12900 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8428), .ZN(n15557) );
  OAI22_X1 U12901 ( .A1(n11238), .A2(n13237), .B1(n11350), .B2(n13225), .ZN(
        n11050) );
  AOI211_X1 U12902 ( .C1(n11242), .C2(n13206), .A(n15557), .B(n11050), .ZN(
        n11052) );
  NAND2_X1 U12903 ( .A1(n13239), .A2(n11241), .ZN(n11051) );
  OAI211_X1 U12904 ( .C1(n11053), .C2(n13229), .A(n11052), .B(n11051), .ZN(
        P3_U3167) );
  INV_X1 U12905 ( .A(n11062), .ZN(n11189) );
  INV_X1 U12906 ( .A(n15937), .ZN(n13552) );
  INV_X1 U12907 ( .A(n15721), .ZN(n13643) );
  AOI22_X1 U12908 ( .A1(n13643), .A2(n13261), .B1(n13259), .B2(n13642), .ZN(
        n11061) );
  AND2_X1 U12909 ( .A1(n11056), .A2(n11057), .ZN(n11059) );
  OAI211_X1 U12910 ( .C1(n11059), .C2(n12575), .A(n11058), .B(n13640), .ZN(
        n11060) );
  OAI211_X1 U12911 ( .C1(n11189), .C2(n13552), .A(n11061), .B(n11060), .ZN(
        n11184) );
  AOI21_X1 U12912 ( .B1(n15931), .B2(n11062), .A(n11184), .ZN(n11247) );
  INV_X1 U12913 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n11063) );
  OAI22_X1 U12914 ( .A1(n13794), .A2(n11249), .B1(n15944), .B2(n11063), .ZN(
        n11064) );
  INV_X1 U12915 ( .A(n11064), .ZN(n11065) );
  OAI21_X1 U12916 ( .B1(n11247), .B2(n15941), .A(n11065), .ZN(P3_U3399) );
  NAND2_X1 U12917 ( .A1(n12828), .A2(n14018), .ZN(n11066) );
  NAND2_X1 U12918 ( .A1(n15860), .A2(n11066), .ZN(n11071) );
  OR2_X1 U12919 ( .A1(n11067), .A2(n10521), .ZN(n11070) );
  AOI22_X1 U12920 ( .A1(n12336), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n12335), 
        .B2(n11068), .ZN(n11069) );
  XNOR2_X1 U12921 ( .A(n12836), .B(n11293), .ZN(n13004) );
  NAND2_X1 U12922 ( .A1(n11071), .A2(n13004), .ZN(n11122) );
  OR2_X1 U12923 ( .A1(n11071), .A2(n13004), .ZN(n11072) );
  NAND2_X1 U12924 ( .A1(n11122), .A2(n11072), .ZN(n15883) );
  NAND2_X1 U12925 ( .A1(n12828), .A2(n12830), .ZN(n11073) );
  INV_X1 U12926 ( .A(n13004), .ZN(n11075) );
  OAI21_X1 U12927 ( .B1(n11076), .B2(n11075), .A(n11136), .ZN(n11086) );
  NAND2_X1 U12928 ( .A1(n12468), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n11084) );
  NAND2_X1 U12929 ( .A1(n7508), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n11083) );
  INV_X1 U12930 ( .A(n11079), .ZN(n11077) );
  NAND2_X1 U12931 ( .A1(n11077), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n11127) );
  INV_X1 U12932 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n11078) );
  NAND2_X1 U12933 ( .A1(n11079), .A2(n11078), .ZN(n11080) );
  AND2_X1 U12934 ( .A1(n11127), .A2(n11080), .ZN(n11140) );
  NAND2_X1 U12935 ( .A1(n12425), .A2(n11140), .ZN(n11082) );
  NAND2_X1 U12936 ( .A1(n12064), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11081) );
  NAND4_X1 U12937 ( .A1(n11084), .A2(n11083), .A3(n11082), .A4(n11081), .ZN(
        n14016) );
  INV_X1 U12938 ( .A(n14016), .ZN(n12846) );
  OAI22_X1 U12939 ( .A1(n12830), .A2(n14283), .B1(n14285), .B2(n12846), .ZN(
        n11085) );
  AOI21_X1 U12940 ( .B1(n11086), .B2(n14267), .A(n11085), .ZN(n11087) );
  OAI21_X1 U12941 ( .B1(n15778), .B2(n15883), .A(n11087), .ZN(n15886) );
  NAND2_X1 U12942 ( .A1(n15886), .A2(n14275), .ZN(n11095) );
  INV_X1 U12943 ( .A(n11088), .ZN(n11116) );
  OAI22_X1 U12944 ( .A1(n14275), .A2(n11089), .B1(n11116), .B2(n14318), .ZN(
        n11093) );
  INV_X1 U12945 ( .A(n12836), .ZN(n15885) );
  INV_X1 U12946 ( .A(n11090), .ZN(n11091) );
  OAI211_X1 U12947 ( .C1(n15885), .C2(n11091), .A(n11286), .B(n11142), .ZN(
        n15884) );
  NOR2_X1 U12948 ( .A1(n15884), .A2(n14234), .ZN(n11092) );
  AOI211_X1 U12949 ( .C1(n15818), .C2(n12836), .A(n11093), .B(n11092), .ZN(
        n11094) );
  OAI211_X1 U12950 ( .C1(n15883), .C2(n14129), .A(n11095), .B(n11094), .ZN(
        P2_U3256) );
  XNOR2_X1 U12951 ( .A(n11096), .B(n12994), .ZN(n15746) );
  OAI21_X1 U12952 ( .B1(n12994), .B2(n11098), .A(n11097), .ZN(n11100) );
  AOI21_X1 U12953 ( .B1(n11100), .B2(n14309), .A(n11099), .ZN(n15748) );
  INV_X1 U12954 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11101) );
  OAI22_X1 U12955 ( .A1(n15829), .A2(n15748), .B1(n11101), .B2(n14318), .ZN(
        n11106) );
  INV_X1 U12956 ( .A(n11102), .ZN(n11104) );
  OAI211_X1 U12957 ( .C1(n11104), .C2(n15749), .A(n11286), .B(n11103), .ZN(
        n15747) );
  OAI22_X1 U12958 ( .A1(n14301), .A2(n15749), .B1(n15747), .B2(n14234), .ZN(
        n11105) );
  AOI211_X1 U12959 ( .C1(P2_REG2_REG_2__SCAN_IN), .C2(n15817), .A(n11106), .B(
        n11105), .ZN(n11107) );
  OAI21_X1 U12960 ( .B1(n14254), .B2(n15746), .A(n11107), .ZN(P2_U3263) );
  INV_X1 U12961 ( .A(n11108), .ZN(n11109) );
  XNOR2_X1 U12962 ( .A(n12836), .B(n13847), .ZN(n11112) );
  NAND2_X1 U12963 ( .A1(n14017), .A2(n14208), .ZN(n11111) );
  NAND2_X1 U12964 ( .A1(n11112), .A2(n11111), .ZN(n11285) );
  OAI21_X1 U12965 ( .B1(n11112), .B2(n11111), .A(n11285), .ZN(n11113) );
  AOI21_X1 U12966 ( .B1(n11114), .B2(n11113), .A(n7351), .ZN(n11120) );
  OAI21_X1 U12967 ( .B1(n13995), .B2(n11116), .A(n11115), .ZN(n11118) );
  OAI22_X1 U12968 ( .A1(n12830), .A2(n13997), .B1(n13998), .B2(n12846), .ZN(
        n11117) );
  AOI211_X1 U12969 ( .C1(n12836), .C2(n14001), .A(n11118), .B(n11117), .ZN(
        n11119) );
  OAI21_X1 U12970 ( .B1(n11120), .B2(n14003), .A(n11119), .ZN(P2_U3203) );
  NAND2_X1 U12971 ( .A1(n12836), .A2(n14017), .ZN(n11121) );
  AOI22_X1 U12972 ( .A1(n12336), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n11124), 
        .B2(n12335), .ZN(n11125) );
  NAND2_X1 U12973 ( .A1(n12844), .A2(n12846), .ZN(n11126) );
  NAND2_X1 U12974 ( .A1(n11301), .A2(n11126), .ZN(n13005) );
  XNOR2_X1 U12975 ( .A(n11315), .B(n13005), .ZN(n15901) );
  NAND2_X1 U12976 ( .A1(n12064), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n11132) );
  NAND2_X1 U12977 ( .A1(n12468), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n11131) );
  NAND2_X1 U12978 ( .A1(n11127), .A2(n11569), .ZN(n11128) );
  AND2_X1 U12979 ( .A1(n11308), .A2(n11128), .ZN(n11568) );
  NAND2_X1 U12980 ( .A1(n12425), .A2(n11568), .ZN(n11130) );
  NAND2_X1 U12981 ( .A1(n7508), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n11129) );
  NAND4_X1 U12982 ( .A1(n11132), .A2(n11131), .A3(n11130), .A4(n11129), .ZN(
        n14015) );
  AOI22_X1 U12983 ( .A1(n14242), .A2(n14017), .B1(n14262), .B2(n14015), .ZN(
        n11139) );
  INV_X1 U12984 ( .A(n11136), .ZN(n11133) );
  AND2_X1 U12985 ( .A1(n12836), .A2(n11293), .ZN(n11134) );
  OAI21_X1 U12986 ( .B1(n11133), .B2(n11134), .A(n13005), .ZN(n11137) );
  NOR2_X1 U12987 ( .A1(n13005), .A2(n11134), .ZN(n11135) );
  NAND3_X1 U12988 ( .A1(n11137), .A2(n14267), .A3(n11302), .ZN(n11138) );
  OAI211_X1 U12989 ( .C1(n15901), .C2(n15778), .A(n11139), .B(n11138), .ZN(
        n15904) );
  NAND2_X1 U12990 ( .A1(n15904), .A2(n14275), .ZN(n11148) );
  INV_X1 U12991 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11141) );
  INV_X1 U12992 ( .A(n11140), .ZN(n11292) );
  OAI22_X1 U12993 ( .A1(n14275), .A2(n11141), .B1(n11292), .B2(n14318), .ZN(
        n11146) );
  INV_X1 U12994 ( .A(n11142), .ZN(n11144) );
  INV_X1 U12995 ( .A(n11322), .ZN(n11143) );
  OAI211_X1 U12996 ( .C1(n15903), .C2(n11144), .A(n11143), .B(n11286), .ZN(
        n15902) );
  NOR2_X1 U12997 ( .A1(n15902), .A2(n14234), .ZN(n11145) );
  AOI211_X1 U12998 ( .C1(n15818), .C2(n12844), .A(n11146), .B(n11145), .ZN(
        n11147) );
  OAI211_X1 U12999 ( .C1(n15901), .C2(n14129), .A(n11148), .B(n11147), .ZN(
        P2_U3255) );
  OR2_X1 U13000 ( .A1(n11149), .A2(n11159), .ZN(n11150) );
  NAND2_X1 U13001 ( .A1(n11151), .A2(n11150), .ZN(n15841) );
  INV_X1 U13002 ( .A(n11152), .ZN(n11155) );
  NAND2_X1 U13003 ( .A1(n11153), .A2(n15836), .ZN(n11154) );
  NAND2_X1 U13004 ( .A1(n11155), .A2(n11154), .ZN(n15838) );
  INV_X1 U13005 ( .A(n11156), .ZN(n11157) );
  AOI22_X1 U13006 ( .A1(n15061), .A2(n15836), .B1(n15678), .B2(n11157), .ZN(
        n11158) );
  OAI21_X1 U13007 ( .B1(n15838), .B2(n15681), .A(n11158), .ZN(n11166) );
  XNOR2_X1 U13008 ( .A(n11160), .B(n11159), .ZN(n11161) );
  NAND2_X1 U13009 ( .A1(n11161), .A2(n15985), .ZN(n11164) );
  NAND2_X1 U13010 ( .A1(n15841), .A2(n11648), .ZN(n11163) );
  AOI22_X1 U13011 ( .A1(n15033), .A2(n14746), .B1(n14744), .B2(n15034), .ZN(
        n11162) );
  NAND3_X1 U13012 ( .A1(n11164), .A2(n11163), .A3(n11162), .ZN(n15839) );
  MUX2_X1 U13013 ( .A(n15839), .B(P1_REG2_REG_7__SCAN_IN), .S(n15036), .Z(
        n11165) );
  AOI211_X1 U13014 ( .C1(n15684), .C2(n15841), .A(n11166), .B(n11165), .ZN(
        n11167) );
  INV_X1 U13015 ( .A(n11167), .ZN(P1_U3286) );
  INV_X1 U13016 ( .A(n11168), .ZN(n11169) );
  AOI21_X1 U13017 ( .B1(n12576), .B2(n11170), .A(n11169), .ZN(n15694) );
  INV_X1 U13018 ( .A(n15931), .ZN(n15895) );
  OAI21_X1 U13019 ( .B1(n12576), .B2(n11171), .A(n15716), .ZN(n11176) );
  OAI22_X1 U13020 ( .A1(n11173), .A2(n15721), .B1(n11172), .B2(n15723), .ZN(
        n11175) );
  NOR2_X1 U13021 ( .A1(n15694), .A2(n13552), .ZN(n11174) );
  AOI211_X1 U13022 ( .C1(n13640), .C2(n11176), .A(n11175), .B(n11174), .ZN(
        n15698) );
  OAI21_X1 U13023 ( .B1(n15694), .B2(n15895), .A(n15698), .ZN(n11181) );
  INV_X1 U13024 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n11177) );
  OAI22_X1 U13025 ( .A1(n13794), .A2(n15697), .B1(n15944), .B2(n11177), .ZN(
        n11178) );
  AOI21_X1 U13026 ( .B1(n11181), .B2(n15944), .A(n11178), .ZN(n11179) );
  INV_X1 U13027 ( .A(n11179), .ZN(P3_U3393) );
  OAI22_X1 U13028 ( .A1(n13738), .A2(n15697), .B1(n15940), .B2(n10250), .ZN(
        n11180) );
  AOI21_X1 U13029 ( .B1(n11181), .B2(n15940), .A(n11180), .ZN(n11182) );
  INV_X1 U13030 ( .A(n11182), .ZN(P3_U3460) );
  AND2_X1 U13031 ( .A1(n11183), .A2(n12612), .ZN(n15702) );
  NAND2_X1 U13032 ( .A1(n15735), .A2(n15702), .ZN(n12002) );
  INV_X1 U13033 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11406) );
  INV_X1 U13034 ( .A(n11184), .ZN(n11185) );
  MUX2_X1 U13035 ( .A(n11406), .B(n11185), .S(n15735), .Z(n11188) );
  AOI22_X1 U13036 ( .A1(n13663), .A2(n11186), .B1(n13648), .B2(n11880), .ZN(
        n11187) );
  OAI211_X1 U13037 ( .C1(n11189), .C2(n12002), .A(n11188), .B(n11187), .ZN(
        P3_U3230) );
  OAI21_X1 U13038 ( .B1(n11191), .B2(n12626), .A(n11190), .ZN(n15773) );
  INV_X1 U13039 ( .A(n15773), .ZN(n11200) );
  INV_X1 U13040 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11412) );
  XNOR2_X1 U13041 ( .A(n11193), .B(n11192), .ZN(n11195) );
  AOI22_X1 U13042 ( .A1(n13643), .A2(n13260), .B1(n13258), .B2(n13642), .ZN(
        n11194) );
  OAI21_X1 U13043 ( .B1(n11195), .B2(n15719), .A(n11194), .ZN(n11196) );
  AOI21_X1 U13044 ( .B1(n15937), .B2(n15773), .A(n11196), .ZN(n15775) );
  MUX2_X1 U13045 ( .A(n11412), .B(n15775), .S(n15735), .Z(n11199) );
  AOI22_X1 U13046 ( .A1(n13663), .A2(n15772), .B1(n13648), .B2(n11197), .ZN(
        n11198) );
  OAI211_X1 U13047 ( .C1(n11200), .C2(n12002), .A(n11199), .B(n11198), .ZN(
        P3_U3229) );
  INV_X1 U13048 ( .A(n11201), .ZN(n11203) );
  NAND2_X1 U13049 ( .A1(n11377), .A2(n14614), .ZN(n11207) );
  NAND2_X1 U13050 ( .A1(n14744), .A2(n14659), .ZN(n11206) );
  NAND2_X1 U13051 ( .A1(n11207), .A2(n11206), .ZN(n11208) );
  XNOR2_X1 U13052 ( .A(n11208), .B(n14584), .ZN(n11213) );
  NAND2_X1 U13053 ( .A1(n11377), .A2(n14659), .ZN(n11211) );
  NAND2_X1 U13054 ( .A1(n14744), .A2(n14607), .ZN(n11210) );
  NAND2_X1 U13055 ( .A1(n11211), .A2(n11210), .ZN(n11212) );
  NOR2_X1 U13056 ( .A1(n11213), .A2(n11212), .ZN(n11250) );
  AOI21_X1 U13057 ( .B1(n11213), .B2(n11212), .A(n11250), .ZN(n11214) );
  NAND2_X1 U13058 ( .A1(n11215), .A2(n11214), .ZN(n11252) );
  OAI21_X1 U13059 ( .B1(n11215), .B2(n11214), .A(n11252), .ZN(n11216) );
  NAND2_X1 U13060 ( .A1(n11216), .A2(n16036), .ZN(n11222) );
  NOR2_X1 U13061 ( .A1(n16041), .A2(n11217), .ZN(n11220) );
  OAI21_X1 U13062 ( .B1(n14728), .B2(n11485), .A(n11218), .ZN(n11219) );
  AOI211_X1 U13063 ( .C1(n16029), .C2(n14745), .A(n11220), .B(n11219), .ZN(
        n11221) );
  OAI211_X1 U13064 ( .C1(n11339), .C2(n16033), .A(n11222), .B(n11221), .ZN(
        P1_U3221) );
  INV_X1 U13065 ( .A(n11333), .ZN(n11230) );
  XNOR2_X1 U13066 ( .A(n11277), .B(n13109), .ZN(n11347) );
  XNOR2_X1 U13067 ( .A(n11347), .B(n11350), .ZN(n11224) );
  NAND2_X1 U13068 ( .A1(n11225), .A2(n11224), .ZN(n11348) );
  OAI211_X1 U13069 ( .C1(n11225), .C2(n11224), .A(n11348), .B(n13221), .ZN(
        n11229) );
  INV_X1 U13070 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n11802) );
  NOR2_X1 U13071 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11802), .ZN(n15569) );
  OAI22_X1 U13072 ( .A1(n11996), .A2(n13225), .B1(n11226), .B2(n13237), .ZN(
        n11227) );
  AOI211_X1 U13073 ( .C1(n11334), .C2(n13206), .A(n15569), .B(n11227), .ZN(
        n11228) );
  OAI211_X1 U13074 ( .C1(n11230), .C2(n12169), .A(n11229), .B(n11228), .ZN(
        P3_U3179) );
  INV_X1 U13075 ( .A(n11231), .ZN(n11233) );
  OAI222_X1 U13076 ( .A1(n12036), .A2(n11233), .B1(n13810), .B2(n11828), .C1(
        P3_U3151), .C2(n11232), .ZN(P3_U3271) );
  INV_X1 U13077 ( .A(n11234), .ZN(n11235) );
  AOI21_X1 U13078 ( .B1(n12632), .B2(n11236), .A(n11235), .ZN(n11237) );
  OAI222_X1 U13079 ( .A1(n15723), .A2(n11350), .B1(n15721), .B2(n11238), .C1(
        n15719), .C2(n11237), .ZN(n15790) );
  INV_X1 U13080 ( .A(n15790), .ZN(n11246) );
  OAI21_X1 U13081 ( .B1(n11240), .B2(n12632), .A(n11239), .ZN(n15792) );
  OR2_X1 U13082 ( .A1(n15937), .A2(n15702), .ZN(n15734) );
  INV_X1 U13083 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15551) );
  AOI22_X1 U13084 ( .A1(n13663), .A2(n11242), .B1(n13648), .B2(n11241), .ZN(
        n11243) );
  OAI21_X1 U13085 ( .B1(n15551), .B2(n15735), .A(n11243), .ZN(n11244) );
  AOI21_X1 U13086 ( .B1(n15792), .B2(n13667), .A(n11244), .ZN(n11245) );
  OAI21_X1 U13087 ( .B1(n11246), .B2(n13670), .A(n11245), .ZN(P3_U3228) );
  INV_X1 U13088 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11405) );
  MUX2_X1 U13089 ( .A(n11405), .B(n11247), .S(n15940), .Z(n11248) );
  OAI21_X1 U13090 ( .B1(n13738), .B2(n11249), .A(n11248), .ZN(P3_U3462) );
  INV_X1 U13091 ( .A(n11250), .ZN(n11251) );
  NAND2_X1 U13092 ( .A1(n11252), .A2(n11251), .ZN(n11501) );
  NAND2_X1 U13093 ( .A1(n11486), .A2(n14614), .ZN(n11254) );
  NAND2_X1 U13094 ( .A1(n14743), .A2(n14659), .ZN(n11253) );
  NAND2_X1 U13095 ( .A1(n11254), .A2(n11253), .ZN(n11255) );
  XNOR2_X1 U13096 ( .A(n11255), .B(n14661), .ZN(n11259) );
  NAND2_X1 U13097 ( .A1(n11486), .A2(n14659), .ZN(n11257) );
  NAND2_X1 U13098 ( .A1(n14743), .A2(n14607), .ZN(n11256) );
  NAND2_X1 U13099 ( .A1(n11257), .A2(n11256), .ZN(n11258) );
  NAND2_X1 U13100 ( .A1(n11259), .A2(n11258), .ZN(n11500) );
  NAND2_X1 U13101 ( .A1(n7349), .A2(n11500), .ZN(n11260) );
  XNOR2_X1 U13102 ( .A(n11501), .B(n11260), .ZN(n11266) );
  NOR2_X1 U13103 ( .A1(n16041), .A2(n11387), .ZN(n11264) );
  NAND2_X1 U13104 ( .A1(n16031), .A2(n14742), .ZN(n11262) );
  OAI211_X1 U13105 ( .C1(n14701), .C2(n11376), .A(n11262), .B(n11261), .ZN(
        n11263) );
  AOI211_X1 U13106 ( .C1(n11486), .C2(n14731), .A(n11264), .B(n11263), .ZN(
        n11265) );
  OAI21_X1 U13107 ( .B1(n11266), .B2(n14733), .A(n11265), .ZN(P1_U3231) );
  XNOR2_X1 U13108 ( .A(n11267), .B(n12637), .ZN(n11330) );
  NAND2_X1 U13109 ( .A1(n11268), .A2(n13640), .ZN(n11273) );
  AOI21_X1 U13110 ( .B1(n11234), .B2(n11270), .A(n11269), .ZN(n11272) );
  AOI22_X1 U13111 ( .A1(n13258), .A2(n13643), .B1(n13642), .B2(n13256), .ZN(
        n11271) );
  OAI21_X1 U13112 ( .B1(n11273), .B2(n11272), .A(n11271), .ZN(n11331) );
  AOI21_X1 U13113 ( .B1(n11330), .B2(n15912), .A(n11331), .ZN(n11280) );
  INV_X1 U13114 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11459) );
  OAI22_X1 U13115 ( .A1(n13738), .A2(n11277), .B1(n15940), .B2(n11459), .ZN(
        n11274) );
  INV_X1 U13116 ( .A(n11274), .ZN(n11275) );
  OAI21_X1 U13117 ( .B1(n11280), .B2(n15939), .A(n11275), .ZN(P3_U3465) );
  INV_X1 U13118 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n11276) );
  OAI22_X1 U13119 ( .A1(n13794), .A2(n11277), .B1(n15944), .B2(n11276), .ZN(
        n11278) );
  INV_X1 U13120 ( .A(n11278), .ZN(n11279) );
  OAI21_X1 U13121 ( .B1(n11280), .B2(n15941), .A(n11279), .ZN(P3_U3408) );
  INV_X1 U13122 ( .A(n14814), .ZN(n14808) );
  OAI222_X1 U13123 ( .A1(n15210), .A2(n11281), .B1(n15215), .B2(n11283), .C1(
        n14808), .C2(P1_U3086), .ZN(P1_U3337) );
  XNOR2_X1 U13124 ( .A(n11282), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14060) );
  INV_X1 U13125 ( .A(n14060), .ZN(n14068) );
  OAI222_X1 U13126 ( .A1(n14509), .A2(n11284), .B1(n14506), .B2(n11283), .C1(
        n14068), .C2(P2_U3088), .ZN(P2_U3309) );
  XNOR2_X1 U13127 ( .A(n12844), .B(n13847), .ZN(n11288) );
  NAND2_X1 U13128 ( .A1(n14016), .A2(n14295), .ZN(n11287) );
  NAND2_X1 U13129 ( .A1(n11288), .A2(n11287), .ZN(n11566) );
  OAI21_X1 U13130 ( .B1(n11288), .B2(n11287), .A(n11566), .ZN(n11289) );
  AOI21_X1 U13131 ( .B1(n11290), .B2(n11289), .A(n11567), .ZN(n11297) );
  OAI21_X1 U13132 ( .B1(n13995), .B2(n11292), .A(n11291), .ZN(n11295) );
  INV_X1 U13133 ( .A(n14015), .ZN(n11963) );
  OAI22_X1 U13134 ( .A1(n11293), .A2(n13997), .B1(n13998), .B2(n11963), .ZN(
        n11294) );
  AOI211_X1 U13135 ( .C1(n12844), .C2(n14001), .A(n11295), .B(n11294), .ZN(
        n11296) );
  OAI21_X1 U13136 ( .B1(n11297), .B2(n14003), .A(n11296), .ZN(P2_U3189) );
  NAND2_X1 U13137 ( .A1(n11298), .A2(n12959), .ZN(n11300) );
  AOI22_X1 U13138 ( .A1(n11361), .A2(n12335), .B1(n12336), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n11299) );
  XNOR2_X1 U13139 ( .A(n12851), .B(n14015), .ZN(n13006) );
  INV_X1 U13140 ( .A(n13006), .ZN(n11305) );
  INV_X1 U13141 ( .A(n11529), .ZN(n11303) );
  AOI21_X1 U13142 ( .B1(n11305), .B2(n11304), .A(n11303), .ZN(n11321) );
  NAND2_X1 U13143 ( .A1(n12468), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n11313) );
  NAND2_X1 U13144 ( .A1(n7508), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n11312) );
  INV_X1 U13145 ( .A(n11308), .ZN(n11306) );
  NAND2_X1 U13146 ( .A1(n11306), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n11521) );
  INV_X1 U13147 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n11307) );
  NAND2_X1 U13148 ( .A1(n11308), .A2(n11307), .ZN(n11309) );
  AND2_X1 U13149 ( .A1(n11521), .A2(n11309), .ZN(n11966) );
  NAND2_X1 U13150 ( .A1(n12425), .A2(n11966), .ZN(n11311) );
  NAND2_X1 U13151 ( .A1(n12064), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n11310) );
  NAND4_X1 U13152 ( .A1(n11313), .A2(n11312), .A3(n11311), .A4(n11310), .ZN(
        n14014) );
  AOI22_X1 U13153 ( .A1(n14242), .A2(n14016), .B1(n14262), .B2(n14014), .ZN(
        n11320) );
  INV_X1 U13154 ( .A(n13005), .ZN(n11314) );
  NAND2_X1 U13155 ( .A1(n15903), .A2(n12846), .ZN(n11316) );
  NAND2_X1 U13156 ( .A1(n11317), .A2(n13006), .ZN(n11318) );
  NAND2_X1 U13157 ( .A1(n15928), .A2(n15812), .ZN(n11319) );
  OAI211_X1 U13158 ( .C1(n11321), .C2(n14289), .A(n11320), .B(n11319), .ZN(
        n15926) );
  INV_X1 U13159 ( .A(n15926), .ZN(n11327) );
  INV_X1 U13160 ( .A(n12851), .ZN(n15925) );
  OAI211_X1 U13161 ( .C1(n15925), .C2(n11322), .A(n11286), .B(n11535), .ZN(
        n15924) );
  AOI22_X1 U13162 ( .A1(n15829), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11568), 
        .B2(n15816), .ZN(n11324) );
  NAND2_X1 U13163 ( .A1(n12851), .A2(n15818), .ZN(n11323) );
  OAI211_X1 U13164 ( .C1(n15924), .C2(n14234), .A(n11324), .B(n11323), .ZN(
        n11325) );
  AOI21_X1 U13165 ( .B1(n15928), .B2(n15824), .A(n11325), .ZN(n11326) );
  OAI21_X1 U13166 ( .B1(n11327), .B2(n15817), .A(n11326), .ZN(P2_U3254) );
  OAI222_X1 U13167 ( .A1(n12036), .A2(n11329), .B1(n13810), .B2(n11713), .C1(
        P3_U3151), .C2(n11328), .ZN(P3_U3270) );
  INV_X1 U13168 ( .A(n11330), .ZN(n11337) );
  INV_X1 U13169 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11423) );
  INV_X1 U13170 ( .A(n11331), .ZN(n11332) );
  MUX2_X1 U13171 ( .A(n11423), .B(n11332), .S(n15735), .Z(n11336) );
  AOI22_X1 U13172 ( .A1(n13663), .A2(n11334), .B1(n13648), .B2(n11333), .ZN(
        n11335) );
  OAI211_X1 U13173 ( .C1(n11337), .C2(n13653), .A(n11336), .B(n11335), .ZN(
        P3_U3227) );
  INV_X1 U13174 ( .A(n11338), .ZN(n11343) );
  OAI22_X1 U13175 ( .A1(n11340), .A2(n16009), .B1(n11339), .B2(n15954), .ZN(
        n11342) );
  AOI211_X1 U13176 ( .C1(n15881), .C2(n11343), .A(n11342), .B(n11341), .ZN(
        n11345) );
  OR2_X1 U13177 ( .A1(n11345), .A2(n16023), .ZN(n11344) );
  OAI21_X1 U13178 ( .B1(n15961), .B2(n9092), .A(n11344), .ZN(P1_U3483) );
  OR2_X1 U13179 ( .A1(n11345), .A2(n16021), .ZN(n11346) );
  OAI21_X1 U13180 ( .B1(n15922), .B2(n7665), .A(n11346), .ZN(P1_U3536) );
  INV_X1 U13181 ( .A(n11347), .ZN(n11349) );
  XNOR2_X1 U13182 ( .A(n13109), .B(n15830), .ZN(n11575) );
  XNOR2_X1 U13183 ( .A(n11575), .B(n11996), .ZN(n11576) );
  XNOR2_X1 U13184 ( .A(n11577), .B(n11576), .ZN(n11354) );
  INV_X1 U13185 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n11876) );
  NOR2_X1 U13186 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11876), .ZN(n15591) );
  OAI22_X1 U13187 ( .A1(n12009), .A2(n13225), .B1(n11350), .B2(n13237), .ZN(
        n11351) );
  AOI211_X1 U13188 ( .C1(n11639), .C2(n13206), .A(n15591), .B(n11351), .ZN(
        n11353) );
  NAND2_X1 U13189 ( .A1(n13239), .A2(n11638), .ZN(n11352) );
  OAI211_X1 U13190 ( .C1(n11354), .C2(n13229), .A(n11353), .B(n11352), .ZN(
        P3_U3153) );
  INV_X1 U13191 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11356) );
  MUX2_X1 U13192 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n11356), .S(n15422), .Z(
        n15417) );
  OAI21_X1 U13193 ( .B1(n15422), .B2(P2_REG1_REG_12__SCAN_IN), .A(n15416), 
        .ZN(n11359) );
  INV_X1 U13194 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n12152) );
  NOR2_X1 U13195 ( .A1(n11701), .A2(n12152), .ZN(n11357) );
  AOI21_X1 U13196 ( .B1(n12152), .B2(n11701), .A(n11357), .ZN(n11358) );
  NOR2_X1 U13197 ( .A1(n11358), .A2(n11359), .ZN(n11695) );
  AOI211_X1 U13198 ( .C1(n11359), .C2(n11358), .A(n11695), .B(n15387), .ZN(
        n11371) );
  OAI21_X1 U13199 ( .B1(n11361), .B2(P2_REG2_REG_11__SCAN_IN), .A(n11360), 
        .ZN(n15414) );
  NOR2_X1 U13200 ( .A1(n15422), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n11362) );
  AOI21_X1 U13201 ( .B1(n15422), .B2(P2_REG2_REG_12__SCAN_IN), .A(n11362), 
        .ZN(n15415) );
  NAND2_X1 U13202 ( .A1(n15414), .A2(n15415), .ZN(n15413) );
  OAI21_X1 U13203 ( .B1(n15422), .B2(P2_REG2_REG_12__SCAN_IN), .A(n15413), 
        .ZN(n11366) );
  INV_X1 U13204 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11364) );
  NOR2_X1 U13205 ( .A1(n11701), .A2(n11364), .ZN(n11363) );
  AOI21_X1 U13206 ( .B1(n11701), .B2(n11364), .A(n11363), .ZN(n11365) );
  NOR2_X1 U13207 ( .A1(n11365), .A2(n11366), .ZN(n11700) );
  AOI211_X1 U13208 ( .C1(n11366), .C2(n11365), .A(n11700), .B(n15406), .ZN(
        n11370) );
  NAND2_X1 U13209 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n12099)
         );
  NAND2_X1 U13210 ( .A1(n15341), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n11367) );
  OAI211_X1 U13211 ( .C1(n14074), .C2(n11368), .A(n12099), .B(n11367), .ZN(
        n11369) );
  OR3_X1 U13212 ( .A1(n11371), .A2(n11370), .A3(n11369), .ZN(P2_U3227) );
  NAND2_X1 U13213 ( .A1(n11377), .A2(n14744), .ZN(n11372) );
  AND2_X1 U13214 ( .A1(n11374), .A2(n11372), .ZN(n11375) );
  AND2_X1 U13215 ( .A1(n11380), .A2(n11372), .ZN(n11373) );
  NAND2_X1 U13216 ( .A1(n11374), .A2(n11373), .ZN(n11556) );
  OAI21_X1 U13217 ( .B1(n11375), .B2(n11380), .A(n11556), .ZN(n15880) );
  INV_X1 U13218 ( .A(n15880), .ZN(n11392) );
  OR2_X1 U13219 ( .A1(n11377), .A2(n11376), .ZN(n11378) );
  INV_X1 U13220 ( .A(n11380), .ZN(n11381) );
  XNOR2_X1 U13221 ( .A(n11484), .B(n11381), .ZN(n11384) );
  NAND2_X1 U13222 ( .A1(n15880), .A2(n11648), .ZN(n11383) );
  AOI22_X1 U13223 ( .A1(n15033), .A2(n14744), .B1(n14742), .B2(n15034), .ZN(
        n11382) );
  OAI211_X1 U13224 ( .C1(n11384), .C2(n16016), .A(n11383), .B(n11382), .ZN(
        n15878) );
  MUX2_X1 U13225 ( .A(n15878), .B(P1_REG2_REG_9__SCAN_IN), .S(n15036), .Z(
        n11385) );
  INV_X1 U13226 ( .A(n11385), .ZN(n11390) );
  AOI211_X1 U13227 ( .C1(n11486), .C2(n11386), .A(n16009), .B(n11478), .ZN(
        n15875) );
  NOR2_X1 U13228 ( .A1(n15020), .A2(n9348), .ZN(n14917) );
  OAI22_X1 U13229 ( .A1(n15877), .A2(n15680), .B1(n15035), .B2(n11387), .ZN(
        n11388) );
  AOI21_X1 U13230 ( .B1(n15875), .B2(n14917), .A(n11388), .ZN(n11389) );
  OAI211_X1 U13231 ( .C1(n11392), .C2(n11391), .A(n11390), .B(n11389), .ZN(
        P1_U3284) );
  INV_X1 U13232 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11404) );
  NOR2_X1 U13233 ( .A1(n15511), .A2(n11406), .ZN(n15510) );
  AOI21_X1 U13234 ( .B1(n11456), .B2(n11394), .A(n15510), .ZN(n15529) );
  MUX2_X1 U13235 ( .A(n11412), .B(P3_REG2_REG_4__SCAN_IN), .S(n15540), .Z(
        n11395) );
  INV_X1 U13236 ( .A(n11395), .ZN(n15528) );
  MUX2_X1 U13237 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n11423), .S(n11460), .Z(
        n11396) );
  INV_X1 U13238 ( .A(n11396), .ZN(n15567) );
  INV_X1 U13239 ( .A(n11397), .ZN(n11398) );
  INV_X1 U13240 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n15590) );
  INV_X1 U13241 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U13242 ( .A1(n11463), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n11399), 
        .B2(n15617), .ZN(n15610) );
  NOR2_X1 U13243 ( .A1(n11438), .A2(n11400), .ZN(n11401) );
  INV_X1 U13244 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15630) );
  XNOR2_X1 U13245 ( .A(n11400), .B(n11438), .ZN(n15629) );
  NOR2_X1 U13246 ( .A1(n15630), .A2(n15629), .ZN(n15628) );
  NAND2_X1 U13247 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n15658), .ZN(n11402) );
  OAI21_X1 U13248 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n15658), .A(n11402), 
        .ZN(n15648) );
  AOI21_X1 U13249 ( .B1(n11404), .B2(n11403), .A(n11668), .ZN(n11474) );
  NAND2_X1 U13250 ( .A1(n15517), .A2(n15516), .ZN(n11410) );
  MUX2_X1 U13251 ( .A(n11406), .B(n11405), .S(n13408), .Z(n11407) );
  NAND2_X1 U13252 ( .A1(n11407), .A2(n15521), .ZN(n15535) );
  INV_X1 U13253 ( .A(n11407), .ZN(n11408) );
  NAND2_X1 U13254 ( .A1(n11408), .A2(n11456), .ZN(n11409) );
  AND2_X1 U13255 ( .A1(n15535), .A2(n11409), .ZN(n15514) );
  NAND2_X1 U13256 ( .A1(n11410), .A2(n15514), .ZN(n15536) );
  NAND2_X1 U13257 ( .A1(n15536), .A2(n15535), .ZN(n11417) );
  INV_X1 U13258 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11411) );
  MUX2_X1 U13259 ( .A(n11412), .B(n11411), .S(n13408), .Z(n11413) );
  NAND2_X1 U13260 ( .A1(n11413), .A2(n15540), .ZN(n15554) );
  INV_X1 U13261 ( .A(n11413), .ZN(n11415) );
  NAND2_X1 U13262 ( .A1(n11415), .A2(n11414), .ZN(n11416) );
  AND2_X1 U13263 ( .A1(n15554), .A2(n11416), .ZN(n15533) );
  NAND2_X1 U13264 ( .A1(n11417), .A2(n15533), .ZN(n15555) );
  NAND2_X1 U13265 ( .A1(n15555), .A2(n15554), .ZN(n11422) );
  INV_X1 U13266 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n11418) );
  MUX2_X1 U13267 ( .A(n15551), .B(n11418), .S(n13408), .Z(n11419) );
  NAND2_X1 U13268 ( .A1(n11419), .A2(n11457), .ZN(n15574) );
  INV_X1 U13269 ( .A(n11419), .ZN(n11420) );
  NAND2_X1 U13270 ( .A1(n11420), .A2(n7678), .ZN(n11421) );
  AND2_X1 U13271 ( .A1(n15574), .A2(n11421), .ZN(n15552) );
  NAND2_X1 U13272 ( .A1(n11422), .A2(n15552), .ZN(n15575) );
  NAND2_X1 U13273 ( .A1(n15575), .A2(n15574), .ZN(n11427) );
  MUX2_X1 U13274 ( .A(n11423), .B(n11459), .S(n13408), .Z(n11424) );
  INV_X1 U13275 ( .A(n11460), .ZN(n15579) );
  NAND2_X1 U13276 ( .A1(n11424), .A2(n15579), .ZN(n15596) );
  INV_X1 U13277 ( .A(n11424), .ZN(n11425) );
  NAND2_X1 U13278 ( .A1(n11425), .A2(n11460), .ZN(n11426) );
  AND2_X1 U13279 ( .A1(n15596), .A2(n11426), .ZN(n15572) );
  NAND2_X1 U13280 ( .A1(n11427), .A2(n15572), .ZN(n15597) );
  NAND2_X1 U13281 ( .A1(n15597), .A2(n15596), .ZN(n11431) );
  INV_X1 U13282 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15603) );
  MUX2_X1 U13283 ( .A(n15590), .B(n15603), .S(n13408), .Z(n11428) );
  NAND2_X1 U13284 ( .A1(n11428), .A2(n15601), .ZN(n15611) );
  INV_X1 U13285 ( .A(n11428), .ZN(n11429) );
  NAND2_X1 U13286 ( .A1(n11429), .A2(n11461), .ZN(n11430) );
  AND2_X1 U13287 ( .A1(n15611), .A2(n11430), .ZN(n15594) );
  NAND2_X1 U13288 ( .A1(n11431), .A2(n15594), .ZN(n15615) );
  NAND2_X1 U13289 ( .A1(n15615), .A2(n15611), .ZN(n11436) );
  INV_X1 U13290 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11432) );
  MUX2_X1 U13291 ( .A(n11399), .B(n11432), .S(n13408), .Z(n11433) );
  NAND2_X1 U13292 ( .A1(n11433), .A2(n11463), .ZN(n15631) );
  INV_X1 U13293 ( .A(n11433), .ZN(n11434) );
  NAND2_X1 U13294 ( .A1(n11434), .A2(n15617), .ZN(n11435) );
  AND2_X1 U13295 ( .A1(n15631), .A2(n11435), .ZN(n15613) );
  NAND2_X1 U13296 ( .A1(n15635), .A2(n15631), .ZN(n11442) );
  INV_X1 U13297 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11437) );
  MUX2_X1 U13298 ( .A(n15630), .B(n11437), .S(n13408), .Z(n11439) );
  NAND2_X1 U13299 ( .A1(n11439), .A2(n11438), .ZN(n15650) );
  INV_X1 U13300 ( .A(n11439), .ZN(n11440) );
  NAND2_X1 U13301 ( .A1(n11440), .A2(n15637), .ZN(n11441) );
  AND2_X1 U13302 ( .A1(n15650), .A2(n11441), .ZN(n15633) );
  NAND2_X1 U13303 ( .A1(n11442), .A2(n15633), .ZN(n15655) );
  NAND2_X1 U13304 ( .A1(n15655), .A2(n15650), .ZN(n11448) );
  INV_X1 U13305 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11444) );
  INV_X1 U13306 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11443) );
  MUX2_X1 U13307 ( .A(n11444), .B(n11443), .S(n13408), .Z(n11445) );
  NAND2_X1 U13308 ( .A1(n11445), .A2(n11452), .ZN(n11449) );
  INV_X1 U13309 ( .A(n11445), .ZN(n11446) );
  NAND2_X1 U13310 ( .A1(n11446), .A2(n15658), .ZN(n11447) );
  AND2_X1 U13311 ( .A1(n11449), .A2(n11447), .ZN(n15652) );
  NAND2_X1 U13312 ( .A1(n11448), .A2(n15652), .ZN(n15653) );
  NAND2_X1 U13313 ( .A1(n15653), .A2(n11449), .ZN(n11451) );
  MUX2_X1 U13314 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13408), .Z(n11681) );
  XNOR2_X1 U13315 ( .A(n11681), .B(n11682), .ZN(n11450) );
  OAI21_X1 U13316 ( .B1(n11451), .B2(n11450), .A(n11687), .ZN(n11472) );
  NAND2_X1 U13317 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n15658), .ZN(n11466) );
  AOI22_X1 U13318 ( .A1(n11452), .A2(n11443), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n15658), .ZN(n15665) );
  AOI22_X1 U13319 ( .A1(n11463), .A2(n11432), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n15617), .ZN(n15622) );
  OAI21_X1 U13320 ( .B1(n11454), .B2(n10305), .A(n11453), .ZN(n11455) );
  XNOR2_X1 U13321 ( .A(n11455), .B(n15521), .ZN(n15522) );
  AOI22_X1 U13322 ( .A1(n15522), .A2(P3_REG1_REG_3__SCAN_IN), .B1(n11456), 
        .B2(n11455), .ZN(n15544) );
  MUX2_X1 U13323 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n11411), .S(n15540), .Z(
        n15543) );
  OR2_X1 U13324 ( .A1(n15544), .A2(n15543), .ZN(n15541) );
  OAI21_X1 U13325 ( .B1(n15540), .B2(n11411), .A(n15541), .ZN(n11458) );
  XNOR2_X1 U13326 ( .A(n11458), .B(n11457), .ZN(n15561) );
  AOI22_X1 U13327 ( .A1(n15561), .A2(P3_REG1_REG_5__SCAN_IN), .B1(n7678), .B2(
        n11458), .ZN(n15582) );
  MUX2_X1 U13328 ( .A(n11459), .B(P3_REG1_REG_6__SCAN_IN), .S(n11460), .Z(
        n15581) );
  NOR2_X1 U13329 ( .A1(n15582), .A2(n15581), .ZN(n15580) );
  AOI21_X1 U13330 ( .B1(n11460), .B2(P3_REG1_REG_6__SCAN_IN), .A(n15580), .ZN(
        n11462) );
  OAI21_X1 U13331 ( .B1(n11463), .B2(n11432), .A(n15621), .ZN(n11464) );
  NAND2_X1 U13332 ( .A1(n15637), .A2(n11464), .ZN(n11465) );
  XNOR2_X1 U13333 ( .A(n11682), .B(n11673), .ZN(n11467) );
  NAND2_X1 U13334 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n11467), .ZN(n11675) );
  OAI21_X1 U13335 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n11467), .A(n11675), 
        .ZN(n11468) );
  NAND2_X1 U13336 ( .A1(n11468), .A2(n15667), .ZN(n11470) );
  INV_X1 U13337 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11813) );
  NOR2_X1 U13338 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11813), .ZN(n12248) );
  AOI21_X1 U13339 ( .B1(n15663), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n12248), 
        .ZN(n11469) );
  OAI211_X1 U13340 ( .C1(n15657), .C2(n11674), .A(n11470), .B(n11469), .ZN(
        n11471) );
  AOI21_X1 U13341 ( .B1(n13412), .B2(n11472), .A(n11471), .ZN(n11473) );
  OAI21_X1 U13342 ( .B1(n11474), .B2(n15671), .A(n11473), .ZN(P3_U3193) );
  OR2_X1 U13343 ( .A1(n11486), .A2(n14743), .ZN(n11551) );
  NAND2_X1 U13344 ( .A1(n11556), .A2(n11551), .ZN(n11476) );
  NAND2_X1 U13345 ( .A1(n11476), .A2(n11553), .ZN(n11475) );
  OAI21_X1 U13346 ( .B1(n11476), .B2(n11553), .A(n11475), .ZN(n11477) );
  INV_X1 U13347 ( .A(n11477), .ZN(n11499) );
  OAI211_X1 U13348 ( .C1(n11544), .C2(n11478), .A(n11559), .B(n15796), .ZN(
        n11482) );
  NAND2_X1 U13349 ( .A1(n14741), .A2(n15034), .ZN(n11480) );
  NAND2_X1 U13350 ( .A1(n14743), .A2(n15033), .ZN(n11479) );
  NAND2_X1 U13351 ( .A1(n11480), .A2(n11479), .ZN(n11511) );
  INV_X1 U13352 ( .A(n11511), .ZN(n11481) );
  NAND2_X1 U13353 ( .A1(n11482), .A2(n11481), .ZN(n11496) );
  AOI21_X1 U13354 ( .B1(n16014), .B2(n11550), .A(n11496), .ZN(n11489) );
  NAND2_X1 U13355 ( .A1(n11486), .A2(n11485), .ZN(n11483) );
  OR2_X1 U13356 ( .A1(n11486), .A2(n11485), .ZN(n11487) );
  XNOR2_X1 U13357 ( .A(n11543), .B(n11553), .ZN(n11488) );
  NAND2_X1 U13358 ( .A1(n11488), .A2(n15985), .ZN(n11494) );
  OAI211_X1 U13359 ( .C1(n11499), .C2(n15799), .A(n11489), .B(n11494), .ZN(
        n11491) );
  NAND2_X1 U13360 ( .A1(n11491), .A2(n15922), .ZN(n11490) );
  OAI21_X1 U13361 ( .B1(n15922), .B2(n10067), .A(n11490), .ZN(P1_U3538) );
  NAND2_X1 U13362 ( .A1(n11491), .A2(n15961), .ZN(n11492) );
  OAI21_X1 U13363 ( .B1(n15961), .B2(n9146), .A(n11492), .ZN(P1_U3489) );
  INV_X1 U13364 ( .A(n15025), .ZN(n14920) );
  MUX2_X1 U13365 ( .A(n11494), .B(n11493), .S(n15036), .Z(n11498) );
  OAI22_X1 U13366 ( .A1(n11544), .A2(n15680), .B1(n11508), .B2(n15035), .ZN(
        n11495) );
  AOI21_X1 U13367 ( .B1(n11496), .B2(n14917), .A(n11495), .ZN(n11497) );
  OAI211_X1 U13368 ( .C1(n14920), .C2(n11499), .A(n11498), .B(n11497), .ZN(
        P1_U3283) );
  NAND2_X1 U13369 ( .A1(n11550), .A2(n14614), .ZN(n11503) );
  NAND2_X1 U13370 ( .A1(n14742), .A2(n14659), .ZN(n11502) );
  NAND2_X1 U13371 ( .A1(n11503), .A2(n11502), .ZN(n11504) );
  XNOR2_X1 U13372 ( .A(n11504), .B(n14584), .ZN(n11931) );
  AND2_X1 U13373 ( .A1(n14742), .A2(n14607), .ZN(n11505) );
  AOI21_X1 U13374 ( .B1(n11550), .B2(n14659), .A(n11505), .ZN(n11933) );
  XNOR2_X1 U13375 ( .A(n11931), .B(n11933), .ZN(n11506) );
  OAI211_X1 U13376 ( .C1(n11507), .C2(n11506), .A(n11932), .B(n16036), .ZN(
        n11513) );
  NOR2_X1 U13377 ( .A1(n16041), .A2(n11508), .ZN(n11509) );
  AOI211_X1 U13378 ( .C1(n14691), .C2(n11511), .A(n11510), .B(n11509), .ZN(
        n11512) );
  OAI211_X1 U13379 ( .C1(n11544), .C2(n16033), .A(n11513), .B(n11512), .ZN(
        P1_U3217) );
  NAND2_X1 U13380 ( .A1(n11514), .A2(n12959), .ZN(n11516) );
  AOI22_X1 U13381 ( .A1(n12336), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n12335), 
        .B2(n15422), .ZN(n11515) );
  INV_X1 U13382 ( .A(n14014), .ZN(n12859) );
  NAND2_X1 U13383 ( .A1(n12857), .A2(n12859), .ZN(n11617) );
  OR2_X1 U13384 ( .A1(n12857), .A2(n12859), .ZN(n11517) );
  NAND2_X1 U13385 ( .A1(n12851), .A2(n14015), .ZN(n11518) );
  XOR2_X1 U13386 ( .A(n13008), .B(n11607), .Z(n11534) );
  NAND2_X1 U13387 ( .A1(n12064), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11526) );
  NAND2_X1 U13388 ( .A1(n12468), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11525) );
  INV_X1 U13389 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11520) );
  NAND2_X1 U13390 ( .A1(n11521), .A2(n11520), .ZN(n11522) );
  AND2_X1 U13391 ( .A1(n11972), .A2(n11522), .ZN(n12103) );
  NAND2_X1 U13392 ( .A1(n12425), .A2(n12103), .ZN(n11524) );
  NAND2_X1 U13393 ( .A1(n7508), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n11523) );
  NAND4_X1 U13394 ( .A1(n11526), .A2(n11525), .A3(n11524), .A4(n11523), .ZN(
        n14013) );
  AOI22_X1 U13395 ( .A1(n14242), .A2(n14015), .B1(n14262), .B2(n14013), .ZN(
        n11533) );
  NAND2_X1 U13396 ( .A1(n12851), .A2(n11963), .ZN(n11527) );
  INV_X1 U13397 ( .A(n11618), .ZN(n11531) );
  INV_X1 U13398 ( .A(n13008), .ZN(n11528) );
  AND3_X1 U13399 ( .A1(n11529), .A2(n11528), .A3(n11527), .ZN(n11530) );
  OAI21_X1 U13400 ( .B1(n11531), .B2(n11530), .A(n14267), .ZN(n11532) );
  OAI211_X1 U13401 ( .C1(n11534), .C2(n15778), .A(n11533), .B(n11532), .ZN(
        n15947) );
  INV_X1 U13402 ( .A(n15947), .ZN(n11541) );
  INV_X1 U13403 ( .A(n11534), .ZN(n15949) );
  INV_X1 U13404 ( .A(n11535), .ZN(n11536) );
  INV_X1 U13405 ( .A(n12857), .ZN(n15946) );
  OAI211_X1 U13406 ( .C1(n11536), .C2(n15946), .A(n11286), .B(n11623), .ZN(
        n15945) );
  AOI22_X1 U13407 ( .A1(n15829), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11966), 
        .B2(n15816), .ZN(n11538) );
  NAND2_X1 U13408 ( .A1(n12857), .A2(n15818), .ZN(n11537) );
  OAI211_X1 U13409 ( .C1(n15945), .C2(n14234), .A(n11538), .B(n11537), .ZN(
        n11539) );
  AOI21_X1 U13410 ( .B1(n15949), .B2(n15824), .A(n11539), .ZN(n11540) );
  OAI21_X1 U13411 ( .B1(n11541), .B2(n15817), .A(n11540), .ZN(P2_U3253) );
  NAND2_X1 U13412 ( .A1(n11543), .A2(n11542), .ZN(n11546) );
  NAND2_X1 U13413 ( .A1(n11544), .A2(n14742), .ZN(n11545) );
  NAND2_X1 U13414 ( .A1(n11546), .A2(n11545), .ZN(n11650) );
  XNOR2_X1 U13415 ( .A(n11650), .B(n7994), .ZN(n11547) );
  NAND2_X1 U13416 ( .A1(n11547), .A2(n15985), .ZN(n11549) );
  AOI22_X1 U13417 ( .A1(n15033), .A2(n14742), .B1(n14740), .B2(n15034), .ZN(
        n11548) );
  NAND2_X1 U13418 ( .A1(n11549), .A2(n11548), .ZN(n15920) );
  INV_X1 U13419 ( .A(n15920), .ZN(n11565) );
  OR2_X1 U13420 ( .A1(n11550), .A2(n14742), .ZN(n11552) );
  AND2_X1 U13421 ( .A1(n11551), .A2(n11552), .ZN(n11555) );
  INV_X1 U13422 ( .A(n11552), .ZN(n11554) );
  INV_X1 U13423 ( .A(n11645), .ZN(n11557) );
  AOI21_X1 U13424 ( .B1(n11649), .B2(n11558), .A(n11557), .ZN(n15921) );
  NAND2_X1 U13425 ( .A1(n15917), .A2(n11559), .ZN(n11560) );
  NAND2_X1 U13426 ( .A1(n11659), .A2(n11560), .ZN(n15918) );
  AOI22_X1 U13427 ( .A1(n15020), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n11939), 
        .B2(n15678), .ZN(n11562) );
  NAND2_X1 U13428 ( .A1(n15917), .A2(n15061), .ZN(n11561) );
  OAI211_X1 U13429 ( .C1(n15918), .C2(n15681), .A(n11562), .B(n11561), .ZN(
        n11563) );
  AOI21_X1 U13430 ( .B1(n15921), .B2(n15048), .A(n11563), .ZN(n11564) );
  OAI21_X1 U13431 ( .B1(n15036), .B2(n11565), .A(n11564), .ZN(P1_U3282) );
  XNOR2_X1 U13432 ( .A(n12851), .B(n7532), .ZN(n11954) );
  NAND2_X1 U13433 ( .A1(n14015), .A2(n14295), .ZN(n11952) );
  XNOR2_X1 U13434 ( .A(n11954), .B(n11952), .ZN(n11956) );
  XNOR2_X1 U13435 ( .A(n11957), .B(n11956), .ZN(n11574) );
  INV_X1 U13436 ( .A(n11568), .ZN(n11570) );
  OAI22_X1 U13437 ( .A1(n13995), .A2(n11570), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11569), .ZN(n11572) );
  OAI22_X1 U13438 ( .A1(n12846), .A2(n13997), .B1(n13998), .B2(n12859), .ZN(
        n11571) );
  AOI211_X1 U13439 ( .C1(n12851), .C2(n14001), .A(n11572), .B(n11571), .ZN(
        n11573) );
  OAI21_X1 U13440 ( .B1(n11574), .B2(n14003), .A(n11573), .ZN(P2_U3208) );
  XNOR2_X1 U13441 ( .A(n7543), .B(n15854), .ZN(n12004) );
  XNOR2_X1 U13442 ( .A(n12004), .B(n12009), .ZN(n12006) );
  XNOR2_X1 U13443 ( .A(n12007), .B(n12006), .ZN(n11582) );
  NOR2_X1 U13444 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11890), .ZN(n15620) );
  OAI22_X1 U13445 ( .A1(n11996), .A2(n13237), .B1(n12163), .B2(n13225), .ZN(
        n11579) );
  AOI211_X1 U13446 ( .C1(n15854), .C2(n13206), .A(n15620), .B(n11579), .ZN(
        n11581) );
  NAND2_X1 U13447 ( .A1(n13239), .A2(n11999), .ZN(n11580) );
  OAI211_X1 U13448 ( .C1(n11582), .C2(n13229), .A(n11581), .B(n11580), .ZN(
        P3_U3161) );
  INV_X1 U13449 ( .A(n12334), .ZN(n11584) );
  OAI222_X1 U13450 ( .A1(n15210), .A2(n11583), .B1(n15215), .B2(n11584), .C1(
        P1_U3086), .C2(n14825), .ZN(P1_U3336) );
  OAI222_X1 U13451 ( .A1(n14509), .A2(n11585), .B1(n14506), .B2(n11584), .C1(
        n14073), .C2(P2_U3088), .ZN(P2_U3308) );
  NAND2_X1 U13452 ( .A1(n11589), .A2(n15433), .ZN(n11590) );
  INV_X1 U13453 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15995) );
  NAND2_X1 U13454 ( .A1(n15429), .A2(n15995), .ZN(n15428) );
  NAND2_X1 U13455 ( .A1(n11590), .A2(n15428), .ZN(n11593) );
  INV_X1 U13456 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n16022) );
  NOR2_X1 U13457 ( .A1(n12112), .A2(n16022), .ZN(n11591) );
  AOI21_X1 U13458 ( .B1(n12112), .B2(n16022), .A(n11591), .ZN(n11592) );
  NOR2_X1 U13459 ( .A1(n11592), .A2(n11593), .ZN(n12111) );
  AOI211_X1 U13460 ( .C1(n11593), .C2(n11592), .A(n12111), .B(n14823), .ZN(
        n11605) );
  AOI21_X1 U13461 ( .B1(n11595), .B2(P1_REG2_REG_14__SCAN_IN), .A(n11594), 
        .ZN(n11596) );
  XNOR2_X1 U13462 ( .A(n11596), .B(n15433), .ZN(n15431) );
  NOR2_X1 U13463 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n15431), .ZN(n15430) );
  AOI21_X1 U13464 ( .B1(n11596), .B2(n15433), .A(n15430), .ZN(n11599) );
  NAND2_X1 U13465 ( .A1(n12112), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n12107) );
  INV_X1 U13466 ( .A(n12107), .ZN(n11597) );
  AOI21_X1 U13467 ( .B1(n15056), .B2(n11603), .A(n11597), .ZN(n11598) );
  NAND2_X1 U13468 ( .A1(n11598), .A2(n11599), .ZN(n12106) );
  OAI211_X1 U13469 ( .C1(n11599), .C2(n11598), .A(n14819), .B(n12106), .ZN(
        n11602) );
  NAND2_X1 U13470 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n16006)
         );
  INV_X1 U13471 ( .A(n16006), .ZN(n11600) );
  AOI21_X1 U13472 ( .B1(n14791), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11600), 
        .ZN(n11601) );
  OAI211_X1 U13473 ( .C1(n15432), .C2(n11603), .A(n11602), .B(n11601), .ZN(
        n11604) );
  OR2_X1 U13474 ( .A1(n11605), .A2(n11604), .ZN(P1_U3259) );
  OR2_X1 U13475 ( .A1(n12857), .A2(n14014), .ZN(n11606) );
  NAND2_X1 U13476 ( .A1(n12857), .A2(n14014), .ZN(n11608) );
  OR2_X1 U13477 ( .A1(n11609), .A2(n10521), .ZN(n11611) );
  AOI22_X1 U13478 ( .A1(n12336), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n12335), 
        .B2(n11701), .ZN(n11610) );
  XNOR2_X1 U13479 ( .A(n12865), .B(n14013), .ZN(n13009) );
  XNOR2_X1 U13480 ( .A(n11984), .B(n11616), .ZN(n12145) );
  NAND2_X1 U13481 ( .A1(n12064), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11615) );
  NAND2_X1 U13482 ( .A1(n12468), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n11614) );
  XNOR2_X1 U13483 ( .A(n11972), .B(P2_REG3_REG_14__SCAN_IN), .ZN(n12220) );
  NAND2_X1 U13484 ( .A1(n12425), .A2(n12220), .ZN(n11613) );
  NAND2_X1 U13485 ( .A1(n7508), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n11612) );
  NAND4_X1 U13486 ( .A1(n11615), .A2(n11614), .A3(n11613), .A4(n11612), .ZN(
        n14012) );
  AOI22_X1 U13487 ( .A1(n14242), .A2(n14014), .B1(n14262), .B2(n14012), .ZN(
        n11622) );
  INV_X1 U13488 ( .A(n11979), .ZN(n11620) );
  AND3_X1 U13489 ( .A1(n11618), .A2(n11616), .A3(n11617), .ZN(n11619) );
  OAI21_X1 U13490 ( .B1(n11620), .B2(n11619), .A(n14309), .ZN(n11621) );
  OAI211_X1 U13491 ( .C1(n12145), .C2(n15778), .A(n11622), .B(n11621), .ZN(
        n12146) );
  NAND2_X1 U13492 ( .A1(n12146), .A2(n14275), .ZN(n11627) );
  AOI211_X1 U13493 ( .C1(n12865), .C2(n11623), .A(n14208), .B(n11985), .ZN(
        n12147) );
  AOI22_X1 U13494 ( .A1(n15829), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12103), 
        .B2(n15816), .ZN(n11624) );
  OAI21_X1 U13495 ( .B1(n12154), .B2(n14301), .A(n11624), .ZN(n11625) );
  AOI21_X1 U13496 ( .B1(n12147), .B2(n15823), .A(n11625), .ZN(n11626) );
  OAI211_X1 U13497 ( .C1(n12145), .C2(n14129), .A(n11627), .B(n11626), .ZN(
        P2_U3252) );
  INV_X1 U13498 ( .A(n11628), .ZN(n11629) );
  OAI222_X1 U13499 ( .A1(P3_U3151), .A2(n11630), .B1(n12036), .B2(n11629), 
        .C1(n11714), .C2(n13810), .ZN(P3_U3269) );
  XNOR2_X1 U13500 ( .A(n11632), .B(n11631), .ZN(n11637) );
  OAI21_X1 U13501 ( .B1(n11634), .B2(n12642), .A(n11633), .ZN(n15833) );
  NAND2_X1 U13502 ( .A1(n15833), .A2(n15937), .ZN(n11636) );
  AOI22_X1 U13503 ( .A1(n13642), .A2(n13255), .B1(n13257), .B2(n13643), .ZN(
        n11635) );
  OAI211_X1 U13504 ( .C1(n15719), .C2(n11637), .A(n11636), .B(n11635), .ZN(
        n15831) );
  INV_X1 U13505 ( .A(n15831), .ZN(n11643) );
  INV_X1 U13506 ( .A(n12002), .ZN(n13558) );
  AOI22_X1 U13507 ( .A1(n13663), .A2(n11639), .B1(n13648), .B2(n11638), .ZN(
        n11640) );
  OAI21_X1 U13508 ( .B1(n15590), .B2(n15735), .A(n11640), .ZN(n11641) );
  AOI21_X1 U13509 ( .B1(n15833), .B2(n13558), .A(n11641), .ZN(n11642) );
  OAI21_X1 U13510 ( .B1(n11643), .B2(n13670), .A(n11642), .ZN(P3_U3226) );
  NAND2_X1 U13511 ( .A1(n15917), .A2(n14741), .ZN(n11644) );
  INV_X1 U13512 ( .A(n11654), .ZN(n12020) );
  AND2_X1 U13513 ( .A1(n11646), .A2(n12020), .ZN(n11647) );
  NAND2_X1 U13514 ( .A1(n15173), .A2(n11648), .ZN(n11658) );
  AOI22_X1 U13515 ( .A1(n15033), .A2(n14741), .B1(n14739), .B2(n15034), .ZN(
        n11657) );
  NAND2_X1 U13516 ( .A1(n11650), .A2(n11649), .ZN(n11653) );
  INV_X1 U13517 ( .A(n14741), .ZN(n11651) );
  OR2_X1 U13518 ( .A1(n15917), .A2(n11651), .ZN(n11652) );
  NAND2_X1 U13519 ( .A1(n11653), .A2(n11652), .ZN(n12021) );
  XNOR2_X1 U13520 ( .A(n12021), .B(n11654), .ZN(n11655) );
  NAND2_X1 U13521 ( .A1(n11655), .A2(n15985), .ZN(n11656) );
  AND2_X1 U13522 ( .A1(n12127), .A2(n11659), .ZN(n11660) );
  OR2_X1 U13523 ( .A1(n11660), .A2(n12017), .ZN(n15171) );
  OAI22_X1 U13524 ( .A1(n15055), .A2(n9181), .B1(n12130), .B2(n15035), .ZN(
        n11661) );
  AOI21_X1 U13525 ( .B1(n12127), .B2(n15061), .A(n11661), .ZN(n11662) );
  OAI21_X1 U13526 ( .B1(n15171), .B2(n15681), .A(n11662), .ZN(n11663) );
  AOI21_X1 U13527 ( .B1(n15173), .B2(n15684), .A(n11663), .ZN(n11664) );
  OAI21_X1 U13528 ( .B1(n15175), .B2(n15036), .A(n11664), .ZN(P1_U3281) );
  INV_X1 U13529 ( .A(n12348), .ZN(n12015) );
  OAI222_X1 U13530 ( .A1(n15210), .A2(n11666), .B1(n15215), .B2(n12015), .C1(
        n11665), .C2(P1_U3086), .ZN(P1_U3335) );
  NOR2_X1 U13531 ( .A1(n11682), .A2(n11667), .ZN(n11669) );
  INV_X1 U13532 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U13533 ( .A1(n13269), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n11670), 
        .B2(n13276), .ZN(n11671) );
  NOR2_X1 U13534 ( .A1(n11672), .A2(n11671), .ZN(n13265) );
  AOI21_X1 U13535 ( .B1(n11672), .B2(n11671), .A(n13265), .ZN(n11694) );
  NAND2_X1 U13536 ( .A1(n11674), .A2(n11673), .ZN(n11676) );
  INV_X1 U13537 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n11677) );
  MUX2_X1 U13538 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n11677), .S(n13276), .Z(
        n11678) );
  OAI21_X1 U13539 ( .B1(n11679), .B2(n11678), .A(n13268), .ZN(n11692) );
  NAND2_X1 U13540 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_U3151), .ZN(n12047)
         );
  NAND2_X1 U13541 ( .A1(n15663), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n11680) );
  OAI211_X1 U13542 ( .C1(n15657), .C2(n13276), .A(n12047), .B(n11680), .ZN(
        n11691) );
  MUX2_X1 U13543 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13408), .Z(n13277) );
  XNOR2_X1 U13544 ( .A(n13277), .B(n13269), .ZN(n11685) );
  INV_X1 U13545 ( .A(n11681), .ZN(n11683) );
  NAND2_X1 U13546 ( .A1(n11683), .A2(n11682), .ZN(n11686) );
  AND2_X1 U13547 ( .A1(n11685), .A2(n11686), .ZN(n11684) );
  NAND2_X1 U13548 ( .A1(n11687), .A2(n11684), .ZN(n13281) );
  INV_X1 U13549 ( .A(n13281), .ZN(n11689) );
  AOI21_X1 U13550 ( .B1(n11687), .B2(n11686), .A(n11685), .ZN(n11688) );
  NOR3_X1 U13551 ( .A1(n11689), .A2(n11688), .A3(n15659), .ZN(n11690) );
  AOI211_X1 U13552 ( .C1(n15667), .C2(n11692), .A(n11691), .B(n11690), .ZN(
        n11693) );
  OAI21_X1 U13553 ( .B1(n11694), .B2(n15671), .A(n11693), .ZN(P3_U3194) );
  INV_X1 U13554 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n11707) );
  INV_X1 U13555 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n15969) );
  NOR2_X1 U13556 ( .A1(n14027), .A2(n15969), .ZN(n11696) );
  AOI21_X1 U13557 ( .B1(n14027), .B2(n15969), .A(n11696), .ZN(n11697) );
  AOI211_X1 U13558 ( .C1(n11698), .C2(n11697), .A(n14026), .B(n15387), .ZN(
        n11699) );
  INV_X1 U13559 ( .A(n11699), .ZN(n11706) );
  NAND2_X1 U13560 ( .A1(n14027), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n14038) );
  OAI21_X1 U13561 ( .B1(n14027), .B2(P2_REG2_REG_14__SCAN_IN), .A(n14038), 
        .ZN(n11703) );
  OAI21_X1 U13562 ( .B1(n14039), .B2(n11703), .A(n15423), .ZN(n11702) );
  AOI21_X1 U13563 ( .B1(n14039), .B2(n11703), .A(n11702), .ZN(n11704) );
  AND2_X1 U13564 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n12219) );
  AOI211_X1 U13565 ( .C1(n15421), .C2(n14027), .A(n11704), .B(n12219), .ZN(
        n11705) );
  OAI211_X1 U13566 ( .C1(n15427), .C2(n11707), .A(n11706), .B(n11705), .ZN(
        P2_U3228) );
  INV_X1 U13567 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n11811) );
  AOI22_X1 U13568 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(keyinput_121), .B1(
        n11813), .B2(keyinput_122), .ZN(n11708) );
  OAI221_X1 U13569 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_121), .C1(
        n11813), .C2(keyinput_122), .A(n11708), .ZN(n11798) );
  INV_X1 U13570 ( .A(keyinput_120), .ZN(n11796) );
  INV_X1 U13571 ( .A(keyinput_119), .ZN(n11794) );
  INV_X1 U13572 ( .A(keyinput_115), .ZN(n11785) );
  INV_X1 U13573 ( .A(keyinput_114), .ZN(n11783) );
  OAI22_X1 U13574 ( .A1(n11892), .A2(keyinput_109), .B1(keyinput_108), .B2(
        P3_REG3_REG_1__SCAN_IN), .ZN(n11709) );
  AOI221_X1 U13575 ( .B1(n11892), .B2(keyinput_109), .C1(
        P3_REG3_REG_1__SCAN_IN), .C2(keyinput_108), .A(n11709), .ZN(n11776) );
  INV_X1 U13576 ( .A(keyinput_107), .ZN(n11774) );
  INV_X1 U13577 ( .A(keyinput_106), .ZN(n11772) );
  INV_X1 U13578 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n11886) );
  XOR2_X1 U13579 ( .A(P3_REG3_REG_14__SCAN_IN), .B(keyinput_101), .Z(n11770)
         );
  INV_X1 U13580 ( .A(keyinput_84), .ZN(n11743) );
  INV_X1 U13581 ( .A(keyinput_83), .ZN(n11741) );
  OAI22_X1 U13582 ( .A1(n11711), .A2(keyinput_81), .B1(n11818), .B2(
        keyinput_82), .ZN(n11710) );
  AOI221_X1 U13583 ( .B1(n11711), .B2(keyinput_81), .C1(keyinput_82), .C2(
        n11818), .A(n11710), .ZN(n11738) );
  INV_X1 U13584 ( .A(keyinput_79), .ZN(n11736) );
  OAI22_X1 U13585 ( .A1(n11714), .A2(keyinput_70), .B1(n11713), .B2(
        keyinput_71), .ZN(n11712) );
  AOI221_X1 U13586 ( .B1(n11714), .B2(keyinput_70), .C1(keyinput_71), .C2(
        n11713), .A(n11712), .ZN(n11726) );
  INV_X1 U13587 ( .A(keyinput_69), .ZN(n11721) );
  INV_X1 U13588 ( .A(SI_30_), .ZN(n13807) );
  OAI22_X1 U13589 ( .A1(n13807), .A2(keyinput_66), .B1(keyinput_67), .B2(
        SI_29_), .ZN(n11715) );
  AOI221_X1 U13590 ( .B1(n13807), .B2(keyinput_66), .C1(SI_29_), .C2(
        keyinput_67), .A(n11715), .ZN(n11718) );
  AOI22_X1 U13591 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput_64), .B1(SI_31_), 
        .B2(keyinput_65), .ZN(n11716) );
  OAI221_X1 U13592 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput_64), .C1(SI_31_), 
        .C2(keyinput_65), .A(n11716), .ZN(n11717) );
  AOI22_X1 U13593 ( .A1(n11718), .A2(n11717), .B1(keyinput_68), .B2(SI_28_), 
        .ZN(n11719) );
  OAI21_X1 U13594 ( .B1(keyinput_68), .B2(SI_28_), .A(n11719), .ZN(n11720) );
  OAI221_X1 U13595 ( .B1(SI_27_), .B2(keyinput_69), .C1(n12031), .C2(n11721), 
        .A(n11720), .ZN(n11725) );
  AOI22_X1 U13596 ( .A1(n11723), .A2(keyinput_73), .B1(n11828), .B2(
        keyinput_72), .ZN(n11722) );
  OAI221_X1 U13597 ( .B1(n11723), .B2(keyinput_73), .C1(n11828), .C2(
        keyinput_72), .A(n11722), .ZN(n11724) );
  AOI21_X1 U13598 ( .B1(n11726), .B2(n11725), .A(n11724), .ZN(n11734) );
  XNOR2_X1 U13599 ( .A(SI_22_), .B(keyinput_74), .ZN(n11733) );
  INV_X1 U13600 ( .A(SI_20_), .ZN(n11729) );
  OAI22_X1 U13601 ( .A1(n11729), .A2(keyinput_76), .B1(n11728), .B2(
        keyinput_77), .ZN(n11727) );
  AOI221_X1 U13602 ( .B1(n11729), .B2(keyinput_76), .C1(keyinput_77), .C2(
        n11728), .A(n11727), .ZN(n11732) );
  OAI22_X1 U13603 ( .A1(SI_21_), .A2(keyinput_75), .B1(SI_18_), .B2(
        keyinput_78), .ZN(n11730) );
  AOI221_X1 U13604 ( .B1(SI_21_), .B2(keyinput_75), .C1(keyinput_78), .C2(
        SI_18_), .A(n11730), .ZN(n11731) );
  OAI211_X1 U13605 ( .C1(n11734), .C2(n11733), .A(n11732), .B(n11731), .ZN(
        n11735) );
  OAI221_X1 U13606 ( .B1(SI_17_), .B2(keyinput_79), .C1(n11840), .C2(n11736), 
        .A(n11735), .ZN(n11737) );
  OAI211_X1 U13607 ( .C1(SI_16_), .C2(keyinput_80), .A(n11738), .B(n11737), 
        .ZN(n11739) );
  AOI21_X1 U13608 ( .B1(SI_16_), .B2(keyinput_80), .A(n11739), .ZN(n11740) );
  AOI221_X1 U13609 ( .B1(SI_13_), .B2(keyinput_83), .C1(n11848), .C2(n11741), 
        .A(n11740), .ZN(n11742) );
  AOI221_X1 U13610 ( .B1(SI_12_), .B2(keyinput_84), .C1(n11850), .C2(n11743), 
        .A(n11742), .ZN(n11746) );
  XOR2_X1 U13611 ( .A(SI_10_), .B(keyinput_86), .Z(n11745) );
  XNOR2_X1 U13612 ( .A(SI_11_), .B(keyinput_85), .ZN(n11744) );
  NOR3_X1 U13613 ( .A1(n11746), .A2(n11745), .A3(n11744), .ZN(n11754) );
  XOR2_X1 U13614 ( .A(SI_9_), .B(keyinput_87), .Z(n11753) );
  AOI22_X1 U13615 ( .A1(SI_6_), .A2(keyinput_90), .B1(SI_7_), .B2(keyinput_89), 
        .ZN(n11747) );
  OAI221_X1 U13616 ( .B1(SI_6_), .B2(keyinput_90), .C1(SI_7_), .C2(keyinput_89), .A(n11747), .ZN(n11751) );
  XOR2_X1 U13617 ( .A(SI_5_), .B(keyinput_91), .Z(n11750) );
  XNOR2_X1 U13618 ( .A(SI_4_), .B(keyinput_92), .ZN(n11749) );
  XNOR2_X1 U13619 ( .A(SI_8_), .B(keyinput_88), .ZN(n11748) );
  NOR4_X1 U13620 ( .A1(n11751), .A2(n11750), .A3(n11749), .A4(n11748), .ZN(
        n11752) );
  OAI21_X1 U13621 ( .B1(n11754), .B2(n11753), .A(n11752), .ZN(n11755) );
  OAI21_X1 U13622 ( .B1(SI_3_), .B2(keyinput_93), .A(n11755), .ZN(n11758) );
  OAI22_X1 U13623 ( .A1(SI_1_), .A2(keyinput_95), .B1(keyinput_96), .B2(SI_0_), 
        .ZN(n11756) );
  AOI221_X1 U13624 ( .B1(SI_1_), .B2(keyinput_95), .C1(SI_0_), .C2(keyinput_96), .A(n11756), .ZN(n11757) );
  OAI221_X1 U13625 ( .B1(n11758), .B2(keyinput_93), .C1(n11758), .C2(SI_3_), 
        .A(n11757), .ZN(n11761) );
  INV_X1 U13626 ( .A(P3_RD_REG_SCAN_IN), .ZN(n15673) );
  AOI22_X1 U13627 ( .A1(keyinput_94), .A2(SI_2_), .B1(n15673), .B2(keyinput_97), .ZN(n11759) );
  OAI221_X1 U13628 ( .B1(keyinput_94), .B2(SI_2_), .C1(n15673), .C2(
        keyinput_97), .A(n11759), .ZN(n11760) );
  OAI22_X1 U13629 ( .A1(P3_STATE_REG_SCAN_IN), .A2(keyinput_98), .B1(n11761), 
        .B2(n11760), .ZN(n11764) );
  OAI22_X1 U13630 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(keyinput_100), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(keyinput_99), .ZN(n11762) );
  AOI221_X1 U13631 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_100), .C1(
        keyinput_99), .C2(P3_REG3_REG_7__SCAN_IN), .A(n11762), .ZN(n11763) );
  OAI221_X1 U13632 ( .B1(n11764), .B2(keyinput_98), .C1(n11764), .C2(
        P3_STATE_REG_SCAN_IN), .A(n11763), .ZN(n11769) );
  INV_X1 U13633 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n11878) );
  OAI22_X1 U13634 ( .A1(n11878), .A2(keyinput_102), .B1(keyinput_103), .B2(
        P3_REG3_REG_10__SCAN_IN), .ZN(n11765) );
  AOI221_X1 U13635 ( .B1(n11878), .B2(keyinput_102), .C1(
        P3_REG3_REG_10__SCAN_IN), .C2(keyinput_103), .A(n11765), .ZN(n11768)
         );
  OAI22_X1 U13636 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(keyinput_105), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(keyinput_104), .ZN(n11766) );
  AOI221_X1 U13637 ( .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_105), .C1(
        keyinput_104), .C2(P3_REG3_REG_3__SCAN_IN), .A(n11766), .ZN(n11767) );
  OAI211_X1 U13638 ( .C1(n11770), .C2(n11769), .A(n11768), .B(n11767), .ZN(
        n11771) );
  OAI221_X1 U13639 ( .B1(P3_REG3_REG_28__SCAN_IN), .B2(n11772), .C1(n11886), 
        .C2(keyinput_106), .A(n11771), .ZN(n11773) );
  OAI221_X1 U13640 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .C1(
        n11890), .C2(n11774), .A(n11773), .ZN(n11775) );
  OAI211_X1 U13641 ( .C1(P3_REG3_REG_12__SCAN_IN), .C2(keyinput_110), .A(
        n11776), .B(n11775), .ZN(n11777) );
  AOI21_X1 U13642 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_110), .A(n11777), .ZN(n11780) );
  AOI22_X1 U13643 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(keyinput_111), .B1(n8428), .B2(keyinput_113), .ZN(n11778) );
  OAI221_X1 U13644 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(keyinput_111), .C1(
        n8428), .C2(keyinput_113), .A(n11778), .ZN(n11779) );
  AOI211_X1 U13645 ( .C1(P3_REG3_REG_16__SCAN_IN), .C2(keyinput_112), .A(
        n11780), .B(n11779), .ZN(n11781) );
  OAI21_X1 U13646 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput_112), .A(n11781), .ZN(n11782) );
  OAI221_X1 U13647 ( .B1(P3_REG3_REG_17__SCAN_IN), .B2(n11783), .C1(n11901), 
        .C2(keyinput_114), .A(n11782), .ZN(n11784) );
  OAI221_X1 U13648 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(n11785), .C1(n13186), 
        .C2(keyinput_115), .A(n11784), .ZN(n11791) );
  XNOR2_X1 U13649 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_118), .ZN(n11790)
         );
  XNOR2_X1 U13650 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput_116), .ZN(n11789)
         );
  INV_X1 U13651 ( .A(keyinput_117), .ZN(n11786) );
  NAND2_X1 U13652 ( .A1(n11787), .A2(n11786), .ZN(n11788) );
  NAND4_X1 U13653 ( .A1(n11791), .A2(n11790), .A3(n11789), .A4(n11788), .ZN(
        n11792) );
  AOI21_X1 U13654 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_117), .A(n11792), 
        .ZN(n11793) );
  AOI221_X1 U13655 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_119), .C1(
        n11913), .C2(n11794), .A(n11793), .ZN(n11795) );
  AOI221_X1 U13656 ( .B1(P3_REG3_REG_13__SCAN_IN), .B2(n11796), .C1(n11915), 
        .C2(keyinput_120), .A(n11795), .ZN(n11797) );
  OAI22_X1 U13657 ( .A1(n11798), .A2(n11797), .B1(keyinput_123), .B2(
        P3_REG3_REG_2__SCAN_IN), .ZN(n11799) );
  AOI21_X1 U13658 ( .B1(keyinput_123), .B2(P3_REG3_REG_2__SCAN_IN), .A(n11799), 
        .ZN(n11804) );
  AOI22_X1 U13659 ( .A1(n11802), .A2(keyinput_125), .B1(n11801), .B2(
        keyinput_124), .ZN(n11800) );
  OAI221_X1 U13660 ( .B1(n11802), .B2(keyinput_125), .C1(n11801), .C2(
        keyinput_124), .A(n11800), .ZN(n11803) );
  AOI211_X1 U13661 ( .C1(n11811), .C2(keyinput_126), .A(n11804), .B(n11803), 
        .ZN(n11805) );
  OAI21_X1 U13662 ( .B1(n11811), .B2(keyinput_126), .A(n11805), .ZN(n11807) );
  AOI21_X1 U13663 ( .B1(keyinput_127), .B2(n11807), .A(keyinput_63), .ZN(
        n11809) );
  INV_X1 U13664 ( .A(keyinput_127), .ZN(n11806) );
  AOI21_X1 U13665 ( .B1(n11807), .B2(n11806), .A(n13234), .ZN(n11808) );
  AOI22_X1 U13666 ( .A1(n13234), .A2(n11809), .B1(keyinput_63), .B2(n11808), 
        .ZN(n11924) );
  OAI22_X1 U13667 ( .A1(n11811), .A2(keyinput_62), .B1(keyinput_60), .B2(
        P3_REG3_REG_18__SCAN_IN), .ZN(n11810) );
  AOI221_X1 U13668 ( .B1(n11811), .B2(keyinput_62), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_60), .A(n11810), .ZN(n11921) );
  OAI22_X1 U13669 ( .A1(n11814), .A2(keyinput_57), .B1(n11813), .B2(
        keyinput_58), .ZN(n11812) );
  AOI221_X1 U13670 ( .B1(n11814), .B2(keyinput_57), .C1(keyinput_58), .C2(
        n11813), .A(n11812), .ZN(n11918) );
  INV_X1 U13671 ( .A(keyinput_56), .ZN(n11916) );
  INV_X1 U13672 ( .A(keyinput_55), .ZN(n11912) );
  INV_X1 U13673 ( .A(keyinput_51), .ZN(n11903) );
  INV_X1 U13674 ( .A(keyinput_50), .ZN(n11900) );
  OAI22_X1 U13675 ( .A1(n11816), .A2(keyinput_48), .B1(keyinput_49), .B2(
        P3_REG3_REG_5__SCAN_IN), .ZN(n11815) );
  AOI221_X1 U13676 ( .B1(n11816), .B2(keyinput_48), .C1(P3_REG3_REG_5__SCAN_IN), .C2(keyinput_49), .A(n11815), .ZN(n11897) );
  INV_X1 U13677 ( .A(keyinput_43), .ZN(n11889) );
  INV_X1 U13678 ( .A(keyinput_42), .ZN(n11887) );
  INV_X1 U13679 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n11874) );
  XOR2_X1 U13680 ( .A(keyinput_34), .B(P3_STATE_REG_SCAN_IN), .Z(n11872) );
  INV_X1 U13681 ( .A(keyinput_20), .ZN(n11851) );
  INV_X1 U13682 ( .A(keyinput_19), .ZN(n11847) );
  OAI22_X1 U13683 ( .A1(n11818), .A2(keyinput_18), .B1(SI_15_), .B2(
        keyinput_17), .ZN(n11817) );
  AOI221_X1 U13684 ( .B1(n11818), .B2(keyinput_18), .C1(keyinput_17), .C2(
        SI_15_), .A(n11817), .ZN(n11843) );
  INV_X1 U13685 ( .A(keyinput_15), .ZN(n11841) );
  OAI22_X1 U13686 ( .A1(SI_26_), .A2(keyinput_6), .B1(keyinput_7), .B2(SI_25_), 
        .ZN(n11819) );
  AOI221_X1 U13687 ( .B1(SI_26_), .B2(keyinput_6), .C1(SI_25_), .C2(keyinput_7), .A(n11819), .ZN(n11831) );
  INV_X1 U13688 ( .A(keyinput_5), .ZN(n11826) );
  OAI22_X1 U13689 ( .A1(SI_29_), .A2(keyinput_3), .B1(SI_30_), .B2(keyinput_2), 
        .ZN(n11820) );
  AOI221_X1 U13690 ( .B1(SI_29_), .B2(keyinput_3), .C1(keyinput_2), .C2(SI_30_), .A(n11820), .ZN(n11823) );
  AOI22_X1 U13691 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput_0), .B1(SI_31_), .B2(
        keyinput_1), .ZN(n11821) );
  OAI221_X1 U13692 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput_0), .C1(SI_31_), 
        .C2(keyinput_1), .A(n11821), .ZN(n11822) );
  AOI22_X1 U13693 ( .A1(n11823), .A2(n11822), .B1(keyinput_4), .B2(SI_28_), 
        .ZN(n11824) );
  OAI21_X1 U13694 ( .B1(keyinput_4), .B2(SI_28_), .A(n11824), .ZN(n11825) );
  OAI221_X1 U13695 ( .B1(SI_27_), .B2(keyinput_5), .C1(n12031), .C2(n11826), 
        .A(n11825), .ZN(n11830) );
  AOI22_X1 U13696 ( .A1(SI_23_), .A2(keyinput_9), .B1(n11828), .B2(keyinput_8), 
        .ZN(n11827) );
  OAI221_X1 U13697 ( .B1(SI_23_), .B2(keyinput_9), .C1(n11828), .C2(keyinput_8), .A(n11827), .ZN(n11829) );
  AOI21_X1 U13698 ( .B1(n11831), .B2(n11830), .A(n11829), .ZN(n11838) );
  XNOR2_X1 U13699 ( .A(SI_22_), .B(keyinput_10), .ZN(n11837) );
  OAI22_X1 U13700 ( .A1(n11833), .A2(keyinput_14), .B1(keyinput_11), .B2(
        SI_21_), .ZN(n11832) );
  AOI221_X1 U13701 ( .B1(n11833), .B2(keyinput_14), .C1(SI_21_), .C2(
        keyinput_11), .A(n11832), .ZN(n11836) );
  OAI22_X1 U13702 ( .A1(SI_20_), .A2(keyinput_12), .B1(keyinput_13), .B2(
        SI_19_), .ZN(n11834) );
  AOI221_X1 U13703 ( .B1(SI_20_), .B2(keyinput_12), .C1(SI_19_), .C2(
        keyinput_13), .A(n11834), .ZN(n11835) );
  OAI211_X1 U13704 ( .C1(n11838), .C2(n11837), .A(n11836), .B(n11835), .ZN(
        n11839) );
  OAI221_X1 U13705 ( .B1(SI_17_), .B2(n11841), .C1(n11840), .C2(keyinput_15), 
        .A(n11839), .ZN(n11842) );
  OAI211_X1 U13706 ( .C1(n11845), .C2(keyinput_16), .A(n11843), .B(n11842), 
        .ZN(n11844) );
  AOI21_X1 U13707 ( .B1(n11845), .B2(keyinput_16), .A(n11844), .ZN(n11846) );
  AOI221_X1 U13708 ( .B1(SI_13_), .B2(keyinput_19), .C1(n11848), .C2(n11847), 
        .A(n11846), .ZN(n11849) );
  AOI221_X1 U13709 ( .B1(SI_12_), .B2(n11851), .C1(n11850), .C2(keyinput_20), 
        .A(n11849), .ZN(n11854) );
  XOR2_X1 U13710 ( .A(SI_10_), .B(keyinput_22), .Z(n11853) );
  XNOR2_X1 U13711 ( .A(SI_11_), .B(keyinput_21), .ZN(n11852) );
  NOR3_X1 U13712 ( .A1(n11854), .A2(n11853), .A3(n11852), .ZN(n11863) );
  XOR2_X1 U13713 ( .A(SI_9_), .B(keyinput_23), .Z(n11862) );
  AOI22_X1 U13714 ( .A1(SI_4_), .A2(keyinput_28), .B1(SI_8_), .B2(keyinput_24), 
        .ZN(n11855) );
  OAI221_X1 U13715 ( .B1(SI_4_), .B2(keyinput_28), .C1(SI_8_), .C2(keyinput_24), .A(n11855), .ZN(n11858) );
  AOI22_X1 U13716 ( .A1(SI_6_), .A2(keyinput_26), .B1(SI_7_), .B2(keyinput_25), 
        .ZN(n11856) );
  OAI221_X1 U13717 ( .B1(SI_6_), .B2(keyinput_26), .C1(SI_7_), .C2(keyinput_25), .A(n11856), .ZN(n11857) );
  AOI211_X1 U13718 ( .C1(keyinput_27), .C2(SI_5_), .A(n11858), .B(n11857), 
        .ZN(n11859) );
  OAI21_X1 U13719 ( .B1(keyinput_27), .B2(SI_5_), .A(n11859), .ZN(n11860) );
  INV_X1 U13720 ( .A(n11860), .ZN(n11861) );
  OAI21_X1 U13721 ( .B1(n11863), .B2(n11862), .A(n11861), .ZN(n11870) );
  XNOR2_X1 U13722 ( .A(SI_3_), .B(keyinput_29), .ZN(n11869) );
  XOR2_X1 U13723 ( .A(keyinput_33), .B(n15673), .Z(n11867) );
  XNOR2_X1 U13724 ( .A(SI_0_), .B(keyinput_32), .ZN(n11866) );
  XNOR2_X1 U13725 ( .A(SI_1_), .B(keyinput_31), .ZN(n11865) );
  XNOR2_X1 U13726 ( .A(SI_2_), .B(keyinput_30), .ZN(n11864) );
  NAND4_X1 U13727 ( .A1(n11867), .A2(n11866), .A3(n11865), .A4(n11864), .ZN(
        n11868) );
  AOI21_X1 U13728 ( .B1(n11870), .B2(n11869), .A(n11868), .ZN(n11871) );
  OAI22_X1 U13729 ( .A1(n11872), .A2(n11871), .B1(n11874), .B2(keyinput_36), 
        .ZN(n11873) );
  AOI21_X1 U13730 ( .B1(n11874), .B2(keyinput_36), .A(n11873), .ZN(n11884) );
  OAI22_X1 U13731 ( .A1(n11876), .A2(keyinput_35), .B1(keyinput_37), .B2(
        P3_REG3_REG_14__SCAN_IN), .ZN(n11875) );
  AOI221_X1 U13732 ( .B1(n11876), .B2(keyinput_35), .C1(
        P3_REG3_REG_14__SCAN_IN), .C2(keyinput_37), .A(n11875), .ZN(n11883) );
  INV_X1 U13733 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U13734 ( .A1(n11878), .A2(keyinput_38), .B1(keyinput_39), .B2(
        n12162), .ZN(n11877) );
  OAI221_X1 U13735 ( .B1(n11878), .B2(keyinput_38), .C1(n12162), .C2(
        keyinput_39), .A(n11877), .ZN(n11882) );
  AOI22_X1 U13736 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(keyinput_41), .B1(n11880), .B2(keyinput_40), .ZN(n11879) );
  OAI221_X1 U13737 ( .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_41), .C1(
        n11880), .C2(keyinput_40), .A(n11879), .ZN(n11881) );
  AOI211_X1 U13738 ( .C1(n11884), .C2(n11883), .A(n11882), .B(n11881), .ZN(
        n11885) );
  AOI221_X1 U13739 ( .B1(P3_REG3_REG_28__SCAN_IN), .B2(n11887), .C1(n11886), 
        .C2(keyinput_42), .A(n11885), .ZN(n11888) );
  AOI221_X1 U13740 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput_43), .C1(n11890), .C2(n11889), .A(n11888), .ZN(n11894) );
  AOI22_X1 U13741 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_44), .B1(n11892), 
        .B2(keyinput_45), .ZN(n11891) );
  OAI221_X1 U13742 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_44), .C1(n11892), .C2(keyinput_45), .A(n11891), .ZN(n11893) );
  AOI211_X1 U13743 ( .C1(P3_REG3_REG_12__SCAN_IN), .C2(keyinput_46), .A(n11894), .B(n11893), .ZN(n11895) );
  OAI21_X1 U13744 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_46), .A(n11895), 
        .ZN(n11896) );
  OAI211_X1 U13745 ( .C1(P3_REG3_REG_25__SCAN_IN), .C2(keyinput_47), .A(n11897), .B(n11896), .ZN(n11898) );
  AOI21_X1 U13746 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(keyinput_47), .A(n11898), 
        .ZN(n11899) );
  AOI221_X1 U13747 ( .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput_50), .C1(
        n11901), .C2(n11900), .A(n11899), .ZN(n11902) );
  AOI221_X1 U13748 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .C1(
        n13186), .C2(n11903), .A(n11902), .ZN(n11909) );
  INV_X1 U13749 ( .A(keyinput_52), .ZN(n11904) );
  XNOR2_X1 U13750 ( .A(n11904), .B(P3_REG3_REG_4__SCAN_IN), .ZN(n11907) );
  XNOR2_X1 U13751 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_54), .ZN(n11906)
         );
  NAND2_X1 U13752 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(keyinput_53), .ZN(n11905)
         );
  NAND3_X1 U13753 ( .A1(n11907), .A2(n11906), .A3(n11905), .ZN(n11908) );
  NOR2_X1 U13754 ( .A1(n11909), .A2(n11908), .ZN(n11910) );
  OAI21_X1 U13755 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_53), .A(n11910), 
        .ZN(n11911) );
  OAI221_X1 U13756 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_55), .C1(
        n11913), .C2(n11912), .A(n11911), .ZN(n11914) );
  OAI221_X1 U13757 ( .B1(P3_REG3_REG_13__SCAN_IN), .B2(n11916), .C1(n11915), 
        .C2(keyinput_56), .A(n11914), .ZN(n11917) );
  AOI22_X1 U13758 ( .A1(n11918), .A2(n11917), .B1(keyinput_59), .B2(
        P3_REG3_REG_2__SCAN_IN), .ZN(n11919) );
  OAI21_X1 U13759 ( .B1(keyinput_59), .B2(P3_REG3_REG_2__SCAN_IN), .A(n11919), 
        .ZN(n11920) );
  OAI211_X1 U13760 ( .C1(P3_REG3_REG_6__SCAN_IN), .C2(keyinput_61), .A(n11921), 
        .B(n11920), .ZN(n11922) );
  AOI21_X1 U13761 ( .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_61), .A(n11922), 
        .ZN(n11923) );
  NOR2_X1 U13762 ( .A1(n11924), .A2(n11923), .ZN(n11929) );
  OAI21_X1 U13763 ( .B1(n11925), .B2(P2_IR_REG_15__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n11926) );
  XNOR2_X1 U13764 ( .A(n11926), .B(P2_IR_REG_16__SCAN_IN), .ZN(n14056) );
  AOI222_X1 U13765 ( .A1(n12170), .A2(n14500), .B1(n14056), .B2(
        P2_STATE_REG_SCAN_IN), .C1(P1_DATAO_REG_16__SCAN_IN), .C2(n11927), 
        .ZN(n11928) );
  XNOR2_X1 U13766 ( .A(n11929), .B(n11928), .ZN(P2_U3311) );
  AOI22_X1 U13767 ( .A1(n15917), .A2(n14614), .B1(n14659), .B2(n14741), .ZN(
        n11930) );
  XNOR2_X1 U13768 ( .A(n11930), .B(n14584), .ZN(n12122) );
  AOI22_X1 U13769 ( .A1(n15917), .A2(n14659), .B1(n14607), .B2(n14741), .ZN(
        n12123) );
  XNOR2_X1 U13770 ( .A(n12122), .B(n12123), .ZN(n11935) );
  AOI21_X1 U13771 ( .B1(n11935), .B2(n11934), .A(n12121), .ZN(n11942) );
  INV_X1 U13772 ( .A(n16041), .ZN(n14722) );
  NAND2_X1 U13773 ( .A1(n16029), .A2(n14742), .ZN(n11937) );
  OAI211_X1 U13774 ( .C1(n12124), .C2(n14728), .A(n11937), .B(n11936), .ZN(
        n11938) );
  AOI21_X1 U13775 ( .B1(n11939), .B2(n14722), .A(n11938), .ZN(n11941) );
  NAND2_X1 U13776 ( .A1(n15917), .A2(n14731), .ZN(n11940) );
  OAI211_X1 U13777 ( .C1(n11942), .C2(n14733), .A(n11941), .B(n11940), .ZN(
        P1_U3236) );
  INV_X1 U13778 ( .A(n12656), .ZN(n11943) );
  OR2_X1 U13779 ( .A1(n11943), .A2(n12654), .ZN(n11948) );
  XNOR2_X1 U13780 ( .A(n11944), .B(n11948), .ZN(n11945) );
  AOI222_X1 U13781 ( .A1(n13640), .A2(n11945), .B1(n13254), .B2(n13642), .C1(
        n13255), .C2(n13643), .ZN(n15869) );
  INV_X1 U13782 ( .A(n12011), .ZN(n11946) );
  OAI22_X1 U13783 ( .A1(n13650), .A2(n15870), .B1(n11946), .B2(n15727), .ZN(
        n11947) );
  AOI21_X1 U13784 ( .B1(n13670), .B2(P3_REG2_REG_9__SCAN_IN), .A(n11947), .ZN(
        n11951) );
  INV_X1 U13785 ( .A(n11948), .ZN(n12652) );
  XNOR2_X1 U13786 ( .A(n11949), .B(n12652), .ZN(n15872) );
  NAND2_X1 U13787 ( .A1(n15872), .A2(n13667), .ZN(n11950) );
  OAI211_X1 U13788 ( .C1(n15869), .C2(n13670), .A(n11951), .B(n11950), .ZN(
        P3_U3224) );
  INV_X1 U13789 ( .A(n11952), .ZN(n11953) );
  AND2_X1 U13790 ( .A1(n14014), .A2(n12208), .ZN(n11959) );
  XNOR2_X1 U13791 ( .A(n12857), .B(n7532), .ZN(n11958) );
  NOR2_X1 U13792 ( .A1(n11958), .A2(n11959), .ZN(n12093) );
  AOI21_X1 U13793 ( .B1(n11959), .B2(n11958), .A(n12093), .ZN(n11960) );
  OAI21_X1 U13794 ( .B1(n11961), .B2(n11960), .A(n12095), .ZN(n11962) );
  NAND2_X1 U13795 ( .A1(n11962), .A2(n13966), .ZN(n11968) );
  NAND2_X1 U13796 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n15425)
         );
  INV_X1 U13797 ( .A(n15425), .ZN(n11965) );
  INV_X1 U13798 ( .A(n14013), .ZN(n12217) );
  OAI22_X1 U13799 ( .A1(n11963), .A2(n13997), .B1(n13998), .B2(n12217), .ZN(
        n11964) );
  AOI211_X1 U13800 ( .C1(n11966), .C2(n13971), .A(n11965), .B(n11964), .ZN(
        n11967) );
  OAI211_X1 U13801 ( .C1(n15946), .C2(n13974), .A(n11968), .B(n11967), .ZN(
        P2_U3196) );
  NAND2_X1 U13802 ( .A1(n12468), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n11977) );
  NAND2_X1 U13803 ( .A1(n12064), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n11976) );
  INV_X1 U13804 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11970) );
  INV_X1 U13805 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11969) );
  OAI21_X1 U13806 ( .B1(n11972), .B2(n11970), .A(n11969), .ZN(n11973) );
  NAND2_X1 U13807 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .ZN(n11971) );
  AND2_X1 U13808 ( .A1(n11973), .A2(n12061), .ZN(n12258) );
  NAND2_X1 U13809 ( .A1(n12425), .A2(n12258), .ZN(n11975) );
  NAND2_X1 U13810 ( .A1(n7508), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n11974) );
  NAND4_X1 U13811 ( .A1(n11977), .A2(n11976), .A3(n11975), .A4(n11974), .ZN(
        n14011) );
  INV_X1 U13812 ( .A(n14011), .ZN(n12879) );
  NAND2_X1 U13813 ( .A1(n12865), .A2(n12217), .ZN(n11978) );
  NAND2_X1 U13814 ( .A1(n11980), .A2(n12959), .ZN(n11982) );
  AOI22_X1 U13815 ( .A1(n12336), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n12335), 
        .B2(n14027), .ZN(n11981) );
  INV_X1 U13816 ( .A(n14012), .ZN(n12100) );
  XNOR2_X1 U13817 ( .A(n12873), .B(n12100), .ZN(n13011) );
  XNOR2_X1 U13818 ( .A(n12054), .B(n13011), .ZN(n11983) );
  OAI222_X1 U13819 ( .A1(n14285), .A2(n12879), .B1(n14283), .B2(n12217), .C1(
        n14289), .C2(n11983), .ZN(n15965) );
  INV_X1 U13820 ( .A(n15965), .ZN(n11990) );
  INV_X1 U13821 ( .A(n13011), .ZN(n12070) );
  XNOR2_X1 U13822 ( .A(n12071), .B(n12070), .ZN(n15967) );
  NAND2_X1 U13823 ( .A1(n15964), .A2(n11985), .ZN(n12076) );
  OAI211_X1 U13824 ( .C1(n15964), .C2(n11985), .A(n11286), .B(n12076), .ZN(
        n15962) );
  AOI22_X1 U13825 ( .A1(n15829), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n12220), 
        .B2(n15816), .ZN(n11987) );
  NAND2_X1 U13826 ( .A1(n12873), .A2(n15818), .ZN(n11986) );
  OAI211_X1 U13827 ( .C1(n15962), .C2(n14234), .A(n11987), .B(n11986), .ZN(
        n11988) );
  AOI21_X1 U13828 ( .B1(n15967), .B2(n14315), .A(n11988), .ZN(n11989) );
  OAI21_X1 U13829 ( .B1(n11990), .B2(n15817), .A(n11989), .ZN(P2_U3251) );
  OAI21_X1 U13830 ( .B1(n11992), .B2(n12647), .A(n11991), .ZN(n15855) );
  INV_X1 U13831 ( .A(n15855), .ZN(n12003) );
  NAND2_X1 U13832 ( .A1(n11993), .A2(n12647), .ZN(n11994) );
  AOI21_X1 U13833 ( .B1(n11995), .B2(n11994), .A(n15719), .ZN(n11998) );
  OAI22_X1 U13834 ( .A1(n11996), .A2(n15721), .B1(n12163), .B2(n15723), .ZN(
        n11997) );
  AOI211_X1 U13835 ( .C1(n15855), .C2(n15937), .A(n11998), .B(n11997), .ZN(
        n15857) );
  MUX2_X1 U13836 ( .A(n11399), .B(n15857), .S(n15735), .Z(n12001) );
  AOI22_X1 U13837 ( .A1(n13663), .A2(n15854), .B1(n13648), .B2(n11999), .ZN(
        n12000) );
  OAI211_X1 U13838 ( .C1(n12003), .C2(n12002), .A(n12001), .B(n12000), .ZN(
        P3_U3225) );
  INV_X1 U13839 ( .A(n12004), .ZN(n12005) );
  XNOR2_X1 U13840 ( .A(n13109), .B(n15870), .ZN(n12037) );
  INV_X1 U13841 ( .A(n12037), .ZN(n12039) );
  XNOR2_X1 U13842 ( .A(n12039), .B(n12163), .ZN(n12008) );
  NOR2_X1 U13843 ( .A1(n7341), .A2(n12008), .ZN(n12159) );
  AOI21_X1 U13844 ( .B1(n7341), .B2(n12008), .A(n12159), .ZN(n12014) );
  AND2_X1 U13845 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n15640) );
  OAI22_X1 U13846 ( .A1(n12246), .A2(n13225), .B1(n12009), .B2(n13237), .ZN(
        n12010) );
  AOI211_X1 U13847 ( .C1(n7905), .C2(n13206), .A(n15640), .B(n12010), .ZN(
        n12013) );
  NAND2_X1 U13848 ( .A1(n13239), .A2(n12011), .ZN(n12012) );
  OAI211_X1 U13849 ( .C1(n12014), .C2(n13229), .A(n12013), .B(n12012), .ZN(
        P3_U3171) );
  OAI222_X1 U13850 ( .A1(n14509), .A2(n12349), .B1(P2_U3088), .B2(n10408), 
        .C1(n14506), .C2(n12015), .ZN(P2_U3307) );
  AOI21_X1 U13851 ( .B1(n12016), .B2(n12230), .A(n12224), .ZN(n15953) );
  OAI22_X1 U13852 ( .A1(n15055), .A2(n9218), .B1(n12272), .B2(n15035), .ZN(
        n12019) );
  OAI21_X1 U13853 ( .B1(n15955), .B2(n12017), .A(n12280), .ZN(n15956) );
  NOR2_X1 U13854 ( .A1(n15956), .A2(n15681), .ZN(n12018) );
  AOI211_X1 U13855 ( .C1(n15061), .C2(n12269), .A(n12019), .B(n12018), .ZN(
        n12029) );
  NAND2_X1 U13856 ( .A1(n12021), .A2(n12020), .ZN(n12023) );
  OR2_X1 U13857 ( .A1(n12127), .A2(n12124), .ZN(n12022) );
  NAND2_X1 U13858 ( .A1(n12023), .A2(n12022), .ZN(n12231) );
  INV_X1 U13859 ( .A(n12230), .ZN(n12024) );
  XNOR2_X1 U13860 ( .A(n12231), .B(n12024), .ZN(n12025) );
  NAND2_X1 U13861 ( .A1(n12025), .A2(n15985), .ZN(n12027) );
  AOI22_X1 U13862 ( .A1(n15033), .A2(n14740), .B1(n15978), .B2(n15034), .ZN(
        n12026) );
  NAND2_X1 U13863 ( .A1(n12027), .A2(n12026), .ZN(n15958) );
  NAND2_X1 U13864 ( .A1(n15958), .A2(n15055), .ZN(n12028) );
  OAI211_X1 U13865 ( .C1(n15953), .C2(n14988), .A(n12029), .B(n12028), .ZN(
        P1_U3280) );
  INV_X1 U13866 ( .A(n12030), .ZN(n12032) );
  OAI222_X1 U13867 ( .A1(P3_U3151), .A2(n13408), .B1(n12036), .B2(n12032), 
        .C1(n12031), .C2(n13810), .ZN(P3_U3268) );
  INV_X1 U13868 ( .A(n12033), .ZN(n12035) );
  XNOR2_X1 U13869 ( .A(n12664), .B(n13109), .ZN(n12245) );
  XNOR2_X1 U13870 ( .A(n15892), .B(n13109), .ZN(n12156) );
  NOR2_X1 U13871 ( .A1(n12156), .A2(n12246), .ZN(n12242) );
  AOI21_X1 U13872 ( .B1(n7907), .B2(n12037), .A(n12242), .ZN(n12038) );
  NAND2_X1 U13873 ( .A1(n12039), .A2(n12163), .ZN(n12155) );
  NAND2_X1 U13874 ( .A1(n12156), .A2(n12246), .ZN(n12040) );
  OAI211_X1 U13875 ( .C1(n12242), .C2(n12155), .A(n12245), .B(n12040), .ZN(
        n12041) );
  OAI21_X1 U13876 ( .B1(n12164), .B2(n12245), .A(n12041), .ZN(n12042) );
  XNOR2_X1 U13877 ( .A(n7543), .B(n12316), .ZN(n12043) );
  NOR2_X1 U13878 ( .A1(n12043), .A2(n13252), .ZN(n12082) );
  NAND2_X1 U13879 ( .A1(n12043), .A2(n13252), .ZN(n12083) );
  INV_X1 U13880 ( .A(n12083), .ZN(n12044) );
  NOR2_X1 U13881 ( .A1(n12082), .A2(n12044), .ZN(n12045) );
  XNOR2_X1 U13882 ( .A(n12084), .B(n12045), .ZN(n12046) );
  NAND2_X1 U13883 ( .A1(n12046), .A2(n13221), .ZN(n12051) );
  NOR2_X1 U13884 ( .A1(n12164), .A2(n13237), .ZN(n12049) );
  OAI21_X1 U13885 ( .B1(n12306), .B2(n13225), .A(n12047), .ZN(n12048) );
  AOI211_X1 U13886 ( .C1(n12313), .C2(n13239), .A(n12049), .B(n12048), .ZN(
        n12050) );
  OAI211_X1 U13887 ( .C1(n13242), .C2(n15934), .A(n12051), .B(n12050), .ZN(
        P3_U3164) );
  INV_X1 U13888 ( .A(n12361), .ZN(n12500) );
  OAI222_X1 U13889 ( .A1(n15210), .A2(n12053), .B1(n15215), .B2(n12500), .C1(
        P1_U3086), .C2(n12052), .ZN(P1_U3334) );
  INV_X1 U13890 ( .A(n12058), .ZN(n12059) );
  NAND2_X1 U13891 ( .A1(n12055), .A2(n12959), .ZN(n12057) );
  AOI22_X1 U13892 ( .A1(n12336), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n12335), 
        .B2(n15393), .ZN(n12056) );
  XNOR2_X1 U13893 ( .A(n12877), .B(n14011), .ZN(n13012) );
  INV_X1 U13894 ( .A(n13012), .ZN(n12074) );
  OAI211_X1 U13895 ( .C1(n12059), .C2(n13012), .A(n14309), .B(n12176), .ZN(
        n12069) );
  INV_X1 U13896 ( .A(n12061), .ZN(n12060) );
  NAND2_X1 U13897 ( .A1(n12060), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n12180) );
  INV_X1 U13898 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n14033) );
  NAND2_X1 U13899 ( .A1(n12061), .A2(n14033), .ZN(n12062) );
  NAND2_X1 U13900 ( .A1(n12180), .A2(n12062), .ZN(n13917) );
  INV_X1 U13901 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n12063) );
  OAI22_X1 U13902 ( .A1(n13917), .A2(n12458), .B1(n12471), .B2(n12063), .ZN(
        n12068) );
  INV_X1 U13903 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n12065) );
  INV_X1 U13904 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12189) );
  OAI22_X1 U13905 ( .A1(n12066), .A2(n12065), .B1(n10460), .B2(n12189), .ZN(
        n12067) );
  AOI22_X1 U13906 ( .A1(n14242), .A2(n14012), .B1(n14262), .B2(n14010), .ZN(
        n12256) );
  NAND2_X1 U13907 ( .A1(n12069), .A2(n12256), .ZN(n12289) );
  INV_X1 U13908 ( .A(n12289), .ZN(n12081) );
  OR2_X1 U13909 ( .A1(n12873), .A2(n14012), .ZN(n12072) );
  NAND2_X1 U13910 ( .A1(n12073), .A2(n12072), .ZN(n12075) );
  NAND2_X1 U13911 ( .A1(n12075), .A2(n12074), .ZN(n12196) );
  OAI21_X1 U13912 ( .B1(n12075), .B2(n12074), .A(n12196), .ZN(n12291) );
  INV_X1 U13913 ( .A(n12877), .ZN(n12296) );
  AOI211_X1 U13914 ( .C1(n12877), .C2(n12076), .A(n14295), .B(n12190), .ZN(
        n12290) );
  NAND2_X1 U13915 ( .A1(n12290), .A2(n15823), .ZN(n12078) );
  AOI22_X1 U13916 ( .A1(n15829), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n12258), 
        .B2(n15816), .ZN(n12077) );
  OAI211_X1 U13917 ( .C1(n12296), .C2(n14301), .A(n12078), .B(n12077), .ZN(
        n12079) );
  AOI21_X1 U13918 ( .B1(n14315), .B2(n12291), .A(n12079), .ZN(n12080) );
  OAI21_X1 U13919 ( .B1(n15817), .B2(n12081), .A(n12080), .ZN(P2_U3250) );
  XNOR2_X1 U13920 ( .A(n13665), .B(n13109), .ZN(n12297) );
  OAI211_X1 U13921 ( .C1(n12085), .C2(n12297), .A(n12300), .B(n13221), .ZN(
        n12090) );
  NAND2_X1 U13922 ( .A1(P3_REG3_REG_13__SCAN_IN), .A2(P3_U3151), .ZN(n13272)
         );
  NAND2_X1 U13923 ( .A1(n13252), .A2(n13223), .ZN(n12086) );
  OAI211_X1 U13924 ( .C1(n13656), .C2(n13225), .A(n13272), .B(n12086), .ZN(
        n12088) );
  NOR2_X1 U13925 ( .A1(n13742), .A2(n13242), .ZN(n12087) );
  AOI211_X1 U13926 ( .C1(n13660), .C2(n13239), .A(n12088), .B(n12087), .ZN(
        n12089) );
  NAND2_X1 U13927 ( .A1(n12090), .A2(n12089), .ZN(P3_U3174) );
  AND2_X1 U13928 ( .A1(n14013), .A2(n14295), .ZN(n12092) );
  XNOR2_X1 U13929 ( .A(n12865), .B(n7532), .ZN(n12091) );
  NOR2_X1 U13930 ( .A1(n12091), .A2(n12092), .ZN(n12211) );
  AOI21_X1 U13931 ( .B1(n12092), .B2(n12091), .A(n12211), .ZN(n12097) );
  INV_X1 U13932 ( .A(n12093), .ZN(n12094) );
  OAI21_X1 U13933 ( .B1(n12097), .B2(n12096), .A(n12213), .ZN(n12098) );
  NAND2_X1 U13934 ( .A1(n12098), .A2(n13966), .ZN(n12105) );
  INV_X1 U13935 ( .A(n12099), .ZN(n12102) );
  OAI22_X1 U13936 ( .A1(n12859), .A2(n13997), .B1(n13998), .B2(n12100), .ZN(
        n12101) );
  AOI211_X1 U13937 ( .C1(n12103), .C2(n13971), .A(n12102), .B(n12101), .ZN(
        n12104) );
  OAI211_X1 U13938 ( .C1(n12154), .C2(n13974), .A(n12105), .B(n12104), .ZN(
        P2_U3206) );
  NAND2_X1 U13939 ( .A1(n12107), .A2(n12106), .ZN(n12110) );
  NOR2_X1 U13940 ( .A1(n14803), .A2(n15032), .ZN(n12108) );
  AOI21_X1 U13941 ( .B1(n15032), .B2(n14803), .A(n12108), .ZN(n12109) );
  NAND2_X1 U13942 ( .A1(n12109), .A2(n12110), .ZN(n14802) );
  OAI211_X1 U13943 ( .C1(n12110), .C2(n12109), .A(n14819), .B(n14802), .ZN(
        n12120) );
  AOI21_X1 U13944 ( .B1(n12112), .B2(P1_REG1_REG_16__SCAN_IN), .A(n12111), 
        .ZN(n12114) );
  XNOR2_X1 U13945 ( .A(n14797), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n12113) );
  NOR2_X1 U13946 ( .A1(n12114), .A2(n12113), .ZN(n14796) );
  AOI211_X1 U13947 ( .C1(n12114), .C2(n12113), .A(n14796), .B(n14823), .ZN(
        n12118) );
  NAND2_X1 U13948 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3086), .ZN(n16038)
         );
  INV_X1 U13949 ( .A(n16038), .ZN(n12115) );
  AOI21_X1 U13950 ( .B1(n14791), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n12115), 
        .ZN(n12116) );
  OAI21_X1 U13951 ( .B1(n15432), .B2(n14803), .A(n12116), .ZN(n12117) );
  NOR2_X1 U13952 ( .A1(n12118), .A2(n12117), .ZN(n12119) );
  NAND2_X1 U13953 ( .A1(n12120), .A2(n12119), .ZN(P1_U3260) );
  OAI22_X1 U13954 ( .A1(n15170), .A2(n14583), .B1(n12124), .B2(n14582), .ZN(
        n12125) );
  XNOR2_X1 U13955 ( .A(n12125), .B(n14584), .ZN(n12262) );
  AND2_X1 U13956 ( .A1(n14740), .A2(n14607), .ZN(n12126) );
  AOI21_X1 U13957 ( .B1(n12127), .B2(n14659), .A(n12126), .ZN(n12263) );
  XNOR2_X1 U13958 ( .A(n12262), .B(n12263), .ZN(n12128) );
  OAI211_X1 U13959 ( .C1(n12129), .C2(n12128), .A(n12265), .B(n16036), .ZN(
        n12134) );
  NOR2_X1 U13960 ( .A1(n16041), .A2(n12130), .ZN(n12132) );
  INV_X1 U13961 ( .A(n14739), .ZN(n12266) );
  OAI22_X1 U13962 ( .A1(n14728), .A2(n12266), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9175), .ZN(n12131) );
  AOI211_X1 U13963 ( .C1(n16029), .C2(n14741), .A(n12132), .B(n12131), .ZN(
        n12133) );
  OAI211_X1 U13964 ( .C1(n15170), .C2(n16033), .A(n12134), .B(n12133), .ZN(
        P1_U3224) );
  AOI21_X1 U13965 ( .B1(n12135), .B2(n12658), .A(n15719), .ZN(n12138) );
  OAI22_X1 U13966 ( .A1(n12164), .A2(n15723), .B1(n12163), .B2(n15721), .ZN(
        n12136) );
  AOI21_X1 U13967 ( .B1(n12138), .B2(n12137), .A(n12136), .ZN(n15894) );
  XNOR2_X1 U13968 ( .A(n12139), .B(n12658), .ZN(n15896) );
  INV_X1 U13969 ( .A(n15896), .ZN(n15898) );
  NAND2_X1 U13970 ( .A1(n15898), .A2(n13667), .ZN(n12144) );
  INV_X1 U13971 ( .A(n15892), .ZN(n12141) );
  INV_X1 U13972 ( .A(n12140), .ZN(n12168) );
  OAI22_X1 U13973 ( .A1(n13650), .A2(n12141), .B1(n12168), .B2(n15727), .ZN(
        n12142) );
  AOI21_X1 U13974 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n13670), .A(n12142), 
        .ZN(n12143) );
  OAI211_X1 U13975 ( .C1(n13670), .C2(n15894), .A(n12144), .B(n12143), .ZN(
        P3_U3223) );
  INV_X1 U13976 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n12149) );
  INV_X1 U13977 ( .A(n12145), .ZN(n12148) );
  AOI211_X1 U13978 ( .C1(n15950), .C2(n12148), .A(n12147), .B(n12146), .ZN(
        n12151) );
  MUX2_X1 U13979 ( .A(n12149), .B(n12151), .S(n15974), .Z(n12150) );
  OAI21_X1 U13980 ( .B1(n12154), .B2(n14467), .A(n12150), .ZN(P2_U3469) );
  MUX2_X1 U13981 ( .A(n12152), .B(n12151), .S(n15970), .Z(n12153) );
  OAI21_X1 U13982 ( .B1(n12154), .B2(n14417), .A(n12153), .ZN(P2_U3512) );
  INV_X1 U13983 ( .A(n12155), .ZN(n12158) );
  XNOR2_X1 U13984 ( .A(n12156), .B(n12246), .ZN(n12157) );
  NOR3_X1 U13985 ( .A1(n12159), .A2(n12158), .A3(n12157), .ZN(n12243) );
  INV_X1 U13986 ( .A(n12243), .ZN(n12161) );
  OAI21_X1 U13987 ( .B1(n12159), .B2(n12158), .A(n12157), .ZN(n12160) );
  NAND3_X1 U13988 ( .A1(n12161), .A2(n13221), .A3(n12160), .ZN(n12167) );
  NOR2_X1 U13989 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12162), .ZN(n15662) );
  OAI22_X1 U13990 ( .A1(n12164), .A2(n13225), .B1(n12163), .B2(n13237), .ZN(
        n12165) );
  AOI211_X1 U13991 ( .C1(n15892), .C2(n13206), .A(n15662), .B(n12165), .ZN(
        n12166) );
  OAI211_X1 U13992 ( .C1(n12169), .C2(n12168), .A(n12167), .B(n12166), .ZN(
        P3_U3157) );
  NAND2_X1 U13993 ( .A1(n12170), .A2(n12959), .ZN(n12172) );
  AOI22_X1 U13994 ( .A1(n12336), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n12335), 
        .B2(n14056), .ZN(n12171) );
  INV_X1 U13995 ( .A(n14010), .ZN(n12173) );
  OR2_X1 U13996 ( .A1(n14471), .A2(n12173), .ZN(n14305) );
  NAND2_X1 U13997 ( .A1(n14471), .A2(n12173), .ZN(n12174) );
  OR2_X1 U13998 ( .A1(n12877), .A2(n12879), .ZN(n12175) );
  OAI211_X1 U13999 ( .C1(n13014), .C2(n12177), .A(n14307), .B(n14267), .ZN(
        n12188) );
  INV_X1 U14000 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14465) );
  INV_X1 U14001 ( .A(n12180), .ZN(n12178) );
  NAND2_X1 U14002 ( .A1(n12178), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n12327) );
  INV_X1 U14003 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n12179) );
  NAND2_X1 U14004 ( .A1(n12180), .A2(n12179), .ZN(n12181) );
  NAND2_X1 U14005 ( .A1(n12327), .A2(n12181), .ZN(n14317) );
  OR2_X1 U14006 ( .A1(n14317), .A2(n12458), .ZN(n12185) );
  NAND2_X1 U14007 ( .A1(n12064), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n12183) );
  NAND2_X1 U14008 ( .A1(n12468), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n12182) );
  AND2_X1 U14009 ( .A1(n12183), .A2(n12182), .ZN(n12184) );
  OAI211_X1 U14010 ( .C1(n12471), .C2(n14465), .A(n12185), .B(n12184), .ZN(
        n14009) );
  NAND2_X1 U14011 ( .A1(n14009), .A2(n14262), .ZN(n12187) );
  NAND2_X1 U14012 ( .A1(n14242), .A2(n14011), .ZN(n12186) );
  AND2_X1 U14013 ( .A1(n12187), .A2(n12186), .ZN(n13918) );
  OAI22_X1 U14014 ( .A1(n14275), .A2(n12189), .B1(n13917), .B2(n14318), .ZN(
        n12195) );
  INV_X1 U14015 ( .A(n14471), .ZN(n12191) );
  AOI21_X1 U14016 ( .B1(n14471), .B2(n12192), .A(n14295), .ZN(n12193) );
  NAND2_X1 U14017 ( .A1(n14321), .A2(n12193), .ZN(n14418) );
  NOR2_X1 U14018 ( .A1(n14418), .A2(n14234), .ZN(n12194) );
  AOI211_X1 U14019 ( .C1(n15818), .C2(n14471), .A(n12195), .B(n12194), .ZN(
        n12200) );
  INV_X1 U14020 ( .A(n13014), .ZN(n12197) );
  OAI21_X1 U14021 ( .B1(n12198), .B2(n12197), .A(n12480), .ZN(n14420) );
  OR2_X1 U14022 ( .A1(n14420), .A2(n14254), .ZN(n12199) );
  OAI211_X1 U14023 ( .C1(n14419), .C2(n15817), .A(n12200), .B(n12199), .ZN(
        P2_U3249) );
  XNOR2_X1 U14024 ( .A(n12201), .B(n12664), .ZN(n12202) );
  AOI222_X1 U14025 ( .A1(n13640), .A2(n12202), .B1(n13254), .B2(n13643), .C1(
        n13252), .C2(n13642), .ZN(n15909) );
  INV_X1 U14026 ( .A(n12249), .ZN(n12203) );
  OAI22_X1 U14027 ( .A1(n13650), .A2(n15910), .B1(n12203), .B2(n15727), .ZN(
        n12204) );
  AOI21_X1 U14028 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n13670), .A(n12204), 
        .ZN(n12207) );
  XNOR2_X1 U14029 ( .A(n12205), .B(n12664), .ZN(n15913) );
  NAND2_X1 U14030 ( .A1(n15913), .A2(n13667), .ZN(n12206) );
  OAI211_X1 U14031 ( .C1(n15909), .C2(n13670), .A(n12207), .B(n12206), .ZN(
        P3_U3222) );
  AND2_X1 U14032 ( .A1(n14012), .A2(n14208), .ZN(n12210) );
  XNOR2_X1 U14033 ( .A(n12873), .B(n7532), .ZN(n12209) );
  NOR2_X1 U14034 ( .A1(n12209), .A2(n12210), .ZN(n12253) );
  AOI21_X1 U14035 ( .B1(n12210), .B2(n12209), .A(n12253), .ZN(n12215) );
  INV_X1 U14036 ( .A(n12211), .ZN(n12212) );
  OAI21_X1 U14037 ( .B1(n12215), .B2(n12214), .A(n12255), .ZN(n12216) );
  NAND2_X1 U14038 ( .A1(n12216), .A2(n13966), .ZN(n12222) );
  OAI22_X1 U14039 ( .A1(n12217), .A2(n13997), .B1(n13998), .B2(n12879), .ZN(
        n12218) );
  AOI211_X1 U14040 ( .C1(n12220), .C2(n13971), .A(n12219), .B(n12218), .ZN(
        n12221) );
  OAI211_X1 U14041 ( .C1(n15964), .C2(n13974), .A(n12222), .B(n12221), .ZN(
        P2_U3187) );
  XNOR2_X1 U14042 ( .A(n12517), .B(n12236), .ZN(n15994) );
  INV_X1 U14043 ( .A(n15994), .ZN(n12241) );
  INV_X1 U14044 ( .A(n16028), .ZN(n14532) );
  OAI22_X1 U14045 ( .A1(n14520), .A2(n15049), .B1(n14532), .B2(n15051), .ZN(
        n15988) );
  INV_X1 U14046 ( .A(n15984), .ZN(n12225) );
  AOI22_X1 U14047 ( .A1(n15988), .A2(n15055), .B1(n12225), .B2(n15678), .ZN(
        n12226) );
  OAI21_X1 U14048 ( .B1(n12227), .B2(n15055), .A(n12226), .ZN(n12229) );
  OAI21_X1 U14049 ( .B1(n7715), .B2(n7352), .A(n7717), .ZN(n15992) );
  NOR2_X1 U14050 ( .A1(n15992), .A2(n15681), .ZN(n12228) );
  AOI211_X1 U14051 ( .C1(n15061), .C2(n15989), .A(n12229), .B(n12228), .ZN(
        n12240) );
  NAND2_X1 U14052 ( .A1(n12231), .A2(n12230), .ZN(n12233) );
  OR2_X1 U14053 ( .A1(n12269), .A2(n12266), .ZN(n12232) );
  NOR2_X1 U14054 ( .A1(n15165), .A2(n14520), .ZN(n12234) );
  NAND2_X1 U14055 ( .A1(n15165), .A2(n14520), .ZN(n12235) );
  NAND2_X1 U14056 ( .A1(n12238), .A2(n12237), .ZN(n15986) );
  INV_X1 U14057 ( .A(n15064), .ZN(n14985) );
  NAND3_X1 U14058 ( .A1(n15987), .A2(n15986), .A3(n14985), .ZN(n12239) );
  OAI211_X1 U14059 ( .C1(n12241), .C2(n14988), .A(n12240), .B(n12239), .ZN(
        P1_U3278) );
  NOR2_X1 U14060 ( .A1(n12243), .A2(n12242), .ZN(n12244) );
  XOR2_X1 U14061 ( .A(n12245), .B(n12244), .Z(n12252) );
  INV_X1 U14062 ( .A(n13225), .ZN(n13235) );
  OAI22_X1 U14063 ( .A1(n12246), .A2(n13237), .B1(n13242), .B2(n15910), .ZN(
        n12247) );
  AOI211_X1 U14064 ( .C1(n13235), .C2(n13252), .A(n12248), .B(n12247), .ZN(
        n12251) );
  NAND2_X1 U14065 ( .A1(n13239), .A2(n12249), .ZN(n12250) );
  OAI211_X1 U14066 ( .C1(n12252), .C2(n13229), .A(n12251), .B(n12250), .ZN(
        P3_U3176) );
  INV_X1 U14067 ( .A(n12253), .ZN(n12254) );
  NAND2_X1 U14068 ( .A1(n14011), .A2(n12208), .ZN(n13816) );
  XOR2_X1 U14069 ( .A(n13816), .B(n13815), .Z(n13818) );
  XNOR2_X1 U14070 ( .A(n13819), .B(n13818), .ZN(n12261) );
  AND2_X1 U14071 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n15392) );
  NOR2_X1 U14072 ( .A1(n13939), .A2(n12256), .ZN(n12257) );
  AOI211_X1 U14073 ( .C1(n13971), .C2(n12258), .A(n15392), .B(n12257), .ZN(
        n12260) );
  NAND2_X1 U14074 ( .A1(n12877), .A2(n14001), .ZN(n12259) );
  OAI211_X1 U14075 ( .C1(n12261), .C2(n14003), .A(n12260), .B(n12259), .ZN(
        P2_U3213) );
  INV_X1 U14076 ( .A(n12262), .ZN(n12264) );
  NAND2_X1 U14077 ( .A1(n12265), .A2(n8256), .ZN(n12271) );
  OAI22_X1 U14078 ( .A1(n15955), .A2(n14583), .B1(n12266), .B2(n14582), .ZN(
        n12267) );
  XNOR2_X1 U14079 ( .A(n12267), .B(n14584), .ZN(n14515) );
  AND2_X1 U14080 ( .A1(n14739), .A2(n14607), .ZN(n12268) );
  AOI21_X1 U14081 ( .B1(n12269), .B2(n14659), .A(n12268), .ZN(n14516) );
  XNOR2_X1 U14082 ( .A(n14515), .B(n14516), .ZN(n12270) );
  OAI211_X1 U14083 ( .C1(n12271), .C2(n12270), .A(n14518), .B(n16036), .ZN(
        n12277) );
  NOR2_X1 U14084 ( .A1(n16041), .A2(n12272), .ZN(n12275) );
  OAI22_X1 U14085 ( .A1(n14728), .A2(n14520), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12273), .ZN(n12274) );
  AOI211_X1 U14086 ( .C1(n16029), .C2(n14740), .A(n12275), .B(n12274), .ZN(
        n12276) );
  OAI211_X1 U14087 ( .C1(n15955), .C2(n16033), .A(n12277), .B(n12276), .ZN(
        P1_U3234) );
  XNOR2_X1 U14088 ( .A(n12278), .B(n12284), .ZN(n12279) );
  AOI222_X1 U14089 ( .A1(n14739), .A2(n15033), .B1(n15985), .B2(n12279), .C1(
        n16000), .C2(n15034), .ZN(n15168) );
  XNOR2_X1 U14090 ( .A(n14521), .B(n12280), .ZN(n15166) );
  INV_X1 U14091 ( .A(n14636), .ZN(n12281) );
  AOI22_X1 U14092 ( .A1(n15020), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n12281), 
        .B2(n15678), .ZN(n12282) );
  OAI21_X1 U14093 ( .B1(n14521), .B2(n15680), .A(n12282), .ZN(n12287) );
  OAI21_X1 U14094 ( .B1(n12285), .B2(n12284), .A(n12283), .ZN(n15169) );
  NOR2_X1 U14095 ( .A1(n15169), .A2(n14988), .ZN(n12286) );
  AOI211_X1 U14096 ( .C1(n15166), .C2(n15018), .A(n12287), .B(n12286), .ZN(
        n12288) );
  OAI21_X1 U14097 ( .B1(n15036), .B2(n15168), .A(n12288), .ZN(P1_U3279) );
  INV_X1 U14098 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n12292) );
  INV_X1 U14099 ( .A(n15847), .ZN(n15968) );
  AOI211_X1 U14100 ( .C1(n15968), .C2(n12291), .A(n12290), .B(n12289), .ZN(
        n12294) );
  MUX2_X1 U14101 ( .A(n12292), .B(n12294), .S(n15974), .Z(n12293) );
  OAI21_X1 U14102 ( .B1(n12296), .B2(n14467), .A(n12293), .ZN(P2_U3475) );
  INV_X1 U14103 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n15389) );
  MUX2_X1 U14104 ( .A(n15389), .B(n12294), .S(n15970), .Z(n12295) );
  OAI21_X1 U14105 ( .B1(n12296), .B2(n14417), .A(n12295), .ZN(P2_U3514) );
  XNOR2_X1 U14106 ( .A(n13793), .B(n13109), .ZN(n13062) );
  XNOR2_X1 U14107 ( .A(n13062), .B(n13627), .ZN(n12304) );
  INV_X1 U14108 ( .A(n12297), .ZN(n12298) );
  NAND2_X1 U14109 ( .A1(n12298), .A2(n13644), .ZN(n12299) );
  INV_X1 U14110 ( .A(n13064), .ZN(n12302) );
  AOI21_X1 U14111 ( .B1(n12304), .B2(n12303), .A(n12302), .ZN(n12310) );
  NAND2_X1 U14112 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(P3_U3151), .ZN(n13298)
         );
  NAND2_X1 U14113 ( .A1(n13235), .A2(n13641), .ZN(n12305) );
  OAI211_X1 U14114 ( .C1(n12306), .C2(n13237), .A(n13298), .B(n12305), .ZN(
        n12308) );
  NOR2_X1 U14115 ( .A1(n13793), .A2(n13242), .ZN(n12307) );
  AOI211_X1 U14116 ( .C1(n13647), .C2(n13239), .A(n12308), .B(n12307), .ZN(
        n12309) );
  OAI21_X1 U14117 ( .B1(n12310), .B2(n13229), .A(n12309), .ZN(P3_U3155) );
  XNOR2_X1 U14118 ( .A(n12311), .B(n12581), .ZN(n12312) );
  AOI222_X1 U14119 ( .A1(n13640), .A2(n12312), .B1(n13644), .B2(n13642), .C1(
        n13253), .C2(n13643), .ZN(n15933) );
  INV_X1 U14120 ( .A(n12313), .ZN(n12314) );
  OAI22_X1 U14121 ( .A1(n15735), .A2(n11670), .B1(n12314), .B2(n15727), .ZN(
        n12315) );
  AOI21_X1 U14122 ( .B1(n12316), .B2(n13663), .A(n12315), .ZN(n12319) );
  XNOR2_X1 U14123 ( .A(n12317), .B(n12581), .ZN(n15938) );
  NAND2_X1 U14124 ( .A1(n15938), .A2(n13667), .ZN(n12318) );
  OAI211_X1 U14125 ( .C1(n15933), .C2(n13670), .A(n12319), .B(n12318), .ZN(
        P3_U3221) );
  NAND2_X1 U14126 ( .A1(n12320), .A2(n12959), .ZN(n12322) );
  AOI22_X1 U14127 ( .A1(n12336), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n12335), 
        .B2(n15404), .ZN(n12321) );
  XNOR2_X1 U14128 ( .A(n14320), .B(n14009), .ZN(n14313) );
  INV_X1 U14129 ( .A(n14009), .ZN(n14284) );
  OR2_X1 U14130 ( .A1(n14320), .A2(n14284), .ZN(n12323) );
  AOI22_X1 U14131 ( .A1(n12336), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n12335), 
        .B2(n14060), .ZN(n12324) );
  NAND2_X1 U14132 ( .A1(n12327), .A2(n12326), .ZN(n12328) );
  NAND2_X1 U14133 ( .A1(n12340), .A2(n12328), .ZN(n14297) );
  AOI22_X1 U14134 ( .A1(n12468), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n12064), 
        .B2(P2_REG2_REG_18__SCAN_IN), .ZN(n12330) );
  NAND2_X1 U14135 ( .A1(n7508), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n12329) );
  OAI211_X1 U14136 ( .C1(n14297), .C2(n12458), .A(n12330), .B(n12329), .ZN(
        n14008) );
  INV_X1 U14137 ( .A(n14008), .ZN(n14265) );
  NAND2_X1 U14138 ( .A1(n14408), .A2(n14265), .ZN(n12331) );
  INV_X1 U14139 ( .A(n14408), .ZN(n14302) );
  NAND2_X1 U14140 ( .A1(n14302), .A2(n14008), .ZN(n12332) );
  NAND2_X1 U14141 ( .A1(n12334), .A2(n12959), .ZN(n12338) );
  AOI22_X1 U14142 ( .A1(n12336), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n12335), 
        .B2(n14078), .ZN(n12337) );
  INV_X1 U14143 ( .A(n12340), .ZN(n12339) );
  NAND2_X1 U14144 ( .A1(n12339), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n12352) );
  INV_X1 U14145 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n14072) );
  NAND2_X1 U14146 ( .A1(n12340), .A2(n14072), .ZN(n12341) );
  NAND2_X1 U14147 ( .A1(n12352), .A2(n12341), .ZN(n14273) );
  OR2_X1 U14148 ( .A1(n14273), .A2(n12458), .ZN(n12346) );
  INV_X1 U14149 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14274) );
  NAND2_X1 U14150 ( .A1(n12468), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n12343) );
  NAND2_X1 U14151 ( .A1(n7508), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n12342) );
  OAI211_X1 U14152 ( .C1(n10460), .C2(n14274), .A(n12343), .B(n12342), .ZN(
        n12344) );
  INV_X1 U14153 ( .A(n12344), .ZN(n12345) );
  NAND2_X1 U14154 ( .A1(n12346), .A2(n12345), .ZN(n14243) );
  XNOR2_X1 U14155 ( .A(n14461), .B(n14243), .ZN(n13016) );
  INV_X1 U14156 ( .A(n14243), .ZN(n14286) );
  NAND2_X1 U14157 ( .A1(n14461), .A2(n14286), .ZN(n12347) );
  NAND2_X1 U14158 ( .A1(n12348), .A2(n12959), .ZN(n12351) );
  OR2_X1 U14159 ( .A1(n12960), .A2(n12349), .ZN(n12350) );
  NAND2_X1 U14160 ( .A1(n12352), .A2(n13968), .ZN(n12353) );
  AND2_X1 U14161 ( .A1(n12365), .A2(n12353), .ZN(n14248) );
  NAND2_X1 U14162 ( .A1(n14248), .A2(n12425), .ZN(n12359) );
  INV_X1 U14163 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n12356) );
  NAND2_X1 U14164 ( .A1(n12468), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n12355) );
  NAND2_X1 U14165 ( .A1(n12064), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n12354) );
  OAI211_X1 U14166 ( .C1(n12356), .C2(n12471), .A(n12355), .B(n12354), .ZN(
        n12357) );
  INV_X1 U14167 ( .A(n12357), .ZN(n12358) );
  NAND2_X1 U14168 ( .A1(n12359), .A2(n12358), .ZN(n14263) );
  XNOR2_X1 U14169 ( .A(n14396), .B(n14263), .ZN(n14240) );
  INV_X1 U14170 ( .A(n14263), .ZN(n14222) );
  NAND2_X1 U14171 ( .A1(n14396), .A2(n14222), .ZN(n12360) );
  NAND2_X1 U14172 ( .A1(n12361), .A2(n12959), .ZN(n12363) );
  OR2_X1 U14173 ( .A1(n12960), .A2(n12501), .ZN(n12362) );
  INV_X1 U14174 ( .A(n12365), .ZN(n12364) );
  NAND2_X1 U14175 ( .A1(n12364), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n12381) );
  INV_X1 U14176 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13900) );
  NAND2_X1 U14177 ( .A1(n12365), .A2(n13900), .ZN(n12366) );
  NAND2_X1 U14178 ( .A1(n12381), .A2(n12366), .ZN(n14231) );
  OR2_X1 U14179 ( .A1(n14231), .A2(n12458), .ZN(n12372) );
  INV_X1 U14180 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n12369) );
  NAND2_X1 U14181 ( .A1(n12468), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n12368) );
  NAND2_X1 U14182 ( .A1(n12064), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n12367) );
  OAI211_X1 U14183 ( .C1(n12369), .C2(n12471), .A(n12368), .B(n12367), .ZN(
        n12370) );
  INV_X1 U14184 ( .A(n12370), .ZN(n12371) );
  NAND2_X1 U14185 ( .A1(n12372), .A2(n12371), .ZN(n14244) );
  INV_X1 U14186 ( .A(n14244), .ZN(n13979) );
  XNOR2_X1 U14187 ( .A(n14456), .B(n13979), .ZN(n14220) );
  OR2_X1 U14188 ( .A1(n14456), .A2(n13979), .ZN(n12373) );
  INV_X1 U14189 ( .A(n12374), .ZN(n12376) );
  NAND2_X1 U14190 ( .A1(n12376), .A2(n12375), .ZN(n12377) );
  NAND2_X1 U14191 ( .A1(n12378), .A2(n12377), .ZN(n14505) );
  OR2_X1 U14192 ( .A1(n12960), .A2(n14508), .ZN(n12379) );
  INV_X1 U14193 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13977) );
  NAND2_X1 U14194 ( .A1(n12381), .A2(n13977), .ZN(n12382) );
  AND2_X1 U14195 ( .A1(n12393), .A2(n12382), .ZN(n14210) );
  NAND2_X1 U14196 ( .A1(n14210), .A2(n12425), .ZN(n12388) );
  INV_X1 U14197 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n12385) );
  NAND2_X1 U14198 ( .A1(n12468), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n12384) );
  NAND2_X1 U14199 ( .A1(n12064), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n12383) );
  OAI211_X1 U14200 ( .C1(n12385), .C2(n12471), .A(n12384), .B(n12383), .ZN(
        n12386) );
  INV_X1 U14201 ( .A(n12386), .ZN(n12387) );
  NAND2_X1 U14202 ( .A1(n15211), .A2(n12959), .ZN(n12390) );
  OR2_X1 U14203 ( .A1(n12960), .A2(n14504), .ZN(n12389) );
  INV_X1 U14204 ( .A(n12393), .ZN(n12391) );
  NAND2_X1 U14205 ( .A1(n12391), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n12405) );
  INV_X1 U14206 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n12392) );
  NAND2_X1 U14207 ( .A1(n12393), .A2(n12392), .ZN(n12394) );
  NAND2_X1 U14208 ( .A1(n12405), .A2(n12394), .ZN(n14197) );
  OR2_X1 U14209 ( .A1(n14197), .A2(n12458), .ZN(n12399) );
  INV_X1 U14210 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n14450) );
  NAND2_X1 U14211 ( .A1(n12468), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n12396) );
  NAND2_X1 U14212 ( .A1(n12064), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n12395) );
  OAI211_X1 U14213 ( .C1(n12471), .C2(n14450), .A(n12396), .B(n12395), .ZN(
        n12397) );
  INV_X1 U14214 ( .A(n12397), .ZN(n12398) );
  NAND2_X1 U14215 ( .A1(n12399), .A2(n12398), .ZN(n14204) );
  INV_X1 U14216 ( .A(n14204), .ZN(n14171) );
  NAND2_X1 U14217 ( .A1(n14497), .A2(n12959), .ZN(n12402) );
  OR2_X1 U14218 ( .A1(n12960), .A2(n14499), .ZN(n12401) );
  INV_X1 U14219 ( .A(n14372), .ZN(n12924) );
  INV_X1 U14220 ( .A(n12405), .ZN(n12403) );
  INV_X1 U14221 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n12404) );
  NAND2_X1 U14222 ( .A1(n12405), .A2(n12404), .ZN(n12406) );
  NAND2_X1 U14223 ( .A1(n12423), .A2(n12406), .ZN(n14178) );
  OR2_X1 U14224 ( .A1(n14178), .A2(n12458), .ZN(n12411) );
  INV_X1 U14225 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n14447) );
  NAND2_X1 U14226 ( .A1(n12468), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n12408) );
  NAND2_X1 U14227 ( .A1(n12064), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n12407) );
  OAI211_X1 U14228 ( .C1(n12471), .C2(n14447), .A(n12408), .B(n12407), .ZN(
        n12409) );
  INV_X1 U14229 ( .A(n12409), .ZN(n12410) );
  XNOR2_X1 U14230 ( .A(n12924), .B(n14006), .ZN(n13021) );
  INV_X1 U14231 ( .A(n13021), .ZN(n14174) );
  OR2_X1 U14232 ( .A1(n14372), .A2(n14006), .ZN(n14147) );
  NAND2_X1 U14233 ( .A1(n14494), .A2(n12959), .ZN(n12413) );
  OR2_X1 U14234 ( .A1(n12960), .A2(n14496), .ZN(n12412) );
  XNOR2_X1 U14235 ( .A(n12423), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n14161) );
  NAND2_X1 U14236 ( .A1(n14161), .A2(n12425), .ZN(n12418) );
  INV_X1 U14237 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14443) );
  NAND2_X1 U14238 ( .A1(n12468), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n12415) );
  NAND2_X1 U14239 ( .A1(n12064), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n12414) );
  OAI211_X1 U14240 ( .C1(n14443), .C2(n12471), .A(n12415), .B(n12414), .ZN(
        n12416) );
  INV_X1 U14241 ( .A(n12416), .ZN(n12417) );
  NAND2_X1 U14242 ( .A1(n12418), .A2(n12417), .ZN(n14169) );
  NAND2_X1 U14243 ( .A1(n14158), .A2(n14134), .ZN(n12420) );
  OR2_X1 U14244 ( .A1(n14158), .A2(n14134), .ZN(n12419) );
  NAND2_X1 U14245 ( .A1(n12420), .A2(n12419), .ZN(n14148) );
  NAND2_X1 U14246 ( .A1(n14491), .A2(n12959), .ZN(n12422) );
  OR2_X1 U14247 ( .A1(n12960), .A2(n14492), .ZN(n12421) );
  INV_X1 U14248 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13907) );
  INV_X1 U14249 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13994) );
  OAI21_X1 U14250 ( .B1(n12423), .B2(n13907), .A(n13994), .ZN(n12424) );
  AND2_X1 U14251 ( .A1(n12424), .A2(n12435), .ZN(n14141) );
  NAND2_X1 U14252 ( .A1(n14141), .A2(n12425), .ZN(n12431) );
  INV_X1 U14253 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n12428) );
  NAND2_X1 U14254 ( .A1(n12468), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n12427) );
  NAND2_X1 U14255 ( .A1(n12064), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n12426) );
  OAI211_X1 U14256 ( .C1(n12428), .C2(n12471), .A(n12427), .B(n12426), .ZN(
        n12429) );
  INV_X1 U14257 ( .A(n12429), .ZN(n12430) );
  NAND2_X1 U14258 ( .A1(n14363), .A2(n14151), .ZN(n14115) );
  OR2_X1 U14259 ( .A1(n14363), .A2(n14151), .ZN(n12432) );
  NAND2_X1 U14260 ( .A1(n12498), .A2(n12959), .ZN(n12434) );
  OR2_X1 U14261 ( .A1(n12960), .A2(n14489), .ZN(n12433) );
  INV_X1 U14262 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13864) );
  NOR2_X1 U14263 ( .A1(n12435), .A2(n13864), .ZN(n12444) );
  INV_X1 U14264 ( .A(n12444), .ZN(n12445) );
  NAND2_X1 U14265 ( .A1(n12435), .A2(n13864), .ZN(n12436) );
  NAND2_X1 U14266 ( .A1(n12445), .A2(n12436), .ZN(n14123) );
  OR2_X1 U14267 ( .A1(n14123), .A2(n12458), .ZN(n12441) );
  INV_X1 U14268 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n14435) );
  NAND2_X1 U14269 ( .A1(n12468), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n12438) );
  NAND2_X1 U14270 ( .A1(n12064), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n12437) );
  OAI211_X1 U14271 ( .C1(n14435), .C2(n12471), .A(n12438), .B(n12437), .ZN(
        n12439) );
  INV_X1 U14272 ( .A(n12439), .ZN(n12440) );
  XNOR2_X1 U14273 ( .A(n14122), .B(n14101), .ZN(n13025) );
  NAND2_X1 U14274 ( .A1(n14483), .A2(n12959), .ZN(n12443) );
  OR2_X1 U14275 ( .A1(n12960), .A2(n14486), .ZN(n12442) );
  NAND2_X1 U14276 ( .A1(n12444), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n12478) );
  INV_X1 U14277 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n13892) );
  NAND2_X1 U14278 ( .A1(n12445), .A2(n13892), .ZN(n12446) );
  NAND2_X1 U14279 ( .A1(n12478), .A2(n12446), .ZN(n14105) );
  INV_X1 U14280 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n12449) );
  NAND2_X1 U14281 ( .A1(n12468), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n12448) );
  NAND2_X1 U14282 ( .A1(n12064), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n12447) );
  OAI211_X1 U14283 ( .C1(n12449), .C2(n12471), .A(n12448), .B(n12447), .ZN(
        n12450) );
  INV_X1 U14284 ( .A(n12450), .ZN(n12451) );
  INV_X1 U14285 ( .A(n14114), .ZN(n13865) );
  NAND2_X1 U14286 ( .A1(n14341), .A2(n13865), .ZN(n12453) );
  OR2_X1 U14287 ( .A1(n14437), .A2(n14101), .ZN(n14096) );
  AND2_X1 U14288 ( .A1(n14094), .A2(n14096), .ZN(n12454) );
  NAND2_X1 U14289 ( .A1(n14480), .A2(n12959), .ZN(n12457) );
  OR2_X1 U14290 ( .A1(n12960), .A2(n14481), .ZN(n12456) );
  OR2_X1 U14291 ( .A1(n12478), .A2(n12458), .ZN(n12464) );
  INV_X1 U14292 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n12461) );
  NAND2_X1 U14293 ( .A1(n12468), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n12460) );
  NAND2_X1 U14294 ( .A1(n12064), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n12459) );
  OAI211_X1 U14295 ( .C1(n12461), .C2(n12471), .A(n12460), .B(n12459), .ZN(
        n12462) );
  INV_X1 U14296 ( .A(n12462), .ZN(n12463) );
  NAND2_X1 U14297 ( .A1(n12464), .A2(n12463), .ZN(n14100) );
  XNOR2_X1 U14298 ( .A(n14337), .B(n14100), .ZN(n13022) );
  NAND2_X1 U14299 ( .A1(n14114), .A2(n14242), .ZN(n12473) );
  OR2_X1 U14300 ( .A1(n14487), .A2(n12466), .ZN(n12467) );
  AND2_X1 U14301 ( .A1(n14262), .A2(n12467), .ZN(n14086) );
  INV_X1 U14302 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14430) );
  NAND2_X1 U14303 ( .A1(n12468), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n12470) );
  NAND2_X1 U14304 ( .A1(n12064), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n12469) );
  OAI211_X1 U14305 ( .C1(n12471), .C2(n14430), .A(n12470), .B(n12469), .ZN(
        n14005) );
  NAND2_X1 U14306 ( .A1(n14086), .A2(n14005), .ZN(n12472) );
  NAND2_X1 U14307 ( .A1(n14302), .A2(n14324), .ZN(n14293) );
  NAND2_X1 U14308 ( .A1(n14196), .A2(n14372), .ZN(n14181) );
  OR2_X2 U14309 ( .A1(n14181), .A2(n14158), .ZN(n14159) );
  AOI21_X1 U14310 ( .B1(n7267), .B2(n14337), .A(n14295), .ZN(n12475) );
  AND2_X1 U14311 ( .A1(n12475), .A2(n7311), .ZN(n14336) );
  NAND2_X1 U14312 ( .A1(n14337), .A2(n15818), .ZN(n12477) );
  NAND2_X1 U14313 ( .A1(n15829), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n12476) );
  OAI211_X1 U14314 ( .C1(n14318), .C2(n12478), .A(n12477), .B(n12476), .ZN(
        n12496) );
  NAND2_X1 U14315 ( .A1(n14471), .A2(n14010), .ZN(n12479) );
  OR2_X1 U14316 ( .A1(n14320), .A2(n14009), .ZN(n12481) );
  NAND2_X1 U14317 ( .A1(n12482), .A2(n12481), .ZN(n14282) );
  XNOR2_X1 U14318 ( .A(n14408), .B(n14265), .ZN(n14288) );
  NAND2_X1 U14319 ( .A1(n14302), .A2(n14265), .ZN(n12483) );
  NAND2_X1 U14320 ( .A1(n14396), .A2(n14263), .ZN(n12484) );
  NAND2_X1 U14321 ( .A1(n14238), .A2(n12484), .ZN(n12486) );
  OR2_X1 U14322 ( .A1(n14396), .A2(n14263), .ZN(n12485) );
  NOR2_X1 U14323 ( .A1(n14456), .A2(n14244), .ZN(n12487) );
  NAND2_X1 U14324 ( .A1(n14456), .A2(n14244), .ZN(n12488) );
  OR2_X1 U14325 ( .A1(n14193), .A2(n14204), .ZN(n12991) );
  NAND2_X1 U14326 ( .A1(n14185), .A2(n12991), .ZN(n12489) );
  NAND2_X1 U14327 ( .A1(n14193), .A2(n14204), .ZN(n12990) );
  NAND2_X1 U14328 ( .A1(n12489), .A2(n12990), .ZN(n14175) );
  OR2_X1 U14329 ( .A1(n14372), .A2(n14188), .ZN(n12490) );
  OR2_X1 U14330 ( .A1(n14158), .A2(n14169), .ZN(n12491) );
  NAND2_X1 U14331 ( .A1(n14157), .A2(n12491), .ZN(n14130) );
  AND2_X1 U14332 ( .A1(n14441), .A2(n14151), .ZN(n12492) );
  OR2_X1 U14333 ( .A1(n14441), .A2(n14151), .ZN(n12493) );
  INV_X1 U14334 ( .A(n13025), .ZN(n14116) );
  INV_X1 U14335 ( .A(n14094), .ZN(n14097) );
  XNOR2_X1 U14336 ( .A(n12494), .B(n13022), .ZN(n14340) );
  NOR2_X1 U14337 ( .A1(n14340), .A2(n14254), .ZN(n12495) );
  OAI21_X1 U14338 ( .B1(n14339), .B2(n15817), .A(n12497), .ZN(P2_U3236) );
  INV_X1 U14339 ( .A(n12498), .ZN(n14488) );
  OAI222_X1 U14340 ( .A1(n15210), .A2(n12499), .B1(n15215), .B2(n14488), .C1(
        P1_U3086), .C2(n12531), .ZN(P1_U3328) );
  OAI222_X1 U14341 ( .A1(n14509), .A2(n12501), .B1(n14506), .B2(n12500), .C1(
        n7526), .C2(P2_U3088), .ZN(P2_U3306) );
  INV_X1 U14342 ( .A(n15107), .ZN(n14912) );
  OR2_X1 U14343 ( .A1(n15989), .A2(n15050), .ZN(n12502) );
  NAND2_X1 U14344 ( .A1(n15987), .A2(n12502), .ZN(n15044) );
  INV_X1 U14345 ( .A(n15044), .ZN(n12504) );
  NAND2_X1 U14346 ( .A1(n12504), .A2(n12503), .ZN(n15042) );
  NAND2_X1 U14347 ( .A1(n16013), .A2(n14532), .ZN(n12505) );
  NAND2_X1 U14348 ( .A1(n15042), .A2(n12505), .ZN(n15028) );
  INV_X1 U14349 ( .A(n16001), .ZN(n15052) );
  AND2_X1 U14350 ( .A1(n16027), .A2(n15052), .ZN(n12506) );
  NAND2_X1 U14351 ( .A1(n15007), .A2(n15006), .ZN(n15005) );
  NAND2_X1 U14352 ( .A1(n15023), .A2(n16030), .ZN(n12507) );
  NAND2_X1 U14353 ( .A1(n15145), .A2(n14719), .ZN(n12508) );
  OR2_X1 U14354 ( .A1(n14562), .A2(n12520), .ZN(n12509) );
  OR2_X1 U14355 ( .A1(n14961), .A2(n14573), .ZN(n12510) );
  INV_X1 U14356 ( .A(n14923), .ZN(n14937) );
  AND2_X1 U14357 ( .A1(n15117), .A2(n12511), .ZN(n12512) );
  INV_X1 U14358 ( .A(n14895), .ZN(n15100) );
  NOR2_X1 U14359 ( .A1(n14884), .A2(n14896), .ZN(n12513) );
  INV_X1 U14360 ( .A(n14896), .ZN(n14870) );
  INV_X1 U14361 ( .A(n14857), .ZN(n14868) );
  INV_X1 U14362 ( .A(n14877), .ZN(n14841) );
  INV_X1 U14363 ( .A(n14737), .ZN(n14871) );
  NAND2_X1 U14364 ( .A1(n14843), .A2(n12514), .ZN(n12516) );
  XNOR2_X1 U14365 ( .A(n12516), .B(n12515), .ZN(n15080) );
  NAND2_X1 U14366 ( .A1(n15047), .A2(n15046), .ZN(n15045) );
  INV_X1 U14367 ( .A(n15006), .ZN(n15012) );
  INV_X1 U14368 ( .A(n14942), .ZN(n14947) );
  INV_X1 U14369 ( .A(n14954), .ZN(n15123) );
  NAND2_X1 U14370 ( .A1(n14954), .A2(n14927), .ZN(n12521) );
  NAND2_X1 U14371 ( .A1(n15117), .A2(n14738), .ZN(n12522) );
  INV_X1 U14372 ( .A(n12525), .ZN(n14846) );
  XNOR2_X1 U14373 ( .A(n12528), .B(n12515), .ZN(n15072) );
  NAND2_X1 U14374 ( .A1(n15072), .A2(n15048), .ZN(n12540) );
  INV_X1 U14375 ( .A(n16013), .ZN(n16003) );
  NAND2_X1 U14376 ( .A1(n15023), .A2(n15014), .ZN(n15017) );
  XNOR2_X1 U14377 ( .A(n14849), .B(n12529), .ZN(n15077) );
  NOR2_X1 U14378 ( .A1(n12531), .A2(n12530), .ZN(n12532) );
  NOR2_X1 U14379 ( .A1(n15051), .A2(n12532), .ZN(n14829) );
  NAND2_X1 U14380 ( .A1(n14735), .A2(n14829), .ZN(n15074) );
  OAI22_X1 U14381 ( .A1(n12534), .A2(n15074), .B1(n12533), .B2(n15035), .ZN(
        n12536) );
  NAND2_X1 U14382 ( .A1(n14737), .A2(n15033), .ZN(n15073) );
  NOR2_X1 U14383 ( .A1(n15036), .A2(n15073), .ZN(n12535) );
  AOI211_X1 U14384 ( .C1(n15020), .C2(P1_REG2_REG_29__SCAN_IN), .A(n12536), 
        .B(n12535), .ZN(n12537) );
  OAI21_X1 U14385 ( .B1(n15075), .B2(n15680), .A(n12537), .ZN(n12538) );
  AOI21_X1 U14386 ( .B1(n15077), .B2(n15018), .A(n12538), .ZN(n12539) );
  OAI211_X1 U14387 ( .C1(n15064), .C2(n15080), .A(n12540), .B(n12539), .ZN(
        P1_U3356) );
  INV_X1 U14388 ( .A(n12541), .ZN(n12542) );
  NAND2_X1 U14389 ( .A1(n12543), .A2(n12542), .ZN(n12545) );
  NAND2_X1 U14390 ( .A1(n15198), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12544) );
  NAND2_X1 U14391 ( .A1(n12545), .A2(n12544), .ZN(n12559) );
  XNOR2_X1 U14392 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n12557) );
  NAND2_X1 U14393 ( .A1(n12559), .A2(n12557), .ZN(n12547) );
  INV_X1 U14394 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13060) );
  NAND2_X1 U14395 ( .A1(n13060), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12546) );
  NAND2_X1 U14396 ( .A1(n12547), .A2(n12546), .ZN(n12549) );
  INV_X1 U14397 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n14479) );
  XNOR2_X1 U14398 ( .A(n14479), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n12548) );
  XNOR2_X1 U14399 ( .A(n12549), .B(n12548), .ZN(n13799) );
  NAND2_X1 U14400 ( .A1(n13799), .A2(n12560), .ZN(n12551) );
  INV_X1 U14401 ( .A(SI_31_), .ZN(n13804) );
  OR2_X1 U14402 ( .A1(n7221), .A2(n13804), .ZN(n12550) );
  NAND2_X1 U14403 ( .A1(n12552), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12555) );
  NAND2_X1 U14404 ( .A1(n8520), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12554) );
  NAND2_X1 U14405 ( .A1(n8759), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12553) );
  INV_X1 U14406 ( .A(n12557), .ZN(n12558) );
  XNOR2_X1 U14407 ( .A(n12559), .B(n12558), .ZN(n13805) );
  NAND2_X1 U14408 ( .A1(n13805), .A2(n12560), .ZN(n12562) );
  OR2_X1 U14409 ( .A1(n7221), .A2(n13807), .ZN(n12561) );
  NAND2_X1 U14410 ( .A1(n12562), .A2(n12561), .ZN(n12566) );
  NAND2_X1 U14411 ( .A1(n12566), .A2(n12565), .ZN(n12563) );
  INV_X1 U14412 ( .A(n13423), .ZN(n13243) );
  NOR2_X1 U14413 ( .A1(n13748), .A2(n13243), .ZN(n12601) );
  INV_X1 U14414 ( .A(n12735), .ZN(n12564) );
  NAND2_X1 U14415 ( .A1(n12612), .A2(n13407), .ZN(n12597) );
  NOR4_X1 U14416 ( .A1(n12600), .A2(n12601), .A3(n12564), .A4(n12597), .ZN(
        n12571) );
  OR2_X1 U14417 ( .A1(n12566), .A2(n12565), .ZN(n12740) );
  NAND2_X1 U14418 ( .A1(n12740), .A2(n13243), .ZN(n12567) );
  AND2_X1 U14419 ( .A1(n12567), .A2(n13421), .ZN(n12598) );
  NAND3_X1 U14420 ( .A1(n12740), .A2(n13407), .A3(n13243), .ZN(n12568) );
  OAI211_X1 U14421 ( .C1(n13421), .C2(n13419), .A(n12568), .B(n12612), .ZN(
        n12569) );
  AOI21_X1 U14422 ( .B1(n13419), .B2(n12598), .A(n12569), .ZN(n12570) );
  NAND2_X1 U14423 ( .A1(n12603), .A2(n12572), .ZN(n13471) );
  INV_X1 U14424 ( .A(n13478), .ZN(n13481) );
  NOR2_X1 U14425 ( .A1(n13471), .A2(n13481), .ZN(n12573) );
  INV_X1 U14426 ( .A(n13532), .ZN(n12589) );
  NAND2_X1 U14427 ( .A1(n12701), .A2(n12702), .ZN(n13565) );
  NOR3_X1 U14428 ( .A1(n12576), .A2(n12575), .A3(n12574), .ZN(n12577) );
  NAND3_X1 U14429 ( .A1(n12577), .A2(n12647), .A3(n12652), .ZN(n12580) );
  INV_X1 U14430 ( .A(n12664), .ZN(n12579) );
  NAND4_X1 U14431 ( .A1(n15715), .A2(n12626), .A3(n12637), .A4(n12632), .ZN(
        n12578) );
  NOR3_X1 U14432 ( .A1(n12580), .A2(n12579), .A3(n12578), .ZN(n12582) );
  NAND4_X1 U14433 ( .A1(n12582), .A2(n12658), .A3(n12642), .A4(n12581), .ZN(
        n12585) );
  NOR4_X1 U14434 ( .A1(n12585), .A2(n12584), .A3(n7395), .A4(n12583), .ZN(
        n12586) );
  NAND4_X1 U14435 ( .A1(n13578), .A2(n13611), .A3(n13599), .A4(n12586), .ZN(
        n12587) );
  NOR4_X1 U14436 ( .A1(n12589), .A2(n12588), .A3(n13565), .A4(n12587), .ZN(
        n12590) );
  NAND4_X1 U14437 ( .A1(n13493), .A2(n13505), .A3(n12590), .A4(n13524), .ZN(
        n12591) );
  NOR4_X1 U14438 ( .A1(n12732), .A2(n13437), .A3(n12611), .A4(n12591), .ZN(
        n12592) );
  NAND2_X1 U14439 ( .A1(n13421), .A2(n13423), .ZN(n12741) );
  NAND4_X1 U14440 ( .A1(n12743), .A2(n12592), .A3(n12741), .A4(n12740), .ZN(
        n12593) );
  MUX2_X1 U14441 ( .A(n13407), .B(n12594), .S(n12593), .Z(n12595) );
  INV_X1 U14442 ( .A(n12736), .ZN(n12596) );
  NAND3_X1 U14443 ( .A1(n12735), .A2(n12612), .A3(n13419), .ZN(n12599) );
  INV_X1 U14444 ( .A(n12603), .ZN(n12605) );
  OAI21_X1 U14445 ( .B1(n12606), .B2(n12605), .A(n12604), .ZN(n12608) );
  NAND2_X1 U14446 ( .A1(n12608), .A2(n12607), .ZN(n12610) );
  INV_X1 U14447 ( .A(n12611), .ZN(n12725) );
  NAND3_X1 U14448 ( .A1(n12618), .A2(n12617), .A3(n12612), .ZN(n12613) );
  NAND2_X1 U14449 ( .A1(n12613), .A2(n12738), .ZN(n12616) );
  NAND2_X1 U14450 ( .A1(n12623), .A2(n12614), .ZN(n12615) );
  AOI22_X1 U14451 ( .A1(n15715), .A2(n12616), .B1(n12738), .B2(n12615), .ZN(
        n12621) );
  NAND2_X1 U14452 ( .A1(n12618), .A2(n12617), .ZN(n12619) );
  AOI21_X1 U14453 ( .B1(n15712), .B2(n12621), .A(n12620), .ZN(n12628) );
  AOI21_X1 U14454 ( .B1(n12624), .B2(n12622), .A(n12738), .ZN(n12627) );
  MUX2_X1 U14455 ( .A(n12624), .B(n12623), .S(n12727), .Z(n12625) );
  OAI211_X1 U14456 ( .C1(n12628), .C2(n12627), .A(n12626), .B(n12625), .ZN(
        n12633) );
  MUX2_X1 U14457 ( .A(n12630), .B(n12629), .S(n12738), .Z(n12631) );
  NAND3_X1 U14458 ( .A1(n12633), .A2(n12632), .A3(n12631), .ZN(n12638) );
  MUX2_X1 U14459 ( .A(n12635), .B(n12634), .S(n12727), .Z(n12636) );
  NAND3_X1 U14460 ( .A1(n12638), .A2(n12637), .A3(n12636), .ZN(n12643) );
  MUX2_X1 U14461 ( .A(n12640), .B(n12639), .S(n12738), .Z(n12641) );
  NAND3_X1 U14462 ( .A1(n12643), .A2(n12642), .A3(n12641), .ZN(n12648) );
  OR2_X1 U14463 ( .A1(n15830), .A2(n12738), .ZN(n12645) );
  NAND2_X1 U14464 ( .A1(n15830), .A2(n12738), .ZN(n12644) );
  MUX2_X1 U14465 ( .A(n12645), .B(n12644), .S(n13256), .Z(n12646) );
  NAND3_X1 U14466 ( .A1(n12648), .A2(n12647), .A3(n12646), .ZN(n12653) );
  MUX2_X1 U14467 ( .A(n12650), .B(n12649), .S(n12738), .Z(n12651) );
  NAND3_X1 U14468 ( .A1(n12653), .A2(n12652), .A3(n12651), .ZN(n12659) );
  INV_X1 U14469 ( .A(n12654), .ZN(n12655) );
  MUX2_X1 U14470 ( .A(n12656), .B(n12655), .S(n12727), .Z(n12657) );
  NAND3_X1 U14471 ( .A1(n12659), .A2(n12658), .A3(n12657), .ZN(n12663) );
  NAND2_X1 U14472 ( .A1(n15892), .A2(n12738), .ZN(n12661) );
  OR2_X1 U14473 ( .A1(n15892), .A2(n12738), .ZN(n12660) );
  MUX2_X1 U14474 ( .A(n12661), .B(n12660), .S(n13254), .Z(n12662) );
  NAND2_X1 U14475 ( .A1(n12663), .A2(n12662), .ZN(n12665) );
  NAND2_X1 U14476 ( .A1(n12665), .A2(n12664), .ZN(n12669) );
  NAND3_X1 U14477 ( .A1(n12669), .A2(n12666), .A3(n12672), .ZN(n12667) );
  NAND2_X1 U14478 ( .A1(n12667), .A2(n12670), .ZN(n12675) );
  NAND2_X1 U14479 ( .A1(n12669), .A2(n12668), .ZN(n12673) );
  INV_X1 U14480 ( .A(n12670), .ZN(n12671) );
  AOI21_X1 U14481 ( .B1(n12673), .B2(n12672), .A(n12671), .ZN(n12674) );
  MUX2_X1 U14482 ( .A(n12675), .B(n12674), .S(n12727), .Z(n12679) );
  MUX2_X1 U14483 ( .A(n12677), .B(n12676), .S(n12738), .Z(n12678) );
  OAI211_X1 U14484 ( .C1(n12679), .C2(n7395), .A(n13638), .B(n12678), .ZN(
        n12683) );
  NAND2_X1 U14485 ( .A1(n13793), .A2(n13627), .ZN(n12680) );
  MUX2_X1 U14486 ( .A(n12681), .B(n12680), .S(n12738), .Z(n12682) );
  NAND3_X1 U14487 ( .A1(n12683), .A2(n13624), .A3(n12682), .ZN(n12687) );
  MUX2_X1 U14488 ( .A(n12685), .B(n12684), .S(n12738), .Z(n12686) );
  NAND3_X1 U14489 ( .A1(n12687), .A2(n13611), .A3(n12686), .ZN(n12692) );
  AND2_X1 U14490 ( .A1(n12693), .A2(n12688), .ZN(n12689) );
  MUX2_X1 U14491 ( .A(n12690), .B(n12689), .S(n12727), .Z(n12691) );
  NAND4_X1 U14492 ( .A1(n12692), .A2(n13599), .A3(n13561), .A4(n12691), .ZN(
        n12700) );
  INV_X1 U14493 ( .A(n12693), .ZN(n12695) );
  OAI211_X1 U14494 ( .C1(n12695), .C2(n12694), .A(n12701), .B(n13561), .ZN(
        n12696) );
  INV_X1 U14495 ( .A(n12696), .ZN(n12697) );
  MUX2_X1 U14496 ( .A(n12698), .B(n12697), .S(n12727), .Z(n12699) );
  NAND2_X1 U14497 ( .A1(n12700), .A2(n12699), .ZN(n12704) );
  MUX2_X1 U14498 ( .A(n12702), .B(n12701), .S(n12738), .Z(n12703) );
  NAND3_X1 U14499 ( .A1(n12704), .A2(n13546), .A3(n12703), .ZN(n12708) );
  MUX2_X1 U14500 ( .A(n12706), .B(n12705), .S(n12727), .Z(n12707) );
  NAND3_X1 U14501 ( .A1(n12708), .A2(n13532), .A3(n12707), .ZN(n12712) );
  MUX2_X1 U14502 ( .A(n12710), .B(n12709), .S(n12738), .Z(n12711) );
  NAND3_X1 U14503 ( .A1(n12712), .A2(n13524), .A3(n12711), .ZN(n12716) );
  NAND2_X1 U14504 ( .A1(n13509), .A2(n12727), .ZN(n12714) );
  NAND2_X1 U14505 ( .A1(n13534), .A2(n12738), .ZN(n12713) );
  MUX2_X1 U14506 ( .A(n12714), .B(n12713), .S(n13525), .Z(n12715) );
  NAND3_X1 U14507 ( .A1(n12716), .A2(n13505), .A3(n12715), .ZN(n12720) );
  MUX2_X1 U14508 ( .A(n12718), .B(n12717), .S(n12738), .Z(n12719) );
  NAND2_X1 U14509 ( .A1(n12720), .A2(n12719), .ZN(n12721) );
  NAND2_X1 U14510 ( .A1(n12721), .A2(n13493), .ZN(n12723) );
  NAND3_X1 U14511 ( .A1(n13181), .A2(n13486), .A3(n12727), .ZN(n12722) );
  NAND2_X1 U14512 ( .A1(n12723), .A2(n12722), .ZN(n12724) );
  AOI21_X1 U14513 ( .B1(n12725), .B2(n12724), .A(n13437), .ZN(n12726) );
  MUX2_X1 U14514 ( .A(n12729), .B(n12728), .S(n12727), .Z(n12730) );
  INV_X1 U14515 ( .A(n12730), .ZN(n12731) );
  NOR2_X1 U14516 ( .A1(n12732), .A2(n12731), .ZN(n12733) );
  NAND2_X1 U14517 ( .A1(n12734), .A2(n12733), .ZN(n12737) );
  NAND2_X1 U14518 ( .A1(n12737), .A2(n12735), .ZN(n12739) );
  INV_X1 U14519 ( .A(n12741), .ZN(n12742) );
  NAND3_X1 U14520 ( .A1(n12752), .A2(n12751), .A3(n13408), .ZN(n12753) );
  OAI211_X1 U14521 ( .C1(n12754), .C2(n12756), .A(n12753), .B(P3_B_REG_SCAN_IN), .ZN(n12755) );
  OAI21_X1 U14522 ( .B1(n12757), .B2(n12756), .A(n12755), .ZN(P3_U3296) );
  INV_X1 U14523 ( .A(n14483), .ZN(n12759) );
  OAI222_X1 U14524 ( .A1(n15210), .A2(n12760), .B1(n15215), .B2(n12759), .C1(
        P1_U3086), .C2(n12758), .ZN(P1_U3327) );
  AND2_X4 U14525 ( .A1(n12761), .A2(n14507), .ZN(n12781) );
  NAND2_X1 U14526 ( .A1(n14023), .A2(n12920), .ZN(n12763) );
  NAND2_X1 U14527 ( .A1(n12795), .A2(n12794), .ZN(n12762) );
  NAND2_X1 U14528 ( .A1(n12763), .A2(n12762), .ZN(n12797) );
  NAND2_X1 U14529 ( .A1(n12765), .A2(n12764), .ZN(n12784) );
  NAND2_X1 U14530 ( .A1(n12772), .A2(n12768), .ZN(n12769) );
  NAND2_X1 U14531 ( .A1(n14507), .A2(n14078), .ZN(n12767) );
  NAND3_X1 U14532 ( .A1(n12773), .A2(n12772), .A3(n12848), .ZN(n12774) );
  AOI21_X1 U14533 ( .B1(n12784), .B2(n12785), .A(n12777), .ZN(n12789) );
  NAND2_X1 U14534 ( .A1(n12848), .A2(n12780), .ZN(n12778) );
  NAND2_X1 U14535 ( .A1(n12781), .A2(n12780), .ZN(n12782) );
  NAND2_X1 U14536 ( .A1(n14022), .A2(n12795), .ZN(n12791) );
  NAND2_X1 U14537 ( .A1(n13958), .A2(n12848), .ZN(n12790) );
  AND2_X1 U14538 ( .A1(n12791), .A2(n12790), .ZN(n12800) );
  NAND2_X1 U14539 ( .A1(n13958), .A2(n12795), .ZN(n12793) );
  NAND2_X1 U14540 ( .A1(n14022), .A2(n12920), .ZN(n12792) );
  NAND2_X1 U14541 ( .A1(n12793), .A2(n12792), .ZN(n12799) );
  AOI22_X1 U14542 ( .A1(n12795), .A2(n14023), .B1(n12920), .B2(n12794), .ZN(
        n12796) );
  AOI21_X1 U14543 ( .B1(n12798), .B2(n12797), .A(n12796), .ZN(n12802) );
  NAND2_X1 U14544 ( .A1(n12800), .A2(n12799), .ZN(n12801) );
  NAND2_X1 U14545 ( .A1(n15804), .A2(n12795), .ZN(n12805) );
  NAND2_X1 U14546 ( .A1(n14021), .A2(n12920), .ZN(n12804) );
  NAND2_X1 U14547 ( .A1(n15804), .A2(n12920), .ZN(n12806) );
  INV_X1 U14548 ( .A(n12810), .ZN(n12811) );
  NAND2_X1 U14549 ( .A1(n15819), .A2(n12920), .ZN(n12813) );
  NAND2_X1 U14550 ( .A1(n14020), .A2(n12795), .ZN(n12812) );
  INV_X1 U14551 ( .A(n12781), .ZN(n12920) );
  NAND2_X1 U14552 ( .A1(n15819), .A2(n12795), .ZN(n12814) );
  OAI21_X1 U14553 ( .B1(n12815), .B2(n12956), .A(n12814), .ZN(n12816) );
  INV_X1 U14554 ( .A(n12817), .ZN(n12818) );
  NAND2_X1 U14555 ( .A1(n15844), .A2(n12781), .ZN(n12821) );
  NAND2_X1 U14556 ( .A1(n14019), .A2(n12965), .ZN(n12820) );
  NAND2_X1 U14557 ( .A1(n12821), .A2(n12820), .ZN(n12824) );
  AOI22_X1 U14558 ( .A1(n15844), .A2(n12965), .B1(n12956), .B2(n14019), .ZN(
        n12822) );
  NAND2_X1 U14559 ( .A1(n12828), .A2(n12920), .ZN(n12827) );
  NAND2_X1 U14560 ( .A1(n14018), .A2(n12781), .ZN(n12826) );
  NAND2_X1 U14561 ( .A1(n12827), .A2(n12826), .ZN(n12832) );
  NAND2_X1 U14562 ( .A1(n12828), .A2(n12795), .ZN(n12829) );
  OAI21_X1 U14563 ( .B1(n12830), .B2(n12795), .A(n12829), .ZN(n12831) );
  INV_X1 U14564 ( .A(n12832), .ZN(n12833) );
  NAND2_X1 U14565 ( .A1(n12836), .A2(n12795), .ZN(n12835) );
  NAND2_X1 U14566 ( .A1(n14017), .A2(n12965), .ZN(n12834) );
  NAND2_X1 U14567 ( .A1(n12835), .A2(n12834), .ZN(n12838) );
  AOI22_X1 U14568 ( .A1(n12836), .A2(n12965), .B1(n12795), .B2(n14017), .ZN(
        n12837) );
  NAND2_X1 U14569 ( .A1(n12844), .A2(n12920), .ZN(n12843) );
  NAND2_X1 U14570 ( .A1(n14016), .A2(n12781), .ZN(n12842) );
  NAND2_X1 U14571 ( .A1(n12844), .A2(n12781), .ZN(n12845) );
  OAI21_X1 U14572 ( .B1(n12846), .B2(n12781), .A(n12845), .ZN(n12847) );
  NAND2_X1 U14573 ( .A1(n12851), .A2(n12956), .ZN(n12850) );
  NAND2_X1 U14574 ( .A1(n14015), .A2(n12965), .ZN(n12849) );
  NAND2_X1 U14575 ( .A1(n12850), .A2(n12849), .ZN(n12853) );
  AOI22_X1 U14576 ( .A1(n12851), .A2(n12965), .B1(n12781), .B2(n14015), .ZN(
        n12852) );
  NAND2_X1 U14577 ( .A1(n12857), .A2(n12965), .ZN(n12856) );
  NAND2_X1 U14578 ( .A1(n14014), .A2(n12781), .ZN(n12855) );
  NAND2_X1 U14579 ( .A1(n12856), .A2(n12855), .ZN(n12861) );
  NAND2_X1 U14580 ( .A1(n12857), .A2(n12781), .ZN(n12858) );
  OAI21_X1 U14581 ( .B1(n12859), .B2(n12956), .A(n12858), .ZN(n12860) );
  INV_X1 U14582 ( .A(n12861), .ZN(n12862) );
  NAND2_X1 U14583 ( .A1(n12865), .A2(n12781), .ZN(n12864) );
  NAND2_X1 U14584 ( .A1(n14013), .A2(n12965), .ZN(n12863) );
  NAND2_X1 U14585 ( .A1(n12864), .A2(n12863), .ZN(n12867) );
  AOI22_X1 U14586 ( .A1(n12865), .A2(n12965), .B1(n12795), .B2(n14013), .ZN(
        n12866) );
  NAND2_X1 U14587 ( .A1(n12873), .A2(n12965), .ZN(n12872) );
  NAND2_X1 U14588 ( .A1(n14012), .A2(n12795), .ZN(n12871) );
  AOI22_X1 U14590 ( .A1(n12873), .A2(n12956), .B1(n14012), .B2(n12965), .ZN(
        n12874) );
  NAND2_X1 U14591 ( .A1(n12877), .A2(n12781), .ZN(n12876) );
  NAND2_X1 U14592 ( .A1(n14011), .A2(n12965), .ZN(n12875) );
  NAND2_X1 U14593 ( .A1(n12876), .A2(n12875), .ZN(n12881) );
  NAND2_X1 U14594 ( .A1(n12877), .A2(n12965), .ZN(n12878) );
  OAI21_X1 U14595 ( .B1(n12879), .B2(n12920), .A(n12878), .ZN(n12880) );
  NAND2_X1 U14596 ( .A1(n14471), .A2(n12965), .ZN(n12883) );
  NAND2_X1 U14597 ( .A1(n14010), .A2(n12795), .ZN(n12882) );
  NAND2_X1 U14598 ( .A1(n12883), .A2(n12882), .ZN(n12885) );
  AOI22_X1 U14599 ( .A1(n14471), .A2(n12956), .B1(n14010), .B2(n12965), .ZN(
        n12884) );
  NAND2_X1 U14600 ( .A1(n14320), .A2(n12956), .ZN(n12888) );
  NAND2_X1 U14601 ( .A1(n14009), .A2(n12965), .ZN(n12887) );
  NAND2_X1 U14602 ( .A1(n14320), .A2(n12920), .ZN(n12889) );
  OAI21_X1 U14603 ( .B1(n14284), .B2(n12965), .A(n12889), .ZN(n12890) );
  NAND2_X1 U14604 ( .A1(n14408), .A2(n12920), .ZN(n12892) );
  NAND2_X1 U14605 ( .A1(n14008), .A2(n12795), .ZN(n12891) );
  NAND2_X1 U14606 ( .A1(n12892), .A2(n12891), .ZN(n12894) );
  NAND2_X1 U14607 ( .A1(n14461), .A2(n12956), .ZN(n12896) );
  NAND2_X1 U14608 ( .A1(n14243), .A2(n12965), .ZN(n12895) );
  NAND2_X1 U14609 ( .A1(n12896), .A2(n12895), .ZN(n12899) );
  NAND2_X1 U14610 ( .A1(n14461), .A2(n12965), .ZN(n12897) );
  OAI21_X1 U14611 ( .B1(n14286), .B2(n12920), .A(n12897), .ZN(n12898) );
  NAND2_X1 U14612 ( .A1(n14396), .A2(n12965), .ZN(n12902) );
  NAND2_X1 U14613 ( .A1(n14263), .A2(n12781), .ZN(n12901) );
  NAND2_X1 U14614 ( .A1(n12902), .A2(n12901), .ZN(n12907) );
  AOI22_X1 U14615 ( .A1(n14396), .A2(n12781), .B1(n14263), .B2(n12965), .ZN(
        n12903) );
  INV_X1 U14616 ( .A(n12903), .ZN(n12904) );
  INV_X1 U14617 ( .A(n12906), .ZN(n12909) );
  INV_X1 U14618 ( .A(n12907), .ZN(n12908) );
  NAND2_X1 U14619 ( .A1(n12909), .A2(n12908), .ZN(n12910) );
  NAND2_X1 U14620 ( .A1(n14456), .A2(n12781), .ZN(n12912) );
  NAND2_X1 U14621 ( .A1(n14244), .A2(n12920), .ZN(n12911) );
  NAND2_X1 U14622 ( .A1(n12912), .A2(n12911), .ZN(n12914) );
  AOI22_X1 U14623 ( .A1(n14456), .A2(n12965), .B1(n12956), .B2(n14244), .ZN(
        n12913) );
  AOI22_X1 U14624 ( .A1(n14386), .A2(n12795), .B1(n14007), .B2(n12965), .ZN(
        n12916) );
  INV_X1 U14625 ( .A(n12918), .ZN(n12919) );
  AOI22_X1 U14626 ( .A1(n14193), .A2(n12795), .B1(n14204), .B2(n12965), .ZN(
        n12923) );
  OAI22_X1 U14627 ( .A1(n14452), .A2(n12956), .B1(n14171), .B2(n12965), .ZN(
        n12921) );
  INV_X1 U14628 ( .A(n12921), .ZN(n12922) );
  NAND2_X1 U14629 ( .A1(n12928), .A2(n12929), .ZN(n12927) );
  AOI22_X1 U14630 ( .A1(n12924), .A2(n12781), .B1(n14006), .B2(n12965), .ZN(
        n12925) );
  INV_X1 U14631 ( .A(n12928), .ZN(n12931) );
  INV_X1 U14632 ( .A(n12929), .ZN(n12930) );
  NAND2_X1 U14633 ( .A1(n12931), .A2(n12930), .ZN(n12932) );
  AOI22_X1 U14634 ( .A1(n14158), .A2(n12795), .B1(n14169), .B2(n12965), .ZN(
        n12935) );
  OAI22_X1 U14635 ( .A1(n14445), .A2(n12795), .B1(n14134), .B2(n12920), .ZN(
        n12933) );
  OAI22_X1 U14636 ( .A1(n14441), .A2(n12781), .B1(n14151), .B2(n12920), .ZN(
        n12938) );
  INV_X1 U14637 ( .A(n14151), .ZN(n14113) );
  AOI22_X1 U14638 ( .A1(n14363), .A2(n12781), .B1(n14113), .B2(n12965), .ZN(
        n12937) );
  INV_X1 U14639 ( .A(n12938), .ZN(n12939) );
  OAI22_X1 U14640 ( .A1(n14437), .A2(n12920), .B1(n14135), .B2(n12956), .ZN(
        n12954) );
  AND2_X1 U14641 ( .A1(n14114), .A2(n12920), .ZN(n12941) );
  AOI21_X1 U14642 ( .B1(n14341), .B2(n12781), .A(n12941), .ZN(n12975) );
  NAND2_X1 U14643 ( .A1(n14341), .A2(n12920), .ZN(n12943) );
  NAND2_X1 U14644 ( .A1(n14114), .A2(n12956), .ZN(n12942) );
  NAND2_X1 U14645 ( .A1(n12943), .A2(n12942), .ZN(n12973) );
  AND2_X1 U14646 ( .A1(n14100), .A2(n12965), .ZN(n12944) );
  AOI21_X1 U14647 ( .B1(n14337), .B2(n12781), .A(n12944), .ZN(n12969) );
  NAND2_X1 U14648 ( .A1(n14337), .A2(n12965), .ZN(n12946) );
  NAND2_X1 U14649 ( .A1(n14100), .A2(n12956), .ZN(n12945) );
  NAND2_X1 U14650 ( .A1(n12946), .A2(n12945), .ZN(n12968) );
  AND2_X1 U14651 ( .A1(n12969), .A2(n12968), .ZN(n12974) );
  NAND2_X1 U14652 ( .A1(n15194), .A2(n12959), .ZN(n12948) );
  OR2_X1 U14653 ( .A1(n12960), .A2(n14479), .ZN(n12947) );
  NAND2_X1 U14654 ( .A1(n12468), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n12951) );
  NAND2_X1 U14655 ( .A1(n12064), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n12950) );
  NAND2_X1 U14656 ( .A1(n7508), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n12949) );
  AND3_X1 U14657 ( .A1(n12951), .A2(n12950), .A3(n12949), .ZN(n12958) );
  XNOR2_X1 U14658 ( .A(n14330), .B(n12958), .ZN(n12972) );
  AOI211_X1 U14659 ( .C1(n12975), .C2(n12973), .A(n12974), .B(n12972), .ZN(
        n12952) );
  AOI22_X1 U14660 ( .A1(n14122), .A2(n12965), .B1(n12781), .B2(n14101), .ZN(
        n12953) );
  MUX2_X1 U14661 ( .A(n14085), .B(n12956), .S(n14330), .Z(n12957) );
  OAI21_X1 U14662 ( .B1(n12958), .B2(n12920), .A(n12957), .ZN(n12971) );
  NAND2_X1 U14663 ( .A1(n13059), .A2(n12959), .ZN(n12962) );
  INV_X1 U14664 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13120) );
  OR2_X1 U14665 ( .A1(n12960), .A2(n13120), .ZN(n12961) );
  NAND2_X1 U14666 ( .A1(n12965), .A2(n14085), .ZN(n12986) );
  NAND2_X1 U14667 ( .A1(n13057), .A2(n12963), .ZN(n13033) );
  NAND4_X1 U14668 ( .A1(n12986), .A2(n13030), .A3(n13053), .A4(n13033), .ZN(
        n12964) );
  AOI22_X1 U14669 ( .A1(n14334), .A2(n12781), .B1(n14005), .B2(n12964), .ZN(
        n13035) );
  NAND2_X1 U14670 ( .A1(n14334), .A2(n12965), .ZN(n12967) );
  NAND2_X1 U14671 ( .A1(n14005), .A2(n12781), .ZN(n12966) );
  NAND2_X1 U14672 ( .A1(n12967), .A2(n12966), .ZN(n13034) );
  OAI22_X1 U14673 ( .A1(n13035), .A2(n13034), .B1(n12969), .B2(n12968), .ZN(
        n12970) );
  NAND2_X1 U14674 ( .A1(n12971), .A2(n12970), .ZN(n12980) );
  INV_X1 U14675 ( .A(n12972), .ZN(n13027) );
  INV_X1 U14676 ( .A(n12973), .ZN(n12978) );
  INV_X1 U14677 ( .A(n12974), .ZN(n12977) );
  INV_X1 U14678 ( .A(n12975), .ZN(n12976) );
  NAND4_X1 U14679 ( .A1(n13027), .A2(n12978), .A3(n12977), .A4(n12976), .ZN(
        n12979) );
  NAND2_X1 U14680 ( .A1(n14507), .A2(n12981), .ZN(n12982) );
  NAND2_X1 U14681 ( .A1(n12982), .A2(n14078), .ZN(n12984) );
  NAND2_X1 U14682 ( .A1(n12984), .A2(n12983), .ZN(n13039) );
  INV_X1 U14683 ( .A(n13039), .ZN(n12985) );
  INV_X1 U14684 ( .A(n12986), .ZN(n12988) );
  NOR2_X1 U14685 ( .A1(n14330), .A2(n14085), .ZN(n12987) );
  AOI211_X1 U14686 ( .C1(n12795), .C2(n14330), .A(n12988), .B(n12987), .ZN(
        n13045) );
  INV_X1 U14687 ( .A(n13045), .ZN(n12989) );
  XNOR2_X1 U14688 ( .A(n14334), .B(n14005), .ZN(n13024) );
  NAND2_X1 U14689 ( .A1(n12991), .A2(n12990), .ZN(n14186) );
  NOR2_X1 U14690 ( .A1(n12992), .A2(n10408), .ZN(n12995) );
  NAND4_X1 U14691 ( .A1(n12995), .A2(n15689), .A3(n12994), .A4(n12993), .ZN(
        n12997) );
  NOR2_X1 U14692 ( .A1(n12997), .A2(n12996), .ZN(n13000) );
  NAND4_X1 U14693 ( .A1(n13001), .A2(n13000), .A3(n12999), .A4(n12998), .ZN(
        n13002) );
  NOR4_X1 U14694 ( .A1(n13005), .A2(n13004), .A3(n13003), .A4(n13002), .ZN(
        n13007) );
  NAND4_X1 U14695 ( .A1(n13009), .A2(n13008), .A3(n13007), .A4(n13006), .ZN(
        n13010) );
  NOR2_X1 U14696 ( .A1(n13011), .A2(n13010), .ZN(n13013) );
  NAND4_X1 U14697 ( .A1(n14313), .A2(n13014), .A3(n13013), .A4(n13012), .ZN(
        n13015) );
  NOR2_X1 U14698 ( .A1(n14288), .A2(n13015), .ZN(n13017) );
  NAND3_X1 U14699 ( .A1(n14240), .A2(n13017), .A3(n13016), .ZN(n13018) );
  NOR2_X1 U14700 ( .A1(n14220), .A2(n13018), .ZN(n13019) );
  NAND4_X1 U14701 ( .A1(n14186), .A2(n14133), .A3(n13019), .A4(n14213), .ZN(
        n13020) );
  NOR2_X1 U14702 ( .A1(n14148), .A2(n13020), .ZN(n13023) );
  AND4_X1 U14703 ( .A1(n13024), .A2(n13023), .A3(n13022), .A4(n13021), .ZN(
        n13026) );
  NAND4_X1 U14704 ( .A1(n13027), .A2(n14094), .A3(n13026), .A4(n13025), .ZN(
        n13028) );
  XNOR2_X1 U14705 ( .A(n13028), .B(n14078), .ZN(n13029) );
  AND2_X1 U14706 ( .A1(n13029), .A2(n7526), .ZN(n13043) );
  NOR2_X1 U14707 ( .A1(n10408), .A2(n14073), .ZN(n13031) );
  NAND2_X1 U14708 ( .A1(n13031), .A2(n13030), .ZN(n13032) );
  NAND2_X1 U14709 ( .A1(n13033), .A2(n13032), .ZN(n13037) );
  NAND2_X1 U14710 ( .A1(n13035), .A2(n13034), .ZN(n13038) );
  INV_X1 U14711 ( .A(n13037), .ZN(n13042) );
  INV_X1 U14712 ( .A(n13038), .ZN(n13040) );
  NAND2_X1 U14713 ( .A1(n13040), .A2(n12985), .ZN(n13041) );
  MUX2_X1 U14714 ( .A(n13042), .B(n13041), .S(n12989), .Z(n13047) );
  OAI21_X1 U14715 ( .B1(n13045), .B2(n13044), .A(n13043), .ZN(n13046) );
  OR2_X1 U14716 ( .A1(n13051), .A2(P2_U3088), .ZN(n14501) );
  INV_X1 U14717 ( .A(n14501), .ZN(n13052) );
  INV_X1 U14718 ( .A(n14487), .ZN(n13055) );
  INV_X1 U14719 ( .A(n13053), .ZN(n13054) );
  NAND4_X1 U14720 ( .A1(n15340), .A2(n13055), .A3(n13054), .A4(n14242), .ZN(
        n13056) );
  OAI211_X1 U14721 ( .C1(n13057), .C2(n14501), .A(n13056), .B(P2_B_REG_SCAN_IN), .ZN(n13058) );
  INV_X1 U14722 ( .A(n13059), .ZN(n13121) );
  OAI222_X1 U14723 ( .A1(n15215), .A2(n13121), .B1(P1_U3086), .B2(n8888), .C1(
        n13060), .C2(n15210), .ZN(P1_U3325) );
  XNOR2_X1 U14724 ( .A(n13784), .B(n13109), .ZN(n13070) );
  XNOR2_X1 U14725 ( .A(n13789), .B(n13109), .ZN(n13065) );
  INV_X1 U14726 ( .A(n13065), .ZN(n13066) );
  XNOR2_X1 U14727 ( .A(n13065), .B(n13641), .ZN(n13230) );
  XNOR2_X1 U14728 ( .A(n13726), .B(n13109), .ZN(n13067) );
  XNOR2_X1 U14729 ( .A(n13067), .B(n13626), .ZN(n13166) );
  NAND2_X1 U14730 ( .A1(n13167), .A2(n13166), .ZN(n13165) );
  INV_X1 U14731 ( .A(n13067), .ZN(n13068) );
  NAND2_X1 U14732 ( .A1(n13068), .A2(n13626), .ZN(n13069) );
  NAND2_X1 U14733 ( .A1(n13165), .A2(n13069), .ZN(n13174) );
  XNOR2_X1 U14734 ( .A(n13070), .B(n13251), .ZN(n13175) );
  XNOR2_X1 U14735 ( .A(n13717), .B(n13109), .ZN(n13072) );
  XNOR2_X1 U14736 ( .A(n13072), .B(n13590), .ZN(n13209) );
  XNOR2_X1 U14737 ( .A(n13713), .B(n13109), .ZN(n13077) );
  XNOR2_X1 U14738 ( .A(n13077), .B(n13249), .ZN(n13137) );
  INV_X1 U14739 ( .A(n13137), .ZN(n13074) );
  OR2_X1 U14740 ( .A1(n13209), .A2(n13074), .ZN(n13071) );
  INV_X1 U14741 ( .A(n13072), .ZN(n13073) );
  NAND2_X1 U14742 ( .A1(n13073), .A2(n13250), .ZN(n13135) );
  OR2_X1 U14743 ( .A1(n13074), .A2(n13135), .ZN(n13075) );
  INV_X1 U14744 ( .A(n13075), .ZN(n13076) );
  INV_X1 U14745 ( .A(n13077), .ZN(n13078) );
  XNOR2_X1 U14746 ( .A(n13554), .B(n13109), .ZN(n13079) );
  XNOR2_X1 U14747 ( .A(n13079), .B(n13568), .ZN(n13194) );
  XNOR2_X1 U14748 ( .A(n13539), .B(n13106), .ZN(n13081) );
  NAND2_X1 U14749 ( .A1(n13081), .A2(n13247), .ZN(n13145) );
  INV_X1 U14750 ( .A(n13145), .ZN(n13080) );
  OR2_X1 U14751 ( .A1(n13194), .A2(n13080), .ZN(n13085) );
  NAND2_X1 U14752 ( .A1(n13079), .A2(n13568), .ZN(n13144) );
  OR2_X1 U14753 ( .A1(n13080), .A2(n13144), .ZN(n13083) );
  INV_X1 U14754 ( .A(n13081), .ZN(n13082) );
  NAND2_X1 U14755 ( .A1(n13082), .A2(n13548), .ZN(n13146) );
  XNOR2_X1 U14756 ( .A(n13525), .B(n13109), .ZN(n13086) );
  NAND2_X1 U14757 ( .A1(n13087), .A2(n13086), .ZN(n13090) );
  NAND2_X1 U14758 ( .A1(n13200), .A2(n13090), .ZN(n13095) );
  XNOR2_X1 U14759 ( .A(n13514), .B(n7218), .ZN(n13094) );
  INV_X1 U14760 ( .A(n13094), .ZN(n13091) );
  OR2_X1 U14761 ( .A1(n13509), .A2(n13091), .ZN(n13089) );
  OR2_X1 U14762 ( .A1(n13091), .A2(n13090), .ZN(n13092) );
  AND2_X2 U14763 ( .A1(n13093), .A2(n13092), .ZN(n13182) );
  XNOR2_X1 U14764 ( .A(n13181), .B(n13109), .ZN(n13096) );
  INV_X1 U14765 ( .A(n13096), .ZN(n13097) );
  NAND2_X1 U14766 ( .A1(n13097), .A2(n13508), .ZN(n13098) );
  NAND2_X1 U14767 ( .A1(n13154), .A2(n13155), .ZN(n13102) );
  XNOR2_X1 U14768 ( .A(n13688), .B(n7218), .ZN(n13099) );
  NAND2_X1 U14769 ( .A1(n13099), .A2(n13495), .ZN(n13103) );
  INV_X1 U14770 ( .A(n13099), .ZN(n13100) );
  NAND2_X1 U14771 ( .A1(n13100), .A2(n13245), .ZN(n13101) );
  NAND2_X1 U14772 ( .A1(n13102), .A2(n13156), .ZN(n13158) );
  XNOR2_X1 U14773 ( .A(n13217), .B(n13106), .ZN(n13104) );
  NOR2_X1 U14774 ( .A1(n13104), .A2(n13483), .ZN(n13105) );
  AOI21_X1 U14775 ( .B1(n13104), .B2(n13483), .A(n13105), .ZN(n13220) );
  XNOR2_X1 U14776 ( .A(n13680), .B(n13106), .ZN(n13107) );
  NOR2_X1 U14777 ( .A1(n13107), .A2(n13244), .ZN(n13108) );
  AOI21_X1 U14778 ( .B1(n13107), .B2(n13244), .A(n13108), .ZN(n13122) );
  XNOR2_X1 U14779 ( .A(n7769), .B(n13109), .ZN(n13110) );
  XNOR2_X1 U14780 ( .A(n13111), .B(n13110), .ZN(n13112) );
  NAND2_X1 U14781 ( .A1(n13112), .A2(n13221), .ZN(n13118) );
  AOI22_X1 U14782 ( .A1(n13244), .A2(n13223), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13114) );
  NAND2_X1 U14783 ( .A1(n13239), .A2(n13444), .ZN(n13113) );
  OAI211_X1 U14784 ( .C1(n13439), .C2(n13225), .A(n13114), .B(n13113), .ZN(
        n13115) );
  AOI21_X1 U14785 ( .B1(n13116), .B2(n13206), .A(n13115), .ZN(n13117) );
  NAND2_X1 U14786 ( .A1(n13118), .A2(n13117), .ZN(P3_U3160) );
  OAI222_X1 U14787 ( .A1(n14506), .A2(n13121), .B1(P2_U3088), .B2(n13119), 
        .C1(n13120), .C2(n14503), .ZN(P2_U3297) );
  INV_X1 U14788 ( .A(n13680), .ZN(n13128) );
  NAND2_X1 U14789 ( .A1(n13123), .A2(n13221), .ZN(n13127) );
  AOI22_X1 U14790 ( .A1(n13483), .A2(n13223), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13124) );
  OAI21_X1 U14791 ( .B1(n13456), .B2(n13225), .A(n13124), .ZN(n13125) );
  AOI21_X1 U14792 ( .B1(n13458), .B2(n13239), .A(n13125), .ZN(n13126) );
  OAI211_X1 U14793 ( .C1(n13128), .C2(n13242), .A(n13127), .B(n13126), .ZN(
        P3_U3154) );
  AOI21_X1 U14794 ( .B1(n13246), .B2(n13129), .A(n7233), .ZN(n13134) );
  AOI22_X1 U14795 ( .A1(n13509), .A2(n13223), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13131) );
  NAND2_X1 U14796 ( .A1(n13239), .A2(n13515), .ZN(n13130) );
  OAI211_X1 U14797 ( .C1(n13486), .C2(n13225), .A(n13131), .B(n13130), .ZN(
        n13132) );
  AOI21_X1 U14798 ( .B1(n13514), .B2(n13206), .A(n13132), .ZN(n13133) );
  OAI21_X1 U14799 ( .B1(n13134), .B2(n13229), .A(n13133), .ZN(P3_U3156) );
  OR2_X1 U14800 ( .A1(n13210), .A2(n13209), .ZN(n13211) );
  NAND2_X1 U14801 ( .A1(n13211), .A2(n13135), .ZN(n13138) );
  OAI211_X1 U14802 ( .C1(n13138), .C2(n13137), .A(n13136), .B(n13221), .ZN(
        n13142) );
  NAND2_X1 U14803 ( .A1(n13250), .A2(n13223), .ZN(n13139) );
  NAND2_X1 U14804 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13418)
         );
  OAI211_X1 U14805 ( .C1(n13568), .C2(n13225), .A(n13139), .B(n13418), .ZN(
        n13140) );
  AOI21_X1 U14806 ( .B1(n13569), .B2(n13239), .A(n13140), .ZN(n13141) );
  OAI211_X1 U14807 ( .C1(n13143), .C2(n13242), .A(n13142), .B(n13141), .ZN(
        P3_U3159) );
  OR2_X1 U14808 ( .A1(n13193), .A2(n13194), .ZN(n13191) );
  NAND2_X1 U14809 ( .A1(n13191), .A2(n13144), .ZN(n13148) );
  NAND2_X1 U14810 ( .A1(n13146), .A2(n13145), .ZN(n13147) );
  XNOR2_X1 U14811 ( .A(n13148), .B(n13147), .ZN(n13153) );
  AOI22_X1 U14812 ( .A1(n13248), .A2(n13223), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13150) );
  NAND2_X1 U14813 ( .A1(n13239), .A2(n13540), .ZN(n13149) );
  OAI211_X1 U14814 ( .C1(n13534), .C2(n13225), .A(n13150), .B(n13149), .ZN(
        n13151) );
  AOI21_X1 U14815 ( .B1(n13539), .B2(n13206), .A(n13151), .ZN(n13152) );
  OAI21_X1 U14816 ( .B1(n13153), .B2(n13229), .A(n13152), .ZN(P3_U3163) );
  INV_X1 U14817 ( .A(n13688), .ZN(n13489) );
  INV_X1 U14818 ( .A(n13154), .ZN(n13184) );
  INV_X1 U14819 ( .A(n13155), .ZN(n13157) );
  NOR3_X1 U14820 ( .A1(n13184), .A2(n13157), .A3(n13156), .ZN(n13160) );
  INV_X1 U14821 ( .A(n13158), .ZN(n13159) );
  OAI21_X1 U14822 ( .B1(n13160), .B2(n13159), .A(n13221), .ZN(n13164) );
  AOI22_X1 U14823 ( .A1(n13235), .A2(n13483), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13161) );
  OAI21_X1 U14824 ( .B1(n13486), .B2(n13237), .A(n13161), .ZN(n13162) );
  AOI21_X1 U14825 ( .B1(n13487), .B2(n13239), .A(n13162), .ZN(n13163) );
  OAI211_X1 U14826 ( .C1(n13489), .C2(n13242), .A(n13164), .B(n13163), .ZN(
        P3_U3165) );
  INV_X1 U14827 ( .A(n13726), .ZN(n13617) );
  OAI211_X1 U14828 ( .C1(n13167), .C2(n13166), .A(n13165), .B(n13221), .ZN(
        n13171) );
  NAND2_X1 U14829 ( .A1(n13641), .A2(n13223), .ZN(n13168) );
  NAND2_X1 U14830 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13345)
         );
  OAI211_X1 U14831 ( .C1(n13614), .C2(n13225), .A(n13168), .B(n13345), .ZN(
        n13169) );
  AOI21_X1 U14832 ( .B1(n13615), .B2(n13239), .A(n13169), .ZN(n13170) );
  OAI211_X1 U14833 ( .C1(n13617), .C2(n13242), .A(n13171), .B(n13170), .ZN(
        P3_U3166) );
  INV_X1 U14834 ( .A(n13172), .ZN(n13173) );
  AOI21_X1 U14835 ( .B1(n13175), .B2(n13174), .A(n13173), .ZN(n13180) );
  INV_X1 U14836 ( .A(n13784), .ZN(n13598) );
  AND2_X1 U14837 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13361) );
  AOI21_X1 U14838 ( .B1(n13250), .B2(n13235), .A(n13361), .ZN(n13177) );
  NAND2_X1 U14839 ( .A1(n13239), .A2(n13595), .ZN(n13176) );
  OAI211_X1 U14840 ( .C1(n13591), .C2(n13237), .A(n13177), .B(n13176), .ZN(
        n13178) );
  AOI21_X1 U14841 ( .B1(n13598), .B2(n13206), .A(n13178), .ZN(n13179) );
  OAI21_X1 U14842 ( .B1(n13180), .B2(n13229), .A(n13179), .ZN(P3_U3168) );
  NOR3_X1 U14843 ( .A1(n7233), .A2(n8135), .A3(n13183), .ZN(n13185) );
  OAI21_X1 U14844 ( .B1(n13185), .B2(n13184), .A(n13221), .ZN(n13190) );
  NOR2_X1 U14845 ( .A1(n13522), .A2(n13237), .ZN(n13188) );
  OAI22_X1 U14846 ( .A1(n13495), .A2(n13225), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13186), .ZN(n13187) );
  AOI211_X1 U14847 ( .C1(n13500), .C2(n13239), .A(n13188), .B(n13187), .ZN(
        n13189) );
  OAI211_X1 U14848 ( .C1(n13762), .C2(n13242), .A(n13190), .B(n13189), .ZN(
        P3_U3169) );
  INV_X1 U14849 ( .A(n13191), .ZN(n13192) );
  AOI21_X1 U14850 ( .B1(n13194), .B2(n13193), .A(n13192), .ZN(n13199) );
  AOI22_X1 U14851 ( .A1(n13235), .A2(n13247), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13196) );
  NAND2_X1 U14852 ( .A1(n13239), .A2(n13555), .ZN(n13195) );
  OAI211_X1 U14853 ( .C1(n13580), .C2(n13237), .A(n13196), .B(n13195), .ZN(
        n13197) );
  AOI21_X1 U14854 ( .B1(n13554), .B2(n13206), .A(n13197), .ZN(n13198) );
  OAI21_X1 U14855 ( .B1(n13199), .B2(n13229), .A(n13198), .ZN(P3_U3173) );
  INV_X1 U14856 ( .A(n13200), .ZN(n13201) );
  AOI21_X1 U14857 ( .B1(n13509), .B2(n13202), .A(n13201), .ZN(n13208) );
  AOI22_X1 U14858 ( .A1(n13247), .A2(n13223), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13204) );
  NAND2_X1 U14859 ( .A1(n13239), .A2(n13526), .ZN(n13203) );
  OAI211_X1 U14860 ( .C1(n13522), .C2(n13225), .A(n13204), .B(n13203), .ZN(
        n13205) );
  AOI21_X1 U14861 ( .B1(n13525), .B2(n13206), .A(n13205), .ZN(n13207) );
  OAI21_X1 U14862 ( .B1(n13208), .B2(n13229), .A(n13207), .ZN(P3_U3175) );
  INV_X1 U14863 ( .A(n13717), .ZN(n13583) );
  AOI21_X1 U14864 ( .B1(n13210), .B2(n13209), .A(n13229), .ZN(n13212) );
  NAND2_X1 U14865 ( .A1(n13212), .A2(n13211), .ZN(n13216) );
  NAND2_X1 U14866 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13388)
         );
  NAND2_X1 U14867 ( .A1(n13251), .A2(n13223), .ZN(n13213) );
  OAI211_X1 U14868 ( .C1(n13580), .C2(n13225), .A(n13388), .B(n13213), .ZN(
        n13214) );
  AOI21_X1 U14869 ( .B1(n13581), .B2(n13239), .A(n13214), .ZN(n13215) );
  OAI211_X1 U14870 ( .C1(n13583), .C2(n13242), .A(n13216), .B(n13215), .ZN(
        P3_U3178) );
  OAI21_X1 U14871 ( .B1(n13220), .B2(n13219), .A(n13218), .ZN(n13222) );
  NAND2_X1 U14872 ( .A1(n13222), .A2(n13221), .ZN(n13228) );
  AOI22_X1 U14873 ( .A1(n13245), .A2(n13223), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13224) );
  OAI21_X1 U14874 ( .B1(n13467), .B2(n13225), .A(n13224), .ZN(n13226) );
  AOI21_X1 U14875 ( .B1(n13472), .B2(n13239), .A(n13226), .ZN(n13227) );
  OAI211_X1 U14876 ( .C1(n13757), .C2(n13242), .A(n13228), .B(n13227), .ZN(
        P3_U3180) );
  AOI21_X1 U14877 ( .B1(n13231), .B2(n13230), .A(n13229), .ZN(n13233) );
  NAND2_X1 U14878 ( .A1(n13233), .A2(n13232), .ZN(n13241) );
  NOR2_X1 U14879 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13234), .ZN(n13316) );
  AOI21_X1 U14880 ( .B1(n13626), .B2(n13235), .A(n13316), .ZN(n13236) );
  OAI21_X1 U14881 ( .B1(n13656), .B2(n13237), .A(n13236), .ZN(n13238) );
  AOI21_X1 U14882 ( .B1(n13630), .B2(n13239), .A(n13238), .ZN(n13240) );
  OAI211_X1 U14883 ( .C1(n13242), .C2(n13789), .A(n13241), .B(n13240), .ZN(
        P3_U3181) );
  MUX2_X1 U14884 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n13243), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14885 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13244), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14886 ( .A(n13483), .B(P3_DATAO_REG_26__SCAN_IN), .S(n13263), .Z(
        P3_U3517) );
  MUX2_X1 U14887 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n13245), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14888 ( .A(n13508), .B(P3_DATAO_REG_24__SCAN_IN), .S(n13263), .Z(
        P3_U3515) );
  MUX2_X1 U14889 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n13246), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14890 ( .A(n13509), .B(P3_DATAO_REG_22__SCAN_IN), .S(n13263), .Z(
        P3_U3513) );
  MUX2_X1 U14891 ( .A(n13247), .B(P3_DATAO_REG_21__SCAN_IN), .S(n13263), .Z(
        P3_U3512) );
  MUX2_X1 U14892 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13248), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14893 ( .A(n13249), .B(P3_DATAO_REG_19__SCAN_IN), .S(n13263), .Z(
        P3_U3510) );
  MUX2_X1 U14894 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13250), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14895 ( .A(n13251), .B(P3_DATAO_REG_17__SCAN_IN), .S(n13263), .Z(
        P3_U3508) );
  MUX2_X1 U14896 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13626), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14897 ( .A(n13641), .B(P3_DATAO_REG_15__SCAN_IN), .S(n13263), .Z(
        P3_U3506) );
  MUX2_X1 U14898 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n13627), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14899 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n13644), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14900 ( .A(n13252), .B(P3_DATAO_REG_12__SCAN_IN), .S(n13263), .Z(
        P3_U3503) );
  MUX2_X1 U14901 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n13253), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14902 ( .A(n13254), .B(P3_DATAO_REG_10__SCAN_IN), .S(n13263), .Z(
        P3_U3501) );
  MUX2_X1 U14903 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n7907), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14904 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n13255), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14905 ( .A(n13256), .B(P3_DATAO_REG_7__SCAN_IN), .S(n13263), .Z(
        P3_U3498) );
  MUX2_X1 U14906 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13257), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14907 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13258), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14908 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n13259), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14909 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n13260), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14910 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13261), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14911 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n13262), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14912 ( .A(n13264), .B(P3_DATAO_REG_0__SCAN_IN), .S(n13263), .Z(
        P3_U3491) );
  INV_X1 U14913 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13267) );
  INV_X1 U14914 ( .A(n13299), .ZN(n13287) );
  AOI21_X1 U14915 ( .B1(n13267), .B2(n13266), .A(n13288), .ZN(n13285) );
  NAND2_X1 U14916 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n13270), .ZN(n13293) );
  OAI21_X1 U14917 ( .B1(n13270), .B2(P3_REG1_REG_13__SCAN_IN), .A(n13293), 
        .ZN(n13271) );
  INV_X1 U14918 ( .A(n13271), .ZN(n13274) );
  NAND2_X1 U14919 ( .A1(n15663), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n13273) );
  OAI211_X1 U14920 ( .C1(n15583), .C2(n13274), .A(n13273), .B(n13272), .ZN(
        n13275) );
  AOI21_X1 U14921 ( .B1(n13287), .B2(n15602), .A(n13275), .ZN(n13284) );
  NAND2_X1 U14922 ( .A1(n13277), .A2(n13276), .ZN(n13278) );
  MUX2_X1 U14923 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13408), .Z(n13300) );
  XNOR2_X1 U14924 ( .A(n13300), .B(n13287), .ZN(n13279) );
  AOI21_X1 U14925 ( .B1(n13281), .B2(n13278), .A(n13279), .ZN(n13282) );
  AND2_X1 U14926 ( .A1(n13279), .A2(n13278), .ZN(n13280) );
  OAI21_X1 U14927 ( .B1(n13282), .B2(n13302), .A(n13412), .ZN(n13283) );
  OAI211_X1 U14928 ( .C1(n13285), .C2(n15671), .A(n13284), .B(n13283), .ZN(
        P3_U3195) );
  NOR2_X1 U14929 ( .A1(n13287), .A2(n13286), .ZN(n13289) );
  NAND2_X1 U14930 ( .A1(P3_REG2_REG_14__SCAN_IN), .A2(n13321), .ZN(n13290) );
  OAI21_X1 U14931 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n13321), .A(n13290), 
        .ZN(n13291) );
  AOI21_X1 U14932 ( .B1(n7343), .B2(n13291), .A(n13310), .ZN(n13309) );
  NAND2_X1 U14933 ( .A1(n13299), .A2(n13292), .ZN(n13294) );
  NAND2_X1 U14934 ( .A1(n13294), .A2(n13293), .ZN(n13296) );
  INV_X1 U14935 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13736) );
  XNOR2_X1 U14936 ( .A(n13321), .B(n13736), .ZN(n13295) );
  NAND2_X1 U14937 ( .A1(n13295), .A2(n13296), .ZN(n13313) );
  OAI21_X1 U14938 ( .B1(n13296), .B2(n13295), .A(n13313), .ZN(n13307) );
  NAND2_X1 U14939 ( .A1(n15663), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n13297) );
  OAI211_X1 U14940 ( .C1(n15657), .C2(n13321), .A(n13298), .B(n13297), .ZN(
        n13306) );
  MUX2_X1 U14941 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n13408), .Z(n13322) );
  XNOR2_X1 U14942 ( .A(n13322), .B(n13321), .ZN(n13304) );
  NOR2_X1 U14943 ( .A1(n13300), .A2(n13299), .ZN(n13301) );
  OR2_X1 U14944 ( .A1(n13302), .A2(n13301), .ZN(n13303) );
  AOI211_X1 U14945 ( .C1(n13304), .C2(n13303), .A(n15659), .B(n13320), .ZN(
        n13305) );
  AOI211_X1 U14946 ( .C1(n15667), .C2(n13307), .A(n13306), .B(n13305), .ZN(
        n13308) );
  OAI21_X1 U14947 ( .B1(n13309), .B2(n15671), .A(n13308), .ZN(P3_U3196) );
  INV_X1 U14948 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13312) );
  INV_X1 U14949 ( .A(n13340), .ZN(n13337) );
  XNOR2_X1 U14950 ( .A(n13328), .B(n13337), .ZN(n13311) );
  AOI21_X1 U14951 ( .B1(n13312), .B2(n13311), .A(n13329), .ZN(n13327) );
  NAND2_X1 U14952 ( .A1(P3_REG1_REG_14__SCAN_IN), .A2(n13321), .ZN(n13314) );
  OAI21_X1 U14953 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n13315), .A(n13341), 
        .ZN(n13319) );
  AOI21_X1 U14954 ( .B1(n15663), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n13316), 
        .ZN(n13317) );
  OAI21_X1 U14955 ( .B1(n15657), .B2(n13340), .A(n13317), .ZN(n13318) );
  AOI21_X1 U14956 ( .B1(n13319), .B2(n15667), .A(n13318), .ZN(n13326) );
  AOI21_X1 U14957 ( .B1(n13322), .B2(n13321), .A(n13320), .ZN(n13336) );
  XNOR2_X1 U14958 ( .A(n13336), .B(n13340), .ZN(n13324) );
  MUX2_X1 U14959 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n13408), .Z(n13323) );
  NAND2_X1 U14960 ( .A1(n13324), .A2(n13323), .ZN(n13335) );
  OAI211_X1 U14961 ( .C1(n13324), .C2(n13323), .A(n13335), .B(n13412), .ZN(
        n13325) );
  OAI211_X1 U14962 ( .C1(n13327), .C2(n15671), .A(n13326), .B(n13325), .ZN(
        P3_U3197) );
  NOR2_X1 U14963 ( .A1(n13337), .A2(n13328), .ZN(n13330) );
  INV_X1 U14964 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13331) );
  NOR2_X1 U14965 ( .A1(n13348), .A2(n13331), .ZN(n13363) );
  INV_X1 U14966 ( .A(n13363), .ZN(n13332) );
  OAI21_X1 U14967 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n13372), .A(n13332), 
        .ZN(n13333) );
  AOI21_X1 U14968 ( .B1(n7282), .B2(n13333), .A(n13362), .ZN(n13354) );
  MUX2_X1 U14969 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n13408), .Z(n13371) );
  NOR2_X1 U14970 ( .A1(n13371), .A2(n13372), .ZN(n13373) );
  INV_X1 U14971 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13343) );
  NOR2_X1 U14972 ( .A1(n13348), .A2(n13343), .ZN(n13355) );
  MUX2_X1 U14973 ( .A(n13363), .B(n13355), .S(n13408), .Z(n13334) );
  NOR2_X1 U14974 ( .A1(n13373), .A2(n13334), .ZN(n13338) );
  OAI21_X1 U14975 ( .B1(n13337), .B2(n13336), .A(n13335), .ZN(n13370) );
  XOR2_X1 U14976 ( .A(n13338), .B(n13370), .Z(n13352) );
  NAND2_X1 U14977 ( .A1(n13340), .A2(n13339), .ZN(n13342) );
  NAND2_X1 U14978 ( .A1(n13348), .A2(n13343), .ZN(n13356) );
  OAI21_X1 U14979 ( .B1(n13348), .B2(n13343), .A(n13356), .ZN(n13344) );
  XNOR2_X1 U14980 ( .A(n13357), .B(n13344), .ZN(n13350) );
  INV_X1 U14981 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n13346) );
  OAI21_X1 U14982 ( .B1(n15593), .B2(n13346), .A(n13345), .ZN(n13347) );
  AOI21_X1 U14983 ( .B1(n13348), .B2(n15602), .A(n13347), .ZN(n13349) );
  OAI21_X1 U14984 ( .B1(n13350), .B2(n15583), .A(n13349), .ZN(n13351) );
  AOI21_X1 U14985 ( .B1(n13412), .B2(n13352), .A(n13351), .ZN(n13353) );
  OAI21_X1 U14986 ( .B1(n13354), .B2(n15671), .A(n13353), .ZN(P3_U3198) );
  AOI21_X1 U14987 ( .B1(n13357), .B2(n13356), .A(n13355), .ZN(n13359) );
  INV_X1 U14988 ( .A(n13379), .ZN(n13358) );
  OAI21_X1 U14989 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n13360), .A(n13395), 
        .ZN(n13377) );
  AOI21_X1 U14990 ( .B1(n15663), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n13361), 
        .ZN(n13369) );
  OR2_X1 U14991 ( .A1(n13364), .A2(n13379), .ZN(n13365) );
  OAI21_X1 U14992 ( .B1(P3_REG2_REG_17__SCAN_IN), .B2(n13366), .A(n13386), 
        .ZN(n13367) );
  MUX2_X1 U14993 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13408), .Z(n13380) );
  XNOR2_X1 U14994 ( .A(n13380), .B(n13379), .ZN(n13375) );
  NOR2_X1 U14995 ( .A1(n13374), .A2(n13375), .ZN(n13378) );
  AOI211_X1 U14996 ( .C1(n13375), .C2(n13374), .A(n15659), .B(n13378), .ZN(
        n13376) );
  MUX2_X1 U14997 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13408), .Z(n13382) );
  AOI21_X1 U14998 ( .B1(n13380), .B2(n13379), .A(n13378), .ZN(n13406) );
  XNOR2_X1 U14999 ( .A(n13406), .B(n13405), .ZN(n13381) );
  NOR2_X1 U15000 ( .A1(n13381), .A2(n13382), .ZN(n13404) );
  AOI21_X1 U15001 ( .B1(n13382), .B2(n13381), .A(n13404), .ZN(n13399) );
  INV_X1 U15002 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13383) );
  OR2_X1 U15003 ( .A1(n13405), .A2(n13383), .ZN(n13414) );
  NAND2_X1 U15004 ( .A1(n13405), .A2(n13383), .ZN(n13384) );
  NAND3_X1 U15005 ( .A1(n13386), .A2(n13385), .A3(n7359), .ZN(n13387) );
  AND2_X1 U15006 ( .A1(n13415), .A2(n13387), .ZN(n13390) );
  NAND2_X1 U15007 ( .A1(n15663), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n13389) );
  OAI211_X1 U15008 ( .C1(n15671), .C2(n13390), .A(n13389), .B(n13388), .ZN(
        n13391) );
  AOI21_X1 U15009 ( .B1(n13405), .B2(n15602), .A(n13391), .ZN(n13398) );
  INV_X1 U15010 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13392) );
  OR2_X1 U15011 ( .A1(n13405), .A2(n13392), .ZN(n13400) );
  NAND2_X1 U15012 ( .A1(n13405), .A2(n13392), .ZN(n13393) );
  NAND2_X1 U15013 ( .A1(n13400), .A2(n13393), .ZN(n13394) );
  AND3_X1 U15014 ( .A1(n13395), .A2(n7269), .A3(n13394), .ZN(n13396) );
  OAI21_X1 U15015 ( .B1(n13402), .B2(n13396), .A(n15667), .ZN(n13397) );
  OAI211_X1 U15016 ( .C1(n13399), .C2(n15659), .A(n13398), .B(n13397), .ZN(
        P3_U3200) );
  XNOR2_X1 U15017 ( .A(n13407), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13409) );
  INV_X1 U15018 ( .A(n13400), .ZN(n13401) );
  NOR2_X1 U15019 ( .A1(n13402), .A2(n13401), .ZN(n13403) );
  XNOR2_X1 U15020 ( .A(n13407), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13416) );
  MUX2_X1 U15021 ( .A(n13416), .B(n13409), .S(n13408), .Z(n13410) );
  XNOR2_X1 U15022 ( .A(n13411), .B(n13410), .ZN(n13413) );
  NAND2_X1 U15023 ( .A1(n13413), .A2(n13412), .ZN(n13420) );
  NAND2_X1 U15024 ( .A1(n13415), .A2(n13414), .ZN(n13417) );
  NOR2_X1 U15025 ( .A1(n13423), .A2(n13422), .ZN(n13743) );
  NOR2_X1 U15026 ( .A1(n15727), .A2(n13424), .ZN(n13432) );
  NOR3_X1 U15027 ( .A1(n13743), .A2(n13670), .A3(n13432), .ZN(n13427) );
  NOR2_X1 U15028 ( .A1(n15735), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13425) );
  OAI22_X1 U15029 ( .A1(n13745), .A2(n13650), .B1(n13427), .B2(n13425), .ZN(
        P3_U3202) );
  NOR2_X1 U15030 ( .A1(n15735), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13426) );
  OAI22_X1 U15031 ( .A1(n13748), .A2(n13650), .B1(n13427), .B2(n13426), .ZN(
        P3_U3203) );
  INV_X1 U15032 ( .A(n13428), .ZN(n13435) );
  NAND2_X1 U15033 ( .A1(n13429), .A2(n15735), .ZN(n13434) );
  NOR2_X1 U15034 ( .A1(n13430), .A2(n13650), .ZN(n13431) );
  AOI211_X1 U15035 ( .C1(n13670), .C2(P3_REG2_REG_29__SCAN_IN), .A(n13432), 
        .B(n13431), .ZN(n13433) );
  OAI211_X1 U15036 ( .C1(n13435), .C2(n13653), .A(n13434), .B(n13433), .ZN(
        P3_U3204) );
  OAI211_X1 U15037 ( .C1(n13438), .C2(n13437), .A(n13436), .B(n13640), .ZN(
        n13442) );
  OAI22_X1 U15038 ( .A1(n13439), .A2(n15723), .B1(n13467), .B2(n15721), .ZN(
        n13440) );
  INV_X1 U15039 ( .A(n13440), .ZN(n13441) );
  XNOR2_X1 U15040 ( .A(n13443), .B(n7769), .ZN(n13674) );
  AOI22_X1 U15041 ( .A1(n13670), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n13648), 
        .B2(n13444), .ZN(n13445) );
  OAI21_X1 U15042 ( .B1(n13752), .B2(n13650), .A(n13445), .ZN(n13446) );
  AOI21_X1 U15043 ( .B1(n13674), .B2(n13667), .A(n13446), .ZN(n13447) );
  OAI21_X1 U15044 ( .B1(n13676), .B2(n13670), .A(n13447), .ZN(P3_U3205) );
  XNOR2_X1 U15045 ( .A(n13448), .B(n13454), .ZN(n13682) );
  NAND2_X1 U15046 ( .A1(n13452), .A2(n13450), .ZN(n13453) );
  AOI21_X1 U15047 ( .B1(n13454), .B2(n13453), .A(n8260), .ZN(n13455) );
  OAI222_X1 U15048 ( .A1(n15721), .A2(n13457), .B1(n15723), .B2(n13456), .C1(
        n15719), .C2(n13455), .ZN(n13679) );
  NAND2_X1 U15049 ( .A1(n13679), .A2(n15735), .ZN(n13463) );
  INV_X1 U15050 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n13460) );
  INV_X1 U15051 ( .A(n13458), .ZN(n13459) );
  OAI22_X1 U15052 ( .A1(n15735), .A2(n13460), .B1(n13459), .B2(n15727), .ZN(
        n13461) );
  AOI21_X1 U15053 ( .B1(n13680), .B2(n13663), .A(n13461), .ZN(n13462) );
  OAI211_X1 U15054 ( .C1(n13682), .C2(n13653), .A(n13463), .B(n13462), .ZN(
        P3_U3206) );
  XNOR2_X1 U15055 ( .A(n13465), .B(n13471), .ZN(n13466) );
  OAI222_X1 U15056 ( .A1(n15723), .A2(n13467), .B1(n15721), .B2(n13495), .C1(
        n13466), .C2(n15719), .ZN(n13683) );
  INV_X1 U15057 ( .A(n13683), .ZN(n13476) );
  NAND2_X1 U15058 ( .A1(n13469), .A2(n13468), .ZN(n13470) );
  XOR2_X1 U15059 ( .A(n13471), .B(n13470), .Z(n13684) );
  AOI22_X1 U15060 ( .A1(n13670), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n13472), 
        .B2(n13648), .ZN(n13473) );
  OAI21_X1 U15061 ( .B1(n13757), .B2(n13650), .A(n13473), .ZN(n13474) );
  AOI21_X1 U15062 ( .B1(n13684), .B2(n13667), .A(n13474), .ZN(n13475) );
  OAI21_X1 U15063 ( .B1(n13476), .B2(n13670), .A(n13475), .ZN(P3_U3207) );
  XNOR2_X1 U15064 ( .A(n13477), .B(n13478), .ZN(n13690) );
  INV_X1 U15065 ( .A(n13479), .ZN(n13482) );
  OAI211_X1 U15066 ( .C1(n13482), .C2(n13481), .A(n13480), .B(n13640), .ZN(
        n13485) );
  NAND2_X1 U15067 ( .A1(n13483), .A2(n13642), .ZN(n13484) );
  OAI211_X1 U15068 ( .C1(n13486), .C2(n15721), .A(n13485), .B(n13484), .ZN(
        n13687) );
  AOI22_X1 U15069 ( .A1(n13670), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n13648), 
        .B2(n13487), .ZN(n13488) );
  OAI21_X1 U15070 ( .B1(n13489), .B2(n13650), .A(n13488), .ZN(n13490) );
  AOI21_X1 U15071 ( .B1(n13687), .B2(n15735), .A(n13490), .ZN(n13491) );
  OAI21_X1 U15072 ( .B1(n13690), .B2(n13653), .A(n13491), .ZN(P3_U3208) );
  XNOR2_X1 U15073 ( .A(n13492), .B(n13493), .ZN(n13499) );
  XNOR2_X1 U15074 ( .A(n13494), .B(n13493), .ZN(n13497) );
  OAI22_X1 U15075 ( .A1(n13522), .A2(n15721), .B1(n13495), .B2(n15723), .ZN(
        n13496) );
  AOI21_X1 U15076 ( .B1(n13497), .B2(n13640), .A(n13496), .ZN(n13498) );
  OAI21_X1 U15077 ( .B1(n13552), .B2(n13499), .A(n13498), .ZN(n13691) );
  INV_X1 U15078 ( .A(n13691), .ZN(n13504) );
  INV_X1 U15079 ( .A(n13499), .ZN(n13692) );
  AOI22_X1 U15080 ( .A1(n13670), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n13648), 
        .B2(n13500), .ZN(n13501) );
  OAI21_X1 U15081 ( .B1(n13762), .B2(n13650), .A(n13501), .ZN(n13502) );
  AOI21_X1 U15082 ( .B1(n13692), .B2(n13558), .A(n13502), .ZN(n13503) );
  OAI21_X1 U15083 ( .B1(n13504), .B2(n13670), .A(n13503), .ZN(P3_U3209) );
  XNOR2_X1 U15084 ( .A(n13506), .B(n13505), .ZN(n13507) );
  NAND2_X1 U15085 ( .A1(n13507), .A2(n13640), .ZN(n13511) );
  AOI22_X1 U15086 ( .A1(n13643), .A2(n13509), .B1(n13508), .B2(n13642), .ZN(
        n13510) );
  NAND2_X1 U15087 ( .A1(n13511), .A2(n13510), .ZN(n13697) );
  INV_X1 U15088 ( .A(n13697), .ZN(n13519) );
  XNOR2_X1 U15089 ( .A(n13512), .B(n13513), .ZN(n13695) );
  INV_X1 U15090 ( .A(n13514), .ZN(n13766) );
  AOI22_X1 U15091 ( .A1(n13670), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n13648), 
        .B2(n13515), .ZN(n13516) );
  OAI21_X1 U15092 ( .B1(n13766), .B2(n13650), .A(n13516), .ZN(n13517) );
  AOI21_X1 U15093 ( .B1(n13695), .B2(n13667), .A(n13517), .ZN(n13518) );
  OAI21_X1 U15094 ( .B1(n13519), .B2(n13670), .A(n13518), .ZN(P3_U3210) );
  XNOR2_X1 U15095 ( .A(n13520), .B(n13524), .ZN(n13521) );
  OAI222_X1 U15096 ( .A1(n15721), .A2(n13548), .B1(n15723), .B2(n13522), .C1(
        n13521), .C2(n15719), .ZN(n13700) );
  INV_X1 U15097 ( .A(n13700), .ZN(n13530) );
  XOR2_X1 U15098 ( .A(n13524), .B(n13523), .Z(n13701) );
  INV_X1 U15099 ( .A(n13525), .ZN(n13770) );
  AOI22_X1 U15100 ( .A1(n13670), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n13648), 
        .B2(n13526), .ZN(n13527) );
  OAI21_X1 U15101 ( .B1(n13770), .B2(n13650), .A(n13527), .ZN(n13528) );
  AOI21_X1 U15102 ( .B1(n13701), .B2(n13667), .A(n13528), .ZN(n13529) );
  OAI21_X1 U15103 ( .B1(n13530), .B2(n13670), .A(n13529), .ZN(P3_U3211) );
  XNOR2_X1 U15104 ( .A(n13531), .B(n13532), .ZN(n13538) );
  XNOR2_X1 U15105 ( .A(n13533), .B(n13532), .ZN(n13536) );
  OAI22_X1 U15106 ( .A1(n13534), .A2(n15723), .B1(n13568), .B2(n15721), .ZN(
        n13535) );
  AOI21_X1 U15107 ( .B1(n13536), .B2(n13640), .A(n13535), .ZN(n13537) );
  OAI21_X1 U15108 ( .B1(n13552), .B2(n13538), .A(n13537), .ZN(n13704) );
  INV_X1 U15109 ( .A(n13704), .ZN(n13544) );
  INV_X1 U15110 ( .A(n13538), .ZN(n13705) );
  INV_X1 U15111 ( .A(n13539), .ZN(n13774) );
  AOI22_X1 U15112 ( .A1(n13670), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n13648), 
        .B2(n13540), .ZN(n13541) );
  OAI21_X1 U15113 ( .B1(n13774), .B2(n13650), .A(n13541), .ZN(n13542) );
  AOI21_X1 U15114 ( .B1(n13705), .B2(n13558), .A(n13542), .ZN(n13543) );
  OAI21_X1 U15115 ( .B1(n13544), .B2(n13670), .A(n13543), .ZN(P3_U3212) );
  XNOR2_X1 U15116 ( .A(n13545), .B(n13546), .ZN(n13553) );
  XNOR2_X1 U15117 ( .A(n13547), .B(n13546), .ZN(n13550) );
  OAI22_X1 U15118 ( .A1(n13580), .A2(n15721), .B1(n13548), .B2(n15723), .ZN(
        n13549) );
  AOI21_X1 U15119 ( .B1(n13550), .B2(n13640), .A(n13549), .ZN(n13551) );
  OAI21_X1 U15120 ( .B1(n13552), .B2(n13553), .A(n13551), .ZN(n13708) );
  INV_X1 U15121 ( .A(n13708), .ZN(n13560) );
  INV_X1 U15122 ( .A(n13553), .ZN(n13709) );
  INV_X1 U15123 ( .A(n13554), .ZN(n13778) );
  AOI22_X1 U15124 ( .A1(n13670), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n13648), 
        .B2(n13555), .ZN(n13556) );
  OAI21_X1 U15125 ( .B1(n13778), .B2(n13650), .A(n13556), .ZN(n13557) );
  AOI21_X1 U15126 ( .B1(n13709), .B2(n13558), .A(n13557), .ZN(n13559) );
  OAI21_X1 U15127 ( .B1(n13560), .B2(n13670), .A(n13559), .ZN(P3_U3213) );
  INV_X1 U15128 ( .A(n13602), .ZN(n13563) );
  OAI21_X1 U15129 ( .B1(n13563), .B2(n13562), .A(n13561), .ZN(n13564) );
  XOR2_X1 U15130 ( .A(n13565), .B(n13564), .Z(n13715) );
  XOR2_X1 U15131 ( .A(n13566), .B(n13565), .Z(n13567) );
  OAI222_X1 U15132 ( .A1(n15723), .A2(n13568), .B1(n15721), .B2(n13590), .C1(
        n15719), .C2(n13567), .ZN(n13712) );
  NAND2_X1 U15133 ( .A1(n13712), .A2(n15735), .ZN(n13574) );
  INV_X1 U15134 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13571) );
  INV_X1 U15135 ( .A(n13569), .ZN(n13570) );
  OAI22_X1 U15136 ( .A1(n15735), .A2(n13571), .B1(n13570), .B2(n15727), .ZN(
        n13572) );
  AOI21_X1 U15137 ( .B1(n13713), .B2(n13663), .A(n13572), .ZN(n13573) );
  OAI211_X1 U15138 ( .C1(n13715), .C2(n13653), .A(n13574), .B(n13573), .ZN(
        P3_U3214) );
  NAND2_X1 U15139 ( .A1(n13602), .A2(n13575), .ZN(n13576) );
  XOR2_X1 U15140 ( .A(n13578), .B(n13576), .Z(n13719) );
  AOI21_X1 U15141 ( .B1(n13578), .B2(n13577), .A(n7344), .ZN(n13579) );
  OAI222_X1 U15142 ( .A1(n15723), .A2(n13580), .B1(n15721), .B2(n13614), .C1(
        n15719), .C2(n13579), .ZN(n13716) );
  AOI22_X1 U15143 ( .A1(n13670), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n13648), 
        .B2(n13581), .ZN(n13582) );
  OAI21_X1 U15144 ( .B1(n13583), .B2(n13650), .A(n13582), .ZN(n13584) );
  AOI21_X1 U15145 ( .B1(n13716), .B2(n15735), .A(n13584), .ZN(n13585) );
  OAI21_X1 U15146 ( .B1(n13653), .B2(n13719), .A(n13585), .ZN(P3_U3215) );
  NAND2_X1 U15147 ( .A1(n13608), .A2(n13586), .ZN(n13587) );
  NAND2_X1 U15148 ( .A1(n13587), .A2(n13599), .ZN(n13589) );
  NAND3_X1 U15149 ( .A1(n13589), .A2(n13640), .A3(n13588), .ZN(n13594) );
  OAI22_X1 U15150 ( .A1(n13591), .A2(n15721), .B1(n13590), .B2(n15723), .ZN(
        n13592) );
  INV_X1 U15151 ( .A(n13592), .ZN(n13593) );
  INV_X1 U15152 ( .A(n13595), .ZN(n13596) );
  OAI22_X1 U15153 ( .A1(n15735), .A2(n7952), .B1(n13596), .B2(n15727), .ZN(
        n13597) );
  AOI21_X1 U15154 ( .B1(n13598), .B2(n13663), .A(n13597), .ZN(n13604) );
  OR2_X1 U15155 ( .A1(n13600), .A2(n13599), .ZN(n13601) );
  NAND2_X1 U15156 ( .A1(n13602), .A2(n13601), .ZN(n13720) );
  NAND2_X1 U15157 ( .A1(n13720), .A2(n13667), .ZN(n13603) );
  OAI211_X1 U15158 ( .C1(n13721), .C2(n13670), .A(n13604), .B(n13603), .ZN(
        P3_U3216) );
  XOR2_X1 U15159 ( .A(n13611), .B(n13605), .Z(n13728) );
  NAND2_X1 U15160 ( .A1(n13606), .A2(n13607), .ZN(n13610) );
  INV_X1 U15161 ( .A(n13608), .ZN(n13609) );
  AOI21_X1 U15162 ( .B1(n13611), .B2(n13610), .A(n13609), .ZN(n13612) );
  OAI222_X1 U15163 ( .A1(n15723), .A2(n13614), .B1(n15721), .B2(n13613), .C1(
        n15719), .C2(n13612), .ZN(n13725) );
  AOI22_X1 U15164 ( .A1(n13670), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n13648), 
        .B2(n13615), .ZN(n13616) );
  OAI21_X1 U15165 ( .B1(n13617), .B2(n13650), .A(n13616), .ZN(n13618) );
  AOI21_X1 U15166 ( .B1(n13725), .B2(n15735), .A(n13618), .ZN(n13619) );
  OAI21_X1 U15167 ( .B1(n13653), .B2(n13728), .A(n13619), .ZN(P3_U3217) );
  OAI21_X1 U15168 ( .B1(n13621), .B2(n13624), .A(n13620), .ZN(n13731) );
  INV_X1 U15169 ( .A(n13731), .ZN(n13634) );
  NAND3_X1 U15170 ( .A1(n13622), .A2(n13624), .A3(n13623), .ZN(n13625) );
  NAND3_X1 U15171 ( .A1(n13606), .A2(n13640), .A3(n13625), .ZN(n13629) );
  AOI22_X1 U15172 ( .A1(n13643), .A2(n13627), .B1(n13626), .B2(n13642), .ZN(
        n13628) );
  NAND2_X1 U15173 ( .A1(n13629), .A2(n13628), .ZN(n13730) );
  AOI22_X1 U15174 ( .A1(n13670), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n13630), 
        .B2(n13648), .ZN(n13631) );
  OAI21_X1 U15175 ( .B1(n13789), .B2(n13650), .A(n13631), .ZN(n13632) );
  AOI21_X1 U15176 ( .B1(n13730), .B2(n15735), .A(n13632), .ZN(n13633) );
  OAI21_X1 U15177 ( .B1(n13634), .B2(n13653), .A(n13633), .ZN(P3_U3218) );
  XNOR2_X1 U15178 ( .A(n13635), .B(n13638), .ZN(n13735) );
  INV_X1 U15179 ( .A(n13735), .ZN(n13654) );
  NAND3_X1 U15180 ( .A1(n13636), .A2(n13638), .A3(n13637), .ZN(n13639) );
  NAND3_X1 U15181 ( .A1(n13622), .A2(n13640), .A3(n13639), .ZN(n13646) );
  AOI22_X1 U15182 ( .A1(n13644), .A2(n13643), .B1(n13642), .B2(n13641), .ZN(
        n13645) );
  NAND2_X1 U15183 ( .A1(n13646), .A2(n13645), .ZN(n13734) );
  AOI22_X1 U15184 ( .A1(n13670), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n13648), 
        .B2(n13647), .ZN(n13649) );
  OAI21_X1 U15185 ( .B1(n13793), .B2(n13650), .A(n13649), .ZN(n13651) );
  AOI21_X1 U15186 ( .B1(n13734), .B2(n15735), .A(n13651), .ZN(n13652) );
  OAI21_X1 U15187 ( .B1(n13654), .B2(n13653), .A(n13652), .ZN(P3_U3219) );
  AOI21_X1 U15188 ( .B1(n13655), .B2(n13665), .A(n15719), .ZN(n13659) );
  OAI22_X1 U15189 ( .A1(n13657), .A2(n15721), .B1(n13656), .B2(n15723), .ZN(
        n13658) );
  AOI21_X1 U15190 ( .B1(n13659), .B2(n13636), .A(n13658), .ZN(n13740) );
  INV_X1 U15191 ( .A(n13660), .ZN(n13661) );
  OAI22_X1 U15192 ( .A1(n15735), .A2(n13267), .B1(n13661), .B2(n15727), .ZN(
        n13662) );
  AOI21_X1 U15193 ( .B1(n13664), .B2(n13663), .A(n13662), .ZN(n13669) );
  XNOR2_X1 U15194 ( .A(n13666), .B(n13665), .ZN(n13739) );
  NAND2_X1 U15195 ( .A1(n13739), .A2(n13667), .ZN(n13668) );
  OAI211_X1 U15196 ( .C1(n13740), .C2(n13670), .A(n13669), .B(n13668), .ZN(
        P3_U3220) );
  NAND2_X1 U15197 ( .A1(n15939), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13671) );
  NAND2_X1 U15198 ( .A1(n13743), .A2(n15940), .ZN(n13673) );
  OAI211_X1 U15199 ( .C1(n13745), .C2(n13738), .A(n13671), .B(n13673), .ZN(
        P3_U3490) );
  NAND2_X1 U15200 ( .A1(n15939), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13672) );
  OAI211_X1 U15201 ( .C1(n13748), .C2(n13738), .A(n13673), .B(n13672), .ZN(
        P3_U3489) );
  NAND2_X1 U15202 ( .A1(n13674), .A2(n15912), .ZN(n13675) );
  NAND2_X1 U15203 ( .A1(n13676), .A2(n13675), .ZN(n13749) );
  MUX2_X1 U15204 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n13749), .S(n15940), .Z(
        n13677) );
  INV_X1 U15205 ( .A(n13677), .ZN(n13678) );
  OAI21_X1 U15206 ( .B1(n13752), .B2(n13738), .A(n13678), .ZN(P3_U3487) );
  OAI21_X1 U15207 ( .B1(n13729), .B2(n13682), .A(n13681), .ZN(n13753) );
  MUX2_X1 U15208 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13753), .S(n15940), .Z(
        P3_U3486) );
  INV_X1 U15209 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13685) );
  AOI21_X1 U15210 ( .B1(n13684), .B2(n15912), .A(n13683), .ZN(n13754) );
  OAI21_X1 U15211 ( .B1(n13757), .B2(n13738), .A(n13686), .ZN(P3_U3485) );
  AOI21_X1 U15212 ( .B1(n15891), .B2(n13688), .A(n13687), .ZN(n13689) );
  OAI21_X1 U15213 ( .B1(n13729), .B2(n13690), .A(n13689), .ZN(n13758) );
  MUX2_X1 U15214 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13758), .S(n15940), .Z(
        P3_U3484) );
  INV_X1 U15215 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13693) );
  AOI21_X1 U15216 ( .B1(n15931), .B2(n13692), .A(n13691), .ZN(n13759) );
  MUX2_X1 U15217 ( .A(n13693), .B(n13759), .S(n15940), .Z(n13694) );
  OAI21_X1 U15218 ( .B1(n13762), .B2(n13738), .A(n13694), .ZN(P3_U3483) );
  INV_X1 U15219 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13698) );
  AND2_X1 U15220 ( .A1(n13695), .A2(n15912), .ZN(n13696) );
  NOR2_X1 U15221 ( .A1(n13697), .A2(n13696), .ZN(n13763) );
  MUX2_X1 U15222 ( .A(n13698), .B(n13763), .S(n15940), .Z(n13699) );
  OAI21_X1 U15223 ( .B1(n13766), .B2(n13738), .A(n13699), .ZN(P3_U3482) );
  INV_X1 U15224 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13702) );
  AOI21_X1 U15225 ( .B1(n13701), .B2(n15912), .A(n13700), .ZN(n13767) );
  MUX2_X1 U15226 ( .A(n13702), .B(n13767), .S(n15940), .Z(n13703) );
  OAI21_X1 U15227 ( .B1(n13770), .B2(n13738), .A(n13703), .ZN(P3_U3481) );
  INV_X1 U15228 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13706) );
  AOI21_X1 U15229 ( .B1(n15931), .B2(n13705), .A(n13704), .ZN(n13771) );
  MUX2_X1 U15230 ( .A(n13706), .B(n13771), .S(n15940), .Z(n13707) );
  OAI21_X1 U15231 ( .B1(n13774), .B2(n13738), .A(n13707), .ZN(P3_U3480) );
  INV_X1 U15232 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13710) );
  AOI21_X1 U15233 ( .B1(n15931), .B2(n13709), .A(n13708), .ZN(n13775) );
  MUX2_X1 U15234 ( .A(n13710), .B(n13775), .S(n15940), .Z(n13711) );
  OAI21_X1 U15235 ( .B1(n13778), .B2(n13738), .A(n13711), .ZN(P3_U3479) );
  AOI21_X1 U15236 ( .B1(n15891), .B2(n13713), .A(n13712), .ZN(n13714) );
  OAI21_X1 U15237 ( .B1(n13729), .B2(n13715), .A(n13714), .ZN(n13779) );
  MUX2_X1 U15238 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n13779), .S(n15940), .Z(
        P3_U3478) );
  AOI21_X1 U15239 ( .B1(n15891), .B2(n13717), .A(n13716), .ZN(n13718) );
  OAI21_X1 U15240 ( .B1(n13729), .B2(n13719), .A(n13718), .ZN(n13780) );
  MUX2_X1 U15241 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n13780), .S(n15940), .Z(
        P3_U3477) );
  NAND2_X1 U15242 ( .A1(n13720), .A2(n15912), .ZN(n13722) );
  NAND2_X1 U15243 ( .A1(n13722), .A2(n13721), .ZN(n13781) );
  MUX2_X1 U15244 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13781), .S(n15940), .Z(
        n13723) );
  INV_X1 U15245 ( .A(n13723), .ZN(n13724) );
  OAI21_X1 U15246 ( .B1(n13738), .B2(n13784), .A(n13724), .ZN(P3_U3476) );
  AOI21_X1 U15247 ( .B1(n15891), .B2(n13726), .A(n13725), .ZN(n13727) );
  OAI21_X1 U15248 ( .B1(n13729), .B2(n13728), .A(n13727), .ZN(n13785) );
  MUX2_X1 U15249 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n13785), .S(n15940), .Z(
        P3_U3475) );
  INV_X1 U15250 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13732) );
  AOI21_X1 U15251 ( .B1(n15912), .B2(n13731), .A(n13730), .ZN(n13786) );
  MUX2_X1 U15252 ( .A(n13732), .B(n13786), .S(n15940), .Z(n13733) );
  OAI21_X1 U15253 ( .B1(n13738), .B2(n13789), .A(n13733), .ZN(P3_U3474) );
  AOI21_X1 U15254 ( .B1(n15912), .B2(n13735), .A(n13734), .ZN(n13790) );
  MUX2_X1 U15255 ( .A(n13736), .B(n13790), .S(n15940), .Z(n13737) );
  OAI21_X1 U15256 ( .B1(n13738), .B2(n13793), .A(n13737), .ZN(P3_U3473) );
  NAND2_X1 U15257 ( .A1(n13739), .A2(n15912), .ZN(n13741) );
  OAI211_X1 U15258 ( .C1(n15935), .C2(n13742), .A(n13741), .B(n13740), .ZN(
        n13795) );
  MUX2_X1 U15259 ( .A(P3_REG1_REG_13__SCAN_IN), .B(n13795), .S(n15940), .Z(
        P3_U3472) );
  NAND2_X1 U15260 ( .A1(n15941), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13744) );
  NAND2_X1 U15261 ( .A1(n13743), .A2(n15944), .ZN(n13747) );
  OAI211_X1 U15262 ( .C1(n13745), .C2(n13794), .A(n13744), .B(n13747), .ZN(
        P3_U3458) );
  NAND2_X1 U15263 ( .A1(n15941), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n13746) );
  OAI211_X1 U15264 ( .C1(n13748), .C2(n13794), .A(n13747), .B(n13746), .ZN(
        P3_U3457) );
  MUX2_X1 U15265 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n13749), .S(n15944), .Z(
        n13750) );
  INV_X1 U15266 ( .A(n13750), .ZN(n13751) );
  OAI21_X1 U15267 ( .B1(n13752), .B2(n13794), .A(n13751), .ZN(P3_U3455) );
  MUX2_X1 U15268 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n13753), .S(n15944), .Z(
        P3_U3454) );
  INV_X1 U15269 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13755) );
  OAI21_X1 U15270 ( .B1(n13757), .B2(n13794), .A(n13756), .ZN(P3_U3453) );
  MUX2_X1 U15271 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n13758), .S(n15944), .Z(
        P3_U3452) );
  INV_X1 U15272 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13760) );
  MUX2_X1 U15273 ( .A(n13760), .B(n13759), .S(n15944), .Z(n13761) );
  OAI21_X1 U15274 ( .B1(n13762), .B2(n13794), .A(n13761), .ZN(P3_U3451) );
  INV_X1 U15275 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13764) );
  MUX2_X1 U15276 ( .A(n13764), .B(n13763), .S(n15944), .Z(n13765) );
  OAI21_X1 U15277 ( .B1(n13766), .B2(n13794), .A(n13765), .ZN(P3_U3450) );
  INV_X1 U15278 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13768) );
  MUX2_X1 U15279 ( .A(n13768), .B(n13767), .S(n15944), .Z(n13769) );
  OAI21_X1 U15280 ( .B1(n13770), .B2(n13794), .A(n13769), .ZN(P3_U3449) );
  INV_X1 U15281 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13772) );
  MUX2_X1 U15282 ( .A(n13772), .B(n13771), .S(n15944), .Z(n13773) );
  OAI21_X1 U15283 ( .B1(n13774), .B2(n13794), .A(n13773), .ZN(P3_U3448) );
  INV_X1 U15284 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13776) );
  MUX2_X1 U15285 ( .A(n13776), .B(n13775), .S(n15944), .Z(n13777) );
  OAI21_X1 U15286 ( .B1(n13778), .B2(n13794), .A(n13777), .ZN(P3_U3447) );
  MUX2_X1 U15287 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n13779), .S(n15944), .Z(
        P3_U3446) );
  MUX2_X1 U15288 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n13780), .S(n15944), .Z(
        P3_U3444) );
  MUX2_X1 U15289 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13781), .S(n15944), .Z(
        n13782) );
  INV_X1 U15290 ( .A(n13782), .ZN(n13783) );
  OAI21_X1 U15291 ( .B1(n13794), .B2(n13784), .A(n13783), .ZN(P3_U3441) );
  MUX2_X1 U15292 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n13785), .S(n15944), .Z(
        P3_U3438) );
  INV_X1 U15293 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13787) );
  MUX2_X1 U15294 ( .A(n13787), .B(n13786), .S(n15944), .Z(n13788) );
  OAI21_X1 U15295 ( .B1(n13794), .B2(n13789), .A(n13788), .ZN(P3_U3435) );
  INV_X1 U15296 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13791) );
  MUX2_X1 U15297 ( .A(n13791), .B(n13790), .S(n15944), .Z(n13792) );
  OAI21_X1 U15298 ( .B1(n13794), .B2(n13793), .A(n13792), .ZN(P3_U3432) );
  MUX2_X1 U15299 ( .A(P3_REG0_REG_13__SCAN_IN), .B(n13795), .S(n15944), .Z(
        P3_U3429) );
  MUX2_X1 U15300 ( .A(P3_D_REG_1__SCAN_IN), .B(n13797), .S(n13796), .Z(
        P3_U3377) );
  NAND2_X1 U15301 ( .A1(n13799), .A2(n13798), .ZN(n13803) );
  OR4_X1 U15302 ( .A1(n13801), .A2(P3_IR_REG_30__SCAN_IN), .A3(n8554), .A4(
        P3_U3151), .ZN(n13802) );
  OAI211_X1 U15303 ( .C1(n13804), .C2(n13810), .A(n13803), .B(n13802), .ZN(
        P3_U3264) );
  INV_X1 U15304 ( .A(n13805), .ZN(n13806) );
  OAI222_X1 U15305 ( .A1(n13808), .A2(P3_U3151), .B1(n13810), .B2(n13807), 
        .C1(n12036), .C2(n13806), .ZN(P3_U3265) );
  INV_X1 U15306 ( .A(n13809), .ZN(n13813) );
  OAI222_X1 U15307 ( .A1(n12036), .A2(n13813), .B1(P3_U3151), .B2(n13812), 
        .C1(n13811), .C2(n13810), .ZN(P3_U3266) );
  MUX2_X1 U15308 ( .A(n13814), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  INV_X1 U15309 ( .A(n13815), .ZN(n13817) );
  XNOR2_X1 U15310 ( .A(n14471), .B(n13847), .ZN(n13821) );
  NAND2_X1 U15311 ( .A1(n14010), .A2(n12208), .ZN(n13820) );
  NAND2_X1 U15312 ( .A1(n13821), .A2(n13820), .ZN(n13822) );
  OAI21_X1 U15313 ( .B1(n13821), .B2(n13820), .A(n13822), .ZN(n13916) );
  AND2_X1 U15314 ( .A1(n14009), .A2(n14295), .ZN(n13824) );
  XNOR2_X1 U15315 ( .A(n14320), .B(n7532), .ZN(n13823) );
  NOR2_X1 U15316 ( .A1(n13823), .A2(n13824), .ZN(n13825) );
  AOI21_X1 U15317 ( .B1(n13824), .B2(n13823), .A(n13825), .ZN(n13937) );
  INV_X1 U15318 ( .A(n13825), .ZN(n13826) );
  NAND2_X1 U15319 ( .A1(n14008), .A2(n12208), .ZN(n13827) );
  XNOR2_X1 U15320 ( .A(n13829), .B(n13827), .ZN(n13985) );
  INV_X1 U15321 ( .A(n13827), .ZN(n13828) );
  NAND2_X1 U15322 ( .A1(n13829), .A2(n13828), .ZN(n13830) );
  XNOR2_X1 U15323 ( .A(n14461), .B(n7532), .ZN(n13832) );
  NAND2_X1 U15324 ( .A1(n14243), .A2(n12208), .ZN(n13831) );
  XNOR2_X1 U15325 ( .A(n13832), .B(n13831), .ZN(n13878) );
  INV_X1 U15326 ( .A(n13831), .ZN(n13833) );
  AND2_X1 U15327 ( .A1(n14263), .A2(n14208), .ZN(n13835) );
  XNOR2_X1 U15328 ( .A(n14396), .B(n7532), .ZN(n13834) );
  NOR2_X1 U15329 ( .A1(n13834), .A2(n13835), .ZN(n13836) );
  AOI21_X1 U15330 ( .B1(n13835), .B2(n13834), .A(n13836), .ZN(n13964) );
  INV_X1 U15331 ( .A(n13836), .ZN(n13837) );
  NAND2_X1 U15332 ( .A1(n13963), .A2(n13837), .ZN(n13899) );
  NAND2_X1 U15333 ( .A1(n14244), .A2(n12208), .ZN(n13838) );
  XNOR2_X1 U15334 ( .A(n14456), .B(n7532), .ZN(n13840) );
  XOR2_X1 U15335 ( .A(n13838), .B(n13840), .Z(n13898) );
  INV_X1 U15336 ( .A(n13838), .ZN(n13839) );
  NAND2_X1 U15337 ( .A1(n13840), .A2(n13839), .ZN(n13841) );
  XNOR2_X1 U15338 ( .A(n14212), .B(n7532), .ZN(n13842) );
  NOR2_X1 U15339 ( .A1(n14223), .A2(n11286), .ZN(n13975) );
  INV_X1 U15340 ( .A(n13842), .ZN(n13843) );
  NAND2_X1 U15341 ( .A1(n13844), .A2(n13843), .ZN(n13845) );
  XNOR2_X1 U15342 ( .A(n14193), .B(n13847), .ZN(n13849) );
  NAND2_X1 U15343 ( .A1(n14204), .A2(n12208), .ZN(n13871) );
  INV_X1 U15344 ( .A(n13848), .ZN(n13850) );
  NOR2_X1 U15345 ( .A1(n14188), .A2(n11286), .ZN(n13853) );
  XNOR2_X1 U15346 ( .A(n14372), .B(n7532), .ZN(n13852) );
  XOR2_X1 U15347 ( .A(n13853), .B(n13852), .Z(n13944) );
  INV_X1 U15348 ( .A(n13852), .ZN(n13854) );
  NAND2_X1 U15349 ( .A1(n13854), .A2(n13853), .ZN(n13855) );
  XNOR2_X1 U15350 ( .A(n14158), .B(n7188), .ZN(n13858) );
  NAND2_X1 U15351 ( .A1(n14169), .A2(n12208), .ZN(n13856) );
  INV_X1 U15352 ( .A(n13856), .ZN(n13857) );
  NAND2_X1 U15353 ( .A1(n13858), .A2(n13857), .ZN(n13859) );
  XNOR2_X1 U15354 ( .A(n14441), .B(n7188), .ZN(n13862) );
  NAND2_X1 U15355 ( .A1(n14113), .A2(n12208), .ZN(n13861) );
  OAI21_X1 U15356 ( .B1(n13862), .B2(n13861), .A(n13863), .ZN(n13993) );
  XNOR2_X1 U15357 ( .A(n14437), .B(n7532), .ZN(n13885) );
  NAND2_X1 U15358 ( .A1(n14101), .A2(n12208), .ZN(n13884) );
  XNOR2_X1 U15359 ( .A(n13885), .B(n13884), .ZN(n13886) );
  XNOR2_X1 U15360 ( .A(n13887), .B(n13886), .ZN(n13869) );
  OAI22_X1 U15361 ( .A1(n14123), .A2(n13995), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13864), .ZN(n13867) );
  OAI22_X1 U15362 ( .A1(n13865), .A2(n13998), .B1(n14151), .B2(n13997), .ZN(
        n13866) );
  AOI211_X1 U15363 ( .C1(n14122), .C2(n14001), .A(n13867), .B(n13866), .ZN(
        n13868) );
  OAI21_X1 U15364 ( .B1(n13869), .B2(n14003), .A(n13868), .ZN(P2_U3186) );
  OAI21_X1 U15365 ( .B1(n13872), .B2(n13871), .A(n13870), .ZN(n13873) );
  NAND2_X1 U15366 ( .A1(n13873), .A2(n13966), .ZN(n13877) );
  NOR2_X1 U15367 ( .A1(n13995), .A2(n14197), .ZN(n13875) );
  OAI22_X1 U15368 ( .A1(n14223), .A2(n13997), .B1(n13998), .B2(n14188), .ZN(
        n13874) );
  AOI211_X1 U15369 ( .C1(P2_REG3_REG_23__SCAN_IN), .C2(P2_U3088), .A(n13875), 
        .B(n13874), .ZN(n13876) );
  OAI211_X1 U15370 ( .C1(n14452), .C2(n13974), .A(n13877), .B(n13876), .ZN(
        P2_U3188) );
  XNOR2_X1 U15371 ( .A(n13879), .B(n13878), .ZN(n13883) );
  OAI22_X1 U15372 ( .A1(n13995), .A2(n14273), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14072), .ZN(n13881) );
  OAI22_X1 U15373 ( .A1(n14265), .A2(n13997), .B1(n13998), .B2(n14222), .ZN(
        n13880) );
  AOI211_X1 U15374 ( .C1(n14461), .C2(n14001), .A(n13881), .B(n13880), .ZN(
        n13882) );
  OAI21_X1 U15375 ( .B1(n13883), .B2(n14003), .A(n13882), .ZN(P2_U3191) );
  NAND2_X1 U15376 ( .A1(n14114), .A2(n12208), .ZN(n13888) );
  XNOR2_X1 U15377 ( .A(n13888), .B(n7188), .ZN(n13889) );
  XNOR2_X1 U15378 ( .A(n14341), .B(n13889), .ZN(n13890) );
  XNOR2_X1 U15379 ( .A(n13891), .B(n13890), .ZN(n13897) );
  OAI22_X1 U15380 ( .A1(n14105), .A2(n13995), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13892), .ZN(n13895) );
  INV_X1 U15381 ( .A(n14100), .ZN(n13893) );
  OAI22_X1 U15382 ( .A1(n13893), .A2(n13998), .B1(n14135), .B2(n13997), .ZN(
        n13894) );
  AOI211_X1 U15383 ( .C1(n14341), .C2(n14001), .A(n13895), .B(n13894), .ZN(
        n13896) );
  OAI21_X1 U15384 ( .B1(n13897), .B2(n14003), .A(n13896), .ZN(P2_U3192) );
  XNOR2_X1 U15385 ( .A(n13899), .B(n13898), .ZN(n13904) );
  OAI22_X1 U15386 ( .A1(n13995), .A2(n14231), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13900), .ZN(n13902) );
  OAI22_X1 U15387 ( .A1(n14223), .A2(n13998), .B1(n13997), .B2(n14222), .ZN(
        n13901) );
  AOI211_X1 U15388 ( .C1(n14456), .C2(n14001), .A(n13902), .B(n13901), .ZN(
        n13903) );
  OAI21_X1 U15389 ( .B1(n13904), .B2(n14003), .A(n13903), .ZN(P2_U3195) );
  XNOR2_X1 U15390 ( .A(n13906), .B(n13905), .ZN(n13912) );
  INV_X1 U15391 ( .A(n14161), .ZN(n13908) );
  OAI22_X1 U15392 ( .A1(n13908), .A2(n13995), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13907), .ZN(n13910) );
  OAI22_X1 U15393 ( .A1(n14151), .A2(n13998), .B1(n14188), .B2(n13997), .ZN(
        n13909) );
  AOI211_X1 U15394 ( .C1(n14158), .C2(n14001), .A(n13910), .B(n13909), .ZN(
        n13911) );
  OAI21_X1 U15395 ( .B1(n13912), .B2(n14003), .A(n13911), .ZN(P2_U3197) );
  INV_X1 U15396 ( .A(n13913), .ZN(n13914) );
  AOI21_X1 U15397 ( .B1(n13916), .B2(n13915), .A(n13914), .ZN(n13922) );
  NOR2_X1 U15398 ( .A1(n13995), .A2(n13917), .ZN(n13920) );
  OAI22_X1 U15399 ( .A1(n13939), .A2(n13918), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14033), .ZN(n13919) );
  AOI211_X1 U15400 ( .C1(n14471), .C2(n14001), .A(n13920), .B(n13919), .ZN(
        n13921) );
  OAI21_X1 U15401 ( .B1(n13922), .B2(n14003), .A(n13921), .ZN(P2_U3198) );
  OAI21_X1 U15402 ( .B1(n13925), .B2(n13924), .A(n13923), .ZN(n13926) );
  NAND2_X1 U15403 ( .A1(n13926), .A2(n13966), .ZN(n13934) );
  INV_X1 U15404 ( .A(n13927), .ZN(n13930) );
  INV_X1 U15405 ( .A(n13928), .ZN(n13929) );
  AOI21_X1 U15406 ( .B1(n13957), .B2(n13930), .A(n13929), .ZN(n13933) );
  AOI22_X1 U15407 ( .A1(n13971), .A2(n13931), .B1(n14001), .B2(n15804), .ZN(
        n13932) );
  NAND3_X1 U15408 ( .A1(n13934), .A2(n13933), .A3(n13932), .ZN(P2_U3199) );
  OAI21_X1 U15409 ( .B1(n13937), .B2(n13936), .A(n13935), .ZN(n13938) );
  NAND2_X1 U15410 ( .A1(n13938), .A2(n13966), .ZN(n13943) );
  INV_X1 U15411 ( .A(n14317), .ZN(n13941) );
  AND2_X1 U15412 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n15403) );
  AOI22_X1 U15413 ( .A1(n14008), .A2(n14262), .B1(n14242), .B2(n14010), .ZN(
        n14311) );
  NOR2_X1 U15414 ( .A1(n13939), .A2(n14311), .ZN(n13940) );
  AOI211_X1 U15415 ( .C1(n13971), .C2(n13941), .A(n15403), .B(n13940), .ZN(
        n13942) );
  OAI211_X1 U15416 ( .C1(n14468), .C2(n13974), .A(n13943), .B(n13942), .ZN(
        P2_U3200) );
  AOI21_X1 U15417 ( .B1(n13945), .B2(n13944), .A(n14003), .ZN(n13947) );
  NAND2_X1 U15418 ( .A1(n13947), .A2(n13946), .ZN(n13951) );
  NOR2_X1 U15419 ( .A1(n13995), .A2(n14178), .ZN(n13949) );
  OAI22_X1 U15420 ( .A1(n14134), .A2(n13998), .B1(n14171), .B2(n13997), .ZN(
        n13948) );
  AOI211_X1 U15421 ( .C1(P2_REG3_REG_24__SCAN_IN), .C2(P2_U3088), .A(n13949), 
        .B(n13948), .ZN(n13950) );
  OAI211_X1 U15422 ( .C1(n14372), .C2(n13974), .A(n13951), .B(n13950), .ZN(
        P2_U3201) );
  OAI21_X1 U15423 ( .B1(n13954), .B2(n13953), .A(n13952), .ZN(n13955) );
  NAND2_X1 U15424 ( .A1(n13955), .A2(n13966), .ZN(n13962) );
  AOI22_X1 U15425 ( .A1(n13957), .A2(n13956), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13961) );
  AOI22_X1 U15426 ( .A1(n13971), .A2(n13959), .B1(n14001), .B2(n13958), .ZN(
        n13960) );
  NAND3_X1 U15427 ( .A1(n13962), .A2(n13961), .A3(n13960), .ZN(P2_U3202) );
  OAI21_X1 U15428 ( .B1(n13965), .B2(n13964), .A(n13963), .ZN(n13967) );
  NAND2_X1 U15429 ( .A1(n13967), .A2(n13966), .ZN(n13973) );
  NOR2_X1 U15430 ( .A1(n13968), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13970) );
  OAI22_X1 U15431 ( .A1(n14286), .A2(n13997), .B1(n13998), .B2(n13979), .ZN(
        n13969) );
  AOI211_X1 U15432 ( .C1(n13971), .C2(n14248), .A(n13970), .B(n13969), .ZN(
        n13972) );
  OAI211_X1 U15433 ( .C1(n7838), .C2(n13974), .A(n13973), .B(n13972), .ZN(
        P2_U3205) );
  XNOR2_X1 U15434 ( .A(n13976), .B(n13975), .ZN(n13983) );
  INV_X1 U15435 ( .A(n14210), .ZN(n13978) );
  OAI22_X1 U15436 ( .A1(n13995), .A2(n13978), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13977), .ZN(n13981) );
  OAI22_X1 U15437 ( .A1(n14171), .A2(n13998), .B1(n13997), .B2(n13979), .ZN(
        n13980) );
  AOI211_X1 U15438 ( .C1(n14386), .C2(n14001), .A(n13981), .B(n13980), .ZN(
        n13982) );
  OAI21_X1 U15439 ( .B1(n13983), .B2(n14003), .A(n13982), .ZN(P2_U3207) );
  XNOR2_X1 U15440 ( .A(n13984), .B(n13985), .ZN(n13989) );
  NAND2_X1 U15441 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14054)
         );
  OAI21_X1 U15442 ( .B1(n13995), .B2(n14297), .A(n14054), .ZN(n13987) );
  OAI22_X1 U15443 ( .A1(n14284), .A2(n13997), .B1(n13998), .B2(n14286), .ZN(
        n13986) );
  AOI211_X1 U15444 ( .C1(n14408), .C2(n14001), .A(n13987), .B(n13986), .ZN(
        n13988) );
  OAI21_X1 U15445 ( .B1(n13989), .B2(n14003), .A(n13988), .ZN(P2_U3210) );
  INV_X1 U15446 ( .A(n13990), .ZN(n13991) );
  AOI21_X1 U15447 ( .B1(n13993), .B2(n13992), .A(n13991), .ZN(n14004) );
  INV_X1 U15448 ( .A(n14141), .ZN(n13996) );
  OAI22_X1 U15449 ( .A1(n13996), .A2(n13995), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13994), .ZN(n14000) );
  OAI22_X1 U15450 ( .A1(n14135), .A2(n13998), .B1(n14134), .B2(n13997), .ZN(
        n13999) );
  AOI211_X1 U15451 ( .C1(n14363), .C2(n14001), .A(n14000), .B(n13999), .ZN(
        n14002) );
  OAI21_X1 U15452 ( .B1(n14004), .B2(n14003), .A(n14002), .ZN(P2_U3212) );
  MUX2_X1 U15453 ( .A(n14085), .B(P2_DATAO_REG_31__SCAN_IN), .S(n14025), .Z(
        P2_U3562) );
  MUX2_X1 U15454 ( .A(n14005), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14025), .Z(
        P2_U3561) );
  MUX2_X1 U15455 ( .A(n14100), .B(P2_DATAO_REG_29__SCAN_IN), .S(n14025), .Z(
        P2_U3560) );
  MUX2_X1 U15456 ( .A(n14114), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14025), .Z(
        P2_U3559) );
  MUX2_X1 U15457 ( .A(n14101), .B(P2_DATAO_REG_27__SCAN_IN), .S(n14025), .Z(
        P2_U3558) );
  MUX2_X1 U15458 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n14113), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15459 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n14169), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15460 ( .A(n14006), .B(P2_DATAO_REG_24__SCAN_IN), .S(n14025), .Z(
        P2_U3555) );
  MUX2_X1 U15461 ( .A(n14204), .B(P2_DATAO_REG_23__SCAN_IN), .S(n14025), .Z(
        P2_U3554) );
  MUX2_X1 U15462 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n14007), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U15463 ( .A(n14244), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14025), .Z(
        P2_U3552) );
  MUX2_X1 U15464 ( .A(n14263), .B(P2_DATAO_REG_20__SCAN_IN), .S(n14025), .Z(
        P2_U3551) );
  MUX2_X1 U15465 ( .A(n14243), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14025), .Z(
        P2_U3550) );
  MUX2_X1 U15466 ( .A(n14008), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14025), .Z(
        P2_U3549) );
  MUX2_X1 U15467 ( .A(n14009), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14025), .Z(
        P2_U3548) );
  MUX2_X1 U15468 ( .A(n14010), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14025), .Z(
        P2_U3547) );
  MUX2_X1 U15469 ( .A(n14011), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14025), .Z(
        P2_U3546) );
  MUX2_X1 U15470 ( .A(n14012), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14025), .Z(
        P2_U3545) );
  MUX2_X1 U15471 ( .A(n14013), .B(P2_DATAO_REG_13__SCAN_IN), .S(n14025), .Z(
        P2_U3544) );
  MUX2_X1 U15472 ( .A(n14014), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14025), .Z(
        P2_U3543) );
  MUX2_X1 U15473 ( .A(n14015), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14025), .Z(
        P2_U3542) );
  MUX2_X1 U15474 ( .A(n14016), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14025), .Z(
        P2_U3541) );
  MUX2_X1 U15475 ( .A(n14017), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14025), .Z(
        P2_U3540) );
  MUX2_X1 U15476 ( .A(n14018), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14025), .Z(
        P2_U3539) );
  MUX2_X1 U15477 ( .A(n14019), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14025), .Z(
        P2_U3538) );
  MUX2_X1 U15478 ( .A(n14020), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14025), .Z(
        P2_U3537) );
  MUX2_X1 U15479 ( .A(n14021), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14025), .Z(
        P2_U3536) );
  MUX2_X1 U15480 ( .A(n14022), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14025), .Z(
        P2_U3535) );
  MUX2_X1 U15481 ( .A(n14023), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14025), .Z(
        P2_U3534) );
  MUX2_X1 U15482 ( .A(n14024), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14025), .Z(
        P2_U3533) );
  MUX2_X1 U15483 ( .A(n12772), .B(P2_DATAO_REG_0__SCAN_IN), .S(n14025), .Z(
        P2_U3531) );
  NOR2_X1 U15484 ( .A1(n14028), .A2(n14040), .ZN(n14029) );
  XNOR2_X1 U15485 ( .A(n14040), .B(n14028), .ZN(n15390) );
  NOR2_X1 U15486 ( .A1(n15389), .A2(n15390), .ZN(n15388) );
  XNOR2_X1 U15487 ( .A(n14056), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14030) );
  NAND2_X1 U15488 ( .A1(n14031), .A2(n14030), .ZN(n14032) );
  NAND3_X1 U15489 ( .A1(n14032), .A2(n15419), .A3(n14057), .ZN(n14049) );
  NOR2_X1 U15490 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14033), .ZN(n14035) );
  INV_X1 U15491 ( .A(n14056), .ZN(n14044) );
  NOR2_X1 U15492 ( .A1(n14074), .A2(n14044), .ZN(n14034) );
  AOI211_X1 U15493 ( .C1(P2_ADDR_REG_16__SCAN_IN), .C2(n15341), .A(n14035), 
        .B(n14034), .ZN(n14048) );
  INV_X1 U15494 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n14036) );
  AOI22_X1 U15495 ( .A1(n14039), .A2(n14038), .B1(n14037), .B2(n14036), .ZN(
        n14041) );
  NAND2_X1 U15496 ( .A1(n15393), .A2(n14041), .ZN(n14042) );
  XNOR2_X1 U15497 ( .A(n14041), .B(n14040), .ZN(n15395) );
  NAND2_X1 U15498 ( .A1(n14042), .A2(n15394), .ZN(n14046) );
  NAND2_X1 U15499 ( .A1(n14056), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n14051) );
  INV_X1 U15500 ( .A(n14051), .ZN(n14043) );
  AOI21_X1 U15501 ( .B1(n12189), .B2(n14044), .A(n14043), .ZN(n14045) );
  NAND2_X1 U15502 ( .A1(n14045), .A2(n14046), .ZN(n14050) );
  OAI211_X1 U15503 ( .C1(n14046), .C2(n14045), .A(n15423), .B(n14050), .ZN(
        n14047) );
  NAND3_X1 U15504 ( .A1(n14049), .A2(n14048), .A3(n14047), .ZN(P2_U3230) );
  INV_X1 U15505 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n14052) );
  MUX2_X1 U15506 ( .A(n14052), .B(P2_REG2_REG_17__SCAN_IN), .S(n15404), .Z(
        n15408) );
  NOR2_X1 U15507 ( .A1(n15407), .A2(n15408), .ZN(n15405) );
  AOI21_X1 U15508 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n15404), .A(n15405), 
        .ZN(n14069) );
  XOR2_X1 U15509 ( .A(n14060), .B(n14069), .Z(n14053) );
  NOR2_X1 U15510 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n14053), .ZN(n14067) );
  AOI21_X1 U15511 ( .B1(n14053), .B2(P2_REG2_REG_18__SCAN_IN), .A(n14067), 
        .ZN(n14066) );
  OAI21_X1 U15512 ( .B1(n14074), .B2(n14068), .A(n14054), .ZN(n14055) );
  AOI21_X1 U15513 ( .B1(n15341), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n14055), 
        .ZN(n14065) );
  NAND2_X1 U15514 ( .A1(n14056), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n14058) );
  NAND2_X1 U15515 ( .A1(n14058), .A2(n14057), .ZN(n15399) );
  INV_X1 U15516 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14415) );
  XNOR2_X1 U15517 ( .A(n15404), .B(n14415), .ZN(n15400) );
  NAND2_X1 U15518 ( .A1(n15399), .A2(n15400), .ZN(n15398) );
  NAND2_X1 U15519 ( .A1(n15404), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n14059) );
  NAND2_X1 U15520 ( .A1(n15398), .A2(n14059), .ZN(n14061) );
  NAND2_X1 U15521 ( .A1(n14061), .A2(n14060), .ZN(n14076) );
  NAND2_X1 U15522 ( .A1(n14063), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n14077) );
  OAI211_X1 U15523 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n14063), .A(n15419), 
        .B(n14077), .ZN(n14064) );
  OAI211_X1 U15524 ( .C1(n14066), .C2(n15406), .A(n14065), .B(n14064), .ZN(
        P2_U3232) );
  MUX2_X1 U15525 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n14274), .S(n14078), .Z(
        n14070) );
  XNOR2_X1 U15526 ( .A(n14071), .B(n14070), .ZN(n14083) );
  OAI22_X1 U15527 ( .A1(n14074), .A2(n14073), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14072), .ZN(n14075) );
  AOI21_X1 U15528 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(n15341), .A(n14075), 
        .ZN(n14082) );
  NAND2_X1 U15529 ( .A1(n14077), .A2(n14076), .ZN(n14080) );
  XNOR2_X1 U15530 ( .A(n14078), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n14079) );
  XNOR2_X1 U15531 ( .A(n14080), .B(n14079), .ZN(n14081) );
  XNOR2_X1 U15532 ( .A(n14089), .B(n14427), .ZN(n14084) );
  NAND2_X1 U15533 ( .A1(n14084), .A2(n11286), .ZN(n14329) );
  NAND2_X1 U15534 ( .A1(n14086), .A2(n14085), .ZN(n14331) );
  NOR2_X1 U15535 ( .A1(n15817), .A2(n14331), .ZN(n14092) );
  NOR2_X1 U15536 ( .A1(n14427), .A2(n14301), .ZN(n14087) );
  AOI211_X1 U15537 ( .C1(n15829), .C2(P2_REG2_REG_31__SCAN_IN), .A(n14092), 
        .B(n14087), .ZN(n14088) );
  OAI21_X1 U15538 ( .B1(n14329), .B2(n14234), .A(n14088), .ZN(P2_U3234) );
  AOI21_X1 U15539 ( .B1(n7311), .B2(n14334), .A(n14295), .ZN(n14090) );
  NAND2_X1 U15540 ( .A1(n14090), .A2(n14089), .ZN(n14332) );
  NOR2_X1 U15541 ( .A1(n7842), .A2(n14301), .ZN(n14091) );
  AOI211_X1 U15542 ( .C1(n15829), .C2(P2_REG2_REG_30__SCAN_IN), .A(n14092), 
        .B(n14091), .ZN(n14093) );
  OAI21_X1 U15543 ( .B1(n14332), .B2(n14234), .A(n14093), .ZN(P2_U3235) );
  XNOR2_X1 U15544 ( .A(n14095), .B(n14094), .ZN(n14342) );
  INV_X1 U15545 ( .A(n14342), .ZN(n14111) );
  NAND2_X1 U15546 ( .A1(n14342), .A2(n15812), .ZN(n14103) );
  NAND2_X1 U15547 ( .A1(n14117), .A2(n14096), .ZN(n14098) );
  AOI22_X1 U15548 ( .A1(n14101), .A2(n14242), .B1(n14262), .B2(n14100), .ZN(
        n14102) );
  INV_X1 U15549 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n14104) );
  OAI22_X1 U15550 ( .A1(n14105), .A2(n14318), .B1(n14104), .B2(n14275), .ZN(
        n14108) );
  AOI21_X1 U15551 ( .B1(n14119), .B2(n14341), .A(n14295), .ZN(n14106) );
  NAND2_X1 U15552 ( .A1(n14106), .A2(n7267), .ZN(n14343) );
  NOR2_X1 U15553 ( .A1(n14343), .A2(n14234), .ZN(n14107) );
  AOI211_X1 U15554 ( .C1(n15818), .C2(n14341), .A(n14108), .B(n14107), .ZN(
        n14109) );
  OAI211_X1 U15555 ( .C1(n14129), .C2(n14111), .A(n14110), .B(n14109), .ZN(
        P2_U3237) );
  XNOR2_X1 U15556 ( .A(n14112), .B(n14116), .ZN(n14347) );
  AOI22_X1 U15557 ( .A1(n14114), .A2(n14262), .B1(n14113), .B2(n14242), .ZN(
        n14118) );
  NAND2_X1 U15558 ( .A1(n14353), .A2(n14275), .ZN(n14128) );
  INV_X1 U15559 ( .A(n14140), .ZN(n14121) );
  INV_X1 U15560 ( .A(n14119), .ZN(n14120) );
  AOI211_X1 U15561 ( .C1(n14122), .C2(n14121), .A(n14208), .B(n14120), .ZN(
        n14349) );
  INV_X1 U15562 ( .A(n14123), .ZN(n14124) );
  AOI22_X1 U15563 ( .A1(n14124), .A2(n15816), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n15829), .ZN(n14125) );
  OAI21_X1 U15564 ( .B1(n14437), .B2(n14301), .A(n14125), .ZN(n14126) );
  AOI21_X1 U15565 ( .B1(n14349), .B2(n15823), .A(n14126), .ZN(n14127) );
  OAI211_X1 U15566 ( .C1(n14347), .C2(n14129), .A(n14128), .B(n14127), .ZN(
        P2_U3238) );
  XNOR2_X1 U15567 ( .A(n14130), .B(n14133), .ZN(n14361) );
  OAI21_X1 U15568 ( .B1(n14133), .B2(n14132), .A(n14131), .ZN(n14137) );
  OAI22_X1 U15569 ( .A1(n14135), .A2(n14285), .B1(n14134), .B2(n14283), .ZN(
        n14136) );
  INV_X1 U15570 ( .A(n14360), .ZN(n14145) );
  NAND2_X1 U15571 ( .A1(n14159), .A2(n14363), .ZN(n14138) );
  NAND2_X1 U15572 ( .A1(n14138), .A2(n11286), .ZN(n14139) );
  OR2_X1 U15573 ( .A1(n14140), .A2(n14139), .ZN(n14359) );
  NOR2_X1 U15574 ( .A1(n14359), .A2(n14234), .ZN(n14144) );
  AOI22_X1 U15575 ( .A1(n14141), .A2(n15816), .B1(n15829), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n14142) );
  OAI21_X1 U15576 ( .B1(n14441), .B2(n14301), .A(n14142), .ZN(n14143) );
  AOI211_X1 U15577 ( .C1(n14145), .C2(n14275), .A(n14144), .B(n14143), .ZN(
        n14146) );
  OAI21_X1 U15578 ( .B1(n14254), .B2(n14361), .A(n14146), .ZN(P2_U3239) );
  NAND3_X1 U15579 ( .A1(n14168), .A2(n14148), .A3(n14147), .ZN(n14149) );
  NAND2_X1 U15580 ( .A1(n14150), .A2(n14149), .ZN(n14153) );
  OAI22_X1 U15581 ( .A1(n14151), .A2(n14285), .B1(n14188), .B2(n14283), .ZN(
        n14152) );
  AOI21_X1 U15582 ( .B1(n14153), .B2(n14309), .A(n14152), .ZN(n14367) );
  NAND2_X1 U15583 ( .A1(n14155), .A2(n14154), .ZN(n14156) );
  NAND2_X1 U15584 ( .A1(n14157), .A2(n14156), .ZN(n14366) );
  AOI21_X1 U15585 ( .B1(n14181), .B2(n14158), .A(n14295), .ZN(n14160) );
  AND2_X1 U15586 ( .A1(n14160), .A2(n14159), .ZN(n14365) );
  NAND2_X1 U15587 ( .A1(n14365), .A2(n15823), .ZN(n14163) );
  AOI22_X1 U15588 ( .A1(n14161), .A2(n15816), .B1(n15829), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n14162) );
  OAI211_X1 U15589 ( .C1(n14445), .C2(n14301), .A(n14163), .B(n14162), .ZN(
        n14164) );
  AOI21_X1 U15590 ( .B1(n14366), .B2(n14315), .A(n14164), .ZN(n14165) );
  OAI21_X1 U15591 ( .B1(n14367), .B2(n15817), .A(n14165), .ZN(P2_U3240) );
  NAND2_X1 U15592 ( .A1(n14166), .A2(n14174), .ZN(n14167) );
  NAND2_X1 U15593 ( .A1(n14168), .A2(n14167), .ZN(n14173) );
  NAND2_X1 U15594 ( .A1(n14169), .A2(n14262), .ZN(n14170) );
  OAI21_X1 U15595 ( .B1(n14171), .B2(n14283), .A(n14170), .ZN(n14172) );
  AOI21_X1 U15596 ( .B1(n14173), .B2(n14309), .A(n14172), .ZN(n14375) );
  OR2_X1 U15597 ( .A1(n14175), .A2(n14174), .ZN(n14176) );
  AND2_X1 U15598 ( .A1(n14177), .A2(n14176), .ZN(n14374) );
  INV_X1 U15599 ( .A(n14178), .ZN(n14179) );
  AOI22_X1 U15600 ( .A1(n15829), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n14179), 
        .B2(n15816), .ZN(n14180) );
  OAI21_X1 U15601 ( .B1(n14372), .B2(n14301), .A(n14180), .ZN(n14183) );
  OAI211_X1 U15602 ( .C1(n14196), .C2(n14372), .A(n11286), .B(n14181), .ZN(
        n14371) );
  NOR2_X1 U15603 ( .A1(n14371), .A2(n14234), .ZN(n14182) );
  AOI211_X1 U15604 ( .C1(n14374), .C2(n14315), .A(n14183), .B(n14182), .ZN(
        n14184) );
  OAI21_X1 U15605 ( .B1(n15817), .B2(n14375), .A(n14184), .ZN(P2_U3241) );
  XNOR2_X1 U15606 ( .A(n14185), .B(n14186), .ZN(n14380) );
  NAND2_X1 U15607 ( .A1(n14380), .A2(n15812), .ZN(n14192) );
  XNOR2_X1 U15608 ( .A(n14187), .B(n14186), .ZN(n14190) );
  OAI22_X1 U15609 ( .A1(n14188), .A2(n14285), .B1(n14223), .B2(n14283), .ZN(
        n14189) );
  AOI21_X1 U15610 ( .B1(n14190), .B2(n14309), .A(n14189), .ZN(n14191) );
  NAND2_X1 U15611 ( .A1(n14193), .A2(n14206), .ZN(n14194) );
  NAND2_X1 U15612 ( .A1(n14194), .A2(n11286), .ZN(n14195) );
  NOR2_X1 U15613 ( .A1(n14196), .A2(n14195), .ZN(n14379) );
  NAND2_X1 U15614 ( .A1(n14379), .A2(n15823), .ZN(n14200) );
  INV_X1 U15615 ( .A(n14197), .ZN(n14198) );
  AOI22_X1 U15616 ( .A1(n15817), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n14198), 
        .B2(n15816), .ZN(n14199) );
  OAI211_X1 U15617 ( .C1(n14452), .C2(n14301), .A(n14200), .B(n14199), .ZN(
        n14201) );
  AOI21_X1 U15618 ( .B1(n15824), .B2(n14380), .A(n14201), .ZN(n14202) );
  OAI21_X1 U15619 ( .B1(n14382), .B2(n15817), .A(n14202), .ZN(P2_U3242) );
  XOR2_X1 U15620 ( .A(n14203), .B(n14213), .Z(n14205) );
  AOI222_X1 U15621 ( .A1(n14309), .A2(n14205), .B1(n14244), .B2(n14242), .C1(
        n14204), .C2(n14262), .ZN(n14388) );
  INV_X1 U15622 ( .A(n14228), .ZN(n14209) );
  INV_X1 U15623 ( .A(n14206), .ZN(n14207) );
  AOI211_X1 U15624 ( .C1(n14386), .C2(n14209), .A(n14208), .B(n14207), .ZN(
        n14385) );
  AOI22_X1 U15625 ( .A1(n15817), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n14210), 
        .B2(n15816), .ZN(n14211) );
  OAI21_X1 U15626 ( .B1(n14212), .B2(n14301), .A(n14211), .ZN(n14216) );
  XNOR2_X1 U15627 ( .A(n14214), .B(n14213), .ZN(n14389) );
  NOR2_X1 U15628 ( .A1(n14389), .A2(n14254), .ZN(n14215) );
  AOI211_X1 U15629 ( .C1(n14385), .C2(n15823), .A(n14216), .B(n14215), .ZN(
        n14217) );
  OAI21_X1 U15630 ( .B1(n14388), .B2(n15817), .A(n14217), .ZN(P2_U3243) );
  INV_X1 U15631 ( .A(n14220), .ZN(n14218) );
  XNOR2_X1 U15632 ( .A(n14219), .B(n14218), .ZN(n14392) );
  AOI21_X1 U15633 ( .B1(n14221), .B2(n14220), .A(n14289), .ZN(n14226) );
  OAI22_X1 U15634 ( .A1(n14223), .A2(n14285), .B1(n14222), .B2(n14283), .ZN(
        n14224) );
  AOI21_X1 U15635 ( .B1(n14226), .B2(n14225), .A(n14224), .ZN(n14391) );
  INV_X1 U15636 ( .A(n14391), .ZN(n14236) );
  NAND2_X1 U15637 ( .A1(n14456), .A2(n14247), .ZN(n14227) );
  NAND2_X1 U15638 ( .A1(n14227), .A2(n11286), .ZN(n14229) );
  OR2_X1 U15639 ( .A1(n14229), .A2(n14228), .ZN(n14390) );
  NAND2_X1 U15640 ( .A1(n15829), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n14230) );
  OAI21_X1 U15641 ( .B1(n14318), .B2(n14231), .A(n14230), .ZN(n14232) );
  AOI21_X1 U15642 ( .B1(n14456), .B2(n15818), .A(n14232), .ZN(n14233) );
  OAI21_X1 U15643 ( .B1(n14390), .B2(n14234), .A(n14233), .ZN(n14235) );
  AOI21_X1 U15644 ( .B1(n14236), .B2(n14275), .A(n14235), .ZN(n14237) );
  OAI21_X1 U15645 ( .B1(n14254), .B2(n14392), .A(n14237), .ZN(P2_U3244) );
  XNOR2_X1 U15646 ( .A(n14238), .B(n14240), .ZN(n14399) );
  OAI21_X1 U15647 ( .B1(n14241), .B2(n14240), .A(n14239), .ZN(n14245) );
  AOI222_X1 U15648 ( .A1(n14309), .A2(n14245), .B1(n14244), .B2(n14262), .C1(
        n14243), .C2(n14242), .ZN(n14398) );
  INV_X1 U15649 ( .A(n14398), .ZN(n14252) );
  AOI21_X1 U15650 ( .B1(n14396), .B2(n14271), .A(n14295), .ZN(n14246) );
  AND2_X1 U15651 ( .A1(n14247), .A2(n14246), .ZN(n14395) );
  NAND2_X1 U15652 ( .A1(n14395), .A2(n15823), .ZN(n14250) );
  AOI22_X1 U15653 ( .A1(n15829), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14248), 
        .B2(n15816), .ZN(n14249) );
  OAI211_X1 U15654 ( .C1(n7838), .C2(n14301), .A(n14250), .B(n14249), .ZN(
        n14251) );
  AOI21_X1 U15655 ( .B1(n14252), .B2(n14275), .A(n14251), .ZN(n14253) );
  OAI21_X1 U15656 ( .B1(n14254), .B2(n14399), .A(n14253), .ZN(P2_U3245) );
  OR2_X1 U15657 ( .A1(n14255), .A2(n14258), .ZN(n14257) );
  NAND2_X1 U15658 ( .A1(n14257), .A2(n14256), .ZN(n14401) );
  NAND2_X1 U15659 ( .A1(n14401), .A2(n15812), .ZN(n14270) );
  NAND2_X1 U15660 ( .A1(n14259), .A2(n14258), .ZN(n14260) );
  NAND2_X1 U15661 ( .A1(n14261), .A2(n14260), .ZN(n14268) );
  NAND2_X1 U15662 ( .A1(n14263), .A2(n14262), .ZN(n14264) );
  OAI21_X1 U15663 ( .B1(n14265), .B2(n14283), .A(n14264), .ZN(n14266) );
  AOI21_X1 U15664 ( .B1(n14268), .B2(n14267), .A(n14266), .ZN(n14269) );
  AOI21_X1 U15665 ( .B1(n14293), .B2(n14461), .A(n14295), .ZN(n14272) );
  AND2_X1 U15666 ( .A1(n14272), .A2(n14271), .ZN(n14400) );
  OAI22_X1 U15667 ( .A1(n14275), .A2(n14274), .B1(n14273), .B2(n14318), .ZN(
        n14278) );
  INV_X1 U15668 ( .A(n14461), .ZN(n14276) );
  NOR2_X1 U15669 ( .A1(n14276), .A2(n14301), .ZN(n14277) );
  AOI211_X1 U15670 ( .C1(n14400), .C2(n15823), .A(n14278), .B(n14277), .ZN(
        n14280) );
  NAND2_X1 U15671 ( .A1(n14401), .A2(n15824), .ZN(n14279) );
  OAI211_X1 U15672 ( .C1(n14403), .C2(n15817), .A(n14280), .B(n14279), .ZN(
        P2_U3246) );
  OAI21_X1 U15673 ( .B1(n14282), .B2(n14288), .A(n14281), .ZN(n14406) );
  OAI22_X1 U15674 ( .A1(n14286), .A2(n14285), .B1(n14284), .B2(n14283), .ZN(
        n14292) );
  XOR2_X1 U15675 ( .A(n14287), .B(n14288), .Z(n14290) );
  NOR2_X1 U15676 ( .A1(n14290), .A2(n14289), .ZN(n14291) );
  AOI211_X1 U15677 ( .C1(n15812), .C2(n14406), .A(n14292), .B(n14291), .ZN(
        n14410) );
  INV_X1 U15678 ( .A(n14324), .ZN(n14296) );
  INV_X1 U15679 ( .A(n14293), .ZN(n14294) );
  AOI211_X1 U15680 ( .C1(n14408), .C2(n14296), .A(n14295), .B(n14294), .ZN(
        n14407) );
  NAND2_X1 U15681 ( .A1(n14407), .A2(n15823), .ZN(n14300) );
  INV_X1 U15682 ( .A(n14297), .ZN(n14298) );
  AOI22_X1 U15683 ( .A1(n15829), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14298), 
        .B2(n15816), .ZN(n14299) );
  OAI211_X1 U15684 ( .C1(n14302), .C2(n14301), .A(n14300), .B(n14299), .ZN(
        n14303) );
  AOI21_X1 U15685 ( .B1(n15824), .B2(n14406), .A(n14303), .ZN(n14304) );
  OAI21_X1 U15686 ( .B1(n14410), .B2(n15817), .A(n14304), .ZN(P2_U3247) );
  INV_X1 U15687 ( .A(n14313), .ZN(n14306) );
  NAND3_X1 U15688 ( .A1(n14307), .A2(n14306), .A3(n14305), .ZN(n14308) );
  NAND3_X1 U15689 ( .A1(n14310), .A2(n14309), .A3(n14308), .ZN(n14312) );
  NAND2_X1 U15690 ( .A1(n14312), .A2(n14311), .ZN(n14412) );
  NAND2_X1 U15691 ( .A1(n14412), .A2(n14275), .ZN(n14328) );
  XNOR2_X1 U15692 ( .A(n14314), .B(n14313), .ZN(n14414) );
  NAND2_X1 U15693 ( .A1(n14414), .A2(n14315), .ZN(n14327) );
  NAND2_X1 U15694 ( .A1(n15829), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n14316) );
  OAI21_X1 U15695 ( .B1(n14318), .B2(n14317), .A(n14316), .ZN(n14319) );
  AOI21_X1 U15696 ( .B1(n14320), .B2(n15818), .A(n14319), .ZN(n14326) );
  NAND2_X1 U15697 ( .A1(n14321), .A2(n14320), .ZN(n14322) );
  NAND2_X1 U15698 ( .A1(n14322), .A2(n11286), .ZN(n14323) );
  NOR2_X1 U15699 ( .A1(n14324), .A2(n14323), .ZN(n14413) );
  NAND2_X1 U15700 ( .A1(n14413), .A2(n15823), .ZN(n14325) );
  NAND4_X1 U15701 ( .A1(n14328), .A2(n14327), .A3(n14326), .A4(n14325), .ZN(
        P2_U3248) );
  NAND2_X1 U15702 ( .A1(n14332), .A2(n14331), .ZN(n14428) );
  MUX2_X1 U15703 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14428), .S(n15970), .Z(
        n14333) );
  AOI21_X1 U15704 ( .B1(n14422), .B2(n14334), .A(n14333), .ZN(n14335) );
  INV_X1 U15705 ( .A(n14335), .ZN(P2_U3529) );
  AOI21_X1 U15706 ( .B1(n15845), .B2(n14337), .A(n14336), .ZN(n14338) );
  OAI211_X1 U15707 ( .C1(n15847), .C2(n14340), .A(n14339), .B(n14338), .ZN(
        n14432) );
  MUX2_X1 U15708 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14432), .S(n15970), .Z(
        P2_U3528) );
  INV_X1 U15709 ( .A(n14341), .ZN(n14345) );
  NAND2_X1 U15710 ( .A1(n14342), .A2(n15950), .ZN(n14344) );
  OAI211_X1 U15711 ( .C1(n14345), .C2(n15963), .A(n14344), .B(n14343), .ZN(
        n14346) );
  INV_X1 U15712 ( .A(n14347), .ZN(n14348) );
  INV_X1 U15713 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n14354) );
  NAND2_X1 U15714 ( .A1(n14355), .A2(n14354), .ZN(n14356) );
  OAI21_X1 U15715 ( .B1(n14437), .B2(n14417), .A(n14358), .ZN(P2_U3526) );
  INV_X1 U15716 ( .A(n14364), .ZN(P2_U3525) );
  INV_X1 U15717 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14369) );
  AOI21_X1 U15718 ( .B1(n14366), .B2(n15968), .A(n14365), .ZN(n14368) );
  AND2_X1 U15719 ( .A1(n14368), .A2(n14367), .ZN(n14442) );
  MUX2_X1 U15720 ( .A(n14369), .B(n14442), .S(n15970), .Z(n14370) );
  OAI21_X1 U15721 ( .B1(n14445), .B2(n14417), .A(n14370), .ZN(P2_U3524) );
  INV_X1 U15722 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n14377) );
  OAI21_X1 U15723 ( .B1(n14372), .B2(n15963), .A(n14371), .ZN(n14373) );
  AOI21_X1 U15724 ( .B1(n14374), .B2(n15968), .A(n14373), .ZN(n14376) );
  AND2_X1 U15725 ( .A1(n14376), .A2(n14375), .ZN(n14446) );
  MUX2_X1 U15726 ( .A(n14377), .B(n14446), .S(n15970), .Z(n14378) );
  INV_X1 U15727 ( .A(n14378), .ZN(P2_U3523) );
  INV_X1 U15728 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n14383) );
  AOI21_X1 U15729 ( .B1(n14380), .B2(n15950), .A(n14379), .ZN(n14381) );
  AND2_X1 U15730 ( .A1(n14382), .A2(n14381), .ZN(n14449) );
  MUX2_X1 U15731 ( .A(n14383), .B(n14449), .S(n15970), .Z(n14384) );
  OAI21_X1 U15732 ( .B1(n14452), .B2(n14417), .A(n14384), .ZN(P2_U3522) );
  AOI21_X1 U15733 ( .B1(n15845), .B2(n14386), .A(n14385), .ZN(n14387) );
  OAI211_X1 U15734 ( .C1(n15847), .C2(n14389), .A(n14388), .B(n14387), .ZN(
        n14453) );
  MUX2_X1 U15735 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14453), .S(n15970), .Z(
        P2_U3521) );
  OAI211_X1 U15736 ( .C1(n14392), .C2(n15847), .A(n14391), .B(n14390), .ZN(
        n14454) );
  MUX2_X1 U15737 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14454), .S(n15970), .Z(
        n14393) );
  AOI21_X1 U15738 ( .B1(n14422), .B2(n14456), .A(n14393), .ZN(n14394) );
  INV_X1 U15739 ( .A(n14394), .ZN(P2_U3520) );
  AOI21_X1 U15740 ( .B1(n15845), .B2(n14396), .A(n14395), .ZN(n14397) );
  OAI211_X1 U15741 ( .C1(n15847), .C2(n14399), .A(n14398), .B(n14397), .ZN(
        n14458) );
  MUX2_X1 U15742 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14458), .S(n15970), .Z(
        P2_U3519) );
  AOI21_X1 U15743 ( .B1(n14401), .B2(n15950), .A(n14400), .ZN(n14402) );
  NAND2_X1 U15744 ( .A1(n14403), .A2(n14402), .ZN(n14459) );
  MUX2_X1 U15745 ( .A(n14459), .B(P2_REG1_REG_19__SCAN_IN), .S(n14355), .Z(
        n14404) );
  AOI21_X1 U15746 ( .B1(n14422), .B2(n14461), .A(n14404), .ZN(n14405) );
  INV_X1 U15747 ( .A(n14405), .ZN(P2_U3518) );
  INV_X1 U15748 ( .A(n14406), .ZN(n14411) );
  AOI21_X1 U15749 ( .B1(n15845), .B2(n14408), .A(n14407), .ZN(n14409) );
  OAI211_X1 U15750 ( .C1(n14411), .C2(n15807), .A(n14410), .B(n14409), .ZN(
        n14463) );
  MUX2_X1 U15751 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14463), .S(n15970), .Z(
        P2_U3517) );
  AOI211_X1 U15752 ( .C1(n15968), .C2(n14414), .A(n14413), .B(n14412), .ZN(
        n14464) );
  MUX2_X1 U15753 ( .A(n14415), .B(n14464), .S(n15970), .Z(n14416) );
  OAI21_X1 U15754 ( .B1(n14468), .B2(n14417), .A(n14416), .ZN(P2_U3516) );
  OAI211_X1 U15755 ( .C1(n14420), .C2(n15847), .A(n14419), .B(n14418), .ZN(
        n14469) );
  MUX2_X1 U15756 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14469), .S(n15970), .Z(
        n14421) );
  AOI21_X1 U15757 ( .B1(n14422), .B2(n14471), .A(n14421), .ZN(n14423) );
  INV_X1 U15758 ( .A(n14423), .ZN(P2_U3515) );
  MUX2_X1 U15759 ( .A(n14424), .B(P2_REG0_REG_31__SCAN_IN), .S(n15971), .Z(
        n14425) );
  INV_X1 U15760 ( .A(n14425), .ZN(n14426) );
  OAI21_X1 U15761 ( .B1(n14427), .B2(n14467), .A(n14426), .ZN(P2_U3498) );
  INV_X1 U15762 ( .A(n14428), .ZN(n14429) );
  MUX2_X1 U15763 ( .A(n14430), .B(n14429), .S(n15974), .Z(n14431) );
  OAI21_X1 U15764 ( .B1(n7842), .B2(n14467), .A(n14431), .ZN(P2_U3497) );
  MUX2_X1 U15765 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n14432), .S(n15974), .Z(
        P2_U3496) );
  OAI21_X1 U15766 ( .B1(n14437), .B2(n14467), .A(n14436), .ZN(P2_U3494) );
  MUX2_X1 U15767 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14438), .S(n15974), .Z(
        n14439) );
  INV_X1 U15768 ( .A(n14439), .ZN(n14440) );
  OAI21_X1 U15769 ( .B1(n14441), .B2(n14467), .A(n14440), .ZN(P2_U3493) );
  MUX2_X1 U15770 ( .A(n14443), .B(n14442), .S(n15974), .Z(n14444) );
  OAI21_X1 U15771 ( .B1(n14445), .B2(n14467), .A(n14444), .ZN(P2_U3492) );
  MUX2_X1 U15772 ( .A(n14447), .B(n14446), .S(n15974), .Z(n14448) );
  INV_X1 U15773 ( .A(n14448), .ZN(P2_U3491) );
  MUX2_X1 U15774 ( .A(n14450), .B(n14449), .S(n15974), .Z(n14451) );
  OAI21_X1 U15775 ( .B1(n14452), .B2(n14467), .A(n14451), .ZN(P2_U3490) );
  MUX2_X1 U15776 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14453), .S(n15974), .Z(
        P2_U3489) );
  INV_X1 U15777 ( .A(n14467), .ZN(n14472) );
  MUX2_X1 U15778 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14454), .S(n15974), .Z(
        n14455) );
  AOI21_X1 U15779 ( .B1(n14472), .B2(n14456), .A(n14455), .ZN(n14457) );
  INV_X1 U15780 ( .A(n14457), .ZN(P2_U3488) );
  MUX2_X1 U15781 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14458), .S(n15974), .Z(
        P2_U3487) );
  MUX2_X1 U15782 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14459), .S(n15974), .Z(
        n14460) );
  AOI21_X1 U15783 ( .B1(n14472), .B2(n14461), .A(n14460), .ZN(n14462) );
  INV_X1 U15784 ( .A(n14462), .ZN(P2_U3486) );
  MUX2_X1 U15785 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14463), .S(n15974), .Z(
        P2_U3484) );
  MUX2_X1 U15786 ( .A(n14465), .B(n14464), .S(n15974), .Z(n14466) );
  OAI21_X1 U15787 ( .B1(n14468), .B2(n14467), .A(n14466), .ZN(P2_U3481) );
  MUX2_X1 U15788 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14469), .S(n15974), .Z(
        n14470) );
  AOI21_X1 U15789 ( .B1(n14472), .B2(n14471), .A(n14470), .ZN(n14473) );
  INV_X1 U15790 ( .A(n14473), .ZN(P2_U3478) );
  NAND2_X1 U15791 ( .A1(n15194), .A2(n14500), .ZN(n14478) );
  NAND4_X1 U15792 ( .A1(n14476), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .A4(n14475), .ZN(n14477) );
  OAI211_X1 U15793 ( .C1(n14503), .C2(n14479), .A(n14478), .B(n14477), .ZN(
        P2_U3296) );
  INV_X1 U15794 ( .A(n14480), .ZN(n15199) );
  OAI222_X1 U15795 ( .A1(n14506), .A2(n15199), .B1(P2_U3088), .B2(n14482), 
        .C1(n14481), .C2(n14503), .ZN(P2_U3298) );
  NAND2_X1 U15796 ( .A1(n14483), .A2(n14500), .ZN(n14485) );
  OAI211_X1 U15797 ( .C1(n14486), .C2(n14503), .A(n14485), .B(n14484), .ZN(
        P2_U3299) );
  OAI222_X1 U15798 ( .A1(n14509), .A2(n14489), .B1(n14506), .B2(n14488), .C1(
        P2_U3088), .C2(n14487), .ZN(P2_U3300) );
  INV_X1 U15799 ( .A(n14490), .ZN(n14493) );
  INV_X1 U15800 ( .A(n14491), .ZN(n15202) );
  OAI222_X1 U15801 ( .A1(P2_U3088), .A2(n14493), .B1(n14506), .B2(n15202), 
        .C1(n14492), .C2(n14503), .ZN(P2_U3301) );
  INV_X1 U15802 ( .A(n14494), .ZN(n15206) );
  OAI222_X1 U15803 ( .A1(n14509), .A2(n14496), .B1(n14506), .B2(n15206), .C1(
        P2_U3088), .C2(n14495), .ZN(P2_U3302) );
  INV_X1 U15804 ( .A(n14497), .ZN(n15208) );
  OAI222_X1 U15805 ( .A1(n14509), .A2(n14499), .B1(n14506), .B2(n15208), .C1(
        P2_U3088), .C2(n14498), .ZN(P2_U3303) );
  NAND2_X1 U15806 ( .A1(n15211), .A2(n14500), .ZN(n14502) );
  OAI211_X1 U15807 ( .C1(n14504), .C2(n14503), .A(n14502), .B(n14501), .ZN(
        P2_U3304) );
  OAI222_X1 U15808 ( .A1(n14509), .A2(n14508), .B1(P2_U3088), .B2(n14507), 
        .C1(n14506), .C2(n14505), .ZN(P2_U3305) );
  INV_X1 U15809 ( .A(n14510), .ZN(n14511) );
  MUX2_X1 U15810 ( .A(n14511), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI22_X1 U15811 ( .A1(n14861), .A2(n14582), .B1(n14841), .B2(n14613), .ZN(
        n14655) );
  NAND2_X1 U15812 ( .A1(n15087), .A2(n9735), .ZN(n14513) );
  NAND2_X1 U15813 ( .A1(n14877), .A2(n14659), .ZN(n14512) );
  NAND2_X1 U15814 ( .A1(n14513), .A2(n14512), .ZN(n14514) );
  XNOR2_X1 U15815 ( .A(n14514), .B(n14661), .ZN(n14654) );
  XOR2_X1 U15816 ( .A(n14655), .B(n14654), .Z(n14658) );
  INV_X1 U15817 ( .A(n14515), .ZN(n14517) );
  OAI22_X1 U15818 ( .A1(n14521), .A2(n14583), .B1(n14520), .B2(n14582), .ZN(
        n14519) );
  XNOR2_X1 U15819 ( .A(n14519), .B(n14584), .ZN(n14524) );
  OAI22_X1 U15820 ( .A1(n14521), .A2(n7189), .B1(n14520), .B2(n14613), .ZN(
        n14523) );
  XNOR2_X1 U15821 ( .A(n14524), .B(n14523), .ZN(n14632) );
  OR2_X1 U15822 ( .A1(n14524), .A2(n14523), .ZN(n14525) );
  NAND2_X1 U15823 ( .A1(n15989), .A2(n14614), .ZN(n14527) );
  NAND2_X1 U15824 ( .A1(n16000), .A2(n14659), .ZN(n14526) );
  NAND2_X1 U15825 ( .A1(n14527), .A2(n14526), .ZN(n14528) );
  XNOR2_X1 U15826 ( .A(n14528), .B(n14661), .ZN(n14530) );
  AOI22_X1 U15827 ( .A1(n15989), .A2(n14659), .B1(n14607), .B2(n16000), .ZN(
        n15977) );
  NAND2_X1 U15828 ( .A1(n15976), .A2(n15977), .ZN(n15975) );
  INV_X1 U15829 ( .A(n14529), .ZN(n14531) );
  NAND2_X1 U15830 ( .A1(n15975), .A2(n8261), .ZN(n15997) );
  OAI22_X1 U15831 ( .A1(n16003), .A2(n14582), .B1(n14532), .B2(n14613), .ZN(
        n14536) );
  NAND2_X1 U15832 ( .A1(n16013), .A2(n14614), .ZN(n14534) );
  NAND2_X1 U15833 ( .A1(n16028), .A2(n14659), .ZN(n14533) );
  NAND2_X1 U15834 ( .A1(n14534), .A2(n14533), .ZN(n14535) );
  XNOR2_X1 U15835 ( .A(n14535), .B(n14661), .ZN(n14537) );
  XOR2_X1 U15836 ( .A(n14536), .B(n14537), .Z(n15999) );
  NAND2_X1 U15837 ( .A1(n15997), .A2(n15999), .ZN(n14539) );
  OR2_X1 U15838 ( .A1(n14537), .A2(n14536), .ZN(n14538) );
  NAND2_X1 U15839 ( .A1(n14539), .A2(n14538), .ZN(n16025) );
  NAND2_X1 U15840 ( .A1(n16027), .A2(n14614), .ZN(n14541) );
  NAND2_X1 U15841 ( .A1(n16001), .A2(n14659), .ZN(n14540) );
  NAND2_X1 U15842 ( .A1(n14541), .A2(n14540), .ZN(n14542) );
  XNOR2_X1 U15843 ( .A(n14542), .B(n14661), .ZN(n14545) );
  AOI22_X1 U15844 ( .A1(n16027), .A2(n14615), .B1(n14607), .B2(n16001), .ZN(
        n14543) );
  XNOR2_X1 U15845 ( .A(n14545), .B(n14543), .ZN(n16026) );
  NAND2_X1 U15846 ( .A1(n16025), .A2(n16026), .ZN(n14547) );
  INV_X1 U15847 ( .A(n14543), .ZN(n14544) );
  NAND2_X1 U15848 ( .A1(n15153), .A2(n14614), .ZN(n14549) );
  NAND2_X1 U15849 ( .A1(n16030), .A2(n14659), .ZN(n14548) );
  NAND2_X1 U15850 ( .A1(n14549), .A2(n14548), .ZN(n14550) );
  XNOR2_X1 U15851 ( .A(n14550), .B(n14661), .ZN(n14553) );
  AOI22_X1 U15852 ( .A1(n15153), .A2(n14659), .B1(n14607), .B2(n16030), .ZN(
        n14551) );
  XNOR2_X1 U15853 ( .A(n14553), .B(n14551), .ZN(n14717) );
  INV_X1 U15854 ( .A(n14551), .ZN(n14552) );
  OR2_X1 U15855 ( .A1(n14553), .A2(n14552), .ZN(n14554) );
  NAND2_X1 U15856 ( .A1(n15145), .A2(n14614), .ZN(n14556) );
  NAND2_X1 U15857 ( .A1(n15008), .A2(n14659), .ZN(n14555) );
  NAND2_X1 U15858 ( .A1(n14556), .A2(n14555), .ZN(n14557) );
  XNOR2_X1 U15859 ( .A(n14557), .B(n14661), .ZN(n14558) );
  AOI22_X1 U15860 ( .A1(n15145), .A2(n14659), .B1(n14607), .B2(n15008), .ZN(
        n14559) );
  XNOR2_X1 U15861 ( .A(n14558), .B(n14559), .ZN(n14647) );
  INV_X1 U15862 ( .A(n14558), .ZN(n14560) );
  INV_X1 U15863 ( .A(n14697), .ZN(n14567) );
  AND2_X1 U15864 ( .A1(n14963), .A2(n14607), .ZN(n14561) );
  AOI21_X1 U15865 ( .B1(n14562), .B2(n14659), .A(n14561), .ZN(n14568) );
  NAND2_X1 U15866 ( .A1(n14562), .A2(n14614), .ZN(n14564) );
  NAND2_X1 U15867 ( .A1(n14963), .A2(n14615), .ZN(n14563) );
  NAND2_X1 U15868 ( .A1(n14564), .A2(n14563), .ZN(n14565) );
  XNOR2_X1 U15869 ( .A(n14565), .B(n14661), .ZN(n14570) );
  XOR2_X1 U15870 ( .A(n14568), .B(n14570), .Z(n14696) );
  INV_X1 U15871 ( .A(n14696), .ZN(n14566) );
  INV_X1 U15872 ( .A(n14568), .ZN(n14569) );
  NAND2_X1 U15873 ( .A1(n14570), .A2(n14569), .ZN(n14571) );
  OAI22_X1 U15874 ( .A1(n15129), .A2(n14583), .B1(n14573), .B2(n7189), .ZN(
        n14572) );
  XNOR2_X1 U15875 ( .A(n14572), .B(n14661), .ZN(n14575) );
  OAI22_X1 U15876 ( .A1(n15129), .A2(n7189), .B1(n14573), .B2(n14613), .ZN(
        n14576) );
  XNOR2_X1 U15877 ( .A(n14575), .B(n14576), .ZN(n14674) );
  INV_X1 U15878 ( .A(n14674), .ZN(n14574) );
  INV_X1 U15879 ( .A(n14575), .ZN(n14578) );
  INV_X1 U15880 ( .A(n14576), .ZN(n14577) );
  NAND2_X1 U15881 ( .A1(n14578), .A2(n14577), .ZN(n14579) );
  OR2_X1 U15882 ( .A1(n14954), .A2(n7189), .ZN(n14581) );
  NAND2_X1 U15883 ( .A1(n14962), .A2(n14607), .ZN(n14580) );
  NAND2_X1 U15884 ( .A1(n14581), .A2(n14580), .ZN(n14587) );
  OAI22_X1 U15885 ( .A1(n14954), .A2(n14583), .B1(n14927), .B2(n14582), .ZN(
        n14585) );
  XNOR2_X1 U15886 ( .A(n14585), .B(n14584), .ZN(n14586) );
  XOR2_X1 U15887 ( .A(n14587), .B(n14586), .Z(n14708) );
  NAND2_X1 U15888 ( .A1(n14707), .A2(n14708), .ZN(n14706) );
  INV_X1 U15889 ( .A(n14586), .ZN(n14589) );
  INV_X1 U15890 ( .A(n14587), .ZN(n14588) );
  NAND2_X1 U15891 ( .A1(n14589), .A2(n14588), .ZN(n14590) );
  NAND2_X1 U15892 ( .A1(n15117), .A2(n14614), .ZN(n14592) );
  NAND2_X1 U15893 ( .A1(n14738), .A2(n14659), .ZN(n14591) );
  NAND2_X1 U15894 ( .A1(n14592), .A2(n14591), .ZN(n14593) );
  XNOR2_X1 U15895 ( .A(n14593), .B(n14661), .ZN(n14594) );
  AOI22_X1 U15896 ( .A1(n15117), .A2(n14659), .B1(n14607), .B2(n14738), .ZN(
        n14595) );
  XNOR2_X1 U15897 ( .A(n14594), .B(n14595), .ZN(n14641) );
  INV_X1 U15898 ( .A(n14594), .ZN(n14596) );
  NAND2_X1 U15899 ( .A1(n14596), .A2(n14595), .ZN(n14597) );
  NAND2_X1 U15900 ( .A1(n15107), .A2(n14614), .ZN(n14599) );
  NAND2_X1 U15901 ( .A1(n14925), .A2(n14659), .ZN(n14598) );
  NAND2_X1 U15902 ( .A1(n14599), .A2(n14598), .ZN(n14600) );
  XNOR2_X1 U15903 ( .A(n14600), .B(n14661), .ZN(n14601) );
  AOI22_X1 U15904 ( .A1(n15107), .A2(n14659), .B1(n14607), .B2(n14925), .ZN(
        n14602) );
  XNOR2_X1 U15905 ( .A(n14601), .B(n14602), .ZN(n14688) );
  INV_X1 U15906 ( .A(n14601), .ZN(n14603) );
  NAND2_X1 U15907 ( .A1(n14895), .A2(n14614), .ZN(n14605) );
  NAND2_X1 U15908 ( .A1(n14876), .A2(n14659), .ZN(n14604) );
  NAND2_X1 U15909 ( .A1(n14605), .A2(n14604), .ZN(n14606) );
  XNOR2_X1 U15910 ( .A(n14606), .B(n14661), .ZN(n14608) );
  AOI22_X1 U15911 ( .A1(n14895), .A2(n14659), .B1(n14607), .B2(n14876), .ZN(
        n14609) );
  XNOR2_X1 U15912 ( .A(n14608), .B(n14609), .ZN(n14681) );
  NAND2_X1 U15913 ( .A1(n14680), .A2(n14681), .ZN(n14612) );
  INV_X1 U15914 ( .A(n14608), .ZN(n14610) );
  NAND2_X1 U15915 ( .A1(n14610), .A2(n14609), .ZN(n14611) );
  OAI22_X1 U15916 ( .A1(n14884), .A2(n7189), .B1(n14870), .B2(n14613), .ZN(
        n14620) );
  NAND2_X1 U15917 ( .A1(n15092), .A2(n14614), .ZN(n14617) );
  NAND2_X1 U15918 ( .A1(n14896), .A2(n14615), .ZN(n14616) );
  NAND2_X1 U15919 ( .A1(n14617), .A2(n14616), .ZN(n14618) );
  XNOR2_X1 U15920 ( .A(n14618), .B(n14661), .ZN(n14619) );
  XOR2_X1 U15921 ( .A(n14620), .B(n14619), .Z(n14726) );
  INV_X1 U15922 ( .A(n14619), .ZN(n14622) );
  INV_X1 U15923 ( .A(n14620), .ZN(n14621) );
  NAND2_X1 U15924 ( .A1(n14622), .A2(n14621), .ZN(n14623) );
  NOR2_X1 U15925 ( .A1(n16041), .A2(n14862), .ZN(n14626) );
  AOI22_X1 U15926 ( .A1(n16029), .A2(n14896), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14624) );
  OAI21_X1 U15927 ( .B1(n14871), .B2(n14728), .A(n14624), .ZN(n14625) );
  AOI211_X1 U15928 ( .C1(n15087), .C2(n14731), .A(n14626), .B(n14625), .ZN(
        n14627) );
  OAI21_X1 U15929 ( .B1(n14628), .B2(n14733), .A(n14627), .ZN(P1_U3214) );
  INV_X1 U15930 ( .A(n14629), .ZN(n14630) );
  AOI21_X1 U15931 ( .B1(n14632), .B2(n14631), .A(n14630), .ZN(n14639) );
  OAI21_X1 U15932 ( .B1(n14728), .B2(n15050), .A(n14633), .ZN(n14634) );
  AOI21_X1 U15933 ( .B1(n16029), .B2(n14739), .A(n14634), .ZN(n14635) );
  OAI21_X1 U15934 ( .B1(n14636), .B2(n16041), .A(n14635), .ZN(n14637) );
  AOI21_X1 U15935 ( .B1(n15165), .B2(n14731), .A(n14637), .ZN(n14638) );
  OAI21_X1 U15936 ( .B1(n14639), .B2(n14733), .A(n14638), .ZN(P1_U3215) );
  XOR2_X1 U15937 ( .A(n14640), .B(n14641), .Z(n14646) );
  AOI22_X1 U15938 ( .A1(n16029), .A2(n14962), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14643) );
  NAND2_X1 U15939 ( .A1(n16031), .A2(n14925), .ZN(n14642) );
  OAI211_X1 U15940 ( .C1(n16041), .C2(n14928), .A(n14643), .B(n14642), .ZN(
        n14644) );
  AOI21_X1 U15941 ( .B1(n15117), .B2(n14731), .A(n14644), .ZN(n14645) );
  OAI21_X1 U15942 ( .B1(n14646), .B2(n14733), .A(n14645), .ZN(P1_U3216) );
  XOR2_X1 U15943 ( .A(n14648), .B(n14647), .Z(n14653) );
  NOR2_X1 U15944 ( .A1(n16041), .A2(n14989), .ZN(n14651) );
  AND2_X1 U15945 ( .A1(n16030), .A2(n15033), .ZN(n14649) );
  AOI21_X1 U15946 ( .B1(n14963), .B2(n15034), .A(n14649), .ZN(n14990) );
  INV_X1 U15947 ( .A(n14691), .ZN(n14712) );
  NAND2_X1 U15948 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14827)
         );
  OAI21_X1 U15949 ( .B1(n14990), .B2(n14712), .A(n14827), .ZN(n14650) );
  AOI211_X1 U15950 ( .C1(n15145), .C2(n14731), .A(n14651), .B(n14650), .ZN(
        n14652) );
  OAI21_X1 U15951 ( .B1(n14653), .B2(n14733), .A(n14652), .ZN(P1_U3219) );
  INV_X1 U15952 ( .A(n14654), .ZN(n14657) );
  INV_X1 U15953 ( .A(n14655), .ZN(n14656) );
  AOI22_X1 U15954 ( .A1(n15081), .A2(n9735), .B1(n14659), .B2(n14737), .ZN(
        n14664) );
  AOI22_X1 U15955 ( .A1(n15081), .A2(n14659), .B1(n14607), .B2(n14737), .ZN(
        n14662) );
  XNOR2_X1 U15956 ( .A(n14662), .B(n14661), .ZN(n14663) );
  XOR2_X1 U15957 ( .A(n14664), .B(n14663), .Z(n14665) );
  NOR2_X1 U15958 ( .A1(n16041), .A2(n14851), .ZN(n14668) );
  AOI22_X1 U15959 ( .A1(n16029), .A2(n14877), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14666) );
  OAI21_X1 U15960 ( .B1(n14840), .B2(n14728), .A(n14666), .ZN(n14667) );
  AOI211_X1 U15961 ( .C1(n15081), .C2(n14731), .A(n14668), .B(n14667), .ZN(
        n14669) );
  OAI21_X1 U15962 ( .B1(n14670), .B2(n14733), .A(n14669), .ZN(P1_U3220) );
  INV_X1 U15963 ( .A(n14671), .ZN(n14672) );
  AOI21_X1 U15964 ( .B1(n14674), .B2(n14673), .A(n14672), .ZN(n14679) );
  AOI22_X1 U15965 ( .A1(n16031), .A2(n14962), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14676) );
  NAND2_X1 U15966 ( .A1(n14963), .A2(n16029), .ZN(n14675) );
  OAI211_X1 U15967 ( .C1(n16041), .C2(n14964), .A(n14676), .B(n14675), .ZN(
        n14677) );
  AOI21_X1 U15968 ( .B1(n14961), .B2(n14731), .A(n14677), .ZN(n14678) );
  OAI21_X1 U15969 ( .B1(n14679), .B2(n14733), .A(n14678), .ZN(P1_U3223) );
  XOR2_X1 U15970 ( .A(n14681), .B(n14680), .Z(n14686) );
  NOR2_X1 U15971 ( .A1(n16041), .A2(n14897), .ZN(n14684) );
  AOI22_X1 U15972 ( .A1(n16029), .A2(n14925), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14682) );
  OAI21_X1 U15973 ( .B1(n14870), .B2(n14728), .A(n14682), .ZN(n14683) );
  AOI211_X1 U15974 ( .C1(n14895), .C2(n14731), .A(n14684), .B(n14683), .ZN(
        n14685) );
  OAI21_X1 U15975 ( .B1(n14686), .B2(n14733), .A(n14685), .ZN(P1_U3225) );
  XOR2_X1 U15976 ( .A(n14688), .B(n14687), .Z(n14695) );
  NAND2_X1 U15977 ( .A1(n14738), .A2(n15033), .ZN(n14690) );
  NAND2_X1 U15978 ( .A1(n14876), .A2(n15034), .ZN(n14689) );
  NAND2_X1 U15979 ( .A1(n14690), .A2(n14689), .ZN(n15106) );
  AOI22_X1 U15980 ( .A1(n15106), .A2(n14691), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14692) );
  OAI21_X1 U15981 ( .B1(n14908), .B2(n16041), .A(n14692), .ZN(n14693) );
  AOI21_X1 U15982 ( .B1(n15107), .B2(n14731), .A(n14693), .ZN(n14694) );
  OAI21_X1 U15983 ( .B1(n14695), .B2(n14733), .A(n14694), .ZN(P1_U3229) );
  AOI21_X1 U15984 ( .B1(n14697), .B2(n14696), .A(n14733), .ZN(n14699) );
  NAND2_X1 U15985 ( .A1(n14699), .A2(n14698), .ZN(n14705) );
  INV_X1 U15986 ( .A(n14977), .ZN(n14703) );
  AOI22_X1 U15987 ( .A1(n14976), .A2(n16031), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14700) );
  OAI21_X1 U15988 ( .B1(n14719), .B2(n14701), .A(n14700), .ZN(n14702) );
  AOI21_X1 U15989 ( .B1(n14703), .B2(n14722), .A(n14702), .ZN(n14704) );
  OAI211_X1 U15990 ( .C1(n15137), .C2(n16033), .A(n14705), .B(n14704), .ZN(
        P1_U3233) );
  OAI21_X1 U15991 ( .B1(n14708), .B2(n14707), .A(n14706), .ZN(n14709) );
  NAND2_X1 U15992 ( .A1(n14709), .A2(n16036), .ZN(n14715) );
  INV_X1 U15993 ( .A(n14710), .ZN(n14951) );
  AOI22_X1 U15994 ( .A1(n14976), .A2(n15033), .B1(n15034), .B2(n14738), .ZN(
        n14943) );
  INV_X1 U15995 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14711) );
  OAI22_X1 U15996 ( .A1(n14943), .A2(n14712), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14711), .ZN(n14713) );
  AOI21_X1 U15997 ( .B1(n14951), .B2(n14722), .A(n14713), .ZN(n14714) );
  OAI211_X1 U15998 ( .C1(n16033), .C2(n14954), .A(n14715), .B(n14714), .ZN(
        P1_U3235) );
  XOR2_X1 U15999 ( .A(n7542), .B(n14717), .Z(n14724) );
  NAND2_X1 U16000 ( .A1(n16029), .A2(n16001), .ZN(n14718) );
  NAND2_X1 U16001 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14792)
         );
  OAI211_X1 U16002 ( .C1(n14719), .C2(n14728), .A(n14718), .B(n14792), .ZN(
        n14721) );
  NOR2_X1 U16003 ( .A1(n15023), .A2(n16033), .ZN(n14720) );
  AOI211_X1 U16004 ( .C1(n14722), .C2(n15019), .A(n14721), .B(n14720), .ZN(
        n14723) );
  OAI21_X1 U16005 ( .B1(n14724), .B2(n14733), .A(n14723), .ZN(P1_U3238) );
  XOR2_X1 U16006 ( .A(n14726), .B(n14725), .Z(n14734) );
  NOR2_X1 U16007 ( .A1(n16041), .A2(n14881), .ZN(n14730) );
  AOI22_X1 U16008 ( .A1(n16029), .A2(n14876), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14727) );
  OAI21_X1 U16009 ( .B1(n14841), .B2(n14728), .A(n14727), .ZN(n14729) );
  AOI211_X1 U16010 ( .C1(n15092), .C2(n14731), .A(n14730), .B(n14729), .ZN(
        n14732) );
  OAI21_X1 U16011 ( .B1(n14734), .B2(n14733), .A(n14732), .ZN(P1_U3240) );
  MUX2_X1 U16012 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14830), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16013 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14735), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16014 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14736), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16015 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14737), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16016 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14877), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16017 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14896), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16018 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14876), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16019 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14925), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16020 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14738), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16021 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14962), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16022 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14976), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16023 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14963), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16024 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n15008), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16025 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n16030), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16026 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n16001), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16027 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n16028), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16028 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n16000), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16029 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n15978), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16030 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14739), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16031 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14740), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16032 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14741), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16033 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14742), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16034 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14743), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16035 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14744), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16036 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14745), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16037 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14746), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16038 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14747), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16039 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14748), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16040 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14749), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16041 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n10604), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16042 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9700), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16043 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14750), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U16044 ( .C1(n14753), .C2(n14752), .A(n15437), .B(n14751), .ZN(
        n14761) );
  OAI211_X1 U16045 ( .C1(n14756), .C2(n14755), .A(n14819), .B(n14754), .ZN(
        n14760) );
  NAND2_X1 U16046 ( .A1(n14795), .A2(n14757), .ZN(n14759) );
  AOI22_X1 U16047 ( .A1(n14791), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14758) );
  NAND4_X1 U16048 ( .A1(n14761), .A2(n14760), .A3(n14759), .A4(n14758), .ZN(
        P1_U3244) );
  OAI211_X1 U16049 ( .C1(n14764), .C2(n14763), .A(n15437), .B(n14762), .ZN(
        n14774) );
  NOR2_X1 U16050 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10606), .ZN(n14765) );
  AOI21_X1 U16051 ( .B1(n14791), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n14765), .ZN(
        n14773) );
  NAND2_X1 U16052 ( .A1(n14795), .A2(n14766), .ZN(n14772) );
  MUX2_X1 U16053 ( .A(n9955), .B(P1_REG2_REG_3__SCAN_IN), .S(n14766), .Z(
        n14769) );
  NAND3_X1 U16054 ( .A1(n14769), .A2(n14768), .A3(n14767), .ZN(n14770) );
  NAND3_X1 U16055 ( .A1(n14819), .A2(n14778), .A3(n14770), .ZN(n14771) );
  NAND4_X1 U16056 ( .A1(n14774), .A2(n14773), .A3(n14772), .A4(n14771), .ZN(
        P1_U3246) );
  INV_X1 U16057 ( .A(n14775), .ZN(n14790) );
  AOI22_X1 U16058 ( .A1(n14791), .A2(P1_ADDR_REG_4__SCAN_IN), .B1(
        P1_REG3_REG_4__SCAN_IN), .B2(P1_U3086), .ZN(n14789) );
  MUX2_X1 U16059 ( .A(n9958), .B(P1_REG2_REG_4__SCAN_IN), .S(n14782), .Z(
        n14776) );
  NAND3_X1 U16060 ( .A1(n14778), .A2(n14777), .A3(n14776), .ZN(n14779) );
  AND2_X1 U16061 ( .A1(n14780), .A2(n14779), .ZN(n14781) );
  AOI22_X1 U16062 ( .A1(n14795), .A2(n14782), .B1(n14819), .B2(n14781), .ZN(
        n14788) );
  INV_X1 U16063 ( .A(n14783), .ZN(n14784) );
  OAI211_X1 U16064 ( .C1(n14786), .C2(n14785), .A(n15437), .B(n14784), .ZN(
        n14787) );
  NAND4_X1 U16065 ( .A1(n14790), .A2(n14789), .A3(n14788), .A4(n14787), .ZN(
        P1_U3247) );
  INV_X1 U16066 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14793) );
  OAI21_X1 U16067 ( .B1(n15440), .B2(n14793), .A(n14792), .ZN(n14794) );
  AOI21_X1 U16068 ( .B1(n14814), .B2(n14795), .A(n14794), .ZN(n14807) );
  AOI21_X1 U16069 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n14797), .A(n14796), 
        .ZN(n14809) );
  XNOR2_X1 U16070 ( .A(n14808), .B(n14809), .ZN(n14798) );
  INV_X1 U16071 ( .A(n14798), .ZN(n14801) );
  NOR2_X1 U16072 ( .A1(n14799), .A2(n14798), .ZN(n14810) );
  INV_X1 U16073 ( .A(n14810), .ZN(n14800) );
  OAI211_X1 U16074 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n14801), .A(n15437), 
        .B(n14800), .ZN(n14806) );
  OAI21_X1 U16075 ( .B1(n15032), .B2(n14803), .A(n14802), .ZN(n14813) );
  XNOR2_X1 U16076 ( .A(n14808), .B(n14813), .ZN(n14804) );
  NAND2_X1 U16077 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14804), .ZN(n14816) );
  OAI211_X1 U16078 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n14804), .A(n14819), 
        .B(n14816), .ZN(n14805) );
  NAND3_X1 U16079 ( .A1(n14807), .A2(n14806), .A3(n14805), .ZN(P1_U3261) );
  NOR2_X1 U16080 ( .A1(n14809), .A2(n14808), .ZN(n14811) );
  NOR2_X1 U16081 ( .A1(n14811), .A2(n14810), .ZN(n14812) );
  XOR2_X1 U16082 ( .A(n14812), .B(P1_REG1_REG_19__SCAN_IN), .Z(n14824) );
  INV_X1 U16083 ( .A(n14824), .ZN(n14821) );
  NAND2_X1 U16084 ( .A1(n14814), .A2(n14813), .ZN(n14815) );
  NAND2_X1 U16085 ( .A1(n14816), .A2(n14815), .ZN(n14818) );
  XOR2_X1 U16086 ( .A(n14818), .B(n14817), .Z(n14822) );
  NAND2_X1 U16087 ( .A1(n14822), .A2(n14819), .ZN(n14820) );
  OAI211_X1 U16088 ( .C1(n14821), .C2(n14823), .A(n15432), .B(n14820), .ZN(
        n14826) );
  NAND2_X1 U16089 ( .A1(n14849), .A2(n15075), .ZN(n14834) );
  XNOR2_X1 U16090 ( .A(n14833), .B(n14828), .ZN(n15065) );
  NAND2_X1 U16091 ( .A1(n15065), .A2(n15018), .ZN(n14832) );
  NAND2_X1 U16092 ( .A1(n14830), .A2(n14829), .ZN(n15069) );
  NOR2_X1 U16093 ( .A1(n15020), .A2(n15069), .ZN(n14836) );
  AOI21_X1 U16094 ( .B1(n15020), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14836), 
        .ZN(n14831) );
  OAI211_X1 U16095 ( .C1(n15067), .C2(n15680), .A(n14832), .B(n14831), .ZN(
        P1_U3263) );
  INV_X1 U16096 ( .A(n14835), .ZN(n15071) );
  AOI21_X1 U16097 ( .B1(n14835), .B2(n14834), .A(n14833), .ZN(n15068) );
  NAND2_X1 U16098 ( .A1(n15068), .A2(n15018), .ZN(n14838) );
  AOI21_X1 U16099 ( .B1(n15020), .B2(P1_REG2_REG_30__SCAN_IN), .A(n14836), 
        .ZN(n14837) );
  OAI211_X1 U16100 ( .C1(n15071), .C2(n15680), .A(n14838), .B(n14837), .ZN(
        P1_U3264) );
  AOI21_X1 U16101 ( .B1(n14839), .B2(n14846), .A(n16016), .ZN(n14844) );
  OAI22_X1 U16102 ( .A1(n14841), .A2(n15049), .B1(n14840), .B2(n15051), .ZN(
        n14842) );
  AOI21_X1 U16103 ( .B1(n14844), .B2(n14843), .A(n14842), .ZN(n15084) );
  OAI21_X1 U16104 ( .B1(n14847), .B2(n14846), .A(n14845), .ZN(n15085) );
  INV_X1 U16105 ( .A(n15085), .ZN(n14848) );
  NAND2_X1 U16106 ( .A1(n14848), .A2(n15025), .ZN(n14856) );
  AOI21_X1 U16107 ( .B1(n15081), .B2(n14858), .A(n14849), .ZN(n15082) );
  INV_X1 U16108 ( .A(n15081), .ZN(n14850) );
  NOR2_X1 U16109 ( .A1(n14850), .A2(n15680), .ZN(n14854) );
  OAI22_X1 U16110 ( .A1(n15055), .A2(n14852), .B1(n14851), .B2(n15035), .ZN(
        n14853) );
  AOI211_X1 U16111 ( .C1(n15082), .C2(n15018), .A(n14854), .B(n14853), .ZN(
        n14855) );
  OAI211_X1 U16112 ( .C1(n15036), .C2(n15084), .A(n14856), .B(n14855), .ZN(
        P1_U3265) );
  INV_X1 U16113 ( .A(n14880), .ZN(n14860) );
  INV_X1 U16114 ( .A(n14858), .ZN(n14859) );
  AOI211_X1 U16115 ( .C1(n15087), .C2(n14860), .A(n16009), .B(n14859), .ZN(
        n15089) );
  NOR2_X1 U16116 ( .A1(n14861), .A2(n15680), .ZN(n14865) );
  OAI22_X1 U16117 ( .A1(n15055), .A2(n14863), .B1(n14862), .B2(n15035), .ZN(
        n14864) );
  AOI21_X1 U16118 ( .B1(n14868), .B2(n14867), .A(n14866), .ZN(n14869) );
  OAI222_X1 U16119 ( .A1(n15051), .A2(n14871), .B1(n15049), .B2(n14870), .C1(
        n14869), .C2(n16016), .ZN(n15090) );
  NAND2_X1 U16120 ( .A1(n15090), .A2(n15055), .ZN(n14872) );
  OAI211_X1 U16121 ( .C1(n15086), .C2(n14988), .A(n14873), .B(n14872), .ZN(
        P1_U3266) );
  XNOR2_X1 U16122 ( .A(n14875), .B(n14874), .ZN(n14878) );
  AOI222_X1 U16123 ( .A1(n14878), .A2(n15985), .B1(n14877), .B2(n15034), .C1(
        n14876), .C2(n15033), .ZN(n15095) );
  NOR2_X1 U16124 ( .A1(n14894), .A2(n14884), .ZN(n14879) );
  NOR2_X1 U16125 ( .A1(n14880), .A2(n14879), .ZN(n15093) );
  INV_X1 U16126 ( .A(n14881), .ZN(n14882) );
  AOI22_X1 U16127 ( .A1(n15020), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n14882), 
        .B2(n15678), .ZN(n14883) );
  OAI21_X1 U16128 ( .B1(n14884), .B2(n15680), .A(n14883), .ZN(n14888) );
  XNOR2_X1 U16129 ( .A(n14886), .B(n14885), .ZN(n15096) );
  NOR2_X1 U16130 ( .A1(n15096), .A2(n14988), .ZN(n14887) );
  AOI211_X1 U16131 ( .C1(n15093), .C2(n15018), .A(n14888), .B(n14887), .ZN(
        n14889) );
  OAI21_X1 U16132 ( .B1(n15020), .B2(n15095), .A(n14889), .ZN(P1_U3267) );
  OAI21_X1 U16133 ( .B1(n7276), .B2(n8000), .A(n14890), .ZN(n15104) );
  OAI21_X1 U16134 ( .B1(n14893), .B2(n14892), .A(n14891), .ZN(n15102) );
  AOI21_X1 U16135 ( .B1(n14895), .B2(n14906), .A(n14894), .ZN(n15097) );
  NAND2_X1 U16136 ( .A1(n15097), .A2(n15018), .ZN(n14900) );
  AOI22_X1 U16137 ( .A1(n15033), .A2(n14925), .B1(n14896), .B2(n15034), .ZN(
        n15098) );
  OAI22_X1 U16138 ( .A1(n15098), .A2(n15020), .B1(n14897), .B2(n15035), .ZN(
        n14898) );
  AOI21_X1 U16139 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(n15020), .A(n14898), 
        .ZN(n14899) );
  OAI211_X1 U16140 ( .C1(n15100), .C2(n15680), .A(n14900), .B(n14899), .ZN(
        n14901) );
  AOI21_X1 U16141 ( .B1(n15102), .B2(n14985), .A(n14901), .ZN(n14902) );
  OAI21_X1 U16142 ( .B1(n15104), .B2(n14988), .A(n14902), .ZN(P1_U3268) );
  INV_X1 U16143 ( .A(n14913), .ZN(n14904) );
  OAI21_X1 U16144 ( .B1(n14905), .B2(n14904), .A(n14903), .ZN(n15105) );
  INV_X1 U16145 ( .A(n15105), .ZN(n14921) );
  AOI21_X1 U16146 ( .B1(n14933), .B2(n15107), .A(n16009), .ZN(n14907) );
  NAND2_X1 U16147 ( .A1(n14907), .A2(n14906), .ZN(n15110) );
  INV_X1 U16148 ( .A(n15110), .ZN(n14918) );
  INV_X1 U16149 ( .A(n15106), .ZN(n14909) );
  OAI22_X1 U16150 ( .A1(n14909), .A2(n15020), .B1(n14908), .B2(n15035), .ZN(
        n14910) );
  AOI21_X1 U16151 ( .B1(P1_REG2_REG_24__SCAN_IN), .B2(n15020), .A(n14910), 
        .ZN(n14911) );
  OAI21_X1 U16152 ( .B1(n14912), .B2(n15680), .A(n14911), .ZN(n14916) );
  NOR2_X1 U16153 ( .A1(n14914), .A2(n14913), .ZN(n15109) );
  NOR3_X1 U16154 ( .A1(n15109), .A2(n15108), .A3(n15064), .ZN(n14915) );
  AOI211_X1 U16155 ( .C1(n14918), .C2(n14917), .A(n14916), .B(n14915), .ZN(
        n14919) );
  OAI21_X1 U16156 ( .B1(n14921), .B2(n14920), .A(n14919), .ZN(P1_U3269) );
  OAI21_X1 U16157 ( .B1(n14924), .B2(n14923), .A(n14922), .ZN(n15121) );
  NAND2_X1 U16158 ( .A1(n14925), .A2(n15034), .ZN(n14926) );
  OAI21_X1 U16159 ( .B1(n14927), .B2(n15049), .A(n14926), .ZN(n15116) );
  NOR2_X1 U16160 ( .A1(n15035), .A2(n14928), .ZN(n14929) );
  AOI21_X1 U16161 ( .B1(n15055), .B2(n15116), .A(n14929), .ZN(n14930) );
  OAI21_X1 U16162 ( .B1(n14931), .B2(n15055), .A(n14930), .ZN(n14936) );
  INV_X1 U16163 ( .A(n15117), .ZN(n14934) );
  INV_X1 U16164 ( .A(n14932), .ZN(n14949) );
  OAI21_X1 U16165 ( .B1(n14934), .B2(n14949), .A(n14933), .ZN(n15114) );
  NOR2_X1 U16166 ( .A1(n15114), .A2(n15681), .ZN(n14935) );
  AOI211_X1 U16167 ( .C1(n15061), .C2(n15117), .A(n14936), .B(n14935), .ZN(
        n14940) );
  XNOR2_X1 U16168 ( .A(n14938), .B(n14937), .ZN(n15118) );
  NAND2_X1 U16169 ( .A1(n15118), .A2(n14985), .ZN(n14939) );
  OAI211_X1 U16170 ( .C1(n15121), .C2(n14988), .A(n14940), .B(n14939), .ZN(
        P1_U3270) );
  OAI21_X1 U16171 ( .B1(n14942), .B2(n7333), .A(n14941), .ZN(n14945) );
  INV_X1 U16172 ( .A(n14943), .ZN(n14944) );
  AOI21_X1 U16173 ( .B1(n14945), .B2(n15985), .A(n14944), .ZN(n15126) );
  OAI21_X1 U16174 ( .B1(n14948), .B2(n14947), .A(n14946), .ZN(n15122) );
  INV_X1 U16175 ( .A(n14959), .ZN(n14950) );
  AOI21_X1 U16176 ( .B1(n15123), .B2(n14950), .A(n14949), .ZN(n15124) );
  NAND2_X1 U16177 ( .A1(n15124), .A2(n15018), .ZN(n14953) );
  AOI22_X1 U16178 ( .A1(n15020), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14951), 
        .B2(n15678), .ZN(n14952) );
  OAI211_X1 U16179 ( .C1(n15680), .C2(n14954), .A(n14953), .B(n14952), .ZN(
        n14955) );
  AOI21_X1 U16180 ( .B1(n15122), .B2(n15048), .A(n14955), .ZN(n14956) );
  OAI21_X1 U16181 ( .B1(n15020), .B2(n15126), .A(n14956), .ZN(P1_U3271) );
  XNOR2_X1 U16182 ( .A(n14958), .B(n14957), .ZN(n15135) );
  AOI21_X1 U16183 ( .B1(n14961), .B2(n14960), .A(n14959), .ZN(n15133) );
  AOI22_X1 U16184 ( .A1(n14963), .A2(n15033), .B1(n15034), .B2(n14962), .ZN(
        n15128) );
  OAI22_X1 U16185 ( .A1(n15128), .A2(n15036), .B1(n14964), .B2(n15035), .ZN(
        n14965) );
  AOI21_X1 U16186 ( .B1(P1_REG2_REG_21__SCAN_IN), .B2(n15036), .A(n14965), 
        .ZN(n14966) );
  OAI21_X1 U16187 ( .B1(n15129), .B2(n15680), .A(n14966), .ZN(n14971) );
  OAI21_X1 U16188 ( .B1(n14969), .B2(n14968), .A(n14967), .ZN(n15130) );
  NOR2_X1 U16189 ( .A1(n15130), .A2(n15064), .ZN(n14970) );
  AOI211_X1 U16190 ( .C1(n15133), .C2(n15018), .A(n14971), .B(n14970), .ZN(
        n14972) );
  OAI21_X1 U16191 ( .B1(n15135), .B2(n14988), .A(n14972), .ZN(P1_U3272) );
  OAI21_X1 U16192 ( .B1(n14974), .B2(n14984), .A(n14973), .ZN(n15143) );
  XNOR2_X1 U16193 ( .A(n15137), .B(n15000), .ZN(n15139) );
  AND2_X1 U16194 ( .A1(n15008), .A2(n15033), .ZN(n14975) );
  AOI21_X1 U16195 ( .B1(n14976), .B2(n15034), .A(n14975), .ZN(n15136) );
  OAI22_X1 U16196 ( .A1(n15136), .A2(n15036), .B1(n14977), .B2(n15035), .ZN(
        n14978) );
  AOI21_X1 U16197 ( .B1(P1_REG2_REG_20__SCAN_IN), .B2(n15036), .A(n14978), 
        .ZN(n14979) );
  OAI21_X1 U16198 ( .B1(n15137), .B2(n15680), .A(n14979), .ZN(n14980) );
  AOI21_X1 U16199 ( .B1(n15139), .B2(n15018), .A(n14980), .ZN(n14987) );
  INV_X1 U16200 ( .A(n14981), .ZN(n14982) );
  AOI21_X1 U16201 ( .B1(n14984), .B2(n14983), .A(n14982), .ZN(n15140) );
  NAND2_X1 U16202 ( .A1(n15140), .A2(n14985), .ZN(n14986) );
  OAI211_X1 U16203 ( .C1(n15143), .C2(n14988), .A(n14987), .B(n14986), .ZN(
        P1_U3273) );
  INV_X1 U16204 ( .A(n14989), .ZN(n14995) );
  INV_X1 U16205 ( .A(n14990), .ZN(n15144) );
  INV_X1 U16206 ( .A(n14991), .ZN(n14992) );
  AOI21_X1 U16207 ( .B1(n14997), .B2(n14993), .A(n14992), .ZN(n15151) );
  NOR2_X1 U16208 ( .A1(n15151), .A2(n15064), .ZN(n14994) );
  AOI211_X1 U16209 ( .C1(n15678), .C2(n14995), .A(n15144), .B(n14994), .ZN(
        n15004) );
  OAI21_X1 U16210 ( .B1(n14998), .B2(n14997), .A(n14996), .ZN(n15149) );
  NAND2_X1 U16211 ( .A1(n15017), .A2(n15145), .ZN(n14999) );
  NAND2_X1 U16212 ( .A1(n15000), .A2(n14999), .ZN(n15147) );
  AOI22_X1 U16213 ( .A1(n15145), .A2(n15061), .B1(n15020), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n15001) );
  OAI21_X1 U16214 ( .B1(n15147), .B2(n15681), .A(n15001), .ZN(n15002) );
  AOI21_X1 U16215 ( .B1(n15149), .B2(n15048), .A(n15002), .ZN(n15003) );
  OAI21_X1 U16216 ( .B1(n15036), .B2(n15004), .A(n15003), .ZN(P1_U3274) );
  OAI211_X1 U16217 ( .C1(n15007), .C2(n15006), .A(n15005), .B(n15985), .ZN(
        n15010) );
  AOI22_X1 U16218 ( .A1(n15008), .A2(n15034), .B1(n15033), .B2(n16001), .ZN(
        n15009) );
  AND2_X1 U16219 ( .A1(n15010), .A2(n15009), .ZN(n15156) );
  OAI21_X1 U16220 ( .B1(n15013), .B2(n15012), .A(n15011), .ZN(n15152) );
  INV_X1 U16221 ( .A(n15014), .ZN(n15015) );
  NAND2_X1 U16222 ( .A1(n15153), .A2(n15015), .ZN(n15016) );
  AND2_X1 U16223 ( .A1(n15017), .A2(n15016), .ZN(n15154) );
  NAND2_X1 U16224 ( .A1(n15154), .A2(n15018), .ZN(n15022) );
  AOI22_X1 U16225 ( .A1(n15020), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n15019), 
        .B2(n15678), .ZN(n15021) );
  OAI211_X1 U16226 ( .C1(n15023), .C2(n15680), .A(n15022), .B(n15021), .ZN(
        n15024) );
  AOI21_X1 U16227 ( .B1(n15152), .B2(n15025), .A(n15024), .ZN(n15026) );
  OAI21_X1 U16228 ( .B1(n15036), .B2(n15156), .A(n15026), .ZN(P1_U3275) );
  INV_X1 U16229 ( .A(n15031), .ZN(n15027) );
  XNOR2_X1 U16230 ( .A(n15028), .B(n15027), .ZN(n15164) );
  AOI21_X1 U16231 ( .B1(n15031), .B2(n15030), .A(n15029), .ZN(n15162) );
  XNOR2_X1 U16232 ( .A(n15057), .B(n16027), .ZN(n15160) );
  NOR2_X1 U16233 ( .A1(n15055), .A2(n15032), .ZN(n15038) );
  AOI22_X1 U16234 ( .A1(n16030), .A2(n15034), .B1(n16028), .B2(n15033), .ZN(
        n15159) );
  OAI22_X1 U16235 ( .A1(n15159), .A2(n15036), .B1(n16040), .B2(n15035), .ZN(
        n15037) );
  AOI211_X1 U16236 ( .C1(n16027), .C2(n15061), .A(n15038), .B(n15037), .ZN(
        n15039) );
  OAI21_X1 U16237 ( .B1(n15160), .B2(n15681), .A(n15039), .ZN(n15040) );
  AOI21_X1 U16238 ( .B1(n15162), .B2(n15048), .A(n15040), .ZN(n15041) );
  OAI21_X1 U16239 ( .B1(n15164), .B2(n15064), .A(n15041), .ZN(P1_U3276) );
  INV_X1 U16240 ( .A(n15042), .ZN(n15043) );
  AOI21_X1 U16241 ( .B1(n15046), .B2(n15044), .A(n15043), .ZN(n16017) );
  OAI21_X1 U16242 ( .B1(n15047), .B2(n15046), .A(n15045), .ZN(n16020) );
  NAND2_X1 U16243 ( .A1(n16020), .A2(n15048), .ZN(n15063) );
  OAI22_X1 U16244 ( .A1(n15052), .A2(n15051), .B1(n15050), .B2(n15049), .ZN(
        n16012) );
  INV_X1 U16245 ( .A(n16008), .ZN(n15053) );
  AOI22_X1 U16246 ( .A1(n16012), .A2(n15055), .B1(n15053), .B2(n15678), .ZN(
        n15054) );
  OAI21_X1 U16247 ( .B1(n15056), .B2(n15055), .A(n15054), .ZN(n15060) );
  OAI21_X1 U16248 ( .B1(n16003), .B2(n15058), .A(n15057), .ZN(n16010) );
  NOR2_X1 U16249 ( .A1(n16010), .A2(n15681), .ZN(n15059) );
  AOI211_X1 U16250 ( .C1(n15061), .C2(n16013), .A(n15060), .B(n15059), .ZN(
        n15062) );
  OAI211_X1 U16251 ( .C1(n16017), .C2(n15064), .A(n15063), .B(n15062), .ZN(
        P1_U3277) );
  NAND2_X1 U16252 ( .A1(n15065), .A2(n15796), .ZN(n15066) );
  OAI211_X1 U16253 ( .C1(n15067), .C2(n15954), .A(n15066), .B(n15069), .ZN(
        n15176) );
  MUX2_X1 U16254 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15176), .S(n15922), .Z(
        P1_U3559) );
  NAND2_X1 U16255 ( .A1(n15068), .A2(n15796), .ZN(n15070) );
  OAI211_X1 U16256 ( .C1(n15071), .C2(n15954), .A(n15070), .B(n15069), .ZN(
        n15177) );
  MUX2_X1 U16257 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15177), .S(n15922), .Z(
        P1_U3558) );
  NAND2_X1 U16258 ( .A1(n15072), .A2(n16019), .ZN(n15079) );
  OAI211_X1 U16259 ( .C1(n15075), .C2(n15954), .A(n15074), .B(n15073), .ZN(
        n15076) );
  AOI21_X1 U16260 ( .B1(n15077), .B2(n15796), .A(n15076), .ZN(n15078) );
  OAI211_X1 U16261 ( .C1(n16016), .C2(n15080), .A(n15079), .B(n15078), .ZN(
        n15178) );
  MUX2_X1 U16262 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n15178), .S(n15922), .Z(
        P1_U3557) );
  AOI22_X1 U16263 ( .A1(n15082), .A2(n15796), .B1(n16014), .B2(n15081), .ZN(
        n15083) );
  OAI211_X1 U16264 ( .C1(n15085), .C2(n15799), .A(n15084), .B(n15083), .ZN(
        n15179) );
  MUX2_X1 U16265 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15179), .S(n15922), .Z(
        P1_U3556) );
  MUX2_X1 U16266 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15180), .S(n15922), .Z(
        P1_U3555) );
  AOI22_X1 U16267 ( .A1(n15093), .A2(n15796), .B1(n16014), .B2(n15092), .ZN(
        n15094) );
  OAI211_X1 U16268 ( .C1(n15096), .C2(n15799), .A(n15095), .B(n15094), .ZN(
        n15181) );
  MUX2_X1 U16269 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15181), .S(n15922), .Z(
        P1_U3554) );
  NAND2_X1 U16270 ( .A1(n15097), .A2(n15796), .ZN(n15099) );
  OAI211_X1 U16271 ( .C1(n15100), .C2(n15954), .A(n15099), .B(n15098), .ZN(
        n15101) );
  AOI21_X1 U16272 ( .B1(n15102), .B2(n15985), .A(n15101), .ZN(n15103) );
  OAI21_X1 U16273 ( .B1(n15104), .B2(n15799), .A(n15103), .ZN(n15182) );
  MUX2_X1 U16274 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15182), .S(n15922), .Z(
        P1_U3553) );
  NAND2_X1 U16275 ( .A1(n15105), .A2(n16019), .ZN(n15113) );
  AOI21_X1 U16276 ( .B1(n15107), .B2(n16014), .A(n15106), .ZN(n15112) );
  OR3_X1 U16277 ( .A1(n15109), .A2(n15108), .A3(n16016), .ZN(n15111) );
  NAND4_X1 U16278 ( .A1(n15113), .A2(n15112), .A3(n15111), .A4(n15110), .ZN(
        n15183) );
  MUX2_X1 U16279 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15183), .S(n15922), .Z(
        P1_U3552) );
  NOR2_X1 U16280 ( .A1(n15114), .A2(n16009), .ZN(n15115) );
  AOI211_X1 U16281 ( .C1(n16014), .C2(n15117), .A(n15116), .B(n15115), .ZN(
        n15120) );
  NAND2_X1 U16282 ( .A1(n15118), .A2(n15985), .ZN(n15119) );
  OAI211_X1 U16283 ( .C1(n15121), .C2(n15799), .A(n15120), .B(n15119), .ZN(
        n15184) );
  MUX2_X1 U16284 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15184), .S(n15922), .Z(
        P1_U3551) );
  INV_X1 U16285 ( .A(n15122), .ZN(n15127) );
  AOI22_X1 U16286 ( .A1(n15124), .A2(n15796), .B1(n15123), .B2(n16014), .ZN(
        n15125) );
  OAI211_X1 U16287 ( .C1(n15127), .C2(n15799), .A(n15126), .B(n15125), .ZN(
        n15185) );
  MUX2_X1 U16288 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15185), .S(n15922), .Z(
        P1_U3550) );
  OAI21_X1 U16289 ( .B1(n15129), .B2(n15954), .A(n15128), .ZN(n15132) );
  NOR2_X1 U16290 ( .A1(n15130), .A2(n16016), .ZN(n15131) );
  AOI211_X1 U16291 ( .C1(n15796), .C2(n15133), .A(n15132), .B(n15131), .ZN(
        n15134) );
  OAI21_X1 U16292 ( .B1(n15135), .B2(n15799), .A(n15134), .ZN(n15186) );
  MUX2_X1 U16293 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15186), .S(n15922), .Z(
        P1_U3549) );
  OAI21_X1 U16294 ( .B1(n15137), .B2(n15954), .A(n15136), .ZN(n15138) );
  AOI21_X1 U16295 ( .B1(n15139), .B2(n15796), .A(n15138), .ZN(n15142) );
  NAND2_X1 U16296 ( .A1(n15140), .A2(n15985), .ZN(n15141) );
  OAI211_X1 U16297 ( .C1(n15143), .C2(n15799), .A(n15142), .B(n15141), .ZN(
        n15187) );
  MUX2_X1 U16298 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15187), .S(n15922), .Z(
        P1_U3548) );
  AOI21_X1 U16299 ( .B1(n15145), .B2(n16014), .A(n15144), .ZN(n15146) );
  OAI21_X1 U16300 ( .B1(n15147), .B2(n16009), .A(n15146), .ZN(n15148) );
  AOI21_X1 U16301 ( .B1(n15149), .B2(n16019), .A(n15148), .ZN(n15150) );
  OAI21_X1 U16302 ( .B1(n16016), .B2(n15151), .A(n15150), .ZN(n15188) );
  MUX2_X1 U16303 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15188), .S(n15922), .Z(
        P1_U3547) );
  INV_X1 U16304 ( .A(n15152), .ZN(n15157) );
  AOI22_X1 U16305 ( .A1(n15154), .A2(n15796), .B1(n16014), .B2(n15153), .ZN(
        n15155) );
  OAI211_X1 U16306 ( .C1(n15157), .C2(n15799), .A(n15156), .B(n15155), .ZN(
        n15189) );
  MUX2_X1 U16307 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15189), .S(n15922), .Z(
        P1_U3546) );
  NAND2_X1 U16308 ( .A1(n16027), .A2(n16014), .ZN(n15158) );
  OAI211_X1 U16309 ( .C1(n15160), .C2(n16009), .A(n15159), .B(n15158), .ZN(
        n15161) );
  AOI21_X1 U16310 ( .B1(n15162), .B2(n16019), .A(n15161), .ZN(n15163) );
  OAI21_X1 U16311 ( .B1(n16016), .B2(n15164), .A(n15163), .ZN(n15190) );
  MUX2_X1 U16312 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15190), .S(n15922), .Z(
        P1_U3545) );
  AOI22_X1 U16313 ( .A1(n15166), .A2(n15796), .B1(n16014), .B2(n15165), .ZN(
        n15167) );
  OAI211_X1 U16314 ( .C1(n15169), .C2(n15799), .A(n15168), .B(n15167), .ZN(
        n15191) );
  MUX2_X1 U16315 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15191), .S(n15922), .Z(
        P1_U3542) );
  OAI22_X1 U16316 ( .A1(n15171), .A2(n16009), .B1(n15170), .B2(n15954), .ZN(
        n15172) );
  AOI21_X1 U16317 ( .B1(n15173), .B2(n15881), .A(n15172), .ZN(n15174) );
  NAND2_X1 U16318 ( .A1(n15175), .A2(n15174), .ZN(n15192) );
  MUX2_X1 U16319 ( .A(n15192), .B(P1_REG1_REG_12__SCAN_IN), .S(n16021), .Z(
        P1_U3540) );
  MUX2_X1 U16320 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15176), .S(n15961), .Z(
        P1_U3527) );
  MUX2_X1 U16321 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15177), .S(n15961), .Z(
        P1_U3526) );
  MUX2_X1 U16322 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n15178), .S(n15961), .Z(
        P1_U3525) );
  MUX2_X1 U16323 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15179), .S(n15961), .Z(
        P1_U3524) );
  MUX2_X1 U16324 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15180), .S(n15961), .Z(
        P1_U3523) );
  MUX2_X1 U16325 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15181), .S(n15961), .Z(
        P1_U3522) );
  MUX2_X1 U16326 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15182), .S(n15961), .Z(
        P1_U3521) );
  MUX2_X1 U16327 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15183), .S(n15961), .Z(
        P1_U3520) );
  MUX2_X1 U16328 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15184), .S(n15961), .Z(
        P1_U3519) );
  MUX2_X1 U16329 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15185), .S(n15961), .Z(
        P1_U3518) );
  MUX2_X1 U16330 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15186), .S(n15961), .Z(
        P1_U3517) );
  MUX2_X1 U16331 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15187), .S(n15961), .Z(
        P1_U3516) );
  MUX2_X1 U16332 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15188), .S(n15961), .Z(
        P1_U3515) );
  MUX2_X1 U16333 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15189), .S(n15961), .Z(
        P1_U3513) );
  MUX2_X1 U16334 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15190), .S(n15961), .Z(
        P1_U3510) );
  MUX2_X1 U16335 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15191), .S(n15961), .Z(
        P1_U3501) );
  MUX2_X1 U16336 ( .A(n15192), .B(P1_REG0_REG_12__SCAN_IN), .S(n16023), .Z(
        P1_U3495) );
  MUX2_X1 U16337 ( .A(n15193), .B(P1_D_REG_1__SCAN_IN), .S(n15332), .Z(
        P1_U3446) );
  INV_X1 U16338 ( .A(n15194), .ZN(n15197) );
  NOR4_X1 U16339 ( .A1(n8885), .A2(P1_IR_REG_30__SCAN_IN), .A3(n8880), .A4(
        P1_U3086), .ZN(n15195) );
  AOI21_X1 U16340 ( .B1(n15212), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15195), 
        .ZN(n15196) );
  OAI21_X1 U16341 ( .B1(n15197), .B2(n15215), .A(n15196), .ZN(P1_U3324) );
  OAI222_X1 U16342 ( .A1(P1_U3086), .A2(n15200), .B1(n15215), .B2(n15199), 
        .C1(n15198), .C2(n15210), .ZN(P1_U3326) );
  OAI222_X1 U16343 ( .A1(P1_U3086), .A2(n15203), .B1(n15215), .B2(n15202), 
        .C1(n15201), .C2(n15210), .ZN(P1_U3329) );
  AOI22_X1 U16344 ( .A1(n15204), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n15212), .ZN(n15205) );
  OAI21_X1 U16345 ( .B1(n15206), .B2(n15215), .A(n15205), .ZN(P1_U3330) );
  INV_X1 U16346 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n15209) );
  OAI222_X1 U16347 ( .A1(n15210), .A2(n15209), .B1(n15215), .B2(n15208), .C1(
        P1_U3086), .C2(n15207), .ZN(P1_U3331) );
  INV_X1 U16348 ( .A(n15211), .ZN(n15216) );
  NAND2_X1 U16349 ( .A1(n15212), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n15214) );
  OAI211_X1 U16350 ( .C1(n15216), .C2(n15215), .A(n15214), .B(n15213), .ZN(
        P1_U3332) );
  MUX2_X1 U16351 ( .A(n15218), .B(n15217), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16352 ( .A(n15219), .ZN(n15220) );
  MUX2_X1 U16353 ( .A(n15220), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16354 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15250) );
  NOR2_X1 U16355 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n15250), .ZN(n15221) );
  AOI21_X1 U16356 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n15250), .A(n15221), 
        .ZN(n15257) );
  INV_X1 U16357 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15246) );
  XOR2_X1 U16358 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n15309) );
  INV_X1 U16359 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15244) );
  XOR2_X1 U16360 ( .A(n15244), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n15304) );
  INV_X1 U16361 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n15241) );
  INV_X1 U16362 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n15239) );
  XOR2_X1 U16363 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n15239), .Z(n15297) );
  XOR2_X1 U16364 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n15237), .Z(n15293) );
  INV_X1 U16365 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15232) );
  AND2_X1 U16366 ( .A1(n15284), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n15231) );
  XOR2_X1 U16367 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n15226), .Z(n15267) );
  INV_X1 U16368 ( .A(n15271), .ZN(n15222) );
  NAND2_X1 U16369 ( .A1(n15222), .A2(n15269), .ZN(n15223) );
  OAI21_X1 U16370 ( .B1(P1_ADDR_REG_1__SCAN_IN), .B2(n15224), .A(n15223), .ZN(
        n15268) );
  NAND2_X1 U16371 ( .A1(n15267), .A2(n15268), .ZN(n15225) );
  NAND2_X1 U16372 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n15227), .ZN(n15228) );
  AOI22_X1 U16373 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n15262), .B1(n15263), 
        .B2(n15229), .ZN(n15279) );
  OR2_X1 U16374 ( .A1(n15278), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n15230) );
  AOI22_X1 U16375 ( .A1(n15279), .A2(n15230), .B1(P1_ADDR_REG_5__SCAN_IN), 
        .B2(n15278), .ZN(n15285) );
  OAI22_X1 U16376 ( .A1(n15231), .A2(n15285), .B1(P3_ADDR_REG_6__SCAN_IN), 
        .B2(n15284), .ZN(n15233) );
  NOR2_X1 U16377 ( .A1(n15232), .A2(n15233), .ZN(n15235) );
  XOR2_X1 U16378 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n15233), .Z(n15289) );
  NOR2_X1 U16379 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n15289), .ZN(n15234) );
  NAND2_X1 U16380 ( .A1(n15293), .A2(n15292), .ZN(n15236) );
  NAND2_X1 U16381 ( .A1(n15297), .A2(n15298), .ZN(n15238) );
  XNOR2_X1 U16382 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n15241), .ZN(n15260) );
  NOR2_X1 U16383 ( .A1(n15261), .A2(n15260), .ZN(n15240) );
  INV_X1 U16384 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15300) );
  OR2_X1 U16385 ( .A1(n15300), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n15242) );
  AOI22_X1 U16386 ( .A1(n15301), .A2(n15242), .B1(P1_ADDR_REG_11__SCAN_IN), 
        .B2(n15300), .ZN(n15303) );
  NAND2_X1 U16387 ( .A1(n15304), .A2(n15303), .ZN(n15243) );
  NOR2_X1 U16388 ( .A1(n15309), .A2(n15308), .ZN(n15245) );
  AOI21_X1 U16389 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n15246), .A(n15245), 
        .ZN(n15259) );
  XNOR2_X1 U16390 ( .A(n15248), .B(P1_ADDR_REG_14__SCAN_IN), .ZN(n15258) );
  NOR2_X1 U16391 ( .A1(n15259), .A2(n15258), .ZN(n15247) );
  AOI21_X1 U16392 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n15248), .A(n15247), 
        .ZN(n15256) );
  NAND2_X1 U16393 ( .A1(n15257), .A2(n15256), .ZN(n15249) );
  INV_X1 U16394 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15252) );
  NOR2_X1 U16395 ( .A1(n15251), .A2(n15252), .ZN(n15254) );
  XNOR2_X1 U16396 ( .A(n15252), .B(n15251), .ZN(n15255) );
  NOR2_X1 U16397 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n15255), .ZN(n15253) );
  NOR2_X1 U16398 ( .A1(n15254), .A2(n15253), .ZN(n15316) );
  XOR2_X1 U16399 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n15316), .Z(n15317) );
  XOR2_X1 U16400 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n15317), .Z(n15313) );
  AND2_X1 U16401 ( .A1(n15313), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n15314) );
  XOR2_X1 U16402 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n15255), .Z(n15312) );
  XOR2_X1 U16403 ( .A(n15257), .B(n15256), .Z(n15488) );
  XNOR2_X1 U16404 ( .A(n15259), .B(n15258), .ZN(n15485) );
  XOR2_X1 U16405 ( .A(n15261), .B(n15260), .Z(n15468) );
  INV_X1 U16406 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n15375) );
  NOR2_X1 U16407 ( .A1(n15264), .A2(n15375), .ZN(n15277) );
  XOR2_X1 U16408 ( .A(n15264), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n15452) );
  XOR2_X1 U16409 ( .A(n15268), .B(n15267), .Z(n15445) );
  XNOR2_X1 U16410 ( .A(n15271), .B(n15269), .ZN(n15270) );
  NOR2_X1 U16411 ( .A1(n15270), .A2(n7505), .ZN(n15273) );
  OAI21_X1 U16412 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n15272), .A(n15271), .ZN(
        n15442) );
  NAND2_X1 U16413 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15442), .ZN(n15508) );
  NAND2_X1 U16414 ( .A1(n15445), .A2(n15444), .ZN(n15443) );
  NAND2_X1 U16415 ( .A1(n15274), .A2(n15275), .ZN(n15276) );
  INV_X1 U16416 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15448) );
  NAND2_X1 U16417 ( .A1(n15449), .A2(n15448), .ZN(n15447) );
  NAND2_X1 U16418 ( .A1(n15276), .A2(n15447), .ZN(n15451) );
  XOR2_X1 U16419 ( .A(n15278), .B(P1_ADDR_REG_5__SCAN_IN), .Z(n15280) );
  XNOR2_X1 U16420 ( .A(n15280), .B(n15279), .ZN(n15282) );
  NOR2_X1 U16421 ( .A1(n15281), .A2(n15282), .ZN(n15283) );
  XOR2_X1 U16422 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(n15284), .Z(n15286) );
  XOR2_X1 U16423 ( .A(n15286), .B(n15285), .Z(n15287) );
  NAND2_X1 U16424 ( .A1(n15288), .A2(n15287), .ZN(n15504) );
  INV_X1 U16425 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n15506) );
  NOR2_X1 U16426 ( .A1(n15290), .A2(n7745), .ZN(n15291) );
  XOR2_X1 U16427 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n15289), .Z(n15458) );
  XNOR2_X1 U16428 ( .A(n15293), .B(n15292), .ZN(n15295) );
  NOR2_X1 U16429 ( .A1(n15294), .A2(n15295), .ZN(n15296) );
  XNOR2_X1 U16430 ( .A(n15295), .B(n15294), .ZN(n15461) );
  XNOR2_X1 U16431 ( .A(n15298), .B(n15297), .ZN(n15464) );
  NAND2_X1 U16432 ( .A1(n15468), .A2(n15467), .ZN(n15299) );
  XOR2_X1 U16433 ( .A(n15300), .B(P1_ADDR_REG_11__SCAN_IN), .Z(n15302) );
  XNOR2_X1 U16434 ( .A(n15302), .B(n15301), .ZN(n15472) );
  XOR2_X1 U16435 ( .A(n15304), .B(n15303), .Z(n15305) );
  NAND2_X1 U16436 ( .A1(n15306), .A2(n15305), .ZN(n15307) );
  INV_X1 U16437 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15477) );
  XNOR2_X1 U16438 ( .A(n15309), .B(n15308), .ZN(n15480) );
  NAND2_X1 U16439 ( .A1(n15485), .A2(n15484), .ZN(n15483) );
  INV_X1 U16440 ( .A(n15492), .ZN(n15493) );
  INV_X1 U16441 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15495) );
  NAND2_X1 U16442 ( .A1(n15493), .A2(n15491), .ZN(n15498) );
  INV_X1 U16443 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15412) );
  XOR2_X1 U16444 ( .A(n15313), .B(n15412), .Z(n15497) );
  INV_X1 U16445 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15315) );
  NOR2_X1 U16446 ( .A1(n15316), .A2(n15315), .ZN(n15319) );
  NOR2_X1 U16447 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n15317), .ZN(n15318) );
  NOR2_X1 U16448 ( .A1(n15319), .A2(n15318), .ZN(n15323) );
  INV_X1 U16449 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15325) );
  NAND2_X1 U16450 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n15325), .ZN(n15320) );
  OAI21_X1 U16451 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15325), .A(n15320), 
        .ZN(n15322) );
  XNOR2_X1 U16452 ( .A(n15323), .B(n15322), .ZN(n15500) );
  NAND2_X1 U16453 ( .A1(n15501), .A2(n15500), .ZN(n15321) );
  AOI21_X1 U16454 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n15321), .A(n15499), 
        .ZN(n15331) );
  NOR2_X1 U16455 ( .A1(n15323), .A2(n15322), .ZN(n15324) );
  AOI21_X1 U16456 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15325), .A(n15324), 
        .ZN(n15329) );
  XNOR2_X1 U16457 ( .A(n15326), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n15327) );
  XNOR2_X1 U16458 ( .A(n15327), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n15328) );
  XNOR2_X1 U16459 ( .A(n15329), .B(n15328), .ZN(n15330) );
  XNOR2_X1 U16460 ( .A(n15331), .B(n15330), .ZN(SUB_1596_U4) );
  AND2_X1 U16461 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15332), .ZN(P1_U3323) );
  AND2_X1 U16462 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15332), .ZN(P1_U3322) );
  AND2_X1 U16463 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15332), .ZN(P1_U3321) );
  AND2_X1 U16464 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15332), .ZN(P1_U3320) );
  AND2_X1 U16465 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15332), .ZN(P1_U3319) );
  AND2_X1 U16466 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15332), .ZN(P1_U3318) );
  AND2_X1 U16467 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15332), .ZN(P1_U3317) );
  AND2_X1 U16468 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15332), .ZN(P1_U3316) );
  AND2_X1 U16469 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15332), .ZN(P1_U3315) );
  AND2_X1 U16470 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15332), .ZN(P1_U3314) );
  AND2_X1 U16471 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15332), .ZN(P1_U3313) );
  AND2_X1 U16472 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15332), .ZN(P1_U3312) );
  AND2_X1 U16473 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15332), .ZN(P1_U3311) );
  AND2_X1 U16474 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15332), .ZN(P1_U3310) );
  AND2_X1 U16475 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15332), .ZN(P1_U3309) );
  AND2_X1 U16476 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15332), .ZN(P1_U3308) );
  AND2_X1 U16477 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15332), .ZN(P1_U3307) );
  AND2_X1 U16478 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15332), .ZN(P1_U3306) );
  AND2_X1 U16479 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15332), .ZN(P1_U3305) );
  AND2_X1 U16480 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15332), .ZN(P1_U3304) );
  AND2_X1 U16481 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15332), .ZN(P1_U3303) );
  AND2_X1 U16482 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15332), .ZN(P1_U3302) );
  AND2_X1 U16483 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15332), .ZN(P1_U3301) );
  AND2_X1 U16484 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15332), .ZN(P1_U3300) );
  AND2_X1 U16485 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15332), .ZN(P1_U3299) );
  AND2_X1 U16486 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15332), .ZN(P1_U3298) );
  AND2_X1 U16487 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15332), .ZN(P1_U3297) );
  AND2_X1 U16488 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15332), .ZN(P1_U3296) );
  AND2_X1 U16489 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15332), .ZN(P1_U3295) );
  AND2_X1 U16490 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15332), .ZN(P1_U3294) );
  INV_X1 U16491 ( .A(n15340), .ZN(n15337) );
  AOI21_X1 U16492 ( .B1(n15334), .B2(n15337), .A(n15333), .ZN(P2_U3417) );
  AND2_X1 U16493 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15336), .ZN(P2_U3295) );
  AND2_X1 U16494 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15336), .ZN(P2_U3294) );
  AND2_X1 U16495 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15336), .ZN(P2_U3293) );
  AND2_X1 U16496 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15336), .ZN(P2_U3292) );
  AND2_X1 U16497 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15336), .ZN(P2_U3291) );
  AND2_X1 U16498 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15336), .ZN(P2_U3290) );
  AND2_X1 U16499 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15336), .ZN(P2_U3289) );
  AND2_X1 U16500 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15336), .ZN(P2_U3288) );
  AND2_X1 U16501 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15336), .ZN(P2_U3287) );
  AND2_X1 U16502 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15336), .ZN(P2_U3286) );
  AND2_X1 U16503 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15336), .ZN(P2_U3285) );
  AND2_X1 U16504 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15336), .ZN(P2_U3284) );
  AND2_X1 U16505 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15336), .ZN(P2_U3283) );
  AND2_X1 U16506 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15336), .ZN(P2_U3282) );
  AND2_X1 U16507 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15336), .ZN(P2_U3281) );
  AND2_X1 U16508 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15336), .ZN(P2_U3280) );
  AND2_X1 U16509 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15336), .ZN(P2_U3279) );
  AND2_X1 U16510 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15336), .ZN(P2_U3278) );
  AND2_X1 U16511 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15336), .ZN(P2_U3277) );
  AND2_X1 U16512 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15336), .ZN(P2_U3276) );
  AND2_X1 U16513 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15336), .ZN(P2_U3275) );
  AND2_X1 U16514 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15336), .ZN(P2_U3274) );
  AND2_X1 U16515 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15336), .ZN(P2_U3273) );
  AND2_X1 U16516 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15336), .ZN(P2_U3272) );
  AND2_X1 U16517 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15336), .ZN(P2_U3271) );
  AND2_X1 U16518 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15336), .ZN(P2_U3270) );
  AND2_X1 U16519 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15336), .ZN(P2_U3269) );
  AND2_X1 U16520 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15336), .ZN(P2_U3268) );
  AND2_X1 U16521 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15336), .ZN(P2_U3267) );
  AND2_X1 U16522 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15336), .ZN(P2_U3266) );
  NOR2_X1 U16523 ( .A1(n15341), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U16524 ( .A1(P3_U3897), .A2(n15663), .ZN(P3_U3150) );
  AOI22_X1 U16525 ( .A1(n15340), .A2(n15339), .B1(n15338), .B2(n15337), .ZN(
        P2_U3416) );
  AOI22_X1 U16526 ( .A1(n15341), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n15352) );
  NAND2_X1 U16527 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15344) );
  AOI211_X1 U16528 ( .C1(n15344), .C2(n15343), .A(n15342), .B(n15406), .ZN(
        n15349) );
  NAND2_X1 U16529 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15347) );
  AOI211_X1 U16530 ( .C1(n15347), .C2(n15346), .A(n15345), .B(n15387), .ZN(
        n15348) );
  AOI211_X1 U16531 ( .C1(n15421), .C2(n15350), .A(n15349), .B(n15348), .ZN(
        n15351) );
  NAND2_X1 U16532 ( .A1(n15352), .A2(n15351), .ZN(P2_U3215) );
  AOI211_X1 U16533 ( .C1(n15355), .C2(n15354), .A(n15353), .B(n15406), .ZN(
        n15360) );
  AOI211_X1 U16534 ( .C1(n15358), .C2(n15357), .A(n15356), .B(n15387), .ZN(
        n15359) );
  AOI211_X1 U16535 ( .C1(n15421), .C2(n15361), .A(n15360), .B(n15359), .ZN(
        n15363) );
  NAND2_X1 U16536 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n15362) );
  OAI211_X1 U16537 ( .C1(n15427), .C2(n15448), .A(n15363), .B(n15362), .ZN(
        P2_U3217) );
  AOI211_X1 U16538 ( .C1(n15366), .C2(n15365), .A(n15364), .B(n15406), .ZN(
        n15371) );
  AOI211_X1 U16539 ( .C1(n15369), .C2(n15368), .A(n15367), .B(n15387), .ZN(
        n15370) );
  AOI211_X1 U16540 ( .C1(n15421), .C2(n15372), .A(n15371), .B(n15370), .ZN(
        n15374) );
  NAND2_X1 U16541 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n15373) );
  OAI211_X1 U16542 ( .C1(n15427), .C2(n15375), .A(n15374), .B(n15373), .ZN(
        P2_U3218) );
  AOI211_X1 U16543 ( .C1(n15378), .C2(n15377), .A(n15387), .B(n15376), .ZN(
        n15383) );
  AOI211_X1 U16544 ( .C1(n15381), .C2(n15380), .A(n15406), .B(n15379), .ZN(
        n15382) );
  AOI211_X1 U16545 ( .C1(n15421), .C2(n15384), .A(n15383), .B(n15382), .ZN(
        n15386) );
  NAND2_X1 U16546 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n15385) );
  OAI211_X1 U16547 ( .C1(n15427), .C2(n15506), .A(n15386), .B(n15385), .ZN(
        P2_U3220) );
  AOI211_X1 U16548 ( .C1(n15390), .C2(n15389), .A(n15388), .B(n15387), .ZN(
        n15391) );
  AOI211_X1 U16549 ( .C1(n15393), .C2(n15421), .A(n15392), .B(n15391), .ZN(
        n15397) );
  OAI211_X1 U16550 ( .C1(n15395), .C2(P2_REG2_REG_15__SCAN_IN), .A(n15423), 
        .B(n15394), .ZN(n15396) );
  OAI211_X1 U16551 ( .C1(n15427), .C2(n7742), .A(n15397), .B(n15396), .ZN(
        P2_U3229) );
  OAI211_X1 U16552 ( .C1(n15400), .C2(n15399), .A(n15419), .B(n15398), .ZN(
        n15401) );
  INV_X1 U16553 ( .A(n15401), .ZN(n15402) );
  AOI211_X1 U16554 ( .C1(n15404), .C2(n15421), .A(n15403), .B(n15402), .ZN(
        n15411) );
  AOI211_X1 U16555 ( .C1(n15408), .C2(n15407), .A(n15406), .B(n15405), .ZN(
        n15409) );
  INV_X1 U16556 ( .A(n15409), .ZN(n15410) );
  OAI211_X1 U16557 ( .C1(n15427), .C2(n15412), .A(n15411), .B(n15410), .ZN(
        P2_U3231) );
  OAI21_X1 U16558 ( .B1(n15415), .B2(n15414), .A(n15413), .ZN(n15424) );
  OAI21_X1 U16559 ( .B1(n15418), .B2(n15417), .A(n15416), .ZN(n15420) );
  AOI222_X1 U16560 ( .A1(n15424), .A2(n15423), .B1(n15422), .B2(n15421), .C1(
        n15420), .C2(n15419), .ZN(n15426) );
  OAI211_X1 U16561 ( .C1(n15477), .C2(n15427), .A(n15426), .B(n15425), .ZN(
        P2_U3226) );
  INV_X1 U16562 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15441) );
  OAI21_X1 U16563 ( .B1(n15429), .B2(n15995), .A(n15428), .ZN(n15438) );
  AOI21_X1 U16564 ( .B1(n15431), .B2(P1_REG2_REG_15__SCAN_IN), .A(n15430), 
        .ZN(n15435) );
  OAI22_X1 U16565 ( .A1(n15435), .A2(n15434), .B1(n15433), .B2(n15432), .ZN(
        n15436) );
  AOI21_X1 U16566 ( .B1(n15438), .B2(n15437), .A(n15436), .ZN(n15439) );
  NAND2_X1 U16567 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n15982)
         );
  OAI211_X1 U16568 ( .C1(n15441), .C2(n15440), .A(n15439), .B(n15982), .ZN(
        P1_U3258) );
  XOR2_X1 U16569 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15442), .Z(SUB_1596_U53) );
  OAI21_X1 U16570 ( .B1(n15445), .B2(n15444), .A(n15443), .ZN(n15446) );
  XNOR2_X1 U16571 ( .A(n15446), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  OAI21_X1 U16572 ( .B1(n15449), .B2(n15448), .A(n15447), .ZN(SUB_1596_U60) );
  AOI21_X1 U16573 ( .B1(n15452), .B2(n15451), .A(n15450), .ZN(SUB_1596_U59) );
  AOI21_X1 U16574 ( .B1(n15455), .B2(n15454), .A(n15453), .ZN(SUB_1596_U58) );
  AOI21_X1 U16575 ( .B1(n15458), .B2(n15457), .A(n15456), .ZN(SUB_1596_U56) );
  AOI21_X1 U16576 ( .B1(n15461), .B2(n15460), .A(n15459), .ZN(SUB_1596_U55) );
  OAI21_X1 U16577 ( .B1(n15464), .B2(n15463), .A(n15462), .ZN(n15465) );
  XOR2_X1 U16578 ( .A(n15465), .B(n7743), .Z(SUB_1596_U54) );
  AOI21_X1 U16579 ( .B1(n15468), .B2(n15467), .A(n15466), .ZN(n15469) );
  XNOR2_X1 U16580 ( .A(n15470), .B(n15469), .ZN(SUB_1596_U70) );
  AOI21_X1 U16581 ( .B1(n15473), .B2(n15472), .A(n15471), .ZN(n15474) );
  XNOR2_X1 U16582 ( .A(n15475), .B(n15474), .ZN(SUB_1596_U69) );
  OAI21_X1 U16583 ( .B1(n15478), .B2(n15477), .A(n15476), .ZN(SUB_1596_U68) );
  OAI21_X1 U16584 ( .B1(n15481), .B2(n15480), .A(n15479), .ZN(n15482) );
  XNOR2_X1 U16585 ( .A(n15482), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  OAI21_X1 U16586 ( .B1(n15485), .B2(n15484), .A(n15483), .ZN(n15486) );
  XNOR2_X1 U16587 ( .A(n15486), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI21_X1 U16588 ( .B1(n15489), .B2(n15488), .A(n15487), .ZN(n15490) );
  XOR2_X1 U16589 ( .A(n15490), .B(n7742), .Z(SUB_1596_U65) );
  OAI222_X1 U16590 ( .A1(n15495), .A2(n15494), .B1(n15495), .B2(n15493), .C1(
        n15492), .C2(n15491), .ZN(SUB_1596_U64) );
  AOI21_X1 U16591 ( .B1(n15498), .B2(n15497), .A(n15496), .ZN(SUB_1596_U63) );
  INV_X1 U16592 ( .A(n15504), .ZN(n15503) );
  OAI222_X1 U16593 ( .A1(n15506), .A2(n15505), .B1(n15506), .B2(n15504), .C1(
        n15503), .C2(n15502), .ZN(SUB_1596_U57) );
  AOI21_X1 U16594 ( .B1(n15509), .B2(n15508), .A(n15507), .ZN(SUB_1596_U5) );
  AOI21_X1 U16595 ( .B1(n11406), .B2(n15511), .A(n15510), .ZN(n15526) );
  INV_X1 U16596 ( .A(n15512), .ZN(n15513) );
  OAI21_X1 U16597 ( .B1(n15593), .B2(n7737), .A(n15513), .ZN(n15520) );
  INV_X1 U16598 ( .A(n15514), .ZN(n15515) );
  NAND3_X1 U16599 ( .A1(n15517), .A2(n15516), .A3(n15515), .ZN(n15518) );
  AOI21_X1 U16600 ( .B1(n15536), .B2(n15518), .A(n15659), .ZN(n15519) );
  AOI211_X1 U16601 ( .C1(n15602), .C2(n15521), .A(n15520), .B(n15519), .ZN(
        n15525) );
  XNOR2_X1 U16602 ( .A(n15522), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n15523) );
  NAND2_X1 U16603 ( .A1(n15667), .A2(n15523), .ZN(n15524) );
  OAI211_X1 U16604 ( .C1(n15526), .C2(n15671), .A(n15525), .B(n15524), .ZN(
        P3_U3185) );
  AOI21_X1 U16605 ( .B1(n15529), .B2(n15528), .A(n15527), .ZN(n15548) );
  INV_X1 U16606 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15532) );
  INV_X1 U16607 ( .A(n15530), .ZN(n15531) );
  OAI21_X1 U16608 ( .B1(n15593), .B2(n15532), .A(n15531), .ZN(n15539) );
  INV_X1 U16609 ( .A(n15533), .ZN(n15534) );
  NAND3_X1 U16610 ( .A1(n15536), .A2(n15535), .A3(n15534), .ZN(n15537) );
  AOI21_X1 U16611 ( .B1(n15555), .B2(n15537), .A(n15659), .ZN(n15538) );
  AOI211_X1 U16612 ( .C1(n15602), .C2(n15540), .A(n15539), .B(n15538), .ZN(
        n15547) );
  INV_X1 U16613 ( .A(n15541), .ZN(n15542) );
  AOI21_X1 U16614 ( .B1(n15544), .B2(n15543), .A(n15542), .ZN(n15545) );
  OR2_X1 U16615 ( .A1(n15583), .A2(n15545), .ZN(n15546) );
  OAI211_X1 U16616 ( .C1(n15548), .C2(n15671), .A(n15547), .B(n15546), .ZN(
        P3_U3186) );
  AOI21_X1 U16617 ( .B1(n15551), .B2(n15550), .A(n15549), .ZN(n15565) );
  INV_X1 U16618 ( .A(n15552), .ZN(n15553) );
  NAND3_X1 U16619 ( .A1(n15555), .A2(n15554), .A3(n15553), .ZN(n15556) );
  AOI21_X1 U16620 ( .B1(n15575), .B2(n15556), .A(n15659), .ZN(n15560) );
  AOI21_X1 U16621 ( .B1(n15663), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n15557), .ZN(
        n15558) );
  OAI21_X1 U16622 ( .B1(n15657), .B2(n7678), .A(n15558), .ZN(n15559) );
  NOR2_X1 U16623 ( .A1(n15560), .A2(n15559), .ZN(n15564) );
  XNOR2_X1 U16624 ( .A(n15561), .B(P3_REG1_REG_5__SCAN_IN), .ZN(n15562) );
  NAND2_X1 U16625 ( .A1(n15667), .A2(n15562), .ZN(n15563) );
  OAI211_X1 U16626 ( .C1(n15565), .C2(n15671), .A(n15564), .B(n15563), .ZN(
        P3_U3187) );
  AOI21_X1 U16627 ( .B1(n15568), .B2(n15567), .A(n15566), .ZN(n15587) );
  INV_X1 U16628 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15571) );
  INV_X1 U16629 ( .A(n15569), .ZN(n15570) );
  OAI21_X1 U16630 ( .B1(n15593), .B2(n15571), .A(n15570), .ZN(n15578) );
  INV_X1 U16631 ( .A(n15572), .ZN(n15573) );
  NAND3_X1 U16632 ( .A1(n15575), .A2(n15574), .A3(n15573), .ZN(n15576) );
  AOI21_X1 U16633 ( .B1(n15597), .B2(n15576), .A(n15659), .ZN(n15577) );
  AOI211_X1 U16634 ( .C1(n15602), .C2(n15579), .A(n15578), .B(n15577), .ZN(
        n15586) );
  AOI21_X1 U16635 ( .B1(n15582), .B2(n15581), .A(n15580), .ZN(n15584) );
  OR2_X1 U16636 ( .A1(n15584), .A2(n15583), .ZN(n15585) );
  OAI211_X1 U16637 ( .C1(n15587), .C2(n15671), .A(n15586), .B(n15585), .ZN(
        P3_U3188) );
  AOI21_X1 U16638 ( .B1(n15590), .B2(n15589), .A(n15588), .ZN(n15608) );
  INV_X1 U16639 ( .A(n15591), .ZN(n15592) );
  OAI21_X1 U16640 ( .B1(n15593), .B2(n15232), .A(n15592), .ZN(n15600) );
  INV_X1 U16641 ( .A(n15594), .ZN(n15595) );
  NAND3_X1 U16642 ( .A1(n15597), .A2(n15596), .A3(n15595), .ZN(n15598) );
  AOI21_X1 U16643 ( .B1(n15615), .B2(n15598), .A(n15659), .ZN(n15599) );
  AOI211_X1 U16644 ( .C1(n15602), .C2(n15601), .A(n15600), .B(n15599), .ZN(
        n15607) );
  XNOR2_X1 U16645 ( .A(n15604), .B(n15603), .ZN(n15605) );
  NAND2_X1 U16646 ( .A1(n15605), .A2(n15667), .ZN(n15606) );
  OAI211_X1 U16647 ( .C1(n15608), .C2(n15671), .A(n15607), .B(n15606), .ZN(
        P3_U3189) );
  AOI21_X1 U16648 ( .B1(n7360), .B2(n15610), .A(n15609), .ZN(n15627) );
  INV_X1 U16649 ( .A(n15611), .ZN(n15612) );
  NOR2_X1 U16650 ( .A1(n15613), .A2(n15612), .ZN(n15616) );
  INV_X1 U16651 ( .A(n15635), .ZN(n15614) );
  AOI21_X1 U16652 ( .B1(n15616), .B2(n15615), .A(n15614), .ZN(n15618) );
  OAI22_X1 U16653 ( .A1(n15618), .A2(n15659), .B1(n15617), .B2(n15657), .ZN(
        n15619) );
  AOI211_X1 U16654 ( .C1(P3_ADDR_REG_8__SCAN_IN), .C2(n15663), .A(n15620), .B(
        n15619), .ZN(n15626) );
  OAI21_X1 U16655 ( .B1(n15623), .B2(n15622), .A(n15621), .ZN(n15624) );
  NAND2_X1 U16656 ( .A1(n15624), .A2(n15667), .ZN(n15625) );
  OAI211_X1 U16657 ( .C1(n15627), .C2(n15671), .A(n15626), .B(n15625), .ZN(
        P3_U3190) );
  AOI21_X1 U16658 ( .B1(n15630), .B2(n15629), .A(n15628), .ZN(n15646) );
  INV_X1 U16659 ( .A(n15631), .ZN(n15632) );
  NOR2_X1 U16660 ( .A1(n15633), .A2(n15632), .ZN(n15636) );
  INV_X1 U16661 ( .A(n15655), .ZN(n15634) );
  AOI21_X1 U16662 ( .B1(n15636), .B2(n15635), .A(n15634), .ZN(n15638) );
  OAI22_X1 U16663 ( .A1(n15638), .A2(n15659), .B1(n15637), .B2(n15657), .ZN(
        n15639) );
  AOI211_X1 U16664 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15663), .A(n15640), .B(
        n15639), .ZN(n15645) );
  OAI21_X1 U16665 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15642), .A(n15641), .ZN(
        n15643) );
  NAND2_X1 U16666 ( .A1(n15643), .A2(n15667), .ZN(n15644) );
  OAI211_X1 U16667 ( .C1(n15646), .C2(n15671), .A(n15645), .B(n15644), .ZN(
        P3_U3191) );
  AOI21_X1 U16668 ( .B1(n15649), .B2(n15648), .A(n15647), .ZN(n15672) );
  INV_X1 U16669 ( .A(n15650), .ZN(n15651) );
  NOR2_X1 U16670 ( .A1(n15652), .A2(n15651), .ZN(n15656) );
  INV_X1 U16671 ( .A(n15653), .ZN(n15654) );
  AOI21_X1 U16672 ( .B1(n15656), .B2(n15655), .A(n15654), .ZN(n15660) );
  OAI22_X1 U16673 ( .A1(n15660), .A2(n15659), .B1(n15658), .B2(n15657), .ZN(
        n15661) );
  AOI211_X1 U16674 ( .C1(P3_ADDR_REG_10__SCAN_IN), .C2(n15663), .A(n15662), 
        .B(n15661), .ZN(n15670) );
  OAI21_X1 U16675 ( .B1(n15666), .B2(n15665), .A(n15664), .ZN(n15668) );
  NAND2_X1 U16676 ( .A1(n15668), .A2(n15667), .ZN(n15669) );
  OAI211_X1 U16677 ( .C1(n15672), .C2(n15671), .A(n15670), .B(n15669), .ZN(
        P3_U3192) );
  INV_X1 U16678 ( .A(P1_RD_REG_SCAN_IN), .ZN(n15674) );
  OAI221_X1 U16679 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(
        n15675), .C2(n15674), .A(n15673), .ZN(U29) );
  INV_X1 U16680 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15676) );
  AOI22_X1 U16681 ( .A1(n15961), .A2(n15677), .B1(n15676), .B2(n16023), .ZN(
        P1_U3459) );
  AOI22_X1 U16682 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(n15020), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n15678), .ZN(n15686) );
  AOI21_X1 U16683 ( .B1(n15681), .B2(n15680), .A(n15679), .ZN(n15682) );
  AOI21_X1 U16684 ( .B1(n15684), .B2(n15683), .A(n15682), .ZN(n15685) );
  OAI211_X1 U16685 ( .C1(n15020), .C2(n15687), .A(n15686), .B(n15685), .ZN(
        P1_U3293) );
  OAI211_X1 U16686 ( .C1(n15689), .C2(n15807), .A(n7201), .B(n15688), .ZN(
        n15690) );
  INV_X1 U16687 ( .A(n15690), .ZN(n15693) );
  AOI22_X1 U16688 ( .A1(n15970), .A2(n15693), .B1(n15691), .B2(n14355), .ZN(
        P2_U3499) );
  INV_X1 U16689 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15692) );
  AOI22_X1 U16690 ( .A1(n15974), .A2(n15693), .B1(n15692), .B2(n15971), .ZN(
        P2_U3430) );
  INV_X1 U16691 ( .A(n15694), .ZN(n15701) );
  INV_X1 U16692 ( .A(n15695), .ZN(n15729) );
  OAI22_X1 U16693 ( .A1(n15697), .A2(n15729), .B1(n15696), .B2(n15727), .ZN(
        n15700) );
  INV_X1 U16694 ( .A(n15698), .ZN(n15699) );
  AOI211_X1 U16695 ( .C1(n15702), .C2(n15701), .A(n15700), .B(n15699), .ZN(
        n15703) );
  AOI22_X1 U16696 ( .A1(n13670), .A2(n10251), .B1(n15703), .B2(n15735), .ZN(
        P3_U3232) );
  OAI22_X1 U16697 ( .A1(n15704), .A2(n16009), .B1(n9699), .B2(n15954), .ZN(
        n15706) );
  AOI211_X1 U16698 ( .C1(n15881), .C2(n15707), .A(n15706), .B(n15705), .ZN(
        n15709) );
  INV_X1 U16699 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15708) );
  AOI22_X1 U16700 ( .A1(n15922), .A2(n15709), .B1(n15708), .B2(n16021), .ZN(
        P1_U3529) );
  AOI22_X1 U16701 ( .A1(n15961), .A2(n15709), .B1(n8938), .B2(n16023), .ZN(
        P1_U3462) );
  INV_X1 U16702 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15710) );
  AOI22_X1 U16703 ( .A1(n15974), .A2(n15711), .B1(n15710), .B2(n15971), .ZN(
        P2_U3433) );
  OAI21_X1 U16704 ( .B1(n15713), .B2(n15715), .A(n15712), .ZN(n15733) );
  NOR2_X1 U16705 ( .A1(n15730), .A2(n15935), .ZN(n15724) );
  NAND3_X1 U16706 ( .A1(n15716), .A2(n15715), .A3(n15714), .ZN(n15717) );
  AND2_X1 U16707 ( .A1(n11056), .A2(n15717), .ZN(n15718) );
  OAI222_X1 U16708 ( .A1(n15723), .A2(n15722), .B1(n15721), .B2(n15720), .C1(
        n15719), .C2(n15718), .ZN(n15731) );
  AOI211_X1 U16709 ( .C1(n15912), .C2(n15733), .A(n15724), .B(n15731), .ZN(
        n15726) );
  AOI22_X1 U16710 ( .A1(n15940), .A2(n15726), .B1(n10305), .B2(n15939), .ZN(
        P3_U3461) );
  INV_X1 U16711 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15725) );
  AOI22_X1 U16712 ( .A1(n15944), .A2(n15726), .B1(n15725), .B2(n15941), .ZN(
        P3_U3396) );
  OAI22_X1 U16713 ( .A1(n15730), .A2(n15729), .B1(n15728), .B2(n15727), .ZN(
        n15732) );
  AOI211_X1 U16714 ( .C1(n15734), .C2(n15733), .A(n15732), .B(n15731), .ZN(
        n15736) );
  AOI22_X1 U16715 ( .A1(n13670), .A2(n15737), .B1(n15736), .B2(n15735), .ZN(
        P3_U3231) );
  INV_X1 U16716 ( .A(n15738), .ZN(n15743) );
  OAI22_X1 U16717 ( .A1(n15740), .A2(n16009), .B1(n15739), .B2(n15954), .ZN(
        n15742) );
  AOI211_X1 U16718 ( .C1(n15881), .C2(n15743), .A(n15742), .B(n15741), .ZN(
        n15745) );
  INV_X1 U16719 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n15744) );
  AOI22_X1 U16720 ( .A1(n15922), .A2(n15745), .B1(n15744), .B2(n16021), .ZN(
        P1_U3530) );
  AOI22_X1 U16721 ( .A1(n15961), .A2(n15745), .B1(n8889), .B2(n16023), .ZN(
        P1_U3465) );
  INV_X1 U16722 ( .A(n15746), .ZN(n15752) );
  NOR2_X1 U16723 ( .A1(n15746), .A2(n15778), .ZN(n15751) );
  OAI211_X1 U16724 ( .C1(n15749), .C2(n15963), .A(n15748), .B(n15747), .ZN(
        n15750) );
  AOI211_X1 U16725 ( .C1(n15950), .C2(n15752), .A(n15751), .B(n15750), .ZN(
        n15755) );
  INV_X1 U16726 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n15753) );
  AOI22_X1 U16727 ( .A1(n15970), .A2(n15755), .B1(n15753), .B2(n14355), .ZN(
        P2_U3501) );
  INV_X1 U16728 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15754) );
  AOI22_X1 U16729 ( .A1(n15974), .A2(n15755), .B1(n15754), .B2(n15971), .ZN(
        P2_U3436) );
  OAI22_X1 U16730 ( .A1(n15757), .A2(n16009), .B1(n15756), .B2(n15954), .ZN(
        n15759) );
  AOI211_X1 U16731 ( .C1(n15760), .C2(n16019), .A(n15759), .B(n15758), .ZN(
        n15761) );
  AOI22_X1 U16732 ( .A1(n15922), .A2(n15761), .B1(n9941), .B2(n16021), .ZN(
        P1_U3531) );
  AOI22_X1 U16733 ( .A1(n15961), .A2(n15761), .B1(n8966), .B2(n16023), .ZN(
        P1_U3468) );
  INV_X1 U16734 ( .A(n15762), .ZN(n15763) );
  OAI21_X1 U16735 ( .B1(n15764), .B2(n15963), .A(n15763), .ZN(n15767) );
  INV_X1 U16736 ( .A(n15765), .ZN(n15766) );
  AOI211_X1 U16737 ( .C1(n15950), .C2(n15768), .A(n15767), .B(n15766), .ZN(
        n15771) );
  INV_X1 U16738 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n15769) );
  AOI22_X1 U16739 ( .A1(n15970), .A2(n15771), .B1(n15769), .B2(n14355), .ZN(
        P2_U3502) );
  INV_X1 U16740 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15770) );
  AOI22_X1 U16741 ( .A1(n15974), .A2(n15771), .B1(n15770), .B2(n15971), .ZN(
        P2_U3439) );
  AOI22_X1 U16742 ( .A1(n15773), .A2(n15931), .B1(n15772), .B2(n15891), .ZN(
        n15774) );
  AND2_X1 U16743 ( .A1(n15775), .A2(n15774), .ZN(n15777) );
  AOI22_X1 U16744 ( .A1(n15940), .A2(n15777), .B1(n11411), .B2(n15939), .ZN(
        P3_U3463) );
  INV_X1 U16745 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15776) );
  AOI22_X1 U16746 ( .A1(n15944), .A2(n15777), .B1(n15776), .B2(n15941), .ZN(
        P3_U3402) );
  NOR2_X1 U16747 ( .A1(n15779), .A2(n15778), .ZN(n15784) );
  OAI211_X1 U16748 ( .C1(n15782), .C2(n15963), .A(n15781), .B(n15780), .ZN(
        n15783) );
  AOI211_X1 U16749 ( .C1(n15785), .C2(n15950), .A(n15784), .B(n15783), .ZN(
        n15788) );
  INV_X1 U16750 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n15786) );
  AOI22_X1 U16751 ( .A1(n15970), .A2(n15788), .B1(n15786), .B2(n14355), .ZN(
        P2_U3503) );
  INV_X1 U16752 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15787) );
  AOI22_X1 U16753 ( .A1(n15974), .A2(n15788), .B1(n15787), .B2(n15971), .ZN(
        P2_U3442) );
  NOR2_X1 U16754 ( .A1(n15789), .A2(n15935), .ZN(n15791) );
  AOI211_X1 U16755 ( .C1(n15912), .C2(n15792), .A(n15791), .B(n15790), .ZN(
        n15794) );
  AOI22_X1 U16756 ( .A1(n15940), .A2(n15794), .B1(n11418), .B2(n15939), .ZN(
        P3_U3464) );
  INV_X1 U16757 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15793) );
  AOI22_X1 U16758 ( .A1(n15944), .A2(n15794), .B1(n15793), .B2(n15941), .ZN(
        P3_U3405) );
  AOI22_X1 U16759 ( .A1(n15797), .A2(n15796), .B1(n16014), .B2(n15795), .ZN(
        n15798) );
  OAI21_X1 U16760 ( .B1(n15800), .B2(n15799), .A(n15798), .ZN(n15801) );
  NOR2_X1 U16761 ( .A1(n15802), .A2(n15801), .ZN(n15803) );
  AOI22_X1 U16762 ( .A1(n15922), .A2(n15803), .B1(n9943), .B2(n16021), .ZN(
        P1_U3533) );
  AOI22_X1 U16763 ( .A1(n15961), .A2(n15803), .B1(n9033), .B2(n16023), .ZN(
        P1_U3474) );
  INV_X1 U16764 ( .A(n15808), .ZN(n15811) );
  NAND2_X1 U16765 ( .A1(n15804), .A2(n15845), .ZN(n15805) );
  OAI211_X1 U16766 ( .C1(n15808), .C2(n15807), .A(n15806), .B(n15805), .ZN(
        n15810) );
  AOI211_X1 U16767 ( .C1(n15812), .C2(n15811), .A(n15810), .B(n15809), .ZN(
        n15814) );
  AOI22_X1 U16768 ( .A1(n15970), .A2(n15814), .B1(n10185), .B2(n14355), .ZN(
        P2_U3504) );
  INV_X1 U16769 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15813) );
  AOI22_X1 U16770 ( .A1(n15974), .A2(n15814), .B1(n15813), .B2(n15971), .ZN(
        P2_U3445) );
  AOI222_X1 U16771 ( .A1(n15819), .A2(n15818), .B1(P2_REG2_REG_6__SCAN_IN), 
        .B2(n15817), .C1(n15816), .C2(n15815), .ZN(n15827) );
  INV_X1 U16772 ( .A(n15820), .ZN(n15825) );
  INV_X1 U16773 ( .A(n15821), .ZN(n15822) );
  AOI22_X1 U16774 ( .A1(n15825), .A2(n15824), .B1(n15823), .B2(n15822), .ZN(
        n15826) );
  OAI211_X1 U16775 ( .C1(n15829), .C2(n15828), .A(n15827), .B(n15826), .ZN(
        P2_U3259) );
  NOR2_X1 U16776 ( .A1(n15830), .A2(n15935), .ZN(n15832) );
  AOI211_X1 U16777 ( .C1(n15931), .C2(n15833), .A(n15832), .B(n15831), .ZN(
        n15835) );
  AOI22_X1 U16778 ( .A1(n15940), .A2(n15835), .B1(n15603), .B2(n15939), .ZN(
        P3_U3466) );
  INV_X1 U16779 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15834) );
  AOI22_X1 U16780 ( .A1(n15944), .A2(n15835), .B1(n15834), .B2(n15941), .ZN(
        P3_U3411) );
  INV_X1 U16781 ( .A(n15836), .ZN(n15837) );
  OAI22_X1 U16782 ( .A1(n15838), .A2(n16009), .B1(n15837), .B2(n15954), .ZN(
        n15840) );
  AOI211_X1 U16783 ( .C1(n15881), .C2(n15841), .A(n15840), .B(n15839), .ZN(
        n15842) );
  AOI22_X1 U16784 ( .A1(n15922), .A2(n15842), .B1(n9945), .B2(n16021), .ZN(
        P1_U3535) );
  AOI22_X1 U16785 ( .A1(n15961), .A2(n15842), .B1(n9073), .B2(n16023), .ZN(
        P1_U3480) );
  AOI21_X1 U16786 ( .B1(n15845), .B2(n15844), .A(n15843), .ZN(n15846) );
  OAI21_X1 U16787 ( .B1(n15848), .B2(n15847), .A(n15846), .ZN(n15850) );
  NOR2_X1 U16788 ( .A1(n15850), .A2(n15849), .ZN(n15853) );
  INV_X1 U16789 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n15851) );
  AOI22_X1 U16790 ( .A1(n15970), .A2(n15853), .B1(n15851), .B2(n14355), .ZN(
        P2_U3506) );
  INV_X1 U16791 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15852) );
  AOI22_X1 U16792 ( .A1(n15974), .A2(n15853), .B1(n15852), .B2(n15971), .ZN(
        P2_U3451) );
  AOI22_X1 U16793 ( .A1(n15855), .A2(n15931), .B1(n15891), .B2(n15854), .ZN(
        n15856) );
  AND2_X1 U16794 ( .A1(n15857), .A2(n15856), .ZN(n15859) );
  AOI22_X1 U16795 ( .A1(n15940), .A2(n15859), .B1(n11432), .B2(n15939), .ZN(
        P3_U3467) );
  INV_X1 U16796 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15858) );
  AOI22_X1 U16797 ( .A1(n15944), .A2(n15859), .B1(n15858), .B2(n15941), .ZN(
        P3_U3414) );
  NAND3_X1 U16798 ( .A1(n15861), .A2(n15860), .A3(n15968), .ZN(n15863) );
  OAI211_X1 U16799 ( .C1(n15864), .C2(n15963), .A(n15863), .B(n15862), .ZN(
        n15865) );
  NOR2_X1 U16800 ( .A1(n15866), .A2(n15865), .ZN(n15868) );
  AOI22_X1 U16801 ( .A1(n15970), .A2(n15868), .B1(n10186), .B2(n14355), .ZN(
        P2_U3507) );
  INV_X1 U16802 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15867) );
  AOI22_X1 U16803 ( .A1(n15974), .A2(n15868), .B1(n15867), .B2(n15971), .ZN(
        P2_U3454) );
  OAI21_X1 U16804 ( .B1(n15870), .B2(n15935), .A(n15869), .ZN(n15871) );
  AOI21_X1 U16805 ( .B1(n15872), .B2(n15912), .A(n15871), .ZN(n15874) );
  AOI22_X1 U16806 ( .A1(n15940), .A2(n15874), .B1(n11437), .B2(n15939), .ZN(
        P3_U3468) );
  INV_X1 U16807 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15873) );
  AOI22_X1 U16808 ( .A1(n15944), .A2(n15874), .B1(n15873), .B2(n15941), .ZN(
        P3_U3417) );
  INV_X1 U16809 ( .A(n15875), .ZN(n15876) );
  OAI21_X1 U16810 ( .B1(n15877), .B2(n15954), .A(n15876), .ZN(n15879) );
  AOI211_X1 U16811 ( .C1(n15881), .C2(n15880), .A(n15879), .B(n15878), .ZN(
        n15882) );
  AOI22_X1 U16812 ( .A1(n15922), .A2(n15882), .B1(n10020), .B2(n16021), .ZN(
        P1_U3537) );
  AOI22_X1 U16813 ( .A1(n15961), .A2(n15882), .B1(n9117), .B2(n16023), .ZN(
        P1_U3486) );
  INV_X1 U16814 ( .A(n15883), .ZN(n15888) );
  OAI21_X1 U16815 ( .B1(n15885), .B2(n15963), .A(n15884), .ZN(n15887) );
  AOI211_X1 U16816 ( .C1(n15950), .C2(n15888), .A(n15887), .B(n15886), .ZN(
        n15890) );
  AOI22_X1 U16817 ( .A1(n15970), .A2(n15890), .B1(n10319), .B2(n14355), .ZN(
        P2_U3508) );
  INV_X1 U16818 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n15889) );
  AOI22_X1 U16819 ( .A1(n15974), .A2(n15890), .B1(n15889), .B2(n15971), .ZN(
        P2_U3457) );
  NAND2_X1 U16820 ( .A1(n15892), .A2(n15891), .ZN(n15893) );
  OAI211_X1 U16821 ( .C1(n15896), .C2(n15895), .A(n15894), .B(n15893), .ZN(
        n15897) );
  AOI21_X1 U16822 ( .B1(n15937), .B2(n15898), .A(n15897), .ZN(n15900) );
  AOI22_X1 U16823 ( .A1(n15940), .A2(n15900), .B1(n11443), .B2(n15939), .ZN(
        P3_U3469) );
  INV_X1 U16824 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15899) );
  AOI22_X1 U16825 ( .A1(n15944), .A2(n15900), .B1(n15899), .B2(n15941), .ZN(
        P3_U3420) );
  INV_X1 U16826 ( .A(n15901), .ZN(n15906) );
  OAI21_X1 U16827 ( .B1(n15903), .B2(n15963), .A(n15902), .ZN(n15905) );
  AOI211_X1 U16828 ( .C1(n15950), .C2(n15906), .A(n15905), .B(n15904), .ZN(
        n15908) );
  AOI22_X1 U16829 ( .A1(n15970), .A2(n15908), .B1(n10673), .B2(n14355), .ZN(
        P2_U3509) );
  INV_X1 U16830 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15907) );
  AOI22_X1 U16831 ( .A1(n15974), .A2(n15908), .B1(n15907), .B2(n15971), .ZN(
        P2_U3460) );
  OAI21_X1 U16832 ( .B1(n15910), .B2(n15935), .A(n15909), .ZN(n15911) );
  AOI21_X1 U16833 ( .B1(n15913), .B2(n15912), .A(n15911), .ZN(n15916) );
  INV_X1 U16834 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n15914) );
  AOI22_X1 U16835 ( .A1(n15940), .A2(n15916), .B1(n15914), .B2(n15939), .ZN(
        P3_U3470) );
  INV_X1 U16836 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n15915) );
  AOI22_X1 U16837 ( .A1(n15944), .A2(n15916), .B1(n15915), .B2(n15941), .ZN(
        P3_U3423) );
  OAI22_X1 U16838 ( .A1(n15918), .A2(n16009), .B1(n7721), .B2(n15954), .ZN(
        n15919) );
  AOI211_X1 U16839 ( .C1(n15921), .C2(n16019), .A(n15920), .B(n15919), .ZN(
        n15923) );
  AOI22_X1 U16840 ( .A1(n15922), .A2(n15923), .B1(n10096), .B2(n16021), .ZN(
        P1_U3539) );
  AOI22_X1 U16841 ( .A1(n15961), .A2(n15923), .B1(n9159), .B2(n16023), .ZN(
        P1_U3492) );
  OAI21_X1 U16842 ( .B1(n15925), .B2(n15963), .A(n15924), .ZN(n15927) );
  AOI211_X1 U16843 ( .C1(n15950), .C2(n15928), .A(n15927), .B(n15926), .ZN(
        n15930) );
  AOI22_X1 U16844 ( .A1(n15970), .A2(n15930), .B1(n10904), .B2(n14355), .ZN(
        P2_U3510) );
  INV_X1 U16845 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n15929) );
  AOI22_X1 U16846 ( .A1(n15974), .A2(n15930), .B1(n15929), .B2(n15971), .ZN(
        P2_U3463) );
  NAND2_X1 U16847 ( .A1(n15938), .A2(n15931), .ZN(n15932) );
  OAI211_X1 U16848 ( .C1(n15935), .C2(n15934), .A(n15933), .B(n15932), .ZN(
        n15936) );
  AOI21_X1 U16849 ( .B1(n15938), .B2(n15937), .A(n15936), .ZN(n15943) );
  AOI22_X1 U16850 ( .A1(n15940), .A2(n15943), .B1(n11677), .B2(n15939), .ZN(
        P3_U3471) );
  INV_X1 U16851 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n15942) );
  AOI22_X1 U16852 ( .A1(n15944), .A2(n15943), .B1(n15942), .B2(n15941), .ZN(
        P3_U3426) );
  OAI21_X1 U16853 ( .B1(n15946), .B2(n15963), .A(n15945), .ZN(n15948) );
  AOI211_X1 U16854 ( .C1(n15950), .C2(n15949), .A(n15948), .B(n15947), .ZN(
        n15952) );
  AOI22_X1 U16855 ( .A1(n15970), .A2(n15952), .B1(n11356), .B2(n14355), .ZN(
        P2_U3511) );
  INV_X1 U16856 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n15951) );
  AOI22_X1 U16857 ( .A1(n15974), .A2(n15952), .B1(n15951), .B2(n15971), .ZN(
        P2_U3466) );
  INV_X1 U16858 ( .A(n15953), .ZN(n15959) );
  OAI22_X1 U16859 ( .A1(n15956), .A2(n16009), .B1(n15955), .B2(n15954), .ZN(
        n15957) );
  AOI211_X1 U16860 ( .C1(n15959), .C2(n16019), .A(n15958), .B(n15957), .ZN(
        n15960) );
  AOI22_X1 U16861 ( .A1(n15922), .A2(n15960), .B1(n10631), .B2(n16021), .ZN(
        P1_U3541) );
  AOI22_X1 U16862 ( .A1(n15961), .A2(n15960), .B1(n9219), .B2(n16023), .ZN(
        P1_U3498) );
  OAI21_X1 U16863 ( .B1(n15964), .B2(n15963), .A(n15962), .ZN(n15966) );
  AOI211_X1 U16864 ( .C1(n15968), .C2(n15967), .A(n15966), .B(n15965), .ZN(
        n15973) );
  AOI22_X1 U16865 ( .A1(n15970), .A2(n15973), .B1(n15969), .B2(n14355), .ZN(
        P2_U3513) );
  INV_X1 U16866 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n15972) );
  AOI22_X1 U16867 ( .A1(n15974), .A2(n15973), .B1(n15972), .B2(n15971), .ZN(
        P2_U3472) );
  OAI21_X1 U16868 ( .B1(n15977), .B2(n15976), .A(n15975), .ZN(n15981) );
  AOI22_X1 U16869 ( .A1(n16031), .A2(n16028), .B1(n16029), .B2(n15978), .ZN(
        n15979) );
  OAI21_X1 U16870 ( .B1(n7715), .B2(n16033), .A(n15979), .ZN(n15980) );
  AOI21_X1 U16871 ( .B1(n15981), .B2(n16036), .A(n15980), .ZN(n15983) );
  OAI211_X1 U16872 ( .C1(n16041), .C2(n15984), .A(n15983), .B(n15982), .ZN(
        P1_U3241) );
  NAND3_X1 U16873 ( .A1(n15987), .A2(n15986), .A3(n15985), .ZN(n15991) );
  AOI21_X1 U16874 ( .B1(n15989), .B2(n16014), .A(n15988), .ZN(n15990) );
  OAI211_X1 U16875 ( .C1(n16009), .C2(n15992), .A(n15991), .B(n15990), .ZN(
        n15993) );
  AOI21_X1 U16876 ( .B1(n15994), .B2(n16019), .A(n15993), .ZN(n15996) );
  AOI22_X1 U16877 ( .A1(n15922), .A2(n15996), .B1(n15995), .B2(n16021), .ZN(
        P1_U3543) );
  AOI22_X1 U16878 ( .A1(n15961), .A2(n15996), .B1(n9252), .B2(n16023), .ZN(
        P1_U3504) );
  XNOR2_X1 U16879 ( .A(n15998), .B(n15999), .ZN(n16005) );
  AOI22_X1 U16880 ( .A1(n16031), .A2(n16001), .B1(n16029), .B2(n16000), .ZN(
        n16002) );
  OAI21_X1 U16881 ( .B1(n16003), .B2(n16033), .A(n16002), .ZN(n16004) );
  AOI21_X1 U16882 ( .B1(n16005), .B2(n16036), .A(n16004), .ZN(n16007) );
  OAI211_X1 U16883 ( .C1(n16041), .C2(n16008), .A(n16007), .B(n16006), .ZN(
        P1_U3226) );
  NOR2_X1 U16884 ( .A1(n16010), .A2(n16009), .ZN(n16011) );
  AOI211_X1 U16885 ( .C1(n16014), .C2(n16013), .A(n16012), .B(n16011), .ZN(
        n16015) );
  OAI21_X1 U16886 ( .B1(n16017), .B2(n16016), .A(n16015), .ZN(n16018) );
  AOI21_X1 U16887 ( .B1(n16020), .B2(n16019), .A(n16018), .ZN(n16024) );
  AOI22_X1 U16888 ( .A1(n15922), .A2(n16024), .B1(n16022), .B2(n16021), .ZN(
        P1_U3544) );
  AOI22_X1 U16889 ( .A1(n15961), .A2(n16024), .B1(n9278), .B2(n16023), .ZN(
        P1_U3507) );
  XNOR2_X1 U16890 ( .A(n16025), .B(n16026), .ZN(n16037) );
  INV_X1 U16891 ( .A(n16027), .ZN(n16034) );
  AOI22_X1 U16892 ( .A1(n16031), .A2(n16030), .B1(n16029), .B2(n16028), .ZN(
        n16032) );
  OAI21_X1 U16893 ( .B1(n16034), .B2(n16033), .A(n16032), .ZN(n16035) );
  AOI21_X1 U16894 ( .B1(n16037), .B2(n16036), .A(n16035), .ZN(n16039) );
  OAI211_X1 U16895 ( .C1(n16041), .C2(n16040), .A(n16039), .B(n16038), .ZN(
        P1_U3228) );
  AOI21_X1 U16896 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16042) );
  OAI21_X1 U16897 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16042), 
        .ZN(U28) );
  CLKBUF_X1 U7297 ( .A(n9267), .Z(n9538) );
  AND2_X1 U7306 ( .A1(n14507), .A2(n7526), .ZN(n8259) );
  CLKBUF_X1 U7310 ( .A(n7250), .Z(n8759) );
  CLKBUF_X3 U7372 ( .A(n8521), .Z(n12552) );
  NAND2_X1 U7542 ( .A1(n13600), .A2(n13599), .ZN(n13602) );
  CLKBUF_X2 U7595 ( .A(n9031), .Z(n9544) );
  CLKBUF_X1 U8613 ( .A(n8959), .Z(n9891) );
  CLKBUF_X1 U8735 ( .A(n7642), .Z(n8885) );
  INV_X1 U9102 ( .A(n12848), .ZN(n12956) );
endmodule

