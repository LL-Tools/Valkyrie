

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620;

  INV_X4 U7530 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U7531 ( .A1(n12253), .A2(n12254), .ZN(n12463) );
  INV_X2 U7532 ( .A(n14827), .ZN(n14919) );
  INV_X1 U7533 ( .A(n14863), .ZN(n11755) );
  INV_X1 U7534 ( .A(n7458), .ZN(n7460) );
  INV_X2 U7535 ( .A(n9817), .ZN(n9770) );
  BUF_X2 U7536 ( .A(n9311), .Z(n7814) );
  NAND2_X1 U7537 ( .A1(n15761), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9212) );
  OR2_X1 U7538 ( .A1(n14148), .A2(n14147), .ZN(n14155) );
  INV_X1 U7539 ( .A(n14235), .ZN(n14256) );
  AND2_X1 U7540 ( .A1(n10949), .A2(n10948), .ZN(n11080) );
  INV_X1 U7541 ( .A(n12731), .ZN(n12728) );
  INV_X1 U7542 ( .A(n11208), .ZN(n14917) );
  INV_X1 U7543 ( .A(n7458), .ZN(n7459) );
  INV_X1 U7544 ( .A(n9814), .ZN(n11433) );
  XNOR2_X1 U7545 ( .A(n14763), .B(n14133), .ZN(n14307) );
  CLKBUF_X2 U7546 ( .A(n7490), .Z(n7437) );
  INV_X1 U7548 ( .A(n16396), .ZN(n9625) );
  AND2_X1 U7549 ( .A1(n12726), .A2(n12722), .ZN(n13104) );
  INV_X1 U7550 ( .A(n11026), .ZN(n7779) );
  BUF_X1 U7551 ( .A(n14218), .Z(n8851) );
  CLKBUF_X3 U7552 ( .A(n9147), .Z(n7431) );
  INV_X1 U7553 ( .A(n15213), .ZN(n15783) );
  OR2_X1 U7554 ( .A1(n14051), .A2(n14050), .ZN(n7429) );
  OAI21_X1 U7555 ( .B1(n14970), .B2(n14968), .A(n14966), .ZN(n15004) );
  AOI21_X2 U7556 ( .B1(n8231), .B2(n8233), .A(n7477), .ZN(n8229) );
  NAND2_X2 U7557 ( .A1(n14286), .A2(n14320), .ZN(n7685) );
  NAND2_X2 U7559 ( .A1(n12064), .A2(n15236), .ZN(n16422) );
  XNOR2_X2 U7560 ( .A(n7749), .B(n11831), .ZN(n11818) );
  NAND2_X2 U7561 ( .A1(n11663), .A2(n11662), .ZN(n7749) );
  NOR2_X2 U7562 ( .A1(n7453), .A2(n7452), .ZN(n9456) );
  OAI222_X1 U7563 ( .A1(n15780), .A2(n15768), .B1(P1_U3086), .B2(n15767), .C1(
        n15766), .C2(n15777), .ZN(P1_U3325) );
  BUF_X2 U7564 ( .A(n10269), .Z(n7430) );
  XNOR2_X2 U7565 ( .A(n8593), .B(SI_2_), .ZN(n8592) );
  OAI22_X1 U7566 ( .A1(n8334), .A2(n8331), .B1(n14070), .B2(n14069), .ZN(
        n14078) );
  XNOR2_X2 U7567 ( .A(n9755), .B(P3_IR_REG_30__SCAN_IN), .ZN(n9760) );
  XNOR2_X2 U7568 ( .A(n7698), .B(n8550), .ZN(n9149) );
  XNOR2_X2 U7569 ( .A(n9214), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9216) );
  NAND2_X2 U7570 ( .A1(n7444), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9214) );
  AOI21_X2 U7571 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(n16023), .A(n16022), .ZN(
        n16034) );
  INV_X4 U7572 ( .A(n8586), .ZN(n8612) );
  NAND2_X4 U7573 ( .A1(n8867), .A2(n8866), .ZN(n14763) );
  XNOR2_X1 U7574 ( .A(n9769), .B(n9768), .ZN(n7432) );
  INV_X8 U7575 ( .A(n10990), .ZN(n13036) );
  NOR2_X1 U7576 ( .A1(n15681), .A2(n8106), .ZN(n8105) );
  INV_X1 U7577 ( .A(n15260), .ZN(n7434) );
  OAI21_X1 U7578 ( .B1(n15630), .B2(n8286), .A(n8285), .ZN(n15593) );
  NAND2_X1 U7579 ( .A1(n9570), .A2(n9569), .ZN(n15664) );
  AND2_X1 U7580 ( .A1(n12305), .A2(n8168), .ZN(n12390) );
  CLKBUF_X2 U7581 ( .A(n14716), .Z(n7757) );
  OR2_X1 U7582 ( .A1(n10158), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n10171) );
  NAND2_X1 U7583 ( .A1(n8728), .A2(n8727), .ZN(n14073) );
  INV_X4 U7584 ( .A(n15211), .ZN(n15065) );
  INV_X1 U7585 ( .A(n15323), .ZN(n11466) );
  CLKBUF_X1 U7586 ( .A(n11576), .Z(n15327) );
  INV_X2 U7587 ( .A(n10884), .ZN(n7433) );
  INV_X1 U7588 ( .A(n15195), .ZN(n9254) );
  BUF_X2 U7589 ( .A(n9318), .Z(n15206) );
  NOR2_X1 U7590 ( .A1(n8158), .A2(n8156), .ZN(n9287) );
  AND2_X1 U7591 ( .A1(n9261), .A2(n8156), .ZN(n9318) );
  INV_X1 U7592 ( .A(n14006), .ZN(n11365) );
  CLKBUF_X2 U7593 ( .A(n8575), .Z(n9039) );
  NAND2_X2 U7594 ( .A1(n15772), .A2(n15885), .ZN(n9261) );
  INV_X2 U7595 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n13843) );
  AND2_X1 U7596 ( .A1(n9683), .A2(n9682), .ZN(n7777) );
  INV_X1 U7597 ( .A(n9680), .ZN(n12777) );
  AOI21_X1 U7598 ( .B1(n15466), .B2(n16536), .A(n15465), .ZN(n15666) );
  NAND2_X1 U7599 ( .A1(n15447), .A2(n9676), .ZN(n7447) );
  AOI21_X1 U7600 ( .B1(n13320), .B2(n16597), .A(n13319), .ZN(n13388) );
  AND2_X1 U7601 ( .A1(n8124), .A2(n12769), .ZN(n7776) );
  NAND2_X1 U7602 ( .A1(n15446), .A2(n15445), .ZN(n15447) );
  OR2_X1 U7603 ( .A1(n14738), .A2(n16561), .ZN(n7806) );
  NOR2_X1 U7604 ( .A1(n15450), .A2(n15256), .ZN(n9675) );
  OAI21_X1 U7605 ( .B1(n8139), .B2(n7790), .A(n12578), .ZN(n12579) );
  AOI21_X1 U7606 ( .B1(n14950), .B2(n14951), .A(n8511), .ZN(n15014) );
  OR2_X1 U7607 ( .A1(n12734), .A2(n12733), .ZN(n8123) );
  NAND2_X1 U7608 ( .A1(n15520), .A2(n7451), .ZN(n15497) );
  AND2_X1 U7609 ( .A1(n15520), .A2(n9671), .ZN(n15499) );
  NAND2_X1 U7610 ( .A1(n8292), .A2(n8291), .ZN(n15520) );
  AOI21_X1 U7611 ( .B1(n8049), .B2(n16195), .A(n8048), .ZN(n8047) );
  NAND2_X1 U7612 ( .A1(n15525), .A2(n15528), .ZN(n8292) );
  NAND2_X1 U7613 ( .A1(n15542), .A2(n9669), .ZN(n15525) );
  AOI22_X1 U7614 ( .A1(n9738), .A2(n14312), .B1(n14193), .B2(n14341), .ZN(
        n9106) );
  NOR2_X1 U7615 ( .A1(n13062), .A2(n13061), .ZN(n13073) );
  NAND2_X1 U7616 ( .A1(n7442), .A2(n8277), .ZN(n15542) );
  NAND2_X1 U7617 ( .A1(n13885), .A2(n8519), .ZN(n13943) );
  NAND2_X1 U7618 ( .A1(n7441), .A2(n7439), .ZN(n7442) );
  NAND2_X1 U7619 ( .A1(n7441), .A2(n9664), .ZN(n15571) );
  OAI21_X1 U7620 ( .B1(n14489), .B2(n14313), .A(n7691), .ZN(n14465) );
  NOR2_X1 U7621 ( .A1(n16257), .A2(n13060), .ZN(n13062) );
  NAND2_X1 U7622 ( .A1(n7809), .A2(n8216), .ZN(n14489) );
  NAND2_X1 U7623 ( .A1(n9139), .A2(n9138), .ZN(n14506) );
  NAND2_X1 U7624 ( .A1(n9663), .A2(n8517), .ZN(n7441) );
  OR2_X1 U7625 ( .A1(n15482), .A2(n15664), .ZN(n15470) );
  NAND2_X1 U7626 ( .A1(n7658), .A2(n9136), .ZN(n14521) );
  OAI22_X1 U7627 ( .A1(n12500), .A2(n15249), .B1(n15314), .B2(n15732), .ZN(
        n15630) );
  OAI21_X1 U7628 ( .B1(n14566), .B2(n8213), .A(n8211), .ZN(n7658) );
  NAND2_X1 U7629 ( .A1(n12490), .A2(n9660), .ZN(n12500) );
  NAND2_X1 U7630 ( .A1(n14562), .A2(n8220), .ZN(n14680) );
  NAND2_X1 U7631 ( .A1(n8197), .A2(n8195), .ZN(n14583) );
  NAND2_X1 U7632 ( .A1(n12288), .A2(n7445), .ZN(n12490) );
  AND2_X1 U7633 ( .A1(n15498), .A2(n9671), .ZN(n7451) );
  AND2_X1 U7634 ( .A1(n12288), .A2(n9659), .ZN(n7446) );
  OR2_X1 U7635 ( .A1(n12514), .A2(n8200), .ZN(n8197) );
  AND2_X1 U7636 ( .A1(n8212), .A2(n14541), .ZN(n8211) );
  NAND2_X1 U7637 ( .A1(n16214), .A2(n13019), .ZN(n13021) );
  NAND2_X1 U7638 ( .A1(n9557), .A2(n9556), .ZN(n15681) );
  NAND2_X1 U7639 ( .A1(n12463), .A2(n7521), .ZN(n14943) );
  NOR2_X1 U7640 ( .A1(n8279), .A2(n7440), .ZN(n7439) );
  NAND2_X1 U7641 ( .A1(n12367), .A2(n9125), .ZN(n12430) );
  NAND2_X1 U7642 ( .A1(n14610), .A2(n14609), .ZN(n14608) );
  NAND2_X1 U7643 ( .A1(n12001), .A2(n9655), .ZN(n11955) );
  AOI21_X1 U7644 ( .B1(n9124), .B2(n7473), .A(n7532), .ZN(n12368) );
  OR2_X1 U7645 ( .A1(n14066), .A2(n14065), .ZN(n8334) );
  INV_X1 U7646 ( .A(n9664), .ZN(n7440) );
  AND2_X1 U7647 ( .A1(n12491), .A2(n9659), .ZN(n7445) );
  XNOR2_X1 U7648 ( .A(n13015), .B(n13047), .ZN(n16160) );
  NAND2_X1 U7649 ( .A1(n7784), .A2(n7783), .ZN(n11879) );
  NAND2_X1 U7650 ( .A1(n9488), .A2(n9487), .ZN(n15715) );
  NAND2_X1 U7651 ( .A1(n9474), .A2(n9473), .ZN(n15725) );
  OAI21_X1 U7652 ( .B1(n11382), .B2(n14294), .A(n9118), .ZN(n11608) );
  NAND2_X1 U7653 ( .A1(n8850), .A2(n8849), .ZN(n14122) );
  XNOR2_X1 U7654 ( .A(n8432), .B(n7595), .ZN(n11263) );
  CLKBUF_X2 U7655 ( .A(n14101), .Z(n7765) );
  NAND2_X1 U7656 ( .A1(n11867), .A2(n12744), .ZN(n11866) );
  NAND2_X1 U7657 ( .A1(n9398), .A2(n9397), .ZN(n16572) );
  NAND2_X1 U7658 ( .A1(n8775), .A2(n8774), .ZN(n14094) );
  NAND2_X1 U7659 ( .A1(n8784), .A2(n8514), .ZN(n8786) );
  INV_X2 U7660 ( .A(n16579), .ZN(n7435) );
  NAND2_X1 U7661 ( .A1(n8767), .A2(n8766), .ZN(n8784) );
  NAND2_X1 U7662 ( .A1(n8745), .A2(n8444), .ZN(n8767) );
  NAND2_X1 U7663 ( .A1(n10774), .A2(n9113), .ZN(n10355) );
  NAND2_X1 U7664 ( .A1(n9367), .A2(n9366), .ZN(n16531) );
  NAND2_X1 U7665 ( .A1(n8708), .A2(n8707), .ZN(n14629) );
  NAND2_X1 U7666 ( .A1(n9641), .A2(n9640), .ZN(n12106) );
  NAND2_X2 U7667 ( .A1(n11283), .A2(P1_STATE_REG_SCAN_IN), .ZN(n16619) );
  NOR2_X1 U7668 ( .A1(n15895), .A2(n15345), .ZN(n16294) );
  INV_X1 U7669 ( .A(n9648), .ZN(n7449) );
  INV_X1 U7670 ( .A(n11988), .ZN(n15234) );
  AND2_X1 U7671 ( .A1(n15041), .A2(n15044), .ZN(n11987) );
  AND2_X1 U7672 ( .A1(n12608), .A2(n12607), .ZN(n12740) );
  INV_X1 U7673 ( .A(n16425), .ZN(n15055) );
  XNOR2_X1 U7674 ( .A(n15325), .B(n16425), .ZN(n15236) );
  INV_X2 U7675 ( .A(n11080), .ZN(n12821) );
  NAND2_X1 U7676 ( .A1(n7747), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7769) );
  INV_X1 U7677 ( .A(n16465), .ZN(n7436) );
  NAND2_X1 U7678 ( .A1(n9295), .A2(n9294), .ZN(n16425) );
  NOR2_X1 U7679 ( .A1(n11126), .A2(n11125), .ZN(n11128) );
  NAND2_X1 U7680 ( .A1(n9269), .A2(n9268), .ZN(n15045) );
  OR2_X1 U7681 ( .A1(n8118), .A2(n8119), .ZN(n12997) );
  XNOR2_X1 U7682 ( .A(n15326), .B(n16396), .ZN(n15235) );
  AND2_X2 U7683 ( .A1(n11977), .A2(n15212), .ZN(n16473) );
  AND4_X1 U7684 ( .A1(n9299), .A2(n9298), .A3(n9297), .A4(n9296), .ZN(n15056)
         );
  AND4_X1 U7685 ( .A1(n9843), .A2(n9842), .A3(n9841), .A4(n9840), .ZN(n11926)
         );
  INV_X1 U7686 ( .A(n16374), .ZN(n7812) );
  AND4_X1 U7687 ( .A1(n9821), .A2(n9820), .A3(n9819), .A4(n9818), .ZN(n11738)
         );
  NAND4_X1 U7688 ( .A1(n9271), .A2(n9272), .A3(n9273), .A4(n9270), .ZN(n9639)
         );
  NAND2_X1 U7689 ( .A1(n8299), .A2(n9291), .ZN(n16396) );
  AOI21_X1 U7690 ( .B1(n8087), .B2(n11101), .A(n11030), .ZN(n11105) );
  XNOR2_X2 U7691 ( .A(n14366), .B(n11365), .ZN(n14287) );
  INV_X1 U7692 ( .A(n9287), .ZN(n7458) );
  NAND2_X1 U7693 ( .A1(n7684), .A2(n14424), .ZN(n11636) );
  NAND4_X1 U7694 ( .A1(n8567), .A2(n8565), .A3(n8566), .A4(n8568), .ZN(n14366)
         );
  OR2_X1 U7695 ( .A1(n9311), .A2(n15332), .ZN(n7456) );
  NAND2_X1 U7696 ( .A1(n8180), .A2(n8598), .ZN(n14027) );
  NAND2_X2 U7697 ( .A1(n7904), .A2(n9761), .ZN(n9814) );
  NAND2_X1 U7698 ( .A1(n15767), .A2(n15769), .ZN(n9282) );
  NAND2_X1 U7699 ( .A1(n9216), .A2(n15767), .ZN(n15195) );
  NAND2_X1 U7700 ( .A1(n7984), .A2(n7983), .ZN(n8624) );
  NAND2_X1 U7701 ( .A1(n9216), .A2(n9217), .ZN(n9311) );
  INV_X1 U7702 ( .A(n9477), .ZN(n7818) );
  INV_X1 U7703 ( .A(n13854), .ZN(n9761) );
  XNOR2_X1 U7704 ( .A(n9686), .B(P1_IR_REG_24__SCAN_IN), .ZN(n9704) );
  INV_X2 U7705 ( .A(n9860), .ZN(n10088) );
  OAI21_X1 U7706 ( .B1(n9709), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9685) );
  XNOR2_X1 U7708 ( .A(n9623), .B(n13801), .ZN(n15212) );
  XNOR2_X1 U7709 ( .A(n9769), .B(n9768), .ZN(n10270) );
  NAND2_X1 U7710 ( .A1(n9756), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9758) );
  NAND2_X1 U7711 ( .A1(n8535), .A2(n8534), .ZN(n14286) );
  NAND2_X1 U7712 ( .A1(n10488), .A2(n8156), .ZN(n8921) );
  NAND2_X1 U7713 ( .A1(n9202), .A2(n7557), .ZN(n7444) );
  OR2_X1 U7714 ( .A1(n9890), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9913) );
  XNOR2_X1 U7715 ( .A(n8538), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9147) );
  XNOR2_X1 U7716 ( .A(n8533), .B(P2_IR_REG_21__SCAN_IN), .ZN(n14320) );
  AND3_X1 U7717 ( .A1(n8494), .A2(n8076), .A3(n9861), .ZN(n9767) );
  OR2_X1 U7718 ( .A1(n9159), .A2(n14772), .ZN(n8537) );
  NAND2_X1 U7719 ( .A1(n9210), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9204) );
  INV_X1 U7720 ( .A(n9205), .ZN(n9202) );
  XNOR2_X1 U7721 ( .A(n8275), .B(SI_1_), .ZN(n8585) );
  NOR2_X1 U7722 ( .A1(n8077), .A2(n8151), .ZN(n8076) );
  NOR2_X1 U7723 ( .A1(n8536), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n9159) );
  XNOR2_X1 U7724 ( .A(n7660), .B(n8558), .ZN(n12791) );
  NAND2_X1 U7725 ( .A1(n8459), .A2(n7443), .ZN(n9205) );
  INV_X2 U7726 ( .A(n7626), .ZN(n14787) );
  AND2_X1 U7727 ( .A1(n7640), .A2(n9301), .ZN(n7443) );
  NAND2_X1 U7728 ( .A1(n7851), .A2(n7461), .ZN(n8077) );
  NAND2_X1 U7729 ( .A1(n8155), .A2(SI_0_), .ZN(n10420) );
  OAI21_X1 U7730 ( .B1(P1_ADDR_REG_1__SCAN_IN), .B2(n15940), .A(n15939), .ZN(
        n15949) );
  NAND2_X1 U7731 ( .A1(n8094), .A2(n8093), .ZN(n11026) );
  BUF_X4 U7732 ( .A(n10419), .Z(n8156) );
  NOR2_X1 U7733 ( .A1(n8495), .A2(P3_IR_REG_24__SCAN_IN), .ZN(n8494) );
  AND2_X1 U7734 ( .A1(n7642), .A2(n7641), .ZN(n7640) );
  NAND2_X2 U7735 ( .A1(n10419), .A2(P1_U3086), .ZN(n15780) );
  NAND2_X2 U7736 ( .A1(n8403), .A2(n8401), .ZN(n10419) );
  NAND4_X1 U7737 ( .A1(n15421), .A2(n10404), .A3(n8404), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n8403) );
  NAND4_X1 U7738 ( .A1(n13084), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(n8402), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n8401) );
  AND4_X1 U7739 ( .A1(n7653), .A2(n7652), .A3(n7651), .A4(n7650), .ZN(n8524)
         );
  AND2_X1 U7740 ( .A1(n8581), .A2(n8522), .ZN(n8596) );
  AND2_X1 U7741 ( .A1(n13770), .A2(n7890), .ZN(n7889) );
  INV_X1 U7742 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n13584) );
  NOR2_X1 U7743 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n9196) );
  NOR2_X1 U7744 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n9197) );
  NOR2_X1 U7745 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n9198) );
  INV_X1 U7746 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n13589) );
  INV_X1 U7747 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n13789) );
  INV_X1 U7748 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9211) );
  INV_X1 U7749 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9335) );
  INV_X4 U7750 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7751 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9884) );
  INV_X4 U7752 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7753 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9441) );
  NOR2_X1 U7754 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n7455) );
  INV_X1 U7755 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n7454) );
  INV_X1 U7756 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n13581) );
  INV_X1 U7757 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n13582) );
  INV_X1 U7758 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n13583) );
  INV_X1 U7759 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7891) );
  INV_X1 U7760 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n10009) );
  NOR2_X1 U7761 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7653) );
  NOR2_X1 U7762 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n7652) );
  NOR2_X1 U7763 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7651) );
  OAI211_X1 U7764 ( .C1(n12830), .C2(n7838), .A(n7837), .B(1'b1), .ZN(n12835)
         );
  XNOR2_X2 U7766 ( .A(n7447), .B(n7434), .ZN(n9680) );
  NAND2_X1 U7767 ( .A1(n9649), .A2(n9648), .ZN(n11972) );
  OAI21_X1 U7768 ( .B1(n9649), .B2(n15323), .A(n7448), .ZN(n9651) );
  AOI21_X1 U7769 ( .B1(n7449), .B2(n11466), .A(n7436), .ZN(n7448) );
  NAND3_X1 U7770 ( .A1(n9650), .A2(n16477), .A3(n9651), .ZN(n8293) );
  NAND2_X1 U7771 ( .A1(n7450), .A2(n15323), .ZN(n9650) );
  INV_X1 U7772 ( .A(n11972), .ZN(n7450) );
  OAI21_X2 U7773 ( .B1(n15497), .B2(n8290), .A(n7541), .ZN(n15468) );
  NAND4_X1 U7774 ( .A1(n13581), .A2(n13582), .A3(n13583), .A4(n9335), .ZN(
        n7452) );
  NAND4_X1 U7775 ( .A1(n7455), .A2(n13589), .A3(n7454), .A4(n9441), .ZN(n7453)
         );
  NAND4_X2 U7776 ( .A1(n7456), .A2(n9258), .A3(n9259), .A4(n9257), .ZN(n9636)
         );
  INV_X2 U7777 ( .A(n9636), .ZN(n9269) );
  INV_X1 U7778 ( .A(n9498), .ZN(n9499) );
  OAI21_X2 U7779 ( .B1(n8551), .B2(P2_IR_REG_27__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7698) );
  NOR2_X2 U7780 ( .A1(n15527), .A2(n15528), .ZN(n15526) );
  INV_X1 U7781 ( .A(n9477), .ZN(n7457) );
  AND2_X4 U7782 ( .A1(n7904), .A2(n13854), .ZN(n9813) );
  AND3_X2 U7783 ( .A1(n9280), .A2(n9279), .A3(n9278), .ZN(n16374) );
  NOR2_X1 U7784 ( .A1(n9131), .A2(n8202), .ZN(n8201) );
  INV_X1 U7785 ( .A(n9130), .ZN(n8202) );
  NAND2_X1 U7786 ( .A1(n8010), .A2(n8008), .ZN(n9010) );
  AOI21_X1 U7787 ( .B1(n8012), .B2(n8014), .A(n8009), .ZN(n8008) );
  INV_X1 U7788 ( .A(n8993), .ZN(n8009) );
  NAND2_X1 U7789 ( .A1(n10297), .A2(n10946), .ZN(n10949) );
  AND2_X1 U7790 ( .A1(n13380), .A2(n13091), .ZN(n12764) );
  NOR2_X1 U7791 ( .A1(n9845), .A2(n7725), .ZN(n7724) );
  INV_X1 U7792 ( .A(n9824), .ZN(n7725) );
  NAND2_X1 U7793 ( .A1(n10488), .A2(n8155), .ZN(n8586) );
  OR2_X1 U7794 ( .A1(n9075), .A2(n9074), .ZN(n9091) );
  NAND2_X1 U7795 ( .A1(n10272), .A2(n12728), .ZN(n16352) );
  OR2_X1 U7796 ( .A1(n14193), .A2(n9088), .ZN(n9145) );
  NAND2_X1 U7797 ( .A1(n14581), .A2(n8910), .ZN(n14564) );
  NAND2_X1 U7798 ( .A1(n14030), .A2(n7514), .ZN(n8342) );
  NOR2_X1 U7799 ( .A1(n14097), .A2(n7468), .ZN(n8329) );
  AOI21_X1 U7800 ( .B1(n8323), .B2(n8327), .A(n14102), .ZN(n8322) );
  INV_X1 U7801 ( .A(n14190), .ZN(n8310) );
  AND2_X1 U7802 ( .A1(n10009), .A2(n9957), .ZN(n7858) );
  AND2_X1 U7803 ( .A1(n8596), .A2(n7687), .ZN(n7976) );
  AND2_X1 U7804 ( .A1(n8523), .A2(n8544), .ZN(n7687) );
  INV_X1 U7805 ( .A(n8032), .ZN(n8031) );
  OAI21_X1 U7806 ( .B1(n8034), .B2(n8033), .A(n9067), .ZN(n8032) );
  AOI21_X1 U7807 ( .B1(n8021), .B2(n8023), .A(n8020), .ZN(n8019) );
  INV_X1 U7808 ( .A(n8844), .ZN(n8020) );
  INV_X1 U7809 ( .A(n8026), .ZN(n8021) );
  AOI21_X1 U7810 ( .B1(n8843), .B2(n8842), .A(n8841), .ZN(n8844) );
  INV_X1 U7811 ( .A(n8023), .ZN(n8022) );
  AOI21_X1 U7812 ( .B1(n8702), .B2(n8400), .A(n7539), .ZN(n8399) );
  INV_X1 U7813 ( .A(n8681), .ZN(n8400) );
  NOR2_X1 U7814 ( .A1(n8701), .A2(n8677), .ZN(n7992) );
  NOR2_X1 U7815 ( .A1(n8275), .A2(n13650), .ZN(n8583) );
  INV_X1 U7816 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15940) );
  NAND2_X1 U7817 ( .A1(n15937), .A2(n15938), .ZN(n15939) );
  NAND2_X1 U7818 ( .A1(n12848), .A2(n7875), .ZN(n7874) );
  NAND2_X1 U7819 ( .A1(n8497), .A2(n8499), .ZN(n7875) );
  OR2_X1 U7820 ( .A1(n13384), .A2(n12574), .ZN(n12576) );
  INV_X1 U7821 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8502) );
  OR2_X1 U7822 ( .A1(n13113), .A2(n13125), .ZN(n12726) );
  AOI21_X1 U7823 ( .B1(n7466), .B2(n10192), .A(n7533), .ZN(n7939) );
  NAND2_X1 U7824 ( .A1(n13138), .A2(n12983), .ZN(n12716) );
  OR2_X1 U7825 ( .A1(n13330), .A2(n12915), .ZN(n12711) );
  OR2_X1 U7826 ( .A1(n13164), .A2(n12891), .ZN(n10294) );
  OR2_X1 U7827 ( .A1(n10142), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n10158) );
  OR2_X1 U7828 ( .A1(n13216), .A2(n13227), .ZN(n12700) );
  AND2_X1 U7829 ( .A1(n11377), .A2(n10303), .ZN(n10297) );
  AND4_X1 U7830 ( .A1(n9920), .A2(n9885), .A3(n9897), .A4(n9884), .ZN(n7461)
         );
  AND2_X1 U7831 ( .A1(n7850), .A2(n9789), .ZN(n7857) );
  AND2_X1 U7832 ( .A1(n9790), .A2(n9746), .ZN(n7850) );
  NAND2_X1 U7833 ( .A1(n10411), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9798) );
  NAND2_X1 U7834 ( .A1(n8185), .A2(n8184), .ZN(n9733) );
  AOI21_X1 U7835 ( .B1(n8186), .B2(n8189), .A(n7556), .ZN(n8184) );
  NAND2_X1 U7836 ( .A1(n14542), .A2(n7948), .ZN(n7810) );
  NAND2_X1 U7837 ( .A1(n7948), .A2(n7467), .ZN(n7947) );
  AOI21_X1 U7838 ( .B1(n8199), .B2(n8201), .A(n7543), .ZN(n8198) );
  INV_X1 U7839 ( .A(n9129), .ZN(n8199) );
  INV_X1 U7840 ( .A(n8201), .ZN(n8200) );
  NOR2_X1 U7841 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n7649) );
  INV_X1 U7842 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8541) );
  NOR2_X1 U7843 ( .A1(n15451), .A2(n8413), .ZN(n8412) );
  NAND2_X1 U7844 ( .A1(n9676), .A2(n9603), .ZN(n15258) );
  OR2_X1 U7845 ( .A1(n15651), .A2(n15301), .ZN(n9603) );
  NAND2_X1 U7846 ( .A1(n8440), .A2(n8438), .ZN(n8437) );
  INV_X1 U7847 ( .A(n15498), .ZN(n8438) );
  NOR2_X1 U7848 ( .A1(n15601), .A2(n8430), .ZN(n8429) );
  INV_X1 U7849 ( .A(n9497), .ZN(n8430) );
  NAND2_X1 U7850 ( .A1(n9012), .A2(n9011), .ZN(n9017) );
  NAND2_X1 U7851 ( .A1(n9007), .A2(SI_24_), .ZN(n9012) );
  OR2_X2 U7852 ( .A1(n9017), .A2(n9016), .ZN(n9032) );
  INV_X1 U7853 ( .A(n9620), .ZN(n9616) );
  NAND2_X1 U7854 ( .A1(n9614), .A2(n13801), .ZN(n9620) );
  NAND2_X1 U7855 ( .A1(n9499), .A2(n9500), .ZN(n9509) );
  XNOR2_X1 U7856 ( .A(n8801), .B(n13629), .ZN(n8800) );
  INV_X1 U7857 ( .A(n8740), .ZN(n8741) );
  XNOR2_X1 U7858 ( .A(n8610), .B(SI_3_), .ZN(n8609) );
  AOI21_X1 U7859 ( .B1(n7846), .B2(n12794), .A(n7559), .ZN(n7845) );
  INV_X1 U7860 ( .A(n12845), .ZN(n7863) );
  NAND2_X1 U7861 ( .A1(n12914), .A2(n13188), .ZN(n7839) );
  AND2_X1 U7862 ( .A1(n8141), .A2(n13118), .ZN(n7790) );
  AND2_X1 U7863 ( .A1(n8142), .A2(n12581), .ZN(n8141) );
  AND3_X1 U7864 ( .A1(n7564), .A2(n7807), .A3(n7782), .ZN(n12766) );
  NOR2_X1 U7865 ( .A1(n12764), .A2(n12765), .ZN(n7782) );
  INV_X1 U7866 ( .A(n11031), .ZN(n7747) );
  NAND2_X1 U7867 ( .A1(n11524), .A2(n11534), .ZN(n8075) );
  NOR2_X1 U7868 ( .A1(n13016), .A2(n16159), .ZN(n16177) );
  NOR2_X1 U7869 ( .A1(n13125), .A2(n16350), .ZN(n10273) );
  AND2_X1 U7870 ( .A1(n10287), .A2(n12662), .ZN(n8132) );
  OR2_X1 U7871 ( .A1(n16593), .A2(n12733), .ZN(n10809) );
  AND2_X1 U7872 ( .A1(n10264), .A2(n12580), .ZN(n16349) );
  NAND2_X1 U7873 ( .A1(n10090), .A2(n10089), .ZN(n12875) );
  INV_X1 U7874 ( .A(n12569), .ZN(n12562) );
  INV_X1 U7875 ( .A(n9800), .ZN(n12568) );
  NAND2_X1 U7876 ( .A1(n10320), .A2(n10332), .ZN(n12527) );
  OR2_X1 U7877 ( .A1(n13841), .A2(n13843), .ZN(n9755) );
  OAI21_X1 U7878 ( .B1(n10241), .B2(n10240), .A(n10243), .ZN(n12556) );
  NOR2_X1 U7879 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n9752) );
  AND2_X1 U7880 ( .A1(n9751), .A2(n10255), .ZN(n8120) );
  NAND2_X1 U7881 ( .A1(n10133), .A2(n7614), .ZN(n10150) );
  INV_X1 U7882 ( .A(n10136), .ZN(n7793) );
  INV_X1 U7883 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7877) );
  AOI21_X1 U7884 ( .B1(n7743), .B2(n7745), .A(n7617), .ZN(n7741) );
  XNOR2_X1 U7885 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n9901) );
  NAND2_X1 U7886 ( .A1(n10448), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9882) );
  NAND2_X1 U7887 ( .A1(n9863), .A2(n9848), .ZN(n9864) );
  NAND2_X1 U7888 ( .A1(n10446), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n9848) );
  AOI21_X1 U7889 ( .B1(n7724), .B2(n7722), .A(n7549), .ZN(n7721) );
  INV_X1 U7890 ( .A(n9822), .ZN(n7722) );
  INV_X1 U7891 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9847) );
  XNOR2_X1 U7892 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n9844) );
  NAND2_X1 U7893 ( .A1(n10408), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9824) );
  NAND2_X1 U7894 ( .A1(n13924), .A2(n8161), .ZN(n8160) );
  INV_X1 U7895 ( .A(n12549), .ZN(n8162) );
  AOI21_X1 U7896 ( .B1(n13924), .B2(n12549), .A(n8165), .ZN(n8164) );
  INV_X1 U7897 ( .A(n13857), .ZN(n8165) );
  NOR2_X1 U7898 ( .A1(n7536), .A2(n7675), .ZN(n7674) );
  NOR2_X1 U7899 ( .A1(n13932), .A2(n13869), .ZN(n7675) );
  INV_X1 U7900 ( .A(n8599), .ZN(n14219) );
  INV_X1 U7901 ( .A(n8831), .ZN(n9153) );
  NAND2_X2 U7902 ( .A1(n8561), .A2(n12791), .ZN(n8831) );
  INV_X1 U7903 ( .A(n8831), .ZN(n7946) );
  NAND2_X1 U7904 ( .A1(n14776), .A2(n8562), .ZN(n14218) );
  NAND2_X1 U7905 ( .A1(n8529), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8538) );
  NOR3_X1 U7906 ( .A1(n14495), .A2(n7958), .A3(n14234), .ZN(n14439) );
  NAND2_X1 U7907 ( .A1(n9145), .A2(n9089), .ZN(n14312) );
  AND2_X1 U7908 ( .A1(n8223), .A2(n7692), .ZN(n7691) );
  NOR2_X1 U7909 ( .A1(n14462), .A2(n8224), .ZN(n8223) );
  NAND2_X1 U7910 ( .A1(n14478), .A2(n7693), .ZN(n7692) );
  NAND2_X1 U7911 ( .A1(n14489), .A2(n9030), .ZN(n14477) );
  OR2_X1 U7912 ( .A1(n14688), .A2(n13958), .ZN(n9133) );
  NAND2_X1 U7913 ( .A1(n14608), .A2(n8893), .ZN(n14582) );
  XNOR2_X1 U7914 ( .A(n14326), .B(n7685), .ZN(n7684) );
  NAND2_X1 U7915 ( .A1(n14233), .A2(n14232), .ZN(n14435) );
  AND2_X1 U7916 ( .A1(n14785), .A2(n9169), .ZN(n15819) );
  NAND2_X1 U7917 ( .A1(n9707), .A2(n9706), .ZN(n11177) );
  AND2_X1 U7918 ( .A1(n9704), .A2(n9716), .ZN(n9707) );
  AND2_X1 U7919 ( .A1(n8377), .A2(n8371), .ZN(n8370) );
  INV_X1 U7920 ( .A(n8378), .ZN(n8377) );
  NAND2_X1 U7921 ( .A1(n8375), .A2(n8372), .ZN(n8371) );
  OAI21_X1 U7922 ( .B1(n15015), .B2(n8380), .A(n8379), .ZN(n8378) );
  NAND2_X1 U7923 ( .A1(n16609), .A2(n14812), .ZN(n14814) );
  NAND2_X1 U7924 ( .A1(n15651), .A2(n15301), .ZN(n9676) );
  OR2_X1 U7925 ( .A1(n15464), .A2(n8415), .ZN(n8408) );
  NAND2_X1 U7926 ( .A1(n15464), .A2(n8412), .ZN(n8411) );
  NAND2_X1 U7927 ( .A1(n15664), .A2(n14952), .ZN(n8423) );
  XNOR2_X1 U7928 ( .A(n15675), .B(n14953), .ZN(n15498) );
  OR2_X1 U7929 ( .A1(n15694), .A2(n9553), .ZN(n9554) );
  NAND2_X1 U7930 ( .A1(n8281), .A2(n9668), .ZN(n8280) );
  INV_X1 U7931 ( .A(n8283), .ZN(n8281) );
  OR2_X1 U7932 ( .A1(n15699), .A2(n14934), .ZN(n9542) );
  NAND2_X1 U7933 ( .A1(n15734), .A2(n8450), .ZN(n15624) );
  AND2_X1 U7934 ( .A1(n15625), .A2(n9471), .ZN(n8450) );
  XNOR2_X1 U7935 ( .A(n15732), .B(n15314), .ZN(n15249) );
  INV_X1 U7936 ( .A(n9261), .ZN(n8158) );
  NAND2_X1 U7937 ( .A1(n9091), .A2(n9076), .ZN(n14778) );
  NOR2_X1 U7938 ( .A1(n16009), .A2(n16008), .ZN(n16015) );
  AND2_X1 U7939 ( .A1(n16007), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n16008) );
  OAI22_X1 U7940 ( .A1(n16034), .A2(n7627), .B1(n16033), .B2(n7630), .ZN(n7629) );
  AND2_X1 U7941 ( .A1(n16033), .A2(n7630), .ZN(n7627) );
  INV_X1 U7942 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7630) );
  OAI21_X1 U7943 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n16032), .A(n16031), .ZN(
        n16038) );
  INV_X1 U7944 ( .A(n12992), .ZN(n12133) );
  NAND2_X1 U7945 ( .A1(n13112), .A2(n13111), .ZN(n13319) );
  OR2_X1 U7946 ( .A1(n13107), .A2(n7572), .ZN(n13112) );
  NAND2_X1 U7947 ( .A1(n11897), .A2(n7683), .ZN(n12305) );
  NAND2_X1 U7948 ( .A1(n7978), .A2(n7680), .ZN(n7683) );
  AND2_X1 U7949 ( .A1(n8170), .A2(n7563), .ZN(n7978) );
  NAND2_X1 U7950 ( .A1(n7681), .A2(n11879), .ZN(n7680) );
  INV_X1 U7951 ( .A(n8174), .ZN(n8173) );
  OAI21_X1 U7952 ( .B1(n8176), .B2(n8175), .A(n13893), .ZN(n8174) );
  INV_X1 U7953 ( .A(n12541), .ZN(n8175) );
  NAND2_X1 U7954 ( .A1(n7801), .A2(n7800), .ZN(n7799) );
  NAND2_X1 U7955 ( .A1(n16001), .A2(n16000), .ZN(n16004) );
  NAND2_X1 U7956 ( .A1(n16016), .A2(n16017), .ZN(n16018) );
  NOR2_X1 U7957 ( .A1(n16020), .A2(n16021), .ZN(n16022) );
  INV_X1 U7958 ( .A(n14035), .ZN(n7763) );
  OAI21_X1 U7959 ( .B1(n15059), .B2(n15058), .A(n15057), .ZN(n15061) );
  NAND2_X1 U7960 ( .A1(n14058), .A2(n7511), .ZN(n8345) );
  NAND2_X1 U7961 ( .A1(n15089), .A2(n15087), .ZN(n7899) );
  NOR2_X1 U7962 ( .A1(n8471), .A2(n15091), .ZN(n8472) );
  NAND2_X1 U7963 ( .A1(n8471), .A2(n15091), .ZN(n8470) );
  NOR2_X1 U7964 ( .A1(n8327), .A2(n14103), .ZN(n8326) );
  NAND2_X1 U7965 ( .A1(n8321), .A2(n8320), .ZN(n8319) );
  INV_X1 U7966 ( .A(n8326), .ZN(n8320) );
  INV_X1 U7967 ( .A(n8322), .ZN(n8321) );
  NAND2_X1 U7968 ( .A1(n8329), .A2(n8328), .ZN(n8325) );
  NAND2_X1 U7969 ( .A1(n15104), .A2(n15102), .ZN(n7894) );
  NAND2_X1 U7970 ( .A1(n15103), .A2(n7895), .ZN(n7893) );
  NAND2_X1 U7971 ( .A1(n15117), .A2(n15119), .ZN(n7901) );
  NOR2_X1 U7972 ( .A1(n15120), .A2(n15123), .ZN(n8466) );
  NAND2_X1 U7973 ( .A1(n15123), .A2(n15120), .ZN(n8465) );
  NAND2_X1 U7974 ( .A1(n15131), .A2(n15134), .ZN(n7882) );
  NAND2_X1 U7975 ( .A1(n7497), .A2(n7881), .ZN(n7880) );
  AND2_X1 U7976 ( .A1(n15133), .A2(n7883), .ZN(n7881) );
  AND2_X1 U7977 ( .A1(n15151), .A2(n15142), .ZN(n8456) );
  INV_X1 U7978 ( .A(n8955), .ZN(n8014) );
  NOR2_X1 U7979 ( .A1(n8845), .A2(n8024), .ZN(n8023) );
  INV_X1 U7980 ( .A(n8802), .ZN(n8024) );
  NAND2_X1 U7981 ( .A1(n8513), .A2(n8842), .ZN(n8845) );
  INV_X1 U7982 ( .A(n7731), .ZN(n7730) );
  OAI21_X1 U7983 ( .B1(n10082), .B2(n7732), .A(n10102), .ZN(n7731) );
  INV_X1 U7984 ( .A(n10084), .ZN(n7732) );
  AND2_X1 U7985 ( .A1(n8309), .A2(n8306), .ZN(n8303) );
  INV_X1 U7986 ( .A(n8307), .ZN(n8306) );
  OR2_X1 U7987 ( .A1(n8309), .A2(n8312), .ZN(n8302) );
  INV_X1 U7988 ( .A(n11273), .ZN(n8354) );
  INV_X1 U7989 ( .A(n15179), .ZN(n7888) );
  NAND2_X1 U7990 ( .A1(n15176), .A2(n15178), .ZN(n8477) );
  NAND2_X1 U7991 ( .A1(n15179), .A2(n7887), .ZN(n7886) );
  NAND2_X1 U7992 ( .A1(n8746), .A2(n13437), .ZN(n8766) );
  AND2_X1 U7993 ( .A1(n8399), .A2(n7999), .ZN(n7997) );
  INV_X1 U7994 ( .A(n8622), .ZN(n8623) );
  OAI21_X1 U7995 ( .B1(n8595), .B2(n8609), .A(n8611), .ZN(n7985) );
  NAND2_X1 U7996 ( .A1(n7635), .A2(n15952), .ZN(n15955) );
  NAND2_X1 U7997 ( .A1(n15951), .A2(n15950), .ZN(n7635) );
  NAND2_X1 U7998 ( .A1(n7826), .A2(n12819), .ZN(n7824) );
  OR2_X1 U7999 ( .A1(n16117), .A2(n11003), .ZN(n8087) );
  INV_X1 U8000 ( .A(n16121), .ZN(n8056) );
  INV_X1 U8001 ( .A(n16122), .ZN(n8053) );
  NAND2_X1 U8002 ( .A1(n16138), .A2(n11254), .ZN(n7748) );
  NAND2_X1 U8003 ( .A1(n16133), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8037) );
  OAI21_X1 U8004 ( .B1(n16133), .B2(P3_REG2_REG_6__SCAN_IN), .A(n16143), .ZN(
        n8038) );
  NAND2_X1 U8005 ( .A1(n13013), .A2(n13012), .ZN(n13015) );
  INV_X1 U8006 ( .A(n10270), .ZN(n10990) );
  NOR2_X1 U8007 ( .A1(n10239), .A2(n13123), .ZN(n7912) );
  INV_X1 U8008 ( .A(n7913), .ZN(n7910) );
  NOR2_X1 U8009 ( .A1(n13104), .A2(n7914), .ZN(n7913) );
  INV_X1 U8010 ( .A(n10226), .ZN(n7914) );
  OR2_X1 U8011 ( .A1(n10225), .A2(n8270), .ZN(n10226) );
  INV_X1 U8012 ( .A(n10179), .ZN(n7938) );
  NAND2_X1 U8013 ( .A1(n8271), .A2(n8270), .ZN(n12717) );
  INV_X1 U8014 ( .A(n10178), .ZN(n7940) );
  INV_X1 U8015 ( .A(n13162), .ZN(n12585) );
  NAND2_X1 U8016 ( .A1(n10293), .A2(n10148), .ZN(n13182) );
  OR2_X1 U8017 ( .A1(n13349), .A2(n12945), .ZN(n12820) );
  INV_X1 U8018 ( .A(n8138), .ZN(n8136) );
  NOR2_X1 U8019 ( .A1(n7921), .A2(n7918), .ZN(n7917) );
  INV_X1 U8020 ( .A(n10052), .ZN(n7918) );
  INV_X1 U8021 ( .A(n7922), .ZN(n7921) );
  NOR2_X1 U8022 ( .A1(n13239), .A2(n7923), .ZN(n7922) );
  INV_X1 U8023 ( .A(n10068), .ZN(n7923) );
  NOR2_X1 U8024 ( .A1(n10288), .A2(n12684), .ZN(n8138) );
  NAND2_X1 U8025 ( .A1(n9994), .A2(n13690), .ZN(n10013) );
  INV_X1 U8026 ( .A(n9995), .ZN(n9994) );
  INV_X1 U8027 ( .A(n9963), .ZN(n7927) );
  AND2_X1 U8028 ( .A1(n12194), .A2(n9930), .ZN(n7930) );
  NAND2_X1 U8029 ( .A1(n8117), .A2(n8115), .ZN(n12597) );
  INV_X1 U8030 ( .A(n8119), .ZN(n8117) );
  NOR2_X1 U8031 ( .A1(n8118), .A2(n8116), .ZN(n8115) );
  NAND2_X1 U8032 ( .A1(n8116), .A2(n12997), .ZN(n12591) );
  INV_X1 U8033 ( .A(n11377), .ZN(n12594) );
  NAND2_X1 U8034 ( .A1(n12597), .A2(n12591), .ZN(n12739) );
  NAND2_X1 U8035 ( .A1(n12223), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n10195) );
  INV_X1 U8036 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n9750) );
  INV_X1 U8037 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8496) );
  INV_X1 U8038 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n10255) );
  INV_X1 U8039 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9986) );
  INV_X1 U8040 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9954) );
  NOR2_X1 U8041 ( .A1(n9903), .A2(n8266), .ZN(n8265) );
  INV_X1 U8042 ( .A(n9882), .ZN(n8266) );
  INV_X1 U8043 ( .A(n9901), .ZN(n9903) );
  NAND2_X1 U8044 ( .A1(n10460), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n9925) );
  NAND2_X1 U8045 ( .A1(n9789), .A2(n9790), .ZN(n9801) );
  AND2_X1 U8046 ( .A1(n8997), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n9021) );
  XNOR2_X1 U8047 ( .A(n7433), .B(n11348), .ZN(n10374) );
  NOR2_X1 U8048 ( .A1(n9134), .A2(n8215), .ZN(n8214) );
  INV_X1 U8049 ( .A(n9133), .ZN(n8215) );
  NOR2_X1 U8050 ( .A1(n12513), .A2(n8237), .ZN(n8236) );
  INV_X1 U8051 ( .A(n8857), .ZN(n8237) );
  NOR2_X1 U8052 ( .A1(n14061), .A2(n7961), .ZN(n7960) );
  INV_X1 U8053 ( .A(n7962), .ZN(n7961) );
  INV_X1 U8054 ( .A(n8183), .ZN(n14285) );
  NAND2_X1 U8055 ( .A1(n7686), .A2(n8330), .ZN(n8536) );
  AND2_X1 U8056 ( .A1(n7976), .A2(n7975), .ZN(n7686) );
  NOR2_X1 U8057 ( .A1(n7523), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n7975) );
  INV_X1 U8058 ( .A(n8627), .ZN(n8647) );
  INV_X1 U8059 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8523) );
  INV_X1 U8060 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8522) );
  NOR2_X1 U8061 ( .A1(n15015), .A2(n8376), .ZN(n8375) );
  INV_X1 U8062 ( .A(n14951), .ZN(n8376) );
  NOR2_X1 U8063 ( .A1(n11268), .A2(n8354), .ZN(n8350) );
  INV_X1 U8064 ( .A(n11278), .ZN(n8355) );
  NOR2_X1 U8065 ( .A1(n16399), .A2(n8354), .ZN(n8353) );
  XNOR2_X1 U8066 ( .A(n15427), .B(n15424), .ZN(n15231) );
  XNOR2_X1 U8067 ( .A(n15659), .B(n15302), .ZN(n15256) );
  NOR2_X1 U8068 ( .A1(n9662), .A2(n8288), .ZN(n8287) );
  INV_X1 U8069 ( .A(n9661), .ZN(n8288) );
  NOR2_X1 U8070 ( .A1(n16531), .A2(n15078), .ZN(n8109) );
  AND2_X1 U8071 ( .A1(n16475), .A2(n16493), .ZN(n11772) );
  OR2_X1 U8072 ( .A1(n15573), .A2(n15699), .ZN(n15565) );
  NAND2_X1 U8073 ( .A1(n8029), .A2(n8028), .ZN(n9075) );
  AOI21_X1 U8074 ( .B1(n8031), .B2(n8033), .A(n7619), .ZN(n8028) );
  INV_X1 U8075 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9201) );
  XNOR2_X1 U8076 ( .A(n9010), .B(n9008), .ZN(n9007) );
  INV_X1 U8077 ( .A(n8397), .ZN(n8395) );
  NAND2_X1 U8078 ( .A1(n8940), .A2(n8939), .ZN(n8953) );
  OR2_X1 U8079 ( .A1(n8938), .A2(n7989), .ZN(n8939) );
  NAND2_X1 U8080 ( .A1(n8937), .A2(n8936), .ZN(n8940) );
  NAND2_X1 U8081 ( .A1(n8885), .A2(n8884), .ZN(n8914) );
  NAND2_X1 U8082 ( .A1(n8025), .A2(n8802), .ZN(n8820) );
  XNOR2_X1 U8083 ( .A(n8820), .B(SI_14_), .ZN(n8819) );
  OAI21_X1 U8084 ( .B1(n8723), .B2(n8722), .A(n8721), .ZN(n8742) );
  NAND2_X1 U8085 ( .A1(n8426), .A2(n8428), .ZN(n8679) );
  AOI21_X1 U8086 ( .B1(n8662), .B2(n7477), .A(n7538), .ZN(n8428) );
  INV_X1 U8087 ( .A(n8626), .ZN(n8233) );
  NAND2_X1 U8088 ( .A1(n8230), .A2(n8626), .ZN(n8645) );
  NAND2_X1 U8089 ( .A1(n8624), .A2(n8623), .ZN(n8230) );
  XNOR2_X1 U8090 ( .A(n15955), .B(n16130), .ZN(n15957) );
  AOI22_X1 U8091 ( .A1(n15987), .A2(n15986), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n16150), .ZN(n15995) );
  AOI21_X1 U8092 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n16040), .A(n16039), .ZN(
        n16053) );
  INV_X1 U8093 ( .A(n12841), .ZN(n7869) );
  AOI21_X1 U8094 ( .B1(n7832), .B2(n11687), .A(n7831), .ZN(n7830) );
  NAND2_X1 U8095 ( .A1(n10122), .A2(n13666), .ZN(n10142) );
  INV_X1 U8096 ( .A(n10123), .ZN(n10122) );
  OAI21_X1 U8097 ( .B1(n12203), .B2(n8482), .A(n12396), .ZN(n8481) );
  INV_X1 U8098 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n13679) );
  AOI22_X1 U8099 ( .A1(n12136), .A2(n12135), .B1(n12134), .B2(n12993), .ZN(
        n12137) );
  NAND2_X1 U8100 ( .A1(n7849), .A2(n7848), .ZN(n7847) );
  NAND2_X1 U8101 ( .A1(n7847), .A2(n7846), .ZN(n12935) );
  INV_X1 U8102 ( .A(n12811), .ZN(n8488) );
  NOR2_X1 U8103 ( .A1(n8488), .A2(n8485), .ZN(n8484) );
  INV_X1 U8104 ( .A(n12809), .ZN(n8485) );
  NOR2_X1 U8105 ( .A1(n11513), .A2(n7500), .ZN(n8491) );
  AOI21_X1 U8106 ( .B1(n7551), .B2(n8142), .A(n7788), .ZN(n8140) );
  AND2_X1 U8107 ( .A1(n7704), .A2(n7702), .ZN(n12734) );
  AOI21_X1 U8108 ( .B1(n7789), .B2(n7703), .A(n12764), .ZN(n7702) );
  INV_X1 U8109 ( .A(n12576), .ZN(n7703) );
  INV_X1 U8110 ( .A(n9813), .ZN(n11436) );
  AND3_X1 U8111 ( .A1(n10146), .A2(n10145), .A3(n10144), .ZN(n12867) );
  AND4_X1 U8112 ( .A1(n9972), .A2(n9971), .A3(n9970), .A4(n9969), .ZN(n12228)
         );
  AND4_X1 U8113 ( .A1(n9950), .A2(n9949), .A3(n9948), .A4(n9947), .ZN(n12267)
         );
  OAI22_X1 U8114 ( .A1(n9814), .A2(n10991), .B1(n7904), .B2(n7903), .ZN(n8119)
         );
  NAND2_X1 U8115 ( .A1(n13854), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7903) );
  NAND2_X1 U8116 ( .A1(n8040), .A2(n8039), .ZN(n11245) );
  OAI21_X1 U8117 ( .B1(n11100), .B2(P3_REG2_REG_4__SCAN_IN), .A(n11113), .ZN(
        n8040) );
  NAND2_X1 U8118 ( .A1(n7769), .A2(n7508), .ZN(n8082) );
  NAND2_X1 U8119 ( .A1(n8082), .A2(n8081), .ZN(n16138) );
  INV_X1 U8120 ( .A(n16135), .ZN(n8081) );
  XNOR2_X1 U8121 ( .A(n7748), .B(n11526), .ZN(n11255) );
  NOR2_X1 U8122 ( .A1(n9877), .A2(n11255), .ZN(n11535) );
  XNOR2_X1 U8123 ( .A(n11525), .B(n11534), .ZN(n11249) );
  NOR2_X1 U8124 ( .A1(n11244), .A2(n8072), .ZN(n8071) );
  INV_X1 U8125 ( .A(n16139), .ZN(n8072) );
  NOR2_X1 U8126 ( .A1(n8070), .A2(n8069), .ZN(n8068) );
  INV_X1 U8127 ( .A(n8075), .ZN(n8069) );
  INV_X1 U8128 ( .A(n7622), .ZN(n8070) );
  INV_X1 U8129 ( .A(n11669), .ZN(n8065) );
  NOR2_X1 U8130 ( .A1(n8068), .A2(n11669), .ZN(n8064) );
  OR2_X1 U8131 ( .A1(n11824), .A2(n11823), .ZN(n13013) );
  OR2_X1 U8132 ( .A1(n13031), .A2(n16187), .ZN(n8080) );
  AND2_X1 U8133 ( .A1(n13031), .A2(n16187), .ZN(n8079) );
  NOR2_X1 U8134 ( .A1(n16198), .A2(n16600), .ZN(n16197) );
  NAND2_X1 U8135 ( .A1(n16192), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n16191) );
  XNOR2_X1 U8136 ( .A(n13021), .B(n13055), .ZN(n16235) );
  NOR2_X1 U8137 ( .A1(n16232), .A2(n13020), .ZN(n13022) );
  NOR2_X1 U8138 ( .A1(n16227), .A2(n8059), .ZN(n16247) );
  AND2_X1 U8139 ( .A1(n13037), .A2(n13055), .ZN(n8059) );
  OR2_X1 U8140 ( .A1(n16247), .A2(n16246), .ZN(n8058) );
  NOR2_X1 U8141 ( .A1(n16265), .A2(n16264), .ZN(n16262) );
  OR2_X1 U8142 ( .A1(n10234), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n13092) );
  AND2_X1 U8143 ( .A1(n13104), .A2(n12718), .ZN(n8144) );
  NAND2_X1 U8144 ( .A1(n10224), .A2(n13119), .ZN(n13120) );
  INV_X1 U8145 ( .A(n12716), .ZN(n12584) );
  NAND2_X1 U8146 ( .A1(n12716), .A2(n12714), .ZN(n13132) );
  OR2_X1 U8147 ( .A1(n7942), .A2(n7466), .ZN(n13144) );
  OR2_X1 U8148 ( .A1(n13400), .A2(n13188), .ZN(n13158) );
  OAI21_X1 U8149 ( .B1(n10100), .B2(n7933), .A(n7931), .ZN(n13186) );
  INV_X1 U8150 ( .A(n7932), .ZN(n7931) );
  OAI21_X1 U8151 ( .B1(n7495), .B2(n7933), .A(n12820), .ZN(n7932) );
  OR2_X1 U8152 ( .A1(n10128), .A2(n7934), .ZN(n7933) );
  AND2_X1 U8153 ( .A1(n12820), .A2(n12696), .ZN(n13201) );
  NAND2_X1 U8154 ( .A1(n12700), .A2(n12695), .ZN(n13213) );
  NAND2_X1 U8155 ( .A1(n10100), .A2(n7495), .ZN(n13212) );
  INV_X1 U8156 ( .A(n10100), .ZN(n7936) );
  INV_X1 U8157 ( .A(n13252), .ZN(n13226) );
  AND4_X1 U8158 ( .A1(n10097), .A2(n10096), .A3(n10095), .A4(n10094), .ZN(
        n13237) );
  NAND2_X1 U8159 ( .A1(n13265), .A2(n8138), .ZN(n13241) );
  NAND2_X1 U8160 ( .A1(n10286), .A2(n7605), .ZN(n8133) );
  AND2_X1 U8161 ( .A1(n10019), .A2(n12662), .ZN(n13297) );
  OR2_X1 U8162 ( .A1(n16594), .A2(n12990), .ZN(n12658) );
  OAI21_X1 U8163 ( .B1(n12451), .B2(n10002), .A(n12800), .ZN(n13300) );
  AND2_X1 U8164 ( .A1(n12658), .A2(n12799), .ZN(n12796) );
  AND2_X1 U8165 ( .A1(n12651), .A2(n12646), .ZN(n12751) );
  NAND2_X1 U8166 ( .A1(n9931), .A2(n7930), .ZN(n12193) );
  INV_X1 U8167 ( .A(n9931), .ZN(n7929) );
  NAND2_X1 U8168 ( .A1(n9874), .A2(n13460), .ZN(n9890) );
  INV_X1 U8169 ( .A(n9875), .ZN(n9874) );
  OAI21_X1 U8170 ( .B1(n11696), .B2(n7906), .A(n7905), .ZN(n11867) );
  NAND2_X1 U8171 ( .A1(n9873), .A2(n7465), .ZN(n7906) );
  NAND2_X1 U8172 ( .A1(n7907), .A2(n7465), .ZN(n7905) );
  INV_X1 U8173 ( .A(n16349), .ZN(n13299) );
  AND3_X1 U8174 ( .A1(n9805), .A2(n9804), .A3(n9803), .ZN(n11081) );
  INV_X1 U8175 ( .A(n10989), .ZN(n10811) );
  AND4_X1 U8176 ( .A1(n9774), .A2(n9773), .A3(n9772), .A4(n9771), .ZN(n10278)
         );
  OR2_X1 U8177 ( .A1(n9814), .A2(n10996), .ZN(n9771) );
  OR2_X1 U8178 ( .A1(n10272), .A2(n12731), .ZN(n16350) );
  NOR2_X1 U8179 ( .A1(n10278), .A2(n11626), .ZN(n16311) );
  NAND2_X1 U8180 ( .A1(n10246), .A2(n10245), .ZN(n10343) );
  NAND2_X1 U8181 ( .A1(n10233), .A2(n10232), .ZN(n13113) );
  INV_X1 U8182 ( .A(n16593), .ZN(n16544) );
  OAI21_X1 U8183 ( .B1(n12556), .B2(n12555), .A(n12557), .ZN(n12567) );
  AND2_X1 U8184 ( .A1(n8503), .A2(n8150), .ZN(n8149) );
  NOR2_X1 U8185 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_28__SCAN_IN), .ZN(
        n8503) );
  INV_X1 U8186 ( .A(n8151), .ZN(n8150) );
  OAI21_X1 U8187 ( .B1(n10229), .B2(n10228), .A(n10230), .ZN(n10241) );
  OAI21_X1 U8188 ( .B1(n10194), .B2(n10193), .A(n10195), .ZN(n10210) );
  INV_X1 U8189 ( .A(n8077), .ZN(n9749) );
  NOR2_X1 U8190 ( .A1(n7856), .A2(n7855), .ZN(n7854) );
  INV_X1 U8191 ( .A(n7943), .ZN(n7855) );
  NAND2_X1 U8192 ( .A1(n7717), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7716) );
  NAND2_X1 U8193 ( .A1(n10154), .A2(n10153), .ZN(n10166) );
  NAND2_X1 U8194 ( .A1(n10256), .A2(n10255), .ZN(n10306) );
  INV_X1 U8195 ( .A(n10262), .ZN(n10256) );
  NAND2_X1 U8196 ( .A1(n10117), .A2(n10116), .ZN(n10131) );
  AND2_X1 U8197 ( .A1(n10263), .A2(n10262), .ZN(n10303) );
  NAND2_X1 U8198 ( .A1(n10086), .A2(n7878), .ZN(n10260) );
  XNOR2_X1 U8199 ( .A(n10087), .B(P3_IR_REG_19__SCAN_IN), .ZN(n13086) );
  NAND2_X1 U8200 ( .A1(n10086), .A2(n10085), .ZN(n10254) );
  NAND2_X1 U8201 ( .A1(n8253), .A2(n8252), .ZN(n10083) );
  AOI21_X1 U8202 ( .B1(n8255), .B2(n8257), .A(n7618), .ZN(n8252) );
  NAND2_X1 U8203 ( .A1(n10005), .A2(n10004), .ZN(n10006) );
  XNOR2_X1 U8204 ( .A(n10005), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n10003) );
  NOR2_X1 U8205 ( .A1(n9973), .A2(n7739), .ZN(n7738) );
  INV_X1 U8206 ( .A(n9955), .ZN(n7739) );
  OAI22_X1 U8207 ( .A1(n9941), .A2(n9940), .B1(P2_DATAO_REG_9__SCAN_IN), .B2(
        n10473), .ZN(n9953) );
  OR2_X1 U8208 ( .A1(n9899), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9922) );
  NOR2_X1 U8209 ( .A1(n9906), .A2(n8263), .ZN(n8262) );
  INV_X1 U8210 ( .A(n9902), .ZN(n8263) );
  NAND2_X1 U8211 ( .A1(n9883), .A2(n8265), .ZN(n8264) );
  NAND2_X1 U8212 ( .A1(n7721), .A2(n7526), .ZN(n7718) );
  AND2_X1 U8213 ( .A1(n9882), .A2(n9866), .ZN(n9867) );
  INV_X1 U8214 ( .A(n7724), .ZN(n7723) );
  AND2_X1 U8215 ( .A1(n9824), .A2(n9799), .ZN(n9822) );
  OR2_X1 U8216 ( .A1(n8812), .A2(n8811), .ZN(n8829) );
  INV_X1 U8217 ( .A(n11227), .ZN(n7973) );
  NOR2_X1 U8218 ( .A1(n13964), .A2(n8177), .ZN(n8176) );
  INV_X1 U8219 ( .A(n12538), .ZN(n8177) );
  XNOR2_X1 U8220 ( .A(n10884), .B(n14006), .ZN(n10371) );
  AND3_X1 U8221 ( .A1(n8167), .A2(n10377), .A3(n10885), .ZN(n8166) );
  NAND2_X1 U8222 ( .A1(n13951), .A2(n12544), .ZN(n13948) );
  NOR2_X1 U8223 ( .A1(n7668), .A2(n7974), .ZN(n7667) );
  INV_X1 U8224 ( .A(n11881), .ZN(n7783) );
  OR2_X1 U8225 ( .A1(n12306), .A2(n12307), .ZN(n8172) );
  NAND2_X1 U8226 ( .A1(n8827), .A2(n8826), .ZN(n14716) );
  OR2_X1 U8227 ( .A1(n14266), .A2(n14265), .ZN(n14267) );
  AND2_X1 U8228 ( .A1(n8950), .A2(n8949), .ZN(n14165) );
  XNOR2_X1 U8229 ( .A(n14234), .B(n14340), .ZN(n14314) );
  NAND2_X1 U8230 ( .A1(n14465), .A2(n9066), .ZN(n9738) );
  OR2_X1 U8231 ( .A1(n9733), .A2(n14312), .ZN(n9732) );
  NAND2_X1 U8232 ( .A1(n14477), .A2(n14478), .ZN(n14476) );
  AND2_X1 U8233 ( .A1(n8217), .A2(n14491), .ZN(n8216) );
  NAND2_X1 U8234 ( .A1(n7810), .A2(n7527), .ZN(n7809) );
  OR2_X1 U8235 ( .A1(n14505), .A2(n8218), .ZN(n8217) );
  NAND2_X1 U8236 ( .A1(n9142), .A2(n9141), .ZN(n14492) );
  NAND2_X1 U8237 ( .A1(n8219), .A2(n14505), .ZN(n14504) );
  NAND2_X1 U8238 ( .A1(n14559), .A2(n14551), .ZN(n7699) );
  NAND2_X1 U8239 ( .A1(n14680), .A2(n14165), .ZN(n7700) );
  NAND2_X1 U8240 ( .A1(n14562), .A2(n8934), .ZN(n14559) );
  NAND2_X1 U8241 ( .A1(n14566), .A2(n8214), .ZN(n14547) );
  NAND2_X1 U8242 ( .A1(n14564), .A2(n14563), .ZN(n14562) );
  NAND2_X1 U8243 ( .A1(n9128), .A2(n9127), .ZN(n12514) );
  OR2_X1 U8244 ( .A1(n8829), .A2(n8828), .ZN(n8870) );
  NAND2_X1 U8245 ( .A1(n12375), .A2(n8238), .ZN(n12433) );
  NAND2_X1 U8246 ( .A1(n12082), .A2(n8222), .ZN(n12284) );
  AND2_X1 U8247 ( .A1(n14303), .A2(n8799), .ZN(n8222) );
  OAI21_X1 U8248 ( .B1(n9122), .B2(n8208), .A(n8206), .ZN(n12275) );
  INV_X1 U8249 ( .A(n8207), .ZN(n8206) );
  OAI22_X1 U8250 ( .A1(n8208), .A2(n8209), .B1(n12090), .B2(n14354), .ZN(n8207) );
  NAND2_X1 U8251 ( .A1(n7542), .A2(n9123), .ZN(n8208) );
  AOI21_X1 U8252 ( .B1(n11941), .B2(n14301), .A(n7519), .ZN(n12083) );
  NAND2_X1 U8253 ( .A1(n11647), .A2(n14299), .ZN(n9122) );
  OR2_X1 U8254 ( .A1(n14073), .A2(n11639), .ZN(n11652) );
  OR2_X1 U8255 ( .A1(n8710), .A2(n8709), .ZN(n8731) );
  NAND2_X1 U8256 ( .A1(n8652), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8692) );
  NAND2_X1 U8257 ( .A1(n8225), .A2(n8642), .ZN(n7950) );
  NAND2_X1 U8258 ( .A1(n10364), .A2(n8225), .ZN(n7695) );
  NAND2_X1 U8259 ( .A1(n11166), .A2(n9116), .ZN(n11408) );
  NAND2_X1 U8260 ( .A1(n7951), .A2(n8227), .ZN(n8226) );
  INV_X1 U8261 ( .A(n10364), .ZN(n7951) );
  NAND2_X1 U8262 ( .A1(n8226), .A2(n8225), .ZN(n11162) );
  NAND2_X1 U8263 ( .A1(n10777), .A2(n7957), .ZN(n11169) );
  NOR2_X1 U8264 ( .A1(n10778), .A2(n14034), .ZN(n10777) );
  XNOR2_X1 U8265 ( .A(n14027), .B(n14364), .ZN(n14289) );
  OAI21_X1 U8266 ( .B1(n14287), .B2(n10819), .A(n7656), .ZN(n11351) );
  NAND2_X1 U8267 ( .A1(n7657), .A2(n14006), .ZN(n7656) );
  NAND2_X1 U8268 ( .A1(n11351), .A2(n8183), .ZN(n11350) );
  AND2_X1 U8269 ( .A1(n10487), .A2(n9149), .ZN(n14589) );
  NAND2_X1 U8270 ( .A1(n10786), .A2(n10743), .ZN(n10819) );
  INV_X1 U8271 ( .A(n9148), .ZN(n14606) );
  AND2_X1 U8272 ( .A1(n8539), .A2(n14276), .ZN(n10822) );
  NOR2_X1 U8273 ( .A1(n14458), .A2(n8241), .ZN(n8240) );
  INV_X1 U8274 ( .A(n9741), .ZN(n8241) );
  OR2_X1 U8275 ( .A1(n14461), .A2(n11636), .ZN(n8242) );
  OR2_X1 U8276 ( .A1(n14461), .A2(n10825), .ZN(n9739) );
  NAND2_X1 U8277 ( .A1(n8957), .A2(n8956), .ZN(n14675) );
  NAND2_X1 U8278 ( .A1(n8904), .A2(n8903), .ZN(n14596) );
  NAND2_X1 U8279 ( .A1(n8888), .A2(n8887), .ZN(n14698) );
  AND2_X1 U8280 ( .A1(n9190), .A2(n9189), .ZN(n10385) );
  XNOR2_X1 U8281 ( .A(n8560), .B(n8559), .ZN(n8563) );
  NAND2_X1 U8282 ( .A1(n14773), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8560) );
  AND2_X1 U8283 ( .A1(n8548), .A2(n8550), .ZN(n7953) );
  OAI21_X1 U8284 ( .B1(n11208), .B2(n9625), .A(n7638), .ZN(n11274) );
  NAND2_X1 U8285 ( .A1(n15326), .A2(n11755), .ZN(n7638) );
  OAI22_X1 U8286 ( .A1(n14830), .A2(n7639), .B1(n9625), .B2(n14863), .ZN(
        n11275) );
  OR2_X1 U8287 ( .A1(n8370), .A2(n8368), .ZN(n8366) );
  NAND2_X1 U8288 ( .A1(n8375), .A2(n8374), .ZN(n8373) );
  INV_X1 U8289 ( .A(n14977), .ZN(n8374) );
  INV_X1 U8290 ( .A(n14914), .ZN(n8368) );
  INV_X1 U8291 ( .A(n14854), .ZN(n8362) );
  NOR2_X1 U8292 ( .A1(n14879), .A2(n14878), .ZN(n8372) );
  OR2_X1 U8293 ( .A1(n15024), .A2(n15023), .ZN(n8390) );
  NAND2_X1 U8294 ( .A1(n7472), .A2(n14823), .ZN(n8381) );
  INV_X1 U8295 ( .A(n15023), .ZN(n8387) );
  INV_X1 U8296 ( .A(n12034), .ZN(n8394) );
  NAND2_X1 U8297 ( .A1(n11184), .A2(n11183), .ZN(n11194) );
  NAND2_X1 U8298 ( .A1(n15327), .A2(n11755), .ZN(n11184) );
  AND2_X1 U8299 ( .A1(n7645), .A2(n7571), .ZN(n12253) );
  INV_X1 U8300 ( .A(n14814), .ZN(n8382) );
  AOI22_X1 U8301 ( .A1(n15190), .A2(n15189), .B1(n15188), .B2(n15187), .ZN(
        n15229) );
  CLKBUF_X1 U8302 ( .A(n15195), .Z(n7778) );
  CLKBUF_X1 U8303 ( .A(n9282), .Z(n9634) );
  NOR2_X1 U8304 ( .A1(n11492), .A2(n11489), .ZN(n7796) );
  XNOR2_X1 U8305 ( .A(n7798), .B(n7797), .ZN(n15414) );
  INV_X1 U8306 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n7797) );
  NAND2_X1 U8307 ( .A1(n15908), .A2(n15411), .ZN(n7798) );
  NAND2_X1 U8308 ( .A1(n8407), .A2(n8414), .ZN(n8406) );
  INV_X1 U8309 ( .A(n8412), .ZN(n8407) );
  NOR2_X1 U8310 ( .A1(n7434), .A2(n8410), .ZN(n8409) );
  NAND2_X1 U8311 ( .A1(n8414), .A2(n8422), .ZN(n8410) );
  NAND2_X1 U8312 ( .A1(n7434), .A2(n8422), .ZN(n8417) );
  NOR2_X1 U8313 ( .A1(n15258), .A2(n8421), .ZN(n8418) );
  OR2_X1 U8314 ( .A1(n15470), .A2(n15659), .ZN(n15453) );
  NAND2_X1 U8315 ( .A1(n15668), .A2(n15018), .ZN(n7780) );
  OR2_X1 U8316 ( .A1(n7498), .A2(n8290), .ZN(n8289) );
  INV_X1 U8317 ( .A(n9673), .ZN(n8290) );
  INV_X1 U8318 ( .A(n8437), .ZN(n8436) );
  NAND2_X1 U8319 ( .A1(n7781), .A2(n8442), .ZN(n8439) );
  AND2_X1 U8320 ( .A1(n8433), .A2(n7503), .ZN(n8440) );
  OR2_X1 U8321 ( .A1(n15255), .A2(n8441), .ZN(n8433) );
  AND2_X1 U8322 ( .A1(n8106), .A2(n15146), .ZN(n8443) );
  NOR2_X1 U8323 ( .A1(n15565), .A2(n15694), .ZN(n15531) );
  INV_X1 U8324 ( .A(n15524), .ZN(n15528) );
  AND2_X1 U8325 ( .A1(n15580), .A2(n9668), .ZN(n8282) );
  INV_X1 U8326 ( .A(n8280), .ZN(n8279) );
  AOI21_X1 U8327 ( .B1(n8280), .B2(n8278), .A(n15252), .ZN(n8277) );
  INV_X1 U8328 ( .A(n8282), .ZN(n8278) );
  AND2_X1 U8329 ( .A1(n8447), .A2(n15252), .ZN(n8446) );
  OR2_X1 U8330 ( .A1(n8449), .A2(n8448), .ZN(n8447) );
  INV_X1 U8331 ( .A(n9542), .ZN(n8448) );
  NOR2_X1 U8332 ( .A1(n15559), .A2(n9666), .ZN(n8283) );
  NAND2_X1 U8333 ( .A1(n15571), .A2(n15580), .ZN(n8284) );
  NOR2_X1 U8334 ( .A1(n15613), .A2(n15710), .ZN(n15572) );
  NAND2_X1 U8335 ( .A1(n15630), .A2(n15629), .ZN(n15628) );
  NAND2_X1 U8336 ( .A1(n8298), .A2(n9657), .ZN(n8295) );
  AND2_X1 U8337 ( .A1(n15245), .A2(n9657), .ZN(n8296) );
  NAND2_X1 U8338 ( .A1(n11955), .A2(n15245), .ZN(n11954) );
  NAND2_X1 U8339 ( .A1(n7639), .A2(n9625), .ZN(n9643) );
  NOR2_X1 U8340 ( .A1(n15783), .A2(n9714), .ZN(n11977) );
  INV_X1 U8341 ( .A(n15427), .ZN(n15645) );
  NAND2_X1 U8342 ( .A1(n9691), .A2(n9716), .ZN(n10468) );
  XNOR2_X1 U8343 ( .A(n14230), .B(n14229), .ZN(n15207) );
  NAND2_X1 U8344 ( .A1(n8001), .A2(n8002), .ZN(n14230) );
  XNOR2_X1 U8345 ( .A(n9068), .B(n9052), .ZN(n14781) );
  NAND2_X1 U8346 ( .A1(n8030), .A2(n9049), .ZN(n9068) );
  NOR2_X1 U8347 ( .A1(n8397), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n8396) );
  NAND2_X1 U8348 ( .A1(n8011), .A2(n8955), .ZN(n8986) );
  NAND2_X1 U8349 ( .A1(n8953), .A2(n8952), .ZN(n8011) );
  XNOR2_X1 U8350 ( .A(n8804), .B(n8800), .ZN(n10782) );
  XNOR2_X1 U8351 ( .A(n8181), .B(n8609), .ZN(n10405) );
  NAND2_X1 U8352 ( .A1(n8595), .A2(n8424), .ZN(n8181) );
  NAND2_X1 U8353 ( .A1(n15970), .A2(n15969), .ZN(n15978) );
  AND2_X1 U8354 ( .A1(n7632), .A2(n7631), .ZN(n15992) );
  NAND2_X1 U8355 ( .A1(n15985), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7631) );
  AOI21_X1 U8356 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n16027), .A(n16026), .ZN(
        n16029) );
  NOR2_X1 U8357 ( .A1(n16025), .A2(n16024), .ZN(n16026) );
  AND2_X1 U8358 ( .A1(n8245), .A2(n8244), .ZN(n16048) );
  OAI21_X1 U8359 ( .B1(n16056), .B2(n16057), .A(n7634), .ZN(n7633) );
  INV_X1 U8360 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7634) );
  OAI21_X1 U8361 ( .B1(n12838), .B2(n7545), .A(n7862), .ZN(n7859) );
  AOI21_X1 U8362 ( .B1(n7864), .B2(n7867), .A(n7863), .ZN(n7862) );
  NAND2_X1 U8363 ( .A1(n12841), .A2(n7871), .ZN(n7870) );
  NOR2_X1 U8364 ( .A1(n7839), .A2(n12831), .ZN(n7838) );
  XNOR2_X1 U8365 ( .A(n12836), .B(n12984), .ZN(n12890) );
  NAND2_X1 U8366 ( .A1(n10184), .A2(n10183), .ZN(n13330) );
  NAND2_X1 U8367 ( .A1(n7836), .A2(n7834), .ZN(n12898) );
  AOI21_X1 U8368 ( .B1(n12970), .B2(n8510), .A(n7835), .ZN(n7834) );
  INV_X1 U8369 ( .A(n12899), .ZN(n7835) );
  OAI21_X1 U8370 ( .B1(n8489), .B2(n11513), .A(n8492), .ZN(n8493) );
  INV_X1 U8371 ( .A(n11298), .ZN(n8489) );
  NAND2_X1 U8372 ( .A1(n10168), .A2(n10167), .ZN(n13164) );
  NAND2_X1 U8373 ( .A1(n10105), .A2(n10104), .ZN(n13216) );
  NAND2_X1 U8374 ( .A1(n10141), .A2(n10140), .ZN(n13193) );
  NAND4_X1 U8375 ( .A1(n10018), .A2(n10017), .A3(n10016), .A4(n10015), .ZN(
        n12989) );
  INV_X1 U8376 ( .A(n12267), .ZN(n12991) );
  NAND4_X1 U8377 ( .A1(n9937), .A2(n9936), .A3(n9935), .A4(n9934), .ZN(n12640)
         );
  NAND4_X1 U8378 ( .A1(n9919), .A2(n9918), .A3(n9917), .A4(n9916), .ZN(n12992)
         );
  OR2_X1 U8379 ( .A1(n9817), .A2(n10999), .ZN(n9784) );
  XNOR2_X1 U8380 ( .A(n11245), .B(n11251), .ZN(n11022) );
  NAND2_X1 U8381 ( .A1(n8074), .A2(n7622), .ZN(n8073) );
  NAND2_X1 U8382 ( .A1(n8067), .A2(n8075), .ZN(n8066) );
  INV_X1 U8383 ( .A(n8071), .ZN(n8067) );
  NAND2_X1 U8384 ( .A1(n8074), .A2(n8068), .ZN(n8061) );
  OAI21_X1 U8385 ( .B1(n13068), .B2(n16274), .A(n8045), .ZN(n8044) );
  NOR2_X1 U8386 ( .A1(n13067), .A2(n13066), .ZN(n8045) );
  OAI21_X1 U8387 ( .B1(n10276), .B2(n16349), .A(n10275), .ZN(n13101) );
  NOR2_X1 U8388 ( .A1(n10274), .A2(n10273), .ZN(n10275) );
  AND2_X1 U8389 ( .A1(n9984), .A2(n9983), .ZN(n12412) );
  AND3_X1 U8390 ( .A1(n9962), .A2(n9961), .A3(n9960), .ZN(n12272) );
  AND3_X1 U8391 ( .A1(n9832), .A2(n9831), .A3(n9830), .ZN(n11597) );
  OR2_X1 U8392 ( .A1(n16601), .A2(n13321), .ZN(n7752) );
  AND3_X1 U8393 ( .A1(n9889), .A2(n9888), .A3(n9887), .ZN(n11859) );
  AND3_X1 U8394 ( .A1(n9853), .A2(n9852), .A3(n9851), .ZN(n11703) );
  NOR2_X1 U8395 ( .A1(n11441), .A2(n10341), .ZN(n16568) );
  INV_X1 U8396 ( .A(n13318), .ZN(n13320) );
  NAND2_X1 U8397 ( .A1(n10060), .A2(n10059), .ZN(n13824) );
  NAND2_X1 U8398 ( .A1(n10029), .A2(n10028), .ZN(n13832) );
  OR2_X1 U8399 ( .A1(n16605), .A2(n16593), .ZN(n13837) );
  INV_X1 U8400 ( .A(n14361), .ZN(n11311) );
  OAI211_X1 U8401 ( .C1(n7672), .C2(n13860), .A(n7669), .B(n7670), .ZN(n13886)
         );
  NAND2_X1 U8402 ( .A1(n13859), .A2(n7671), .ZN(n7670) );
  NAND2_X1 U8403 ( .A1(n7673), .A2(n13861), .ZN(n7672) );
  NAND2_X1 U8404 ( .A1(n13886), .A2(n7774), .ZN(n13885) );
  NOR2_X1 U8405 ( .A1(n14177), .A2(n14430), .ZN(n7774) );
  NAND2_X1 U8406 ( .A1(n11319), .A2(n11145), .ZN(n8153) );
  NAND2_X1 U8407 ( .A1(n8154), .A2(n11219), .ZN(n11319) );
  AND2_X1 U8408 ( .A1(n11314), .A2(n11142), .ZN(n8154) );
  INV_X1 U8409 ( .A(n13949), .ZN(n7679) );
  AND2_X1 U8410 ( .A1(n13925), .A2(n7677), .ZN(n7676) );
  NAND2_X1 U8411 ( .A1(n7678), .A2(n13949), .ZN(n7677) );
  NAND2_X1 U8412 ( .A1(n9020), .A2(n9019), .ZN(n14497) );
  NOR2_X2 U8413 ( .A1(n12390), .A2(n7977), .ZN(n12427) );
  OR2_X1 U8414 ( .A1(n12314), .A2(n12313), .ZN(n7977) );
  INV_X1 U8415 ( .A(n13994), .ZN(n10786) );
  NAND2_X1 U8416 ( .A1(n8923), .A2(n8922), .ZN(n14688) );
  OAI21_X1 U8417 ( .B1(n13981), .B2(n13963), .A(n7980), .ZN(n7979) );
  INV_X1 U8418 ( .A(n13989), .ZN(n7980) );
  AOI21_X1 U8419 ( .B1(n13931), .B2(n13869), .A(n13932), .ZN(n13930) );
  INV_X1 U8420 ( .A(n14286), .ZN(n14323) );
  NAND2_X1 U8421 ( .A1(n9063), .A2(n9062), .ZN(n14342) );
  NAND2_X1 U8422 ( .A1(n8578), .A2(n7509), .ZN(n14365) );
  OR2_X1 U8423 ( .A1(n8831), .A2(n11353), .ZN(n8579) );
  NAND2_X1 U8424 ( .A1(n7946), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8567) );
  OR2_X1 U8425 ( .A1(n14218), .A2(n8564), .ZN(n8565) );
  NAND2_X1 U8426 ( .A1(n14653), .A2(n14652), .ZN(n14737) );
  OR2_X1 U8427 ( .A1(n14649), .A2(n16386), .ZN(n14653) );
  NAND2_X1 U8428 ( .A1(n7955), .A2(n7954), .ZN(n8204) );
  NOR2_X1 U8429 ( .A1(n14443), .A2(n14449), .ZN(n7954) );
  NAND2_X1 U8430 ( .A1(n9078), .A2(n9077), .ZN(n14193) );
  NAND2_X1 U8431 ( .A1(n7644), .A2(n7522), .ZN(n16609) );
  INV_X1 U8432 ( .A(n16606), .ZN(n7643) );
  NAND2_X1 U8433 ( .A1(n14993), .A2(n14867), .ZN(n14898) );
  AOI22_X1 U8434 ( .A1(n15004), .A2(n15005), .B1(n14839), .B2(n14838), .ZN(
        n14904) );
  NAND2_X1 U8435 ( .A1(n9515), .A2(n9514), .ZN(n15703) );
  NAND2_X1 U8436 ( .A1(n9413), .A2(n9412), .ZN(n15101) );
  NAND2_X1 U8437 ( .A1(n14786), .A2(n15206), .ZN(n9570) );
  NAND2_X1 U8438 ( .A1(n11263), .A2(n15206), .ZN(n9461) );
  NOR2_X1 U8439 ( .A1(n10925), .A2(n10924), .ZN(n10923) );
  NAND2_X1 U8440 ( .A1(n9226), .A2(n9225), .ZN(n15675) );
  NAND2_X1 U8441 ( .A1(n9511), .A2(n9510), .ZN(n8347) );
  NOR2_X1 U8442 ( .A1(n15973), .A2(n15974), .ZN(n15983) );
  NAND2_X1 U8443 ( .A1(n16004), .A2(n16005), .ZN(n16016) );
  INV_X1 U8444 ( .A(n7629), .ZN(n16042) );
  OR2_X1 U8445 ( .A1(n16042), .A2(n16043), .ZN(n8244) );
  XNOR2_X1 U8446 ( .A(n16048), .B(n8243), .ZN(n16046) );
  INV_X1 U8447 ( .A(n16047), .ZN(n8243) );
  NAND2_X1 U8448 ( .A1(n16046), .A2(n16045), .ZN(n16049) );
  NOR2_X1 U8449 ( .A1(n7499), .A2(n16063), .ZN(n16064) );
  NOR2_X1 U8450 ( .A1(n16095), .A2(n16094), .ZN(n16098) );
  NAND2_X1 U8451 ( .A1(n16381), .A2(n14013), .ZN(n14011) );
  AOI21_X1 U8452 ( .B1(n15065), .B2(n7639), .A(n9625), .ZN(n15054) );
  NAND2_X1 U8453 ( .A1(n14044), .A2(n7510), .ZN(n8335) );
  NOR2_X1 U8454 ( .A1(n14044), .A2(n7510), .ZN(n8336) );
  OAI22_X1 U8455 ( .A1(n8454), .A2(n8453), .B1(n15063), .B2(n8452), .ZN(n15068) );
  INV_X1 U8456 ( .A(n15062), .ZN(n8452) );
  NOR2_X1 U8457 ( .A1(n15064), .A2(n15062), .ZN(n8453) );
  INV_X1 U8458 ( .A(n15075), .ZN(n8474) );
  NOR2_X1 U8459 ( .A1(n8333), .A2(n8332), .ZN(n8331) );
  AOI21_X1 U8460 ( .B1(n8472), .B2(n8470), .A(n8469), .ZN(n8468) );
  INV_X1 U8461 ( .A(n15102), .ZN(n7895) );
  NAND2_X1 U8462 ( .A1(n8318), .A2(n8317), .ZN(n14110) );
  AOI21_X1 U8463 ( .B1(n8322), .B2(n8324), .A(n7537), .ZN(n8317) );
  NAND2_X1 U8464 ( .A1(n15106), .A2(n15108), .ZN(n8461) );
  NAND2_X1 U8465 ( .A1(n14119), .A2(n7482), .ZN(n8341) );
  AOI21_X1 U8466 ( .B1(n8466), .B2(n8465), .A(n8464), .ZN(n8463) );
  NAND2_X1 U8467 ( .A1(n15137), .A2(n15135), .ZN(n8475) );
  NAND2_X1 U8468 ( .A1(n14174), .A2(n14175), .ZN(n8313) );
  OAI22_X1 U8469 ( .A1(n15165), .A2(n7897), .B1(n15166), .B2(n7896), .ZN(
        n15170) );
  NOR2_X1 U8470 ( .A1(n15167), .A2(n15164), .ZN(n7897) );
  INV_X1 U8471 ( .A(n15164), .ZN(n7896) );
  NOR2_X1 U8472 ( .A1(n14191), .A2(n8308), .ZN(n8307) );
  INV_X1 U8473 ( .A(n8313), .ZN(n8308) );
  NAND2_X1 U8474 ( .A1(n14164), .A2(n7601), .ZN(n8339) );
  NAND2_X1 U8475 ( .A1(n8316), .A2(n8315), .ZN(n8314) );
  INV_X1 U8476 ( .A(n14175), .ZN(n8315) );
  INV_X1 U8477 ( .A(n14174), .ZN(n8316) );
  NAND2_X1 U8478 ( .A1(n8305), .A2(n8307), .ZN(n8304) );
  INV_X1 U8479 ( .A(n8314), .ZN(n8305) );
  NOR2_X1 U8480 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7650) );
  INV_X1 U8481 ( .A(n8013), .ZN(n8012) );
  OAI21_X1 U8482 ( .B1(n8952), .B2(n8014), .A(n8985), .ZN(n8013) );
  INV_X1 U8483 ( .A(SI_1_), .ZN(n13650) );
  INV_X1 U8484 ( .A(n9975), .ZN(n7736) );
  AND2_X1 U8485 ( .A1(n8188), .A2(n14462), .ZN(n8186) );
  NAND2_X1 U8486 ( .A1(n8193), .A2(n8190), .ZN(n8189) );
  INV_X1 U8487 ( .A(n7596), .ZN(n8190) );
  NOR2_X1 U8488 ( .A1(n14671), .A2(n7965), .ZN(n7964) );
  INV_X1 U8489 ( .A(n7966), .ZN(n7965) );
  INV_X1 U8490 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8526) );
  INV_X1 U8491 ( .A(n9049), .ZN(n8033) );
  INV_X1 U8492 ( .A(n8920), .ZN(n7987) );
  AOI21_X1 U8493 ( .B1(n8019), .B2(n8022), .A(n8877), .ZN(n8018) );
  NOR2_X1 U8494 ( .A1(n8803), .A2(n8027), .ZN(n8026) );
  INV_X1 U8495 ( .A(n8785), .ZN(n8027) );
  INV_X1 U8496 ( .A(n8800), .ZN(n8803) );
  NOR2_X1 U8497 ( .A1(n8661), .A2(n8643), .ZN(n8427) );
  NAND2_X1 U8498 ( .A1(n7759), .A2(n7758), .ZN(n8625) );
  OR2_X1 U8499 ( .A1(n8156), .A2(n7760), .ZN(n7759) );
  NAND2_X1 U8500 ( .A1(n8156), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7758) );
  INV_X1 U8501 ( .A(n12017), .ZN(n7831) );
  AND2_X1 U8502 ( .A1(n8269), .A2(n8268), .ZN(n8267) );
  NOR2_X1 U8503 ( .A1(n13145), .A2(n12585), .ZN(n8269) );
  INV_X1 U8504 ( .A(n13132), .ZN(n8268) );
  NOR2_X1 U8505 ( .A1(n7808), .A2(n12761), .ZN(n7807) );
  OR2_X1 U8506 ( .A1(n16272), .A2(n7625), .ZN(n8088) );
  OR2_X1 U8507 ( .A1(n7488), .A2(n13024), .ZN(n8089) );
  NAND2_X1 U8508 ( .A1(n12581), .A2(n12582), .ZN(n7761) );
  INV_X1 U8509 ( .A(n10113), .ZN(n7934) );
  OR2_X1 U8510 ( .A1(n13193), .A2(n12867), .ZN(n12587) );
  OR2_X1 U8511 ( .A1(n13832), .A2(n12903), .ZN(n12670) );
  OR2_X1 U8512 ( .A1(n10013), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n10031) );
  OAI21_X1 U8513 ( .B1(n9872), .B2(n7908), .A(n12737), .ZN(n7907) );
  INV_X1 U8514 ( .A(n12616), .ZN(n8130) );
  NOR2_X1 U8515 ( .A1(n8129), .A2(n8130), .ZN(n8128) );
  INV_X1 U8516 ( .A(n12612), .ZN(n8129) );
  INV_X1 U8517 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n13475) );
  NAND2_X1 U8518 ( .A1(n16363), .A2(n9794), .ZN(n12599) );
  NAND2_X1 U8519 ( .A1(n9770), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9774) );
  NAND2_X1 U8520 ( .A1(n9754), .A2(n8152), .ZN(n8151) );
  INV_X1 U8521 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n9754) );
  INV_X1 U8522 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8152) );
  OAI21_X1 U8523 ( .B1(n7713), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n7710), .ZN(
        n7709) );
  NAND2_X1 U8524 ( .A1(n10165), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7710) );
  NOR2_X1 U8525 ( .A1(n7714), .A2(n7621), .ZN(n7713) );
  INV_X1 U8526 ( .A(n7716), .ZN(n7714) );
  INV_X1 U8527 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n9751) );
  INV_X1 U8528 ( .A(n7856), .ZN(n7851) );
  NOR2_X1 U8529 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n7878) );
  NAND2_X1 U8530 ( .A1(n7728), .A2(n7727), .ZN(n10115) );
  AOI21_X1 U8531 ( .B1(n7730), .B2(n7732), .A(n7616), .ZN(n7727) );
  INV_X1 U8532 ( .A(n8256), .ZN(n8255) );
  OAI21_X1 U8533 ( .B1(n10055), .B2(n8257), .A(n10069), .ZN(n8256) );
  INV_X1 U8534 ( .A(n10057), .ZN(n8257) );
  AND4_X1 U8535 ( .A1(n7853), .A2(n7858), .A3(n9747), .A4(n7943), .ZN(n7852)
         );
  AND2_X1 U8536 ( .A1(n7592), .A2(n9748), .ZN(n7853) );
  INV_X1 U8537 ( .A(n10024), .ZN(n7745) );
  INV_X1 U8538 ( .A(n7744), .ZN(n7743) );
  OAI21_X1 U8539 ( .B1(n10021), .B2(n7745), .A(n10039), .ZN(n7744) );
  NAND2_X1 U8540 ( .A1(n7735), .A2(n7733), .ZN(n10005) );
  INV_X1 U8541 ( .A(n7734), .ZN(n7733) );
  OR2_X1 U8542 ( .A1(n7791), .A2(n7594), .ZN(n7735) );
  OAI21_X1 U8543 ( .B1(n7738), .B2(n7594), .A(n9987), .ZN(n7734) );
  INV_X1 U8544 ( .A(n8265), .ZN(n8260) );
  INV_X1 U8545 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9920) );
  INV_X1 U8546 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9885) );
  AND2_X1 U8547 ( .A1(n8502), .A2(n9849), .ZN(n7943) );
  INV_X1 U8548 ( .A(n9864), .ZN(n7720) );
  OR2_X1 U8549 ( .A1(n13953), .A2(n12545), .ZN(n12544) );
  NAND2_X1 U8550 ( .A1(n7470), .A2(n8303), .ZN(n8301) );
  INV_X1 U8551 ( .A(n14318), .ZN(n14249) );
  INV_X1 U8552 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8823) );
  NAND2_X1 U8553 ( .A1(n7547), .A2(n14740), .ZN(n7958) );
  AND2_X1 U8554 ( .A1(n9055), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9079) );
  INV_X1 U8555 ( .A(n9030), .ZN(n7693) );
  INV_X1 U8556 ( .A(n9045), .ZN(n8224) );
  INV_X1 U8557 ( .A(n7949), .ZN(n7948) );
  OAI21_X1 U8558 ( .B1(n7467), .B2(n8966), .A(n8982), .ZN(n7949) );
  INV_X1 U8559 ( .A(n9135), .ZN(n8213) );
  OR2_X1 U8560 ( .A1(n8214), .A2(n8213), .ZN(n8212) );
  NOR2_X1 U8561 ( .A1(n14675), .A2(n14681), .ZN(n7966) );
  NOR2_X1 U8562 ( .A1(n12519), .A2(n14763), .ZN(n12520) );
  OR2_X1 U8563 ( .A1(n8778), .A2(n8777), .ZN(n8792) );
  NOR2_X1 U8564 ( .A1(n14301), .A2(n8210), .ZN(n8209) );
  INV_X1 U8565 ( .A(n9121), .ZN(n8210) );
  NOR2_X1 U8566 ( .A1(n14047), .A2(n14055), .ZN(n7962) );
  OR2_X1 U8567 ( .A1(n14492), .A2(n8189), .ZN(n8187) );
  OR2_X1 U8568 ( .A1(n8191), .A2(n9144), .ZN(n8188) );
  AND2_X1 U8569 ( .A1(n14313), .A2(n8192), .ZN(n8191) );
  OR2_X1 U8570 ( .A1(n14310), .A2(n7596), .ZN(n8192) );
  OR2_X1 U8571 ( .A1(n14509), .A2(n14497), .ZN(n14495) );
  NAND2_X1 U8572 ( .A1(n14572), .A2(n7964), .ZN(n14524) );
  INV_X1 U8573 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U8574 ( .A1(n9160), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9165) );
  NAND2_X1 U8575 ( .A1(n8528), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8886) );
  OR2_X1 U8576 ( .A1(n8705), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8706) );
  OR2_X1 U8577 ( .A1(n8647), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n8665) );
  OR2_X1 U8578 ( .A1(n14891), .A2(n14890), .ZN(n8379) );
  NOR2_X1 U8579 ( .A1(n9417), .A2(n9416), .ZN(n9415) );
  NOR2_X1 U8580 ( .A1(n9464), .A2(n11498), .ZN(n9463) );
  AOI21_X1 U8581 ( .B1(n7469), .B2(n7515), .A(n7462), .ZN(n7885) );
  OR2_X1 U8582 ( .A1(n15193), .A2(n8113), .ZN(n8112) );
  NAND2_X1 U8583 ( .A1(n8114), .A2(n15460), .ZN(n8113) );
  NOR2_X1 U8584 ( .A1(n8104), .A2(n15675), .ZN(n8103) );
  INV_X1 U8585 ( .A(n8105), .ZN(n8104) );
  INV_X1 U8586 ( .A(n8443), .ZN(n8441) );
  AND2_X1 U8587 ( .A1(n15559), .A2(n9529), .ZN(n8449) );
  NOR2_X1 U8588 ( .A1(n15631), .A2(n15725), .ZN(n8099) );
  NOR2_X1 U8589 ( .A1(n9309), .A2(n9308), .ZN(n9307) );
  INV_X1 U8590 ( .A(n15322), .ZN(n11768) );
  OR2_X1 U8591 ( .A1(n15326), .A2(n9625), .ZN(n15042) );
  INV_X1 U8592 ( .A(n15038), .ZN(n11575) );
  AND2_X1 U8593 ( .A1(n11174), .A2(n11173), .ZN(n11568) );
  NAND2_X1 U8594 ( .A1(n8101), .A2(n8100), .ZN(n15631) );
  AOI21_X1 U8595 ( .B1(n7464), .B2(n8007), .A(n7624), .ZN(n8002) );
  AOI21_X1 U8596 ( .B1(n9095), .B2(n8006), .A(n8005), .ZN(n8004) );
  INV_X1 U8597 ( .A(n14223), .ZN(n8005) );
  INV_X1 U8598 ( .A(n9090), .ZN(n8006) );
  INV_X1 U8599 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9194) );
  NOR2_X1 U8600 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n7641) );
  NOR2_X1 U8601 ( .A1(n9050), .A2(n8035), .ZN(n8034) );
  INV_X1 U8602 ( .A(n9031), .ZN(n8035) );
  NOR2_X1 U8603 ( .A1(n9200), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n8458) );
  NAND2_X1 U8604 ( .A1(n9615), .A2(n8398), .ZN(n8397) );
  INV_X1 U8605 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8398) );
  INV_X1 U8606 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8346) );
  NAND2_X1 U8607 ( .A1(n8768), .A2(n13436), .ZN(n8785) );
  NOR2_X1 U8608 ( .A1(n8749), .A2(n8445), .ZN(n8444) );
  INV_X1 U8609 ( .A(n8744), .ZN(n8445) );
  XNOR2_X1 U8610 ( .A(n8743), .B(SI_10_), .ZN(n8740) );
  OR2_X1 U8611 ( .A1(n9364), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9381) );
  NAND2_X1 U8612 ( .A1(n7996), .A2(n7998), .ZN(n8723) );
  AND2_X1 U8613 ( .A1(n7995), .A2(n7993), .ZN(n7998) );
  NAND2_X1 U8614 ( .A1(n7994), .A2(SI_9_), .ZN(n7993) );
  OAI21_X1 U8615 ( .B1(n8623), .B2(n8233), .A(n8644), .ZN(n8232) );
  INV_X1 U8616 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n7890) );
  XNOR2_X1 U8617 ( .A(n8625), .B(SI_4_), .ZN(n8622) );
  NAND2_X1 U8618 ( .A1(n8425), .A2(n8592), .ZN(n7983) );
  NOR2_X1 U8619 ( .A1(n8609), .A2(n8590), .ZN(n8425) );
  OAI21_X1 U8620 ( .B1(n10419), .B2(P1_DATAO_REG_1__SCAN_IN), .A(n7991), .ZN(
        n8275) );
  NAND2_X1 U8621 ( .A1(n10419), .A2(n10414), .ZN(n7991) );
  XNOR2_X1 U8622 ( .A(n15949), .B(n15941), .ZN(n15951) );
  NAND2_X1 U8623 ( .A1(n15958), .A2(n15959), .ZN(n15967) );
  XNOR2_X1 U8624 ( .A(n15967), .B(n15960), .ZN(n15968) );
  NAND2_X1 U8625 ( .A1(n15999), .A2(n15998), .ZN(n16006) );
  INV_X1 U8626 ( .A(n11620), .ZN(n7832) );
  OR2_X1 U8627 ( .A1(n12622), .A2(n11686), .ZN(n11687) );
  INV_X1 U8628 ( .A(n12963), .ZN(n8499) );
  AOI21_X1 U8629 ( .B1(n12963), .B2(n8498), .A(n7504), .ZN(n8497) );
  INV_X1 U8630 ( .A(n12837), .ZN(n8498) );
  XNOR2_X1 U8631 ( .A(n12840), .B(n8270), .ZN(n12848) );
  INV_X1 U8632 ( .A(n7874), .ZN(n7871) );
  NAND2_X1 U8633 ( .A1(n7868), .A2(n7872), .ZN(n7867) );
  OR2_X1 U8634 ( .A1(n12841), .A2(n7871), .ZN(n7868) );
  AND2_X1 U8635 ( .A1(n7866), .A2(n7876), .ZN(n7864) );
  NAND2_X1 U8636 ( .A1(n7873), .A2(n7869), .ZN(n7866) );
  NAND2_X1 U8637 ( .A1(n7471), .A2(n7839), .ZN(n7837) );
  NAND2_X1 U8638 ( .A1(n10030), .A2(n13702), .ZN(n10045) );
  INV_X1 U8639 ( .A(n10031), .ZN(n10030) );
  AOI21_X1 U8640 ( .B1(n11512), .B2(n11297), .A(n11515), .ZN(n8492) );
  OR2_X1 U8641 ( .A1(n10045), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n10062) );
  INV_X1 U8642 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n11106) );
  INV_X1 U8643 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n13489) );
  NAND2_X1 U8644 ( .A1(n12876), .A2(n7494), .ZN(n12922) );
  OR2_X1 U8645 ( .A1(n10106), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n10123) );
  NAND2_X1 U8646 ( .A1(n10091), .A2(n13469), .ZN(n10106) );
  INV_X1 U8647 ( .A(n10092), .ZN(n10091) );
  NAND2_X1 U8648 ( .A1(n7823), .A2(n7822), .ZN(n12825) );
  NAND2_X1 U8649 ( .A1(n7481), .A2(n7826), .ZN(n7822) );
  OR2_X1 U8650 ( .A1(n12876), .A2(n7824), .ZN(n7823) );
  NOR2_X1 U8651 ( .A1(n12997), .A2(n10950), .ZN(n10977) );
  OR2_X1 U8652 ( .A1(n10075), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n10092) );
  NAND2_X1 U8653 ( .A1(n10061), .A2(n13680), .ZN(n10075) );
  INV_X1 U8654 ( .A(n10062), .ZN(n10061) );
  OR2_X1 U8655 ( .A1(n12803), .A2(n12989), .ZN(n12804) );
  INV_X1 U8656 ( .A(n10297), .ZN(n12767) );
  AOI21_X1 U8657 ( .B1(n13148), .B2(n10247), .A(n10191), .ZN(n12915) );
  AND2_X1 U8658 ( .A1(n10177), .A2(n10176), .ZN(n12891) );
  OR2_X1 U8659 ( .A1(n11114), .A2(n10991), .ZN(n11116) );
  NAND2_X1 U8660 ( .A1(n8092), .A2(n8091), .ZN(n11050) );
  NAND2_X1 U8661 ( .A1(n11026), .A2(n10998), .ZN(n8091) );
  NAND2_X1 U8662 ( .A1(n7779), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8092) );
  AND2_X1 U8663 ( .A1(n11021), .A2(n11046), .ZN(n11044) );
  XNOR2_X1 U8664 ( .A(n11044), .B(n11028), .ZN(n16115) );
  NAND2_X1 U8665 ( .A1(n7768), .A2(n7767), .ZN(n7766) );
  INV_X1 U8666 ( .A(n11029), .ZN(n7768) );
  NAND2_X1 U8667 ( .A1(n8501), .A2(n9746), .ZN(n9826) );
  INV_X1 U8668 ( .A(n9801), .ZN(n8501) );
  INV_X1 U8669 ( .A(n8087), .ZN(n16116) );
  NAND2_X1 U8670 ( .A1(n8042), .A2(n8041), .ZN(n11100) );
  OR2_X1 U8671 ( .A1(n11044), .A2(n7767), .ZN(n8041) );
  NAND2_X1 U8672 ( .A1(n16115), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8042) );
  NAND2_X1 U8673 ( .A1(n8055), .A2(n8054), .ZN(n16120) );
  OAI211_X1 U8674 ( .C1(n11056), .C2(n8053), .A(n8056), .B(n8052), .ZN(n8055)
         );
  NAND2_X1 U8675 ( .A1(n10997), .A2(n16122), .ZN(n8052) );
  NAND2_X1 U8676 ( .A1(n9746), .A2(n8502), .ZN(n8500) );
  INV_X1 U8677 ( .A(n7748), .ZN(n11533) );
  NAND2_X1 U8678 ( .A1(n11659), .A2(n7520), .ZN(n11830) );
  XNOR2_X1 U8679 ( .A(n13051), .B(n16187), .ZN(n16192) );
  AND2_X1 U8680 ( .A1(n16171), .A2(n13032), .ZN(n16190) );
  NOR2_X1 U8681 ( .A1(n16197), .A2(n13018), .ZN(n16216) );
  NAND2_X1 U8682 ( .A1(n16168), .A2(n13050), .ZN(n13051) );
  NAND2_X1 U8683 ( .A1(n8086), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8084) );
  NAND2_X1 U8684 ( .A1(n13022), .A2(n8086), .ZN(n8085) );
  INV_X1 U8685 ( .A(n16252), .ZN(n8086) );
  NOR2_X1 U8686 ( .A1(n16235), .A2(n16234), .ZN(n16233) );
  NAND2_X1 U8687 ( .A1(n13054), .A2(n13306), .ZN(n7785) );
  OAI21_X1 U8688 ( .B1(n13054), .B2(n13306), .A(n7787), .ZN(n7786) );
  AND2_X1 U8689 ( .A1(n8058), .A2(n8057), .ZN(n16265) );
  NAND2_X1 U8690 ( .A1(n13038), .A2(n13058), .ZN(n8057) );
  NAND2_X1 U8691 ( .A1(n8088), .A2(n8089), .ZN(n13070) );
  INV_X1 U8692 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n13084) );
  NAND3_X1 U8693 ( .A1(n8088), .A2(n8089), .A3(n13069), .ZN(n7816) );
  INV_X1 U8694 ( .A(n13079), .ZN(n7815) );
  INV_X1 U8695 ( .A(n8144), .ZN(n8143) );
  AOI21_X1 U8696 ( .B1(n8144), .B2(n13119), .A(n10296), .ZN(n8142) );
  NAND2_X1 U8697 ( .A1(n7911), .A2(n7909), .ZN(n10253) );
  NAND2_X1 U8698 ( .A1(n7910), .A2(n7915), .ZN(n7909) );
  INV_X1 U8699 ( .A(n7761), .ZN(n12762) );
  NAND2_X1 U8700 ( .A1(n13120), .A2(n10226), .ZN(n13105) );
  NAND2_X1 U8701 ( .A1(n10215), .A2(n13461), .ZN(n10234) );
  INV_X1 U8702 ( .A(n10216), .ZN(n10215) );
  OAI21_X1 U8703 ( .B1(n13153), .B2(n7937), .A(n7939), .ZN(n10208) );
  NAND2_X1 U8704 ( .A1(n10192), .A2(n7938), .ZN(n7937) );
  OR2_X1 U8705 ( .A1(n10199), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n10216) );
  NAND2_X1 U8706 ( .A1(n10170), .A2(n10169), .ZN(n10186) );
  INV_X1 U8707 ( .A(n10171), .ZN(n10170) );
  NAND2_X1 U8708 ( .A1(n10185), .A2(n13675), .ZN(n10199) );
  INV_X1 U8709 ( .A(n10186), .ZN(n10185) );
  AND2_X1 U8710 ( .A1(n12711), .A2(n12710), .ZN(n13142) );
  OR2_X1 U8711 ( .A1(n12585), .A2(n13158), .ZN(n13159) );
  AND2_X1 U8712 ( .A1(n8520), .A2(n12588), .ZN(n8131) );
  AND2_X1 U8713 ( .A1(n10294), .A2(n12709), .ZN(n13162) );
  NAND2_X1 U8714 ( .A1(n13158), .A2(n12706), .ZN(n13176) );
  NAND2_X1 U8715 ( .A1(n12587), .A2(n12588), .ZN(n13185) );
  AND3_X1 U8716 ( .A1(n10127), .A2(n10126), .A3(n10125), .ZN(n13187) );
  AND2_X1 U8717 ( .A1(n10290), .A2(n13250), .ZN(n8137) );
  NAND2_X1 U8718 ( .A1(n8135), .A2(n12736), .ZN(n8134) );
  NAND2_X1 U8719 ( .A1(n8136), .A2(n10290), .ZN(n8135) );
  AND4_X1 U8720 ( .A1(n10112), .A2(n10111), .A3(n10110), .A4(n10109), .ZN(
        n13227) );
  AOI21_X1 U8721 ( .B1(n7922), .B2(n13250), .A(n7920), .ZN(n7919) );
  INV_X1 U8722 ( .A(n12679), .ZN(n7920) );
  AND4_X1 U8723 ( .A1(n10050), .A2(n10049), .A3(n10048), .A4(n10047), .ZN(
        n13254) );
  INV_X1 U8724 ( .A(n13297), .ZN(n13301) );
  NAND2_X1 U8725 ( .A1(n9966), .A2(n9965), .ZN(n9995) );
  INV_X1 U8726 ( .A(n9967), .ZN(n9966) );
  AND2_X1 U8727 ( .A1(n12652), .A2(n12653), .ZN(n12750) );
  INV_X1 U8728 ( .A(n7926), .ZN(n7925) );
  OAI21_X1 U8729 ( .B1(n7930), .B2(n7927), .A(n9964), .ZN(n7926) );
  OR2_X1 U8730 ( .A1(n9945), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9967) );
  NAND2_X1 U8731 ( .A1(n9912), .A2(n13489), .ZN(n9932) );
  INV_X1 U8732 ( .A(n9913), .ZN(n9912) );
  OR2_X1 U8733 ( .A1(n9932), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9945) );
  AND2_X1 U8734 ( .A1(n12631), .A2(n12632), .ZN(n12629) );
  INV_X1 U8735 ( .A(n12629), .ZN(n12744) );
  INV_X1 U8736 ( .A(n16352), .ZN(n13251) );
  NAND2_X1 U8737 ( .A1(n11924), .A2(n9873), .ZN(n11847) );
  AND2_X1 U8738 ( .A1(n12626), .A2(n12627), .ZN(n12624) );
  NAND2_X1 U8739 ( .A1(n11696), .A2(n9872), .ZN(n11924) );
  OR2_X1 U8740 ( .A1(n9854), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9875) );
  INV_X1 U8741 ( .A(n12995), .ZN(n12622) );
  NAND2_X1 U8742 ( .A1(n13475), .A2(n11106), .ZN(n9837) );
  NAND2_X1 U8743 ( .A1(n9836), .A2(n13679), .ZN(n9854) );
  INV_X1 U8744 ( .A(n9837), .ZN(n9836) );
  NAND2_X1 U8745 ( .A1(n11590), .A2(n12612), .ZN(n11695) );
  NAND2_X1 U8746 ( .A1(n11695), .A2(n12746), .ZN(n11917) );
  AND2_X1 U8747 ( .A1(n12612), .A2(n12613), .ZN(n12610) );
  NOR2_X1 U8748 ( .A1(n12740), .A2(n11733), .ZN(n9811) );
  AND3_X1 U8749 ( .A1(n9793), .A2(n9792), .A3(n9791), .ZN(n10976) );
  OR2_X1 U8750 ( .A1(n9800), .A2(n10433), .ZN(n9792) );
  OR2_X1 U8751 ( .A1(n12569), .A2(SI_2_), .ZN(n9793) );
  NAND2_X1 U8752 ( .A1(n12599), .A2(n12600), .ZN(n10277) );
  INV_X1 U8753 ( .A(n10277), .ZN(n10281) );
  INV_X1 U8754 ( .A(n12739), .ZN(n16312) );
  INV_X1 U8755 ( .A(n16311), .ZN(n9779) );
  OR2_X1 U8756 ( .A1(n10335), .A2(n10334), .ZN(n11441) );
  INV_X1 U8757 ( .A(n12412), .ZN(n16583) );
  INV_X1 U8758 ( .A(n16597), .ZN(n16414) );
  NAND2_X1 U8759 ( .A1(n8149), .A2(n9757), .ZN(n8148) );
  AND2_X1 U8760 ( .A1(n10311), .A2(n10310), .ZN(n10332) );
  OAI21_X1 U8761 ( .B1(n10166), .B2(n7711), .A(n7708), .ZN(n10194) );
  NAND2_X1 U8762 ( .A1(n7715), .A2(n10180), .ZN(n7711) );
  NAND2_X1 U8763 ( .A1(n10166), .A2(n7709), .ZN(n7708) );
  NAND2_X1 U8764 ( .A1(n7716), .A2(n12191), .ZN(n7715) );
  NAND2_X1 U8765 ( .A1(n10195), .A2(n10182), .ZN(n10193) );
  XNOR2_X1 U8766 ( .A(n10115), .B(n11707), .ZN(n10114) );
  OR2_X1 U8767 ( .A1(n10008), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n10025) );
  AND2_X1 U8768 ( .A1(n9977), .A2(n9976), .ZN(n9981) );
  NOR2_X1 U8769 ( .A1(n9922), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n9958) );
  XNOR2_X1 U8770 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n9939) );
  OAI21_X1 U8771 ( .B1(n9883), .B2(n8261), .A(n8258), .ZN(n9941) );
  INV_X1 U8772 ( .A(n8262), .ZN(n8261) );
  AOI21_X1 U8773 ( .B1(n8260), .B2(n8262), .A(n8259), .ZN(n8258) );
  INV_X1 U8774 ( .A(n9925), .ZN(n8259) );
  INV_X1 U8775 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n9897) );
  OR2_X1 U8776 ( .A1(n9896), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9899) );
  NAND2_X1 U8777 ( .A1(n7701), .A2(n9787), .ZN(n9797) );
  AND2_X1 U8778 ( .A1(n9798), .A2(n9788), .ZN(n9796) );
  XNOR2_X1 U8779 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9786) );
  NOR2_X1 U8780 ( .A1(n7746), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9785) );
  AND2_X1 U8781 ( .A1(n7803), .A2(n7682), .ZN(n7681) );
  INV_X1 U8782 ( .A(n8171), .ZN(n7682) );
  OR2_X1 U8783 ( .A1(n8171), .A2(n11719), .ZN(n8170) );
  NAND2_X1 U8784 ( .A1(n8790), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8812) );
  INV_X1 U8785 ( .A(n8792), .ZN(n8790) );
  INV_X1 U8786 ( .A(n13859), .ZN(n7673) );
  OR2_X1 U8787 ( .A1(n10891), .A2(n10378), .ZN(n8167) );
  NAND2_X1 U8788 ( .A1(n8928), .A2(n8927), .ZN(n8943) );
  INV_X1 U8789 ( .A(n8926), .ZN(n8928) );
  INV_X1 U8790 ( .A(n12544), .ZN(n7678) );
  XNOR2_X1 U8791 ( .A(n7433), .B(n7981), .ZN(n10966) );
  AND2_X1 U8792 ( .A1(n11910), .A2(n11716), .ZN(n7803) );
  NAND2_X1 U8793 ( .A1(n9153), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n14221) );
  INV_X1 U8794 ( .A(n8851), .ZN(n9154) );
  OR2_X1 U8795 ( .A1(n14218), .A2(n8576), .ZN(n8577) );
  AND2_X1 U8796 ( .A1(n9037), .A2(n9024), .ZN(n14498) );
  OR2_X1 U8797 ( .A1(n8958), .A2(n12550), .ZN(n8974) );
  NAND2_X1 U8798 ( .A1(n14572), .A2(n14551), .ZN(n14550) );
  AND2_X1 U8799 ( .A1(n14595), .A2(n14577), .ZN(n14572) );
  AND2_X1 U8800 ( .A1(n9133), .A2(n8933), .ZN(n14567) );
  AND2_X1 U8801 ( .A1(n8198), .A2(n8196), .ZN(n8195) );
  INV_X1 U8802 ( .A(n14586), .ZN(n8196) );
  NAND2_X1 U8803 ( .A1(n8197), .A2(n8198), .ZN(n14585) );
  NAND2_X1 U8804 ( .A1(n12520), .A2(n9109), .ZN(n14611) );
  OAI21_X1 U8805 ( .B1(n12375), .B2(n8235), .A(n8234), .ZN(n14610) );
  INV_X1 U8806 ( .A(n8870), .ZN(n8869) );
  NAND2_X1 U8807 ( .A1(n12435), .A2(n14769), .ZN(n12519) );
  NOR2_X1 U8808 ( .A1(n12376), .A2(n7757), .ZN(n12435) );
  NAND2_X1 U8809 ( .A1(n7969), .A2(n7968), .ZN(n12376) );
  NAND2_X1 U8810 ( .A1(n11942), .A2(n9123), .ZN(n12085) );
  NAND2_X1 U8811 ( .A1(n9122), .A2(n8209), .ZN(n11942) );
  AOI21_X1 U8812 ( .B1(n11646), .B2(n7690), .A(n7506), .ZN(n7689) );
  INV_X1 U8813 ( .A(n8739), .ZN(n7690) );
  NAND2_X1 U8814 ( .A1(n11607), .A2(n7475), .ZN(n7654) );
  NAND2_X1 U8815 ( .A1(n11607), .A2(n9119), .ZN(n11631) );
  INV_X1 U8816 ( .A(n14629), .ZN(n7959) );
  NAND2_X1 U8817 ( .A1(n9107), .A2(n7960), .ZN(n11605) );
  OR2_X1 U8818 ( .A1(n8692), .A2(n8691), .ZN(n8710) );
  NAND2_X1 U8819 ( .A1(n11406), .A2(n8676), .ZN(n11389) );
  AND2_X1 U8820 ( .A1(n8676), .A2(n8675), .ZN(n14295) );
  NAND2_X1 U8821 ( .A1(n11167), .A2(n8194), .ZN(n11166) );
  NAND2_X1 U8822 ( .A1(n9107), .A2(n11378), .ZN(n11413) );
  XNOR2_X1 U8823 ( .A(n14363), .B(n14034), .ZN(n14290) );
  NAND2_X1 U8824 ( .A1(n7688), .A2(n8589), .ZN(n10753) );
  INV_X1 U8825 ( .A(n14289), .ZN(n10752) );
  NOR2_X1 U8826 ( .A1(n11346), .A2(n16381), .ZN(n11345) );
  NAND2_X1 U8827 ( .A1(n14255), .A2(n14254), .ZN(n14429) );
  CLKBUF_X1 U8828 ( .A(n8921), .Z(n14253) );
  NAND2_X1 U8829 ( .A1(n8789), .A2(n8788), .ZN(n14101) );
  AND2_X1 U8830 ( .A1(n10822), .A2(n10396), .ZN(n16382) );
  AND2_X1 U8831 ( .A1(n8613), .A2(n8615), .ZN(n8627) );
  NOR2_X1 U8832 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n8581) );
  INV_X1 U8833 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9762) );
  INV_X1 U8834 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9340) );
  NAND2_X1 U8835 ( .A1(n9560), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9559) );
  OR2_X1 U8836 ( .A1(n9341), .A2(n9340), .ZN(n9356) );
  INV_X1 U8837 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9355) );
  INV_X1 U8838 ( .A(n9228), .ZN(n9218) );
  NAND2_X1 U8839 ( .A1(n9463), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9490) );
  INV_X1 U8840 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9308) );
  INV_X1 U8841 ( .A(n9559), .ZN(n9229) );
  NAND2_X1 U8842 ( .A1(n9229), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9228) );
  AOI21_X1 U8843 ( .B1(n8350), .B2(n8349), .A(n7496), .ZN(n8348) );
  INV_X1 U8844 ( .A(n11269), .ZN(n8352) );
  NAND2_X1 U8845 ( .A1(n7648), .A2(n11277), .ZN(n7647) );
  NAND2_X1 U8846 ( .A1(n11792), .A2(n11791), .ZN(n12035) );
  OR2_X1 U8847 ( .A1(n9356), .A2(n9355), .ZN(n9371) );
  INV_X1 U8848 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9370) );
  NAND2_X1 U8849 ( .A1(n8360), .A2(n8359), .ZN(n8363) );
  INV_X1 U8850 ( .A(n14988), .ZN(n8360) );
  AND2_X1 U8851 ( .A1(n9516), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9545) );
  NAND2_X1 U8852 ( .A1(n9415), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9448) );
  INV_X1 U8853 ( .A(n14946), .ZN(n12469) );
  NAND2_X1 U8854 ( .A1(n8357), .A2(n8358), .ZN(n14994) );
  AOI21_X1 U8855 ( .B1(n8361), .B2(n14989), .A(n7531), .ZN(n8358) );
  NAND2_X1 U8856 ( .A1(n14994), .A2(n14995), .ZN(n14993) );
  OR2_X1 U8857 ( .A1(n9448), .A2(n9447), .ZN(n9464) );
  INV_X1 U8858 ( .A(n14830), .ZN(n14918) );
  AND3_X1 U8859 ( .A1(n7434), .A2(n15231), .A3(n8015), .ZN(n15261) );
  NOR2_X1 U8860 ( .A1(n8016), .A2(n15259), .ZN(n8015) );
  XNOR2_X1 U8861 ( .A(n15648), .B(n15299), .ZN(n8016) );
  AND4_X1 U8862 ( .A1(n9613), .A2(n9612), .A3(n9611), .A4(n9610), .ZN(n15192)
         );
  NAND4_X1 U8863 ( .A1(n9251), .A2(n9250), .A3(n9249), .A4(n9248), .ZN(n11576)
         );
  OR2_X1 U8864 ( .A1(n15195), .A2(n9246), .ZN(n9249) );
  NOR3_X1 U8865 ( .A1(n10567), .A2(n11580), .A3(n15887), .ZN(n15328) );
  INV_X1 U8866 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n15950) );
  AOI21_X1 U8867 ( .B1(n15371), .B2(n15370), .A(n15369), .ZN(n16282) );
  AOI21_X1 U8868 ( .B1(n16279), .B2(n10623), .A(n10622), .ZN(n10625) );
  OR2_X1 U8869 ( .A1(n10859), .A2(n10858), .ZN(n15382) );
  AOI21_X1 U8870 ( .B1(n15382), .B2(n15381), .A(n15380), .ZN(n15379) );
  OR2_X1 U8871 ( .A1(n10765), .A2(n10764), .ZN(n10766) );
  NOR2_X1 U8872 ( .A1(n15406), .A2(n15405), .ZN(n15920) );
  NOR2_X1 U8873 ( .A1(n15470), .A2(n8112), .ZN(n15430) );
  NAND2_X1 U8874 ( .A1(n8111), .A2(n8110), .ZN(n15429) );
  NOR2_X1 U8875 ( .A1(n15232), .A2(n8112), .ZN(n8110) );
  INV_X1 U8876 ( .A(n15470), .ZN(n8111) );
  INV_X1 U8877 ( .A(n15258), .ZN(n15445) );
  INV_X1 U8878 ( .A(n9572), .ZN(n9573) );
  NAND2_X1 U8879 ( .A1(n8437), .A2(n7493), .ZN(n8434) );
  NAND2_X1 U8880 ( .A1(n15531), .A2(n8105), .ZN(n15511) );
  NAND2_X1 U8881 ( .A1(n15531), .A2(n15688), .ZN(n15530) );
  NAND2_X1 U8882 ( .A1(n15583), .A2(n8449), .ZN(n15555) );
  AOI21_X1 U8883 ( .B1(n8287), .B2(n15625), .A(n7501), .ZN(n8285) );
  INV_X1 U8884 ( .A(n8287), .ZN(n8286) );
  NAND2_X1 U8885 ( .A1(n8099), .A2(n8098), .ZN(n15613) );
  INV_X1 U8886 ( .A(n8099), .ZN(n15632) );
  NAND2_X1 U8887 ( .A1(n12153), .A2(n9658), .ZN(n12289) );
  NOR2_X1 U8888 ( .A1(n8108), .A2(n16572), .ZN(n8107) );
  INV_X1 U8889 ( .A(n8109), .ZN(n8108) );
  AND2_X1 U8890 ( .A1(n9714), .A2(n15212), .ZN(n15038) );
  INV_X1 U8891 ( .A(n15241), .ZN(n9653) );
  NAND2_X1 U8892 ( .A1(n11772), .A2(n16511), .ZN(n12003) );
  INV_X1 U8893 ( .A(n15240), .ZN(n11767) );
  NOR2_X1 U8894 ( .A1(n16439), .A2(n16465), .ZN(n16475) );
  NAND2_X1 U8895 ( .A1(n9307), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9341) );
  NAND2_X1 U8896 ( .A1(n12110), .A2(n15055), .ZN(n16438) );
  NAND2_X1 U8897 ( .A1(n8097), .A2(n8096), .ZN(n16439) );
  INV_X1 U8898 ( .A(n16438), .ZN(n8097) );
  INV_X1 U8899 ( .A(n15016), .ZN(n15008) );
  INV_X1 U8900 ( .A(n15293), .ZN(n15006) );
  NAND2_X1 U8901 ( .A1(n10405), .A2(n9318), .ZN(n8299) );
  NOR2_X1 U8902 ( .A1(n12107), .A2(n16396), .ZN(n12110) );
  AND2_X1 U8903 ( .A1(n15471), .A2(n15470), .ZN(n15663) );
  AND2_X1 U8904 ( .A1(n15497), .A2(n9672), .ZN(n15484) );
  INV_X1 U8905 ( .A(n16473), .ZN(n16437) );
  AND2_X1 U8906 ( .A1(n11977), .A2(n9628), .ZN(n16573) );
  INV_X1 U8907 ( .A(n16573), .ZN(n16476) );
  NOR2_X1 U8908 ( .A1(n15783), .A2(n9679), .ZN(n16486) );
  XNOR2_X1 U8909 ( .A(n14252), .B(n7623), .ZN(n15200) );
  NAND2_X1 U8910 ( .A1(n8003), .A2(n8004), .ZN(n14252) );
  OR2_X1 U8911 ( .A1(n9091), .A2(n8007), .ZN(n8003) );
  NAND2_X1 U8912 ( .A1(n14224), .A2(n9097), .ZN(n12790) );
  NAND2_X1 U8913 ( .A1(n9096), .A2(n9095), .ZN(n14224) );
  OR2_X1 U8914 ( .A1(n9096), .A2(n9095), .ZN(n9097) );
  XNOR2_X1 U8915 ( .A(n9051), .B(n9046), .ZN(n14786) );
  XNOR2_X1 U8916 ( .A(n8994), .B(SI_24_), .ZN(n12104) );
  NAND2_X1 U8917 ( .A1(n9619), .A2(n7489), .ZN(n15213) );
  MUX2_X1 U8918 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9617), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n9619) );
  INV_X1 U8919 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n13801) );
  INV_X1 U8920 ( .A(n9509), .ZN(n9511) );
  XNOR2_X1 U8921 ( .A(n8900), .B(n8899), .ZN(n11600) );
  XNOR2_X1 U8922 ( .A(n8864), .B(n8863), .ZN(n11546) );
  OAI21_X1 U8923 ( .B1(n8819), .B2(n8839), .A(n7480), .ZN(n8432) );
  OAI21_X1 U8924 ( .B1(n9381), .B2(P1_IR_REG_9__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9395) );
  OR2_X1 U8925 ( .A1(n9350), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9364) );
  NAND2_X1 U8926 ( .A1(n8682), .A2(n8681), .ZN(n8703) );
  NAND2_X1 U8927 ( .A1(n8679), .A2(n8678), .ZN(n8682) );
  AND2_X1 U8928 ( .A1(n15932), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n15938) );
  XNOR2_X1 U8929 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n15937) );
  XNOR2_X1 U8930 ( .A(n15968), .B(n16300), .ZN(n15972) );
  AOI21_X1 U8931 ( .B1(n15979), .B2(n15978), .A(n15977), .ZN(n15987) );
  NAND2_X1 U8932 ( .A1(n15993), .A2(n15994), .ZN(n16002) );
  AOI21_X1 U8933 ( .B1(n16015), .B2(n16014), .A(n16013), .ZN(n16025) );
  NOR2_X1 U8934 ( .A1(n7636), .A2(n16064), .ZN(n16073) );
  INV_X1 U8935 ( .A(n16067), .ZN(n7636) );
  OR2_X1 U8936 ( .A1(n7829), .A2(n7828), .ZN(n12018) );
  NOR2_X1 U8937 ( .A1(n7833), .A2(n7832), .ZN(n7829) );
  OAI21_X1 U8938 ( .B1(n8490), .B2(n7832), .A(n11687), .ZN(n7828) );
  AOI21_X1 U8939 ( .B1(n13114), .B2(n10247), .A(n10238), .ZN(n13125) );
  NAND2_X1 U8940 ( .A1(n12935), .A2(n12801), .ZN(n12858) );
  NAND2_X1 U8941 ( .A1(n12204), .A2(n12203), .ZN(n12266) );
  NAND2_X1 U8942 ( .A1(n12878), .A2(n12877), .ZN(n12876) );
  AND4_X1 U8943 ( .A1(n9881), .A2(n9880), .A3(n9879), .A4(n9878), .ZN(n12022)
         );
  NOR2_X1 U8944 ( .A1(n10977), .A2(n10951), .ZN(n10952) );
  AND2_X1 U8945 ( .A1(n12997), .A2(n10950), .ZN(n10951) );
  AOI21_X1 U8946 ( .B1(n11626), .B2(n12821), .A(n16311), .ZN(n10953) );
  NAND2_X1 U8947 ( .A1(n12922), .A2(n12819), .ZN(n12883) );
  INV_X1 U8948 ( .A(n8481), .ZN(n8480) );
  NAND2_X1 U8949 ( .A1(n12972), .A2(n8510), .ZN(n12900) );
  NOR2_X1 U8950 ( .A1(n11514), .A2(n11513), .ZN(n11516) );
  NAND2_X1 U8951 ( .A1(n12908), .A2(n12907), .ZN(n12906) );
  NAND2_X1 U8952 ( .A1(n12898), .A2(n12809), .ZN(n12908) );
  NAND2_X1 U8953 ( .A1(n12865), .A2(n13188), .ZN(n7840) );
  NAND2_X1 U8954 ( .A1(n11293), .A2(n9810), .ZN(n11294) );
  NOR2_X1 U8955 ( .A1(n11298), .A2(n11297), .ZN(n11514) );
  AND4_X1 U8956 ( .A1(n9895), .A2(n9894), .A3(n9893), .A4(n9892), .ZN(n12140)
         );
  NAND2_X1 U8957 ( .A1(n9778), .A2(n9777), .ZN(n10813) );
  NAND2_X1 U8958 ( .A1(n12876), .A2(n12816), .ZN(n12924) );
  NAND2_X1 U8959 ( .A1(n7847), .A2(n12793), .ZN(n12937) );
  XNOR2_X1 U8960 ( .A(n12825), .B(n12826), .ZN(n12943) );
  NAND2_X1 U8961 ( .A1(n8483), .A2(n8486), .ZN(n12951) );
  AND2_X1 U8962 ( .A1(n12952), .A2(n8487), .ZN(n8486) );
  OR2_X1 U8963 ( .A1(n12907), .A2(n8488), .ZN(n8487) );
  NAND2_X1 U8964 ( .A1(n12906), .A2(n12811), .ZN(n12953) );
  NAND2_X1 U8965 ( .A1(n10812), .A2(n16360), .ZN(n12966) );
  XNOR2_X1 U8966 ( .A(n12839), .B(n12983), .ZN(n12963) );
  OR2_X1 U8967 ( .A1(n12971), .A2(n12970), .ZN(n12972) );
  NAND2_X1 U8968 ( .A1(n10802), .A2(n10801), .ZN(n12978) );
  XNOR2_X1 U8969 ( .A(n12579), .B(n13086), .ZN(n8124) );
  NAND2_X1 U8970 ( .A1(n12734), .A2(n10346), .ZN(n8272) );
  AND2_X1 U8971 ( .A1(n11439), .A2(n11438), .ZN(n13091) );
  AND2_X1 U8972 ( .A1(n11439), .A2(n10268), .ZN(n12574) );
  AND2_X1 U8973 ( .A1(n11439), .A2(n10252), .ZN(n13109) );
  INV_X1 U8974 ( .A(n12891), .ZN(n12832) );
  INV_X1 U8975 ( .A(n13254), .ZN(n12988) );
  INV_X1 U8976 ( .A(n12228), .ZN(n12452) );
  NOR2_X1 U8977 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n11452), .ZN(n13008) );
  OAI21_X1 U8978 ( .B1(n16120), .B2(n11094), .A(n11093), .ZN(n11092) );
  INV_X1 U8979 ( .A(n7769), .ZN(n11252) );
  NAND2_X1 U8980 ( .A1(n11247), .A2(n11248), .ZN(n16133) );
  INV_X1 U8981 ( .A(n8082), .ZN(n16136) );
  NAND2_X1 U8982 ( .A1(n8060), .A2(n8062), .ZN(n11671) );
  AOI21_X1 U8983 ( .B1(n8066), .B2(n8064), .A(n8063), .ZN(n8062) );
  NOR2_X1 U8984 ( .A1(n11668), .A2(n11667), .ZN(n8063) );
  XNOR2_X1 U8985 ( .A(n11830), .B(n11817), .ZN(n11661) );
  INV_X1 U8986 ( .A(n7749), .ZN(n11816) );
  INV_X1 U8987 ( .A(n8058), .ZN(n16245) );
  XNOR2_X1 U8988 ( .A(n13082), .B(n8050), .ZN(n8049) );
  INV_X1 U8989 ( .A(n13081), .ZN(n8050) );
  OAI21_X1 U8990 ( .B1(n7478), .B2(n13104), .A(n7553), .ZN(n13318) );
  XNOR2_X1 U8991 ( .A(n13118), .B(n13119), .ZN(n13324) );
  NAND2_X1 U8992 ( .A1(n13144), .A2(n10192), .ZN(n13133) );
  NAND2_X1 U8993 ( .A1(n10119), .A2(n10118), .ZN(n13349) );
  NAND2_X1 U8994 ( .A1(n13212), .A2(n10113), .ZN(n13202) );
  NOR2_X1 U8995 ( .A1(n7936), .A2(n7935), .ZN(n8505) );
  INV_X1 U8996 ( .A(n10099), .ZN(n7935) );
  NAND2_X1 U8997 ( .A1(n7924), .A2(n10068), .ZN(n13235) );
  NAND2_X1 U8998 ( .A1(n13249), .A2(n13263), .ZN(n7924) );
  AND2_X1 U8999 ( .A1(n13265), .A2(n12683), .ZN(n13240) );
  AND2_X1 U9000 ( .A1(n8133), .A2(n12662), .ZN(n13283) );
  NAND2_X1 U9001 ( .A1(n10286), .A2(n12658), .ZN(n13298) );
  NAND2_X1 U9002 ( .A1(n9993), .A2(n9992), .ZN(n16594) );
  NAND2_X1 U9003 ( .A1(n12193), .A2(n9963), .ZN(n12226) );
  NOR2_X1 U9004 ( .A1(n7929), .A2(n7928), .ZN(n8521) );
  INV_X1 U9005 ( .A(n9930), .ZN(n7928) );
  INV_X1 U9006 ( .A(n13313), .ZN(n13266) );
  INV_X1 U9007 ( .A(n10976), .ZN(n16363) );
  NAND2_X1 U9008 ( .A1(n10811), .A2(n10810), .ZN(n16360) );
  NAND2_X1 U9009 ( .A1(n12571), .A2(n12570), .ZN(n13384) );
  NAND2_X1 U9010 ( .A1(n10157), .A2(n10156), .ZN(n13400) );
  AND2_X1 U9011 ( .A1(n10074), .A2(n10073), .ZN(n13820) );
  NAND2_X1 U9012 ( .A1(n10012), .A2(n10011), .ZN(n13836) );
  INV_X1 U9013 ( .A(n11859), .ZN(n11862) );
  XNOR2_X1 U9014 ( .A(n12556), .B(n10244), .ZN(n13849) );
  NAND2_X1 U9015 ( .A1(n8147), .A2(n8149), .ZN(n9756) );
  NAND2_X1 U9016 ( .A1(n10310), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9769) );
  INV_X1 U9017 ( .A(n10332), .ZN(n12031) );
  AND2_X1 U9018 ( .A1(n10316), .A2(n10312), .ZN(n11681) );
  OAI211_X1 U9019 ( .C1(n10166), .C2(n12191), .A(n7716), .B(n7712), .ZN(n10181) );
  NAND2_X1 U9020 ( .A1(n10166), .A2(n7621), .ZN(n7712) );
  NAND2_X1 U9021 ( .A1(n10133), .A2(n10132), .ZN(n10137) );
  XNOR2_X1 U9022 ( .A(n10257), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12773) );
  NAND2_X1 U9023 ( .A1(n10259), .A2(n10306), .ZN(n11377) );
  MUX2_X1 U9024 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10258), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n10259) );
  INV_X1 U9025 ( .A(n10303), .ZN(n11216) );
  NAND2_X1 U9026 ( .A1(n7729), .A2(n10084), .ZN(n10103) );
  NAND2_X1 U9027 ( .A1(n10083), .A2(n10082), .ZN(n7729) );
  NAND2_X1 U9028 ( .A1(n8254), .A2(n10057), .ZN(n10070) );
  NAND2_X1 U9029 ( .A1(n10056), .A2(n10055), .ZN(n8254) );
  NAND2_X1 U9030 ( .A1(n7742), .A2(n10024), .ZN(n10040) );
  NAND2_X1 U9031 ( .A1(n7737), .A2(n9975), .ZN(n9989) );
  NAND2_X1 U9032 ( .A1(n7791), .A2(n7738), .ZN(n7737) );
  NAND2_X1 U9033 ( .A1(n7791), .A2(n9955), .ZN(n9974) );
  NAND2_X1 U9034 ( .A1(n8264), .A2(n8262), .ZN(n9926) );
  NAND2_X1 U9035 ( .A1(n8264), .A2(n9902), .ZN(n9907) );
  NAND2_X1 U9036 ( .A1(n9883), .A2(n9882), .ZN(n9904) );
  NAND2_X1 U9037 ( .A1(P3_U3151), .A2(n8155), .ZN(n13850) );
  OAI21_X1 U9038 ( .B1(n9823), .B2(n7723), .A(n7721), .ZN(n9865) );
  NAND2_X1 U9039 ( .A1(n7726), .A2(n9824), .ZN(n9846) );
  NAND2_X1 U9040 ( .A1(n9823), .A2(n9822), .ZN(n7726) );
  AND2_X1 U9041 ( .A1(n13981), .A2(n13874), .ZN(n13877) );
  NAND2_X1 U9042 ( .A1(n7664), .A2(n7971), .ZN(n7663) );
  INV_X1 U9043 ( .A(n7667), .ZN(n7664) );
  AND2_X1 U9044 ( .A1(n10649), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13985) );
  INV_X1 U9045 ( .A(n13918), .ZN(n13910) );
  NAND2_X1 U9046 ( .A1(n13981), .A2(n8182), .ZN(n13918) );
  AND2_X1 U9047 ( .A1(n13876), .A2(n13874), .ZN(n8182) );
  NOR2_X1 U9048 ( .A1(n13860), .A2(n13859), .ZN(n13862) );
  XNOR2_X1 U9049 ( .A(n10958), .B(n10966), .ZN(n10893) );
  NAND2_X1 U9050 ( .A1(n7970), .A2(n11233), .ZN(n11403) );
  NAND2_X1 U9051 ( .A1(n11237), .A2(n11227), .ZN(n7970) );
  NAND2_X1 U9052 ( .A1(n13948), .A2(n13949), .ZN(n13923) );
  NAND2_X1 U9053 ( .A1(n12542), .A2(n8179), .ZN(n8178) );
  AOI21_X1 U9054 ( .B1(n11915), .B2(n11719), .A(n8171), .ZN(n11899) );
  NAND2_X1 U9055 ( .A1(n11879), .A2(n7803), .ZN(n11915) );
  NAND2_X1 U9056 ( .A1(n7666), .A2(n7665), .ZN(n11880) );
  AOI21_X1 U9057 ( .B1(n7662), .B2(n11399), .A(n7479), .ZN(n7665) );
  NAND2_X1 U9058 ( .A1(n7982), .A2(n10851), .ZN(n10857) );
  NAND2_X1 U9059 ( .A1(n12539), .A2(n12538), .ZN(n13965) );
  NAND2_X1 U9060 ( .A1(n11136), .A2(n11135), .ZN(n11221) );
  NAND2_X1 U9061 ( .A1(n12305), .A2(n8172), .ZN(n12392) );
  INV_X1 U9062 ( .A(n8172), .ZN(n8169) );
  NAND2_X1 U9063 ( .A1(n10394), .A2(n14624), .ZN(n13983) );
  NAND4_X1 U9064 ( .A1(n8659), .A2(n8658), .A3(n8657), .A4(n8656), .ZN(n14361)
         );
  NAND2_X1 U9065 ( .A1(n7946), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8569) );
  XNOR2_X1 U9066 ( .A(n14438), .B(n14732), .ZN(n14431) );
  XNOR2_X1 U9067 ( .A(n9146), .B(n14314), .ZN(n8205) );
  INV_X1 U9068 ( .A(n14314), .ZN(n9105) );
  XNOR2_X1 U9069 ( .A(n9738), .B(n14312), .ZN(n14461) );
  NAND2_X1 U9070 ( .A1(n8242), .A2(n9741), .ZN(n14454) );
  NAND2_X1 U9071 ( .A1(n14476), .A2(n9045), .ZN(n14463) );
  XNOR2_X1 U9072 ( .A(n7655), .B(n14313), .ZN(n14480) );
  AOI21_X1 U9073 ( .B1(n14492), .B2(n14310), .A(n7596), .ZN(n7655) );
  NAND2_X1 U9074 ( .A1(n14504), .A2(n9006), .ZN(n14490) );
  NAND2_X1 U9075 ( .A1(n14542), .A2(n8966), .ZN(n14519) );
  AND2_X1 U9076 ( .A1(n7700), .A2(n7699), .ZN(n14543) );
  NAND2_X1 U9077 ( .A1(n14547), .A2(n9135), .ZN(n14532) );
  NOR2_X1 U9078 ( .A1(n14558), .A2(n8221), .ZN(n8220) );
  INV_X1 U9079 ( .A(n8934), .ZN(n8221) );
  NAND2_X1 U9080 ( .A1(n8203), .A2(n9130), .ZN(n14604) );
  NAND2_X1 U9081 ( .A1(n12514), .A2(n9129), .ZN(n8203) );
  NAND2_X1 U9082 ( .A1(n12433), .A2(n8857), .ZN(n12524) );
  AND2_X1 U9083 ( .A1(n12375), .A2(n8837), .ZN(n12434) );
  NAND2_X1 U9084 ( .A1(n12284), .A2(n8818), .ZN(n12373) );
  AND2_X1 U9085 ( .A1(n12082), .A2(n8799), .ZN(n12282) );
  NAND2_X1 U9086 ( .A1(n7944), .A2(n8739), .ZN(n11645) );
  NAND2_X1 U9087 ( .A1(n8226), .A2(n8641), .ZN(n11164) );
  INV_X1 U9088 ( .A(n7956), .ZN(n10361) );
  OAI21_X1 U9089 ( .B1(n10777), .B2(n7957), .A(n14430), .ZN(n7956) );
  NAND2_X1 U9090 ( .A1(n10405), .A2(n8612), .ZN(n8180) );
  XNOR2_X1 U9091 ( .A(n11344), .B(n8183), .ZN(n16385) );
  OAI21_X1 U9092 ( .B1(n8183), .B2(n11351), .A(n11350), .ZN(n11352) );
  OR2_X1 U9093 ( .A1(n15822), .A2(n10386), .ZN(n14624) );
  NAND2_X1 U9094 ( .A1(n11368), .A2(n10393), .ZN(n14619) );
  AND2_X1 U9095 ( .A1(n11368), .A2(n14424), .ZN(n14632) );
  AND2_X1 U9096 ( .A1(n14638), .A2(n14641), .ZN(n14729) );
  INV_X1 U9097 ( .A(n14429), .ZN(n14736) );
  AOI211_X1 U9098 ( .C1(n14717), .C2(n14656), .A(n14655), .B(n14654), .ZN(
        n14741) );
  AND2_X1 U9099 ( .A1(n7953), .A2(n8558), .ZN(n7952) );
  INV_X1 U9100 ( .A(n8551), .ZN(n8549) );
  OAI21_X1 U9101 ( .B1(n8551), .B2(n7661), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7660) );
  INV_X1 U9102 ( .A(n7953), .ZN(n7661) );
  XNOR2_X1 U9103 ( .A(n8552), .B(n8548), .ZN(n14782) );
  XNOR2_X1 U9104 ( .A(n9164), .B(P2_IR_REG_26__SCAN_IN), .ZN(n14785) );
  NAND2_X1 U9105 ( .A1(n8531), .A2(n8530), .ZN(n8535) );
  NOR2_X1 U9106 ( .A1(n14772), .A2(n8532), .ZN(n8530) );
  INV_X1 U9107 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10473) );
  INV_X1 U9108 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10460) );
  INV_X1 U9109 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10448) );
  INV_X1 U9110 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10444) );
  INV_X1 U9111 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10408) );
  INV_X1 U9112 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10411) );
  NAND2_X1 U9113 ( .A1(n14781), .A2(n15206), .ZN(n9580) );
  NAND2_X1 U9114 ( .A1(n7644), .A2(n14801), .ZN(n16607) );
  AOI21_X1 U9115 ( .B1(n8393), .B2(n11795), .A(n7548), .ZN(n8392) );
  NAND2_X1 U9116 ( .A1(n8356), .A2(n11273), .ZN(n16400) );
  INV_X1 U9117 ( .A(n8364), .ZN(n14924) );
  OR2_X1 U9118 ( .A1(n8373), .A2(n8368), .ZN(n8367) );
  AND2_X1 U9119 ( .A1(n8366), .A2(n7570), .ZN(n8365) );
  NAND2_X1 U9120 ( .A1(n14778), .A2(n15206), .ZN(n9592) );
  NAND2_X1 U9121 ( .A1(n8363), .A2(n8361), .ZN(n14931) );
  NAND2_X1 U9122 ( .A1(n12463), .A2(n12462), .ZN(n14945) );
  INV_X1 U9123 ( .A(n8372), .ZN(n8369) );
  AND2_X1 U9124 ( .A1(n8391), .A2(n8389), .ZN(n8388) );
  NAND2_X1 U9125 ( .A1(n8390), .A2(n8391), .ZN(n14958) );
  NOR2_X1 U9126 ( .A1(n14959), .A2(n8386), .ZN(n8384) );
  OR2_X1 U9127 ( .A1(n14824), .A2(n14815), .ZN(n8383) );
  NAND2_X1 U9128 ( .A1(n12035), .A2(n12034), .ZN(n12216) );
  INV_X1 U9129 ( .A(n8363), .ZN(n14987) );
  NAND2_X1 U9130 ( .A1(n9430), .A2(n9429), .ZN(n15105) );
  OAI22_X1 U9131 ( .A1(n7639), .A2(n15016), .B1(n9269), .B2(n15293), .ZN(
        n11989) );
  INV_X1 U9132 ( .A(n15029), .ZN(n16612) );
  NAND2_X1 U9133 ( .A1(n8391), .A2(n8385), .ZN(n15024) );
  NAND2_X1 U9134 ( .A1(n14814), .A2(n14815), .ZN(n8385) );
  AND2_X1 U9135 ( .A1(n16398), .A2(n16573), .ZN(n16610) );
  OR2_X1 U9136 ( .A1(n11280), .A2(P1_U3086), .ZN(n15294) );
  NAND4_X1 U9137 ( .A1(n9590), .A2(n9589), .A3(n9588), .A4(n9587), .ZN(n15302)
         );
  AOI21_X1 U9138 ( .B1(n10766), .B2(n10575), .A(n10574), .ZN(n10725) );
  AOI21_X1 U9139 ( .B1(n10913), .B2(n10912), .A(n10911), .ZN(n11488) );
  NAND2_X1 U9140 ( .A1(n15209), .A2(n15208), .ZN(n15427) );
  OAI21_X1 U9141 ( .B1(n7434), .B2(n8418), .A(n8417), .ZN(n8416) );
  NAND2_X1 U9142 ( .A1(n8411), .A2(n8409), .ZN(n8420) );
  NAND2_X1 U9143 ( .A1(n8408), .A2(n7476), .ZN(n8419) );
  INV_X1 U9144 ( .A(n8423), .ZN(n8405) );
  NAND2_X1 U9145 ( .A1(n15485), .A2(n9673), .ZN(n15469) );
  NAND2_X1 U9146 ( .A1(n8439), .A2(n8440), .ZN(n15494) );
  AND2_X1 U9147 ( .A1(n8436), .A2(n8439), .ZN(n15493) );
  AND2_X1 U9148 ( .A1(n15255), .A2(n9670), .ZN(n8291) );
  NAND2_X1 U9149 ( .A1(n8292), .A2(n9670), .ZN(n15521) );
  NOR2_X1 U9150 ( .A1(n7781), .A2(n8443), .ZN(n15510) );
  NAND2_X1 U9151 ( .A1(n9544), .A2(n9543), .ZN(n15694) );
  NAND2_X1 U9152 ( .A1(n8276), .A2(n8280), .ZN(n15544) );
  NAND2_X1 U9153 ( .A1(n15571), .A2(n8282), .ZN(n8276) );
  NAND2_X1 U9154 ( .A1(n8284), .A2(n8283), .ZN(n15560) );
  AND2_X1 U9155 ( .A1(n8284), .A2(n9665), .ZN(n15561) );
  NAND2_X1 U9156 ( .A1(n9531), .A2(n9530), .ZN(n15699) );
  NAND2_X1 U9157 ( .A1(n9503), .A2(n9502), .ZN(n15710) );
  NAND2_X1 U9158 ( .A1(n15628), .A2(n9661), .ZN(n15612) );
  AND2_X1 U9159 ( .A1(n15734), .A2(n9471), .ZN(n15626) );
  INV_X1 U9160 ( .A(n15246), .ZN(n9424) );
  NAND2_X1 U9161 ( .A1(n11954), .A2(n8297), .ZN(n12177) );
  AND2_X1 U9162 ( .A1(n11954), .A2(n9656), .ZN(n12179) );
  OR2_X1 U9163 ( .A1(n16522), .A2(n11978), .ZN(n16512) );
  INV_X2 U9164 ( .A(n16580), .ZN(n16540) );
  AND2_X1 U9165 ( .A1(n7557), .A2(n9213), .ZN(n8478) );
  INV_X1 U9166 ( .A(n9216), .ZN(n15769) );
  NAND2_X1 U9167 ( .A1(n9709), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9686) );
  XNOR2_X1 U9168 ( .A(n8970), .B(n8969), .ZN(n12149) );
  AOI21_X1 U9169 ( .B1(n8968), .B2(n8987), .A(n8967), .ZN(n8970) );
  XNOR2_X1 U9170 ( .A(n9236), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15782) );
  INV_X1 U9171 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10463) );
  INV_X1 U9172 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10456) );
  INV_X1 U9173 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10450) );
  INV_X1 U9174 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10446) );
  INV_X1 U9175 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10406) );
  INV_X1 U9176 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10416) );
  NAND2_X1 U9177 ( .A1(n8155), .A2(P1_U3086), .ZN(n15777) );
  NAND2_X1 U9178 ( .A1(n8157), .A2(n7746), .ZN(n9252) );
  NAND2_X1 U9179 ( .A1(n8156), .A2(SI_0_), .ZN(n8157) );
  INV_X1 U9180 ( .A(P1_RD_REG_SCAN_IN), .ZN(n10404) );
  INV_X1 U9181 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15933) );
  XNOR2_X1 U9182 ( .A(n15972), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15966) );
  NAND2_X1 U9183 ( .A1(n15984), .A2(n8247), .ZN(n16107) );
  INV_X1 U9184 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n8248) );
  NOR2_X1 U9185 ( .A1(n16107), .A2(n16108), .ZN(n16106) );
  XNOR2_X1 U9186 ( .A(n15992), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15990) );
  NAND2_X1 U9187 ( .A1(n15990), .A2(n15989), .ZN(n15993) );
  XNOR2_X1 U9188 ( .A(n16002), .B(n8246), .ZN(n16001) );
  INV_X1 U9189 ( .A(n16003), .ZN(n8246) );
  NAND2_X1 U9190 ( .A1(n7637), .A2(n16018), .ZN(n16020) );
  INV_X1 U9191 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7817) );
  NAND2_X1 U9192 ( .A1(n16049), .A2(n16050), .ZN(n16056) );
  NAND2_X1 U9193 ( .A1(n16056), .A2(n16057), .ZN(n16058) );
  NAND2_X1 U9194 ( .A1(n16073), .A2(n16074), .ZN(n16076) );
  NOR2_X1 U9195 ( .A1(n16073), .A2(n16074), .ZN(n16075) );
  NAND2_X1 U9196 ( .A1(n16076), .A2(n16077), .ZN(n16083) );
  NOR2_X1 U9197 ( .A1(n16086), .A2(n16085), .ZN(n16094) );
  NAND2_X1 U9198 ( .A1(n7861), .A2(n7860), .ZN(P3_U3160) );
  NAND2_X1 U9199 ( .A1(n12838), .A2(n7865), .ZN(n7860) );
  NOR2_X1 U9200 ( .A1(n7529), .A2(n12969), .ZN(n7865) );
  NAND2_X1 U9201 ( .A1(n8073), .A2(n16139), .ZN(n11243) );
  NAND2_X1 U9202 ( .A1(n8061), .A2(n8066), .ZN(n11670) );
  NAND2_X1 U9203 ( .A1(n8046), .A2(n8043), .ZN(P3_U3200) );
  OAI21_X1 U9204 ( .B1(n13073), .B2(n7474), .A(n16194), .ZN(n8046) );
  INV_X1 U9205 ( .A(n8044), .ZN(n8043) );
  NOR2_X1 U9206 ( .A1(n7599), .A2(n7773), .ZN(n7772) );
  NOR2_X1 U9207 ( .A1(n16601), .A2(n10342), .ZN(n7773) );
  INV_X1 U9208 ( .A(n7751), .ZN(n7750) );
  OAI21_X1 U9209 ( .B1(n13390), .B2(n13379), .A(n7752), .ZN(n7751) );
  NOR2_X1 U9210 ( .A1(n7600), .A2(n7771), .ZN(n7770) );
  NOR2_X1 U9211 ( .A1(n16602), .A2(n10352), .ZN(n7771) );
  INV_X1 U9212 ( .A(n7755), .ZN(n7754) );
  OAI22_X1 U9213 ( .A1(n13390), .A2(n13837), .B1(n16602), .B2(n13389), .ZN(
        n7755) );
  INV_X1 U9214 ( .A(n7979), .ZN(n13991) );
  OAI22_X1 U9215 ( .A1(n14447), .A2(n14715), .B1(n16560), .B2(n9191), .ZN(
        n9192) );
  INV_X1 U9216 ( .A(n7819), .ZN(P2_U3526) );
  AOI21_X1 U9217 ( .B1(n14737), .B2(n16560), .A(n7820), .ZN(n7819) );
  OAI22_X1 U9218 ( .A1(n14740), .A2(n14715), .B1(n16560), .B2(n7821), .ZN(
        n7820) );
  INV_X1 U9219 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n7821) );
  NAND2_X1 U9220 ( .A1(n8204), .A2(n11936), .ZN(n9731) );
  OAI22_X1 U9221 ( .A1(n14447), .A2(n14768), .B1(n11936), .B2(n9728), .ZN(
        n9729) );
  NAND2_X1 U9222 ( .A1(n7696), .A2(n9745), .ZN(P2_U3495) );
  NAND2_X1 U9223 ( .A1(n7806), .A2(n7804), .ZN(P2_U3494) );
  AOI21_X1 U9224 ( .B1(n14198), .B2(n9744), .A(n7805), .ZN(n7804) );
  NOR2_X1 U9225 ( .A1(n11936), .A2(n14739), .ZN(n7805) );
  NAND2_X1 U9226 ( .A1(n7802), .A2(n7517), .ZN(n15420) );
  NAND2_X1 U9227 ( .A1(n15418), .A2(n15417), .ZN(n7802) );
  NOR2_X1 U9228 ( .A1(n16034), .A2(n16033), .ZN(n16035) );
  INV_X1 U9229 ( .A(n8244), .ZN(n16044) );
  INV_X1 U9230 ( .A(n16064), .ZN(n16068) );
  XNOR2_X1 U9231 ( .A(n16104), .B(n8250), .ZN(n8249) );
  XNOR2_X1 U9232 ( .A(n16105), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n8250) );
  INV_X2 U9233 ( .A(n14013), .ZN(n14235) );
  AND2_X1 U9234 ( .A1(n15182), .A2(n15184), .ZN(n7462) );
  AND2_X1 U9235 ( .A1(n8913), .A2(SI_20_), .ZN(n7463) );
  AND2_X1 U9236 ( .A1(n8004), .A2(n7623), .ZN(n7464) );
  INV_X1 U9237 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n15760) );
  OR2_X1 U9238 ( .A1(n12022), .A2(n11862), .ZN(n7465) );
  OR2_X1 U9239 ( .A1(n13142), .A2(n7940), .ZN(n7466) );
  INV_X1 U9240 ( .A(n15255), .ZN(n8442) );
  NAND2_X1 U9241 ( .A1(n10214), .A2(n10213), .ZN(n10225) );
  AND2_X1 U9242 ( .A1(n14529), .A2(n14177), .ZN(n7467) );
  NAND2_X1 U9243 ( .A1(n15497), .A2(n7498), .ZN(n15485) );
  AND2_X1 U9244 ( .A1(n14093), .A2(n14092), .ZN(n7468) );
  AND2_X1 U9245 ( .A1(n12717), .A2(n12718), .ZN(n13123) );
  XNOR2_X1 U9246 ( .A(n8704), .B(SI_8_), .ZN(n8701) );
  AND2_X1 U9247 ( .A1(n7554), .A2(n7886), .ZN(n7469) );
  AND2_X1 U9248 ( .A1(n7558), .A2(n8302), .ZN(n7470) );
  NAND2_X1 U9249 ( .A1(n14097), .A2(n7468), .ZN(n8328) );
  INV_X1 U9250 ( .A(n8328), .ZN(n8327) );
  OR2_X1 U9251 ( .A1(n7841), .A2(n12831), .ZN(n7471) );
  INV_X1 U9252 ( .A(n16316), .ZN(n8116) );
  INV_X1 U9253 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14772) );
  OR2_X1 U9254 ( .A1(n14959), .A2(n8387), .ZN(n7472) );
  INV_X1 U9255 ( .A(n14989), .ZN(n8359) );
  NAND2_X1 U9256 ( .A1(n9580), .A2(n9579), .ZN(n15659) );
  INV_X1 U9257 ( .A(n8661), .ZN(n8662) );
  XNOR2_X1 U9258 ( .A(n8664), .B(SI_6_), .ZN(n8661) );
  AND2_X1 U9259 ( .A1(n8972), .A2(n8971), .ZN(n14529) );
  INV_X1 U9260 ( .A(n14529), .ZN(n14671) );
  NAND2_X1 U9261 ( .A1(n14725), .A2(n14107), .ZN(n7473) );
  INV_X1 U9262 ( .A(n13123), .ZN(n13119) );
  INV_X1 U9263 ( .A(n12794), .ZN(n7848) );
  AND2_X1 U9264 ( .A1(n10206), .A2(n10205), .ZN(n13126) );
  AND2_X1 U9265 ( .A1(n13062), .A2(n13061), .ZN(n7474) );
  INV_X1 U9266 ( .A(n8324), .ZN(n8323) );
  NAND2_X1 U9267 ( .A1(n8325), .A2(n14103), .ZN(n8324) );
  AND2_X1 U9268 ( .A1(n7550), .A2(n9119), .ZN(n7475) );
  AND2_X1 U9269 ( .A1(n7552), .A2(n8406), .ZN(n7476) );
  AND2_X1 U9270 ( .A1(n8646), .A2(SI_5_), .ZN(n7477) );
  INV_X1 U9271 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n9768) );
  AND2_X1 U9272 ( .A1(n8145), .A2(n12718), .ZN(n7478) );
  AND2_X1 U9273 ( .A1(n11710), .A2(n11709), .ZN(n7479) );
  OR2_X1 U9274 ( .A1(n8820), .A2(SI_14_), .ZN(n7480) );
  INV_X1 U9275 ( .A(n12914), .ZN(n7841) );
  XNOR2_X1 U9276 ( .A(n12833), .B(n12832), .ZN(n12914) );
  NAND2_X1 U9277 ( .A1(n13053), .A2(n16191), .ZN(n16206) );
  NAND2_X1 U9278 ( .A1(n12884), .A2(n7588), .ZN(n7481) );
  AND2_X1 U9279 ( .A1(n14117), .A2(n14116), .ZN(n7482) );
  AND3_X1 U9280 ( .A1(n8702), .A2(n8678), .A3(SI_9_), .ZN(n7483) );
  OR2_X1 U9281 ( .A1(n15074), .A2(n15322), .ZN(n7484) );
  AND2_X1 U9282 ( .A1(n7964), .A2(n7963), .ZN(n7485) );
  NOR2_X1 U9283 ( .A1(n14763), .A2(n14350), .ZN(n7486) );
  INV_X1 U9284 ( .A(n15668), .ZN(n8102) );
  NAND2_X1 U9285 ( .A1(n9461), .A2(n9460), .ZN(n15732) );
  INV_X1 U9286 ( .A(n15732), .ZN(n8100) );
  INV_X1 U9287 ( .A(n14198), .ZN(n14740) );
  NAND2_X1 U9288 ( .A1(n9054), .A2(n9053), .ZN(n14198) );
  AND2_X1 U9289 ( .A1(n7987), .A2(SI_20_), .ZN(n7487) );
  INV_X1 U9290 ( .A(n11233), .ZN(n7974) );
  INV_X1 U9291 ( .A(n9095), .ZN(n8007) );
  AND2_X1 U9292 ( .A1(n10807), .A2(n10806), .ZN(n12969) );
  AND2_X2 U9293 ( .A1(n14332), .A2(n13997), .ZN(n14040) );
  INV_X2 U9294 ( .A(n14040), .ZN(n14013) );
  NAND2_X2 U9295 ( .A1(n9760), .A2(n9761), .ZN(n9815) );
  NAND2_X2 U9296 ( .A1(n7430), .A2(n7432), .ZN(n9860) );
  INV_X1 U9297 ( .A(n11028), .ZN(n7767) );
  OR2_X1 U9298 ( .A1(n13023), .A2(n16268), .ZN(n7488) );
  NAND2_X1 U9299 ( .A1(n9616), .A2(n8395), .ZN(n7489) );
  NAND4_X1 U9300 ( .A1(n9784), .A2(n9783), .A3(n9782), .A4(n9781), .ZN(n9794)
         );
  NAND2_X1 U9301 ( .A1(n11177), .A2(n11575), .ZN(n11208) );
  NAND2_X1 U9302 ( .A1(n10822), .A2(n14286), .ZN(n7490) );
  NOR2_X1 U9303 ( .A1(n13153), .A2(n10179), .ZN(n7942) );
  NAND2_X1 U9304 ( .A1(n9263), .A2(n13770), .ZN(n9276) );
  INV_X1 U9305 ( .A(n14366), .ZN(n7657) );
  AND2_X1 U9306 ( .A1(n15531), .A2(n8103), .ZN(n7491) );
  INV_X1 U9307 ( .A(n13861), .ZN(n7671) );
  AND2_X1 U9308 ( .A1(n10787), .A2(n10370), .ZN(n7492) );
  NAND2_X1 U9309 ( .A1(n9568), .A2(n15305), .ZN(n7493) );
  AND2_X1 U9310 ( .A1(n12817), .A2(n12816), .ZN(n7494) );
  INV_X1 U9311 ( .A(n9760), .ZN(n7904) );
  AND2_X1 U9312 ( .A1(n13213), .A2(n10099), .ZN(n7495) );
  NOR2_X1 U9313 ( .A1(n9801), .A2(n8500), .ZN(n9825) );
  NAND2_X1 U9314 ( .A1(n11277), .A2(n8355), .ZN(n7496) );
  OR2_X1 U9315 ( .A1(n15137), .A2(n15135), .ZN(n7497) );
  AND2_X1 U9316 ( .A1(n7857), .A2(n7943), .ZN(n9861) );
  NAND2_X1 U9317 ( .A1(n13182), .A2(n12588), .ZN(n13157) );
  AND2_X1 U9318 ( .A1(n15483), .A2(n9672), .ZN(n7498) );
  INV_X1 U9319 ( .A(n7685), .ZN(n14332) );
  XNOR2_X1 U9320 ( .A(n15664), .B(n15303), .ZN(n15463) );
  INV_X1 U9321 ( .A(n15463), .ZN(n8413) );
  NAND2_X1 U9322 ( .A1(n9261), .A2(n15782), .ZN(n15688) );
  INV_X1 U9323 ( .A(n15688), .ZN(n8106) );
  OAI21_X1 U9324 ( .B1(n13211), .B2(n13213), .A(n12700), .ZN(n13200) );
  NAND2_X1 U9325 ( .A1(n7840), .A2(n7842), .ZN(n12913) );
  NAND2_X1 U9326 ( .A1(n10225), .A2(n13108), .ZN(n12718) );
  AND2_X1 U9327 ( .A1(n7633), .A2(n16058), .ZN(n7499) );
  AND2_X1 U9328 ( .A1(n11618), .A2(n11926), .ZN(n7500) );
  OR2_X1 U9329 ( .A1(n10343), .A2(n13109), .ZN(n12581) );
  NAND2_X1 U9330 ( .A1(n11177), .A2(n15038), .ZN(n14863) );
  AND2_X1 U9331 ( .A1(n15715), .A2(n15312), .ZN(n7501) );
  OR2_X1 U9332 ( .A1(n11488), .A2(n7796), .ZN(n7502) );
  INV_X1 U9333 ( .A(n12997), .ZN(n9780) );
  AND2_X1 U9334 ( .A1(n9301), .A2(n13775), .ZN(n9500) );
  AND2_X1 U9335 ( .A1(n8942), .A2(n8941), .ZN(n14551) );
  INV_X1 U9336 ( .A(n14551), .ZN(n14681) );
  OR2_X1 U9337 ( .A1(n9567), .A2(n15306), .ZN(n7503) );
  INV_X1 U9338 ( .A(n14959), .ZN(n8389) );
  AND2_X1 U9339 ( .A1(n12839), .A2(n13126), .ZN(n7504) );
  XNOR2_X1 U9340 ( .A(n15193), .B(n15192), .ZN(n15260) );
  NAND2_X1 U9341 ( .A1(n8650), .A2(n8649), .ZN(n14047) );
  INV_X1 U9342 ( .A(n8539), .ZN(n14326) );
  XNOR2_X1 U9343 ( .A(n8537), .B(n9158), .ZN(n8539) );
  INV_X1 U9344 ( .A(n15181), .ZN(n7887) );
  NAND2_X1 U9345 ( .A1(n8431), .A2(n9497), .ZN(n15600) );
  AND2_X1 U9346 ( .A1(n8240), .A2(n16560), .ZN(n7505) );
  AND2_X1 U9347 ( .A1(n14086), .A2(n14356), .ZN(n7506) );
  OR2_X1 U9348 ( .A1(n14495), .A2(n7958), .ZN(n7507) );
  INV_X1 U9349 ( .A(n15252), .ZN(n15543) );
  OR2_X1 U9350 ( .A1(n11251), .A2(n11250), .ZN(n7508) );
  AND3_X1 U9351 ( .A1(n8579), .A2(n8577), .A3(n8580), .ZN(n7509) );
  INV_X1 U9352 ( .A(n13250), .ZN(n13263) );
  AND2_X1 U9353 ( .A1(n12680), .A2(n12683), .ZN(n13250) );
  AND2_X1 U9354 ( .A1(n14039), .A2(n14038), .ZN(n7510) );
  AND2_X1 U9355 ( .A1(n14054), .A2(n14053), .ZN(n7511) );
  NOR2_X1 U9356 ( .A1(n12217), .A2(n8394), .ZN(n8393) );
  NOR2_X1 U9357 ( .A1(n13022), .A2(n16233), .ZN(n7512) );
  AND2_X1 U9358 ( .A1(n12616), .A2(n12617), .ZN(n12746) );
  AND2_X1 U9359 ( .A1(n14566), .A2(n9133), .ZN(n7513) );
  AND2_X1 U9360 ( .A1(n10223), .A2(n10222), .ZN(n13108) );
  INV_X1 U9361 ( .A(n13108), .ZN(n8270) );
  INV_X1 U9362 ( .A(n8642), .ZN(n8227) );
  AND4_X1 U9363 ( .A1(n9809), .A2(n9808), .A3(n9807), .A4(n9806), .ZN(n16351)
         );
  AND2_X1 U9364 ( .A1(n14026), .A2(n14025), .ZN(n7514) );
  XNOR2_X1 U9365 ( .A(n8680), .B(SI_7_), .ZN(n8677) );
  NAND2_X1 U9366 ( .A1(n14572), .A2(n7966), .ZN(n7967) );
  AND2_X1 U9367 ( .A1(n15181), .A2(n7888), .ZN(n7515) );
  AND2_X1 U9368 ( .A1(n8274), .A2(n12728), .ZN(n7516) );
  OR2_X1 U9369 ( .A1(n15412), .A2(n7799), .ZN(n7517) );
  INV_X1 U9370 ( .A(n12265), .ZN(n8482) );
  AND2_X1 U9371 ( .A1(n16178), .A2(n13031), .ZN(n7518) );
  AND2_X1 U9372 ( .A1(n14094), .A2(n14355), .ZN(n7519) );
  INV_X1 U9373 ( .A(n15093), .ZN(n8471) );
  OR2_X1 U9374 ( .A1(n11660), .A2(n11529), .ZN(n7520) );
  AND2_X1 U9375 ( .A1(n12469), .A2(n12462), .ZN(n7521) );
  AND2_X1 U9376 ( .A1(n7643), .A2(n14801), .ZN(n7522) );
  INV_X1 U9377 ( .A(n9006), .ZN(n8218) );
  INV_X1 U9378 ( .A(n8643), .ZN(n8644) );
  XNOR2_X1 U9379 ( .A(n8646), .B(SI_5_), .ZN(n8643) );
  NAND2_X1 U9380 ( .A1(n8541), .A2(n8532), .ZN(n7523) );
  AND2_X1 U9381 ( .A1(n15555), .A2(n9542), .ZN(n7524) );
  AND2_X1 U9382 ( .A1(n9099), .A2(n9098), .ZN(n14447) );
  INV_X1 U9383 ( .A(n14447), .ZN(n14234) );
  OR2_X1 U9384 ( .A1(n15460), .A2(n15302), .ZN(n7525) );
  NAND2_X1 U9385 ( .A1(n9383), .A2(n9382), .ZN(n15090) );
  AND2_X1 U9386 ( .A1(n7723), .A2(n7720), .ZN(n7526) );
  XNOR2_X1 U9387 ( .A(n8986), .B(SI_22_), .ZN(n9235) );
  AND2_X1 U9388 ( .A1(n14293), .A2(n8641), .ZN(n8225) );
  AND2_X1 U9389 ( .A1(n7947), .A2(n9006), .ZN(n7527) );
  AND2_X1 U9390 ( .A1(n8381), .A2(n8383), .ZN(n7528) );
  INV_X1 U9391 ( .A(n10288), .ZN(n10289) );
  OR2_X1 U9392 ( .A1(n12875), .A2(n13237), .ZN(n12736) );
  NAND2_X1 U9393 ( .A1(n7872), .A2(n7869), .ZN(n7529) );
  INV_X1 U9394 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10414) );
  INV_X1 U9395 ( .A(n8422), .ZN(n8421) );
  NAND2_X1 U9396 ( .A1(n15651), .A2(n9604), .ZN(n8422) );
  NOR2_X1 U9397 ( .A1(n16448), .A2(n11467), .ZN(n7530) );
  NOR2_X1 U9398 ( .A1(n14860), .A2(n14859), .ZN(n7531) );
  NOR2_X1 U9399 ( .A1(n14725), .A2(n14107), .ZN(n7532) );
  NOR2_X1 U9400 ( .A1(n13326), .A2(n12983), .ZN(n7533) );
  AND2_X1 U9401 ( .A1(n7941), .A2(n10178), .ZN(n7534) );
  AND4_X1 U9402 ( .A1(n7649), .A2(n8823), .A3(n8525), .A4(n8526), .ZN(n7535)
         );
  INV_X1 U9403 ( .A(n10239), .ZN(n7915) );
  AND2_X1 U9404 ( .A1(n13113), .A2(n12982), .ZN(n10239) );
  OR2_X1 U9405 ( .A1(n13980), .A2(n13871), .ZN(n7536) );
  AND2_X1 U9406 ( .A1(n8326), .A2(n8329), .ZN(n7537) );
  AND2_X1 U9407 ( .A1(n8664), .A2(SI_6_), .ZN(n7538) );
  AND2_X1 U9408 ( .A1(n8704), .A2(SI_8_), .ZN(n7539) );
  NAND2_X1 U9409 ( .A1(n9510), .A2(n8346), .ZN(n7540) );
  AND2_X1 U9410 ( .A1(n8413), .A2(n8289), .ZN(n7541) );
  OR2_X1 U9411 ( .A1(n7765), .A2(n11891), .ZN(n7542) );
  NOR2_X1 U9412 ( .A1(n14698), .A2(n13901), .ZN(n7543) );
  AND2_X1 U9413 ( .A1(n12138), .A2(n12265), .ZN(n7544) );
  INV_X1 U9414 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9765) );
  OR2_X1 U9415 ( .A1(n7870), .A2(n12969), .ZN(n7545) );
  NAND2_X1 U9416 ( .A1(n12840), .A2(n13108), .ZN(n7546) );
  NOR2_X1 U9417 ( .A1(n14193), .A2(n14482), .ZN(n7547) );
  OAI21_X1 U9418 ( .B1(n14542), .B2(n7467), .A(n7948), .ZN(n8983) );
  INV_X1 U9419 ( .A(n8983), .ZN(n8219) );
  INV_X1 U9420 ( .A(n9873), .ZN(n7908) );
  AND2_X1 U9421 ( .A1(n12044), .A2(n12043), .ZN(n7548) );
  AND2_X1 U9422 ( .A1(n9847), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7549) );
  OR2_X1 U9423 ( .A1(n14073), .A2(n14075), .ZN(n7550) );
  AND2_X1 U9424 ( .A1(n8143), .A2(n12581), .ZN(n7551) );
  AND2_X1 U9425 ( .A1(n7434), .A2(n15258), .ZN(n7552) );
  NAND2_X1 U9426 ( .A1(n8145), .A2(n8144), .ZN(n7553) );
  INV_X1 U9427 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10412) );
  INV_X1 U9428 ( .A(n7873), .ZN(n7872) );
  OAI21_X1 U9429 ( .B1(n7874), .B2(n8497), .A(n7546), .ZN(n7873) );
  OR2_X1 U9430 ( .A1(n15184), .A2(n15182), .ZN(n7554) );
  OR2_X1 U9431 ( .A1(n15106), .A2(n15108), .ZN(n7555) );
  NOR2_X1 U9432 ( .A1(n14740), .A2(n14342), .ZN(n7556) );
  AND2_X1 U9433 ( .A1(n9201), .A2(n9203), .ZN(n7557) );
  AND2_X1 U9434 ( .A1(n14189), .A2(n8304), .ZN(n7558) );
  NAND2_X1 U9435 ( .A1(n12802), .A2(n12801), .ZN(n7559) );
  INV_X1 U9436 ( .A(n15131), .ZN(n7883) );
  OR2_X1 U9437 ( .A1(n10312), .A2(P3_IR_REG_25__SCAN_IN), .ZN(n7560) );
  INV_X1 U9438 ( .A(n8298), .ZN(n8297) );
  NAND2_X1 U9439 ( .A1(n12178), .A2(n9656), .ZN(n8298) );
  INV_X1 U9440 ( .A(n14815), .ZN(n8386) );
  INV_X1 U9441 ( .A(n12194), .ZN(n12752) );
  INV_X1 U9442 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8532) );
  AND3_X1 U9443 ( .A1(n12763), .A2(n12582), .A3(n12572), .ZN(n7561) );
  AND2_X1 U9444 ( .A1(n15151), .A2(n15138), .ZN(n7562) );
  OR2_X1 U9445 ( .A1(n11896), .A2(n11890), .ZN(n7563) );
  NOR3_X1 U9446 ( .A1(n12760), .A2(n13176), .A3(n12759), .ZN(n7564) );
  OR2_X1 U9447 ( .A1(n14058), .A2(n7511), .ZN(n7565) );
  AND2_X1 U9448 ( .A1(n15202), .A2(n15201), .ZN(n15648) );
  INV_X1 U9449 ( .A(n15648), .ZN(n15232) );
  AND2_X1 U9450 ( .A1(n7878), .A2(n7877), .ZN(n7566) );
  AND2_X1 U9451 ( .A1(n8504), .A2(n8301), .ZN(n7567) );
  AND2_X1 U9452 ( .A1(n9606), .A2(n9605), .ZN(n15191) );
  INV_X1 U9453 ( .A(n15191), .ZN(n15193) );
  AND2_X1 U9454 ( .A1(n7960), .A2(n7959), .ZN(n7568) );
  INV_X1 U9455 ( .A(n8415), .ZN(n8414) );
  OAI21_X1 U9456 ( .B1(n15451), .B2(n8423), .A(n7525), .ZN(n8415) );
  OR2_X1 U9457 ( .A1(n10315), .A2(n13843), .ZN(n7569) );
  NAND2_X1 U9458 ( .A1(n14913), .A2(n14912), .ZN(n7570) );
  NAND2_X1 U9459 ( .A1(n12250), .A2(n12249), .ZN(n7571) );
  AND2_X1 U9460 ( .A1(n13120), .A2(n7913), .ZN(n7572) );
  AND2_X1 U9461 ( .A1(n8066), .A2(n8065), .ZN(n7573) );
  AND2_X1 U9462 ( .A1(n15583), .A2(n9529), .ZN(n7574) );
  AND2_X1 U9463 ( .A1(n7789), .A2(n12763), .ZN(n7575) );
  INV_X1 U9464 ( .A(n14462), .ZN(n9065) );
  NAND2_X1 U9465 ( .A1(n9066), .A2(n9064), .ZN(n14462) );
  AND2_X1 U9466 ( .A1(n8090), .A2(n7488), .ZN(n7576) );
  NAND2_X1 U9467 ( .A1(n12583), .A2(n12582), .ZN(n7577) );
  AND2_X1 U9468 ( .A1(n8102), .A2(n8103), .ZN(n7578) );
  AND2_X1 U9469 ( .A1(n14295), .A2(n8660), .ZN(n7579) );
  OR2_X1 U9470 ( .A1(n15077), .A2(n15075), .ZN(n7580) );
  OR2_X1 U9471 ( .A1(n15178), .A2(n15176), .ZN(n7581) );
  AND2_X1 U9472 ( .A1(n11767), .A2(n7484), .ZN(n7582) );
  OR2_X1 U9473 ( .A1(n15089), .A2(n15087), .ZN(n7583) );
  OR2_X1 U9474 ( .A1(n15119), .A2(n15117), .ZN(n7584) );
  AND2_X1 U9475 ( .A1(n8442), .A2(n7493), .ZN(n7585) );
  OR2_X1 U9476 ( .A1(n8474), .A2(n15076), .ZN(n7586) );
  AND2_X1 U9477 ( .A1(n7497), .A2(n7882), .ZN(n7587) );
  OR2_X1 U9478 ( .A1(n7494), .A2(n7825), .ZN(n7588) );
  OR2_X1 U9479 ( .A1(n14119), .A2(n7482), .ZN(n7589) );
  AND2_X1 U9480 ( .A1(n7880), .A2(n8475), .ZN(n7590) );
  INV_X1 U9481 ( .A(n9144), .ZN(n8193) );
  AND2_X1 U9482 ( .A1(n12798), .A2(n12793), .ZN(n7846) );
  AND2_X1 U9483 ( .A1(n7555), .A2(n7894), .ZN(n7591) );
  INV_X1 U9484 ( .A(n8239), .ZN(n8238) );
  NAND2_X1 U9485 ( .A1(n8856), .A2(n8837), .ZN(n8239) );
  AND2_X1 U9486 ( .A1(n9750), .A2(n8496), .ZN(n7592) );
  INV_X1 U9487 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n9790) );
  AND2_X1 U9488 ( .A1(n14933), .A2(n8362), .ZN(n8361) );
  NAND2_X1 U9489 ( .A1(n8996), .A2(n8995), .ZN(n14511) );
  INV_X1 U9490 ( .A(n14511), .ZN(n7963) );
  INV_X1 U9491 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n7746) );
  NAND2_X1 U9492 ( .A1(n13262), .A2(n13250), .ZN(n13265) );
  AND2_X1 U9493 ( .A1(n12539), .A2(n8176), .ZN(n7593) );
  NAND2_X1 U9494 ( .A1(n8382), .A2(n8386), .ZN(n8391) );
  NAND2_X1 U9495 ( .A1(n8524), .A2(n8613), .ZN(n8771) );
  NAND2_X1 U9496 ( .A1(n10198), .A2(n10197), .ZN(n13326) );
  OAI22_X1 U9497 ( .A1(n12527), .A2(P3_D_REG_0__SCAN_IN), .B1(n10332), .B2(
        n11681), .ZN(n10945) );
  OAI21_X1 U9498 ( .B1(n9931), .B2(n7927), .A(n7925), .ZN(n12362) );
  AND2_X1 U9499 ( .A1(n8981), .A2(n8980), .ZN(n14177) );
  OR2_X1 U9500 ( .A1(n9988), .A2(n7736), .ZN(n7594) );
  INV_X1 U9501 ( .A(SI_9_), .ZN(n7999) );
  NAND2_X1 U9502 ( .A1(n10053), .A2(n10052), .ZN(n13249) );
  AND2_X1 U9503 ( .A1(n8842), .A2(n8840), .ZN(n7595) );
  NAND2_X1 U9504 ( .A1(n8133), .A2(n8132), .ZN(n13282) );
  AND2_X1 U9505 ( .A1(n14497), .A2(n13977), .ZN(n7596) );
  OR2_X1 U9506 ( .A1(n10041), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n7597) );
  INV_X1 U9507 ( .A(n15097), .ZN(n8469) );
  INV_X1 U9508 ( .A(n15127), .ZN(n8464) );
  NAND2_X1 U9509 ( .A1(n9592), .A2(n9591), .ZN(n15651) );
  INV_X1 U9510 ( .A(n15651), .ZN(n8114) );
  AND2_X1 U9511 ( .A1(n8293), .A2(n7484), .ZN(n11764) );
  OR2_X1 U9512 ( .A1(n14648), .A2(n14715), .ZN(n7598) );
  NOR2_X1 U9513 ( .A1(n13099), .A2(n13379), .ZN(n7599) );
  NOR2_X1 U9514 ( .A1(n13099), .A2(n13837), .ZN(n7600) );
  AND2_X1 U9515 ( .A1(n14162), .A2(n14161), .ZN(n7601) );
  AND2_X1 U9516 ( .A1(n12035), .A2(n8393), .ZN(n7602) );
  AND2_X1 U9517 ( .A1(n8160), .A2(n8163), .ZN(n7603) );
  INV_X1 U9518 ( .A(n12819), .ZN(n7825) );
  AND3_X1 U9519 ( .A1(n10162), .A2(n10161), .A3(n10160), .ZN(n13188) );
  AND2_X1 U9520 ( .A1(n8920), .A2(n7989), .ZN(n7604) );
  AND2_X1 U9521 ( .A1(n10019), .A2(n12658), .ZN(n7605) );
  NAND2_X1 U9522 ( .A1(n7844), .A2(n7845), .ZN(n12856) );
  AND2_X1 U9523 ( .A1(n9122), .A2(n9121), .ZN(n7606) );
  NAND2_X1 U9524 ( .A1(n9209), .A2(n9208), .ZN(n15668) );
  INV_X1 U9525 ( .A(n8839), .ZN(n8838) );
  INV_X1 U9526 ( .A(n8101), .ZN(n12501) );
  NOR2_X1 U9527 ( .A1(n12494), .A2(n16611), .ZN(n8101) );
  INV_X1 U9528 ( .A(n8511), .ZN(n8380) );
  NOR2_X1 U9529 ( .A1(n14172), .A2(n14430), .ZN(n7607) );
  OR2_X1 U9530 ( .A1(n14164), .A2(n7601), .ZN(n7608) );
  AND2_X1 U9531 ( .A1(n8390), .A2(n8388), .ZN(n7609) );
  AND2_X1 U9532 ( .A1(n10350), .A2(n10349), .ZN(n16605) );
  OR2_X1 U9533 ( .A1(n8492), .A2(n7500), .ZN(n7833) );
  NAND2_X1 U9534 ( .A1(n12137), .A2(n12138), .ZN(n12204) );
  OR2_X1 U9535 ( .A1(n11698), .A2(n12746), .ZN(n11696) );
  NAND2_X1 U9536 ( .A1(n12739), .A2(n9779), .ZN(n16309) );
  AND2_X1 U9537 ( .A1(n9107), .A2(n7962), .ZN(n7610) );
  NAND2_X1 U9538 ( .A1(n8153), .A2(n11154), .ZN(n11237) );
  NAND2_X1 U9539 ( .A1(n8330), .A2(n8613), .ZN(n7611) );
  OAI21_X1 U9540 ( .B1(n7944), .B2(n14299), .A(n7689), .ZN(n11941) );
  NAND2_X1 U9541 ( .A1(n12266), .A2(n12265), .ZN(n12397) );
  INV_X1 U9542 ( .A(n15715), .ZN(n8098) );
  NAND2_X2 U9543 ( .A1(n8809), .A2(n8808), .ZN(n14725) );
  INV_X1 U9544 ( .A(n14725), .ZN(n7968) );
  XNOR2_X1 U9545 ( .A(n9685), .B(n9684), .ZN(n9705) );
  INV_X1 U9546 ( .A(n16568), .ZN(n16599) );
  INV_X1 U9547 ( .A(n16599), .ZN(n16601) );
  NAND2_X1 U9548 ( .A1(n11772), .A2(n8109), .ZN(n7612) );
  INV_X1 U9549 ( .A(n7969), .ZN(n12278) );
  NOR2_X1 U9550 ( .A1(n12089), .A2(n7765), .ZN(n7969) );
  NOR2_X1 U9551 ( .A1(n11652), .A2(n14086), .ZN(n11651) );
  AND2_X1 U9552 ( .A1(n9651), .A2(n9650), .ZN(n7613) );
  AND2_X1 U9553 ( .A1(n7793), .A2(n10132), .ZN(n7614) );
  AND2_X1 U9554 ( .A1(n8073), .A2(n8071), .ZN(n7615) );
  AND2_X1 U9555 ( .A1(n11601), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n7616) );
  AND2_X1 U9556 ( .A1(n11264), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7617) );
  AND2_X1 U9557 ( .A1(n11547), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7618) );
  AND2_X1 U9558 ( .A1(n9070), .A2(SI_27_), .ZN(n7619) );
  AND2_X1 U9559 ( .A1(n11162), .A2(n8660), .ZN(n7620) );
  AND2_X1 U9560 ( .A1(n7972), .A2(n11394), .ZN(n7971) );
  INV_X1 U9561 ( .A(n7971), .ZN(n7662) );
  INV_X1 U9562 ( .A(n12969), .ZN(n7876) );
  INV_X1 U9563 ( .A(n16204), .ZN(n7787) );
  INV_X1 U9564 ( .A(n14041), .ZN(n7957) );
  AND2_X1 U9565 ( .A1(n10397), .A2(n10381), .ZN(n13990) );
  INV_X1 U9566 ( .A(n16448), .ZN(n8096) );
  INV_X1 U9567 ( .A(n11154), .ZN(n7668) );
  XNOR2_X1 U9568 ( .A(n14047), .B(n11311), .ZN(n14293) );
  INV_X1 U9569 ( .A(n14293), .ZN(n8194) );
  AND2_X1 U9570 ( .A1(n10165), .A2(n12191), .ZN(n7621) );
  OR2_X1 U9571 ( .A1(n11242), .A2(n16143), .ZN(n7622) );
  NAND2_X1 U9572 ( .A1(n12773), .A2(n12594), .ZN(n12731) );
  XOR2_X1 U9573 ( .A(n14225), .B(SI_30_), .Z(n7623) );
  NAND2_X1 U9574 ( .A1(n8618), .A2(n8617), .ZN(n14034) );
  INV_X1 U9575 ( .A(n14034), .ZN(n7981) );
  NOR2_X1 U9576 ( .A1(n14227), .A2(n14226), .ZN(n7624) );
  OR2_X1 U9577 ( .A1(n13024), .A2(n16271), .ZN(n7625) );
  AND2_X1 U9578 ( .A1(n8156), .A2(P2_U3088), .ZN(n7626) );
  NOR2_X1 U9579 ( .A1(n10312), .A2(n8148), .ZN(n13841) );
  BUF_X1 U9580 ( .A(n8563), .Z(n14776) );
  INV_X1 U9581 ( .A(P2_RD_REG_SCAN_IN), .ZN(n8402) );
  INV_X1 U9582 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7760) );
  NOR2_X1 U9583 ( .A1(n16287), .A2(n15417), .ZN(n7800) );
  NAND2_X1 U9584 ( .A1(n15413), .A2(n16294), .ZN(n7801) );
  NOR2_X4 U9585 ( .A1(n16522), .A2(n11573), .ZN(n16518) );
  OAI21_X1 U9586 ( .B1(n7629), .B2(n7628), .A(P2_ADDR_REG_12__SCAN_IN), .ZN(
        n8245) );
  INV_X1 U9587 ( .A(n16043), .ZN(n7628) );
  INV_X1 U9588 ( .A(n16106), .ZN(n7632) );
  OAI21_X1 U9589 ( .B1(n16016), .B2(n16017), .A(n7817), .ZN(n7637) );
  INV_X1 U9590 ( .A(n15326), .ZN(n7639) );
  AND2_X1 U9591 ( .A1(n7795), .A2(n7640), .ZN(n7794) );
  INV_X1 U9592 ( .A(n9200), .ZN(n7642) );
  NAND2_X1 U9593 ( .A1(n14797), .A2(n14796), .ZN(n7644) );
  INV_X1 U9594 ( .A(n11794), .ZN(n11792) );
  NAND2_X1 U9595 ( .A1(n12252), .A2(n12251), .ZN(n7645) );
  NAND2_X1 U9596 ( .A1(n7646), .A2(n8392), .ZN(n12252) );
  NAND2_X1 U9597 ( .A1(n11794), .A2(n8393), .ZN(n7646) );
  AOI21_X2 U9598 ( .B1(n14898), .B2(n14899), .A(n8512), .ZN(n14976) );
  NAND2_X1 U9599 ( .A1(n7647), .A2(n11278), .ZN(n11322) );
  NAND2_X1 U9600 ( .A1(n8356), .A2(n8353), .ZN(n7648) );
  NAND2_X1 U9601 ( .A1(n11269), .A2(n11268), .ZN(n8356) );
  INV_X1 U9602 ( .A(n15767), .ZN(n9217) );
  OR2_X4 U9603 ( .A1(n9216), .A2(n15767), .ZN(n9477) );
  AND2_X2 U9604 ( .A1(n8524), .A2(n7535), .ZN(n8330) );
  NAND2_X1 U9605 ( .A1(n7654), .A2(n9120), .ZN(n11647) );
  NAND2_X1 U9606 ( .A1(n12430), .A2(n14304), .ZN(n9128) );
  NAND2_X1 U9607 ( .A1(n12368), .A2(n14305), .ZN(n12367) );
  XNOR2_X2 U9608 ( .A(n16381), .B(n14365), .ZN(n8183) );
  NAND2_X2 U9609 ( .A1(n14583), .A2(n9132), .ZN(n14566) );
  NAND2_X1 U9610 ( .A1(n7659), .A2(n9117), .ZN(n11382) );
  NAND2_X1 U9611 ( .A1(n11408), .A2(n11407), .ZN(n7659) );
  OAI211_X1 U9612 ( .C1(n8153), .C2(n7662), .A(n7663), .B(n11399), .ZN(n11711)
         );
  NAND3_X1 U9613 ( .A1(n8153), .A2(n7667), .A3(n11399), .ZN(n7666) );
  INV_X1 U9614 ( .A(n11399), .ZN(n11402) );
  NAND2_X1 U9615 ( .A1(n13860), .A2(n7671), .ZN(n7669) );
  OAI21_X2 U9616 ( .B1(n13931), .B2(n13932), .A(n7674), .ZN(n13981) );
  OAI21_X2 U9617 ( .B1(n13951), .B2(n7679), .A(n7676), .ZN(n13924) );
  NAND2_X2 U9618 ( .A1(n7685), .A2(n11636), .ZN(n10884) );
  AND2_X2 U9619 ( .A1(n8596), .A2(n8523), .ZN(n8613) );
  NAND3_X1 U9620 ( .A1(n11136), .A2(n11135), .A3(n11141), .ZN(n11219) );
  NAND2_X1 U9621 ( .A1(n10753), .A2(n10752), .ZN(n7811) );
  NAND2_X1 U9622 ( .A1(n14285), .A2(n11344), .ZN(n7688) );
  NAND2_X1 U9623 ( .A1(n8574), .A2(n8573), .ZN(n11344) );
  INV_X2 U9624 ( .A(n11348), .ZN(n16381) );
  AND2_X2 U9625 ( .A1(n8588), .A2(n8587), .ZN(n11348) );
  INV_X1 U9626 ( .A(n14305), .ZN(n7694) );
  NAND3_X1 U9627 ( .A1(n7694), .A2(n8818), .A3(n12284), .ZN(n12375) );
  NAND3_X1 U9628 ( .A1(n7695), .A2(n7950), .A3(n7579), .ZN(n11406) );
  NAND2_X1 U9629 ( .A1(n8621), .A2(n8620), .ZN(n10364) );
  NAND3_X1 U9630 ( .A1(n8242), .A2(n9739), .A3(n8240), .ZN(n7697) );
  NAND3_X1 U9631 ( .A1(n7505), .A2(n9739), .A3(n8242), .ZN(n14647) );
  NAND2_X1 U9632 ( .A1(n7697), .A2(n11936), .ZN(n7696) );
  NAND3_X1 U9633 ( .A1(n7700), .A2(n7699), .A3(n8965), .ZN(n14542) );
  NAND2_X1 U9634 ( .A1(n9797), .A2(n9796), .ZN(n7792) );
  NAND2_X1 U9635 ( .A1(n9785), .A2(n9786), .ZN(n7701) );
  NAND3_X1 U9636 ( .A1(n7706), .A2(n7705), .A3(n7575), .ZN(n7704) );
  NAND2_X1 U9637 ( .A1(n8273), .A2(n7516), .ZN(n7705) );
  NAND2_X1 U9638 ( .A1(n7707), .A2(n7577), .ZN(n7706) );
  NAND2_X1 U9639 ( .A1(n8273), .A2(n8274), .ZN(n7707) );
  INV_X1 U9640 ( .A(n10165), .ZN(n7717) );
  NAND3_X1 U9641 ( .A1(n7719), .A2(n9863), .A3(n7718), .ZN(n9868) );
  NAND3_X1 U9642 ( .A1(n9823), .A2(n7721), .A3(n7720), .ZN(n7719) );
  NAND2_X1 U9643 ( .A1(n10083), .A2(n7730), .ZN(n7728) );
  NAND2_X1 U9644 ( .A1(n10022), .A2(n7743), .ZN(n7740) );
  NAND2_X1 U9645 ( .A1(n7740), .A2(n7741), .ZN(n10056) );
  NAND2_X1 U9646 ( .A1(n10022), .A2(n10021), .ZN(n7742) );
  NAND2_X1 U9647 ( .A1(n10150), .A2(n10149), .ZN(n10154) );
  NAND2_X1 U9648 ( .A1(n10212), .A2(n10211), .ZN(n10229) );
  NAND2_X1 U9649 ( .A1(n12154), .A2(n15246), .ZN(n12153) );
  NAND2_X1 U9650 ( .A1(n9654), .A2(n9653), .ZN(n12001) );
  OR2_X1 U9651 ( .A1(n15195), .A2(n10591), .ZN(n9270) );
  NAND2_X1 U9652 ( .A1(n7813), .A2(n7812), .ZN(n15046) );
  NAND2_X1 U9653 ( .A1(n9681), .A2(n7777), .ZN(n9722) );
  NAND2_X1 U9654 ( .A1(n9722), .A2(n16540), .ZN(n9724) );
  NAND2_X1 U9655 ( .A1(n11048), .A2(n11027), .ZN(n11029) );
  NAND2_X1 U9656 ( .A1(n11101), .A2(n7766), .ZN(n16117) );
  AOI21_X1 U9657 ( .B1(P3_REG1_REG_4__SCAN_IN), .B2(n11113), .A(n11105), .ZN(
        n11250) );
  OAI21_X1 U9658 ( .B1(n8084), .B2(n16235), .A(n8085), .ZN(n16251) );
  NOR2_X1 U9659 ( .A1(n11535), .A2(n11536), .ZN(n11539) );
  NOR2_X1 U9660 ( .A1(n8083), .A2(n11819), .ZN(n11824) );
  NAND3_X1 U9661 ( .A1(n7858), .A2(n9747), .A3(n9748), .ZN(n7856) );
  NAND2_X1 U9662 ( .A1(n11590), .A2(n8128), .ZN(n8127) );
  NAND2_X1 U9663 ( .A1(n7753), .A2(n7750), .ZN(P3_U3487) );
  OR2_X1 U9664 ( .A1(n13388), .A2(n16599), .ZN(n7753) );
  NAND2_X1 U9665 ( .A1(n7756), .A2(n7754), .ZN(P3_U3455) );
  OR2_X1 U9666 ( .A1(n13388), .A2(n16605), .ZN(n7756) );
  NOR2_X1 U9667 ( .A1(n12391), .A2(n8169), .ZN(n8168) );
  XNOR2_X1 U9668 ( .A(n8663), .B(n8661), .ZN(n10447) );
  NAND2_X1 U9669 ( .A1(n8160), .A2(n7607), .ZN(n8159) );
  INV_X1 U9670 ( .A(n8232), .ZN(n8231) );
  OAI21_X1 U9671 ( .B1(n12539), .B2(n8175), .A(n8173), .ZN(n13898) );
  OAI21_X1 U9672 ( .B1(n12427), .B2(n12418), .A(n12425), .ZN(n12539) );
  OAI21_X1 U9673 ( .B1(n16100), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n16099), .ZN(
        n8251) );
  NAND2_X1 U9674 ( .A1(n12564), .A2(n12563), .ZN(n13380) );
  AOI21_X1 U9675 ( .B1(n12729), .B2(n12728), .A(n7761), .ZN(n8273) );
  INV_X1 U9676 ( .A(n12765), .ZN(n7789) );
  NAND2_X1 U9677 ( .A1(n7561), .A2(n7789), .ZN(n7788) );
  OR2_X1 U9678 ( .A1(n14091), .A2(n14090), .ZN(n14098) );
  NAND2_X1 U9679 ( .A1(n8338), .A2(n8339), .ZN(n14168) );
  OAI21_X1 U9680 ( .B1(n14037), .B2(n14036), .A(n7762), .ZN(n8337) );
  NAND2_X1 U9681 ( .A1(n7764), .A2(n7763), .ZN(n7762) );
  NAND2_X1 U9682 ( .A1(n14037), .A2(n14036), .ZN(n7764) );
  OAI211_X1 U9683 ( .C1(n7514), .C2(n14030), .A(n14024), .B(n14023), .ZN(n8343) );
  AOI21_X1 U9684 ( .B1(n14171), .B2(n14170), .A(n14169), .ZN(n14176) );
  NAND2_X1 U9685 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8036) );
  NAND2_X1 U9686 ( .A1(n11022), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n11247) );
  XNOR2_X1 U9687 ( .A(n7816), .B(n7815), .ZN(n13089) );
  NAND2_X1 U9688 ( .A1(n11661), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n11832) );
  NAND2_X1 U9689 ( .A1(n11100), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8039) );
  NAND2_X1 U9690 ( .A1(n16170), .A2(n16169), .ZN(n16168) );
  NAND2_X1 U9691 ( .A1(n11120), .A2(n11020), .ZN(n11043) );
  NAND2_X1 U9692 ( .A1(n11531), .A2(n11530), .ZN(n11659) );
  NOR2_X1 U9693 ( .A1(n11818), .A2(n16527), .ZN(n8083) );
  NAND2_X1 U9694 ( .A1(n7786), .A2(n7785), .ZN(n13056) );
  NOR2_X2 U9695 ( .A1(n16160), .A2(n9944), .ZN(n16159) );
  AOI21_X1 U9696 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n13058), .A(n16240), .ZN(
        n13059) );
  NOR2_X1 U9697 ( .A1(n13057), .A2(n16222), .ZN(n16242) );
  NOR2_X1 U9698 ( .A1(n8121), .A2(n7776), .ZN(n12776) );
  OAI21_X1 U9699 ( .B1(n10351), .B2(n16605), .A(n7770), .ZN(P3_U3456) );
  OAI21_X1 U9700 ( .B1(n10351), .B2(n16599), .A(n7772), .ZN(P3_U3488) );
  NAND2_X1 U9701 ( .A1(n7492), .A2(n10650), .ZN(n10852) );
  NAND3_X2 U9702 ( .A1(n8330), .A2(n8547), .A3(n8613), .ZN(n8551) );
  NAND2_X1 U9703 ( .A1(n7775), .A2(n7598), .ZN(P2_U3527) );
  NAND2_X1 U9704 ( .A1(n14647), .A2(n14646), .ZN(n7775) );
  INV_X1 U9705 ( .A(n9498), .ZN(n8459) );
  XNOR2_X1 U9706 ( .A(n16448), .B(n11467), .ZN(n16434) );
  INV_X1 U9707 ( .A(n9639), .ZN(n7813) );
  NAND2_X1 U9708 ( .A1(n10857), .A2(n8166), .ZN(n10886) );
  XNOR2_X1 U9709 ( .A(n11250), .B(n11251), .ZN(n11031) );
  OAI21_X1 U9710 ( .B1(n13089), .B2(n16274), .A(n13087), .ZN(n8048) );
  NAND2_X2 U9711 ( .A1(n15477), .A2(n7780), .ZN(n15464) );
  NAND2_X2 U9712 ( .A1(n8431), .A2(n8429), .ZN(n15602) );
  NAND2_X1 U9713 ( .A1(n10741), .A2(n7490), .ZN(n10787) );
  INV_X1 U9714 ( .A(n11880), .ZN(n7784) );
  NAND3_X1 U9715 ( .A1(n10886), .A2(n10885), .A3(n10893), .ZN(n10967) );
  NAND2_X1 U9716 ( .A1(n13088), .A2(n16194), .ZN(n8051) );
  NAND2_X1 U9717 ( .A1(n8038), .A2(n8037), .ZN(n11525) );
  NAND2_X1 U9718 ( .A1(n16155), .A2(n13049), .ZN(n16170) );
  NAND2_X1 U9719 ( .A1(n11527), .A2(n11528), .ZN(n11531) );
  NAND2_X1 U9720 ( .A1(n10114), .A2(n11617), .ZN(n10117) );
  NAND2_X1 U9721 ( .A1(n12730), .A2(n12731), .ZN(n8274) );
  INV_X1 U9722 ( .A(n10225), .ZN(n8271) );
  NAND2_X1 U9723 ( .A1(n9953), .A2(n9952), .ZN(n7791) );
  NAND2_X1 U9724 ( .A1(n7792), .A2(n9798), .ZN(n9823) );
  OR2_X1 U9725 ( .A1(n12768), .A2(n12767), .ZN(n8122) );
  NAND2_X1 U9726 ( .A1(n10007), .A2(n10006), .ZN(n10022) );
  NAND2_X2 U9727 ( .A1(n15602), .A2(n9528), .ZN(n15583) );
  NAND2_X1 U9728 ( .A1(n9499), .A2(n7794), .ZN(n9210) );
  AND2_X1 U9729 ( .A1(n9301), .A2(n9201), .ZN(n7795) );
  NAND2_X1 U9730 ( .A1(n9425), .A2(n9424), .ZN(n12165) );
  NAND2_X1 U9731 ( .A1(n7945), .A2(n8718), .ZN(n11630) );
  NAND3_X1 U9732 ( .A1(n8123), .A2(n8122), .A3(n8272), .ZN(n8121) );
  XNOR2_X1 U9733 ( .A(n8723), .B(n8719), .ZN(n10472) );
  NAND2_X1 U9734 ( .A1(n8679), .A2(n7483), .ZN(n7995) );
  INV_X1 U9735 ( .A(n7985), .ZN(n7984) );
  NAND2_X1 U9736 ( .A1(n11233), .A2(n7973), .ZN(n7972) );
  NAND2_X1 U9737 ( .A1(n13123), .A2(n8267), .ZN(n12760) );
  NAND2_X1 U9738 ( .A1(n9868), .A2(n9867), .ZN(n9883) );
  NAND2_X1 U9739 ( .A1(n10003), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n10007) );
  NAND3_X1 U9740 ( .A1(n12576), .A2(n12762), .A3(n12763), .ZN(n7808) );
  NAND2_X1 U9741 ( .A1(n7811), .A2(n8604), .ZN(n10773) );
  AND2_X2 U9742 ( .A1(n15049), .A2(n15046), .ZN(n11988) );
  OR2_X2 U9743 ( .A1(n11539), .A2(n11538), .ZN(n11663) );
  NAND2_X1 U9744 ( .A1(n8051), .A2(n8047), .ZN(P3_U3201) );
  NAND2_X1 U9745 ( .A1(n10852), .A2(n10373), .ZN(n7982) );
  NAND2_X1 U9746 ( .A1(n16065), .A2(n16066), .ZN(n16067) );
  OAI21_X1 U9747 ( .B1(n15983), .B2(n15982), .A(n8248), .ZN(n8247) );
  XNOR2_X1 U9748 ( .A(n8251), .B(n8249), .ZN(SUB_1596_U4) );
  NAND2_X1 U9749 ( .A1(n14450), .A2(n14717), .ZN(n7955) );
  INV_X1 U9750 ( .A(n8204), .ZN(n9727) );
  NAND2_X1 U9751 ( .A1(n15610), .A2(n9662), .ZN(n8431) );
  NAND2_X1 U9752 ( .A1(n8411), .A2(n8414), .ZN(n15436) );
  INV_X1 U9753 ( .A(n12509), .ZN(n8451) );
  OAI21_X1 U9754 ( .B1(n10355), .B2(n9115), .A(n9114), .ZN(n11165) );
  NAND2_X1 U9755 ( .A1(n8187), .A2(n8188), .ZN(n14469) );
  NAND2_X1 U9756 ( .A1(n10775), .A2(n14290), .ZN(n10774) );
  INV_X1 U9757 ( .A(n8701), .ZN(n8702) );
  NAND2_X1 U9758 ( .A1(n13898), .A2(n8178), .ZN(n13951) );
  XNOR2_X1 U9759 ( .A(n11888), .B(n11889), .ZN(n8171) );
  INV_X1 U9760 ( .A(n8140), .ZN(n8139) );
  INV_X1 U9761 ( .A(n12824), .ZN(n7826) );
  NAND2_X1 U9762 ( .A1(n7827), .A2(n7830), .ZN(n12019) );
  NAND3_X1 U9763 ( .A1(n8490), .A2(n11687), .A3(n7833), .ZN(n7827) );
  NAND2_X1 U9764 ( .A1(n11621), .A2(n11620), .ZN(n11688) );
  NAND2_X1 U9765 ( .A1(n7833), .A2(n8490), .ZN(n11621) );
  NAND2_X1 U9766 ( .A1(n12971), .A2(n8510), .ZN(n7836) );
  NAND2_X1 U9767 ( .A1(n12830), .A2(n7843), .ZN(n7842) );
  XNOR2_X1 U9768 ( .A(n12830), .B(n12831), .ZN(n12865) );
  INV_X1 U9769 ( .A(n12831), .ZN(n7843) );
  INV_X1 U9770 ( .A(n12795), .ZN(n7849) );
  NAND2_X1 U9771 ( .A1(n12795), .A2(n7846), .ZN(n7844) );
  NAND3_X1 U9772 ( .A1(n7857), .A2(n7461), .A3(n7852), .ZN(n10071) );
  NAND3_X1 U9773 ( .A1(n7857), .A2(n7461), .A3(n7854), .ZN(n10041) );
  INV_X1 U9774 ( .A(n7859), .ZN(n7861) );
  OAI21_X1 U9775 ( .B1(n12838), .B2(n8499), .A(n8497), .ZN(n12850) );
  NAND2_X1 U9776 ( .A1(n10086), .A2(n7566), .ZN(n10262) );
  NAND2_X1 U9777 ( .A1(n15132), .A2(n7587), .ZN(n7879) );
  NAND2_X1 U9778 ( .A1(n7879), .A2(n7590), .ZN(n15140) );
  NOR2_X2 U9779 ( .A1(n9509), .A2(n7540), .ZN(n9614) );
  NAND2_X1 U9780 ( .A1(n15180), .A2(n7469), .ZN(n7884) );
  NAND2_X1 U9781 ( .A1(n7884), .A2(n7885), .ZN(n15185) );
  NAND3_X1 U9782 ( .A1(n7891), .A2(n9263), .A3(n13770), .ZN(n9288) );
  AND3_X2 U9783 ( .A1(n7891), .A2(n9263), .A3(n7889), .ZN(n9301) );
  NAND2_X1 U9784 ( .A1(n7892), .A2(n7591), .ZN(n8460) );
  NAND3_X1 U9785 ( .A1(n15099), .A2(n7893), .A3(n15100), .ZN(n7892) );
  NAND2_X1 U9786 ( .A1(n15170), .A2(n15171), .ZN(n15169) );
  NAND2_X1 U9787 ( .A1(n7898), .A2(n7899), .ZN(n15092) );
  NAND3_X1 U9788 ( .A1(n15086), .A2(n7583), .A3(n15085), .ZN(n7898) );
  NAND2_X1 U9789 ( .A1(n7900), .A2(n7901), .ZN(n15121) );
  NAND3_X1 U9790 ( .A1(n15116), .A2(n7584), .A3(n15115), .ZN(n7900) );
  OR2_X1 U9791 ( .A1(n9815), .A2(n16321), .ZN(n7902) );
  NAND2_X1 U9792 ( .A1(n9759), .A2(n7902), .ZN(n8118) );
  NAND2_X2 U9793 ( .A1(n9760), .A2(n13854), .ZN(n9817) );
  NAND2_X1 U9794 ( .A1(n10224), .A2(n7912), .ZN(n7911) );
  NAND2_X1 U9795 ( .A1(n10053), .A2(n7917), .ZN(n7916) );
  NAND2_X1 U9796 ( .A1(n7916), .A2(n7919), .ZN(n13223) );
  INV_X1 U9797 ( .A(n7942), .ZN(n7941) );
  NAND3_X1 U9798 ( .A1(n9861), .A2(n8494), .A3(n9749), .ZN(n10312) );
  NAND2_X1 U9799 ( .A1(n11630), .A2(n8738), .ZN(n7944) );
  NAND2_X1 U9800 ( .A1(n11604), .A2(n8717), .ZN(n7945) );
  NAND2_X1 U9801 ( .A1(n8549), .A2(n7952), .ZN(n14773) );
  OR3_X1 U9802 ( .A1(n14495), .A2(n14482), .A3(n14198), .ZN(n14466) );
  NOR2_X1 U9803 ( .A1(n14495), .A2(n14482), .ZN(n14481) );
  NAND2_X1 U9804 ( .A1(n7568), .A2(n9107), .ZN(n11639) );
  NAND2_X1 U9805 ( .A1(n14572), .A2(n7485), .ZN(n14509) );
  INV_X1 U9806 ( .A(n7967), .ZN(n14537) );
  NAND2_X2 U9807 ( .A1(n9149), .A2(n14782), .ZN(n10488) );
  NAND2_X1 U9808 ( .A1(n7976), .A2(n8330), .ZN(n8528) );
  NAND2_X1 U9809 ( .A1(n8914), .A2(n8913), .ZN(n7990) );
  NAND2_X1 U9810 ( .A1(n7990), .A2(n7604), .ZN(n7986) );
  NAND2_X1 U9811 ( .A1(n7988), .A2(n7986), .ZN(n8937) );
  AOI21_X1 U9812 ( .B1(n8914), .B2(n7463), .A(n7487), .ZN(n7988) );
  NAND2_X1 U9813 ( .A1(n7990), .A2(n8920), .ZN(n8938) );
  INV_X1 U9814 ( .A(SI_20_), .ZN(n7989) );
  NAND2_X1 U9815 ( .A1(n8679), .A2(n7992), .ZN(n8000) );
  INV_X1 U9816 ( .A(n8399), .ZN(n7994) );
  NAND2_X1 U9817 ( .A1(n8000), .A2(n8399), .ZN(n8720) );
  NAND2_X1 U9818 ( .A1(n8000), .A2(n7997), .ZN(n7996) );
  NAND2_X1 U9819 ( .A1(n9091), .A2(n7464), .ZN(n8001) );
  NAND2_X1 U9820 ( .A1(n9091), .A2(n9090), .ZN(n9096) );
  NAND2_X1 U9821 ( .A1(n8953), .A2(n8012), .ZN(n8010) );
  NAND2_X1 U9822 ( .A1(n8786), .A2(n8019), .ZN(n8017) );
  OAI21_X1 U9823 ( .B1(n8786), .B2(n8022), .A(n8019), .ZN(n8878) );
  NAND2_X1 U9824 ( .A1(n8017), .A2(n8018), .ZN(n8885) );
  NAND2_X1 U9825 ( .A1(n8786), .A2(n8026), .ZN(n8025) );
  NAND2_X1 U9826 ( .A1(n8786), .A2(n8785), .ZN(n8804) );
  NAND2_X1 U9827 ( .A1(n9032), .A2(n8031), .ZN(n8029) );
  NAND2_X1 U9828 ( .A1(n9032), .A2(n8034), .ZN(n8030) );
  NAND2_X1 U9829 ( .A1(n9032), .A2(n9031), .ZN(n9051) );
  XNOR2_X2 U9830 ( .A(n8036), .B(P3_IR_REG_1__SCAN_IN), .ZN(n13855) );
  NOR2_X4 U9831 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n9789) );
  NAND3_X1 U9832 ( .A1(n11128), .A2(n8056), .A3(n11056), .ZN(n8054) );
  OAI21_X1 U9833 ( .B1(n11128), .B2(n11057), .A(n11056), .ZN(n16123) );
  NAND2_X1 U9834 ( .A1(n16141), .A2(n7573), .ZN(n8060) );
  INV_X1 U9835 ( .A(n16141), .ZN(n8074) );
  NAND2_X1 U9836 ( .A1(n16178), .A2(n8079), .ZN(n8078) );
  OAI211_X1 U9837 ( .C1(n16178), .C2(n16187), .A(n8078), .B(n8080), .ZN(n16198) );
  OR2_X1 U9838 ( .A1(n16272), .A2(n16271), .ZN(n8090) );
  INV_X1 U9839 ( .A(n8090), .ZN(n16270) );
  OAI21_X1 U9840 ( .B1(n9789), .B2(n13843), .A(n9790), .ZN(n8093) );
  NAND3_X1 U9841 ( .A1(n8095), .A2(P3_IR_REG_2__SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n8094) );
  INV_X1 U9842 ( .A(n9789), .ZN(n8095) );
  NAND2_X1 U9843 ( .A1(n7578), .A2(n15531), .ZN(n15482) );
  NAND3_X1 U9844 ( .A1(n8107), .A2(n9626), .A3(n11772), .ZN(n12183) );
  NAND3_X1 U9845 ( .A1(n9626), .A2(n11772), .A3(n8109), .ZN(n12182) );
  NOR2_X1 U9846 ( .A1(n8113), .A2(n15470), .ZN(n15439) );
  NAND4_X1 U9847 ( .A1(n7592), .A2(n8120), .A3(n9752), .A4(n9753), .ZN(n8495)
         );
  NAND2_X1 U9848 ( .A1(n8127), .A2(n8125), .ZN(n11919) );
  INV_X1 U9849 ( .A(n8126), .ZN(n8125) );
  OAI21_X1 U9850 ( .B1(n8130), .B2(n12746), .A(n12745), .ZN(n8126) );
  NAND2_X1 U9851 ( .A1(n13182), .A2(n8131), .ZN(n13160) );
  AOI21_X1 U9852 ( .B1(n13262), .B2(n8137), .A(n8134), .ZN(n13211) );
  OAI21_X1 U9853 ( .B1(n13118), .B2(n8143), .A(n8142), .ZN(n8146) );
  NAND2_X1 U9854 ( .A1(n13118), .A2(n13123), .ZN(n8145) );
  INV_X1 U9855 ( .A(n8146), .ZN(n12573) );
  INV_X1 U9856 ( .A(n10312), .ZN(n8147) );
  NAND2_X1 U9857 ( .A1(n11919), .A2(n10284), .ZN(n11846) );
  NAND2_X1 U9858 ( .A1(n13143), .A2(n13142), .ZN(n13141) );
  OAI21_X1 U9859 ( .B1(n12192), .B2(n12194), .A(n12641), .ZN(n12233) );
  NAND2_X1 U9860 ( .A1(n11870), .A2(n12629), .ZN(n11869) );
  NAND2_X1 U9861 ( .A1(n10281), .A2(n10280), .ZN(n16353) );
  OAI21_X2 U9862 ( .B1(n13131), .B2(n12584), .A(n12714), .ZN(n13118) );
  NAND2_X1 U9863 ( .A1(n11869), .A2(n12631), .ZN(n12122) );
  NAND2_X1 U9864 ( .A1(n10282), .A2(n12740), .ZN(n11731) );
  OAI21_X2 U9865 ( .B1(n13269), .B2(n12668), .A(n12673), .ZN(n13262) );
  NAND2_X1 U9866 ( .A1(n10279), .A2(n12591), .ZN(n16355) );
  OAI21_X2 U9867 ( .B1(n12122), .B2(n12121), .A(n12635), .ZN(n12192) );
  NAND2_X2 U9868 ( .A1(n16314), .A2(n10976), .ZN(n12600) );
  INV_X2 U9869 ( .A(n10419), .ZN(n8155) );
  NAND2_X4 U9870 ( .A1(n9860), .A2(n8155), .ZN(n12569) );
  NAND2_X2 U9871 ( .A1(n8155), .A2(P2_U3088), .ZN(n14783) );
  MUX2_X1 U9872 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n10419), .Z(n8610) );
  MUX2_X1 U9873 ( .A(n10411), .B(n10416), .S(n10419), .Z(n8590) );
  MUX2_X1 U9874 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n8156), .Z(n8646) );
  MUX2_X1 U9875 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n8156), .Z(n8664) );
  MUX2_X1 U9876 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n8156), .Z(n8704) );
  MUX2_X1 U9877 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n8156), .Z(n8680) );
  MUX2_X1 U9878 ( .A(n10545), .B(n10543), .S(n8156), .Z(n8746) );
  MUX2_X1 U9879 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n8156), .Z(n8743) );
  MUX2_X1 U9880 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n8156), .Z(n8719) );
  MUX2_X1 U9881 ( .A(n10701), .B(n9986), .S(n8156), .Z(n8768) );
  MUX2_X1 U9882 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n8156), .Z(n8801) );
  MUX2_X1 U9883 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n8156), .Z(n8839) );
  MUX2_X1 U9884 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n8156), .Z(n8821) );
  MUX2_X1 U9885 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n8156), .Z(n8861) );
  MUX2_X1 U9886 ( .A(n11476), .B(n11474), .S(n8156), .Z(n8876) );
  MUX2_X1 U9887 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n8156), .Z(n8897) );
  MUX2_X1 U9888 ( .A(n11586), .B(n11588), .S(n8156), .Z(n8911) );
  MUX2_X1 U9889 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n8156), .Z(n8954) );
  MUX2_X1 U9890 ( .A(n11707), .B(n11617), .S(n8156), .Z(n8935) );
  MUX2_X1 U9891 ( .A(n12152), .B(n10151), .S(n8156), .Z(n8989) );
  MUX2_X1 U9892 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n8156), .Z(n8987) );
  MUX2_X1 U9893 ( .A(n12191), .B(n10180), .S(n8156), .Z(n9008) );
  MUX2_X1 U9894 ( .A(n12223), .B(n12534), .S(n8156), .Z(n9013) );
  MUX2_X1 U9895 ( .A(n14788), .B(n15778), .S(n8156), .Z(n9047) );
  MUX2_X1 U9896 ( .A(n14784), .B(n15776), .S(n8156), .Z(n9069) );
  MUX2_X1 U9897 ( .A(n10242), .B(n15774), .S(n8156), .Z(n9071) );
  MUX2_X1 U9898 ( .A(n12792), .B(n15771), .S(n8156), .Z(n9092) );
  MUX2_X1 U9899 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n8156), .Z(n14225) );
  MUX2_X1 U9900 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n8156), .Z(n14228) );
  MUX2_X1 U9901 ( .A(n9763), .B(SI_1_), .S(n8155), .Z(n13856) );
  NAND2_X1 U9902 ( .A1(n8968), .A2(n8156), .ZN(n9236) );
  NOR2_X2 U9903 ( .A1(n8159), .A2(n8164), .ZN(n13860) );
  NAND2_X1 U9904 ( .A1(n13924), .A2(n12549), .ZN(n13858) );
  NOR2_X1 U9905 ( .A1(n13857), .A2(n8162), .ZN(n8161) );
  INV_X1 U9906 ( .A(n8164), .ZN(n8163) );
  NAND2_X1 U9907 ( .A1(n10885), .A2(n8167), .ZN(n10382) );
  NAND2_X1 U9908 ( .A1(n10857), .A2(n10377), .ZN(n10383) );
  INV_X1 U9909 ( .A(n12543), .ZN(n8179) );
  NAND2_X1 U9910 ( .A1(n14492), .A2(n8186), .ZN(n8185) );
  OAI21_X2 U9911 ( .B1(n8205), .B2(n9148), .A(n9157), .ZN(n14443) );
  NAND2_X1 U9912 ( .A1(n8624), .A2(n8231), .ZN(n8228) );
  NAND2_X1 U9913 ( .A1(n8228), .A2(n8229), .ZN(n8663) );
  AOI21_X1 U9914 ( .B1(n8239), .B2(n8236), .A(n7486), .ZN(n8234) );
  INV_X1 U9915 ( .A(n8236), .ZN(n8235) );
  NAND2_X1 U9916 ( .A1(n10056), .A2(n8255), .ZN(n8253) );
  INV_X1 U9917 ( .A(n15593), .ZN(n9663) );
  NAND2_X1 U9918 ( .A1(n8293), .A2(n7582), .ZN(n11765) );
  NAND2_X1 U9919 ( .A1(n11955), .A2(n8296), .ZN(n8294) );
  NAND2_X1 U9920 ( .A1(n8294), .A2(n8295), .ZN(n12154) );
  NAND2_X1 U9921 ( .A1(n8300), .A2(n7567), .ZN(n14250) );
  NAND2_X1 U9922 ( .A1(n14176), .A2(n7470), .ZN(n8300) );
  OAI21_X1 U9923 ( .B1(n8313), .B2(n8311), .A(n8310), .ZN(n8309) );
  INV_X1 U9924 ( .A(n14191), .ZN(n8311) );
  AND2_X1 U9925 ( .A1(n8314), .A2(n14191), .ZN(n8312) );
  NAND2_X1 U9926 ( .A1(n14098), .A2(n8319), .ZN(n8318) );
  INV_X1 U9927 ( .A(n14070), .ZN(n8332) );
  INV_X1 U9928 ( .A(n14069), .ZN(n8333) );
  OAI21_X2 U9929 ( .B1(n8337), .B2(n8336), .A(n8335), .ZN(n14051) );
  NAND3_X1 U9930 ( .A1(n14160), .A2(n14159), .A3(n7608), .ZN(n8338) );
  NAND2_X1 U9931 ( .A1(n8340), .A2(n8341), .ZN(n14126) );
  NAND3_X1 U9932 ( .A1(n14115), .A2(n7589), .A3(n14114), .ZN(n8340) );
  NAND2_X1 U9933 ( .A1(n8343), .A2(n8342), .ZN(n14037) );
  NAND3_X1 U9934 ( .A1(n14052), .A2(n7429), .A3(n7565), .ZN(n8344) );
  NAND2_X1 U9935 ( .A1(n8344), .A2(n8345), .ZN(n14064) );
  NAND2_X1 U9936 ( .A1(n8347), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9512) );
  INV_X1 U9937 ( .A(n16399), .ZN(n8349) );
  NAND2_X1 U9938 ( .A1(n8351), .A2(n8348), .ZN(n11321) );
  NAND2_X1 U9939 ( .A1(n8352), .A2(n8353), .ZN(n8351) );
  NAND2_X1 U9940 ( .A1(n14988), .A2(n8361), .ZN(n8357) );
  NOR2_X1 U9941 ( .A1(n14987), .A2(n14854), .ZN(n14932) );
  OAI21_X1 U9942 ( .B1(n14976), .B2(n8373), .A(n8370), .ZN(n14915) );
  OAI21_X1 U9943 ( .B1(n14976), .B2(n8367), .A(n8365), .ZN(n8364) );
  OAI21_X1 U9944 ( .B1(n14976), .B2(n14977), .A(n8369), .ZN(n14950) );
  OAI22_X2 U9945 ( .A1(n14814), .A2(n7528), .B1(n8384), .B2(n8381), .ZN(n14970) );
  NAND2_X1 U9946 ( .A1(n9616), .A2(n9615), .ZN(n9618) );
  NAND2_X1 U9947 ( .A1(n9616), .A2(n8396), .ZN(n9709) );
  INV_X1 U9948 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8404) );
  INV_X1 U9949 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n15421) );
  AOI21_X1 U9950 ( .B1(n15464), .B2(n15463), .A(n8405), .ZN(n15452) );
  NAND3_X1 U9951 ( .A1(n8420), .A2(n8419), .A3(n8416), .ZN(n12788) );
  NAND2_X1 U9952 ( .A1(n8592), .A2(n8591), .ZN(n8424) );
  NAND2_X1 U9953 ( .A1(n8645), .A2(n8427), .ZN(n8426) );
  NAND2_X1 U9954 ( .A1(n15526), .A2(n7585), .ZN(n8435) );
  NAND2_X1 U9955 ( .A1(n8435), .A2(n8434), .ZN(n15479) );
  NAND2_X1 U9956 ( .A1(n8745), .A2(n8744), .ZN(n8750) );
  OAI21_X2 U9957 ( .B1(n15583), .B2(n8448), .A(n8446), .ZN(n15540) );
  NAND2_X2 U9958 ( .A1(n8451), .A2(n15249), .ZN(n15734) );
  NAND2_X1 U9959 ( .A1(n15061), .A2(n15060), .ZN(n8454) );
  NAND2_X1 U9960 ( .A1(n15143), .A2(n8456), .ZN(n8455) );
  NAND2_X1 U9961 ( .A1(n15139), .A2(n7562), .ZN(n8457) );
  NAND3_X1 U9962 ( .A1(n8457), .A2(n8455), .A3(n15163), .ZN(n15165) );
  NAND3_X1 U9963 ( .A1(n9499), .A2(n9301), .A3(n8458), .ZN(n9688) );
  NAND2_X1 U9964 ( .A1(n8460), .A2(n8461), .ZN(n15111) );
  NAND2_X1 U9965 ( .A1(n15121), .A2(n8465), .ZN(n8462) );
  OAI21_X1 U9966 ( .B1(n15121), .B2(n8466), .A(n8465), .ZN(n15126) );
  NAND2_X1 U9967 ( .A1(n8462), .A2(n8463), .ZN(n15125) );
  NAND2_X1 U9968 ( .A1(n15092), .A2(n8470), .ZN(n8467) );
  OAI21_X1 U9969 ( .B1(n15092), .B2(n8472), .A(n8470), .ZN(n15096) );
  NAND2_X1 U9970 ( .A1(n8467), .A2(n8468), .ZN(n15095) );
  NAND3_X1 U9971 ( .A1(n15073), .A2(n15072), .A3(n7580), .ZN(n8473) );
  NAND2_X1 U9972 ( .A1(n8473), .A2(n7586), .ZN(n15081) );
  NAND3_X1 U9973 ( .A1(n15175), .A2(n15174), .A3(n7581), .ZN(n8476) );
  NAND2_X1 U9974 ( .A1(n8476), .A2(n8477), .ZN(n15180) );
  NAND2_X1 U9975 ( .A1(n9202), .A2(n8478), .ZN(n15761) );
  NAND2_X1 U9976 ( .A1(n8479), .A2(n8480), .ZN(n12400) );
  NAND2_X1 U9977 ( .A1(n12137), .A2(n7544), .ZN(n8479) );
  NAND2_X1 U9978 ( .A1(n12898), .A2(n8484), .ZN(n8483) );
  NAND2_X1 U9979 ( .A1(n11298), .A2(n8491), .ZN(n8490) );
  INV_X1 U9980 ( .A(n8493), .ZN(n11619) );
  NOR2_X1 U9981 ( .A1(n10041), .A2(n8495), .ZN(n10315) );
  NAND2_X1 U9982 ( .A1(n12838), .A2(n12837), .ZN(n12962) );
  NAND2_X1 U9983 ( .A1(n9767), .A2(n9768), .ZN(n9764) );
  INV_X1 U9984 ( .A(n9705), .ZN(n9706) );
  NAND2_X1 U9985 ( .A1(n14129), .A2(n14128), .ZN(n14136) );
  OR2_X1 U9986 ( .A1(n14009), .A2(n14008), .ZN(n14020) );
  INV_X1 U9987 ( .A(n7431), .ZN(n14424) );
  OR2_X1 U9988 ( .A1(n14218), .A2(n10534), .ZN(n8570) );
  NAND2_X1 U9989 ( .A1(n16331), .A2(n15045), .ZN(n15041) );
  NAND2_X1 U9990 ( .A1(n10278), .A2(n10813), .ZN(n16308) );
  AND3_X1 U9991 ( .A1(n15229), .A2(n15228), .A3(n15227), .ZN(n15291) );
  OR2_X1 U9992 ( .A1(n15446), .A2(n15445), .ZN(n15652) );
  OR2_X1 U9993 ( .A1(n9311), .A2(n11992), .ZN(n9272) );
  OR2_X1 U9994 ( .A1(n9311), .A2(n11579), .ZN(n9250) );
  OR2_X1 U9995 ( .A1(n7814), .A2(n15440), .ZN(n9600) );
  OR2_X1 U9996 ( .A1(n7814), .A2(n15455), .ZN(n9588) );
  NOR2_X1 U9997 ( .A1(n14217), .A2(n14216), .ZN(n8504) );
  INV_X1 U9998 ( .A(n14304), .ZN(n8856) );
  NOR2_X1 U9999 ( .A1(n15308), .A2(n15211), .ZN(n8506) );
  NOR2_X1 U10000 ( .A1(n15659), .A2(n15302), .ZN(n8507) );
  OR2_X1 U10001 ( .A1(n14270), .A2(n14269), .ZN(n8508) );
  NAND2_X1 U10002 ( .A1(n14240), .A2(n14239), .ZN(n8509) );
  OR2_X1 U10003 ( .A1(n12806), .A2(n13274), .ZN(n8510) );
  AND2_X1 U10004 ( .A1(n14885), .A2(n14884), .ZN(n8511) );
  AND2_X1 U10005 ( .A1(n14873), .A2(n14872), .ZN(n8512) );
  OR2_X1 U10006 ( .A1(n8838), .A2(n10465), .ZN(n8513) );
  AND2_X1 U10007 ( .A1(n8785), .A2(n8770), .ZN(n8514) );
  INV_X2 U10008 ( .A(n16559), .ZN(n16560) );
  AND2_X1 U10009 ( .A1(n10493), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15875) );
  INV_X1 U10010 ( .A(n14768), .ZN(n9744) );
  NAND2_X1 U10011 ( .A1(n14242), .A2(n14241), .ZN(n8515) );
  INV_X1 U10012 ( .A(n15559), .ZN(n9667) );
  AND2_X1 U10013 ( .A1(n14278), .A2(n14257), .ZN(n9148) );
  INV_X1 U10014 ( .A(n14094), .ZN(n9108) );
  INV_X1 U10015 ( .A(n7437), .ZN(n14430) );
  AND2_X1 U10016 ( .A1(n13096), .A2(n16597), .ZN(n8516) );
  INV_X1 U10017 ( .A(n13213), .ZN(n13210) );
  INV_X1 U10018 ( .A(n13310), .ZN(n16369) );
  INV_X1 U10019 ( .A(n13292), .ZN(n13307) );
  NAND2_X1 U10020 ( .A1(n15710), .A2(n15311), .ZN(n8517) );
  INV_X1 U10021 ( .A(n14698), .ZN(n9109) );
  OR2_X1 U10022 ( .A1(n15161), .A2(n15688), .ZN(n8518) );
  OR2_X1 U10023 ( .A1(n13862), .A2(n7671), .ZN(n8519) );
  INV_X1 U10024 ( .A(n14541), .ZN(n8965) );
  NAND2_X1 U10025 ( .A1(n9721), .A2(n9720), .ZN(n16580) );
  NAND2_X1 U10026 ( .A1(n9721), .A2(n11567), .ZN(n16579) );
  INV_X1 U10027 ( .A(n12665), .ZN(n10287) );
  NOR2_X1 U10028 ( .A1(n13176), .A2(n12585), .ZN(n8520) );
  INV_X1 U10029 ( .A(n15090), .ZN(n9626) );
  INV_X1 U10030 ( .A(n15238), .ZN(n9333) );
  INV_X1 U10031 ( .A(n15063), .ZN(n15064) );
  AOI21_X1 U10032 ( .B1(n14009), .B2(n14008), .A(n14007), .ZN(n14017) );
  INV_X1 U10033 ( .A(n14079), .ZN(n14080) );
  AND2_X1 U10034 ( .A1(n15162), .A2(n8518), .ZN(n15163) );
  NAND2_X1 U10035 ( .A1(n14141), .A2(n14140), .ZN(n14146) );
  INV_X1 U10036 ( .A(n15177), .ZN(n15178) );
  NAND2_X1 U10037 ( .A1(n8515), .A2(n8509), .ZN(n14217) );
  INV_X1 U10038 ( .A(n14263), .ZN(n14237) );
  AND3_X1 U10039 ( .A1(n9194), .A2(n13793), .A3(n13789), .ZN(n9195) );
  INV_X1 U10040 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n9746) );
  INV_X1 U10041 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8525) );
  INV_X1 U10042 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n13775) );
  OR2_X1 U10043 ( .A1(n13164), .A2(n12832), .ZN(n10178) );
  INV_X1 U10044 ( .A(n16351), .ZN(n9810) );
  AND2_X1 U10045 ( .A1(n14247), .A2(n14246), .ZN(n14248) );
  INV_X1 U10046 ( .A(n12275), .ZN(n9124) );
  OAI21_X1 U10047 ( .B1(n11208), .B2(n16327), .A(n11181), .ZN(n11182) );
  INV_X1 U10048 ( .A(n16339), .ZN(n9268) );
  INV_X1 U10049 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n13793) );
  XNOR2_X1 U10050 ( .A(n11681), .B(n13506), .ZN(n10319) );
  INV_X1 U10051 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9957) );
  XOR2_X1 U10052 ( .A(n14338), .B(n14435), .Z(n14318) );
  AND2_X1 U10053 ( .A1(n9021), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9035) );
  OR2_X1 U10054 ( .A1(n8974), .A2(n8973), .ZN(n8999) );
  INV_X1 U10055 ( .A(n8731), .ZN(n8729) );
  NAND2_X1 U10056 ( .A1(n13994), .A2(n14001), .ZN(n14000) );
  OAI22_X1 U10057 ( .A1(n9269), .A2(n14863), .B1(n11208), .B2(n16339), .ZN(
        n11176) );
  INV_X1 U10058 ( .A(n11182), .ZN(n11183) );
  NOR2_X1 U10059 ( .A1(n9518), .A2(n9517), .ZN(n9516) );
  NAND2_X1 U10060 ( .A1(n15783), .A2(n9714), .ZN(n15033) );
  NOR2_X1 U10061 ( .A1(n9371), .A2(n9370), .ZN(n9369) );
  INV_X1 U10062 ( .A(n8677), .ZN(n8678) );
  NOR2_X2 U10063 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9263) );
  INV_X1 U10064 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n13460) );
  AND2_X1 U10065 ( .A1(n9958), .A2(n9957), .ZN(n9977) );
  INV_X1 U10066 ( .A(n9939), .ZN(n9940) );
  NAND2_X1 U10067 ( .A1(n10444), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9863) );
  OR2_X1 U10068 ( .A1(n12537), .A2(n12536), .ZN(n12538) );
  INV_X1 U10069 ( .A(n9079), .ZN(n9081) );
  OR2_X1 U10070 ( .A1(n8943), .A2(n13926), .ZN(n8958) );
  INV_X1 U10071 ( .A(n12791), .ZN(n8562) );
  NAND2_X1 U10072 ( .A1(n8869), .A2(n8868), .ZN(n8889) );
  NAND2_X1 U10073 ( .A1(n8729), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8759) );
  AND2_X1 U10074 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8632) );
  OR2_X1 U10075 ( .A1(n9174), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n9160) );
  CLKBUF_X3 U10076 ( .A(n11755), .Z(n14916) );
  NAND2_X1 U10077 ( .A1(n9547), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9237) );
  NAND2_X1 U10078 ( .A1(n9218), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9572) );
  INV_X1 U10079 ( .A(n9237), .ZN(n9560) );
  OR2_X1 U10080 ( .A1(n9490), .A2(n9489), .ZN(n9505) );
  OR2_X1 U10081 ( .A1(n9401), .A2(n9400), .ZN(n9417) );
  NAND2_X1 U10082 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n9573), .ZN(n9584) );
  NAND2_X1 U10083 ( .A1(n9636), .A2(n16339), .ZN(n15044) );
  NOR2_X1 U10084 ( .A1(n15101), .A2(n12183), .ZN(n12291) );
  NAND2_X1 U10085 ( .A1(n8821), .A2(SI_15_), .ZN(n8842) );
  NAND2_X1 U10086 ( .A1(n8766), .A2(n8748), .ZN(n8749) );
  NOR2_X1 U10087 ( .A1(n16038), .A2(n16037), .ZN(n16039) );
  OR2_X1 U10088 ( .A1(n13838), .A2(n10353), .ZN(n10989) );
  AND2_X1 U10089 ( .A1(n11085), .A2(n11086), .ZN(n11083) );
  INV_X1 U10090 ( .A(n9815), .ZN(n10247) );
  NAND2_X1 U10091 ( .A1(n13141), .A2(n12711), .ZN(n13131) );
  NAND2_X1 U10092 ( .A1(n11081), .A2(n16351), .ZN(n12608) );
  INV_X1 U10093 ( .A(n10343), .ZN(n13099) );
  AND2_X1 U10094 ( .A1(n10305), .A2(n10336), .ZN(n16541) );
  INV_X1 U10095 ( .A(n11220), .ZN(n11141) );
  NAND2_X1 U10096 ( .A1(n13943), .A2(n13942), .ZN(n13931) );
  INV_X1 U10097 ( .A(n14279), .ZN(n14280) );
  AND2_X1 U10098 ( .A1(n9081), .A2(n9057), .ZN(n14467) );
  OR2_X1 U10099 ( .A1(n8889), .A2(n13969), .ZN(n8926) );
  INV_X1 U10100 ( .A(n10493), .ZN(n10492) );
  AND2_X1 U10101 ( .A1(n10492), .A2(n14779), .ZN(n10511) );
  INV_X1 U10102 ( .A(n14313), .ZN(n14478) );
  INV_X1 U10103 ( .A(n14567), .ZN(n14563) );
  NAND2_X1 U10104 ( .A1(n11651), .A2(n9108), .ZN(n12089) );
  INV_X1 U10105 ( .A(n11651), .ZN(n11947) );
  AOI21_X1 U10106 ( .B1(n9165), .B2(n9161), .A(n14772), .ZN(n9166) );
  AND2_X1 U10107 ( .A1(n9545), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9547) );
  OR2_X1 U10108 ( .A1(n9505), .A2(n9504), .ZN(n9518) );
  OR2_X1 U10109 ( .A1(n9477), .A2(n9255), .ZN(n9258) );
  OR2_X1 U10110 ( .A1(n10929), .A2(n10928), .ZN(n10926) );
  INV_X1 U10111 ( .A(n15243), .ZN(n12178) );
  INV_X1 U10112 ( .A(n16490), .ZN(n16508) );
  NOR2_X1 U10113 ( .A1(n12778), .A2(n9635), .ZN(n9682) );
  OAI21_X1 U10114 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n16062), .A(n16061), 
        .ZN(n16070) );
  INV_X1 U10115 ( .A(n13187), .ZN(n12945) );
  INV_X1 U10116 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n9849) );
  AND2_X1 U10117 ( .A1(n11032), .A2(n11017), .ZN(n16194) );
  INV_X1 U10118 ( .A(n16350), .ZN(n12975) );
  NAND2_X1 U10119 ( .A1(n11450), .A2(n16360), .ZN(n13310) );
  NAND2_X1 U10120 ( .A1(n10299), .A2(n11377), .ZN(n16593) );
  NAND2_X1 U10121 ( .A1(n16541), .A2(n16584), .ZN(n16597) );
  OAI21_X1 U10122 ( .B1(n12527), .B2(P3_D_REG_1__SCAN_IN), .A(n10333), .ZN(
        n11443) );
  XNOR2_X1 U10123 ( .A(n9766), .B(n9765), .ZN(n10269) );
  AND2_X1 U10124 ( .A1(n10491), .A2(n10490), .ZN(n10493) );
  OR2_X1 U10125 ( .A1(n13912), .A2(n9039), .ZN(n9087) );
  INV_X1 U10126 ( .A(n15830), .ZN(n15873) );
  AND2_X1 U10127 ( .A1(n10511), .A2(n14325), .ZN(n15877) );
  AND2_X1 U10128 ( .A1(n10487), .A2(n9150), .ZN(n14588) );
  INV_X1 U10129 ( .A(n14619), .ZN(n14628) );
  INV_X1 U10130 ( .A(n14717), .ZN(n16386) );
  NOR2_X1 U10131 ( .A1(n13996), .A2(n14323), .ZN(n16558) );
  AND3_X1 U10132 ( .A1(n15817), .A2(n10358), .A3(n9187), .ZN(n9726) );
  NAND2_X1 U10133 ( .A1(n8533), .A2(n8532), .ZN(n8534) );
  AND2_X1 U10134 ( .A1(n9245), .A2(n9244), .ZN(n15146) );
  INV_X1 U10135 ( .A(n16285), .ZN(n15415) );
  OR2_X1 U10136 ( .A1(n11572), .A2(n12118), .ZN(n10585) );
  INV_X1 U10137 ( .A(n15256), .ZN(n15451) );
  INV_X1 U10138 ( .A(n15249), .ZN(n12510) );
  INV_X1 U10139 ( .A(n16512), .ZN(n15619) );
  AND2_X1 U10140 ( .A1(n9717), .A2(n15759), .ZN(n11567) );
  INV_X1 U10141 ( .A(n16536), .ZN(n16479) );
  AND2_X1 U10142 ( .A1(n16370), .A2(n16468), .ZN(n16576) );
  INV_X1 U10143 ( .A(n16576), .ZN(n16443) );
  NOR2_X1 U10144 ( .A1(n11174), .A2(n9715), .ZN(n9721) );
  AND2_X1 U10145 ( .A1(n11177), .A2(n10467), .ZN(n11572) );
  AND2_X1 U10146 ( .A1(n11035), .A2(n11034), .ZN(n16259) );
  INV_X1 U10147 ( .A(n12978), .ZN(n12955) );
  INV_X1 U10148 ( .A(n12966), .ZN(n12981) );
  INV_X1 U10149 ( .A(n13126), .ZN(n12983) );
  INV_X1 U10150 ( .A(n13237), .ZN(n12987) );
  INV_X1 U10151 ( .A(n16269), .ZN(n16142) );
  INV_X1 U10152 ( .A(n13310), .ZN(n13292) );
  NAND2_X1 U10153 ( .A1(n13307), .A2(n16367), .ZN(n13313) );
  NAND2_X1 U10154 ( .A1(n16601), .A2(n16544), .ZN(n13379) );
  INV_X2 U10155 ( .A(n16605), .ZN(n16602) );
  OR2_X1 U10156 ( .A1(n12528), .A2(n13838), .ZN(n12530) );
  NAND2_X1 U10157 ( .A1(n10987), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13838) );
  INV_X1 U10158 ( .A(SI_13_), .ZN(n13629) );
  INV_X1 U10159 ( .A(SI_12_), .ZN(n13436) );
  INV_X1 U10160 ( .A(n13990), .ZN(n13963) );
  INV_X1 U10161 ( .A(n14236), .ZN(n14340) );
  INV_X1 U10162 ( .A(n14177), .ZN(n14346) );
  OR2_X1 U10163 ( .A1(n15869), .A2(P2_U3088), .ZN(n15842) );
  INV_X1 U10164 ( .A(n15877), .ZN(n15848) );
  NAND2_X1 U10165 ( .A1(n14431), .A2(n14430), .ZN(n14638) );
  AND2_X2 U10166 ( .A1(n10359), .A2(n14624), .ZN(n14622) );
  INV_X1 U10167 ( .A(n14630), .ZN(n14580) );
  NAND2_X1 U10168 ( .A1(n16560), .A2(n16382), .ZN(n14715) );
  NAND2_X1 U10169 ( .A1(n9726), .A2(n10385), .ZN(n16559) );
  AOI21_X1 U10170 ( .B1(n14193), .B2(n9744), .A(n9743), .ZN(n9745) );
  INV_X1 U10171 ( .A(n14122), .ZN(n14769) );
  NAND2_X1 U10172 ( .A1(n9726), .A2(n9725), .ZN(n16561) );
  OR2_X1 U10173 ( .A1(n15822), .A2(n15819), .ZN(n15820) );
  OR2_X1 U10174 ( .A1(n10390), .A2(P2_U3088), .ZN(n15822) );
  INV_X1 U10175 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10545) );
  NAND2_X1 U10176 ( .A1(n11190), .A2(n11189), .ZN(n15029) );
  OR3_X1 U10177 ( .A1(n9483), .A2(n9482), .A3(n9481), .ZN(n15313) );
  INV_X1 U10178 ( .A(n16287), .ZN(n15928) );
  OR2_X1 U10179 ( .A1(n16522), .A2(n12057), .ZN(n15592) );
  INV_X1 U10180 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11474) );
  INV_X1 U10181 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10543) );
  INV_X1 U10182 ( .A(n12998), .ZN(P3_U3897) );
  INV_X1 U10183 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8527) );
  NAND2_X1 U10184 ( .A1(n8536), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U10185 ( .A1(n8886), .A2(n8527), .ZN(n8529) );
  NAND2_X1 U10186 ( .A1(n8538), .A2(n8541), .ZN(n8531) );
  INV_X1 U10187 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9158) );
  NAND2_X1 U10188 ( .A1(n8539), .A2(n7431), .ZN(n13996) );
  INV_X1 U10189 ( .A(n16558), .ZN(n10825) );
  NAND2_X1 U10190 ( .A1(n11636), .A2(n10825), .ZN(n14717) );
  NOR2_X1 U10191 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n8543) );
  NOR2_X1 U10192 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .ZN(n8542) );
  INV_X1 U10193 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8540) );
  NAND4_X1 U10194 ( .A1(n8543), .A2(n8542), .A3(n8541), .A4(n8540), .ZN(n8546)
         );
  INV_X1 U10195 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9162) );
  NAND4_X1 U10196 ( .A1(n8544), .A2(n8527), .A3(n8532), .A4(n9162), .ZN(n8545)
         );
  NOR2_X1 U10197 ( .A1(n8546), .A2(n8545), .ZN(n8547) );
  INV_X1 U10198 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8548) );
  INV_X1 U10199 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8550) );
  NAND2_X1 U10200 ( .A1(n8551), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8552) );
  INV_X1 U10201 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8554) );
  NAND2_X1 U10202 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8553) );
  XNOR2_X1 U10203 ( .A(n8554), .B(n8553), .ZN(n10498) );
  OR2_X1 U10204 ( .A1(n8921), .A2(n10412), .ZN(n8557) );
  AND2_X1 U10205 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8555) );
  NAND2_X1 U10206 ( .A1(n10419), .A2(n8555), .ZN(n9253) );
  OAI21_X1 U10207 ( .B1(n10420), .B2(n9762), .A(n9253), .ZN(n8584) );
  XNOR2_X1 U10208 ( .A(n8585), .B(n8584), .ZN(n10413) );
  OR2_X1 U10209 ( .A1(n8586), .A2(n10413), .ZN(n8556) );
  OAI211_X2 U10210 ( .C1(n10488), .C2(n10498), .A(n8557), .B(n8556), .ZN(
        n14006) );
  INV_X1 U10211 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8558) );
  INV_X1 U10212 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8559) );
  AND2_X4 U10213 ( .A1(n12791), .A2(n14776), .ZN(n8599) );
  NAND2_X1 U10214 ( .A1(n8599), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8568) );
  INV_X1 U10215 ( .A(n8563), .ZN(n8561) );
  INV_X1 U10216 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11370) );
  NAND2_X1 U10217 ( .A1(n8561), .A2(n8562), .ZN(n8575) );
  INV_X1 U10218 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11364) );
  OR2_X1 U10219 ( .A1(n8575), .A2(n11364), .ZN(n8566) );
  INV_X1 U10220 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n8564) );
  NAND2_X1 U10221 ( .A1(n8599), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8572) );
  INV_X1 U10222 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10937) );
  OR2_X1 U10223 ( .A1(n8575), .A2(n10937), .ZN(n8571) );
  INV_X1 U10224 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10534) );
  INV_X1 U10225 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10940) );
  NAND4_X2 U10226 ( .A1(n8572), .A2(n8569), .A3(n8570), .A4(n8571), .ZN(n13994) );
  INV_X1 U10227 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n14374) );
  XNOR2_X1 U10228 ( .A(n9762), .B(n10420), .ZN(n14791) );
  MUX2_X1 U10229 ( .A(n14374), .B(n14791), .S(n10488), .Z(n14001) );
  INV_X1 U10230 ( .A(n14001), .ZN(n10743) );
  NAND2_X1 U10231 ( .A1(n13994), .A2(n10743), .ZN(n10369) );
  NAND2_X1 U10232 ( .A1(n14287), .A2(n10369), .ZN(n8574) );
  NAND2_X1 U10233 ( .A1(n7657), .A2(n11365), .ZN(n8573) );
  NAND2_X1 U10234 ( .A1(n8599), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8580) );
  INV_X1 U10235 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11353) );
  INV_X1 U10236 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11347) );
  OR2_X1 U10237 ( .A1(n9039), .A2(n11347), .ZN(n8578) );
  INV_X1 U10238 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n8576) );
  INV_X2 U10239 ( .A(n8921), .ZN(n8902) );
  INV_X2 U10240 ( .A(n10488), .ZN(n8901) );
  OR2_X1 U10241 ( .A1(n8581), .A2(n14772), .ZN(n8582) );
  XNOR2_X1 U10242 ( .A(n8582), .B(P2_IR_REG_2__SCAN_IN), .ZN(n14385) );
  AOI22_X1 U10243 ( .A1(n8902), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n8901), .B2(
        n14385), .ZN(n8588) );
  AOI21_X2 U10244 ( .B1(n8585), .B2(n8584), .A(n8583), .ZN(n8593) );
  XNOR2_X1 U10245 ( .A(n8592), .B(n8590), .ZN(n10409) );
  NAND2_X1 U10246 ( .A1(n10409), .A2(n8612), .ZN(n8587) );
  INV_X1 U10247 ( .A(n14365), .ZN(n10648) );
  NAND2_X1 U10248 ( .A1(n10648), .A2(n11348), .ZN(n8589) );
  INV_X1 U10249 ( .A(n8590), .ZN(n8591) );
  INV_X1 U10250 ( .A(n8593), .ZN(n8594) );
  NAND2_X1 U10251 ( .A1(n8594), .A2(SI_2_), .ZN(n8595) );
  OR2_X1 U10252 ( .A1(n8596), .A2(n14772), .ZN(n8597) );
  XNOR2_X1 U10253 ( .A(n8597), .B(P2_IR_REG_3__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U10254 ( .A1(n8902), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8901), .B2(
        n10499), .ZN(n8598) );
  NAND2_X1 U10255 ( .A1(n8599), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8603) );
  INV_X1 U10256 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10481) );
  OR2_X1 U10257 ( .A1(n8831), .A2(n10481), .ZN(n8602) );
  OR2_X1 U10258 ( .A1(n8575), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8601) );
  INV_X1 U10259 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10500) );
  OR2_X1 U10260 ( .A1(n14218), .A2(n10500), .ZN(n8600) );
  NAND4_X1 U10261 ( .A1(n8603), .A2(n8602), .A3(n8601), .A4(n8600), .ZN(n14364) );
  OR2_X1 U10262 ( .A1(n14364), .A2(n14027), .ZN(n8604) );
  NAND2_X1 U10263 ( .A1(n8599), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8608) );
  INV_X1 U10264 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11360) );
  OR2_X1 U10265 ( .A1(n8831), .A2(n11360), .ZN(n8607) );
  XNOR2_X1 U10266 ( .A(P2_REG3_REG_3__SCAN_IN), .B(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n11356) );
  OR2_X1 U10267 ( .A1(n9039), .A2(n11356), .ZN(n8606) );
  INV_X1 U10268 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10501) );
  OR2_X1 U10269 ( .A1(n8851), .A2(n10501), .ZN(n8605) );
  NAND4_X1 U10270 ( .A1(n8608), .A2(n8607), .A3(n8606), .A4(n8605), .ZN(n14363) );
  NAND2_X1 U10271 ( .A1(n8610), .A2(SI_3_), .ZN(n8611) );
  XNOR2_X1 U10272 ( .A(n8624), .B(n8622), .ZN(n10417) );
  NAND2_X1 U10273 ( .A1(n10417), .A2(n8612), .ZN(n8618) );
  NOR2_X1 U10274 ( .A1(n8613), .A2(n14772), .ZN(n8614) );
  MUX2_X1 U10275 ( .A(n14772), .B(n8614), .S(P2_IR_REG_4__SCAN_IN), .Z(n8616)
         );
  INV_X1 U10276 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8615) );
  NOR2_X1 U10277 ( .A1(n8616), .A2(n8627), .ZN(n14401) );
  AOI22_X1 U10278 ( .A1(n8902), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8901), .B2(
        n14401), .ZN(n8617) );
  INV_X1 U10279 ( .A(n14290), .ZN(n8619) );
  NAND2_X1 U10280 ( .A1(n10773), .A2(n8619), .ZN(n8621) );
  OR2_X1 U10281 ( .A1(n14034), .A2(n14363), .ZN(n8620) );
  NAND2_X1 U10282 ( .A1(n8625), .A2(SI_4_), .ZN(n8626) );
  XNOR2_X1 U10283 ( .A(n8645), .B(n8643), .ZN(n10443) );
  NAND2_X1 U10284 ( .A1(n10443), .A2(n8612), .ZN(n8630) );
  NAND2_X1 U10285 ( .A1(n8647), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8628) );
  XNOR2_X1 U10286 ( .A(n8628), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U10287 ( .A1(n8902), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8901), .B2(
        n10503), .ZN(n8629) );
  NAND2_X1 U10288 ( .A1(n8630), .A2(n8629), .ZN(n14041) );
  NAND2_X1 U10289 ( .A1(n8599), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8640) );
  INV_X1 U10290 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n8631) );
  OR2_X1 U10291 ( .A1(n8831), .A2(n8631), .ZN(n8639) );
  NAND2_X1 U10292 ( .A1(n8632), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8654) );
  INV_X1 U10293 ( .A(n8632), .ZN(n8634) );
  INV_X1 U10294 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8633) );
  NAND2_X1 U10295 ( .A1(n8634), .A2(n8633), .ZN(n8635) );
  NAND2_X1 U10296 ( .A1(n8654), .A2(n8635), .ZN(n10965) );
  OR2_X1 U10297 ( .A1(n9039), .A2(n10965), .ZN(n8638) );
  INV_X1 U10298 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n8636) );
  OR2_X1 U10299 ( .A1(n8851), .A2(n8636), .ZN(n8637) );
  NAND4_X1 U10300 ( .A1(n8640), .A2(n8639), .A3(n8638), .A4(n8637), .ZN(n14362) );
  NOR2_X1 U10301 ( .A1(n14041), .A2(n14362), .ZN(n8642) );
  NAND2_X1 U10302 ( .A1(n14041), .A2(n14362), .ZN(n8641) );
  NAND2_X1 U10303 ( .A1(n10447), .A2(n8612), .ZN(n8650) );
  NAND2_X1 U10304 ( .A1(n8665), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8648) );
  XNOR2_X1 U10305 ( .A(n8648), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10504) );
  AOI22_X1 U10306 ( .A1(n8902), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8901), .B2(
        n10504), .ZN(n8649) );
  NAND2_X1 U10307 ( .A1(n9153), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8659) );
  INV_X1 U10308 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n8651) );
  OR2_X1 U10309 ( .A1(n14219), .A2(n8651), .ZN(n8658) );
  INV_X1 U10310 ( .A(n8654), .ZN(n8652) );
  INV_X1 U10311 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U10312 ( .A1(n8654), .A2(n8653), .ZN(n8655) );
  NAND2_X1 U10313 ( .A1(n8692), .A2(n8655), .ZN(n11338) );
  OR2_X1 U10314 ( .A1(n9039), .A2(n11338), .ZN(n8657) );
  INV_X1 U10315 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10505) );
  OR2_X1 U10316 ( .A1(n8851), .A2(n10505), .ZN(n8656) );
  OR2_X1 U10317 ( .A1(n14047), .A2(n14361), .ZN(n8660) );
  XNOR2_X1 U10318 ( .A(n8679), .B(n8677), .ZN(n10455) );
  NAND2_X1 U10319 ( .A1(n10455), .A2(n8612), .ZN(n8670) );
  INV_X1 U10320 ( .A(n8665), .ZN(n8667) );
  INV_X1 U10321 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8666) );
  NAND2_X1 U10322 ( .A1(n8667), .A2(n8666), .ZN(n8683) );
  NAND2_X1 U10323 ( .A1(n8683), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8668) );
  XNOR2_X1 U10324 ( .A(n8668), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U10325 ( .A1(n8902), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8901), .B2(
        n10507), .ZN(n8669) );
  NAND2_X1 U10326 ( .A1(n8670), .A2(n8669), .ZN(n14055) );
  NAND2_X1 U10327 ( .A1(n8599), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8674) );
  INV_X1 U10328 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10483) );
  OR2_X1 U10329 ( .A1(n8831), .A2(n10483), .ZN(n8673) );
  INV_X1 U10330 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8690) );
  XNOR2_X1 U10331 ( .A(n8692), .B(n8690), .ZN(n11416) );
  OR2_X1 U10332 ( .A1(n9039), .A2(n11416), .ZN(n8672) );
  INV_X1 U10333 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10506) );
  OR2_X1 U10334 ( .A1(n8851), .A2(n10506), .ZN(n8671) );
  NAND4_X1 U10335 ( .A1(n8674), .A2(n8673), .A3(n8672), .A4(n8671), .ZN(n14360) );
  NAND2_X1 U10336 ( .A1(n14055), .A2(n14360), .ZN(n8676) );
  OR2_X1 U10337 ( .A1(n14055), .A2(n14360), .ZN(n8675) );
  NAND2_X1 U10338 ( .A1(n8680), .A2(SI_7_), .ZN(n8681) );
  XNOR2_X1 U10339 ( .A(n8703), .B(n8701), .ZN(n10459) );
  NAND2_X1 U10340 ( .A1(n10459), .A2(n8612), .ZN(n8688) );
  INV_X1 U10341 ( .A(n8683), .ZN(n8685) );
  INV_X1 U10342 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8684) );
  NAND2_X1 U10343 ( .A1(n8685), .A2(n8684), .ZN(n8705) );
  NAND2_X1 U10344 ( .A1(n8705), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8686) );
  XNOR2_X1 U10345 ( .A(n8686), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U10346 ( .A1(n8902), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8901), .B2(
        n10508), .ZN(n8687) );
  NAND2_X1 U10347 ( .A1(n8688), .A2(n8687), .ZN(n14061) );
  NAND2_X1 U10348 ( .A1(n8599), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8698) );
  INV_X1 U10349 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11386) );
  OR2_X1 U10350 ( .A1(n8831), .A2(n11386), .ZN(n8697) );
  INV_X1 U10351 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8689) );
  OAI21_X1 U10352 ( .B1(n8692), .B2(n8690), .A(n8689), .ZN(n8693) );
  NAND2_X1 U10353 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .ZN(n8691) );
  NAND2_X1 U10354 ( .A1(n8693), .A2(n8710), .ZN(n11385) );
  OR2_X1 U10355 ( .A1(n9039), .A2(n11385), .ZN(n8696) );
  INV_X1 U10356 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8694) );
  OR2_X1 U10357 ( .A1(n8851), .A2(n8694), .ZN(n8695) );
  NAND4_X1 U10358 ( .A1(n8698), .A2(n8697), .A3(n8696), .A4(n8695), .ZN(n14359) );
  INV_X1 U10359 ( .A(n14359), .ZN(n11234) );
  XNOR2_X1 U10360 ( .A(n14061), .B(n11234), .ZN(n14294) );
  NAND2_X1 U10361 ( .A1(n11389), .A2(n14294), .ZN(n8700) );
  NAND2_X1 U10362 ( .A1(n14061), .A2(n14359), .ZN(n8699) );
  NAND2_X1 U10363 ( .A1(n8700), .A2(n8699), .ZN(n11604) );
  NAND2_X1 U10364 ( .A1(n10472), .A2(n8612), .ZN(n8708) );
  NAND2_X1 U10365 ( .A1(n8706), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8725) );
  XNOR2_X1 U10366 ( .A(n8725), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10676) );
  AOI22_X1 U10367 ( .A1(n8902), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8901), .B2(
        n10676), .ZN(n8707) );
  NAND2_X1 U10368 ( .A1(n8599), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8716) );
  INV_X1 U10369 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n14626) );
  OR2_X1 U10370 ( .A1(n8831), .A2(n14626), .ZN(n8715) );
  INV_X1 U10371 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U10372 ( .A1(n8710), .A2(n8709), .ZN(n8711) );
  NAND2_X1 U10373 ( .A1(n8731), .A2(n8711), .ZN(n14625) );
  OR2_X1 U10374 ( .A1(n9039), .A2(n14625), .ZN(n8714) );
  INV_X1 U10375 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8712) );
  OR2_X1 U10376 ( .A1(n8851), .A2(n8712), .ZN(n8713) );
  NAND4_X1 U10377 ( .A1(n8716), .A2(n8715), .A3(n8714), .A4(n8713), .ZN(n14358) );
  XNOR2_X1 U10378 ( .A(n14629), .B(n14358), .ZN(n14297) );
  INV_X1 U10379 ( .A(n14297), .ZN(n8717) );
  NAND2_X1 U10380 ( .A1(n14629), .A2(n14358), .ZN(n8718) );
  INV_X1 U10381 ( .A(n8719), .ZN(n8722) );
  NAND2_X1 U10382 ( .A1(n8720), .A2(SI_9_), .ZN(n8721) );
  XNOR2_X1 U10383 ( .A(n8742), .B(n8740), .ZN(n10477) );
  NAND2_X1 U10384 ( .A1(n10477), .A2(n8612), .ZN(n8728) );
  INV_X1 U10385 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8724) );
  NAND2_X1 U10386 ( .A1(n8725), .A2(n8724), .ZN(n8726) );
  NAND2_X1 U10387 ( .A1(n8726), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8753) );
  XNOR2_X1 U10388 ( .A(n8753), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10706) );
  AOI22_X1 U10389 ( .A1(n10706), .A2(n8901), .B1(n8902), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n8727) );
  NAND2_X1 U10390 ( .A1(n8599), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8737) );
  INV_X1 U10391 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11638) );
  OR2_X1 U10392 ( .A1(n8831), .A2(n11638), .ZN(n8736) );
  INV_X1 U10393 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8730) );
  NAND2_X1 U10394 ( .A1(n8731), .A2(n8730), .ZN(n8732) );
  NAND2_X1 U10395 ( .A1(n8759), .A2(n8732), .ZN(n11637) );
  OR2_X1 U10396 ( .A1(n9039), .A2(n11637), .ZN(n8735) );
  INV_X1 U10397 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8733) );
  OR2_X1 U10398 ( .A1(n8851), .A2(n8733), .ZN(n8734) );
  NAND4_X1 U10399 ( .A1(n8737), .A2(n8736), .A3(n8735), .A4(n8734), .ZN(n14357) );
  OR2_X1 U10400 ( .A1(n14073), .A2(n14357), .ZN(n8738) );
  NAND2_X1 U10401 ( .A1(n14073), .A2(n14357), .ZN(n8739) );
  NAND2_X1 U10402 ( .A1(n8742), .A2(n8741), .ZN(n8745) );
  NAND2_X1 U10403 ( .A1(n8743), .A2(SI_10_), .ZN(n8744) );
  INV_X1 U10404 ( .A(SI_11_), .ZN(n13437) );
  INV_X1 U10405 ( .A(n8746), .ZN(n8747) );
  NAND2_X1 U10406 ( .A1(n8747), .A2(SI_11_), .ZN(n8748) );
  NAND2_X1 U10407 ( .A1(n8750), .A2(n8749), .ZN(n8751) );
  NAND2_X1 U10408 ( .A1(n8767), .A2(n8751), .ZN(n10541) );
  NAND2_X1 U10409 ( .A1(n10541), .A2(n8612), .ZN(n8757) );
  INV_X1 U10410 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U10411 ( .A1(n8753), .A2(n8752), .ZN(n8754) );
  NAND2_X1 U10412 ( .A1(n8754), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8755) );
  XNOR2_X1 U10413 ( .A(n8755), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10837) );
  AOI22_X1 U10414 ( .A1(n10837), .A2(n8901), .B1(n8902), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8756) );
  NAND2_X2 U10415 ( .A1(n8757), .A2(n8756), .ZN(n14086) );
  NAND2_X1 U10416 ( .A1(n9153), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8765) );
  INV_X1 U10417 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10715) );
  OR2_X1 U10418 ( .A1(n8851), .A2(n10715), .ZN(n8764) );
  INV_X1 U10419 ( .A(n8759), .ZN(n8758) );
  NAND2_X1 U10420 ( .A1(n8758), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8778) );
  INV_X1 U10421 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10710) );
  NAND2_X1 U10422 ( .A1(n8759), .A2(n10710), .ZN(n8760) );
  NAND2_X1 U10423 ( .A1(n8778), .A2(n8760), .ZN(n11875) );
  OR2_X1 U10424 ( .A1(n9039), .A2(n11875), .ZN(n8763) );
  INV_X1 U10425 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8761) );
  OR2_X1 U10426 ( .A1(n14219), .A2(n8761), .ZN(n8762) );
  NAND4_X1 U10427 ( .A1(n8765), .A2(n8764), .A3(n8763), .A4(n8762), .ZN(n14356) );
  XNOR2_X1 U10428 ( .A(n14086), .B(n14356), .ZN(n14299) );
  INV_X1 U10429 ( .A(n14299), .ZN(n11646) );
  INV_X1 U10430 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10701) );
  INV_X1 U10431 ( .A(n8768), .ZN(n8769) );
  NAND2_X1 U10432 ( .A1(n8769), .A2(SI_12_), .ZN(n8770) );
  XNOR2_X1 U10433 ( .A(n8784), .B(n8514), .ZN(n10654) );
  NAND2_X1 U10434 ( .A1(n10654), .A2(n8612), .ZN(n8775) );
  NAND2_X1 U10435 ( .A1(n8771), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8772) );
  MUX2_X1 U10436 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8772), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8773) );
  OR2_X1 U10437 ( .A1(n8771), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8805) );
  AND2_X1 U10438 ( .A1(n8773), .A2(n8805), .ZN(n11072) );
  AOI22_X1 U10439 ( .A1(n8902), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8901), 
        .B2(n11072), .ZN(n8774) );
  NAND2_X1 U10440 ( .A1(n8599), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8783) );
  INV_X1 U10441 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8776) );
  OR2_X1 U10442 ( .A1(n8831), .A2(n8776), .ZN(n8782) );
  INV_X1 U10443 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U10444 ( .A1(n8778), .A2(n8777), .ZN(n8779) );
  NAND2_X1 U10445 ( .A1(n8792), .A2(n8779), .ZN(n11904) );
  OR2_X1 U10446 ( .A1(n9039), .A2(n11904), .ZN(n8781) );
  INV_X1 U10447 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10836) );
  OR2_X1 U10448 ( .A1(n8851), .A2(n10836), .ZN(n8780) );
  NAND4_X1 U10449 ( .A1(n8783), .A2(n8782), .A3(n8781), .A4(n8780), .ZN(n14355) );
  INV_X1 U10450 ( .A(n14355), .ZN(n14096) );
  XNOR2_X1 U10451 ( .A(n14094), .B(n14096), .ZN(n14301) );
  NAND2_X1 U10452 ( .A1(n10782), .A2(n8612), .ZN(n8789) );
  NAND2_X1 U10453 ( .A1(n8805), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8787) );
  XNOR2_X1 U10454 ( .A(n8787), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U10455 ( .A1(n8902), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8901), 
        .B2(n11554), .ZN(n8788) );
  NAND2_X1 U10456 ( .A1(n8599), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8798) );
  INV_X1 U10457 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n12092) );
  OR2_X1 U10458 ( .A1(n8831), .A2(n12092), .ZN(n8797) );
  INV_X1 U10459 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8791) );
  NAND2_X1 U10460 ( .A1(n8792), .A2(n8791), .ZN(n8793) );
  NAND2_X1 U10461 ( .A1(n8812), .A2(n8793), .ZN(n12091) );
  OR2_X1 U10462 ( .A1(n9039), .A2(n12091), .ZN(n8796) );
  INV_X1 U10463 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8794) );
  OR2_X1 U10464 ( .A1(n14218), .A2(n8794), .ZN(n8795) );
  NAND4_X1 U10465 ( .A1(n8798), .A2(n8797), .A3(n8796), .A4(n8795), .ZN(n14354) );
  INV_X1 U10466 ( .A(n14354), .ZN(n11891) );
  XNOR2_X1 U10467 ( .A(n7765), .B(n11891), .ZN(n14302) );
  INV_X1 U10468 ( .A(n14302), .ZN(n12084) );
  NAND2_X1 U10469 ( .A1(n12083), .A2(n14302), .ZN(n12082) );
  OR2_X1 U10470 ( .A1(n7765), .A2(n14354), .ZN(n8799) );
  NAND2_X1 U10471 ( .A1(n8801), .A2(SI_13_), .ZN(n8802) );
  XNOR2_X1 U10472 ( .A(n8819), .B(n8839), .ZN(n11062) );
  NAND2_X1 U10473 ( .A1(n11062), .A2(n8612), .ZN(n8809) );
  NOR2_X1 U10474 ( .A1(n8805), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8824) );
  INV_X1 U10475 ( .A(n8824), .ZN(n8806) );
  NAND2_X1 U10476 ( .A1(n8806), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8807) );
  XNOR2_X1 U10477 ( .A(n8807), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U10478 ( .A1(n8902), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8901), 
        .B2(n11555), .ZN(n8808) );
  NAND2_X1 U10479 ( .A1(n9153), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8817) );
  INV_X1 U10480 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8810) );
  OR2_X1 U10481 ( .A1(n14219), .A2(n8810), .ZN(n8816) );
  INV_X1 U10482 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8811) );
  NAND2_X1 U10483 ( .A1(n8812), .A2(n8811), .ZN(n8813) );
  NAND2_X1 U10484 ( .A1(n8829), .A2(n8813), .ZN(n12279) );
  OR2_X1 U10485 ( .A1(n9039), .A2(n12279), .ZN(n8815) );
  INV_X1 U10486 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11805) );
  OR2_X1 U10487 ( .A1(n8851), .A2(n11805), .ZN(n8814) );
  NAND4_X1 U10488 ( .A1(n8817), .A2(n8816), .A3(n8815), .A4(n8814), .ZN(n14353) );
  INV_X1 U10489 ( .A(n14353), .ZN(n14107) );
  XNOR2_X1 U10490 ( .A(n14725), .B(n14107), .ZN(n14303) );
  NAND2_X1 U10491 ( .A1(n14725), .A2(n14353), .ZN(n8818) );
  INV_X1 U10492 ( .A(n8821), .ZN(n8822) );
  INV_X1 U10493 ( .A(SI_15_), .ZN(n13428) );
  NAND2_X1 U10494 ( .A1(n8822), .A2(n13428), .ZN(n8840) );
  NAND2_X1 U10495 ( .A1(n11263), .A2(n8612), .ZN(n8827) );
  NAND2_X1 U10496 ( .A1(n8824), .A2(n8823), .ZN(n8846) );
  NAND2_X1 U10497 ( .A1(n8846), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8825) );
  XNOR2_X1 U10498 ( .A(n8825), .B(P2_IR_REG_15__SCAN_IN), .ZN(n12349) );
  AOI22_X1 U10499 ( .A1(n8902), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8901), 
        .B2(n12349), .ZN(n8826) );
  NAND2_X1 U10500 ( .A1(n8599), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8836) );
  INV_X1 U10501 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8828) );
  NAND2_X1 U10502 ( .A1(n8829), .A2(n8828), .ZN(n8830) );
  NAND2_X1 U10503 ( .A1(n8870), .A2(n8830), .ZN(n12385) );
  OR2_X1 U10504 ( .A1(n9039), .A2(n12385), .ZN(n8835) );
  INV_X1 U10505 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n12379) );
  OR2_X1 U10506 ( .A1(n8831), .A2(n12379), .ZN(n8834) );
  INV_X1 U10507 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8832) );
  OR2_X1 U10508 ( .A1(n8851), .A2(n8832), .ZN(n8833) );
  NAND4_X1 U10509 ( .A1(n8836), .A2(n8835), .A3(n8834), .A4(n8833), .ZN(n14352) );
  XNOR2_X1 U10510 ( .A(n7757), .B(n14352), .ZN(n14305) );
  OR2_X1 U10511 ( .A1(n7757), .A2(n14352), .ZN(n8837) );
  INV_X1 U10512 ( .A(SI_14_), .ZN(n10465) );
  NOR2_X1 U10513 ( .A1(n8839), .A2(SI_14_), .ZN(n8843) );
  INV_X1 U10514 ( .A(n8840), .ZN(n8841) );
  XNOR2_X1 U10515 ( .A(n8878), .B(SI_16_), .ZN(n8858) );
  INV_X1 U10516 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11476) );
  XNOR2_X1 U10517 ( .A(n8858), .B(n8876), .ZN(n11473) );
  NAND2_X1 U10518 ( .A1(n11473), .A2(n8612), .ZN(n8850) );
  OAI21_X1 U10519 ( .B1(n8846), .B2(P2_IR_REG_15__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8847) );
  MUX2_X1 U10520 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8847), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n8848) );
  AND2_X1 U10521 ( .A1(n8848), .A2(n7611), .ZN(n15859) );
  AOI22_X1 U10522 ( .A1(n8902), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8901), 
        .B2(n15859), .ZN(n8849) );
  INV_X1 U10523 ( .A(n9039), .ZN(n9058) );
  XNOR2_X1 U10524 ( .A(n8870), .B(P2_REG3_REG_16__SCAN_IN), .ZN(n12317) );
  NAND2_X1 U10525 ( .A1(n9058), .A2(n12317), .ZN(n8855) );
  INV_X1 U10526 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n14766) );
  OR2_X1 U10527 ( .A1(n14219), .A2(n14766), .ZN(n8854) );
  INV_X1 U10528 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12437) );
  OR2_X1 U10529 ( .A1(n8831), .A2(n12437), .ZN(n8853) );
  INV_X1 U10530 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n14713) );
  OR2_X1 U10531 ( .A1(n8851), .A2(n14713), .ZN(n8852) );
  NAND4_X1 U10532 ( .A1(n8855), .A2(n8854), .A3(n8853), .A4(n8852), .ZN(n14351) );
  XNOR2_X1 U10533 ( .A(n14122), .B(n14351), .ZN(n14304) );
  NAND2_X1 U10534 ( .A1(n14122), .A2(n14351), .ZN(n8857) );
  INV_X1 U10535 ( .A(n8876), .ZN(n8879) );
  NAND2_X1 U10536 ( .A1(n8858), .A2(n8879), .ZN(n8860) );
  INV_X1 U10537 ( .A(SI_16_), .ZN(n10517) );
  OR2_X1 U10538 ( .A1(n8878), .A2(n10517), .ZN(n8859) );
  NAND2_X1 U10539 ( .A1(n8860), .A2(n8859), .ZN(n8864) );
  NAND2_X1 U10540 ( .A1(n8861), .A2(SI_17_), .ZN(n8882) );
  INV_X1 U10541 ( .A(n8861), .ZN(n8862) );
  INV_X1 U10542 ( .A(SI_17_), .ZN(n10548) );
  NAND2_X1 U10543 ( .A1(n8862), .A2(n10548), .ZN(n8880) );
  NAND2_X1 U10544 ( .A1(n8882), .A2(n8880), .ZN(n8863) );
  NAND2_X1 U10545 ( .A1(n11546), .A2(n8612), .ZN(n8867) );
  NAND2_X1 U10546 ( .A1(n7611), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8865) );
  XNOR2_X1 U10547 ( .A(n8865), .B(P2_IR_REG_17__SCAN_IN), .ZN(n12354) );
  AOI22_X1 U10548 ( .A1(n8902), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8901), 
        .B2(n12354), .ZN(n8866) );
  AND2_X1 U10549 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n8868) );
  INV_X1 U10550 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n12318) );
  INV_X1 U10551 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n12421) );
  OAI21_X1 U10552 ( .B1(n8870), .B2(n12318), .A(n12421), .ZN(n8871) );
  NAND2_X1 U10553 ( .A1(n8889), .A2(n8871), .ZN(n12517) );
  OR2_X1 U10554 ( .A1(n12517), .A2(n9039), .ZN(n8875) );
  NAND2_X1 U10555 ( .A1(n8599), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8874) );
  INV_X1 U10556 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n12518) );
  OR2_X1 U10557 ( .A1(n8831), .A2(n12518), .ZN(n8873) );
  NAND2_X1 U10558 ( .A1(n9154), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8872) );
  NAND4_X1 U10559 ( .A1(n8875), .A2(n8874), .A3(n8873), .A4(n8872), .ZN(n14350) );
  INV_X1 U10560 ( .A(n14350), .ZN(n14133) );
  INV_X1 U10561 ( .A(n14307), .ZN(n12513) );
  OAI21_X1 U10562 ( .B1(n8876), .B2(n10517), .A(n8882), .ZN(n8877) );
  NOR2_X1 U10563 ( .A1(n8879), .A2(SI_16_), .ZN(n8883) );
  INV_X1 U10564 ( .A(n8880), .ZN(n8881) );
  AOI21_X1 U10565 ( .B1(n8883), .B2(n8882), .A(n8881), .ZN(n8884) );
  XNOR2_X1 U10566 ( .A(n8914), .B(SI_18_), .ZN(n8894) );
  INV_X1 U10567 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11588) );
  INV_X1 U10568 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11586) );
  XNOR2_X1 U10569 ( .A(n8894), .B(n8911), .ZN(n11585) );
  NAND2_X1 U10570 ( .A1(n11585), .A2(n8612), .ZN(n8888) );
  XNOR2_X1 U10571 ( .A(n8886), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14413) );
  AOI22_X1 U10572 ( .A1(n8902), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8901), 
        .B2(n14413), .ZN(n8887) );
  INV_X1 U10573 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n13969) );
  NAND2_X1 U10574 ( .A1(n8889), .A2(n13969), .ZN(n8890) );
  NAND2_X1 U10575 ( .A1(n8926), .A2(n8890), .ZN(n14614) );
  AOI22_X1 U10576 ( .A1(n8599), .A2(P2_REG0_REG_18__SCAN_IN), .B1(n9153), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U10577 ( .A1(n9154), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8891) );
  OAI211_X1 U10578 ( .C1(n14614), .C2(n9039), .A(n8892), .B(n8891), .ZN(n14587) );
  INV_X1 U10579 ( .A(n14587), .ZN(n13901) );
  XNOR2_X1 U10580 ( .A(n14698), .B(n13901), .ZN(n14609) );
  OR2_X1 U10581 ( .A1(n14698), .A2(n14587), .ZN(n8893) );
  INV_X1 U10582 ( .A(n8911), .ZN(n8915) );
  NAND2_X1 U10583 ( .A1(n8894), .A2(n8915), .ZN(n8896) );
  INV_X1 U10584 ( .A(SI_18_), .ZN(n10703) );
  OR2_X1 U10585 ( .A1(n8914), .A2(n10703), .ZN(n8895) );
  NAND2_X1 U10586 ( .A1(n8896), .A2(n8895), .ZN(n8900) );
  NAND2_X1 U10587 ( .A1(n8897), .A2(SI_19_), .ZN(n8918) );
  INV_X1 U10588 ( .A(n8897), .ZN(n8898) );
  INV_X1 U10589 ( .A(SI_19_), .ZN(n10877) );
  NAND2_X1 U10590 ( .A1(n8898), .A2(n10877), .ZN(n8916) );
  NAND2_X1 U10591 ( .A1(n8918), .A2(n8916), .ZN(n8899) );
  NAND2_X1 U10592 ( .A1(n11600), .A2(n8612), .ZN(n8904) );
  AOI22_X1 U10593 ( .A1(n8902), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7431), 
        .B2(n8901), .ZN(n8903) );
  XNOR2_X1 U10594 ( .A(n8926), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n14597) );
  NAND2_X1 U10595 ( .A1(n14597), .A2(n9058), .ZN(n8909) );
  NAND2_X1 U10596 ( .A1(n8599), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8906) );
  NAND2_X1 U10597 ( .A1(n9154), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8905) );
  OAI211_X1 U10598 ( .C1(n8831), .C2(n14419), .A(n8906), .B(n8905), .ZN(n8907)
         );
  INV_X1 U10599 ( .A(n8907), .ZN(n8908) );
  NAND2_X1 U10600 ( .A1(n8909), .A2(n8908), .ZN(n14349) );
  INV_X1 U10601 ( .A(n14349), .ZN(n14152) );
  XNOR2_X1 U10602 ( .A(n14596), .B(n14152), .ZN(n14586) );
  NAND2_X1 U10603 ( .A1(n14582), .A2(n14586), .ZN(n14581) );
  OR2_X1 U10604 ( .A1(n14596), .A2(n14349), .ZN(n8910) );
  OAI21_X1 U10605 ( .B1(n8911), .B2(n10703), .A(n8918), .ZN(n8912) );
  INV_X1 U10606 ( .A(n8912), .ZN(n8913) );
  NOR2_X1 U10607 ( .A1(n8915), .A2(SI_18_), .ZN(n8919) );
  INV_X1 U10608 ( .A(n8916), .ZN(n8917) );
  AOI21_X1 U10609 ( .B1(n8919), .B2(n8918), .A(n8917), .ZN(n8920) );
  INV_X1 U10610 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11617) );
  INV_X1 U10611 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11707) );
  XNOR2_X1 U10612 ( .A(n8937), .B(n8935), .ZN(n11616) );
  NAND2_X1 U10613 ( .A1(n11616), .A2(n8612), .ZN(n8923) );
  OR2_X1 U10614 ( .A1(n14253), .A2(n11707), .ZN(n8922) );
  INV_X1 U10615 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8932) );
  INV_X1 U10616 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8925) );
  INV_X1 U10617 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8924) );
  OAI21_X1 U10618 ( .B1(n8926), .B2(n8925), .A(n8924), .ZN(n8929) );
  AND2_X1 U10619 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n8927) );
  NAND2_X1 U10620 ( .A1(n8929), .A2(n8943), .ZN(n13956) );
  OR2_X1 U10621 ( .A1(n13956), .A2(n9039), .ZN(n8931) );
  AOI22_X1 U10622 ( .A1(n8599), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n9153), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n8930) );
  OAI211_X1 U10623 ( .C1(n8851), .C2(n8932), .A(n8931), .B(n8930), .ZN(n14590)
         );
  INV_X1 U10624 ( .A(n14590), .ZN(n13958) );
  NAND2_X1 U10625 ( .A1(n14688), .A2(n13958), .ZN(n8933) );
  OR2_X1 U10626 ( .A1(n14688), .A2(n14590), .ZN(n8934) );
  INV_X1 U10627 ( .A(n8935), .ZN(n8936) );
  XNOR2_X1 U10628 ( .A(n8954), .B(SI_21_), .ZN(n8951) );
  XNOR2_X1 U10629 ( .A(n8953), .B(n8951), .ZN(n11677) );
  NAND2_X1 U10630 ( .A1(n11677), .A2(n8612), .ZN(n8942) );
  INV_X1 U10631 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11680) );
  OR2_X1 U10632 ( .A1(n14253), .A2(n11680), .ZN(n8941) );
  INV_X1 U10633 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13926) );
  NAND2_X1 U10634 ( .A1(n8943), .A2(n13926), .ZN(n8944) );
  NAND2_X1 U10635 ( .A1(n8958), .A2(n8944), .ZN(n14552) );
  OR2_X1 U10636 ( .A1(n14552), .A2(n9039), .ZN(n8950) );
  INV_X1 U10637 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8947) );
  NAND2_X1 U10638 ( .A1(n9153), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8946) );
  NAND2_X1 U10639 ( .A1(n9154), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8945) );
  OAI211_X1 U10640 ( .C1(n14219), .C2(n8947), .A(n8946), .B(n8945), .ZN(n8948)
         );
  INV_X1 U10641 ( .A(n8948), .ZN(n8949) );
  INV_X1 U10642 ( .A(n14165), .ZN(n14348) );
  XNOR2_X1 U10643 ( .A(n14681), .B(n14348), .ZN(n14558) );
  INV_X1 U10644 ( .A(n8951), .ZN(n8952) );
  NAND2_X1 U10645 ( .A1(n8954), .A2(SI_21_), .ZN(n8955) );
  XNOR2_X1 U10646 ( .A(n9235), .B(n8987), .ZN(n11983) );
  NAND2_X1 U10647 ( .A1(n11983), .A2(n8612), .ZN(n8957) );
  INV_X1 U10648 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11985) );
  OR2_X1 U10649 ( .A1(n14253), .A2(n11985), .ZN(n8956) );
  INV_X1 U10650 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n12550) );
  NAND2_X1 U10651 ( .A1(n8958), .A2(n12550), .ZN(n8959) );
  NAND2_X1 U10652 ( .A1(n8974), .A2(n8959), .ZN(n14540) );
  INV_X1 U10653 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U10654 ( .A1(n9153), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8961) );
  NAND2_X1 U10655 ( .A1(n9154), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8960) );
  OAI211_X1 U10656 ( .C1(n14219), .C2(n8962), .A(n8961), .B(n8960), .ZN(n8963)
         );
  INV_X1 U10657 ( .A(n8963), .ZN(n8964) );
  OAI21_X1 U10658 ( .B1(n14540), .B2(n9039), .A(n8964), .ZN(n14347) );
  XNOR2_X1 U10659 ( .A(n14675), .B(n14347), .ZN(n14541) );
  NAND2_X1 U10660 ( .A1(n14675), .A2(n14347), .ZN(n8966) );
  INV_X1 U10661 ( .A(n9235), .ZN(n8968) );
  AND2_X1 U10662 ( .A1(n8986), .A2(SI_22_), .ZN(n8967) );
  INV_X1 U10663 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10151) );
  INV_X1 U10664 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n12152) );
  XNOR2_X1 U10665 ( .A(n8989), .B(SI_23_), .ZN(n8969) );
  NAND2_X1 U10666 ( .A1(n12149), .A2(n8612), .ZN(n8972) );
  OR2_X1 U10667 ( .A1(n14253), .A2(n12152), .ZN(n8971) );
  INV_X1 U10668 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8973) );
  NAND2_X1 U10669 ( .A1(n8974), .A2(n8973), .ZN(n8975) );
  AND2_X1 U10670 ( .A1(n8999), .A2(n8975), .ZN(n14526) );
  NAND2_X1 U10671 ( .A1(n14526), .A2(n9058), .ZN(n8981) );
  INV_X1 U10672 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U10673 ( .A1(n9154), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8977) );
  NAND2_X1 U10674 ( .A1(n9153), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8976) );
  OAI211_X1 U10675 ( .C1(n14219), .C2(n8978), .A(n8977), .B(n8976), .ZN(n8979)
         );
  INV_X1 U10676 ( .A(n8979), .ZN(n8980) );
  OR2_X1 U10677 ( .A1(n14529), .A2(n14177), .ZN(n8982) );
  INV_X1 U10678 ( .A(SI_23_), .ZN(n13614) );
  NAND2_X1 U10679 ( .A1(n8989), .A2(n13614), .ZN(n8991) );
  OAI21_X1 U10680 ( .B1(SI_22_), .B2(n8987), .A(n8991), .ZN(n8984) );
  INV_X1 U10681 ( .A(n8984), .ZN(n8985) );
  INV_X1 U10682 ( .A(n8987), .ZN(n8988) );
  INV_X1 U10683 ( .A(SI_22_), .ZN(n10139) );
  NOR2_X1 U10684 ( .A1(n8988), .A2(n10139), .ZN(n8992) );
  INV_X1 U10685 ( .A(n8989), .ZN(n8990) );
  AOI22_X1 U10686 ( .A1(n8992), .A2(n8991), .B1(n8990), .B2(SI_23_), .ZN(n8993) );
  INV_X1 U10687 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10180) );
  INV_X1 U10688 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12191) );
  INV_X1 U10689 ( .A(n9007), .ZN(n8994) );
  NAND2_X1 U10690 ( .A1(n12104), .A2(n8612), .ZN(n8996) );
  OR2_X1 U10691 ( .A1(n14253), .A2(n12191), .ZN(n8995) );
  INV_X1 U10692 ( .A(n8999), .ZN(n8997) );
  INV_X1 U10693 ( .A(n9021), .ZN(n9023) );
  INV_X1 U10694 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8998) );
  NAND2_X1 U10695 ( .A1(n8999), .A2(n8998), .ZN(n9000) );
  NAND2_X1 U10696 ( .A1(n9023), .A2(n9000), .ZN(n14512) );
  OR2_X1 U10697 ( .A1(n14512), .A2(n9039), .ZN(n9005) );
  INV_X1 U10698 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n14750) );
  NAND2_X1 U10699 ( .A1(n9154), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9002) );
  NAND2_X1 U10700 ( .A1(n9153), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9001) );
  OAI211_X1 U10701 ( .C1(n14219), .C2(n14750), .A(n9002), .B(n9001), .ZN(n9003) );
  INV_X1 U10702 ( .A(n9003), .ZN(n9004) );
  NAND2_X1 U10703 ( .A1(n9005), .A2(n9004), .ZN(n14345) );
  INV_X1 U10704 ( .A(n14345), .ZN(n13933) );
  XNOR2_X1 U10705 ( .A(n14511), .B(n13933), .ZN(n14505) );
  INV_X1 U10706 ( .A(n14505), .ZN(n9140) );
  OR2_X1 U10707 ( .A1(n14511), .A2(n14345), .ZN(n9006) );
  INV_X1 U10708 ( .A(n9008), .ZN(n9009) );
  NAND2_X1 U10709 ( .A1(n9010), .A2(n9009), .ZN(n9011) );
  INV_X1 U10710 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12534) );
  INV_X1 U10711 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12223) );
  INV_X1 U10712 ( .A(SI_25_), .ZN(n13610) );
  NAND2_X1 U10713 ( .A1(n9013), .A2(n13610), .ZN(n9031) );
  INV_X1 U10714 ( .A(n9013), .ZN(n9014) );
  NAND2_X1 U10715 ( .A1(n9014), .A2(SI_25_), .ZN(n9015) );
  NAND2_X1 U10716 ( .A1(n9031), .A2(n9015), .ZN(n9016) );
  NAND2_X1 U10717 ( .A1(n9017), .A2(n9016), .ZN(n9018) );
  NAND2_X1 U10718 ( .A1(n9032), .A2(n9018), .ZN(n12221) );
  NAND2_X1 U10719 ( .A1(n12221), .A2(n8612), .ZN(n9020) );
  OR2_X1 U10720 ( .A1(n14253), .A2(n12223), .ZN(n9019) );
  INV_X1 U10721 ( .A(n9035), .ZN(n9037) );
  INV_X1 U10722 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9022) );
  NAND2_X1 U10723 ( .A1(n9023), .A2(n9022), .ZN(n9024) );
  NAND2_X1 U10724 ( .A1(n14498), .A2(n9058), .ZN(n9029) );
  INV_X1 U10725 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14746) );
  NAND2_X1 U10726 ( .A1(n9154), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n9026) );
  NAND2_X1 U10727 ( .A1(n9153), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9025) );
  OAI211_X1 U10728 ( .C1(n14219), .C2(n14746), .A(n9026), .B(n9025), .ZN(n9027) );
  INV_X1 U10729 ( .A(n9027), .ZN(n9028) );
  NAND2_X1 U10730 ( .A1(n9029), .A2(n9028), .ZN(n14344) );
  XNOR2_X1 U10731 ( .A(n14497), .B(n14344), .ZN(n14310) );
  INV_X1 U10732 ( .A(n14310), .ZN(n14491) );
  OR2_X1 U10733 ( .A1(n14497), .A2(n14344), .ZN(n9030) );
  INV_X1 U10734 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15778) );
  INV_X1 U10735 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14788) );
  XNOR2_X1 U10736 ( .A(n9047), .B(SI_26_), .ZN(n9046) );
  NAND2_X1 U10737 ( .A1(n14786), .A2(n8612), .ZN(n9034) );
  OR2_X1 U10738 ( .A1(n14253), .A2(n14788), .ZN(n9033) );
  NAND2_X2 U10739 ( .A1(n9034), .A2(n9033), .ZN(n14482) );
  NAND2_X1 U10740 ( .A1(n9035), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n9056) );
  INV_X1 U10741 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9036) );
  NAND2_X1 U10742 ( .A1(n9037), .A2(n9036), .ZN(n9038) );
  NAND2_X1 U10743 ( .A1(n9056), .A2(n9038), .ZN(n13984) );
  OR2_X1 U10744 ( .A1(n13984), .A2(n9039), .ZN(n9044) );
  INV_X1 U10745 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n14742) );
  NAND2_X1 U10746 ( .A1(n9153), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9041) );
  NAND2_X1 U10747 ( .A1(n9154), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n9040) );
  OAI211_X1 U10748 ( .C1(n14742), .C2(n14219), .A(n9041), .B(n9040), .ZN(n9042) );
  INV_X1 U10749 ( .A(n9042), .ZN(n9043) );
  NAND2_X1 U10750 ( .A1(n9044), .A2(n9043), .ZN(n14343) );
  XNOR2_X1 U10751 ( .A(n14482), .B(n14343), .ZN(n14313) );
  OR2_X1 U10752 ( .A1(n14482), .A2(n14343), .ZN(n9045) );
  INV_X1 U10753 ( .A(n9046), .ZN(n9050) );
  INV_X1 U10754 ( .A(n9047), .ZN(n9048) );
  NAND2_X1 U10755 ( .A1(n9048), .A2(SI_26_), .ZN(n9049) );
  INV_X1 U10756 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15776) );
  INV_X1 U10757 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14784) );
  XNOR2_X1 U10758 ( .A(n9069), .B(SI_27_), .ZN(n9067) );
  INV_X1 U10759 ( .A(n9067), .ZN(n9052) );
  NAND2_X1 U10760 ( .A1(n14781), .A2(n8612), .ZN(n9054) );
  OR2_X1 U10761 ( .A1(n14253), .A2(n14784), .ZN(n9053) );
  INV_X1 U10762 ( .A(n9056), .ZN(n9055) );
  INV_X1 U10763 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13880) );
  NAND2_X1 U10764 ( .A1(n9056), .A2(n13880), .ZN(n9057) );
  NAND2_X1 U10765 ( .A1(n14467), .A2(n9058), .ZN(n9063) );
  INV_X1 U10766 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n14739) );
  NAND2_X1 U10767 ( .A1(n9154), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9060) );
  NAND2_X1 U10768 ( .A1(n9153), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9059) );
  OAI211_X1 U10769 ( .C1(n14219), .C2(n14739), .A(n9060), .B(n9059), .ZN(n9061) );
  INV_X1 U10770 ( .A(n9061), .ZN(n9062) );
  NAND2_X1 U10771 ( .A1(n14198), .A2(n14342), .ZN(n9066) );
  OR2_X1 U10772 ( .A1(n14198), .A2(n14342), .ZN(n9064) );
  INV_X1 U10773 ( .A(n9069), .ZN(n9070) );
  INV_X1 U10774 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n15774) );
  INV_X1 U10775 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10242) );
  INV_X1 U10776 ( .A(SI_28_), .ZN(n13410) );
  NAND2_X1 U10777 ( .A1(n9071), .A2(n13410), .ZN(n9090) );
  INV_X1 U10778 ( .A(n9071), .ZN(n9072) );
  NAND2_X1 U10779 ( .A1(n9072), .A2(SI_28_), .ZN(n9073) );
  NAND2_X1 U10780 ( .A1(n9090), .A2(n9073), .ZN(n9074) );
  NAND2_X1 U10781 ( .A1(n9075), .A2(n9074), .ZN(n9076) );
  NAND2_X1 U10782 ( .A1(n14778), .A2(n8612), .ZN(n9078) );
  OR2_X1 U10783 ( .A1(n14253), .A2(n10242), .ZN(n9077) );
  NAND2_X1 U10784 ( .A1(n9079), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n14444) );
  INV_X1 U10785 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9080) );
  NAND2_X1 U10786 ( .A1(n9081), .A2(n9080), .ZN(n9082) );
  NAND2_X1 U10787 ( .A1(n14444), .A2(n9082), .ZN(n13912) );
  INV_X1 U10788 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9742) );
  NAND2_X1 U10789 ( .A1(n9153), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U10790 ( .A1(n9154), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9083) );
  OAI211_X1 U10791 ( .C1(n9742), .C2(n14219), .A(n9084), .B(n9083), .ZN(n9085)
         );
  INV_X1 U10792 ( .A(n9085), .ZN(n9086) );
  NAND2_X1 U10793 ( .A1(n9087), .A2(n9086), .ZN(n14341) );
  INV_X1 U10794 ( .A(n14341), .ZN(n9088) );
  NAND2_X1 U10795 ( .A1(n14193), .A2(n9088), .ZN(n9089) );
  INV_X1 U10796 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15771) );
  INV_X1 U10797 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n12792) );
  INV_X1 U10798 ( .A(SI_29_), .ZN(n13851) );
  NAND2_X1 U10799 ( .A1(n9092), .A2(n13851), .ZN(n14223) );
  INV_X1 U10800 ( .A(n9092), .ZN(n9093) );
  NAND2_X1 U10801 ( .A1(n9093), .A2(SI_29_), .ZN(n9094) );
  AND2_X1 U10802 ( .A1(n14223), .A2(n9094), .ZN(n9095) );
  NAND2_X1 U10803 ( .A1(n12790), .A2(n8612), .ZN(n9099) );
  OR2_X1 U10804 ( .A1(n14253), .A2(n12792), .ZN(n9098) );
  OR2_X1 U10805 ( .A1(n14444), .A2(n9039), .ZN(n9104) );
  INV_X1 U10806 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9191) );
  NAND2_X1 U10807 ( .A1(n9153), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U10808 ( .A1(n8599), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9100) );
  OAI211_X1 U10809 ( .C1(n9191), .C2(n8851), .A(n9101), .B(n9100), .ZN(n9102)
         );
  INV_X1 U10810 ( .A(n9102), .ZN(n9103) );
  AND2_X1 U10811 ( .A1(n9104), .A2(n9103), .ZN(n14236) );
  XNOR2_X1 U10812 ( .A(n9106), .B(n9105), .ZN(n14450) );
  INV_X1 U10813 ( .A(n14061), .ZN(n11483) );
  INV_X1 U10814 ( .A(n14047), .ZN(n11378) );
  NAND2_X1 U10815 ( .A1(n11365), .A2(n14001), .ZN(n11346) );
  INV_X1 U10816 ( .A(n14027), .ZN(n10754) );
  NAND2_X1 U10817 ( .A1(n11345), .A2(n10754), .ZN(n10778) );
  INV_X1 U10818 ( .A(n11169), .ZN(n9107) );
  NOR2_X1 U10819 ( .A1(n14611), .A2(n14596), .ZN(n14595) );
  INV_X1 U10820 ( .A(n14688), .ZN(n14577) );
  INV_X1 U10821 ( .A(n14320), .ZN(n14276) );
  AOI211_X1 U10822 ( .C1(n14234), .C2(n7507), .A(n7437), .B(n14439), .ZN(
        n14449) );
  NAND2_X1 U10823 ( .A1(n10648), .A2(n16381), .ZN(n9110) );
  NAND2_X1 U10824 ( .A1(n11350), .A2(n9110), .ZN(n10749) );
  NAND2_X1 U10825 ( .A1(n10749), .A2(n14289), .ZN(n9112) );
  INV_X1 U10826 ( .A(n14364), .ZN(n10889) );
  NAND2_X1 U10827 ( .A1(n10889), .A2(n14027), .ZN(n9111) );
  NAND2_X1 U10828 ( .A1(n9112), .A2(n9111), .ZN(n10775) );
  INV_X1 U10829 ( .A(n14363), .ZN(n10395) );
  NAND2_X1 U10830 ( .A1(n14034), .A2(n10395), .ZN(n9113) );
  INV_X1 U10831 ( .A(n14362), .ZN(n14043) );
  AND2_X1 U10832 ( .A1(n14041), .A2(n14043), .ZN(n9115) );
  OR2_X1 U10833 ( .A1(n14041), .A2(n14043), .ZN(n9114) );
  NAND2_X1 U10834 ( .A1(n14047), .A2(n11311), .ZN(n9116) );
  INV_X1 U10835 ( .A(n14295), .ZN(n11407) );
  INV_X1 U10836 ( .A(n14360), .ZN(n14057) );
  NAND2_X1 U10837 ( .A1(n14055), .A2(n14057), .ZN(n9117) );
  OR2_X1 U10838 ( .A1(n14061), .A2(n11234), .ZN(n9118) );
  NAND2_X1 U10839 ( .A1(n11608), .A2(n14297), .ZN(n11607) );
  INV_X1 U10840 ( .A(n14358), .ZN(n11632) );
  OR2_X1 U10841 ( .A1(n14629), .A2(n11632), .ZN(n9119) );
  INV_X1 U10842 ( .A(n14357), .ZN(n14075) );
  NAND2_X1 U10843 ( .A1(n14073), .A2(n14075), .ZN(n9120) );
  INV_X1 U10844 ( .A(n14356), .ZN(n11906) );
  NAND2_X1 U10845 ( .A1(n14086), .A2(n11906), .ZN(n9121) );
  OR2_X1 U10846 ( .A1(n14094), .A2(n14096), .ZN(n9123) );
  INV_X1 U10847 ( .A(n7765), .ZN(n12090) );
  INV_X1 U10848 ( .A(n14352), .ZN(n12309) );
  NAND2_X1 U10849 ( .A1(n7757), .A2(n12309), .ZN(n9125) );
  INV_X1 U10850 ( .A(n14351), .ZN(n9126) );
  NAND2_X1 U10851 ( .A1(n14122), .A2(n9126), .ZN(n9127) );
  OR2_X1 U10852 ( .A1(n14763), .A2(n14133), .ZN(n9129) );
  NAND2_X1 U10853 ( .A1(n14763), .A2(n14133), .ZN(n9130) );
  AND2_X1 U10854 ( .A1(n14698), .A2(n13901), .ZN(n9131) );
  NAND2_X1 U10855 ( .A1(n14596), .A2(n14152), .ZN(n14568) );
  AND2_X1 U10856 ( .A1(n14567), .A2(n14568), .ZN(n9132) );
  INV_X1 U10857 ( .A(n14558), .ZN(n9134) );
  OR2_X1 U10858 ( .A1(n14551), .A2(n14348), .ZN(n9135) );
  INV_X1 U10859 ( .A(n14347), .ZN(n14172) );
  NAND2_X1 U10860 ( .A1(n14675), .A2(n14172), .ZN(n9136) );
  NAND2_X1 U10861 ( .A1(n14529), .A2(n14346), .ZN(n9137) );
  NAND2_X1 U10862 ( .A1(n14521), .A2(n9137), .ZN(n9139) );
  OR2_X1 U10863 ( .A1(n14529), .A2(n14346), .ZN(n9138) );
  NAND2_X1 U10864 ( .A1(n14506), .A2(n9140), .ZN(n9142) );
  NAND2_X1 U10865 ( .A1(n14511), .A2(n13933), .ZN(n9141) );
  INV_X1 U10866 ( .A(n14344), .ZN(n13977) );
  INV_X1 U10867 ( .A(n14343), .ZN(n9143) );
  AND2_X1 U10868 ( .A1(n14482), .A2(n9143), .ZN(n9144) );
  NAND2_X1 U10869 ( .A1(n9732), .A2(n9145), .ZN(n9146) );
  NAND2_X1 U10870 ( .A1(n14323), .A2(n14320), .ZN(n14278) );
  NAND2_X1 U10871 ( .A1(n14326), .A2(n7431), .ZN(n14257) );
  AND2_X1 U10872 ( .A1(n14326), .A2(n14320), .ZN(n10487) );
  INV_X1 U10873 ( .A(n9149), .ZN(n9150) );
  INV_X1 U10874 ( .A(P2_B_REG_SCAN_IN), .ZN(n9151) );
  OR2_X1 U10875 ( .A1(n14782), .A2(n9151), .ZN(n9152) );
  AND2_X1 U10876 ( .A1(n14589), .A2(n9152), .ZN(n14432) );
  INV_X1 U10877 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14734) );
  NAND2_X1 U10878 ( .A1(n9153), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9156) );
  NAND2_X1 U10879 ( .A1(n9154), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9155) );
  OAI211_X1 U10880 ( .C1(n14219), .C2(n14734), .A(n9156), .B(n9155), .ZN(
        n14339) );
  AOI22_X1 U10881 ( .A1(n14341), .A2(n14588), .B1(n14432), .B2(n14339), .ZN(
        n9157) );
  NAND2_X1 U10882 ( .A1(n9159), .A2(n9158), .ZN(n9174) );
  INV_X1 U10883 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9161) );
  INV_X1 U10884 ( .A(n9166), .ZN(n9163) );
  NAND2_X1 U10885 ( .A1(n9163), .A2(n9162), .ZN(n9167) );
  NAND2_X1 U10886 ( .A1(n9167), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9164) );
  XNOR2_X1 U10887 ( .A(n9165), .B(P2_IR_REG_24__SCAN_IN), .ZN(n9188) );
  INV_X1 U10888 ( .A(n9188), .ZN(n12189) );
  NAND2_X1 U10889 ( .A1(n9166), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n9168) );
  NAND2_X1 U10890 ( .A1(n9168), .A2(n9167), .ZN(n12222) );
  OAI221_X1 U10891 ( .B1(n9188), .B2(P2_B_REG_SCAN_IN), .C1(n12189), .C2(n9151), .A(n12222), .ZN(n9169) );
  INV_X1 U10892 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15818) );
  NAND2_X1 U10893 ( .A1(n15819), .A2(n15818), .ZN(n9172) );
  INV_X1 U10894 ( .A(n12222), .ZN(n9170) );
  OR2_X1 U10895 ( .A1(n14785), .A2(n9170), .ZN(n9171) );
  AND2_X1 U10896 ( .A1(n9172), .A2(n9171), .ZN(n10357) );
  NOR2_X1 U10897 ( .A1(n12222), .A2(n12189), .ZN(n9173) );
  NAND2_X1 U10898 ( .A1(n14785), .A2(n9173), .ZN(n10618) );
  NAND2_X1 U10899 ( .A1(n9174), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9176) );
  INV_X1 U10900 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9175) );
  XNOR2_X1 U10901 ( .A(n9176), .B(n9175), .ZN(n10486) );
  NAND2_X1 U10902 ( .A1(n10618), .A2(n10486), .ZN(n10390) );
  NOR2_X1 U10903 ( .A1(n10357), .A2(n15822), .ZN(n15817) );
  NOR4_X1 U10904 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9180) );
  NOR4_X1 U10905 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9179) );
  NOR4_X1 U10906 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9178) );
  NOR4_X1 U10907 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9177) );
  NAND4_X1 U10908 ( .A1(n9180), .A2(n9179), .A3(n9178), .A4(n9177), .ZN(n9186)
         );
  NOR2_X1 U10909 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n9184) );
  NOR4_X1 U10910 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9183) );
  NOR4_X1 U10911 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9182) );
  NOR4_X1 U10912 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n9181) );
  NAND4_X1 U10913 ( .A1(n9184), .A2(n9183), .A3(n9182), .A4(n9181), .ZN(n9185)
         );
  OAI21_X1 U10914 ( .B1(n9186), .B2(n9185), .A(n15819), .ZN(n10358) );
  NAND2_X1 U10915 ( .A1(n16558), .A2(n14276), .ZN(n10386) );
  NAND2_X1 U10916 ( .A1(n14286), .A2(n14424), .ZN(n10396) );
  AND2_X1 U10917 ( .A1(n10396), .A2(n14320), .ZN(n14259) );
  NAND2_X1 U10918 ( .A1(n14259), .A2(n14326), .ZN(n10388) );
  AND2_X1 U10919 ( .A1(n10386), .A2(n10388), .ZN(n9187) );
  INV_X1 U10920 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15823) );
  NAND2_X1 U10921 ( .A1(n15819), .A2(n15823), .ZN(n9190) );
  OR2_X1 U10922 ( .A1(n14785), .A2(n9188), .ZN(n9189) );
  INV_X1 U10923 ( .A(n9192), .ZN(n9193) );
  OAI21_X1 U10924 ( .B1(n9727), .B2(n16559), .A(n9193), .ZN(P2_U3528) );
  INV_X2 U10925 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n13770) );
  NAND2_X1 U10926 ( .A1(n9456), .A2(n9195), .ZN(n9498) );
  NOR2_X1 U10927 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n9199) );
  NAND4_X1 U10928 ( .A1(n9199), .A2(n9198), .A3(n9197), .A4(n9196), .ZN(n9200)
         );
  INV_X1 U10929 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9203) );
  XNOR2_X2 U10930 ( .A(n9204), .B(n9203), .ZN(n15772) );
  NAND2_X1 U10931 ( .A1(n9205), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9206) );
  MUX2_X1 U10932 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9206), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n9207) );
  NAND2_X2 U10933 ( .A1(n9207), .A2(n9210), .ZN(n15885) );
  NAND2_X1 U10934 ( .A1(n12221), .A2(n15206), .ZN(n9209) );
  NAND2_X1 U10935 ( .A1(n7459), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9208) );
  INV_X1 U10936 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9213) );
  XNOR2_X2 U10937 ( .A(n9212), .B(n9211), .ZN(n15767) );
  INV_X4 U10938 ( .A(n9282), .ZN(n9607) );
  NAND2_X1 U10939 ( .A1(n9607), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9224) );
  INV_X1 U10940 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9215) );
  OR2_X1 U10941 ( .A1(n9477), .A2(n9215), .ZN(n9223) );
  NAND2_X1 U10942 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9309) );
  NAND2_X1 U10943 ( .A1(n9369), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9401) );
  INV_X1 U10944 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9400) );
  INV_X1 U10945 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9416) );
  INV_X1 U10946 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9447) );
  INV_X1 U10947 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n11498) );
  INV_X1 U10948 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9489) );
  INV_X1 U10949 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9504) );
  INV_X1 U10950 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9517) );
  OAI21_X1 U10951 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n9218), .A(n9572), .ZN(
        n15487) );
  OR2_X1 U10952 ( .A1(n7814), .A2(n15487), .ZN(n9222) );
  INV_X1 U10953 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9220) );
  OR2_X1 U10954 ( .A1(n7778), .A2(n9220), .ZN(n9221) );
  NAND4_X1 U10955 ( .A1(n9224), .A2(n9223), .A3(n9222), .A4(n9221), .ZN(n15304) );
  NAND2_X1 U10956 ( .A1(n12104), .A2(n15206), .ZN(n9226) );
  NAND2_X1 U10957 ( .A1(n7459), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9225) );
  INV_X1 U10958 ( .A(n15675), .ZN(n9568) );
  NAND2_X1 U10959 ( .A1(n9607), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9234) );
  INV_X1 U10960 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9227) );
  OR2_X1 U10961 ( .A1(n9477), .A2(n9227), .ZN(n9233) );
  OAI21_X1 U10962 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n9229), .A(n9228), .ZN(
        n15502) );
  OR2_X1 U10963 ( .A1(n7814), .A2(n15502), .ZN(n9232) );
  INV_X1 U10964 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9230) );
  OR2_X1 U10965 ( .A1(n7778), .A2(n9230), .ZN(n9231) );
  NAND4_X1 U10966 ( .A1(n9234), .A2(n9233), .A3(n9232), .A4(n9231), .ZN(n15305) );
  OR2_X1 U10967 ( .A1(n9547), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U10968 ( .A1(n9238), .A2(n9237), .ZN(n15532) );
  INV_X1 U10969 ( .A(n15532), .ZN(n15000) );
  INV_X1 U10970 ( .A(n7814), .ZN(n9239) );
  NAND2_X1 U10971 ( .A1(n15000), .A2(n9239), .ZN(n9245) );
  INV_X1 U10972 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9242) );
  NAND2_X1 U10973 ( .A1(n7818), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9241) );
  NAND2_X1 U10974 ( .A1(n9254), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n9240) );
  OAI211_X1 U10975 ( .C1(n9634), .C2(n9242), .A(n9241), .B(n9240), .ZN(n9243)
         );
  INV_X1 U10976 ( .A(n9243), .ZN(n9244) );
  NAND2_X1 U10977 ( .A1(n7457), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9251) );
  INV_X1 U10978 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11579) );
  INV_X1 U10979 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9246) );
  INV_X1 U10980 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9247) );
  OR2_X1 U10981 ( .A1(n9282), .A2(n9247), .ZN(n9248) );
  INV_X1 U10982 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n15887) );
  NAND2_X1 U10983 ( .A1(n9253), .A2(n9252), .ZN(n15784) );
  MUX2_X1 U10984 ( .A(n15887), .B(n15784), .S(n9261), .Z(n16327) );
  OR2_X1 U10985 ( .A1(n11576), .A2(n16327), .ZN(n16331) );
  NAND2_X1 U10986 ( .A1(n9254), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9259) );
  INV_X1 U10987 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9255) );
  INV_X1 U10988 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9256) );
  OR2_X1 U10989 ( .A1(n9282), .A2(n9256), .ZN(n9257) );
  INV_X1 U10990 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n15332) );
  INV_X1 U10991 ( .A(n10413), .ZN(n9260) );
  NAND2_X1 U10992 ( .A1(n9318), .A2(n9260), .ZN(n9267) );
  NAND2_X1 U10993 ( .A1(n9287), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9266) );
  INV_X4 U10994 ( .A(n9261), .ZN(n10577) );
  NAND2_X1 U10995 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9262) );
  MUX2_X1 U10996 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9262), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9264) );
  INV_X1 U10997 ( .A(n9263), .ZN(n9274) );
  NAND2_X1 U10998 ( .A1(n9264), .A2(n9274), .ZN(n15336) );
  INV_X1 U10999 ( .A(n15336), .ZN(n15335) );
  NAND2_X1 U11000 ( .A1(n10577), .A2(n15335), .ZN(n9265) );
  AND3_X2 U11001 ( .A1(n9267), .A2(n9266), .A3(n9265), .ZN(n16339) );
  INV_X1 U11002 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n15355) );
  OR2_X1 U11003 ( .A1(n9477), .A2(n15355), .ZN(n9273) );
  INV_X1 U11004 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n11992) );
  NAND2_X1 U11005 ( .A1(n9607), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9271) );
  INV_X1 U11006 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10591) );
  NAND2_X1 U11007 ( .A1(n9287), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9280) );
  NAND2_X1 U11008 ( .A1(n9274), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9275) );
  MUX2_X1 U11009 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9275), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n9277) );
  NAND2_X1 U11010 ( .A1(n9277), .A2(n9276), .ZN(n15354) );
  INV_X1 U11011 ( .A(n15354), .ZN(n15351) );
  NAND2_X1 U11012 ( .A1(n10577), .A2(n15351), .ZN(n9279) );
  NAND2_X1 U11013 ( .A1(n10409), .A2(n9318), .ZN(n9278) );
  NAND2_X1 U11014 ( .A1(n9639), .A2(n16374), .ZN(n15049) );
  NAND2_X1 U11015 ( .A1(n11987), .A2(n11988), .ZN(n11986) );
  NAND2_X1 U11016 ( .A1(n11986), .A2(n15046), .ZN(n12115) );
  NAND2_X1 U11017 ( .A1(n7818), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9286) );
  OR2_X1 U11018 ( .A1(n7814), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9285) );
  INV_X1 U11019 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10592) );
  OR2_X1 U11020 ( .A1(n15195), .A2(n10592), .ZN(n9284) );
  INV_X1 U11021 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9281) );
  OR2_X1 U11022 ( .A1(n9282), .A2(n9281), .ZN(n9283) );
  NAND4_X2 U11023 ( .A1(n9286), .A2(n9285), .A3(n9284), .A4(n9283), .ZN(n15326) );
  NAND2_X1 U11024 ( .A1(n9276), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9289) );
  MUX2_X1 U11025 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9289), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9290) );
  AND2_X1 U11026 ( .A1(n9288), .A2(n9290), .ZN(n15364) );
  AOI22_X1 U11027 ( .A1(n9287), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n10577), 
        .B2(n15364), .ZN(n9291) );
  NAND2_X1 U11028 ( .A1(n15326), .A2(n9625), .ZN(n15048) );
  INV_X1 U11029 ( .A(n15042), .ZN(n9292) );
  AOI21_X1 U11030 ( .B1(n12115), .B2(n15048), .A(n9292), .ZN(n12064) );
  NAND2_X1 U11031 ( .A1(n9288), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9293) );
  XNOR2_X1 U11032 ( .A(n9293), .B(P1_IR_REG_4__SCAN_IN), .ZN(n16288) );
  AOI22_X1 U11033 ( .A1(n7460), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n10577), 
        .B2(n16288), .ZN(n9295) );
  NAND2_X1 U11034 ( .A1(n10417), .A2(n9318), .ZN(n9294) );
  NAND2_X1 U11035 ( .A1(n9607), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9299) );
  INV_X1 U11036 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10570) );
  OR2_X1 U11037 ( .A1(n9477), .A2(n10570), .ZN(n9298) );
  INV_X1 U11038 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10595) );
  OR2_X1 U11039 ( .A1(n15195), .A2(n10595), .ZN(n9297) );
  OAI21_X1 U11040 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9309), .ZN(n12058) );
  OR2_X1 U11041 ( .A1(n9311), .A2(n12058), .ZN(n9296) );
  INV_X1 U11042 ( .A(n15056), .ZN(n15325) );
  NAND2_X1 U11043 ( .A1(n15325), .A2(n15055), .ZN(n9300) );
  NAND2_X1 U11044 ( .A1(n10443), .A2(n9318), .ZN(n9305) );
  INV_X1 U11045 ( .A(n9301), .ZN(n9302) );
  NAND2_X1 U11046 ( .A1(n9302), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9303) );
  XNOR2_X1 U11047 ( .A(n9303), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10599) );
  AOI22_X1 U11048 ( .A1(n7459), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n10577), 
        .B2(n10599), .ZN(n9304) );
  NAND2_X1 U11049 ( .A1(n9305), .A2(n9304), .ZN(n16448) );
  NAND2_X1 U11050 ( .A1(n9607), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9316) );
  INV_X1 U11051 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9306) );
  OR2_X1 U11052 ( .A1(n9477), .A2(n9306), .ZN(n9315) );
  INV_X1 U11053 ( .A(n9307), .ZN(n9325) );
  NAND2_X1 U11054 ( .A1(n9309), .A2(n9308), .ZN(n9310) );
  NAND2_X1 U11055 ( .A1(n9325), .A2(n9310), .ZN(n16449) );
  OR2_X1 U11056 ( .A1(n7814), .A2(n16449), .ZN(n9314) );
  INV_X1 U11057 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9312) );
  OR2_X1 U11058 ( .A1(n15195), .A2(n9312), .ZN(n9313) );
  NAND4_X1 U11059 ( .A1(n9316), .A2(n9315), .A3(n9314), .A4(n9313), .ZN(n15324) );
  INV_X1 U11060 ( .A(n15324), .ZN(n11467) );
  NAND2_X1 U11061 ( .A1(n16448), .A2(n11467), .ZN(n9317) );
  AOI21_X2 U11062 ( .B1(n16435), .B2(n9317), .A(n7530), .ZN(n11974) );
  NAND2_X1 U11063 ( .A1(n10447), .A2(n9318), .ZN(n9322) );
  INV_X1 U11064 ( .A(n9500), .ZN(n9319) );
  NAND2_X1 U11065 ( .A1(n9319), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9320) );
  XNOR2_X1 U11066 ( .A(n9320), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10601) );
  AOI22_X1 U11067 ( .A1(n7460), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n10577), 
        .B2(n10601), .ZN(n9321) );
  NAND2_X1 U11068 ( .A1(n9322), .A2(n9321), .ZN(n16465) );
  NAND2_X1 U11069 ( .A1(n7818), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9331) );
  INV_X1 U11070 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9323) );
  OR2_X1 U11071 ( .A1(n7778), .A2(n9323), .ZN(n9330) );
  INV_X1 U11072 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9324) );
  NAND2_X1 U11073 ( .A1(n9325), .A2(n9324), .ZN(n9326) );
  NAND2_X1 U11074 ( .A1(n9341), .A2(n9326), .ZN(n11979) );
  OR2_X1 U11075 ( .A1(n7814), .A2(n11979), .ZN(n9329) );
  INV_X1 U11076 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9327) );
  OR2_X1 U11077 ( .A1(n9634), .A2(n9327), .ZN(n9328) );
  NAND4_X1 U11078 ( .A1(n9331), .A2(n9330), .A3(n9329), .A4(n9328), .ZN(n15323) );
  NAND2_X1 U11079 ( .A1(n16465), .A2(n11466), .ZN(n9334) );
  OR2_X1 U11080 ( .A1(n16465), .A2(n11466), .ZN(n9332) );
  NAND2_X1 U11081 ( .A1(n9334), .A2(n9332), .ZN(n15238) );
  NAND2_X1 U11082 ( .A1(n11974), .A2(n9333), .ZN(n11973) );
  NAND2_X1 U11083 ( .A1(n11973), .A2(n9334), .ZN(n16478) );
  NAND2_X1 U11084 ( .A1(n10455), .A2(n15206), .ZN(n9338) );
  NAND2_X1 U11085 ( .A1(n9500), .A2(n9335), .ZN(n9350) );
  NAND2_X1 U11086 ( .A1(n9350), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9336) );
  XNOR2_X1 U11087 ( .A(n9336), .B(P1_IR_REG_7__SCAN_IN), .ZN(n15385) );
  AOI22_X1 U11088 ( .A1(n7459), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n10577), 
        .B2(n15385), .ZN(n9337) );
  NAND2_X1 U11089 ( .A1(n9338), .A2(n9337), .ZN(n15074) );
  NAND2_X1 U11090 ( .A1(n9607), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9346) );
  INV_X1 U11091 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9339) );
  OR2_X1 U11092 ( .A1(n9477), .A2(n9339), .ZN(n9345) );
  NAND2_X1 U11093 ( .A1(n9341), .A2(n9340), .ZN(n9342) );
  NAND2_X1 U11094 ( .A1(n9356), .A2(n9342), .ZN(n16489) );
  OR2_X1 U11095 ( .A1(n7814), .A2(n16489), .ZN(n9344) );
  INV_X1 U11096 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10602) );
  OR2_X1 U11097 ( .A1(n7778), .A2(n10602), .ZN(n9343) );
  NAND4_X1 U11098 ( .A1(n9346), .A2(n9345), .A3(n9344), .A4(n9343), .ZN(n15322) );
  OR2_X1 U11099 ( .A1(n15074), .A2(n11768), .ZN(n9347) );
  NAND2_X1 U11100 ( .A1(n16478), .A2(n9347), .ZN(n9349) );
  NAND2_X1 U11101 ( .A1(n15074), .A2(n11768), .ZN(n9348) );
  NAND2_X1 U11102 ( .A1(n9349), .A2(n9348), .ZN(n11766) );
  INV_X1 U11103 ( .A(n11766), .ZN(n9362) );
  NAND2_X1 U11104 ( .A1(n10459), .A2(n15206), .ZN(n9353) );
  NAND2_X1 U11105 ( .A1(n9364), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9351) );
  XNOR2_X1 U11106 ( .A(n9351), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10660) );
  AOI22_X1 U11107 ( .A1(n7459), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n10577), 
        .B2(n10660), .ZN(n9352) );
  NAND2_X1 U11108 ( .A1(n9353), .A2(n9352), .ZN(n15078) );
  NAND2_X1 U11109 ( .A1(n9607), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9361) );
  INV_X1 U11110 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10573) );
  OR2_X1 U11111 ( .A1(n9477), .A2(n10573), .ZN(n9360) );
  INV_X1 U11112 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9354) );
  OR2_X1 U11113 ( .A1(n7778), .A2(n9354), .ZN(n9359) );
  NAND2_X1 U11114 ( .A1(n9356), .A2(n9355), .ZN(n9357) );
  NAND2_X1 U11115 ( .A1(n9371), .A2(n9357), .ZN(n16507) );
  OR2_X1 U11116 ( .A1(n7814), .A2(n16507), .ZN(n9358) );
  NAND4_X1 U11117 ( .A1(n9361), .A2(n9360), .A3(n9359), .A4(n9358), .ZN(n15321) );
  XNOR2_X1 U11118 ( .A(n15078), .B(n15321), .ZN(n15240) );
  NAND2_X1 U11119 ( .A1(n9362), .A2(n15240), .ZN(n11770) );
  INV_X1 U11120 ( .A(n15321), .ZN(n11782) );
  OR2_X1 U11121 ( .A1(n15078), .A2(n11782), .ZN(n9363) );
  NAND2_X1 U11122 ( .A1(n11770), .A2(n9363), .ZN(n12013) );
  NAND2_X1 U11123 ( .A1(n10472), .A2(n15206), .ZN(n9367) );
  NAND2_X1 U11124 ( .A1(n9381), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9365) );
  XNOR2_X1 U11125 ( .A(n9365), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U11126 ( .A1(n7459), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n10577), 
        .B2(n10606), .ZN(n9366) );
  NAND2_X1 U11127 ( .A1(n9607), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9377) );
  INV_X1 U11128 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9368) );
  OR2_X1 U11129 ( .A1(n9477), .A2(n9368), .ZN(n9376) );
  INV_X1 U11130 ( .A(n9369), .ZN(n9385) );
  NAND2_X1 U11131 ( .A1(n9371), .A2(n9370), .ZN(n9372) );
  NAND2_X1 U11132 ( .A1(n9385), .A2(n9372), .ZN(n12215) );
  OR2_X1 U11133 ( .A1(n7814), .A2(n12215), .ZN(n9375) );
  INV_X1 U11134 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9373) );
  OR2_X1 U11135 ( .A1(n7778), .A2(n9373), .ZN(n9374) );
  NAND4_X1 U11136 ( .A1(n9377), .A2(n9376), .A3(n9375), .A4(n9374), .ZN(n15320) );
  INV_X1 U11137 ( .A(n15320), .ZN(n12039) );
  NAND2_X1 U11138 ( .A1(n16531), .A2(n12039), .ZN(n9378) );
  NAND2_X1 U11139 ( .A1(n12013), .A2(n9378), .ZN(n9380) );
  OR2_X1 U11140 ( .A1(n16531), .A2(n12039), .ZN(n9379) );
  NAND2_X1 U11141 ( .A1(n9380), .A2(n9379), .ZN(n11957) );
  NAND2_X1 U11142 ( .A1(n10477), .A2(n15206), .ZN(n9383) );
  XNOR2_X1 U11143 ( .A(n9395), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10759) );
  AOI22_X1 U11144 ( .A1(n7459), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n10577), 
        .B2(n10759), .ZN(n9382) );
  NAND2_X1 U11145 ( .A1(n9607), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n9391) );
  INV_X1 U11146 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n12072) );
  OR2_X1 U11147 ( .A1(n9477), .A2(n12072), .ZN(n9390) );
  INV_X1 U11148 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9384) );
  NAND2_X1 U11149 ( .A1(n9385), .A2(n9384), .ZN(n9386) );
  NAND2_X1 U11150 ( .A1(n9401), .A2(n9386), .ZN(n12071) );
  OR2_X1 U11151 ( .A1(n7814), .A2(n12071), .ZN(n9389) );
  INV_X1 U11152 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9387) );
  OR2_X1 U11153 ( .A1(n7778), .A2(n9387), .ZN(n9388) );
  NAND4_X1 U11154 ( .A1(n9391), .A2(n9390), .A3(n9389), .A4(n9388), .ZN(n15319) );
  INV_X1 U11155 ( .A(n15319), .ZN(n12048) );
  XNOR2_X1 U11156 ( .A(n15090), .B(n12048), .ZN(n15245) );
  INV_X1 U11157 ( .A(n15245), .ZN(n9392) );
  NAND2_X1 U11158 ( .A1(n11957), .A2(n9392), .ZN(n9394) );
  OR2_X1 U11159 ( .A1(n15090), .A2(n12048), .ZN(n9393) );
  NAND2_X1 U11160 ( .A1(n9394), .A2(n9393), .ZN(n12173) );
  NAND2_X1 U11161 ( .A1(n10541), .A2(n15206), .ZN(n9398) );
  NAND2_X1 U11162 ( .A1(n9395), .A2(n13584), .ZN(n9396) );
  NAND2_X1 U11163 ( .A1(n9396), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9410) );
  XNOR2_X1 U11164 ( .A(n9410), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10728) );
  AOI22_X1 U11165 ( .A1(n10728), .A2(n10577), .B1(n7460), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n9397) );
  NAND2_X1 U11166 ( .A1(n9607), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9407) );
  INV_X1 U11167 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9399) );
  OR2_X1 U11168 ( .A1(n9477), .A2(n9399), .ZN(n9406) );
  NAND2_X1 U11169 ( .A1(n9401), .A2(n9400), .ZN(n9402) );
  NAND2_X1 U11170 ( .A1(n9417), .A2(n9402), .ZN(n12257) );
  OR2_X1 U11171 ( .A1(n7814), .A2(n12257), .ZN(n9405) );
  INV_X1 U11172 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9403) );
  OR2_X1 U11173 ( .A1(n7778), .A2(n9403), .ZN(n9404) );
  NAND4_X1 U11174 ( .A1(n9407), .A2(n9406), .A3(n9405), .A4(n9404), .ZN(n15318) );
  INV_X1 U11175 ( .A(n15318), .ZN(n12246) );
  NOR2_X1 U11176 ( .A1(n16572), .A2(n12246), .ZN(n9409) );
  NAND2_X1 U11177 ( .A1(n16572), .A2(n12246), .ZN(n9408) );
  OAI21_X2 U11178 ( .B1(n12173), .B2(n9409), .A(n9408), .ZN(n12166) );
  INV_X1 U11179 ( .A(n12166), .ZN(n9425) );
  NAND2_X1 U11180 ( .A1(n10654), .A2(n15206), .ZN(n9413) );
  NAND2_X1 U11181 ( .A1(n9410), .A2(n13589), .ZN(n9411) );
  NAND2_X1 U11182 ( .A1(n9411), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9427) );
  XNOR2_X1 U11183 ( .A(n9427), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10914) );
  AOI22_X1 U11184 ( .A1(n10914), .A2(n10577), .B1(n7460), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n9412) );
  NAND2_X1 U11185 ( .A1(n9607), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9423) );
  INV_X1 U11186 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9414) );
  OR2_X1 U11187 ( .A1(n9477), .A2(n9414), .ZN(n9422) );
  INV_X1 U11188 ( .A(n9415), .ZN(n9433) );
  NAND2_X1 U11189 ( .A1(n9417), .A2(n9416), .ZN(n9418) );
  NAND2_X1 U11190 ( .A1(n9433), .A2(n9418), .ZN(n14942) );
  OR2_X1 U11191 ( .A1(n7814), .A2(n14942), .ZN(n9421) );
  INV_X1 U11192 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9419) );
  OR2_X1 U11193 ( .A1(n7778), .A2(n9419), .ZN(n9420) );
  NAND4_X1 U11194 ( .A1(n9423), .A2(n9422), .A3(n9421), .A4(n9420), .ZN(n15317) );
  INV_X1 U11195 ( .A(n15317), .ZN(n12467) );
  XNOR2_X1 U11196 ( .A(n15101), .B(n12467), .ZN(n15246) );
  OR2_X1 U11197 ( .A1(n15101), .A2(n12467), .ZN(n9426) );
  AND2_X2 U11198 ( .A1(n12165), .A2(n9426), .ZN(n12298) );
  NAND2_X1 U11199 ( .A1(n10782), .A2(n15206), .ZN(n9430) );
  NAND2_X1 U11200 ( .A1(n9427), .A2(n7454), .ZN(n9428) );
  NAND2_X1 U11201 ( .A1(n9428), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9442) );
  XNOR2_X1 U11202 ( .A(n9442), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10930) );
  AOI22_X1 U11203 ( .A1(n10930), .A2(n10577), .B1(n7460), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n9429) );
  NAND2_X1 U11204 ( .A1(n7818), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9439) );
  INV_X1 U11205 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9431) );
  OR2_X1 U11206 ( .A1(n7778), .A2(n9431), .ZN(n9438) );
  INV_X1 U11207 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9432) );
  NAND2_X1 U11208 ( .A1(n9433), .A2(n9432), .ZN(n9434) );
  NAND2_X1 U11209 ( .A1(n9448), .A2(n9434), .ZN(n12482) );
  OR2_X1 U11210 ( .A1(n7814), .A2(n12482), .ZN(n9437) );
  INV_X1 U11211 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9435) );
  OR2_X1 U11212 ( .A1(n9634), .A2(n9435), .ZN(n9436) );
  NAND4_X1 U11213 ( .A1(n9439), .A2(n9438), .A3(n9437), .A4(n9436), .ZN(n15316) );
  INV_X1 U11214 ( .A(n15316), .ZN(n12488) );
  XNOR2_X1 U11215 ( .A(n15105), .B(n12488), .ZN(n15247) );
  INV_X1 U11216 ( .A(n15247), .ZN(n12297) );
  NAND2_X1 U11217 ( .A1(n12298), .A2(n12297), .ZN(n12296) );
  NAND2_X1 U11218 ( .A1(n15105), .A2(n12488), .ZN(n9440) );
  NAND2_X1 U11219 ( .A1(n12296), .A2(n9440), .ZN(n12486) );
  NAND2_X1 U11220 ( .A1(n11062), .A2(n15206), .ZN(n9446) );
  NAND2_X1 U11221 ( .A1(n9442), .A2(n9441), .ZN(n9443) );
  NAND2_X1 U11222 ( .A1(n9443), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9444) );
  XNOR2_X1 U11223 ( .A(n9444), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U11224 ( .A1(n11487), .A2(n10577), .B1(n7460), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9445) );
  NAND2_X2 U11225 ( .A1(n9446), .A2(n9445), .ZN(n16611) );
  NAND2_X1 U11226 ( .A1(n9607), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9453) );
  INV_X1 U11227 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11489) );
  OR2_X1 U11228 ( .A1(n9477), .A2(n11489), .ZN(n9452) );
  INV_X1 U11229 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11494) );
  OR2_X1 U11230 ( .A1(n7778), .A2(n11494), .ZN(n9451) );
  NAND2_X1 U11231 ( .A1(n9448), .A2(n9447), .ZN(n9449) );
  NAND2_X1 U11232 ( .A1(n9464), .A2(n9449), .ZN(n16618) );
  OR2_X1 U11233 ( .A1(n7814), .A2(n16618), .ZN(n9450) );
  NAND4_X1 U11234 ( .A1(n9453), .A2(n9452), .A3(n9451), .A4(n9450), .ZN(n15315) );
  XNOR2_X1 U11235 ( .A(n16611), .B(n15315), .ZN(n15248) );
  NAND2_X1 U11236 ( .A1(n12486), .A2(n15248), .ZN(n9455) );
  INV_X1 U11237 ( .A(n15315), .ZN(n14805) );
  NAND2_X1 U11238 ( .A1(n16611), .A2(n14805), .ZN(n9454) );
  NAND2_X1 U11239 ( .A1(n9455), .A2(n9454), .ZN(n12509) );
  NAND2_X1 U11240 ( .A1(n9500), .A2(n9456), .ZN(n9458) );
  NAND2_X1 U11241 ( .A1(n9458), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9457) );
  MUX2_X1 U11242 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9457), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n9459) );
  OR2_X1 U11243 ( .A1(n9458), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n9485) );
  AND2_X1 U11244 ( .A1(n9459), .A2(n9485), .ZN(n15404) );
  AOI22_X1 U11245 ( .A1(n7460), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n10577), 
        .B2(n15404), .ZN(n9460) );
  NAND2_X1 U11246 ( .A1(n9607), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n9470) );
  INV_X1 U11247 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9462) );
  OR2_X1 U11248 ( .A1(n9477), .A2(n9462), .ZN(n9469) );
  INV_X1 U11249 ( .A(n9463), .ZN(n9479) );
  NAND2_X1 U11250 ( .A1(n9464), .A2(n11498), .ZN(n9465) );
  NAND2_X1 U11251 ( .A1(n9479), .A2(n9465), .ZN(n15026) );
  OR2_X1 U11252 ( .A1(n7814), .A2(n15026), .ZN(n9468) );
  INV_X1 U11253 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9466) );
  OR2_X1 U11254 ( .A1(n7778), .A2(n9466), .ZN(n9467) );
  NAND4_X1 U11255 ( .A1(n9470), .A2(n9469), .A3(n9468), .A4(n9467), .ZN(n15314) );
  INV_X1 U11256 ( .A(n15314), .ZN(n12487) );
  OR2_X1 U11257 ( .A1(n15732), .A2(n12487), .ZN(n9471) );
  NAND2_X1 U11258 ( .A1(n11473), .A2(n15206), .ZN(n9474) );
  NAND2_X1 U11259 ( .A1(n9485), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9472) );
  XNOR2_X1 U11260 ( .A(n9472), .B(P1_IR_REG_16__SCAN_IN), .ZN(n15407) );
  AOI22_X1 U11261 ( .A1(n7460), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n10577), 
        .B2(n15407), .ZN(n9473) );
  INV_X1 U11262 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9476) );
  NAND2_X1 U11263 ( .A1(n9607), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9475) );
  OAI21_X1 U11264 ( .B1(n9477), .B2(n9476), .A(n9475), .ZN(n9483) );
  INV_X1 U11265 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9478) );
  NAND2_X1 U11266 ( .A1(n9479), .A2(n9478), .ZN(n9480) );
  NAND2_X1 U11267 ( .A1(n9490), .A2(n9480), .ZN(n15634) );
  NOR2_X1 U11268 ( .A1(n15634), .A2(n7814), .ZN(n9482) );
  INV_X1 U11269 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n15397) );
  NOR2_X1 U11270 ( .A1(n7778), .A2(n15397), .ZN(n9481) );
  XNOR2_X1 U11271 ( .A(n15725), .B(n15313), .ZN(n15625) );
  INV_X1 U11272 ( .A(n15313), .ZN(n14819) );
  NAND2_X1 U11273 ( .A1(n15725), .A2(n14819), .ZN(n9484) );
  NAND2_X1 U11274 ( .A1(n15624), .A2(n9484), .ZN(n15610) );
  NAND2_X1 U11275 ( .A1(n11546), .A2(n15206), .ZN(n9488) );
  OAI21_X1 U11276 ( .B1(n9485), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9486) );
  XNOR2_X1 U11277 ( .A(n9486), .B(P1_IR_REG_17__SCAN_IN), .ZN(n15403) );
  AOI22_X1 U11278 ( .A1(n7459), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n10577), 
        .B2(n15403), .ZN(n9487) );
  INV_X1 U11279 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n15398) );
  NAND2_X1 U11280 ( .A1(n9490), .A2(n9489), .ZN(n9491) );
  NAND2_X1 U11281 ( .A1(n9505), .A2(n9491), .ZN(n15616) );
  OR2_X1 U11282 ( .A1(n15616), .A2(n7814), .ZN(n9496) );
  INV_X1 U11283 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15615) );
  OR2_X1 U11284 ( .A1(n9477), .A2(n15615), .ZN(n9494) );
  INV_X1 U11285 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9492) );
  OR2_X1 U11286 ( .A1(n9634), .A2(n9492), .ZN(n9493) );
  AND2_X1 U11287 ( .A1(n9494), .A2(n9493), .ZN(n9495) );
  OAI211_X1 U11288 ( .C1(n7778), .C2(n15398), .A(n9496), .B(n9495), .ZN(n15312) );
  INV_X1 U11289 ( .A(n15312), .ZN(n14829) );
  XNOR2_X1 U11290 ( .A(n15715), .B(n14829), .ZN(n15611) );
  INV_X1 U11291 ( .A(n15611), .ZN(n9662) );
  NAND2_X1 U11292 ( .A1(n15715), .A2(n14829), .ZN(n9497) );
  NAND2_X1 U11293 ( .A1(n11585), .A2(n15206), .ZN(n9503) );
  NAND2_X1 U11294 ( .A1(n9509), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9501) );
  XNOR2_X1 U11295 ( .A(n9501), .B(P1_IR_REG_18__SCAN_IN), .ZN(n15410) );
  AOI22_X1 U11296 ( .A1(n7459), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10577), 
        .B2(n15410), .ZN(n9502) );
  NAND2_X1 U11297 ( .A1(n9505), .A2(n9504), .ZN(n9506) );
  NAND2_X1 U11298 ( .A1(n9518), .A2(n9506), .ZN(n15594) );
  AOI22_X1 U11299 ( .A1(n9607), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n7818), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n9508) );
  NAND2_X1 U11300 ( .A1(n9254), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9507) );
  OAI211_X1 U11301 ( .C1(n15594), .C2(n7814), .A(n9508), .B(n9507), .ZN(n15311) );
  INV_X1 U11302 ( .A(n15311), .ZN(n9527) );
  XNOR2_X1 U11303 ( .A(n15710), .B(n9527), .ZN(n15601) );
  NAND2_X1 U11304 ( .A1(n11600), .A2(n15206), .ZN(n9515) );
  INV_X1 U11305 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9510) );
  MUX2_X1 U11306 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9512), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n9513) );
  INV_X1 U11307 ( .A(n9614), .ZN(n9622) );
  NAND2_X1 U11308 ( .A1(n9513), .A2(n9622), .ZN(n15417) );
  INV_X1 U11309 ( .A(n15417), .ZN(n11573) );
  AOI22_X1 U11310 ( .A1(n7459), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n11573), 
        .B2(n10577), .ZN(n9514) );
  INV_X1 U11311 ( .A(n9516), .ZN(n9533) );
  NAND2_X1 U11312 ( .A1(n9518), .A2(n9517), .ZN(n9519) );
  NAND2_X1 U11313 ( .A1(n9533), .A2(n9519), .ZN(n15576) );
  OR2_X1 U11314 ( .A1(n15576), .A2(n7814), .ZN(n9524) );
  INV_X1 U11315 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n15401) );
  NAND2_X1 U11316 ( .A1(n9607), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9521) );
  NAND2_X1 U11317 ( .A1(n7818), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9520) );
  OAI211_X1 U11318 ( .C1(n15401), .C2(n7778), .A(n9521), .B(n9520), .ZN(n9522)
         );
  INV_X1 U11319 ( .A(n9522), .ZN(n9523) );
  NAND2_X1 U11320 ( .A1(n9524), .A2(n9523), .ZN(n15310) );
  INV_X1 U11321 ( .A(n15310), .ZN(n9525) );
  NAND2_X1 U11322 ( .A1(n15703), .A2(n9525), .ZN(n9529) );
  OR2_X1 U11323 ( .A1(n15703), .A2(n9525), .ZN(n9526) );
  NAND2_X1 U11324 ( .A1(n9529), .A2(n9526), .ZN(n15580) );
  NOR2_X1 U11325 ( .A1(n15710), .A2(n9527), .ZN(n15581) );
  NOR2_X1 U11326 ( .A1(n15580), .A2(n15581), .ZN(n9528) );
  NAND2_X1 U11327 ( .A1(n11616), .A2(n15206), .ZN(n9531) );
  NAND2_X1 U11328 ( .A1(n7460), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9530) );
  INV_X1 U11329 ( .A(n9545), .ZN(n9535) );
  INV_X1 U11330 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9532) );
  NAND2_X1 U11331 ( .A1(n9533), .A2(n9532), .ZN(n9534) );
  NAND2_X1 U11332 ( .A1(n9535), .A2(n9534), .ZN(n15563) );
  OR2_X1 U11333 ( .A1(n15563), .A2(n7814), .ZN(n9541) );
  INV_X1 U11334 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9538) );
  NAND2_X1 U11335 ( .A1(n9254), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n9537) );
  NAND2_X1 U11336 ( .A1(n7818), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9536) );
  OAI211_X1 U11337 ( .C1(n9634), .C2(n9538), .A(n9537), .B(n9536), .ZN(n9539)
         );
  INV_X1 U11338 ( .A(n9539), .ZN(n9540) );
  NAND2_X1 U11339 ( .A1(n9541), .A2(n9540), .ZN(n15309) );
  XNOR2_X1 U11340 ( .A(n15699), .B(n15309), .ZN(n15559) );
  INV_X1 U11341 ( .A(n15309), .ZN(n14934) );
  NAND2_X1 U11342 ( .A1(n11677), .A2(n15206), .ZN(n9544) );
  NAND2_X1 U11343 ( .A1(n7460), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9543) );
  NOR2_X1 U11344 ( .A1(n9545), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9546) );
  OR2_X1 U11345 ( .A1(n9547), .A2(n9546), .ZN(n15547) );
  INV_X1 U11346 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9550) );
  NAND2_X1 U11347 ( .A1(n9254), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9549) );
  NAND2_X1 U11348 ( .A1(n7818), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9548) );
  OAI211_X1 U11349 ( .C1(n9634), .C2(n9550), .A(n9549), .B(n9548), .ZN(n9551)
         );
  INV_X1 U11350 ( .A(n9551), .ZN(n9552) );
  OAI21_X1 U11351 ( .B1(n15547), .B2(n7814), .A(n9552), .ZN(n15308) );
  XNOR2_X1 U11352 ( .A(n15694), .B(n15308), .ZN(n15252) );
  INV_X1 U11353 ( .A(n15308), .ZN(n9553) );
  NAND2_X1 U11354 ( .A1(n15540), .A2(n9554), .ZN(n15527) );
  NAND2_X1 U11355 ( .A1(n15688), .A2(n15146), .ZN(n9670) );
  OR2_X1 U11356 ( .A1(n15688), .A2(n15146), .ZN(n9555) );
  NAND2_X1 U11357 ( .A1(n9670), .A2(n9555), .ZN(n15524) );
  NAND2_X1 U11358 ( .A1(n12149), .A2(n15206), .ZN(n9557) );
  NAND2_X1 U11359 ( .A1(n7460), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9556) );
  NAND2_X1 U11360 ( .A1(n7818), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9565) );
  INV_X1 U11361 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9558) );
  OR2_X1 U11362 ( .A1(n7778), .A2(n9558), .ZN(n9564) );
  OAI21_X1 U11363 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n9560), .A(n9559), .ZN(
        n15513) );
  OR2_X1 U11364 ( .A1(n7814), .A2(n15513), .ZN(n9563) );
  INV_X1 U11365 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9561) );
  OR2_X1 U11366 ( .A1(n9634), .A2(n9561), .ZN(n9562) );
  NAND4_X1 U11367 ( .A1(n9565), .A2(n9564), .A3(n9563), .A4(n9562), .ZN(n15306) );
  INV_X1 U11368 ( .A(n15306), .ZN(n9566) );
  XNOR2_X1 U11369 ( .A(n15681), .B(n9566), .ZN(n15255) );
  INV_X1 U11370 ( .A(n15681), .ZN(n9567) );
  INV_X1 U11371 ( .A(n15305), .ZN(n14953) );
  INV_X1 U11372 ( .A(n15304), .ZN(n15018) );
  XNOR2_X1 U11373 ( .A(n15668), .B(n15018), .ZN(n15483) );
  INV_X1 U11374 ( .A(n15483), .ZN(n15478) );
  NAND2_X1 U11375 ( .A1(n15479), .A2(n15478), .ZN(n15477) );
  NAND2_X1 U11376 ( .A1(n7460), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9569) );
  NAND2_X1 U11377 ( .A1(n9607), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9578) );
  INV_X1 U11378 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9571) );
  OR2_X1 U11379 ( .A1(n9477), .A2(n9571), .ZN(n9577) );
  OAI21_X1 U11380 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n9573), .A(n9584), .ZN(
        n15467) );
  OR2_X1 U11381 ( .A1(n7814), .A2(n15467), .ZN(n9576) );
  INV_X1 U11382 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9574) );
  OR2_X1 U11383 ( .A1(n7778), .A2(n9574), .ZN(n9575) );
  NAND4_X1 U11384 ( .A1(n9578), .A2(n9577), .A3(n9576), .A4(n9575), .ZN(n15303) );
  INV_X1 U11385 ( .A(n15303), .ZN(n14952) );
  NAND2_X1 U11386 ( .A1(n7459), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9579) );
  NAND2_X1 U11387 ( .A1(n7818), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9590) );
  INV_X1 U11388 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9581) );
  OR2_X1 U11389 ( .A1(n7778), .A2(n9581), .ZN(n9589) );
  INV_X1 U11390 ( .A(n9584), .ZN(n9582) );
  NAND2_X1 U11391 ( .A1(n9582), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9596) );
  INV_X1 U11392 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9583) );
  NAND2_X1 U11393 ( .A1(n9584), .A2(n9583), .ZN(n9585) );
  NAND2_X1 U11394 ( .A1(n9596), .A2(n9585), .ZN(n15455) );
  INV_X1 U11395 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9586) );
  OR2_X1 U11396 ( .A1(n9634), .A2(n9586), .ZN(n9587) );
  INV_X1 U11397 ( .A(n15659), .ZN(n15460) );
  NAND2_X1 U11398 ( .A1(n7460), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9591) );
  NAND2_X1 U11399 ( .A1(n9607), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9602) );
  INV_X1 U11400 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9593) );
  OR2_X1 U11401 ( .A1(n9477), .A2(n9593), .ZN(n9601) );
  INV_X1 U11402 ( .A(n9596), .ZN(n9594) );
  NAND2_X1 U11403 ( .A1(n9594), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n12779) );
  INV_X1 U11404 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9595) );
  NAND2_X1 U11405 ( .A1(n9596), .A2(n9595), .ZN(n9597) );
  NAND2_X1 U11406 ( .A1(n12779), .A2(n9597), .ZN(n15440) );
  INV_X1 U11407 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9598) );
  OR2_X1 U11408 ( .A1(n7778), .A2(n9598), .ZN(n9599) );
  NAND4_X1 U11409 ( .A1(n9602), .A2(n9601), .A3(n9600), .A4(n9599), .ZN(n15301) );
  INV_X1 U11410 ( .A(n15301), .ZN(n9604) );
  NAND2_X1 U11411 ( .A1(n12790), .A2(n15206), .ZN(n9606) );
  NAND2_X1 U11412 ( .A1(n7459), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9605) );
  NAND2_X1 U11413 ( .A1(n9607), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9613) );
  INV_X1 U11414 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9608) );
  OR2_X1 U11415 ( .A1(n9477), .A2(n9608), .ZN(n9612) );
  OR2_X1 U11416 ( .A1(n7814), .A2(n12779), .ZN(n9611) );
  INV_X1 U11417 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9609) );
  OR2_X1 U11418 ( .A1(n7778), .A2(n9609), .ZN(n9610) );
  INV_X1 U11419 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9615) );
  NAND2_X1 U11420 ( .A1(n9618), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9617) );
  NAND2_X1 U11421 ( .A1(n15783), .A2(n11573), .ZN(n15034) );
  NAND2_X1 U11422 ( .A1(n9620), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9621) );
  XNOR2_X1 U11423 ( .A(n9621), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9714) );
  NAND2_X1 U11424 ( .A1(n9622), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9623) );
  INV_X1 U11425 ( .A(n15212), .ZN(n15217) );
  NAND2_X1 U11426 ( .A1(n9714), .A2(n15217), .ZN(n9624) );
  NAND2_X1 U11427 ( .A1(n15034), .A2(n9624), .ZN(n16536) );
  NAND2_X1 U11428 ( .A1(n12788), .A2(n16536), .ZN(n9683) );
  INV_X1 U11429 ( .A(n15105), .ZN(n12294) );
  NAND2_X1 U11430 ( .A1(n16339), .A2(n16327), .ZN(n16329) );
  OR2_X1 U11431 ( .A1(n16329), .A2(n7812), .ZN(n12107) );
  INV_X1 U11432 ( .A(n15074), .ZN(n16493) );
  INV_X1 U11433 ( .A(n15078), .ZN(n16511) );
  NAND2_X1 U11434 ( .A1(n12294), .A2(n12291), .ZN(n12494) );
  INV_X1 U11435 ( .A(n15703), .ZN(n15579) );
  NAND2_X1 U11436 ( .A1(n15572), .A2(n15579), .ZN(n15573) );
  INV_X1 U11437 ( .A(n15439), .ZN(n9627) );
  AOI211_X1 U11438 ( .C1(n15193), .C2(n9627), .A(n16437), .B(n15430), .ZN(
        n12778) );
  AND2_X1 U11439 ( .A1(n15212), .A2(n15417), .ZN(n9711) );
  INV_X1 U11440 ( .A(n9711), .ZN(n9628) );
  INV_X1 U11441 ( .A(n15033), .ZN(n10579) );
  INV_X1 U11442 ( .A(n15772), .ZN(n15347) );
  NAND2_X1 U11443 ( .A1(n10579), .A2(n15347), .ZN(n15293) );
  NAND2_X1 U11444 ( .A1(n15006), .A2(n15301), .ZN(n12782) );
  NAND2_X1 U11445 ( .A1(n10579), .A2(n15772), .ZN(n15016) );
  INV_X1 U11446 ( .A(P1_B_REG_SCAN_IN), .ZN(n9629) );
  NOR2_X1 U11447 ( .A1(n15885), .A2(n9629), .ZN(n9630) );
  NOR2_X1 U11448 ( .A1(n15016), .A2(n9630), .ZN(n15425) );
  INV_X1 U11449 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9633) );
  NAND2_X1 U11450 ( .A1(n7818), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9632) );
  NAND2_X1 U11451 ( .A1(n9254), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9631) );
  OAI211_X1 U11452 ( .C1(n9634), .C2(n9633), .A(n9632), .B(n9631), .ZN(n15299)
         );
  NAND2_X1 U11453 ( .A1(n15425), .A2(n15299), .ZN(n12780) );
  OAI211_X1 U11454 ( .C1(n15191), .C2(n16476), .A(n12782), .B(n12780), .ZN(
        n9635) );
  NAND2_X1 U11455 ( .A1(n15045), .A2(n15044), .ZN(n15233) );
  INV_X1 U11456 ( .A(n16327), .ZN(n11574) );
  NAND2_X1 U11457 ( .A1(n15327), .A2(n11574), .ZN(n16326) );
  NAND2_X1 U11458 ( .A1(n15233), .A2(n16326), .ZN(n9638) );
  NAND2_X1 U11459 ( .A1(n9269), .A2(n16339), .ZN(n9637) );
  NAND2_X1 U11460 ( .A1(n9638), .A2(n9637), .ZN(n11996) );
  NAND2_X1 U11461 ( .A1(n11996), .A2(n15234), .ZN(n9641) );
  INV_X1 U11462 ( .A(n9639), .ZN(n11210) );
  NAND2_X1 U11463 ( .A1(n11210), .A2(n16374), .ZN(n9640) );
  INV_X1 U11464 ( .A(n15235), .ZN(n9642) );
  NAND2_X1 U11465 ( .A1(n12106), .A2(n9642), .ZN(n9644) );
  NAND2_X1 U11466 ( .A1(n9644), .A2(n9643), .ZN(n12056) );
  INV_X1 U11467 ( .A(n15236), .ZN(n9645) );
  NAND2_X1 U11468 ( .A1(n12056), .A2(n9645), .ZN(n9647) );
  NAND2_X1 U11469 ( .A1(n15055), .A2(n15056), .ZN(n9646) );
  NAND2_X1 U11470 ( .A1(n9647), .A2(n9646), .ZN(n16433) );
  NAND2_X1 U11471 ( .A1(n16433), .A2(n16434), .ZN(n9649) );
  OR2_X1 U11472 ( .A1(n16448), .A2(n15324), .ZN(n9648) );
  XNOR2_X1 U11473 ( .A(n15074), .B(n11768), .ZN(n16477) );
  NAND2_X1 U11474 ( .A1(n15078), .A2(n15321), .ZN(n9652) );
  NAND2_X1 U11475 ( .A1(n11765), .A2(n9652), .ZN(n12000) );
  INV_X1 U11476 ( .A(n12000), .ZN(n9654) );
  XNOR2_X1 U11477 ( .A(n16531), .B(n15320), .ZN(n15241) );
  OR2_X1 U11478 ( .A1(n16531), .A2(n15320), .ZN(n9655) );
  OR2_X1 U11479 ( .A1(n15090), .A2(n15319), .ZN(n9656) );
  XNOR2_X1 U11480 ( .A(n16572), .B(n15318), .ZN(n15243) );
  NAND2_X1 U11481 ( .A1(n16572), .A2(n15318), .ZN(n9657) );
  OR2_X1 U11482 ( .A1(n15101), .A2(n15317), .ZN(n9658) );
  NAND2_X1 U11483 ( .A1(n12289), .A2(n15247), .ZN(n12288) );
  OR2_X1 U11484 ( .A1(n15105), .A2(n15316), .ZN(n9659) );
  INV_X1 U11485 ( .A(n15248), .ZN(n12491) );
  NAND2_X1 U11486 ( .A1(n16611), .A2(n15315), .ZN(n9660) );
  INV_X1 U11487 ( .A(n15625), .ZN(n15629) );
  OR2_X1 U11488 ( .A1(n15725), .A2(n15313), .ZN(n9661) );
  OR2_X1 U11489 ( .A1(n15710), .A2(n15311), .ZN(n9664) );
  OR2_X1 U11490 ( .A1(n15703), .A2(n15310), .ZN(n9665) );
  INV_X1 U11491 ( .A(n9665), .ZN(n9666) );
  NAND2_X1 U11492 ( .A1(n15699), .A2(n15309), .ZN(n9668) );
  OR2_X1 U11493 ( .A1(n15694), .A2(n15308), .ZN(n9669) );
  NAND2_X1 U11494 ( .A1(n15681), .A2(n15306), .ZN(n9671) );
  OR2_X1 U11495 ( .A1(n15675), .A2(n15305), .ZN(n9672) );
  NAND2_X1 U11496 ( .A1(n15668), .A2(n15304), .ZN(n9673) );
  NAND2_X1 U11497 ( .A1(n15664), .A2(n15303), .ZN(n9674) );
  NAND2_X1 U11498 ( .A1(n15468), .A2(n9674), .ZN(n15450) );
  NOR2_X1 U11499 ( .A1(n9675), .A2(n8507), .ZN(n15446) );
  NAND2_X1 U11500 ( .A1(n15783), .A2(n15417), .ZN(n9677) );
  AND2_X2 U11501 ( .A1(n9677), .A2(n11575), .ZN(n14827) );
  AND2_X1 U11502 ( .A1(n15783), .A2(n15038), .ZN(n9678) );
  NOR2_X1 U11503 ( .A1(n14827), .A2(n9678), .ZN(n12070) );
  NAND2_X1 U11504 ( .A1(n12070), .A2(n15417), .ZN(n16370) );
  NAND2_X1 U11505 ( .A1(n15212), .A2(n11573), .ZN(n9679) );
  INV_X1 U11506 ( .A(n16486), .ZN(n16468) );
  NAND2_X1 U11507 ( .A1(n9680), .A2(n16443), .ZN(n9681) );
  INV_X1 U11508 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9684) );
  NAND2_X1 U11509 ( .A1(n9705), .A2(P1_B_REG_SCAN_IN), .ZN(n9687) );
  MUX2_X1 U11510 ( .A(n9687), .B(P1_B_REG_SCAN_IN), .S(n9704), .Z(n9691) );
  NAND2_X1 U11511 ( .A1(n9688), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9689) );
  MUX2_X1 U11512 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9689), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n9690) );
  AND2_X1 U11513 ( .A1(n9205), .A2(n9690), .ZN(n9716) );
  OR2_X1 U11514 ( .A1(n10468), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9692) );
  INV_X1 U11515 ( .A(n9716), .ZN(n15781) );
  NAND2_X1 U11516 ( .A1(n9705), .A2(n15781), .ZN(n10470) );
  AND2_X1 U11517 ( .A1(n9692), .A2(n10470), .ZN(n11174) );
  NOR4_X1 U11518 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n9696) );
  NOR4_X1 U11519 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n9695) );
  NOR4_X1 U11520 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n9694) );
  NOR4_X1 U11521 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n9693) );
  NAND4_X1 U11522 ( .A1(n9696), .A2(n9695), .A3(n9694), .A4(n9693), .ZN(n9702)
         );
  NOR2_X1 U11523 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n9700) );
  NOR4_X1 U11524 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n9699) );
  NOR4_X1 U11525 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9698) );
  NOR4_X1 U11526 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9697) );
  NAND4_X1 U11527 ( .A1(n9700), .A2(n9699), .A3(n9698), .A4(n9697), .ZN(n9701)
         );
  NOR2_X1 U11528 ( .A1(n9702), .A2(n9701), .ZN(n9703) );
  OR2_X1 U11529 ( .A1(n10468), .A2(n9703), .ZN(n11173) );
  NAND2_X1 U11530 ( .A1(n7489), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9708) );
  MUX2_X1 U11531 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9708), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n9710) );
  NAND2_X1 U11532 ( .A1(n9710), .A2(n9709), .ZN(n10578) );
  OAI21_X1 U11533 ( .B1(n15033), .B2(n9711), .A(n10578), .ZN(n9712) );
  INV_X1 U11534 ( .A(n9712), .ZN(n9713) );
  NAND2_X1 U11535 ( .A1(n11177), .A2(n9713), .ZN(n11280) );
  INV_X1 U11536 ( .A(n15294), .ZN(n11175) );
  INV_X1 U11537 ( .A(n9714), .ZN(n15218) );
  NAND2_X1 U11538 ( .A1(n16486), .A2(n15218), .ZN(n11570) );
  NAND3_X1 U11539 ( .A1(n11173), .A2(n11175), .A3(n11570), .ZN(n9715) );
  OR2_X1 U11540 ( .A1(n10468), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9717) );
  OR2_X1 U11541 ( .A1(n9704), .A2(n9716), .ZN(n15759) );
  NAND2_X1 U11542 ( .A1(n9722), .A2(n7435), .ZN(n9719) );
  NAND2_X1 U11543 ( .A1(n16579), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9718) );
  NAND2_X1 U11544 ( .A1(n9719), .A2(n9718), .ZN(P1_U3557) );
  INV_X1 U11545 ( .A(n11567), .ZN(n9720) );
  NAND2_X1 U11546 ( .A1(n16580), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U11547 ( .A1(n9724), .A2(n9723), .ZN(P1_U3525) );
  INV_X1 U11548 ( .A(n10385), .ZN(n9725) );
  INV_X2 U11549 ( .A(n16561), .ZN(n11936) );
  NAND2_X1 U11550 ( .A1(n11936), .A2(n16382), .ZN(n14768) );
  INV_X1 U11551 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9728) );
  INV_X1 U11552 ( .A(n9729), .ZN(n9730) );
  NAND2_X1 U11553 ( .A1(n9731), .A2(n9730), .ZN(P2_U3496) );
  INV_X1 U11554 ( .A(n9732), .ZN(n9737) );
  INV_X1 U11555 ( .A(n9733), .ZN(n9735) );
  INV_X1 U11556 ( .A(n14312), .ZN(n9734) );
  OAI21_X1 U11557 ( .B1(n9735), .B2(n9734), .A(n14606), .ZN(n9736) );
  AOI22_X1 U11558 ( .A1(n14340), .A2(n14589), .B1(n14588), .B2(n14342), .ZN(
        n13914) );
  OAI21_X1 U11559 ( .B1(n9737), .B2(n9736), .A(n13914), .ZN(n14458) );
  INV_X1 U11560 ( .A(n14466), .ZN(n9740) );
  INV_X1 U11561 ( .A(n14193), .ZN(n14648) );
  OAI211_X1 U11562 ( .C1(n9740), .C2(n14648), .A(n7507), .B(n14430), .ZN(n9741) );
  NOR2_X1 U11563 ( .A1(n11936), .A2(n9742), .ZN(n9743) );
  INV_X1 U11564 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n10342) );
  NOR2_X1 U11565 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), 
        .ZN(n9748) );
  NOR2_X1 U11566 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), 
        .ZN(n9747) );
  NOR2_X1 U11567 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n9753) );
  INV_X1 U11568 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n9757) );
  XNOR2_X2 U11569 ( .A(n9758), .B(n9757), .ZN(n13854) );
  INV_X1 U11570 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n16321) );
  NAND2_X1 U11571 ( .A1(n9813), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n9759) );
  INV_X1 U11572 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10992) );
  INV_X1 U11573 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10991) );
  XNOR2_X1 U11574 ( .A(n9785), .B(n9786), .ZN(n9763) );
  NAND2_X1 U11575 ( .A1(n9764), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9766) );
  INV_X1 U11576 ( .A(n9767), .ZN(n10310) );
  MUX2_X1 U11577 ( .A(n13855), .B(n13856), .S(n9860), .Z(n16316) );
  INV_X1 U11578 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10818) );
  OR2_X1 U11579 ( .A1(n9815), .A2(n10818), .ZN(n9773) );
  NAND2_X1 U11580 ( .A1(n9813), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9772) );
  INV_X1 U11581 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10996) );
  INV_X1 U11582 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n13005) );
  MUX2_X1 U11583 ( .A(n13005), .B(n10420), .S(n9860), .Z(n9778) );
  NAND2_X2 U11584 ( .A1(n9860), .A2(n8156), .ZN(n9800) );
  INV_X1 U11585 ( .A(n9785), .ZN(n9776) );
  NAND2_X1 U11586 ( .A1(n7746), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9775) );
  AND2_X1 U11587 ( .A1(n9776), .A2(n9775), .ZN(n10422) );
  OR2_X1 U11588 ( .A1(n9800), .A2(n10422), .ZN(n9777) );
  INV_X1 U11589 ( .A(n10813), .ZN(n11626) );
  NAND2_X1 U11590 ( .A1(n9780), .A2(n8116), .ZN(n16346) );
  NAND2_X1 U11591 ( .A1(n16309), .A2(n16346), .ZN(n9795) );
  INV_X1 U11592 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10999) );
  INV_X1 U11593 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10998) );
  OR2_X1 U11594 ( .A1(n9814), .A2(n10998), .ZN(n9783) );
  NAND2_X1 U11595 ( .A1(n9813), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9782) );
  INV_X1 U11596 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n16361) );
  OR2_X1 U11597 ( .A1(n9815), .A2(n16361), .ZN(n9781) );
  INV_X2 U11598 ( .A(n9794), .ZN(n16314) );
  NAND2_X1 U11599 ( .A1(n10412), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9787) );
  NAND2_X1 U11600 ( .A1(n10416), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n9788) );
  XNOR2_X1 U11601 ( .A(n9797), .B(n9796), .ZN(n10433) );
  NAND2_X1 U11602 ( .A1(n10088), .A2(n11026), .ZN(n9791) );
  NAND2_X1 U11603 ( .A1(n9795), .A2(n10277), .ZN(n11732) );
  OR2_X1 U11604 ( .A1(n12569), .A2(SI_3_), .ZN(n9805) );
  NAND2_X1 U11605 ( .A1(n10406), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n9799) );
  XNOR2_X1 U11606 ( .A(n9823), .B(n9822), .ZN(n10425) );
  OR2_X1 U11607 ( .A1(n9800), .A2(n10425), .ZN(n9804) );
  NAND2_X1 U11608 ( .A1(n9801), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9802) );
  XNOR2_X1 U11609 ( .A(n9802), .B(n9746), .ZN(n11028) );
  NAND2_X1 U11610 ( .A1(n10088), .A2(n11028), .ZN(n9803) );
  NAND2_X1 U11611 ( .A1(n9813), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9809) );
  INV_X1 U11612 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11003) );
  OR2_X1 U11613 ( .A1(n9814), .A2(n11003), .ZN(n9808) );
  INV_X1 U11614 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n16114) );
  OR2_X1 U11615 ( .A1(n9817), .A2(n16114), .ZN(n9807) );
  OR2_X1 U11616 ( .A1(n9815), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n9806) );
  INV_X1 U11617 ( .A(n11081), .ZN(n16390) );
  NAND2_X1 U11618 ( .A1(n9810), .A2(n16390), .ZN(n12607) );
  AND2_X1 U11619 ( .A1(n16314), .A2(n16363), .ZN(n11733) );
  NAND2_X1 U11620 ( .A1(n11732), .A2(n9811), .ZN(n11736) );
  NAND2_X1 U11621 ( .A1(n9810), .A2(n11081), .ZN(n9812) );
  NAND2_X1 U11622 ( .A1(n11736), .A2(n9812), .ZN(n11592) );
  NAND2_X1 U11623 ( .A1(n9813), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9821) );
  INV_X1 U11624 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11008) );
  OR2_X1 U11625 ( .A1(n9814), .A2(n11008), .ZN(n9820) );
  NAND2_X1 U11626 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9816) );
  AND2_X1 U11627 ( .A1(n9837), .A2(n9816), .ZN(n11301) );
  OR2_X1 U11628 ( .A1(n9815), .A2(n11301), .ZN(n9819) );
  INV_X1 U11629 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11595) );
  OR2_X1 U11630 ( .A1(n9817), .A2(n11595), .ZN(n9818) );
  OR2_X1 U11631 ( .A1(n12569), .A2(SI_4_), .ZN(n9832) );
  XNOR2_X1 U11632 ( .A(n9846), .B(n9844), .ZN(n10429) );
  OR2_X1 U11633 ( .A1(n9800), .A2(n10429), .ZN(n9831) );
  INV_X1 U11634 ( .A(n9825), .ZN(n9829) );
  NAND2_X1 U11635 ( .A1(n9826), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9827) );
  MUX2_X1 U11636 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9827), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n9828) );
  NAND2_X1 U11637 ( .A1(n9829), .A2(n9828), .ZN(n11113) );
  NAND2_X1 U11638 ( .A1(n10088), .A2(n11113), .ZN(n9830) );
  NAND2_X1 U11639 ( .A1(n11738), .A2(n11597), .ZN(n12612) );
  INV_X1 U11640 ( .A(n11738), .ZN(n12996) );
  INV_X1 U11641 ( .A(n11597), .ZN(n16413) );
  NAND2_X1 U11642 ( .A1(n12996), .A2(n16413), .ZN(n12613) );
  INV_X1 U11643 ( .A(n12610), .ZN(n12738) );
  NAND2_X1 U11644 ( .A1(n11592), .A2(n12738), .ZN(n9834) );
  NAND2_X1 U11645 ( .A1(n12996), .A2(n11597), .ZN(n9833) );
  NAND2_X1 U11646 ( .A1(n9834), .A2(n9833), .ZN(n11698) );
  NAND2_X1 U11647 ( .A1(n9813), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9843) );
  INV_X1 U11648 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n9835) );
  OR2_X1 U11649 ( .A1(n9814), .A2(n9835), .ZN(n9842) );
  NAND2_X1 U11650 ( .A1(n9837), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n9838) );
  AND2_X1 U11651 ( .A1(n9854), .A2(n9838), .ZN(n11965) );
  OR2_X1 U11652 ( .A1(n9815), .A2(n11965), .ZN(n9841) );
  INV_X1 U11653 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n9839) );
  OR2_X1 U11654 ( .A1(n9817), .A2(n9839), .ZN(n9840) );
  OR2_X1 U11655 ( .A1(n12569), .A2(SI_5_), .ZN(n9853) );
  INV_X1 U11656 ( .A(n9844), .ZN(n9845) );
  XNOR2_X1 U11657 ( .A(n9865), .B(n9864), .ZN(n10431) );
  OR2_X1 U11658 ( .A1(n9800), .A2(n10431), .ZN(n9852) );
  OR2_X1 U11659 ( .A1(n9825), .A2(n13843), .ZN(n9850) );
  XNOR2_X1 U11660 ( .A(n9850), .B(n9849), .ZN(n11246) );
  NAND2_X1 U11661 ( .A1(n10088), .A2(n11246), .ZN(n9851) );
  NAND2_X1 U11662 ( .A1(n11926), .A2(n11703), .ZN(n12616) );
  INV_X1 U11663 ( .A(n11926), .ZN(n10632) );
  INV_X1 U11664 ( .A(n11703), .ZN(n11966) );
  NAND2_X1 U11665 ( .A1(n10632), .A2(n11966), .ZN(n12617) );
  NAND2_X1 U11666 ( .A1(n9813), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9859) );
  NAND2_X1 U11667 ( .A1(n9854), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9855) );
  AND2_X1 U11668 ( .A1(n9875), .A2(n9855), .ZN(n11920) );
  OR2_X1 U11669 ( .A1(n9815), .A2(n11920), .ZN(n9858) );
  INV_X1 U11670 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n16131) );
  OR2_X1 U11671 ( .A1(n9817), .A2(n16131), .ZN(n9857) );
  NAND2_X1 U11672 ( .A1(n11433), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9856) );
  NAND4_X1 U11673 ( .A1(n9859), .A2(n9858), .A3(n9857), .A4(n9856), .ZN(n12995) );
  OR2_X1 U11674 ( .A1(n9861), .A2(n13843), .ZN(n9862) );
  XNOR2_X1 U11675 ( .A(n9862), .B(n9884), .ZN(n16143) );
  NAND2_X1 U11676 ( .A1(n10450), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9866) );
  OR2_X1 U11677 ( .A1(n9868), .A2(n9867), .ZN(n9869) );
  AND2_X1 U11678 ( .A1(n9883), .A2(n9869), .ZN(n10440) );
  OR2_X1 U11679 ( .A1(n9800), .A2(n10440), .ZN(n9871) );
  INV_X1 U11680 ( .A(SI_6_), .ZN(n10439) );
  OR2_X1 U11681 ( .A1(n12569), .A2(n10439), .ZN(n9870) );
  OAI211_X1 U11682 ( .C1(n9860), .C2(n16143), .A(n9871), .B(n9870), .ZN(n12620) );
  XNOR2_X1 U11683 ( .A(n12995), .B(n12620), .ZN(n12745) );
  AND2_X1 U11684 ( .A1(n11926), .A2(n11966), .ZN(n11921) );
  NOR2_X1 U11685 ( .A1(n12745), .A2(n11921), .ZN(n9872) );
  NAND2_X1 U11686 ( .A1(n12995), .A2(n12620), .ZN(n9873) );
  NAND2_X1 U11687 ( .A1(n9813), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9881) );
  INV_X1 U11688 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11851) );
  OR2_X1 U11689 ( .A1(n9817), .A2(n11851), .ZN(n9880) );
  NAND2_X1 U11690 ( .A1(n9875), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9876) );
  AND2_X1 U11691 ( .A1(n9890), .A2(n9876), .ZN(n11689) );
  OR2_X1 U11692 ( .A1(n9815), .A2(n11689), .ZN(n9879) );
  INV_X1 U11693 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n9877) );
  OR2_X1 U11694 ( .A1(n9814), .A2(n9877), .ZN(n9878) );
  OR2_X1 U11695 ( .A1(n12569), .A2(SI_7_), .ZN(n9889) );
  XNOR2_X1 U11696 ( .A(n9904), .B(n9901), .ZN(n10427) );
  OR2_X1 U11697 ( .A1(n9800), .A2(n10427), .ZN(n9888) );
  NAND2_X1 U11698 ( .A1(n9861), .A2(n9884), .ZN(n9896) );
  NAND2_X1 U11699 ( .A1(n9896), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9886) );
  XNOR2_X1 U11700 ( .A(n9886), .B(n9885), .ZN(n11526) );
  NAND2_X1 U11701 ( .A1(n10088), .A2(n11526), .ZN(n9887) );
  NAND2_X1 U11702 ( .A1(n12022), .A2(n11859), .ZN(n12626) );
  INV_X1 U11703 ( .A(n12022), .ZN(n12994) );
  NAND2_X1 U11704 ( .A1(n12994), .A2(n11862), .ZN(n12627) );
  INV_X1 U11705 ( .A(n12624), .ZN(n12737) );
  NAND2_X1 U11706 ( .A1(n9813), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9895) );
  INV_X1 U11707 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11537) );
  OR2_X1 U11708 ( .A1(n9814), .A2(n11537), .ZN(n9894) );
  NAND2_X1 U11709 ( .A1(n9890), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9891) );
  AND2_X1 U11710 ( .A1(n9913), .A2(n9891), .ZN(n12027) );
  OR2_X1 U11711 ( .A1(n9815), .A2(n12027), .ZN(n9893) );
  INV_X1 U11712 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11529) );
  OR2_X1 U11713 ( .A1(n9817), .A2(n11529), .ZN(n9892) );
  NAND2_X1 U11714 ( .A1(n9899), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9898) );
  MUX2_X1 U11715 ( .A(n9898), .B(P3_IR_REG_31__SCAN_IN), .S(n9897), .Z(n9900)
         );
  NAND2_X1 U11716 ( .A1(n9900), .A2(n9922), .ZN(n11667) );
  NAND2_X1 U11717 ( .A1(n10456), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9902) );
  NAND2_X1 U11718 ( .A1(n10463), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9905) );
  NAND2_X1 U11719 ( .A1(n9925), .A2(n9905), .ZN(n9906) );
  NAND2_X1 U11720 ( .A1(n9907), .A2(n9906), .ZN(n9908) );
  AND2_X1 U11721 ( .A1(n9926), .A2(n9908), .ZN(n10438) );
  OR2_X1 U11722 ( .A1(n9800), .A2(n10438), .ZN(n9910) );
  INV_X1 U11723 ( .A(SI_8_), .ZN(n10437) );
  OR2_X1 U11724 ( .A1(n12569), .A2(n10437), .ZN(n9909) );
  OAI211_X1 U11725 ( .C1(n9860), .C2(n11667), .A(n9910), .B(n9909), .ZN(n16501) );
  NAND2_X1 U11726 ( .A1(n12140), .A2(n16501), .ZN(n12631) );
  INV_X1 U11727 ( .A(n12140), .ZN(n12993) );
  INV_X1 U11728 ( .A(n16501), .ZN(n11871) );
  NAND2_X1 U11729 ( .A1(n12993), .A2(n11871), .ZN(n12632) );
  NAND2_X1 U11730 ( .A1(n12140), .A2(n11871), .ZN(n9911) );
  NAND2_X1 U11731 ( .A1(n11866), .A2(n9911), .ZN(n12125) );
  NAND2_X1 U11732 ( .A1(n11433), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9919) );
  NAND2_X1 U11733 ( .A1(n9913), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n9914) );
  AND2_X1 U11734 ( .A1(n9932), .A2(n9914), .ZN(n12147) );
  OR2_X1 U11735 ( .A1(n9815), .A2(n12147), .ZN(n9918) );
  INV_X1 U11736 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n9915) );
  OR2_X1 U11737 ( .A1(n9817), .A2(n9915), .ZN(n9917) );
  NAND2_X1 U11738 ( .A1(n9813), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9916) );
  NAND2_X1 U11739 ( .A1(n9922), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9921) );
  MUX2_X1 U11740 ( .A(n9921), .B(P3_IR_REG_31__SCAN_IN), .S(n9920), .Z(n9924)
         );
  INV_X1 U11741 ( .A(n9958), .ZN(n9923) );
  NAND2_X1 U11742 ( .A1(n9924), .A2(n9923), .ZN(n11831) );
  INV_X1 U11743 ( .A(n11831), .ZN(n11817) );
  OR2_X1 U11744 ( .A1(n12569), .A2(SI_9_), .ZN(n9928) );
  XNOR2_X1 U11745 ( .A(n9941), .B(n9939), .ZN(n10441) );
  OR2_X1 U11746 ( .A1(n9800), .A2(n10441), .ZN(n9927) );
  OAI211_X1 U11747 ( .C1(n11817), .C2(n9860), .A(n9928), .B(n9927), .ZN(n16523) );
  INV_X1 U11748 ( .A(n16523), .ZN(n12144) );
  NAND2_X1 U11749 ( .A1(n12992), .A2(n12144), .ZN(n9929) );
  NAND2_X1 U11750 ( .A1(n12125), .A2(n9929), .ZN(n9931) );
  NAND2_X1 U11751 ( .A1(n12133), .A2(n16523), .ZN(n9930) );
  NAND2_X1 U11752 ( .A1(n11433), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9937) );
  NAND2_X1 U11753 ( .A1(n9813), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9936) );
  NAND2_X1 U11754 ( .A1(n9932), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9933) );
  AND2_X1 U11755 ( .A1(n9945), .A2(n9933), .ZN(n12206) );
  OR2_X1 U11756 ( .A1(n9815), .A2(n12206), .ZN(n9935) );
  NAND2_X1 U11757 ( .A1(n9770), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n9934) );
  OR2_X1 U11758 ( .A1(n9958), .A2(n13843), .ZN(n9938) );
  XNOR2_X1 U11759 ( .A(n9938), .B(P3_IR_REG_10__SCAN_IN), .ZN(n11834) );
  OR2_X1 U11760 ( .A1(n12569), .A2(SI_10_), .ZN(n9943) );
  XNOR2_X1 U11761 ( .A(n9954), .B(P1_DATAO_REG_10__SCAN_IN), .ZN(n9951) );
  XNOR2_X1 U11762 ( .A(n9953), .B(n9951), .ZN(n10435) );
  OR2_X1 U11763 ( .A1(n9800), .A2(n10435), .ZN(n9942) );
  OAI211_X1 U11764 ( .C1(n11834), .C2(n9860), .A(n9943), .B(n9942), .ZN(n12639) );
  XNOR2_X1 U11765 ( .A(n12640), .B(n12639), .ZN(n12194) );
  NAND2_X1 U11766 ( .A1(n9813), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9950) );
  INV_X1 U11767 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n9944) );
  OR2_X1 U11768 ( .A1(n9814), .A2(n9944), .ZN(n9949) );
  NAND2_X1 U11769 ( .A1(n9945), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9946) );
  AND2_X1 U11770 ( .A1(n9967), .A2(n9946), .ZN(n12270) );
  OR2_X1 U11771 ( .A1(n9815), .A2(n12270), .ZN(n9948) );
  INV_X1 U11772 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12231) );
  OR2_X1 U11773 ( .A1(n9817), .A2(n12231), .ZN(n9947) );
  INV_X1 U11774 ( .A(n9951), .ZN(n9952) );
  NAND2_X1 U11775 ( .A1(n9954), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9955) );
  NAND2_X1 U11776 ( .A1(n10545), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9975) );
  NAND2_X1 U11777 ( .A1(n10543), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9956) );
  NAND2_X1 U11778 ( .A1(n9975), .A2(n9956), .ZN(n9973) );
  XNOR2_X1 U11779 ( .A(n9974), .B(n9973), .ZN(n10452) );
  OR2_X1 U11780 ( .A1(n9800), .A2(n10452), .ZN(n9962) );
  OR2_X1 U11781 ( .A1(n12569), .A2(SI_11_), .ZN(n9961) );
  OR2_X1 U11782 ( .A1(n9977), .A2(n13843), .ZN(n9959) );
  INV_X1 U11783 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9976) );
  XNOR2_X1 U11784 ( .A(n9959), .B(n9976), .ZN(n13047) );
  NAND2_X1 U11785 ( .A1(n10088), .A2(n13047), .ZN(n9960) );
  NAND2_X1 U11786 ( .A1(n12267), .A2(n12272), .ZN(n12651) );
  INV_X1 U11787 ( .A(n12272), .ZN(n16565) );
  NAND2_X1 U11788 ( .A1(n12991), .A2(n16565), .ZN(n12646) );
  INV_X1 U11789 ( .A(n12639), .ZN(n16543) );
  AND2_X1 U11790 ( .A1(n12640), .A2(n16543), .ZN(n12224) );
  NOR2_X1 U11791 ( .A1(n12751), .A2(n12224), .ZN(n9963) );
  NAND2_X1 U11792 ( .A1(n12267), .A2(n16565), .ZN(n9964) );
  NAND2_X1 U11793 ( .A1(n9813), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9972) );
  INV_X1 U11794 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n16590) );
  OR2_X1 U11795 ( .A1(n9814), .A2(n16590), .ZN(n9971) );
  INV_X1 U11796 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n9965) );
  NAND2_X1 U11797 ( .A1(n9967), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9968) );
  AND2_X1 U11798 ( .A1(n9995), .A2(n9968), .ZN(n12410) );
  OR2_X1 U11799 ( .A1(n9815), .A2(n12410), .ZN(n9970) );
  INV_X1 U11800 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n13029) );
  OR2_X1 U11801 ( .A1(n9817), .A2(n13029), .ZN(n9969) );
  XNOR2_X1 U11802 ( .A(n9986), .B(P1_DATAO_REG_12__SCAN_IN), .ZN(n9988) );
  XNOR2_X1 U11803 ( .A(n9989), .B(n9988), .ZN(n10451) );
  NAND2_X1 U11804 ( .A1(n10451), .A2(n12568), .ZN(n9984) );
  NOR2_X1 U11805 ( .A1(n9981), .A2(n13843), .ZN(n9978) );
  MUX2_X1 U11806 ( .A(n13843), .B(n9978), .S(P3_IR_REG_12__SCAN_IN), .Z(n9979)
         );
  INV_X1 U11807 ( .A(n9979), .ZN(n9982) );
  INV_X1 U11808 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n9980) );
  NAND2_X1 U11809 ( .A1(n9981), .A2(n9980), .ZN(n10008) );
  NAND2_X1 U11810 ( .A1(n9982), .A2(n10008), .ZN(n16166) );
  AOI22_X1 U11811 ( .A1(n12562), .A2(n13436), .B1(n10088), .B2(n16166), .ZN(
        n9983) );
  NAND2_X1 U11812 ( .A1(n12452), .A2(n12412), .ZN(n12401) );
  NAND2_X1 U11813 ( .A1(n12362), .A2(n12401), .ZN(n9985) );
  NAND2_X1 U11814 ( .A1(n12228), .A2(n16583), .ZN(n12404) );
  NAND2_X1 U11815 ( .A1(n9985), .A2(n12404), .ZN(n12451) );
  NAND2_X1 U11816 ( .A1(n9986), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9987) );
  XNOR2_X1 U11817 ( .A(n10003), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10464) );
  NAND2_X1 U11818 ( .A1(n10464), .A2(n12568), .ZN(n9993) );
  NAND2_X1 U11819 ( .A1(n10008), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9991) );
  INV_X1 U11820 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9990) );
  XNOR2_X1 U11821 ( .A(n9991), .B(n9990), .ZN(n13052) );
  AOI22_X1 U11822 ( .A1(n12562), .A2(n13629), .B1(n10088), .B2(n13052), .ZN(
        n9992) );
  NAND2_X1 U11823 ( .A1(n9813), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n10000) );
  INV_X1 U11824 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12454) );
  OR2_X1 U11825 ( .A1(n9817), .A2(n12454), .ZN(n9999) );
  INV_X1 U11826 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n13690) );
  NAND2_X1 U11827 ( .A1(n9995), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9996) );
  AND2_X1 U11828 ( .A1(n10013), .A2(n9996), .ZN(n12931) );
  OR2_X1 U11829 ( .A1(n9815), .A2(n12931), .ZN(n9998) );
  NAND2_X1 U11830 ( .A1(n11433), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9997) );
  NAND4_X1 U11831 ( .A1(n10000), .A2(n9999), .A3(n9998), .A4(n9997), .ZN(
        n12990) );
  INV_X1 U11832 ( .A(n12990), .ZN(n10001) );
  AND2_X1 U11833 ( .A1(n16594), .A2(n10001), .ZN(n10002) );
  OR2_X1 U11834 ( .A1(n16594), .A2(n10001), .ZN(n12800) );
  INV_X1 U11835 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10004) );
  XNOR2_X1 U11836 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n10021) );
  XNOR2_X1 U11837 ( .A(n10022), .B(n10021), .ZN(n10466) );
  NAND2_X1 U11838 ( .A1(n10466), .A2(n12568), .ZN(n10012) );
  NAND2_X1 U11839 ( .A1(n10025), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10010) );
  XNOR2_X1 U11840 ( .A(n10010), .B(n10009), .ZN(n16204) );
  AOI22_X1 U11841 ( .A1(n12562), .A2(n10465), .B1(n10088), .B2(n16204), .ZN(
        n10011) );
  NAND2_X1 U11842 ( .A1(n11433), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n10018) );
  NAND2_X1 U11843 ( .A1(n10013), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n10014) );
  AND2_X1 U11844 ( .A1(n10031), .A2(n10014), .ZN(n13305) );
  OR2_X1 U11845 ( .A1(n9815), .A2(n13305), .ZN(n10017) );
  INV_X1 U11846 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13306) );
  OR2_X1 U11847 ( .A1(n9817), .A2(n13306), .ZN(n10016) );
  NAND2_X1 U11848 ( .A1(n9813), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n10015) );
  NOR2_X1 U11849 ( .A1(n13836), .A2(n12989), .ZN(n12663) );
  INV_X1 U11850 ( .A(n12663), .ZN(n10019) );
  NAND2_X1 U11851 ( .A1(n13836), .A2(n12989), .ZN(n12662) );
  NAND2_X1 U11852 ( .A1(n13300), .A2(n13301), .ZN(n13284) );
  INV_X1 U11853 ( .A(n12989), .ZN(n10020) );
  OR2_X1 U11854 ( .A1(n13836), .A2(n10020), .ZN(n13285) );
  NAND2_X1 U11855 ( .A1(n13284), .A2(n13285), .ZN(n10037) );
  INV_X1 U11856 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10023) );
  NAND2_X1 U11857 ( .A1(n10023), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n10024) );
  XNOR2_X1 U11858 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n10039) );
  XNOR2_X1 U11859 ( .A(n10040), .B(n10039), .ZN(n10476) );
  NAND2_X1 U11860 ( .A1(n10476), .A2(n12568), .ZN(n10029) );
  OAI21_X1 U11861 ( .B1(n10025), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n10027) );
  INV_X1 U11862 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n10026) );
  XNOR2_X1 U11863 ( .A(n10027), .B(n10026), .ZN(n13055) );
  AOI22_X1 U11864 ( .A1(n12562), .A2(n13428), .B1(n10088), .B2(n13055), .ZN(
        n10028) );
  INV_X1 U11865 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n16234) );
  OR2_X1 U11866 ( .A1(n9814), .A2(n16234), .ZN(n10036) );
  INV_X1 U11867 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n13702) );
  NAND2_X1 U11868 ( .A1(n10031), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n10032) );
  AND2_X1 U11869 ( .A1(n10045), .A2(n10032), .ZN(n12974) );
  OR2_X1 U11870 ( .A1(n9815), .A2(n12974), .ZN(n10035) );
  INV_X1 U11871 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n16224) );
  OR2_X1 U11872 ( .A1(n9817), .A2(n16224), .ZN(n10034) );
  NAND2_X1 U11873 ( .A1(n9813), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n10033) );
  NAND4_X1 U11874 ( .A1(n10036), .A2(n10035), .A3(n10034), .A4(n10033), .ZN(
        n12903) );
  NAND2_X1 U11875 ( .A1(n13832), .A2(n12903), .ZN(n12669) );
  NAND2_X1 U11876 ( .A1(n12670), .A2(n12669), .ZN(n12665) );
  NAND2_X1 U11877 ( .A1(n10037), .A2(n12665), .ZN(n13287) );
  INV_X1 U11878 ( .A(n12903), .ZN(n13274) );
  OR2_X1 U11879 ( .A1(n13832), .A2(n13274), .ZN(n10038) );
  NAND2_X1 U11880 ( .A1(n13287), .A2(n10038), .ZN(n13271) );
  INV_X1 U11881 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11264) );
  XNOR2_X1 U11882 ( .A(n11474), .B(P1_DATAO_REG_16__SCAN_IN), .ZN(n10054) );
  XNOR2_X1 U11883 ( .A(n10056), .B(n10054), .ZN(n10516) );
  NAND2_X1 U11884 ( .A1(n10516), .A2(n12568), .ZN(n10044) );
  NAND2_X1 U11885 ( .A1(n10041), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10042) );
  XNOR2_X1 U11886 ( .A(n10042), .B(P3_IR_REG_16__SCAN_IN), .ZN(n16250) );
  AOI22_X1 U11887 ( .A1(n12562), .A2(SI_16_), .B1(n10088), .B2(n16250), .ZN(
        n10043) );
  NAND2_X1 U11888 ( .A1(n10044), .A2(n10043), .ZN(n12897) );
  NAND2_X1 U11889 ( .A1(n9813), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n10050) );
  INV_X1 U11890 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13370) );
  OR2_X1 U11891 ( .A1(n9814), .A2(n13370), .ZN(n10049) );
  NAND2_X1 U11892 ( .A1(n10045), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n10046) );
  AND2_X1 U11893 ( .A1(n10062), .A2(n10046), .ZN(n13276) );
  OR2_X1 U11894 ( .A1(n9815), .A2(n13276), .ZN(n10048) );
  INV_X1 U11895 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13277) );
  OR2_X1 U11896 ( .A1(n9817), .A2(n13277), .ZN(n10047) );
  OR2_X1 U11897 ( .A1(n12897), .A2(n12988), .ZN(n10051) );
  NAND2_X1 U11898 ( .A1(n13271), .A2(n10051), .ZN(n10053) );
  NAND2_X1 U11899 ( .A1(n12897), .A2(n12988), .ZN(n10052) );
  INV_X1 U11900 ( .A(n10054), .ZN(n10055) );
  NAND2_X1 U11901 ( .A1(n11474), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n10057) );
  XNOR2_X1 U11902 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n10069) );
  XNOR2_X1 U11903 ( .A(n10070), .B(n10069), .ZN(n10549) );
  NAND2_X1 U11904 ( .A1(n10549), .A2(n12568), .ZN(n10060) );
  NAND2_X1 U11905 ( .A1(n7597), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10058) );
  XNOR2_X1 U11906 ( .A(n10058), .B(P3_IR_REG_17__SCAN_IN), .ZN(n16268) );
  INV_X1 U11907 ( .A(n16268), .ZN(n13039) );
  AOI22_X1 U11908 ( .A1(n12562), .A2(n10548), .B1(n10088), .B2(n13039), .ZN(
        n10059) );
  INV_X1 U11909 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13258) );
  OR2_X1 U11910 ( .A1(n9817), .A2(n13258), .ZN(n10067) );
  INV_X1 U11911 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n13680) );
  NAND2_X1 U11912 ( .A1(n10062), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n10063) );
  AND2_X1 U11913 ( .A1(n10075), .A2(n10063), .ZN(n13257) );
  OR2_X1 U11914 ( .A1(n9815), .A2(n13257), .ZN(n10066) );
  INV_X1 U11915 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n16271) );
  OR2_X1 U11916 ( .A1(n9814), .A2(n16271), .ZN(n10065) );
  NAND2_X1 U11917 ( .A1(n9813), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n10064) );
  NAND4_X1 U11918 ( .A1(n10067), .A2(n10066), .A3(n10065), .A4(n10064), .ZN(
        n12958) );
  OR2_X1 U11919 ( .A1(n13824), .A2(n12958), .ZN(n12680) );
  NAND2_X1 U11920 ( .A1(n13824), .A2(n12958), .ZN(n12683) );
  INV_X1 U11921 ( .A(n12958), .ZN(n13275) );
  OR2_X1 U11922 ( .A1(n13824), .A2(n13275), .ZN(n10068) );
  INV_X1 U11923 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11547) );
  XNOR2_X1 U11924 ( .A(n11588), .B(P1_DATAO_REG_18__SCAN_IN), .ZN(n10081) );
  XNOR2_X1 U11925 ( .A(n10083), .B(n10081), .ZN(n10702) );
  NAND2_X1 U11926 ( .A1(n10702), .A2(n12568), .ZN(n10074) );
  NAND2_X1 U11927 ( .A1(n10071), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10072) );
  XNOR2_X1 U11928 ( .A(n10072), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13077) );
  AOI22_X1 U11929 ( .A1(n12562), .A2(SI_18_), .B1(n10088), .B2(n13077), .ZN(
        n10073) );
  NAND2_X1 U11930 ( .A1(n11433), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n10080) );
  NAND2_X1 U11931 ( .A1(n9813), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n10079) );
  NAND2_X1 U11932 ( .A1(n10075), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n10076) );
  AND2_X1 U11933 ( .A1(n10092), .A2(n10076), .ZN(n13243) );
  OR2_X1 U11934 ( .A1(n9815), .A2(n13243), .ZN(n10078) );
  NAND2_X1 U11935 ( .A1(n9770), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n10077) );
  NAND4_X1 U11936 ( .A1(n10080), .A2(n10079), .A3(n10078), .A4(n10077), .ZN(
        n13252) );
  AND2_X1 U11937 ( .A1(n13820), .A2(n13252), .ZN(n10288) );
  INV_X1 U11938 ( .A(n13820), .ZN(n12677) );
  NAND2_X1 U11939 ( .A1(n12677), .A2(n13226), .ZN(n13238) );
  NAND2_X1 U11940 ( .A1(n10289), .A2(n13238), .ZN(n13234) );
  INV_X1 U11941 ( .A(n13234), .ZN(n13239) );
  OR2_X1 U11942 ( .A1(n12677), .A2(n13252), .ZN(n12679) );
  INV_X1 U11943 ( .A(n10081), .ZN(n10082) );
  NAND2_X1 U11944 ( .A1(n11588), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n10084) );
  INV_X1 U11945 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11601) );
  XNOR2_X1 U11946 ( .A(n11601), .B(P1_DATAO_REG_19__SCAN_IN), .ZN(n10101) );
  XNOR2_X1 U11947 ( .A(n10103), .B(n10101), .ZN(n10875) );
  NAND2_X1 U11948 ( .A1(n10875), .A2(n12568), .ZN(n10090) );
  INV_X1 U11949 ( .A(n10071), .ZN(n10086) );
  INV_X1 U11950 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n10085) );
  NAND2_X1 U11951 ( .A1(n10254), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10087) );
  AOI22_X1 U11952 ( .A1(n12562), .A2(SI_19_), .B1(n13086), .B2(n10088), .ZN(
        n10089) );
  NAND2_X1 U11953 ( .A1(n9813), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n10097) );
  INV_X1 U11954 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13358) );
  OR2_X1 U11955 ( .A1(n9814), .A2(n13358), .ZN(n10096) );
  INV_X1 U11956 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n13469) );
  NAND2_X1 U11957 ( .A1(n10092), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n10093) );
  AND2_X1 U11958 ( .A1(n10106), .A2(n10093), .ZN(n13228) );
  OR2_X1 U11959 ( .A1(n9815), .A2(n13228), .ZN(n10095) );
  INV_X1 U11960 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13229) );
  OR2_X1 U11961 ( .A1(n9817), .A2(n13229), .ZN(n10094) );
  NAND2_X1 U11962 ( .A1(n12875), .A2(n12987), .ZN(n10098) );
  NAND2_X1 U11963 ( .A1(n13223), .A2(n10098), .ZN(n10100) );
  OR2_X1 U11964 ( .A1(n12875), .A2(n12987), .ZN(n10099) );
  INV_X1 U11965 ( .A(n10101), .ZN(n10102) );
  XNOR2_X1 U11966 ( .A(n10114), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n11214) );
  NAND2_X1 U11967 ( .A1(n11214), .A2(n12568), .ZN(n10105) );
  OR2_X1 U11968 ( .A1(n12569), .A2(n7989), .ZN(n10104) );
  NAND2_X1 U11969 ( .A1(n10106), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n10107) );
  NAND2_X1 U11970 ( .A1(n10123), .A2(n10107), .ZN(n13217) );
  NAND2_X1 U11971 ( .A1(n10247), .A2(n13217), .ZN(n10112) );
  INV_X1 U11972 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13354) );
  OR2_X1 U11973 ( .A1(n9814), .A2(n13354), .ZN(n10111) );
  INV_X1 U11974 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13810) );
  OR2_X1 U11975 ( .A1(n11436), .A2(n13810), .ZN(n10110) );
  INV_X1 U11976 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n10108) );
  OR2_X1 U11977 ( .A1(n9817), .A2(n10108), .ZN(n10109) );
  NAND2_X1 U11978 ( .A1(n13216), .A2(n13227), .ZN(n12695) );
  INV_X1 U11979 ( .A(n13227), .ZN(n12986) );
  NAND2_X1 U11980 ( .A1(n13216), .A2(n12986), .ZN(n10113) );
  NAND2_X1 U11981 ( .A1(n10115), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n10116) );
  INV_X1 U11982 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11678) );
  XNOR2_X1 U11983 ( .A(n11678), .B(P1_DATAO_REG_21__SCAN_IN), .ZN(n10129) );
  XNOR2_X1 U11984 ( .A(n10131), .B(n10129), .ZN(n11374) );
  NAND2_X1 U11985 ( .A1(n11374), .A2(n12568), .ZN(n10119) );
  INV_X1 U11986 ( .A(SI_21_), .ZN(n11376) );
  OR2_X1 U11987 ( .A1(n12569), .A2(n11376), .ZN(n10118) );
  NAND2_X1 U11988 ( .A1(n11433), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n10121) );
  NAND2_X1 U11989 ( .A1(n9813), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n10120) );
  AND2_X1 U11990 ( .A1(n10121), .A2(n10120), .ZN(n10127) );
  INV_X1 U11991 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n13666) );
  NAND2_X1 U11992 ( .A1(n10123), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n10124) );
  NAND2_X1 U11993 ( .A1(n10142), .A2(n10124), .ZN(n13205) );
  NAND2_X1 U11994 ( .A1(n13205), .A2(n10247), .ZN(n10126) );
  NAND2_X1 U11995 ( .A1(n9770), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n10125) );
  NAND2_X1 U11996 ( .A1(n13349), .A2(n12945), .ZN(n12696) );
  INV_X1 U11997 ( .A(n12696), .ZN(n10128) );
  INV_X1 U11998 ( .A(n10129), .ZN(n10130) );
  NAND2_X1 U11999 ( .A1(n10131), .A2(n10130), .ZN(n10133) );
  NAND2_X1 U12000 ( .A1(n11678), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n10132) );
  NAND2_X1 U12001 ( .A1(n11985), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n10149) );
  INV_X1 U12002 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10134) );
  NAND2_X1 U12003 ( .A1(n10134), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n10135) );
  NAND2_X1 U12004 ( .A1(n10149), .A2(n10135), .ZN(n10136) );
  NAND2_X1 U12005 ( .A1(n10137), .A2(n10136), .ZN(n10138) );
  NAND2_X1 U12006 ( .A1(n10150), .A2(n10138), .ZN(n11290) );
  NAND2_X1 U12007 ( .A1(n11290), .A2(n12568), .ZN(n10141) );
  OR2_X1 U12008 ( .A1(n12569), .A2(n10139), .ZN(n10140) );
  NAND2_X1 U12009 ( .A1(n10142), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n10143) );
  NAND2_X1 U12010 ( .A1(n10158), .A2(n10143), .ZN(n13194) );
  NAND2_X1 U12011 ( .A1(n13194), .A2(n10247), .ZN(n10146) );
  AOI22_X1 U12012 ( .A1(n9813), .A2(P3_REG0_REG_22__SCAN_IN), .B1(n11433), 
        .B2(P3_REG1_REG_22__SCAN_IN), .ZN(n10145) );
  NAND2_X1 U12013 ( .A1(n9770), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n10144) );
  NAND2_X1 U12014 ( .A1(n13193), .A2(n12867), .ZN(n12588) );
  INV_X1 U12015 ( .A(n13185), .ZN(n10148) );
  INV_X1 U12016 ( .A(n12867), .ZN(n12944) );
  NAND2_X1 U12017 ( .A1(n13193), .A2(n12944), .ZN(n10147) );
  OAI21_X1 U12018 ( .B1(n13186), .B2(n10148), .A(n10147), .ZN(n13171) );
  NAND2_X1 U12019 ( .A1(n12152), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n10165) );
  NAND2_X1 U12020 ( .A1(n10151), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n10152) );
  AND2_X1 U12021 ( .A1(n10165), .A2(n10152), .ZN(n10153) );
  OR2_X1 U12022 ( .A1(n10154), .A2(n10153), .ZN(n10155) );
  NAND2_X1 U12023 ( .A1(n10166), .A2(n10155), .ZN(n11551) );
  NAND2_X1 U12024 ( .A1(n11551), .A2(n12568), .ZN(n10157) );
  OR2_X1 U12025 ( .A1(n12569), .A2(n13614), .ZN(n10156) );
  NAND2_X1 U12026 ( .A1(n10158), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n10159) );
  NAND2_X1 U12027 ( .A1(n10171), .A2(n10159), .ZN(n12866) );
  NAND2_X1 U12028 ( .A1(n12866), .A2(n10247), .ZN(n10162) );
  AOI22_X1 U12029 ( .A1(n9813), .A2(P3_REG0_REG_23__SCAN_IN), .B1(n11433), 
        .B2(P3_REG1_REG_23__SCAN_IN), .ZN(n10161) );
  NAND2_X1 U12030 ( .A1(n9770), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n10160) );
  NAND2_X1 U12031 ( .A1(n13400), .A2(n13188), .ZN(n12706) );
  NAND2_X1 U12032 ( .A1(n13171), .A2(n13176), .ZN(n10164) );
  INV_X1 U12033 ( .A(n13188), .ZN(n12985) );
  NAND2_X1 U12034 ( .A1(n13400), .A2(n12985), .ZN(n10163) );
  NAND2_X1 U12035 ( .A1(n10164), .A2(n10163), .ZN(n13153) );
  XNOR2_X1 U12036 ( .A(n10181), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n11682) );
  NAND2_X1 U12037 ( .A1(n11682), .A2(n12568), .ZN(n10168) );
  INV_X1 U12038 ( .A(SI_24_), .ZN(n11683) );
  OR2_X1 U12039 ( .A1(n12569), .A2(n11683), .ZN(n10167) );
  INV_X1 U12040 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n10169) );
  NAND2_X1 U12041 ( .A1(n10171), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n10172) );
  NAND2_X1 U12042 ( .A1(n10186), .A2(n10172), .ZN(n13165) );
  NAND2_X1 U12043 ( .A1(n13165), .A2(n10247), .ZN(n10177) );
  INV_X1 U12044 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13394) );
  NAND2_X1 U12045 ( .A1(n11433), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n10174) );
  NAND2_X1 U12046 ( .A1(n9770), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n10173) );
  OAI211_X1 U12047 ( .C1(n11436), .C2(n13394), .A(n10174), .B(n10173), .ZN(
        n10175) );
  INV_X1 U12048 ( .A(n10175), .ZN(n10176) );
  AND2_X1 U12049 ( .A1(n13164), .A2(n12832), .ZN(n10179) );
  NAND2_X1 U12050 ( .A1(n12534), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n10182) );
  XNOR2_X1 U12051 ( .A(n10194), .B(n10193), .ZN(n11885) );
  NAND2_X1 U12052 ( .A1(n11885), .A2(n12568), .ZN(n10184) );
  OR2_X1 U12053 ( .A1(n12569), .A2(n13610), .ZN(n10183) );
  INV_X1 U12054 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n13675) );
  NAND2_X1 U12055 ( .A1(n10186), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n10187) );
  NAND2_X1 U12056 ( .A1(n10199), .A2(n10187), .ZN(n13148) );
  INV_X1 U12057 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n10190) );
  NAND2_X1 U12058 ( .A1(n11433), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n10189) );
  NAND2_X1 U12059 ( .A1(n9770), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n10188) );
  OAI211_X1 U12060 ( .C1(n11436), .C2(n10190), .A(n10189), .B(n10188), .ZN(
        n10191) );
  NAND2_X1 U12061 ( .A1(n13330), .A2(n12915), .ZN(n12710) );
  INV_X1 U12062 ( .A(n12915), .ZN(n12984) );
  NAND2_X1 U12063 ( .A1(n13330), .A2(n12984), .ZN(n10192) );
  NAND2_X1 U12064 ( .A1(n14788), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n10211) );
  NAND2_X1 U12065 ( .A1(n15778), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n10196) );
  AND2_X1 U12066 ( .A1(n10211), .A2(n10196), .ZN(n10209) );
  XNOR2_X1 U12067 ( .A(n10210), .B(n10209), .ZN(n12028) );
  NAND2_X1 U12068 ( .A1(n12028), .A2(n12568), .ZN(n10198) );
  INV_X1 U12069 ( .A(SI_26_), .ZN(n12030) );
  OR2_X1 U12070 ( .A1(n12569), .A2(n12030), .ZN(n10197) );
  NAND2_X1 U12071 ( .A1(n10199), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n10200) );
  NAND2_X1 U12072 ( .A1(n10216), .A2(n10200), .ZN(n13136) );
  NAND2_X1 U12073 ( .A1(n13136), .A2(n10247), .ZN(n10206) );
  INV_X1 U12074 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n10203) );
  NAND2_X1 U12075 ( .A1(n11433), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n10202) );
  NAND2_X1 U12076 ( .A1(n9770), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n10201) );
  OAI211_X1 U12077 ( .C1(n11436), .C2(n10203), .A(n10202), .B(n10201), .ZN(
        n10204) );
  INV_X1 U12078 ( .A(n10204), .ZN(n10205) );
  NAND2_X1 U12079 ( .A1(n13326), .A2(n12983), .ZN(n10207) );
  NAND2_X1 U12080 ( .A1(n10208), .A2(n10207), .ZN(n13122) );
  INV_X1 U12081 ( .A(n13122), .ZN(n10224) );
  NAND2_X1 U12082 ( .A1(n10210), .A2(n10209), .ZN(n10212) );
  XNOR2_X1 U12083 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n10227) );
  XNOR2_X1 U12084 ( .A(n10229), .B(n10227), .ZN(n12170) );
  NAND2_X1 U12085 ( .A1(n12170), .A2(n12568), .ZN(n10214) );
  INV_X1 U12086 ( .A(SI_27_), .ZN(n12171) );
  OR2_X1 U12087 ( .A1(n12569), .A2(n12171), .ZN(n10213) );
  INV_X1 U12088 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n13461) );
  NAND2_X1 U12089 ( .A1(n10216), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n10217) );
  NAND2_X1 U12090 ( .A1(n10234), .A2(n10217), .ZN(n13127) );
  NAND2_X1 U12091 ( .A1(n13127), .A2(n10247), .ZN(n10223) );
  INV_X1 U12092 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n10220) );
  NAND2_X1 U12093 ( .A1(n11433), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n10219) );
  NAND2_X1 U12094 ( .A1(n9770), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n10218) );
  OAI211_X1 U12095 ( .C1(n11436), .C2(n10220), .A(n10219), .B(n10218), .ZN(
        n10221) );
  INV_X1 U12096 ( .A(n10221), .ZN(n10222) );
  INV_X1 U12097 ( .A(n10227), .ZN(n10228) );
  NAND2_X1 U12098 ( .A1(n15776), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n10230) );
  XNOR2_X1 U12099 ( .A(n10242), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n10231) );
  XNOR2_X1 U12100 ( .A(n10241), .B(n10231), .ZN(n12531) );
  NAND2_X1 U12101 ( .A1(n12531), .A2(n12568), .ZN(n10233) );
  OR2_X1 U12102 ( .A1(n12569), .A2(n13410), .ZN(n10232) );
  NAND2_X1 U12103 ( .A1(n10234), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n10235) );
  NAND2_X1 U12104 ( .A1(n13092), .A2(n10235), .ZN(n13114) );
  INV_X1 U12105 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13389) );
  NAND2_X1 U12106 ( .A1(n9770), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n10237) );
  NAND2_X1 U12107 ( .A1(n11433), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n10236) );
  OAI211_X1 U12108 ( .C1(n11436), .C2(n13389), .A(n10237), .B(n10236), .ZN(
        n10238) );
  NAND2_X1 U12109 ( .A1(n13113), .A2(n13125), .ZN(n12722) );
  INV_X1 U12110 ( .A(n13125), .ZN(n12982) );
  AND2_X1 U12111 ( .A1(n15774), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n10240) );
  NAND2_X1 U12112 ( .A1(n10242), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n10243) );
  XNOR2_X1 U12113 ( .A(n15771), .B(P1_DATAO_REG_29__SCAN_IN), .ZN(n12555) );
  INV_X1 U12114 ( .A(n12555), .ZN(n10244) );
  NAND2_X1 U12115 ( .A1(n13849), .A2(n12568), .ZN(n10246) );
  OR2_X1 U12116 ( .A1(n12569), .A2(n13851), .ZN(n10245) );
  INV_X1 U12117 ( .A(n13092), .ZN(n10248) );
  NAND2_X1 U12118 ( .A1(n10248), .A2(n10247), .ZN(n11439) );
  INV_X1 U12119 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n10352) );
  NAND2_X1 U12120 ( .A1(n11433), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U12121 ( .A1(n9770), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n10249) );
  OAI211_X1 U12122 ( .C1(n11436), .C2(n10352), .A(n10250), .B(n10249), .ZN(
        n10251) );
  INV_X1 U12123 ( .A(n10251), .ZN(n10252) );
  NAND2_X1 U12124 ( .A1(n10343), .A2(n13109), .ZN(n12582) );
  XNOR2_X1 U12125 ( .A(n10253), .B(n12762), .ZN(n10276) );
  NAND2_X1 U12126 ( .A1(n10306), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10257) );
  AND2_X1 U12127 ( .A1(n12773), .A2(n13086), .ZN(n10298) );
  INV_X1 U12128 ( .A(n10298), .ZN(n10264) );
  NAND2_X1 U12129 ( .A1(n10262), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10258) );
  NAND2_X1 U12130 ( .A1(n10260), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10261) );
  MUX2_X1 U12131 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10261), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n10263) );
  NAND2_X1 U12132 ( .A1(n12594), .A2(n10303), .ZN(n12580) );
  INV_X1 U12133 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n13387) );
  NAND2_X1 U12134 ( .A1(n11433), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n10266) );
  NAND2_X1 U12135 ( .A1(n9770), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n10265) );
  OAI211_X1 U12136 ( .C1(n11436), .C2(n13387), .A(n10266), .B(n10265), .ZN(
        n10267) );
  INV_X1 U12137 ( .A(n10267), .ZN(n10268) );
  INV_X1 U12138 ( .A(n7430), .ZN(n12770) );
  NAND2_X1 U12139 ( .A1(n12770), .A2(n10990), .ZN(n11016) );
  NAND2_X1 U12140 ( .A1(n11016), .A2(n9860), .ZN(n10272) );
  INV_X1 U12141 ( .A(P3_B_REG_SCAN_IN), .ZN(n13506) );
  NOR2_X1 U12142 ( .A1(n7430), .A2(n13506), .ZN(n10271) );
  OR2_X1 U12143 ( .A1(n16352), .A2(n10271), .ZN(n13090) );
  NOR2_X1 U12144 ( .A1(n12574), .A2(n13090), .ZN(n10274) );
  NAND2_X1 U12145 ( .A1(n12597), .A2(n16308), .ZN(n10279) );
  INV_X1 U12146 ( .A(n16355), .ZN(n10280) );
  NAND2_X1 U12147 ( .A1(n16353), .A2(n12600), .ZN(n10282) );
  NAND2_X1 U12148 ( .A1(n11731), .A2(n12608), .ZN(n10283) );
  NAND2_X1 U12149 ( .A1(n10283), .A2(n12610), .ZN(n11590) );
  NAND2_X1 U12150 ( .A1(n12622), .A2(n12620), .ZN(n10284) );
  NAND2_X1 U12151 ( .A1(n11846), .A2(n12624), .ZN(n11845) );
  NAND2_X1 U12152 ( .A1(n11845), .A2(n12626), .ZN(n11870) );
  NOR2_X1 U12153 ( .A1(n12992), .A2(n16523), .ZN(n12121) );
  NAND2_X1 U12154 ( .A1(n12992), .A2(n16523), .ZN(n12635) );
  INV_X1 U12155 ( .A(n12640), .ZN(n12229) );
  NAND2_X1 U12156 ( .A1(n12229), .A2(n16543), .ZN(n12641) );
  NAND2_X1 U12157 ( .A1(n12233), .A2(n12751), .ZN(n10285) );
  NAND2_X1 U12158 ( .A1(n10285), .A2(n12651), .ZN(n12361) );
  NAND2_X1 U12159 ( .A1(n12228), .A2(n12412), .ZN(n12652) );
  NAND2_X1 U12160 ( .A1(n12452), .A2(n16583), .ZN(n12653) );
  NAND2_X1 U12161 ( .A1(n12361), .A2(n12750), .ZN(n12360) );
  NAND2_X1 U12162 ( .A1(n12360), .A2(n12652), .ZN(n12450) );
  NAND2_X1 U12163 ( .A1(n16594), .A2(n12990), .ZN(n12799) );
  NAND2_X1 U12164 ( .A1(n12450), .A2(n12796), .ZN(n10286) );
  NAND2_X1 U12165 ( .A1(n13282), .A2(n12670), .ZN(n13269) );
  AND2_X1 U12166 ( .A1(n12897), .A2(n13254), .ZN(n12668) );
  OR2_X1 U12167 ( .A1(n12897), .A2(n13254), .ZN(n12673) );
  NAND2_X1 U12168 ( .A1(n12875), .A2(n13237), .ZN(n12735) );
  AND2_X1 U12169 ( .A1(n13238), .A2(n12735), .ZN(n10290) );
  NAND2_X1 U12170 ( .A1(n13349), .A2(n13187), .ZN(n12586) );
  NAND2_X1 U12171 ( .A1(n13200), .A2(n12586), .ZN(n10292) );
  OR2_X1 U12172 ( .A1(n13349), .A2(n13187), .ZN(n10291) );
  NAND2_X1 U12173 ( .A1(n10292), .A2(n10291), .ZN(n13184) );
  INV_X1 U12174 ( .A(n13184), .ZN(n10293) );
  NAND2_X1 U12175 ( .A1(n13164), .A2(n12891), .ZN(n12709) );
  AND2_X1 U12176 ( .A1(n10294), .A2(n13159), .ZN(n10295) );
  NAND2_X1 U12177 ( .A1(n13160), .A2(n10295), .ZN(n13143) );
  NAND2_X1 U12178 ( .A1(n13326), .A2(n13126), .ZN(n12714) );
  INV_X1 U12179 ( .A(n12726), .ZN(n10296) );
  XNOR2_X1 U12180 ( .A(n12573), .B(n12762), .ZN(n13096) );
  NAND2_X1 U12181 ( .A1(n10298), .A2(n10297), .ZN(n10805) );
  AND2_X1 U12182 ( .A1(n10805), .A2(n12731), .ZN(n10300) );
  INV_X1 U12183 ( .A(n12773), .ZN(n10299) );
  NAND2_X1 U12184 ( .A1(n11216), .A2(n13086), .ZN(n12733) );
  NAND2_X1 U12185 ( .A1(n10300), .A2(n10809), .ZN(n10803) );
  INV_X1 U12186 ( .A(n10803), .ZN(n10302) );
  INV_X1 U12187 ( .A(n13086), .ZN(n10878) );
  NAND2_X1 U12188 ( .A1(n11216), .A2(n10878), .ZN(n12732) );
  INV_X1 U12189 ( .A(n12732), .ZN(n10346) );
  AND2_X1 U12190 ( .A1(n16593), .A2(n10346), .ZN(n10301) );
  NAND2_X1 U12191 ( .A1(n10302), .A2(n10301), .ZN(n10305) );
  AND2_X1 U12192 ( .A1(n10303), .A2(n10878), .ZN(n10304) );
  NAND2_X1 U12193 ( .A1(n12773), .A2(n10304), .ZN(n10336) );
  OR2_X1 U12194 ( .A1(n12773), .A2(n12733), .ZN(n16584) );
  NOR2_X1 U12195 ( .A1(n13101), .A2(n8516), .ZN(n10351) );
  OAI21_X1 U12196 ( .B1(n10306), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n10308) );
  INV_X1 U12197 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n10307) );
  XNOR2_X1 U12198 ( .A(n10308), .B(n10307), .ZN(n10987) );
  NAND2_X1 U12199 ( .A1(n7560), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10309) );
  MUX2_X1 U12200 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10309), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n10311) );
  NAND2_X1 U12201 ( .A1(n10312), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10313) );
  MUX2_X1 U12202 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10313), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n10314) );
  AND2_X1 U12203 ( .A1(n10314), .A2(n7560), .ZN(n10318) );
  MUX2_X1 U12204 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7569), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n10316) );
  NAND2_X1 U12205 ( .A1(n10318), .A2(n11681), .ZN(n10317) );
  NOR2_X1 U12206 ( .A1(n12031), .A2(n10317), .ZN(n10353) );
  INV_X1 U12207 ( .A(n10318), .ZN(n11887) );
  NAND2_X1 U12208 ( .A1(n11887), .A2(n10319), .ZN(n10320) );
  NOR2_X1 U12209 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n10324) );
  NOR4_X1 U12210 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n10323) );
  NOR4_X1 U12211 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n10322) );
  NOR4_X1 U12212 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n10321) );
  NAND4_X1 U12213 ( .A1(n10324), .A2(n10323), .A3(n10322), .A4(n10321), .ZN(
        n10330) );
  NOR4_X1 U12214 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n10328) );
  NOR4_X1 U12215 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n10327) );
  NOR4_X1 U12216 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n10326) );
  NOR4_X1 U12217 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n10325) );
  NAND4_X1 U12218 ( .A1(n10328), .A2(n10327), .A3(n10326), .A4(n10325), .ZN(
        n10329) );
  NOR2_X1 U12219 ( .A1(n10330), .A2(n10329), .ZN(n10331) );
  NOR2_X1 U12220 ( .A1(n12527), .A2(n10331), .ZN(n10344) );
  INV_X1 U12221 ( .A(n10344), .ZN(n10348) );
  NAND2_X1 U12222 ( .A1(n10811), .A2(n10348), .ZN(n10335) );
  NAND2_X1 U12223 ( .A1(n12031), .A2(n11887), .ZN(n10333) );
  XNOR2_X1 U12224 ( .A(n10945), .B(n11443), .ZN(n10334) );
  INV_X1 U12225 ( .A(n11443), .ZN(n13839) );
  NAND2_X1 U12226 ( .A1(n12728), .A2(n12732), .ZN(n10792) );
  NAND2_X1 U12227 ( .A1(n12731), .A2(n10336), .ZN(n10337) );
  NAND2_X1 U12228 ( .A1(n10792), .A2(n10337), .ZN(n11442) );
  NAND2_X1 U12229 ( .A1(n13839), .A2(n11442), .ZN(n10340) );
  INV_X1 U12230 ( .A(n10337), .ZN(n11444) );
  NAND2_X1 U12231 ( .A1(n10809), .A2(n11444), .ZN(n10338) );
  NAND2_X1 U12232 ( .A1(n10338), .A2(n11443), .ZN(n10339) );
  NAND2_X1 U12233 ( .A1(n10340), .A2(n10339), .ZN(n10341) );
  OR2_X1 U12234 ( .A1(n11443), .A2(n10344), .ZN(n10345) );
  NOR2_X1 U12235 ( .A1(n10345), .A2(n10945), .ZN(n10795) );
  AND2_X1 U12236 ( .A1(n10795), .A2(n10811), .ZN(n10808) );
  NAND2_X1 U12237 ( .A1(n12728), .A2(n10346), .ZN(n10879) );
  NAND2_X1 U12238 ( .A1(n10879), .A2(n10805), .ZN(n10347) );
  NAND2_X1 U12239 ( .A1(n10808), .A2(n10347), .ZN(n10350) );
  AND3_X1 U12240 ( .A1(n10945), .A2(n11443), .A3(n10348), .ZN(n10797) );
  NAND2_X1 U12241 ( .A1(n10797), .A2(n10811), .ZN(n10814) );
  OR2_X1 U12242 ( .A1(n10814), .A2(n10803), .ZN(n10349) );
  NAND2_X1 U12243 ( .A1(n10578), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10469) );
  OR2_X1 U12244 ( .A1(n11177), .A2(n10469), .ZN(n12529) );
  INV_X2 U12245 ( .A(n12529), .ZN(P1_U4016) );
  INV_X1 U12246 ( .A(n10353), .ZN(n10791) );
  OR2_X2 U12247 ( .A1(n10791), .A2(n13838), .ZN(n12998) );
  XNOR2_X1 U12248 ( .A(n14041), .B(n14362), .ZN(n14288) );
  XNOR2_X1 U12249 ( .A(n10355), .B(n14288), .ZN(n10356) );
  INV_X1 U12250 ( .A(n14588), .ZN(n13967) );
  INV_X1 U12251 ( .A(n14589), .ZN(n13968) );
  OAI22_X1 U12252 ( .A1(n10395), .A2(n13967), .B1(n11311), .B2(n13968), .ZN(
        n10962) );
  AOI21_X1 U12253 ( .B1(n10356), .B2(n14606), .A(n10962), .ZN(n10871) );
  INV_X1 U12254 ( .A(n10871), .ZN(n10360) );
  AND2_X1 U12255 ( .A1(n10358), .A2(n10357), .ZN(n10384) );
  NOR2_X1 U12256 ( .A1(n10385), .A2(n15822), .ZN(n15821) );
  NAND3_X1 U12257 ( .A1(n10384), .A2(n15821), .A3(n10388), .ZN(n10359) );
  INV_X2 U12258 ( .A(n14622), .ZN(n11368) );
  MUX2_X1 U12259 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10360), .S(n11368), .Z(
        n10368) );
  AND2_X1 U12260 ( .A1(n10361), .A2(n11169), .ZN(n10869) );
  AND2_X1 U12261 ( .A1(n14632), .A2(n10869), .ZN(n10367) );
  AND2_X1 U12262 ( .A1(n14332), .A2(n7431), .ZN(n10362) );
  NAND2_X1 U12263 ( .A1(n11368), .A2(n10362), .ZN(n14602) );
  INV_X1 U12264 ( .A(n11636), .ZN(n14591) );
  NAND2_X1 U12265 ( .A1(n11368), .A2(n14591), .ZN(n10363) );
  NAND2_X1 U12266 ( .A1(n14602), .A2(n10363), .ZN(n14630) );
  XNOR2_X1 U12267 ( .A(n10364), .B(n14288), .ZN(n10872) );
  NOR2_X1 U12268 ( .A1(n14580), .A2(n10872), .ZN(n10366) );
  AND2_X1 U12269 ( .A1(n10822), .A2(n14323), .ZN(n10393) );
  OAI22_X1 U12270 ( .A1(n14619), .A2(n7957), .B1(n10965), .B2(n14624), .ZN(
        n10365) );
  OR4_X1 U12271 ( .A1(n10368), .A2(n10367), .A3(n10366), .A4(n10365), .ZN(
        P2_U3260) );
  INV_X1 U12272 ( .A(n10369), .ZN(n10741) );
  NAND2_X1 U12273 ( .A1(n7433), .A2(n14001), .ZN(n10370) );
  NAND2_X1 U12274 ( .A1(n14366), .A2(n7490), .ZN(n10372) );
  XNOR2_X1 U12275 ( .A(n10371), .B(n10372), .ZN(n10650) );
  INV_X1 U12276 ( .A(n10371), .ZN(n10850) );
  NAND2_X1 U12277 ( .A1(n10850), .A2(n10372), .ZN(n10373) );
  NAND2_X1 U12278 ( .A1(n14365), .A2(n7490), .ZN(n10375) );
  XNOR2_X1 U12279 ( .A(n10374), .B(n10375), .ZN(n10851) );
  INV_X1 U12280 ( .A(n10374), .ZN(n10376) );
  NAND2_X1 U12281 ( .A1(n10376), .A2(n10375), .ZN(n10377) );
  XNOR2_X1 U12282 ( .A(n10884), .B(n14027), .ZN(n10891) );
  AND2_X1 U12283 ( .A1(n14364), .A2(n7437), .ZN(n10378) );
  NAND2_X1 U12284 ( .A1(n10891), .A2(n10378), .ZN(n10885) );
  INV_X1 U12285 ( .A(n10886), .ZN(n10890) );
  INV_X1 U12286 ( .A(n15822), .ZN(n10379) );
  AND2_X1 U12287 ( .A1(n10379), .A2(n10385), .ZN(n10380) );
  AND2_X1 U12288 ( .A1(n10384), .A2(n10380), .ZN(n10397) );
  NOR2_X1 U12289 ( .A1(n16382), .A2(n10487), .ZN(n10381) );
  AOI211_X1 U12290 ( .C1(n10383), .C2(n10382), .A(n10890), .B(n13963), .ZN(
        n10401) );
  NAND2_X1 U12291 ( .A1(n10385), .A2(n10384), .ZN(n10387) );
  NAND2_X1 U12292 ( .A1(n10387), .A2(n10386), .ZN(n10392) );
  INV_X1 U12293 ( .A(n10388), .ZN(n10389) );
  NOR2_X1 U12294 ( .A1(n10390), .A2(n10389), .ZN(n10391) );
  NAND2_X1 U12295 ( .A1(n10392), .A2(n10391), .ZN(n10649) );
  MUX2_X1 U12296 ( .A(n13985), .B(P2_U3088), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n10400) );
  NAND2_X1 U12297 ( .A1(n10397), .A2(n10393), .ZN(n10394) );
  INV_X1 U12298 ( .A(n13983), .ZN(n13975) );
  OAI22_X1 U12299 ( .A1(n10648), .A2(n13967), .B1(n10395), .B2(n13968), .ZN(
        n10750) );
  INV_X1 U12300 ( .A(n10750), .ZN(n10398) );
  INV_X1 U12301 ( .A(n10396), .ZN(n14324) );
  NAND2_X1 U12302 ( .A1(n10397), .A2(n14324), .ZN(n13988) );
  OAI22_X1 U12303 ( .A1(n13975), .A2(n10754), .B1(n10398), .B2(n13988), .ZN(
        n10399) );
  OR3_X1 U12304 ( .A1(n10401), .A2(n10400), .A3(n10399), .ZN(P2_U3190) );
  NAND2_X1 U12305 ( .A1(n8402), .A2(n10404), .ZN(n10403) );
  INV_X1 U12306 ( .A(P3_RD_REG_SCAN_IN), .ZN(n10402) );
  OAI211_X1 U12307 ( .C1(n10404), .C2(n8402), .A(n10403), .B(n10402), .ZN(U29)
         );
  INV_X1 U12308 ( .A(n10405), .ZN(n10407) );
  INV_X1 U12309 ( .A(n15364), .ZN(n15362) );
  OAI222_X1 U12310 ( .A1(n15777), .A2(n10406), .B1(n15780), .B2(n10407), .C1(
        P1_U3086), .C2(n15362), .ZN(P1_U3352) );
  INV_X1 U12311 ( .A(n14783), .ZN(n12148) );
  INV_X1 U12312 ( .A(n10499), .ZN(n15824) );
  OAI222_X1 U12313 ( .A1(n14787), .A2(n10408), .B1(n14783), .B2(n10407), .C1(
        P2_U3088), .C2(n15824), .ZN(P2_U3324) );
  INV_X1 U12314 ( .A(n10409), .ZN(n10415) );
  INV_X1 U12315 ( .A(n14385), .ZN(n10410) );
  OAI222_X1 U12316 ( .A1(n14787), .A2(n10411), .B1(n14783), .B2(n10415), .C1(
        P2_U3088), .C2(n10410), .ZN(P2_U3325) );
  OAI222_X1 U12317 ( .A1(n14787), .A2(n10412), .B1(n14783), .B2(n10413), .C1(
        P2_U3088), .C2(n10498), .ZN(P2_U3326) );
  OAI222_X1 U12318 ( .A1(n15777), .A2(n10414), .B1(n15780), .B2(n10413), .C1(
        P1_U3086), .C2(n15336), .ZN(P1_U3354) );
  OAI222_X1 U12319 ( .A1(n15777), .A2(n10416), .B1(n15780), .B2(n10415), .C1(
        P1_U3086), .C2(n15354), .ZN(P1_U3353) );
  INV_X1 U12320 ( .A(n10417), .ZN(n10424) );
  INV_X1 U12321 ( .A(n15777), .ZN(n15763) );
  AOI22_X1 U12322 ( .A1(n16288), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n15763), .ZN(n10418) );
  OAI21_X1 U12323 ( .B1(n10424), .B2(n15780), .A(n10418), .ZN(P1_U3351) );
  NAND2_X1 U12324 ( .A1(n8156), .A2(P3_U3151), .ZN(n13853) );
  MUX2_X1 U12325 ( .A(n10420), .B(n13005), .S(P3_STATE_REG_SCAN_IN), .Z(n10421) );
  OAI21_X1 U12326 ( .B1(n10422), .B2(n13853), .A(n10421), .ZN(P3_U3295) );
  INV_X1 U12327 ( .A(n14401), .ZN(n10423) );
  OAI222_X1 U12328 ( .A1(n14787), .A2(n7760), .B1(n14783), .B2(n10424), .C1(
        P2_U3088), .C2(n10423), .ZN(P2_U3323) );
  INV_X1 U12329 ( .A(n13853), .ZN(n11550) );
  INV_X1 U12330 ( .A(n13850), .ZN(n13846) );
  AOI222_X1 U12331 ( .A1(n10425), .A2(n11550), .B1(n7767), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_3_), .C2(n13846), .ZN(n10426) );
  INV_X1 U12332 ( .A(n10426), .ZN(P3_U3292) );
  INV_X1 U12333 ( .A(n11526), .ZN(n11534) );
  AOI222_X1 U12334 ( .A1(n10427), .A2(n11550), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11534), .C1(SI_7_), .C2(n13846), .ZN(n10428) );
  INV_X1 U12335 ( .A(n10428), .ZN(P3_U3288) );
  INV_X1 U12336 ( .A(n11113), .ZN(n11097) );
  AOI222_X1 U12337 ( .A1(n10429), .A2(n11550), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11097), .C1(SI_4_), .C2(n13846), .ZN(n10430) );
  INV_X1 U12338 ( .A(n10430), .ZN(P3_U3291) );
  INV_X1 U12339 ( .A(n11246), .ZN(n11251) );
  AOI222_X1 U12340 ( .A1(n10431), .A2(n11550), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11251), .C1(SI_5_), .C2(n13846), .ZN(n10432) );
  INV_X1 U12341 ( .A(n10432), .ZN(P3_U3290) );
  AOI222_X1 U12342 ( .A1(n10433), .A2(n11550), .B1(n7779), .B2(
        P3_STATE_REG_SCAN_IN), .C1(n13846), .C2(SI_2_), .ZN(n10434) );
  INV_X1 U12343 ( .A(n10434), .ZN(P3_U3293) );
  AOI222_X1 U12344 ( .A1(n10435), .A2(n11550), .B1(SI_10_), .B2(n13846), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n11834), .ZN(n10436) );
  INV_X1 U12345 ( .A(n10436), .ZN(P3_U3285) );
  OAI222_X1 U12346 ( .A1(n11667), .A2(P3_U3151), .B1(n13853), .B2(n10438), 
        .C1(n10437), .C2(n13850), .ZN(P3_U3287) );
  OAI222_X1 U12347 ( .A1(n16143), .A2(P3_U3151), .B1(n13853), .B2(n10440), 
        .C1(n10439), .C2(n13850), .ZN(P3_U3289) );
  AOI222_X1 U12348 ( .A1(n10441), .A2(n11550), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11817), .C1(SI_9_), .C2(n13846), .ZN(n10442) );
  INV_X1 U12349 ( .A(n10442), .ZN(P3_U3286) );
  INV_X1 U12350 ( .A(n10443), .ZN(n10445) );
  INV_X1 U12351 ( .A(n10503), .ZN(n10532) );
  OAI222_X1 U12352 ( .A1(n14787), .A2(n10444), .B1(n14783), .B2(n10445), .C1(
        P2_U3088), .C2(n10532), .ZN(P2_U3322) );
  INV_X1 U12353 ( .A(n10599), .ZN(n10631) );
  OAI222_X1 U12354 ( .A1(n15777), .A2(n10446), .B1(n15780), .B2(n10445), .C1(
        P1_U3086), .C2(n10631), .ZN(P1_U3350) );
  INV_X1 U12355 ( .A(n10447), .ZN(n10449) );
  INV_X1 U12356 ( .A(n10504), .ZN(n15841) );
  OAI222_X1 U12357 ( .A1(n14787), .A2(n10448), .B1(n14783), .B2(n10449), .C1(
        P2_U3088), .C2(n15841), .ZN(P2_U3321) );
  INV_X1 U12358 ( .A(n10601), .ZN(n10868) );
  OAI222_X1 U12359 ( .A1(n15777), .A2(n10450), .B1(n15780), .B2(n10449), .C1(
        P1_U3086), .C2(n10868), .ZN(P1_U3349) );
  OAI222_X1 U12360 ( .A1(n16166), .A2(P3_U3151), .B1(n13853), .B2(n10451), 
        .C1(n13436), .C2(n13850), .ZN(P3_U3283) );
  INV_X1 U12361 ( .A(n13047), .ZN(n16152) );
  AOI222_X1 U12362 ( .A1(n10452), .A2(n11550), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n16152), .C1(SI_11_), .C2(n13846), .ZN(n10453) );
  INV_X1 U12363 ( .A(n10453), .ZN(P3_U3284) );
  NAND2_X1 U12364 ( .A1(n13838), .A2(P3_D_REG_0__SCAN_IN), .ZN(n10454) );
  OAI21_X1 U12365 ( .B1(n10945), .B2(n13838), .A(n10454), .ZN(P3_U3376) );
  INV_X1 U12366 ( .A(n10455), .ZN(n10457) );
  INV_X1 U12367 ( .A(n15385), .ZN(n10572) );
  OAI222_X1 U12368 ( .A1(n15777), .A2(n10456), .B1(n15780), .B2(n10457), .C1(
        P1_U3086), .C2(n10572), .ZN(P1_U3348) );
  INV_X1 U12369 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10458) );
  INV_X1 U12370 ( .A(n10507), .ZN(n10647) );
  OAI222_X1 U12371 ( .A1(n14787), .A2(n10458), .B1(n14783), .B2(n10457), .C1(
        P2_U3088), .C2(n10647), .ZN(P2_U3320) );
  INV_X1 U12372 ( .A(n10459), .ZN(n10462) );
  INV_X1 U12373 ( .A(n10508), .ZN(n10562) );
  OAI222_X1 U12374 ( .A1(n14787), .A2(n10460), .B1(n14783), .B2(n10462), .C1(
        P2_U3088), .C2(n10562), .ZN(P2_U3319) );
  INV_X1 U12375 ( .A(n10660), .ZN(n10461) );
  OAI222_X1 U12376 ( .A1(n15777), .A2(n10463), .B1(n15780), .B2(n10462), .C1(
        P1_U3086), .C2(n10461), .ZN(P1_U3347) );
  OAI222_X1 U12377 ( .A1(n13853), .A2(n10464), .B1(n13850), .B2(n13629), .C1(
        n13052), .C2(P3_U3151), .ZN(P3_U3282) );
  OAI222_X1 U12378 ( .A1(n13853), .A2(n10466), .B1(n13850), .B2(n10465), .C1(
        n16204), .C2(P3_U3151), .ZN(P3_U3281) );
  INV_X1 U12379 ( .A(n10469), .ZN(n10467) );
  AND2_X2 U12380 ( .A1(n10468), .A2(n11572), .ZN(n15816) );
  OAI22_X1 U12381 ( .A1(n15816), .A2(P1_D_REG_1__SCAN_IN), .B1(n10470), .B2(
        n10469), .ZN(n10471) );
  INV_X1 U12382 ( .A(n10471), .ZN(P1_U3446) );
  INV_X1 U12383 ( .A(n10472), .ZN(n10474) );
  INV_X1 U12384 ( .A(n10676), .ZN(n10495) );
  OAI222_X1 U12385 ( .A1(n14787), .A2(n10473), .B1(n14783), .B2(n10474), .C1(
        P2_U3088), .C2(n10495), .ZN(P2_U3318) );
  INV_X1 U12386 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10475) );
  INV_X1 U12387 ( .A(n10606), .ZN(n10696) );
  OAI222_X1 U12388 ( .A1(n15777), .A2(n10475), .B1(n15780), .B2(n10474), .C1(
        P1_U3086), .C2(n10696), .ZN(P1_U3346) );
  OAI222_X1 U12389 ( .A1(n13853), .A2(n10476), .B1(n13850), .B2(n13428), .C1(
        n13055), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U12390 ( .A(n10477), .ZN(n10479) );
  AOI22_X1 U12391 ( .A1(n10759), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n15763), .ZN(n10478) );
  OAI21_X1 U12392 ( .B1(n10479), .B2(n15780), .A(n10478), .ZN(P1_U3345) );
  INV_X1 U12393 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10480) );
  INV_X1 U12394 ( .A(n10706), .ZN(n10714) );
  OAI222_X1 U12395 ( .A1(n14787), .A2(n10480), .B1(n14783), .B2(n10479), .C1(
        P2_U3088), .C2(n10714), .ZN(P2_U3317) );
  MUX2_X1 U12396 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n11370), .S(n10498), .Z(
        n14369) );
  NAND2_X1 U12397 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n14370) );
  OR2_X1 U12398 ( .A1(n14369), .A2(n14370), .ZN(n14381) );
  INV_X1 U12399 ( .A(n10498), .ZN(n14372) );
  NAND2_X1 U12400 ( .A1(n14372), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n14380) );
  MUX2_X1 U12401 ( .A(n11353), .B(P2_REG2_REG_2__SCAN_IN), .S(n14385), .Z(
        n14379) );
  AOI21_X1 U12402 ( .B1(n14381), .B2(n14380), .A(n14379), .ZN(n14383) );
  AOI21_X1 U12403 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n14385), .A(n14383), .ZN(
        n15828) );
  MUX2_X1 U12404 ( .A(n10481), .B(P2_REG2_REG_3__SCAN_IN), .S(n10499), .Z(
        n15827) );
  NOR2_X1 U12405 ( .A1(n15828), .A2(n15827), .ZN(n15826) );
  NOR2_X1 U12406 ( .A1(n15824), .A2(n10481), .ZN(n14397) );
  MUX2_X1 U12407 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11360), .S(n14401), .Z(
        n14396) );
  OAI21_X1 U12408 ( .B1(n15826), .B2(n14397), .A(n14396), .ZN(n14395) );
  NAND2_X1 U12409 ( .A1(n14401), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10527) );
  MUX2_X1 U12410 ( .A(n8631), .B(P2_REG2_REG_5__SCAN_IN), .S(n10503), .Z(
        n10526) );
  AOI21_X1 U12411 ( .B1(n14395), .B2(n10527), .A(n10526), .ZN(n10525) );
  AOI21_X1 U12412 ( .B1(n10503), .B2(P2_REG2_REG_5__SCAN_IN), .A(n10525), .ZN(
        n15851) );
  INV_X1 U12413 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10482) );
  MUX2_X1 U12414 ( .A(n10482), .B(P2_REG2_REG_6__SCAN_IN), .S(n10504), .Z(
        n15850) );
  NOR2_X1 U12415 ( .A1(n15851), .A2(n15850), .ZN(n15849) );
  AND2_X1 U12416 ( .A1(n10504), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10641) );
  MUX2_X1 U12417 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10483), .S(n10507), .Z(
        n10640) );
  OAI21_X1 U12418 ( .B1(n15849), .B2(n10641), .A(n10640), .ZN(n10639) );
  NAND2_X1 U12419 ( .A1(n10507), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10557) );
  MUX2_X1 U12420 ( .A(n11386), .B(P2_REG2_REG_8__SCAN_IN), .S(n10508), .Z(
        n10556) );
  AOI21_X1 U12421 ( .B1(n10639), .B2(n10557), .A(n10556), .ZN(n10555) );
  AOI21_X1 U12422 ( .B1(n10508), .B2(P2_REG2_REG_8__SCAN_IN), .A(n10555), .ZN(
        n10485) );
  MUX2_X1 U12423 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n14626), .S(n10676), .Z(
        n10484) );
  NAND2_X1 U12424 ( .A1(n10485), .A2(n10484), .ZN(n10671) );
  OAI21_X1 U12425 ( .B1(n10485), .B2(n10484), .A(n10671), .ZN(n10497) );
  INV_X1 U12426 ( .A(n10486), .ZN(n12150) );
  OR2_X1 U12427 ( .A1(n10618), .A2(n12150), .ZN(n10491) );
  NAND2_X1 U12428 ( .A1(n10487), .A2(n10486), .ZN(n10489) );
  NAND2_X1 U12429 ( .A1(n10489), .A2(n10488), .ZN(n10490) );
  NOR2_X1 U12430 ( .A1(n9149), .A2(P2_U3088), .ZN(n14779) );
  INV_X1 U12431 ( .A(n14782), .ZN(n14325) );
  NAND2_X1 U12432 ( .A1(n10492), .A2(n9149), .ZN(n15869) );
  NAND2_X1 U12433 ( .A1(n15875), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n10494) );
  NAND2_X1 U12434 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n11228) );
  OAI211_X1 U12435 ( .C1(n15842), .C2(n10495), .A(n10494), .B(n11228), .ZN(
        n10496) );
  AOI21_X1 U12436 ( .B1(n10497), .B2(n15877), .A(n10496), .ZN(n10515) );
  MUX2_X1 U12437 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n8564), .S(n10498), .Z(
        n14373) );
  OR3_X1 U12438 ( .A1(n14373), .A2(n10534), .A3(n14374), .ZN(n14389) );
  NAND2_X1 U12439 ( .A1(n14372), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n14388) );
  MUX2_X1 U12440 ( .A(n8576), .B(P2_REG1_REG_2__SCAN_IN), .S(n14385), .Z(
        n14387) );
  AOI21_X1 U12441 ( .B1(n14389), .B2(n14388), .A(n14387), .ZN(n14386) );
  AOI21_X1 U12442 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n14385), .A(n14386), .ZN(
        n15833) );
  MUX2_X1 U12443 ( .A(n10500), .B(P2_REG1_REG_3__SCAN_IN), .S(n10499), .Z(
        n15832) );
  NOR2_X1 U12444 ( .A1(n15833), .A2(n15832), .ZN(n15831) );
  NOR2_X1 U12445 ( .A1(n15824), .A2(n10500), .ZN(n14402) );
  MUX2_X1 U12446 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10501), .S(n14401), .Z(
        n10502) );
  OAI21_X1 U12447 ( .B1(n15831), .B2(n14402), .A(n10502), .ZN(n14405) );
  NAND2_X1 U12448 ( .A1(n14401), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10520) );
  MUX2_X1 U12449 ( .A(n8636), .B(P2_REG1_REG_5__SCAN_IN), .S(n10503), .Z(
        n10519) );
  AOI21_X1 U12450 ( .B1(n14405), .B2(n10520), .A(n10519), .ZN(n10522) );
  AOI21_X1 U12451 ( .B1(n10503), .B2(P2_REG1_REG_5__SCAN_IN), .A(n10522), .ZN(
        n15845) );
  MUX2_X1 U12452 ( .A(n10505), .B(P2_REG1_REG_6__SCAN_IN), .S(n10504), .Z(
        n15844) );
  OR2_X1 U12453 ( .A1(n15845), .A2(n15844), .ZN(n15847) );
  OAI21_X1 U12454 ( .B1(n10505), .B2(n15841), .A(n15847), .ZN(n10637) );
  MUX2_X1 U12455 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10506), .S(n10507), .Z(
        n10636) );
  NAND2_X1 U12456 ( .A1(n10637), .A2(n10636), .ZN(n10635) );
  NAND2_X1 U12457 ( .A1(n10507), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10551) );
  MUX2_X1 U12458 ( .A(n8694), .B(P2_REG1_REG_8__SCAN_IN), .S(n10508), .Z(
        n10550) );
  AOI21_X1 U12459 ( .B1(n10635), .B2(n10551), .A(n10550), .ZN(n10553) );
  AOI21_X1 U12460 ( .B1(n10508), .B2(P2_REG1_REG_8__SCAN_IN), .A(n10553), .ZN(
        n10510) );
  MUX2_X1 U12461 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n8712), .S(n10676), .Z(
        n10509) );
  NAND2_X1 U12462 ( .A1(n10510), .A2(n10509), .ZN(n10675) );
  OAI21_X1 U12463 ( .B1(n10510), .B2(n10509), .A(n10675), .ZN(n10513) );
  INV_X1 U12464 ( .A(n10511), .ZN(n10512) );
  OR2_X1 U12465 ( .A1(n10512), .A2(n14325), .ZN(n15830) );
  NAND2_X1 U12466 ( .A1(n10513), .A2(n15873), .ZN(n10514) );
  NAND2_X1 U12467 ( .A1(n10515), .A2(n10514), .ZN(P2_U3223) );
  INV_X1 U12468 ( .A(n10516), .ZN(n10518) );
  INV_X1 U12469 ( .A(n16250), .ZN(n13058) );
  OAI222_X1 U12470 ( .A1(n13853), .A2(n10518), .B1(n13850), .B2(n10517), .C1(
        n13058), .C2(P3_U3151), .ZN(P3_U3279) );
  NAND2_X1 U12471 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10963) );
  INV_X1 U12472 ( .A(n10963), .ZN(n10524) );
  AND3_X1 U12473 ( .A1(n14405), .A2(n10520), .A3(n10519), .ZN(n10521) );
  NOR3_X1 U12474 ( .A1(n15830), .A2(n10522), .A3(n10521), .ZN(n10523) );
  AOI211_X1 U12475 ( .C1(n15875), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n10524), .B(
        n10523), .ZN(n10531) );
  INV_X1 U12476 ( .A(n10525), .ZN(n10529) );
  NAND3_X1 U12477 ( .A1(n14395), .A2(n10527), .A3(n10526), .ZN(n10528) );
  NAND3_X1 U12478 ( .A1(n15877), .A2(n10529), .A3(n10528), .ZN(n10530) );
  OAI211_X1 U12479 ( .C1(n15842), .C2(n10532), .A(n10531), .B(n10530), .ZN(
        P2_U3219) );
  NAND2_X1 U12480 ( .A1(n15877), .A2(n10940), .ZN(n10533) );
  OAI211_X1 U12481 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15830), .A(n10533), .B(
        n15842), .ZN(n10536) );
  OAI22_X1 U12482 ( .A1(n15848), .A2(n10940), .B1(n10534), .B2(n15830), .ZN(
        n10535) );
  MUX2_X1 U12483 ( .A(n10536), .B(n10535), .S(n14374), .Z(n10540) );
  INV_X1 U12484 ( .A(n15875), .ZN(n10538) );
  INV_X1 U12485 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10537) );
  OAI22_X1 U12486 ( .A1(n10538), .A2(n10537), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10937), .ZN(n10539) );
  OR2_X1 U12487 ( .A1(n10540), .A2(n10539), .ZN(P2_U3214) );
  INV_X1 U12488 ( .A(n10541), .ZN(n10544) );
  INV_X1 U12489 ( .A(n10728), .ZN(n10542) );
  OAI222_X1 U12490 ( .A1(n15777), .A2(n10543), .B1(n15780), .B2(n10544), .C1(
        P1_U3086), .C2(n10542), .ZN(P1_U3344) );
  INV_X1 U12491 ( .A(n10837), .ZN(n10713) );
  OAI222_X1 U12492 ( .A1(n14787), .A2(n10545), .B1(n14783), .B2(n10544), .C1(
        P2_U3088), .C2(n10713), .ZN(P2_U3316) );
  INV_X1 U12493 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n10547) );
  NAND2_X1 U12494 ( .A1(n12958), .A2(P3_U3897), .ZN(n10546) );
  OAI21_X1 U12495 ( .B1(P3_U3897), .B2(n10547), .A(n10546), .ZN(P3_U3508) );
  OAI222_X1 U12496 ( .A1(n13853), .A2(n10549), .B1(n13850), .B2(n10548), .C1(
        n13039), .C2(P3_U3151), .ZN(P3_U3278) );
  AND2_X1 U12497 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n11148) );
  AND3_X1 U12498 ( .A1(n10635), .A2(n10551), .A3(n10550), .ZN(n10552) );
  NOR3_X1 U12499 ( .A1(n10553), .A2(n10552), .A3(n15830), .ZN(n10554) );
  AOI211_X1 U12500 ( .C1(n15875), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n11148), .B(
        n10554), .ZN(n10561) );
  INV_X1 U12501 ( .A(n10555), .ZN(n10559) );
  NAND3_X1 U12502 ( .A1(n10639), .A2(n10557), .A3(n10556), .ZN(n10558) );
  NAND3_X1 U12503 ( .A1(n10559), .A2(n15877), .A3(n10558), .ZN(n10560) );
  OAI211_X1 U12504 ( .C1(n15842), .C2(n10562), .A(n10561), .B(n10560), .ZN(
        P2_U3222) );
  INV_X1 U12505 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n10564) );
  NAND2_X1 U12506 ( .A1(n12903), .A2(P3_U3897), .ZN(n10563) );
  OAI21_X1 U12507 ( .B1(P3_U3897), .B2(n10564), .A(n10563), .ZN(P3_U3506) );
  INV_X1 U12508 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n10566) );
  NAND2_X1 U12509 ( .A1(n12640), .A2(P3_U3897), .ZN(n10565) );
  OAI21_X1 U12510 ( .B1(P3_U3897), .B2(n10566), .A(n10565), .ZN(P3_U3501) );
  MUX2_X1 U12511 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9255), .S(n15336), .Z(
        n10567) );
  AOI21_X1 U12512 ( .B1(n15335), .B2(P1_REG2_REG_1__SCAN_IN), .A(n15328), .ZN(
        n15356) );
  MUX2_X1 U12513 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n15355), .S(n15354), .Z(
        n10568) );
  OR2_X1 U12514 ( .A1(n15356), .A2(n10568), .ZN(n15371) );
  NAND2_X1 U12515 ( .A1(n15351), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n15370) );
  INV_X1 U12516 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10569) );
  MUX2_X1 U12517 ( .A(n10569), .B(P1_REG2_REG_3__SCAN_IN), .S(n15364), .Z(
        n15369) );
  NOR2_X1 U12518 ( .A1(n15362), .A2(n10569), .ZN(n16281) );
  MUX2_X1 U12519 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10570), .S(n16288), .Z(
        n16280) );
  OAI21_X1 U12520 ( .B1(n16282), .B2(n16281), .A(n16280), .ZN(n16279) );
  NAND2_X1 U12521 ( .A1(n16288), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10623) );
  MUX2_X1 U12522 ( .A(n9306), .B(P1_REG2_REG_5__SCAN_IN), .S(n10599), .Z(
        n10622) );
  AOI21_X1 U12523 ( .B1(n10599), .B2(P1_REG2_REG_5__SCAN_IN), .A(n10625), .ZN(
        n10859) );
  INV_X1 U12524 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10571) );
  MUX2_X1 U12525 ( .A(n10571), .B(P1_REG2_REG_6__SCAN_IN), .S(n10601), .Z(
        n10858) );
  NAND2_X1 U12526 ( .A1(n10601), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n15381) );
  MUX2_X1 U12527 ( .A(n9339), .B(P1_REG2_REG_7__SCAN_IN), .S(n15385), .Z(
        n15380) );
  NOR2_X1 U12528 ( .A1(n10572), .A2(n9339), .ZN(n10664) );
  MUX2_X1 U12529 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10573), .S(n10660), .Z(
        n10663) );
  OAI21_X1 U12530 ( .B1(n15379), .B2(n10664), .A(n10663), .ZN(n10686) );
  NAND2_X1 U12531 ( .A1(n10660), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10685) );
  MUX2_X1 U12532 ( .A(n9368), .B(P1_REG2_REG_9__SCAN_IN), .S(n10606), .Z(
        n10684) );
  AOI21_X1 U12533 ( .B1(n10686), .B2(n10685), .A(n10684), .ZN(n10688) );
  AOI21_X1 U12534 ( .B1(n10606), .B2(P1_REG2_REG_9__SCAN_IN), .A(n10688), .ZN(
        n10765) );
  MUX2_X1 U12535 ( .A(n12072), .B(P1_REG2_REG_10__SCAN_IN), .S(n10759), .Z(
        n10764) );
  NAND2_X1 U12536 ( .A1(n10759), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10575) );
  MUX2_X1 U12537 ( .A(n9399), .B(P1_REG2_REG_11__SCAN_IN), .S(n10728), .Z(
        n10574) );
  NAND3_X1 U12538 ( .A1(n10766), .A2(n10575), .A3(n10574), .ZN(n10582) );
  INV_X1 U12539 ( .A(n10578), .ZN(n10576) );
  NAND2_X1 U12540 ( .A1(n10576), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15297) );
  INV_X1 U12541 ( .A(n15297), .ZN(n12118) );
  AOI21_X1 U12542 ( .B1(n10579), .B2(n10578), .A(n10577), .ZN(n10583) );
  NAND2_X1 U12543 ( .A1(n10585), .A2(n10583), .ZN(n15895) );
  INV_X1 U12544 ( .A(n15895), .ZN(n10581) );
  NOR2_X1 U12545 ( .A1(n15772), .A2(n15885), .ZN(n10580) );
  NAND2_X1 U12546 ( .A1(n10581), .A2(n10580), .ZN(n16285) );
  NAND2_X1 U12547 ( .A1(n10582), .A2(n15415), .ZN(n10615) );
  NOR2_X1 U12548 ( .A1(n15895), .A2(n15347), .ZN(n16287) );
  INV_X1 U12549 ( .A(n10583), .ZN(n10584) );
  NAND2_X1 U12550 ( .A1(n10585), .A2(n10584), .ZN(n16301) );
  INV_X1 U12551 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n16032) );
  NAND2_X1 U12552 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n12256)
         );
  OAI21_X1 U12553 ( .B1(n16301), .B2(n16032), .A(n12256), .ZN(n10586) );
  AOI21_X1 U12554 ( .B1(n16287), .B2(n10728), .A(n10586), .ZN(n10614) );
  MUX2_X1 U12555 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9403), .S(n10728), .Z(
        n10611) );
  INV_X1 U12556 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10587) );
  MUX2_X1 U12557 ( .A(n10587), .B(P1_REG1_REG_1__SCAN_IN), .S(n15336), .Z(
        n10589) );
  AND2_X1 U12558 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10588) );
  NAND2_X1 U12559 ( .A1(n10589), .A2(n10588), .ZN(n15339) );
  NAND2_X1 U12560 ( .A1(n15335), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10590) );
  NAND2_X1 U12561 ( .A1(n15339), .A2(n10590), .ZN(n15352) );
  MUX2_X1 U12562 ( .A(n10591), .B(P1_REG1_REG_2__SCAN_IN), .S(n15354), .Z(
        n15353) );
  NAND2_X1 U12563 ( .A1(n15352), .A2(n15353), .ZN(n15366) );
  NAND2_X1 U12564 ( .A1(n15351), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n15365) );
  NAND2_X1 U12565 ( .A1(n15366), .A2(n15365), .ZN(n10594) );
  MUX2_X1 U12566 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10592), .S(n15364), .Z(
        n10593) );
  NAND2_X1 U12567 ( .A1(n10594), .A2(n10593), .ZN(n16291) );
  NAND2_X1 U12568 ( .A1(n15364), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n16290) );
  NAND2_X1 U12569 ( .A1(n16291), .A2(n16290), .ZN(n10597) );
  MUX2_X1 U12570 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10595), .S(n16288), .Z(
        n10596) );
  NAND2_X1 U12571 ( .A1(n10597), .A2(n10596), .ZN(n16293) );
  NAND2_X1 U12572 ( .A1(n16288), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10598) );
  AND2_X1 U12573 ( .A1(n16293), .A2(n10598), .ZN(n10620) );
  MUX2_X1 U12574 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9312), .S(n10599), .Z(
        n10621) );
  NAND2_X1 U12575 ( .A1(n10620), .A2(n10621), .ZN(n10619) );
  OR2_X1 U12576 ( .A1(n10599), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10600) );
  NAND2_X1 U12577 ( .A1(n10619), .A2(n10600), .ZN(n10864) );
  MUX2_X1 U12578 ( .A(n9323), .B(P1_REG1_REG_6__SCAN_IN), .S(n10601), .Z(
        n10863) );
  OR2_X1 U12579 ( .A1(n10864), .A2(n10863), .ZN(n15388) );
  NAND2_X1 U12580 ( .A1(n10601), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n15387) );
  NAND2_X1 U12581 ( .A1(n15388), .A2(n15387), .ZN(n10604) );
  MUX2_X1 U12582 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10602), .S(n15385), .Z(
        n10603) );
  NAND2_X1 U12583 ( .A1(n10604), .A2(n10603), .ZN(n15390) );
  NAND2_X1 U12584 ( .A1(n15385), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10605) );
  AND2_X1 U12585 ( .A1(n15390), .A2(n10605), .ZN(n10658) );
  MUX2_X1 U12586 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9354), .S(n10660), .Z(
        n10659) );
  NAND2_X1 U12587 ( .A1(n10658), .A2(n10659), .ZN(n10692) );
  OR2_X1 U12588 ( .A1(n10660), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10690) );
  NAND2_X1 U12589 ( .A1(n10692), .A2(n10690), .ZN(n10607) );
  MUX2_X1 U12590 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9373), .S(n10606), .Z(
        n10689) );
  NAND2_X1 U12591 ( .A1(n10607), .A2(n10689), .ZN(n10694) );
  NAND2_X1 U12592 ( .A1(n10696), .A2(n9373), .ZN(n10608) );
  NAND2_X1 U12593 ( .A1(n10694), .A2(n10608), .ZN(n10761) );
  MUX2_X1 U12594 ( .A(n9387), .B(P1_REG1_REG_10__SCAN_IN), .S(n10759), .Z(
        n10760) );
  OR2_X1 U12595 ( .A1(n10761), .A2(n10760), .ZN(n10762) );
  NAND2_X1 U12596 ( .A1(n10759), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10609) );
  AND2_X1 U12597 ( .A1(n10762), .A2(n10609), .ZN(n10610) );
  NAND2_X1 U12598 ( .A1(n10610), .A2(n10611), .ZN(n10733) );
  OAI21_X1 U12599 ( .B1(n10611), .B2(n10610), .A(n10733), .ZN(n10612) );
  INV_X1 U12600 ( .A(n15885), .ZN(n15345) );
  NAND2_X1 U12601 ( .A1(n10612), .A2(n16294), .ZN(n10613) );
  OAI211_X1 U12602 ( .C1(n10725), .C2(n10615), .A(n10614), .B(n10613), .ZN(
        P1_U3254) );
  INV_X1 U12603 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n10617) );
  NAND2_X1 U12604 ( .A1(n12452), .A2(P3_U3897), .ZN(n10616) );
  OAI21_X1 U12605 ( .B1(P3_U3897), .B2(n10617), .A(n10616), .ZN(P3_U3503) );
  OR3_X2 U12606 ( .A1(n10618), .A2(n12150), .A3(P2_U3088), .ZN(n14367) );
  INV_X1 U12607 ( .A(n14367), .ZN(P2_U3947) );
  OAI21_X1 U12608 ( .B1(n10621), .B2(n10620), .A(n10619), .ZN(n10627) );
  AND3_X1 U12609 ( .A1(n16279), .A2(n10623), .A3(n10622), .ZN(n10624) );
  NOR3_X1 U12610 ( .A1(n16285), .A2(n10625), .A3(n10624), .ZN(n10626) );
  AOI21_X1 U12611 ( .B1(n16294), .B2(n10627), .A(n10626), .ZN(n10630) );
  INV_X1 U12612 ( .A(n16301), .ZN(n15892) );
  AND2_X1 U12613 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10628) );
  AOI21_X1 U12614 ( .B1(n15892), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10628), .ZN(
        n10629) );
  OAI211_X1 U12615 ( .C1(n10631), .C2(n15928), .A(n10630), .B(n10629), .ZN(
        P1_U3248) );
  INV_X1 U12616 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n10634) );
  NAND2_X1 U12617 ( .A1(n10632), .A2(P3_U3897), .ZN(n10633) );
  OAI21_X1 U12618 ( .B1(P3_U3897), .B2(n10634), .A(n10633), .ZN(P3_U3496) );
  NAND2_X1 U12619 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n11305) );
  OAI211_X1 U12620 ( .C1(n10637), .C2(n10636), .A(n15873), .B(n10635), .ZN(
        n10638) );
  NAND2_X1 U12621 ( .A1(n11305), .A2(n10638), .ZN(n10645) );
  INV_X1 U12622 ( .A(n10639), .ZN(n10643) );
  NOR3_X1 U12623 ( .A1(n15849), .A2(n10641), .A3(n10640), .ZN(n10642) );
  NOR3_X1 U12624 ( .A1(n10643), .A2(n10642), .A3(n15848), .ZN(n10644) );
  AOI211_X1 U12625 ( .C1(n15875), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n10645), .B(
        n10644), .ZN(n10646) );
  OAI21_X1 U12626 ( .B1(n10647), .B2(n15842), .A(n10646), .ZN(P2_U3221) );
  INV_X1 U12627 ( .A(n13988), .ZN(n13972) );
  OAI22_X1 U12628 ( .A1(n10786), .A2(n13967), .B1(n10648), .B2(n13968), .ZN(
        n10744) );
  OR2_X1 U12629 ( .A1(n10649), .A2(P2_U3088), .ZN(n10846) );
  AOI22_X1 U12630 ( .A1(n13972), .A2(n10744), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n10846), .ZN(n10653) );
  OAI21_X1 U12631 ( .B1(n7492), .B2(n10650), .A(n10852), .ZN(n10651) );
  NAND2_X1 U12632 ( .A1(n13990), .A2(n10651), .ZN(n10652) );
  OAI211_X1 U12633 ( .C1(n11365), .C2(n13975), .A(n10653), .B(n10652), .ZN(
        P2_U3194) );
  INV_X1 U12634 ( .A(n10654), .ZN(n10700) );
  AOI22_X1 U12635 ( .A1(n10914), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n15763), .ZN(n10655) );
  OAI21_X1 U12636 ( .B1(n10700), .B2(n15780), .A(n10655), .ZN(P1_U3343) );
  INV_X1 U12637 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n10657) );
  NAND2_X1 U12638 ( .A1(n12945), .A2(P3_U3897), .ZN(n10656) );
  OAI21_X1 U12639 ( .B1(P3_U3897), .B2(n10657), .A(n10656), .ZN(P3_U3512) );
  OAI21_X1 U12640 ( .B1(n10659), .B2(n10658), .A(n10692), .ZN(n10669) );
  INV_X1 U12641 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10662) );
  NAND2_X1 U12642 ( .A1(n16287), .A2(n10660), .ZN(n10661) );
  NAND2_X1 U12643 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11798) );
  OAI211_X1 U12644 ( .C1(n10662), .C2(n16301), .A(n10661), .B(n11798), .ZN(
        n10668) );
  INV_X1 U12645 ( .A(n10686), .ZN(n10666) );
  NOR3_X1 U12646 ( .A1(n15379), .A2(n10664), .A3(n10663), .ZN(n10665) );
  NOR3_X1 U12647 ( .A1(n10666), .A2(n10665), .A3(n16285), .ZN(n10667) );
  AOI211_X1 U12648 ( .C1(n16294), .C2(n10669), .A(n10668), .B(n10667), .ZN(
        n10670) );
  INV_X1 U12649 ( .A(n10670), .ZN(P1_U3251) );
  OAI21_X1 U12650 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n10676), .A(n10671), .ZN(
        n10673) );
  MUX2_X1 U12651 ( .A(n11638), .B(P2_REG2_REG_10__SCAN_IN), .S(n10706), .Z(
        n10672) );
  NOR2_X1 U12652 ( .A1(n10673), .A2(n10672), .ZN(n10705) );
  AOI211_X1 U12653 ( .C1(n10673), .C2(n10672), .A(n15848), .B(n10705), .ZN(
        n10674) );
  INV_X1 U12654 ( .A(n10674), .ZN(n10683) );
  NAND2_X1 U12655 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11395)
         );
  MUX2_X1 U12656 ( .A(n8733), .B(P2_REG1_REG_10__SCAN_IN), .S(n10706), .Z(
        n10678) );
  OAI21_X1 U12657 ( .B1(n10676), .B2(P2_REG1_REG_9__SCAN_IN), .A(n10675), .ZN(
        n10677) );
  NOR2_X1 U12658 ( .A1(n10677), .A2(n10678), .ZN(n10718) );
  AOI211_X1 U12659 ( .C1(n10678), .C2(n10677), .A(n10718), .B(n15830), .ZN(
        n10679) );
  INV_X1 U12660 ( .A(n10679), .ZN(n10680) );
  NAND2_X1 U12661 ( .A1(n11395), .A2(n10680), .ZN(n10681) );
  AOI21_X1 U12662 ( .B1(n15875), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10681), 
        .ZN(n10682) );
  OAI211_X1 U12663 ( .C1(n15842), .C2(n10714), .A(n10683), .B(n10682), .ZN(
        P2_U3224) );
  AND3_X1 U12664 ( .A1(n10686), .A2(n10685), .A3(n10684), .ZN(n10687) );
  NOR3_X1 U12665 ( .A1(n10688), .A2(n10687), .A3(n16285), .ZN(n10699) );
  INV_X1 U12666 ( .A(n10689), .ZN(n10691) );
  NAND3_X1 U12667 ( .A1(n10692), .A2(n10691), .A3(n10690), .ZN(n10693) );
  INV_X1 U12668 ( .A(n16294), .ZN(n15925) );
  AOI21_X1 U12669 ( .B1(n10694), .B2(n10693), .A(n15925), .ZN(n10698) );
  NAND2_X1 U12670 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n12214) );
  NAND2_X1 U12671 ( .A1(n15892), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n10695) );
  OAI211_X1 U12672 ( .C1(n15928), .C2(n10696), .A(n12214), .B(n10695), .ZN(
        n10697) );
  OR3_X1 U12673 ( .A1(n10699), .A2(n10698), .A3(n10697), .ZN(P1_U3252) );
  INV_X1 U12674 ( .A(n11072), .ZN(n10833) );
  OAI222_X1 U12675 ( .A1(n14787), .A2(n10701), .B1(n14783), .B2(n10700), .C1(
        n10833), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U12676 ( .A(n10702), .ZN(n10704) );
  INV_X1 U12677 ( .A(n13077), .ZN(n13065) );
  OAI222_X1 U12678 ( .A1(n13853), .A2(n10704), .B1(n13850), .B2(n10703), .C1(
        n13065), .C2(P3_U3151), .ZN(P3_U3277) );
  AOI21_X1 U12679 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n10706), .A(n10705), 
        .ZN(n10709) );
  INV_X1 U12680 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10707) );
  MUX2_X1 U12681 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10707), .S(n10837), .Z(
        n10708) );
  NAND2_X1 U12682 ( .A1(n10709), .A2(n10708), .ZN(n10830) );
  OAI21_X1 U12683 ( .B1(n10709), .B2(n10708), .A(n10830), .ZN(n10723) );
  NOR2_X1 U12684 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10710), .ZN(n10711) );
  AOI21_X1 U12685 ( .B1(n15875), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n10711), 
        .ZN(n10712) );
  OAI21_X1 U12686 ( .B1(n10713), .B2(n15842), .A(n10712), .ZN(n10722) );
  NOR2_X1 U12687 ( .A1(n10714), .A2(n8733), .ZN(n10717) );
  MUX2_X1 U12688 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10715), .S(n10837), .Z(
        n10716) );
  OAI21_X1 U12689 ( .B1(n10718), .B2(n10717), .A(n10716), .ZN(n10840) );
  INV_X1 U12690 ( .A(n10840), .ZN(n10720) );
  NOR3_X1 U12691 ( .A1(n10718), .A2(n10717), .A3(n10716), .ZN(n10719) );
  NOR3_X1 U12692 ( .A1(n10720), .A2(n10719), .A3(n15830), .ZN(n10721) );
  AOI211_X1 U12693 ( .C1(n15877), .C2(n10723), .A(n10722), .B(n10721), .ZN(
        n10724) );
  INV_X1 U12694 ( .A(n10724), .ZN(P2_U3225) );
  MUX2_X1 U12695 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n9414), .S(n10914), .Z(
        n10727) );
  AOI21_X1 U12696 ( .B1(n10728), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10725), 
        .ZN(n10726) );
  NAND2_X1 U12697 ( .A1(n10726), .A2(n10727), .ZN(n10908) );
  OAI21_X1 U12698 ( .B1(n10727), .B2(n10726), .A(n10908), .ZN(n10739) );
  OR2_X1 U12699 ( .A1(n10728), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10731) );
  NAND2_X1 U12700 ( .A1(n10733), .A2(n10731), .ZN(n10729) );
  MUX2_X1 U12701 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9419), .S(n10914), .Z(
        n10730) );
  NAND2_X1 U12702 ( .A1(n10729), .A2(n10730), .ZN(n10916) );
  INV_X1 U12703 ( .A(n10730), .ZN(n10732) );
  NAND3_X1 U12704 ( .A1(n10733), .A2(n10732), .A3(n10731), .ZN(n10734) );
  AOI21_X1 U12705 ( .B1(n10916), .B2(n10734), .A(n15925), .ZN(n10738) );
  INV_X1 U12706 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n16040) );
  NAND2_X1 U12707 ( .A1(n16287), .A2(n10914), .ZN(n10736) );
  NAND2_X1 U12708 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n10735)
         );
  OAI211_X1 U12709 ( .C1(n16040), .C2(n16301), .A(n10736), .B(n10735), .ZN(
        n10737) );
  AOI211_X1 U12710 ( .C1(n10739), .C2(n15415), .A(n10738), .B(n10737), .ZN(
        n10740) );
  INV_X1 U12711 ( .A(n10740), .ZN(P1_U3255) );
  INV_X1 U12712 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10748) );
  XNOR2_X1 U12713 ( .A(n14287), .B(n10741), .ZN(n11373) );
  INV_X1 U12714 ( .A(n11346), .ZN(n10742) );
  AOI211_X1 U12715 ( .C1(n10743), .C2(n14006), .A(n7437), .B(n10742), .ZN(
        n11367) );
  AOI21_X1 U12716 ( .B1(n16382), .B2(n14006), .A(n11367), .ZN(n10746) );
  XNOR2_X1 U12717 ( .A(n14287), .B(n10819), .ZN(n10745) );
  AOI21_X1 U12718 ( .B1(n10745), .B2(n14606), .A(n10744), .ZN(n11369) );
  OAI211_X1 U12719 ( .C1(n16386), .C2(n11373), .A(n10746), .B(n11369), .ZN(
        n10898) );
  NAND2_X1 U12720 ( .A1(n11936), .A2(n10898), .ZN(n10747) );
  OAI21_X1 U12721 ( .B1(n11936), .B2(n10748), .A(n10747), .ZN(P2_U3433) );
  INV_X1 U12722 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10758) );
  XNOR2_X1 U12723 ( .A(n10749), .B(n14289), .ZN(n10751) );
  AOI21_X1 U12724 ( .B1(n10751), .B2(n14606), .A(n10750), .ZN(n11511) );
  XNOR2_X1 U12725 ( .A(n10753), .B(n10752), .ZN(n11509) );
  INV_X1 U12726 ( .A(n16382), .ZN(n16553) );
  OAI211_X1 U12727 ( .C1(n11345), .C2(n10754), .A(n10778), .B(n14430), .ZN(
        n11507) );
  OAI21_X1 U12728 ( .B1(n10754), .B2(n16553), .A(n11507), .ZN(n10755) );
  AOI21_X1 U12729 ( .B1(n11509), .B2(n14717), .A(n10755), .ZN(n10756) );
  NAND2_X1 U12730 ( .A1(n11511), .A2(n10756), .ZN(n10906) );
  NAND2_X1 U12731 ( .A1(n10906), .A2(n11936), .ZN(n10757) );
  OAI21_X1 U12732 ( .B1(n11936), .B2(n10758), .A(n10757), .ZN(P2_U3439) );
  INV_X1 U12733 ( .A(n10759), .ZN(n10772) );
  AOI21_X1 U12734 ( .B1(n10761), .B2(n10760), .A(n15925), .ZN(n10763) );
  NAND2_X1 U12735 ( .A1(n10763), .A2(n10762), .ZN(n10771) );
  NAND2_X1 U12736 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n12052)
         );
  AOI21_X1 U12737 ( .B1(n10765), .B2(n10764), .A(n16285), .ZN(n10767) );
  NAND2_X1 U12738 ( .A1(n10767), .A2(n10766), .ZN(n10768) );
  NAND2_X1 U12739 ( .A1(n12052), .A2(n10768), .ZN(n10769) );
  AOI21_X1 U12740 ( .B1(n15892), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10769), 
        .ZN(n10770) );
  OAI211_X1 U12741 ( .C1(n15928), .C2(n10772), .A(n10771), .B(n10770), .ZN(
        P1_U3253) );
  INV_X1 U12742 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10781) );
  XNOR2_X1 U12743 ( .A(n10773), .B(n14290), .ZN(n11363) );
  OAI21_X1 U12744 ( .B1(n10775), .B2(n14290), .A(n10774), .ZN(n10776) );
  OAI22_X1 U12745 ( .A1(n10889), .A2(n13967), .B1(n14043), .B2(n13968), .ZN(
        n10887) );
  AOI21_X1 U12746 ( .B1(n10776), .B2(n14606), .A(n10887), .ZN(n11359) );
  AOI211_X1 U12747 ( .C1(n14034), .C2(n10778), .A(n7437), .B(n10777), .ZN(
        n11358) );
  AOI21_X1 U12748 ( .B1(n16382), .B2(n14034), .A(n11358), .ZN(n10779) );
  OAI211_X1 U12749 ( .C1(n16386), .C2(n11363), .A(n11359), .B(n10779), .ZN(
        n10902) );
  NAND2_X1 U12750 ( .A1(n10902), .A2(n11936), .ZN(n10780) );
  OAI21_X1 U12751 ( .B1(n11936), .B2(n10781), .A(n10780), .ZN(P2_U3442) );
  INV_X1 U12752 ( .A(n10782), .ZN(n10828) );
  AOI22_X1 U12753 ( .A1(n10930), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n15763), .ZN(n10783) );
  OAI21_X1 U12754 ( .B1(n10828), .B2(n15780), .A(n10783), .ZN(P1_U3342) );
  INV_X1 U12755 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n10785) );
  NAND2_X1 U12756 ( .A1(n12944), .A2(P3_U3897), .ZN(n10784) );
  OAI21_X1 U12757 ( .B1(P3_U3897), .B2(n10785), .A(n10784), .ZN(P3_U3513) );
  NAND2_X1 U12758 ( .A1(n13990), .A2(n7437), .ZN(n13976) );
  OAI22_X1 U12759 ( .A1(n10786), .A2(n13976), .B1(n13963), .B2(n14001), .ZN(
        n10788) );
  NAND2_X1 U12760 ( .A1(n10788), .A2(n10787), .ZN(n10790) );
  AND2_X1 U12761 ( .A1(n14366), .A2(n14589), .ZN(n10820) );
  AOI22_X1 U12762 ( .A1(n13972), .A2(n10820), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n10846), .ZN(n10789) );
  OAI211_X1 U12763 ( .C1(n13975), .C2(n14001), .A(n10790), .B(n10789), .ZN(
        P2_U3204) );
  AND2_X1 U12764 ( .A1(n10792), .A2(n10791), .ZN(n10794) );
  OR2_X1 U12765 ( .A1(n10797), .A2(n10805), .ZN(n10793) );
  OAI211_X1 U12766 ( .C1(n10795), .C2(n10803), .A(n10794), .B(n10793), .ZN(
        n10796) );
  NAND2_X1 U12767 ( .A1(n10796), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10802) );
  INV_X1 U12768 ( .A(n10797), .ZN(n10800) );
  NOR2_X1 U12769 ( .A1(n10989), .A2(n10879), .ZN(n12771) );
  INV_X1 U12770 ( .A(n10987), .ZN(n10798) );
  NAND2_X1 U12771 ( .A1(n10798), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12775) );
  INV_X1 U12772 ( .A(n12775), .ZN(n10799) );
  AOI21_X1 U12773 ( .B1(n10800), .B2(n12771), .A(n10799), .ZN(n10801) );
  NOR2_X1 U12774 ( .A1(n12978), .A2(P3_U3151), .ZN(n10986) );
  INV_X1 U12775 ( .A(n10278), .ZN(n12999) );
  NAND2_X1 U12776 ( .A1(n12999), .A2(n11626), .ZN(n12595) );
  NAND2_X1 U12777 ( .A1(n16308), .A2(n12595), .ZN(n12743) );
  NOR2_X1 U12778 ( .A1(n10803), .A2(n16544), .ZN(n10804) );
  NAND2_X1 U12779 ( .A1(n10808), .A2(n10804), .ZN(n10807) );
  OR2_X1 U12780 ( .A1(n10814), .A2(n10805), .ZN(n10806) );
  NAND2_X1 U12781 ( .A1(n10808), .A2(n16544), .ZN(n10812) );
  INV_X1 U12782 ( .A(n10809), .ZN(n10810) );
  AOI22_X1 U12783 ( .A1(n12743), .A2(n7876), .B1(n10813), .B2(n12966), .ZN(
        n10817) );
  OR2_X1 U12784 ( .A1(n10814), .A2(n12732), .ZN(n12976) );
  INV_X1 U12785 ( .A(n12976), .ZN(n12870) );
  NAND2_X1 U12786 ( .A1(n12870), .A2(n13251), .ZN(n12954) );
  INV_X1 U12787 ( .A(n12954), .ZN(n10815) );
  NAND2_X1 U12788 ( .A1(n10815), .A2(n12997), .ZN(n10816) );
  OAI211_X1 U12789 ( .C1(n10986), .C2(n10818), .A(n10817), .B(n10816), .ZN(
        P3_U3172) );
  INV_X1 U12790 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10827) );
  NAND2_X1 U12791 ( .A1(n10819), .A2(n14000), .ZN(n14284) );
  INV_X1 U12792 ( .A(n14284), .ZN(n10944) );
  NAND2_X1 U12793 ( .A1(n11636), .A2(n9148), .ZN(n10821) );
  AOI21_X1 U12794 ( .B1(n14284), .B2(n10821), .A(n10820), .ZN(n10936) );
  INV_X1 U12795 ( .A(n10822), .ZN(n10823) );
  NOR2_X1 U12796 ( .A1(n14001), .A2(n10823), .ZN(n10942) );
  INV_X1 U12797 ( .A(n10942), .ZN(n10824) );
  OAI211_X1 U12798 ( .C1(n10944), .C2(n10825), .A(n10936), .B(n10824), .ZN(
        n10900) );
  NAND2_X1 U12799 ( .A1(n11936), .A2(n10900), .ZN(n10826) );
  OAI21_X1 U12800 ( .B1(n11936), .B2(n10827), .A(n10826), .ZN(P2_U3430) );
  INV_X1 U12801 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10829) );
  INV_X1 U12802 ( .A(n11554), .ZN(n11559) );
  OAI222_X1 U12803 ( .A1(n14787), .A2(n10829), .B1(n14783), .B2(n10828), .C1(
        n11559), .C2(P2_U3088), .ZN(P2_U3314) );
  OAI21_X1 U12804 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n10837), .A(n10830), 
        .ZN(n10831) );
  NAND2_X1 U12805 ( .A1(n10831), .A2(n10833), .ZN(n11064) );
  OAI21_X1 U12806 ( .B1(n10831), .B2(n10833), .A(n11064), .ZN(n10832) );
  NOR2_X1 U12807 ( .A1(n10832), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n11066) );
  AOI21_X1 U12808 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n10832), .A(n11066), 
        .ZN(n10845) );
  AND2_X1 U12809 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n10835) );
  NOR2_X1 U12810 ( .A1(n15842), .A2(n10833), .ZN(n10834) );
  AOI211_X1 U12811 ( .C1(n15875), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n10835), 
        .B(n10834), .ZN(n10844) );
  XNOR2_X1 U12812 ( .A(n11072), .B(n10836), .ZN(n10838) );
  NAND2_X1 U12813 ( .A1(n10837), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10839) );
  NAND3_X1 U12814 ( .A1(n10840), .A2(n10838), .A3(n10839), .ZN(n11071) );
  INV_X1 U12815 ( .A(n11071), .ZN(n10842) );
  AOI21_X1 U12816 ( .B1(n10840), .B2(n10839), .A(n10838), .ZN(n10841) );
  OAI21_X1 U12817 ( .B1(n10842), .B2(n10841), .A(n15873), .ZN(n10843) );
  OAI211_X1 U12818 ( .C1(n10845), .C2(n15848), .A(n10844), .B(n10843), .ZN(
        P2_U3226) );
  NOR2_X1 U12819 ( .A1(n13988), .A2(n13968), .ZN(n13904) );
  INV_X1 U12820 ( .A(n10846), .ZN(n10847) );
  OAI22_X1 U12821 ( .A1(n13975), .A2(n11348), .B1(n10847), .B2(n11347), .ZN(
        n10849) );
  NAND2_X1 U12822 ( .A1(n13972), .A2(n14588), .ZN(n13902) );
  NOR2_X1 U12823 ( .A1(n13902), .A2(n7657), .ZN(n10848) );
  AOI211_X1 U12824 ( .C1(n13904), .C2(n14364), .A(n10849), .B(n10848), .ZN(
        n10856) );
  OAI22_X1 U12825 ( .A1(n7657), .A2(n13976), .B1(n13963), .B2(n10850), .ZN(
        n10854) );
  INV_X1 U12826 ( .A(n10851), .ZN(n10853) );
  NAND3_X1 U12827 ( .A1(n10854), .A2(n10853), .A3(n10852), .ZN(n10855) );
  OAI211_X1 U12828 ( .C1(n10857), .C2(n13963), .A(n10856), .B(n10855), .ZN(
        P2_U3209) );
  NAND2_X1 U12829 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n11469) );
  NAND2_X1 U12830 ( .A1(n10859), .A2(n10858), .ZN(n10860) );
  NAND3_X1 U12831 ( .A1(n15415), .A2(n15382), .A3(n10860), .ZN(n10861) );
  NAND2_X1 U12832 ( .A1(n11469), .A2(n10861), .ZN(n10866) );
  INV_X1 U12833 ( .A(n15388), .ZN(n10862) );
  AOI211_X1 U12834 ( .C1(n10864), .C2(n10863), .A(n10862), .B(n15925), .ZN(
        n10865) );
  AOI211_X1 U12835 ( .C1(n15892), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n10866), .B(
        n10865), .ZN(n10867) );
  OAI21_X1 U12836 ( .B1(n10868), .B2(n15928), .A(n10867), .ZN(P1_U3249) );
  INV_X1 U12837 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10874) );
  AOI21_X1 U12838 ( .B1(n16382), .B2(n14041), .A(n10869), .ZN(n10870) );
  OAI211_X1 U12839 ( .C1(n16386), .C2(n10872), .A(n10871), .B(n10870), .ZN(
        n10904) );
  NAND2_X1 U12840 ( .A1(n10904), .A2(n11936), .ZN(n10873) );
  OAI21_X1 U12841 ( .B1(n11936), .B2(n10874), .A(n10873), .ZN(P2_U3445) );
  INV_X1 U12842 ( .A(n10875), .ZN(n10876) );
  OAI222_X1 U12843 ( .A1(P3_U3151), .A2(n10878), .B1(n13850), .B2(n10877), 
        .C1(n13853), .C2(n10876), .ZN(P3_U3276) );
  NAND3_X1 U12844 ( .A1(n12743), .A2(n16593), .A3(n10879), .ZN(n10880) );
  OAI21_X1 U12845 ( .B1(n9780), .B2(n16352), .A(n10880), .ZN(n11628) );
  INV_X1 U12846 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10881) );
  OAI22_X1 U12847 ( .A1(n11626), .A2(n13837), .B1(n16602), .B2(n10881), .ZN(
        n10882) );
  AOI21_X1 U12848 ( .B1(n16602), .B2(n11628), .A(n10882), .ZN(n10883) );
  INV_X1 U12849 ( .A(n10883), .ZN(P3_U3390) );
  NAND2_X1 U12850 ( .A1(n14363), .A2(n7437), .ZN(n10958) );
  INV_X1 U12851 ( .A(n13985), .ZN(n13970) );
  NAND2_X1 U12852 ( .A1(n13972), .A2(n10887), .ZN(n10888) );
  NAND2_X1 U12853 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n14409) );
  OAI211_X1 U12854 ( .C1(n13970), .C2(n11356), .A(n10888), .B(n14409), .ZN(
        n10896) );
  NOR2_X1 U12855 ( .A1(n13976), .A2(n10889), .ZN(n10892) );
  AOI22_X1 U12856 ( .A1(n10892), .A2(n10891), .B1(n13990), .B2(n10890), .ZN(
        n10894) );
  NOR2_X1 U12857 ( .A1(n10894), .A2(n10893), .ZN(n10895) );
  AOI211_X1 U12858 ( .C1(n14034), .C2(n13983), .A(n10896), .B(n10895), .ZN(
        n10897) );
  OAI21_X1 U12859 ( .B1(n13963), .B2(n10967), .A(n10897), .ZN(P2_U3202) );
  NAND2_X1 U12860 ( .A1(n16560), .A2(n10898), .ZN(n10899) );
  OAI21_X1 U12861 ( .B1(n16560), .B2(n8564), .A(n10899), .ZN(P2_U3500) );
  NAND2_X1 U12862 ( .A1(n16560), .A2(n10900), .ZN(n10901) );
  OAI21_X1 U12863 ( .B1(n16560), .B2(n10534), .A(n10901), .ZN(P2_U3499) );
  NAND2_X1 U12864 ( .A1(n10902), .A2(n16560), .ZN(n10903) );
  OAI21_X1 U12865 ( .B1(n16560), .B2(n10501), .A(n10903), .ZN(P2_U3503) );
  NAND2_X1 U12866 ( .A1(n10904), .A2(n16560), .ZN(n10905) );
  OAI21_X1 U12867 ( .B1(n16560), .B2(n8636), .A(n10905), .ZN(P2_U3504) );
  NAND2_X1 U12868 ( .A1(n10906), .A2(n16560), .ZN(n10907) );
  OAI21_X1 U12869 ( .B1(n16560), .B2(n10500), .A(n10907), .ZN(P2_U3502) );
  OAI21_X1 U12870 ( .B1(n10914), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10908), 
        .ZN(n10925) );
  INV_X1 U12871 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10909) );
  MUX2_X1 U12872 ( .A(n10909), .B(P1_REG2_REG_13__SCAN_IN), .S(n10930), .Z(
        n10924) );
  MUX2_X1 U12873 ( .A(n11489), .B(P1_REG2_REG_14__SCAN_IN), .S(n11487), .Z(
        n10911) );
  NAND2_X1 U12874 ( .A1(n10930), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10912) );
  NAND2_X1 U12875 ( .A1(n10911), .A2(n10912), .ZN(n10910) );
  OAI21_X1 U12876 ( .B1(n10923), .B2(n10910), .A(n15415), .ZN(n10922) );
  INV_X1 U12877 ( .A(n10923), .ZN(n10913) );
  AOI22_X1 U12878 ( .A1(n16287), .A2(n11487), .B1(n15892), .B2(
        P1_ADDR_REG_14__SCAN_IN), .ZN(n10921) );
  NAND2_X1 U12879 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n16616)
         );
  OR2_X1 U12880 ( .A1(n10914), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10915) );
  NAND2_X1 U12881 ( .A1(n10916), .A2(n10915), .ZN(n10929) );
  MUX2_X1 U12882 ( .A(n9431), .B(P1_REG1_REG_13__SCAN_IN), .S(n10930), .Z(
        n10928) );
  NAND2_X1 U12883 ( .A1(n10930), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10917) );
  NAND2_X1 U12884 ( .A1(n10926), .A2(n10917), .ZN(n11491) );
  XNOR2_X1 U12885 ( .A(n11491), .B(n11487), .ZN(n11495) );
  XNOR2_X1 U12886 ( .A(n11495), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n10918) );
  NAND2_X1 U12887 ( .A1(n10918), .A2(n16294), .ZN(n10919) );
  AND2_X1 U12888 ( .A1(n16616), .A2(n10919), .ZN(n10920) );
  OAI211_X1 U12889 ( .C1(n10922), .C2(n11488), .A(n10921), .B(n10920), .ZN(
        P1_U3257) );
  AOI211_X1 U12890 ( .C1(n10925), .C2(n10924), .A(n16285), .B(n10923), .ZN(
        n10934) );
  INV_X1 U12891 ( .A(n10926), .ZN(n10927) );
  AOI211_X1 U12892 ( .C1(n10929), .C2(n10928), .A(n15925), .B(n10927), .ZN(
        n10933) );
  INV_X1 U12893 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n16051) );
  NAND2_X1 U12894 ( .A1(n16287), .A2(n10930), .ZN(n10931) );
  NAND2_X1 U12895 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n12481)
         );
  OAI211_X1 U12896 ( .C1(n16051), .C2(n16301), .A(n10931), .B(n12481), .ZN(
        n10932) );
  OR3_X1 U12897 ( .A1(n10934), .A2(n10933), .A3(n10932), .ZN(P1_U3256) );
  NAND2_X1 U12898 ( .A1(n10942), .A2(n14323), .ZN(n10935) );
  OAI211_X1 U12899 ( .C1(n14624), .C2(n10937), .A(n10936), .B(n10935), .ZN(
        n10938) );
  NAND2_X1 U12900 ( .A1(n11368), .A2(n10938), .ZN(n10939) );
  OAI21_X1 U12901 ( .B1(n11368), .B2(n10940), .A(n10939), .ZN(n10941) );
  AOI21_X1 U12902 ( .B1(n14632), .B2(n10942), .A(n10941), .ZN(n10943) );
  OAI21_X1 U12903 ( .B1(n10944), .B2(n14602), .A(n10943), .ZN(P2_U3265) );
  INV_X1 U12904 ( .A(n10945), .ZN(n10946) );
  NAND2_X1 U12905 ( .A1(n11377), .A2(n13086), .ZN(n10947) );
  NAND2_X1 U12906 ( .A1(n10947), .A2(n11216), .ZN(n10948) );
  XNOR2_X1 U12907 ( .A(n16316), .B(n11080), .ZN(n10950) );
  NAND2_X1 U12908 ( .A1(n10952), .A2(n10953), .ZN(n10979) );
  OAI21_X1 U12909 ( .B1(n10953), .B2(n10952), .A(n10979), .ZN(n10954) );
  NAND2_X1 U12910 ( .A1(n10954), .A2(n7876), .ZN(n10957) );
  NOR2_X1 U12911 ( .A1(n12976), .A2(n16350), .ZN(n12959) );
  OAI22_X1 U12912 ( .A1(n12981), .A2(n8116), .B1(n12954), .B2(n16314), .ZN(
        n10955) );
  AOI21_X1 U12913 ( .B1(n12959), .B2(n12999), .A(n10955), .ZN(n10956) );
  OAI211_X1 U12914 ( .C1(n10986), .C2(n16321), .A(n10957), .B(n10956), .ZN(
        P3_U3162) );
  INV_X1 U12915 ( .A(n10966), .ZN(n10959) );
  NAND2_X1 U12916 ( .A1(n10959), .A2(n10958), .ZN(n10960) );
  NAND2_X1 U12917 ( .A1(n10967), .A2(n10960), .ZN(n10961) );
  XNOR2_X1 U12918 ( .A(n14041), .B(n10884), .ZN(n11132) );
  NAND2_X1 U12919 ( .A1(n14362), .A2(n7437), .ZN(n11133) );
  XNOR2_X1 U12920 ( .A(n11132), .B(n11133), .ZN(n10968) );
  NAND2_X1 U12921 ( .A1(n10961), .A2(n10968), .ZN(n11136) );
  NAND2_X1 U12922 ( .A1(n13972), .A2(n10962), .ZN(n10964) );
  OAI211_X1 U12923 ( .C1(n13970), .C2(n10965), .A(n10964), .B(n10963), .ZN(
        n10972) );
  INV_X1 U12924 ( .A(n13976), .ZN(n13894) );
  AOI22_X1 U12925 ( .A1(n13894), .A2(n14363), .B1(n13990), .B2(n10966), .ZN(
        n10970) );
  INV_X1 U12926 ( .A(n10967), .ZN(n10969) );
  NOR3_X1 U12927 ( .A1(n10970), .A2(n10969), .A3(n10968), .ZN(n10971) );
  AOI211_X1 U12928 ( .C1(n14041), .C2(n13983), .A(n10972), .B(n10971), .ZN(
        n10973) );
  OAI21_X1 U12929 ( .B1(n13963), .B2(n11136), .A(n10973), .ZN(P2_U3199) );
  INV_X1 U12930 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n10975) );
  NAND2_X1 U12931 ( .A1(n12832), .A2(P3_U3897), .ZN(n10974) );
  OAI21_X1 U12932 ( .B1(P3_U3897), .B2(n10975), .A(n10974), .ZN(P3_U3515) );
  XNOR2_X1 U12933 ( .A(n10976), .B(n12821), .ZN(n11082) );
  XNOR2_X1 U12934 ( .A(n11082), .B(n9794), .ZN(n10981) );
  INV_X1 U12935 ( .A(n10977), .ZN(n10978) );
  NAND2_X1 U12936 ( .A1(n10979), .A2(n10978), .ZN(n10980) );
  NAND2_X1 U12937 ( .A1(n10980), .A2(n10981), .ZN(n11084) );
  OAI21_X1 U12938 ( .B1(n10981), .B2(n10980), .A(n11084), .ZN(n10982) );
  NAND2_X1 U12939 ( .A1(n10982), .A2(n7876), .ZN(n10985) );
  OAI22_X1 U12940 ( .A1(n12981), .A2(n16363), .B1(n12954), .B2(n16351), .ZN(
        n10983) );
  AOI21_X1 U12941 ( .B1(n12959), .B2(n12997), .A(n10983), .ZN(n10984) );
  OAI211_X1 U12942 ( .C1(n10986), .C2(n16361), .A(n10985), .B(n10984), .ZN(
        P3_U3177) );
  NAND2_X1 U12943 ( .A1(n12728), .A2(n10987), .ZN(n10988) );
  AND2_X1 U12944 ( .A1(n10988), .A2(n9860), .ZN(n11033) );
  NAND2_X1 U12945 ( .A1(n10989), .A2(n12775), .ZN(n11034) );
  AND2_X1 U12946 ( .A1(n11033), .A2(n11034), .ZN(n11032) );
  MUX2_X1 U12947 ( .A(n11032), .B(P3_U3897), .S(n12770), .Z(n16269) );
  MUX2_X1 U12948 ( .A(n10992), .B(n10991), .S(n13036), .Z(n10993) );
  NAND2_X1 U12949 ( .A1(n10993), .A2(n13855), .ZN(n10997) );
  INV_X1 U12950 ( .A(n10993), .ZN(n10994) );
  INV_X1 U12951 ( .A(n13855), .ZN(n11131) );
  NAND2_X1 U12952 ( .A1(n10994), .A2(n11131), .ZN(n10995) );
  NAND2_X1 U12953 ( .A1(n10997), .A2(n10995), .ZN(n11126) );
  INV_X1 U12954 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11452) );
  MUX2_X1 U12955 ( .A(n11452), .B(n10996), .S(n13036), .Z(n13002) );
  NAND2_X1 U12956 ( .A1(n13002), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11125) );
  INV_X1 U12957 ( .A(n10997), .ZN(n11057) );
  MUX2_X1 U12958 ( .A(n10999), .B(n10998), .S(n13036), .Z(n11000) );
  NAND2_X1 U12959 ( .A1(n11000), .A2(n7779), .ZN(n16122) );
  INV_X1 U12960 ( .A(n11000), .ZN(n11001) );
  NAND2_X1 U12961 ( .A1(n11001), .A2(n11026), .ZN(n11002) );
  AND2_X1 U12962 ( .A1(n16122), .A2(n11002), .ZN(n11056) );
  MUX2_X1 U12963 ( .A(n16114), .B(n11003), .S(n13036), .Z(n11004) );
  NAND2_X1 U12964 ( .A1(n11004), .A2(n7767), .ZN(n11007) );
  INV_X1 U12965 ( .A(n11004), .ZN(n11005) );
  NAND2_X1 U12966 ( .A1(n11005), .A2(n11028), .ZN(n11006) );
  NAND2_X1 U12967 ( .A1(n11007), .A2(n11006), .ZN(n16121) );
  INV_X1 U12968 ( .A(n11007), .ZN(n11094) );
  MUX2_X1 U12969 ( .A(n11595), .B(n11008), .S(n13036), .Z(n11009) );
  NAND2_X1 U12970 ( .A1(n11009), .A2(n11097), .ZN(n11012) );
  INV_X1 U12971 ( .A(n11009), .ZN(n11010) );
  NAND2_X1 U12972 ( .A1(n11010), .A2(n11113), .ZN(n11011) );
  AND2_X1 U12973 ( .A1(n11012), .A2(n11011), .ZN(n11093) );
  NAND2_X1 U12974 ( .A1(n11092), .A2(n11012), .ZN(n11014) );
  MUX2_X1 U12975 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13036), .Z(n11241) );
  XNOR2_X1 U12976 ( .A(n11241), .B(n11251), .ZN(n11013) );
  NAND2_X1 U12977 ( .A1(n11014), .A2(n11013), .ZN(n11240) );
  OAI21_X1 U12978 ( .B1(n11014), .B2(n11013), .A(n11240), .ZN(n11015) );
  NAND2_X1 U12979 ( .A1(P3_U3897), .A2(n7430), .ZN(n16263) );
  INV_X1 U12980 ( .A(n16263), .ZN(n16195) );
  NAND2_X1 U12981 ( .A1(n11015), .A2(n16195), .ZN(n11041) );
  INV_X1 U12982 ( .A(n11016), .ZN(n11017) );
  INV_X1 U12983 ( .A(n13008), .ZN(n11018) );
  NAND2_X1 U12984 ( .A1(n13855), .A2(n11018), .ZN(n11019) );
  NAND2_X1 U12985 ( .A1(n9789), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n11020) );
  NAND2_X1 U12986 ( .A1(n11019), .A2(n11020), .ZN(n11118) );
  OR2_X1 U12987 ( .A1(n11118), .A2(n10992), .ZN(n11120) );
  OAI21_X1 U12988 ( .B1(n11026), .B2(P3_REG2_REG_2__SCAN_IN), .A(n11043), .ZN(
        n11021) );
  NAND2_X1 U12989 ( .A1(n11026), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n11046) );
  OAI21_X1 U12990 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n11022), .A(n11247), .ZN(
        n11039) );
  NAND2_X1 U12991 ( .A1(n13005), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n11023) );
  NAND2_X1 U12992 ( .A1(n13855), .A2(n11023), .ZN(n11024) );
  NAND2_X1 U12993 ( .A1(n9789), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n11025) );
  NAND2_X1 U12994 ( .A1(n11024), .A2(n11025), .ZN(n11114) );
  NAND2_X1 U12995 ( .A1(n11116), .A2(n11025), .ZN(n11049) );
  NAND2_X1 U12996 ( .A1(n11050), .A2(n11049), .ZN(n11048) );
  NAND2_X1 U12997 ( .A1(n11026), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n11027) );
  NAND2_X1 U12998 ( .A1(n11029), .A2(n11028), .ZN(n11101) );
  MUX2_X1 U12999 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n11008), .S(n11113), .Z(
        n11103) );
  INV_X1 U13000 ( .A(n11103), .ZN(n11030) );
  AOI21_X1 U13001 ( .B1(n9835), .B2(n11031), .A(n11252), .ZN(n11037) );
  NAND2_X1 U13002 ( .A1(n11032), .A2(n13036), .ZN(n16274) );
  INV_X1 U13003 ( .A(n11033), .ZN(n11035) );
  NOR2_X1 U13004 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13679), .ZN(n11518) );
  AOI21_X1 U13005 ( .B1(n16259), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11518), .ZN(
        n11036) );
  OAI21_X1 U13006 ( .B1(n11037), .B2(n16274), .A(n11036), .ZN(n11038) );
  AOI21_X1 U13007 ( .B1(n16194), .B2(n11039), .A(n11038), .ZN(n11040) );
  OAI211_X1 U13008 ( .C1(n16142), .C2(n11246), .A(n11041), .B(n11040), .ZN(
        P3_U3187) );
  INV_X1 U13009 ( .A(n16194), .ZN(n16277) );
  NOR3_X1 U13010 ( .A1(n16277), .A2(n11043), .A3(P3_REG2_REG_2__SCAN_IN), .ZN(
        n11042) );
  OAI21_X1 U13011 ( .B1(n11042), .B2(n16269), .A(n7779), .ZN(n11055) );
  AOI22_X1 U13012 ( .A1(n16259), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n11054) );
  INV_X1 U13013 ( .A(n11043), .ZN(n11047) );
  INV_X1 U13014 ( .A(n11044), .ZN(n11045) );
  OAI211_X1 U13015 ( .C1(n11047), .C2(n11046), .A(n16194), .B(n11045), .ZN(
        n11053) );
  INV_X1 U13016 ( .A(n16274), .ZN(n16181) );
  OAI21_X1 U13017 ( .B1(n11050), .B2(n11049), .A(n11048), .ZN(n11051) );
  NAND2_X1 U13018 ( .A1(n16181), .A2(n11051), .ZN(n11052) );
  AND4_X1 U13019 ( .A1(n11055), .A2(n11054), .A3(n11053), .A4(n11052), .ZN(
        n11061) );
  INV_X1 U13020 ( .A(n16123), .ZN(n11059) );
  NOR3_X1 U13021 ( .A1(n11128), .A2(n11057), .A3(n11056), .ZN(n11058) );
  OAI21_X1 U13022 ( .B1(n11059), .B2(n11058), .A(n16195), .ZN(n11060) );
  NAND2_X1 U13023 ( .A1(n11061), .A2(n11060), .ZN(P3_U3184) );
  INV_X1 U13024 ( .A(n11062), .ZN(n11160) );
  AOI22_X1 U13025 ( .A1(n11487), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n15763), .ZN(n11063) );
  OAI21_X1 U13026 ( .B1(n11160), .B2(n15780), .A(n11063), .ZN(P1_U3341) );
  INV_X1 U13027 ( .A(n11064), .ZN(n11065) );
  NOR2_X1 U13028 ( .A1(n11066), .A2(n11065), .ZN(n11070) );
  NAND2_X1 U13029 ( .A1(n11554), .A2(n12092), .ZN(n11067) );
  OAI21_X1 U13030 ( .B1(n11554), .B2(n12092), .A(n11067), .ZN(n11069) );
  NAND2_X1 U13031 ( .A1(n11559), .A2(n12092), .ZN(n11068) );
  OAI211_X1 U13032 ( .C1(n11559), .C2(n12092), .A(n11070), .B(n11068), .ZN(
        n11558) );
  OAI211_X1 U13033 ( .C1(n11070), .C2(n11069), .A(n11558), .B(n15877), .ZN(
        n11079) );
  NAND2_X1 U13034 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n11720)
         );
  XNOR2_X1 U13035 ( .A(n11554), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n11074) );
  OAI21_X1 U13036 ( .B1(n11072), .B2(P2_REG1_REG_12__SCAN_IN), .A(n11071), 
        .ZN(n11073) );
  NOR2_X1 U13037 ( .A1(n11073), .A2(n11074), .ZN(n11553) );
  AOI211_X1 U13038 ( .C1(n11074), .C2(n11073), .A(n11553), .B(n15830), .ZN(
        n11075) );
  INV_X1 U13039 ( .A(n11075), .ZN(n11076) );
  NAND2_X1 U13040 ( .A1(n11720), .A2(n11076), .ZN(n11077) );
  AOI21_X1 U13041 ( .B1(n15875), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n11077), 
        .ZN(n11078) );
  OAI211_X1 U13042 ( .C1(n15842), .C2(n11559), .A(n11079), .B(n11078), .ZN(
        P2_U3227) );
  XNOR2_X1 U13043 ( .A(n11081), .B(n11080), .ZN(n11293) );
  XNOR2_X1 U13044 ( .A(n11293), .B(n16351), .ZN(n11085) );
  NAND2_X1 U13045 ( .A1(n11082), .A2(n16314), .ZN(n11086) );
  NAND2_X1 U13046 ( .A1(n11084), .A2(n11083), .ZN(n11295) );
  NAND2_X1 U13047 ( .A1(n11295), .A2(n7876), .ZN(n11091) );
  AOI21_X1 U13048 ( .B1(n11084), .B2(n11086), .A(n11085), .ZN(n11090) );
  MUX2_X1 U13049 ( .A(n12978), .B(P3_U3151), .S(P3_REG3_REG_3__SCAN_IN), .Z(
        n11088) );
  OAI22_X1 U13050 ( .A1(n12981), .A2(n16390), .B1(n12954), .B2(n11738), .ZN(
        n11087) );
  AOI211_X1 U13051 ( .C1(n12959), .C2(n9794), .A(n11088), .B(n11087), .ZN(
        n11089) );
  OAI21_X1 U13052 ( .B1(n11091), .B2(n11090), .A(n11089), .ZN(P3_U3158) );
  INV_X1 U13053 ( .A(n11092), .ZN(n11096) );
  NOR3_X1 U13054 ( .A1(n16120), .A2(n11094), .A3(n11093), .ZN(n11095) );
  OAI21_X1 U13055 ( .B1(n11096), .B2(n11095), .A(n16195), .ZN(n11112) );
  MUX2_X1 U13056 ( .A(n11595), .B(P3_REG2_REG_4__SCAN_IN), .S(n11097), .Z(
        n11099) );
  NAND2_X1 U13057 ( .A1(n11100), .A2(n11099), .ZN(n11098) );
  OAI21_X1 U13058 ( .B1(n11100), .B2(n11099), .A(n11098), .ZN(n11110) );
  INV_X1 U13059 ( .A(n16259), .ZN(n16151) );
  INV_X1 U13060 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15960) );
  INV_X1 U13061 ( .A(n11101), .ZN(n11102) );
  NOR3_X1 U13062 ( .A1(n16116), .A2(n11103), .A3(n11102), .ZN(n11104) );
  OAI21_X1 U13063 ( .B1(n11105), .B2(n11104), .A(n16181), .ZN(n11108) );
  NOR2_X1 U13064 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11106), .ZN(n11300) );
  INV_X1 U13065 ( .A(n11300), .ZN(n11107) );
  OAI211_X1 U13066 ( .C1(n16151), .C2(n15960), .A(n11108), .B(n11107), .ZN(
        n11109) );
  AOI21_X1 U13067 ( .B1(n16194), .B2(n11110), .A(n11109), .ZN(n11111) );
  OAI211_X1 U13068 ( .C1(n16142), .C2(n11113), .A(n11112), .B(n11111), .ZN(
        P3_U3186) );
  AOI22_X1 U13069 ( .A1(n16259), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n11124) );
  NAND2_X1 U13070 ( .A1(n11114), .A2(n10991), .ZN(n11115) );
  NAND2_X1 U13071 ( .A1(n11116), .A2(n11115), .ZN(n11117) );
  NAND2_X1 U13072 ( .A1(n16181), .A2(n11117), .ZN(n11123) );
  NAND2_X1 U13073 ( .A1(n11118), .A2(n10992), .ZN(n11119) );
  NAND2_X1 U13074 ( .A1(n11120), .A2(n11119), .ZN(n11121) );
  NAND2_X1 U13075 ( .A1(n16194), .A2(n11121), .ZN(n11122) );
  AND3_X1 U13076 ( .A1(n11124), .A2(n11123), .A3(n11122), .ZN(n11130) );
  AND2_X1 U13077 ( .A1(n11126), .A2(n11125), .ZN(n11127) );
  OAI21_X1 U13078 ( .B1(n11128), .B2(n11127), .A(n16195), .ZN(n11129) );
  OAI211_X1 U13079 ( .C1(n16142), .C2(n11131), .A(n11130), .B(n11129), .ZN(
        P3_U3183) );
  INV_X1 U13080 ( .A(n11132), .ZN(n11134) );
  NAND2_X1 U13081 ( .A1(n11134), .A2(n11133), .ZN(n11135) );
  XNOR2_X1 U13082 ( .A(n14047), .B(n10884), .ZN(n11137) );
  AND2_X1 U13083 ( .A1(n14361), .A2(n7437), .ZN(n11138) );
  NAND2_X1 U13084 ( .A1(n11137), .A2(n11138), .ZN(n11142) );
  INV_X1 U13085 ( .A(n11137), .ZN(n11310) );
  INV_X1 U13086 ( .A(n11138), .ZN(n11139) );
  NAND2_X1 U13087 ( .A1(n11310), .A2(n11139), .ZN(n11140) );
  NAND2_X1 U13088 ( .A1(n11142), .A2(n11140), .ZN(n11220) );
  XNOR2_X1 U13089 ( .A(n14055), .B(n10884), .ZN(n11155) );
  NAND2_X1 U13090 ( .A1(n14360), .A2(n7437), .ZN(n11143) );
  XNOR2_X1 U13091 ( .A(n11155), .B(n11143), .ZN(n11314) );
  INV_X1 U13092 ( .A(n11155), .ZN(n11144) );
  NAND2_X1 U13093 ( .A1(n11144), .A2(n11143), .ZN(n11145) );
  XNOR2_X1 U13094 ( .A(n14061), .B(n10884), .ZN(n11225) );
  NAND2_X1 U13095 ( .A1(n14359), .A2(n7437), .ZN(n11226) );
  XNOR2_X1 U13096 ( .A(n11225), .B(n11226), .ZN(n11154) );
  NAND2_X1 U13097 ( .A1(n14360), .A2(n14588), .ZN(n11147) );
  NAND2_X1 U13098 ( .A1(n14358), .A2(n14589), .ZN(n11146) );
  NAND2_X1 U13099 ( .A1(n11147), .A2(n11146), .ZN(n11383) );
  INV_X1 U13100 ( .A(n11383), .ZN(n11152) );
  NAND2_X1 U13101 ( .A1(n13983), .A2(n14061), .ZN(n11151) );
  INV_X1 U13102 ( .A(n11385), .ZN(n11149) );
  AOI21_X1 U13103 ( .B1(n13985), .B2(n11149), .A(n11148), .ZN(n11150) );
  OAI211_X1 U13104 ( .C1(n11152), .C2(n13988), .A(n11151), .B(n11150), .ZN(
        n11153) );
  INV_X1 U13105 ( .A(n11153), .ZN(n11159) );
  NAND2_X1 U13106 ( .A1(n13990), .A2(n11155), .ZN(n11156) );
  OAI21_X1 U13107 ( .B1(n13976), .B2(n14057), .A(n11156), .ZN(n11157) );
  NAND3_X1 U13108 ( .A1(n11319), .A2(n7668), .A3(n11157), .ZN(n11158) );
  OAI211_X1 U13109 ( .C1(n11237), .C2(n13963), .A(n11159), .B(n11158), .ZN(
        P2_U3193) );
  INV_X1 U13110 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11161) );
  INV_X1 U13111 ( .A(n11555), .ZN(n11806) );
  OAI222_X1 U13112 ( .A1(n14787), .A2(n11161), .B1(n14783), .B2(n11160), .C1(
        P2_U3088), .C2(n11806), .ZN(P2_U3313) );
  INV_X1 U13113 ( .A(n11162), .ZN(n11163) );
  AOI21_X1 U13114 ( .B1(n8194), .B2(n11164), .A(n11163), .ZN(n11343) );
  INV_X1 U13115 ( .A(n11165), .ZN(n11167) );
  OAI21_X1 U13116 ( .B1(n11167), .B2(n8194), .A(n11166), .ZN(n11168) );
  OAI22_X1 U13117 ( .A1(n14043), .A2(n13967), .B1(n14057), .B2(n13968), .ZN(
        n11217) );
  AOI21_X1 U13118 ( .B1(n11168), .B2(n14606), .A(n11217), .ZN(n11336) );
  AOI21_X1 U13119 ( .B1(n14047), .B2(n11169), .A(n7437), .ZN(n11170) );
  NAND2_X1 U13120 ( .A1(n11413), .A2(n11170), .ZN(n11337) );
  OAI211_X1 U13121 ( .C1(n11343), .C2(n16386), .A(n11336), .B(n11337), .ZN(
        n11380) );
  OAI22_X1 U13122 ( .A1(n14768), .A2(n11378), .B1(n11936), .B2(n8651), .ZN(
        n11171) );
  AOI21_X1 U13123 ( .B1(n11380), .B2(n11936), .A(n11171), .ZN(n11172) );
  INV_X1 U13124 ( .A(n11172), .ZN(P2_U3448) );
  NAND2_X1 U13125 ( .A1(n11568), .A2(n11567), .ZN(n11186) );
  NAND2_X1 U13126 ( .A1(n11186), .A2(n11570), .ZN(n11282) );
  AND2_X1 U13127 ( .A1(n11282), .A2(n11572), .ZN(n16398) );
  INV_X1 U13128 ( .A(n16610), .ZN(n15003) );
  OR2_X1 U13129 ( .A1(n11186), .A2(n15294), .ZN(n15009) );
  INV_X2 U13130 ( .A(n15009), .ZN(n16614) );
  INV_X1 U13131 ( .A(n15327), .ZN(n11179) );
  OAI22_X1 U13132 ( .A1(n11179), .A2(n15293), .B1(n11210), .B2(n15016), .ZN(
        n16334) );
  NAND2_X1 U13133 ( .A1(n11282), .A2(n11175), .ZN(n11200) );
  AOI22_X1 U13134 ( .A1(n16614), .A2(n16334), .B1(n11200), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n11193) );
  XNOR2_X1 U13135 ( .A(n11176), .B(n14827), .ZN(n11205) );
  OR2_X4 U13136 ( .A1(n11208), .A2(n16473), .ZN(n14830) );
  OAI22_X1 U13137 ( .A1(n14830), .A2(n9269), .B1(n16339), .B2(n14863), .ZN(
        n11203) );
  XNOR2_X1 U13138 ( .A(n11205), .B(n11203), .ZN(n11201) );
  INV_X1 U13139 ( .A(n11177), .ZN(n11180) );
  AOI22_X1 U13140 ( .A1(n11755), .A2(n11574), .B1(n11180), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n11178) );
  OAI21_X1 U13141 ( .B1(n14830), .B2(n11179), .A(n11178), .ZN(n11195) );
  NAND2_X1 U13142 ( .A1(n11180), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n11181) );
  NAND2_X1 U13143 ( .A1(n11195), .A2(n11194), .ZN(n11197) );
  OR2_X1 U13144 ( .A1(n11194), .A2(n14919), .ZN(n11185) );
  AND2_X1 U13145 ( .A1(n11197), .A2(n11185), .ZN(n11202) );
  XNOR2_X1 U13146 ( .A(n11201), .B(n11202), .ZN(n11191) );
  INV_X1 U13147 ( .A(n11186), .ZN(n11190) );
  INV_X1 U13148 ( .A(n11572), .ZN(n11188) );
  NAND2_X1 U13149 ( .A1(n16476), .A2(n15033), .ZN(n11187) );
  NOR2_X1 U13150 ( .A1(n11188), .A2(n11187), .ZN(n11189) );
  NAND2_X1 U13151 ( .A1(n11191), .A2(n16612), .ZN(n11192) );
  OAI211_X1 U13152 ( .C1(n15003), .C2(n16339), .A(n11193), .B(n11192), .ZN(
        P1_U3222) );
  OR2_X1 U13153 ( .A1(n11195), .A2(n11194), .ZN(n11196) );
  AND2_X1 U13154 ( .A1(n11197), .A2(n11196), .ZN(n15344) );
  AND2_X1 U13155 ( .A1(n15008), .A2(n9636), .ZN(n11577) );
  AOI22_X1 U13156 ( .A1(n16612), .A2(n15344), .B1(n16614), .B2(n11577), .ZN(
        n11199) );
  NAND2_X1 U13157 ( .A1(n11200), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n11198) );
  OAI211_X1 U13158 ( .C1(n15003), .C2(n16327), .A(n11199), .B(n11198), .ZN(
        P1_U3232) );
  AOI22_X1 U13159 ( .A1(n16614), .A2(n11989), .B1(n11200), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n11213) );
  NAND2_X1 U13160 ( .A1(n11202), .A2(n11201), .ZN(n11207) );
  INV_X1 U13161 ( .A(n11203), .ZN(n11204) );
  NAND2_X1 U13162 ( .A1(n11205), .A2(n11204), .ZN(n11206) );
  NAND2_X1 U13163 ( .A1(n11207), .A2(n11206), .ZN(n11269) );
  OAI22_X1 U13164 ( .A1(n16374), .A2(n11208), .B1(n14863), .B2(n11210), .ZN(
        n11209) );
  XNOR2_X1 U13165 ( .A(n11209), .B(n14827), .ZN(n11272) );
  OAI22_X1 U13166 ( .A1(n14830), .A2(n11210), .B1(n16374), .B2(n14863), .ZN(
        n11270) );
  XNOR2_X1 U13167 ( .A(n11272), .B(n11270), .ZN(n11268) );
  XNOR2_X1 U13168 ( .A(n11269), .B(n11268), .ZN(n11211) );
  NAND2_X1 U13169 ( .A1(n11211), .A2(n16612), .ZN(n11212) );
  OAI211_X1 U13170 ( .C1(n15003), .C2(n16374), .A(n11213), .B(n11212), .ZN(
        P1_U3237) );
  INV_X1 U13171 ( .A(n11214), .ZN(n11215) );
  OAI222_X1 U13172 ( .A1(P3_U3151), .A2(n11216), .B1(n13850), .B2(n7989), .C1(
        n13853), .C2(n11215), .ZN(P3_U3275) );
  NAND2_X1 U13173 ( .A1(n13972), .A2(n11217), .ZN(n11218) );
  NAND2_X1 U13174 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n15840) );
  OAI211_X1 U13175 ( .C1(n13970), .C2(n11338), .A(n11218), .B(n15840), .ZN(
        n11223) );
  INV_X1 U13176 ( .A(n11219), .ZN(n11313) );
  AOI211_X1 U13177 ( .C1(n11221), .C2(n11220), .A(n13963), .B(n11313), .ZN(
        n11222) );
  AOI211_X1 U13178 ( .C1(n14047), .C2(n13983), .A(n11223), .B(n11222), .ZN(
        n11224) );
  INV_X1 U13179 ( .A(n11224), .ZN(P2_U3211) );
  INV_X1 U13180 ( .A(n11225), .ZN(n11235) );
  NAND2_X1 U13181 ( .A1(n11235), .A2(n11226), .ZN(n11227) );
  XNOR2_X1 U13182 ( .A(n14629), .B(n10884), .ZN(n11392) );
  NAND2_X1 U13183 ( .A1(n14358), .A2(n7437), .ZN(n11393) );
  XNOR2_X1 U13184 ( .A(n11392), .B(n11393), .ZN(n11233) );
  OAI21_X1 U13185 ( .B1(n13970), .B2(n14625), .A(n11228), .ZN(n11232) );
  NAND2_X1 U13186 ( .A1(n14359), .A2(n14588), .ZN(n11230) );
  NAND2_X1 U13187 ( .A1(n14357), .A2(n14589), .ZN(n11229) );
  AND2_X1 U13188 ( .A1(n11230), .A2(n11229), .ZN(n11609) );
  NOR2_X1 U13189 ( .A1(n13988), .A2(n11609), .ZN(n11231) );
  AOI211_X1 U13190 ( .C1(n14629), .C2(n13983), .A(n11232), .B(n11231), .ZN(
        n11239) );
  OAI22_X1 U13191 ( .A1(n11235), .A2(n13963), .B1(n13976), .B2(n11234), .ZN(
        n11236) );
  NAND3_X1 U13192 ( .A1(n11237), .A2(n7974), .A3(n11236), .ZN(n11238) );
  OAI211_X1 U13193 ( .C1(n11403), .C2(n13963), .A(n11239), .B(n11238), .ZN(
        P2_U3203) );
  MUX2_X1 U13194 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n13036), .Z(n11523) );
  XNOR2_X1 U13195 ( .A(n11523), .B(n11526), .ZN(n11244) );
  OAI21_X1 U13196 ( .B1(n11241), .B2(n11246), .A(n11240), .ZN(n16141) );
  MUX2_X1 U13197 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n13036), .Z(n11242) );
  NAND2_X1 U13198 ( .A1(n11242), .A2(n16143), .ZN(n16139) );
  AOI21_X1 U13199 ( .B1(n11244), .B2(n11243), .A(n7615), .ZN(n11262) );
  NAND2_X1 U13200 ( .A1(n11246), .A2(n11245), .ZN(n11248) );
  NAND2_X1 U13201 ( .A1(P3_REG2_REG_7__SCAN_IN), .A2(n11249), .ZN(n11527) );
  OAI21_X1 U13202 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n11249), .A(n11527), .ZN(
        n11260) );
  INV_X1 U13203 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11253) );
  MUX2_X1 U13204 ( .A(n11253), .B(P3_REG1_REG_6__SCAN_IN), .S(n16143), .Z(
        n16135) );
  NAND2_X1 U13205 ( .A1(n16143), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n11254) );
  AOI21_X1 U13206 ( .B1(n11255), .B2(n9877), .A(n11535), .ZN(n11258) );
  INV_X1 U13207 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15988) );
  NAND2_X1 U13208 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11690) );
  OAI21_X1 U13209 ( .B1(n16151), .B2(n15988), .A(n11690), .ZN(n11256) );
  AOI21_X1 U13210 ( .B1(n11534), .B2(n16269), .A(n11256), .ZN(n11257) );
  OAI21_X1 U13211 ( .B1(n11258), .B2(n16274), .A(n11257), .ZN(n11259) );
  AOI21_X1 U13212 ( .B1(n16194), .B2(n11260), .A(n11259), .ZN(n11261) );
  OAI21_X1 U13213 ( .B1(n11262), .B2(n16263), .A(n11261), .ZN(P3_U3189) );
  INV_X1 U13214 ( .A(n11263), .ZN(n11266) );
  INV_X1 U13215 ( .A(n15404), .ZN(n11499) );
  OAI222_X1 U13216 ( .A1(n15777), .A2(n11264), .B1(n15780), .B2(n11266), .C1(
        n11499), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U13217 ( .A(n12349), .ZN(n11815) );
  INV_X1 U13218 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11265) );
  OAI222_X1 U13219 ( .A1(P2_U3088), .A2(n11815), .B1(n14783), .B2(n11266), 
        .C1(n11265), .C2(n14787), .ZN(P2_U3312) );
  OAI22_X1 U13220 ( .A1(n15056), .A2(n14863), .B1(n11208), .B2(n15055), .ZN(
        n11267) );
  XNOR2_X1 U13221 ( .A(n11267), .B(n14919), .ZN(n11320) );
  INV_X1 U13222 ( .A(n11270), .ZN(n11271) );
  NAND2_X1 U13223 ( .A1(n11272), .A2(n11271), .ZN(n11273) );
  XNOR2_X1 U13224 ( .A(n11274), .B(n14919), .ZN(n11276) );
  XNOR2_X1 U13225 ( .A(n11276), .B(n11275), .ZN(n16399) );
  NAND2_X1 U13226 ( .A1(n11276), .A2(n11275), .ZN(n11277) );
  OAI22_X1 U13227 ( .A1(n14830), .A2(n15056), .B1(n15055), .B2(n14863), .ZN(
        n11278) );
  NAND2_X1 U13228 ( .A1(n11321), .A2(n11322), .ZN(n11279) );
  XOR2_X1 U13229 ( .A(n11320), .B(n11279), .Z(n11289) );
  INV_X1 U13230 ( .A(n11280), .ZN(n11281) );
  NAND2_X1 U13231 ( .A1(n11282), .A2(n11281), .ZN(n11283) );
  NAND2_X1 U13232 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n16298) );
  NAND2_X1 U13233 ( .A1(n15008), .A2(n15324), .ZN(n11285) );
  NAND2_X1 U13234 ( .A1(n15006), .A2(n15326), .ZN(n11284) );
  NAND2_X1 U13235 ( .A1(n11285), .A2(n11284), .ZN(n16424) );
  NAND2_X1 U13236 ( .A1(n16614), .A2(n16424), .ZN(n11286) );
  OAI211_X1 U13237 ( .C1(n16619), .C2(n12058), .A(n16298), .B(n11286), .ZN(
        n11287) );
  AOI21_X1 U13238 ( .B1(n16610), .B2(n16425), .A(n11287), .ZN(n11288) );
  OAI21_X1 U13239 ( .B1(n11289), .B2(n15029), .A(n11288), .ZN(P1_U3230) );
  INV_X1 U13240 ( .A(n11290), .ZN(n11292) );
  OAI22_X1 U13241 ( .A1(n12773), .A2(P3_U3151), .B1(SI_22_), .B2(n13850), .ZN(
        n11291) );
  AOI21_X1 U13242 ( .B1(n11292), .B2(n11550), .A(n11291), .ZN(P3_U3273) );
  NAND2_X1 U13243 ( .A1(n11295), .A2(n11294), .ZN(n11298) );
  XNOR2_X1 U13244 ( .A(n11597), .B(n12821), .ZN(n11296) );
  NAND2_X1 U13245 ( .A1(n11296), .A2(n11738), .ZN(n11512) );
  OAI21_X1 U13246 ( .B1(n11296), .B2(n11738), .A(n11512), .ZN(n11297) );
  AOI21_X1 U13247 ( .B1(n11298), .B2(n11297), .A(n11514), .ZN(n11304) );
  INV_X1 U13248 ( .A(n12959), .ZN(n12141) );
  OAI22_X1 U13249 ( .A1(n12141), .A2(n16351), .B1(n11926), .B2(n12954), .ZN(
        n11299) );
  AOI211_X1 U13250 ( .C1(n11597), .C2(n12966), .A(n11300), .B(n11299), .ZN(
        n11303) );
  INV_X1 U13251 ( .A(n11301), .ZN(n11596) );
  NAND2_X1 U13252 ( .A1(n12978), .A2(n11596), .ZN(n11302) );
  OAI211_X1 U13253 ( .C1(n11304), .C2(n12969), .A(n11303), .B(n11302), .ZN(
        P3_U3170) );
  NAND2_X1 U13254 ( .A1(n13904), .A2(n14359), .ZN(n11309) );
  INV_X1 U13255 ( .A(n11416), .ZN(n11307) );
  INV_X1 U13256 ( .A(n11305), .ZN(n11306) );
  AOI21_X1 U13257 ( .B1(n13985), .B2(n11307), .A(n11306), .ZN(n11308) );
  OAI211_X1 U13258 ( .C1(n13902), .C2(n11311), .A(n11309), .B(n11308), .ZN(
        n11317) );
  NOR3_X1 U13259 ( .A1(n13976), .A2(n11311), .A3(n11310), .ZN(n11312) );
  AOI21_X1 U13260 ( .B1(n11313), .B2(n13990), .A(n11312), .ZN(n11315) );
  NOR2_X1 U13261 ( .A1(n11315), .A2(n11314), .ZN(n11316) );
  AOI211_X1 U13262 ( .C1(n14055), .C2(n13983), .A(n11317), .B(n11316), .ZN(
        n11318) );
  OAI21_X1 U13263 ( .B1(n13963), .B2(n11319), .A(n11318), .ZN(P2_U3185) );
  NAND2_X1 U13264 ( .A1(n11321), .A2(n11320), .ZN(n11323) );
  NAND2_X1 U13265 ( .A1(n11323), .A2(n11322), .ZN(n11456) );
  NAND2_X1 U13266 ( .A1(n14918), .A2(n15324), .ZN(n11325) );
  NAND2_X1 U13267 ( .A1(n14916), .A2(n16448), .ZN(n11324) );
  AND2_X1 U13268 ( .A1(n11325), .A2(n11324), .ZN(n11454) );
  INV_X1 U13269 ( .A(n11454), .ZN(n11458) );
  NAND2_X1 U13270 ( .A1(n14917), .A2(n16448), .ZN(n11327) );
  NAND2_X1 U13271 ( .A1(n14916), .A2(n15324), .ZN(n11326) );
  NAND2_X1 U13272 ( .A1(n11327), .A2(n11326), .ZN(n11328) );
  XNOR2_X1 U13273 ( .A(n11328), .B(n14827), .ZN(n11457) );
  XNOR2_X1 U13274 ( .A(n11458), .B(n11457), .ZN(n11329) );
  XNOR2_X1 U13275 ( .A(n11456), .B(n11329), .ZN(n11335) );
  AND2_X1 U13276 ( .A1(n16448), .A2(n16573), .ZN(n16441) );
  OR2_X1 U13277 ( .A1(n15056), .A2(n15293), .ZN(n11331) );
  NAND2_X1 U13278 ( .A1(n15008), .A2(n15323), .ZN(n11330) );
  NAND2_X1 U13279 ( .A1(n11331), .A2(n11330), .ZN(n16447) );
  AOI22_X1 U13280 ( .A1(n16614), .A2(n16447), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11332) );
  OAI21_X1 U13281 ( .B1(n16449), .B2(n16619), .A(n11332), .ZN(n11333) );
  AOI21_X1 U13282 ( .B1(n16398), .B2(n16441), .A(n11333), .ZN(n11334) );
  OAI21_X1 U13283 ( .B1(n11335), .B2(n15029), .A(n11334), .ZN(P1_U3227) );
  MUX2_X1 U13284 ( .A(n10482), .B(n11336), .S(n11368), .Z(n11342) );
  INV_X1 U13285 ( .A(n11337), .ZN(n11340) );
  OAI22_X1 U13286 ( .A1(n14619), .A2(n11378), .B1(n14624), .B2(n11338), .ZN(
        n11339) );
  AOI21_X1 U13287 ( .B1(n14632), .B2(n11340), .A(n11339), .ZN(n11341) );
  OAI211_X1 U13288 ( .C1(n14580), .C2(n11343), .A(n11342), .B(n11341), .ZN(
        P2_U3259) );
  AOI211_X1 U13289 ( .C1(n16381), .C2(n11346), .A(n7437), .B(n11345), .ZN(
        n16380) );
  OAI22_X1 U13290 ( .A1(n14619), .A2(n11348), .B1(n14624), .B2(n11347), .ZN(
        n11349) );
  AOI21_X1 U13291 ( .B1(n14632), .B2(n16380), .A(n11349), .ZN(n11355) );
  AOI222_X1 U13292 ( .A1(n14606), .A2(n11352), .B1(n14364), .B2(n14589), .C1(
        n14366), .C2(n14588), .ZN(n16384) );
  MUX2_X1 U13293 ( .A(n11353), .B(n16384), .S(n11368), .Z(n11354) );
  OAI211_X1 U13294 ( .C1(n14580), .C2(n16385), .A(n11355), .B(n11354), .ZN(
        P2_U3263) );
  OAI22_X1 U13295 ( .A1(n14619), .A2(n7981), .B1(n14624), .B2(n11356), .ZN(
        n11357) );
  AOI21_X1 U13296 ( .B1(n14632), .B2(n11358), .A(n11357), .ZN(n11362) );
  MUX2_X1 U13297 ( .A(n11360), .B(n11359), .S(n11368), .Z(n11361) );
  OAI211_X1 U13298 ( .C1(n14580), .C2(n11363), .A(n11362), .B(n11361), .ZN(
        P2_U3261) );
  OAI22_X1 U13299 ( .A1(n14619), .A2(n11365), .B1(n11364), .B2(n14624), .ZN(
        n11366) );
  AOI21_X1 U13300 ( .B1(n14632), .B2(n11367), .A(n11366), .ZN(n11372) );
  MUX2_X1 U13301 ( .A(n11370), .B(n11369), .S(n11368), .Z(n11371) );
  OAI211_X1 U13302 ( .C1(n14580), .C2(n11373), .A(n11372), .B(n11371), .ZN(
        P2_U3264) );
  INV_X1 U13303 ( .A(n11374), .ZN(n11375) );
  OAI222_X1 U13304 ( .A1(P3_U3151), .A2(n11377), .B1(n13850), .B2(n11376), 
        .C1(n13853), .C2(n11375), .ZN(P3_U3274) );
  OAI22_X1 U13305 ( .A1(n14715), .A2(n11378), .B1(n16560), .B2(n10505), .ZN(
        n11379) );
  AOI21_X1 U13306 ( .B1(n11380), .B2(n16560), .A(n11379), .ZN(n11381) );
  INV_X1 U13307 ( .A(n11381), .ZN(P2_U3505) );
  XOR2_X1 U13308 ( .A(n11382), .B(n14294), .Z(n11384) );
  AOI21_X1 U13309 ( .B1(n11384), .B2(n14606), .A(n11383), .ZN(n11478) );
  OAI22_X1 U13310 ( .A1(n11368), .A2(n11386), .B1(n11385), .B2(n14624), .ZN(
        n11388) );
  OAI211_X1 U13311 ( .C1(n11483), .C2(n7610), .A(n14430), .B(n11605), .ZN(
        n11477) );
  INV_X1 U13312 ( .A(n14632), .ZN(n14556) );
  NOR2_X1 U13313 ( .A1(n11477), .A2(n14556), .ZN(n11387) );
  AOI211_X1 U13314 ( .C1(n14628), .C2(n14061), .A(n11388), .B(n11387), .ZN(
        n11391) );
  XNOR2_X1 U13315 ( .A(n11389), .B(n14294), .ZN(n11479) );
  OR2_X1 U13316 ( .A1(n11479), .A2(n14580), .ZN(n11390) );
  OAI211_X1 U13317 ( .C1(n11478), .C2(n14622), .A(n11391), .B(n11390), .ZN(
        P2_U3257) );
  INV_X1 U13318 ( .A(n11392), .ZN(n11400) );
  NAND2_X1 U13319 ( .A1(n11400), .A2(n11393), .ZN(n11394) );
  XNOR2_X1 U13320 ( .A(n14073), .B(n10884), .ZN(n11708) );
  NAND2_X1 U13321 ( .A1(n14357), .A2(n7437), .ZN(n11709) );
  XNOR2_X1 U13322 ( .A(n11708), .B(n11709), .ZN(n11399) );
  NOR2_X1 U13323 ( .A1(n13902), .A2(n11632), .ZN(n11398) );
  NAND2_X1 U13324 ( .A1(n13904), .A2(n14356), .ZN(n11396) );
  OAI211_X1 U13325 ( .C1(n13970), .C2(n11637), .A(n11396), .B(n11395), .ZN(
        n11397) );
  AOI211_X1 U13326 ( .C1(n14073), .C2(n13983), .A(n11398), .B(n11397), .ZN(
        n11405) );
  OAI22_X1 U13327 ( .A1(n11400), .A2(n13963), .B1(n11632), .B2(n13976), .ZN(
        n11401) );
  NAND3_X1 U13328 ( .A1(n11403), .A2(n11402), .A3(n11401), .ZN(n11404) );
  OAI211_X1 U13329 ( .C1(n11711), .C2(n13963), .A(n11405), .B(n11404), .ZN(
        P2_U3189) );
  OAI21_X1 U13330 ( .B1(n7620), .B2(n14295), .A(n11406), .ZN(n11420) );
  AOI22_X1 U13331 ( .A1(n14588), .A2(n14361), .B1(n14359), .B2(n14589), .ZN(
        n11411) );
  XNOR2_X1 U13332 ( .A(n11408), .B(n11407), .ZN(n11409) );
  NAND2_X1 U13333 ( .A1(n11409), .A2(n14606), .ZN(n11410) );
  OAI211_X1 U13334 ( .C1(n11420), .C2(n11636), .A(n11411), .B(n11410), .ZN(
        n11421) );
  MUX2_X1 U13335 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11421), .S(n11368), .Z(
        n11412) );
  INV_X1 U13336 ( .A(n11412), .ZN(n11419) );
  NAND2_X1 U13337 ( .A1(n11413), .A2(n14055), .ZN(n11414) );
  NAND2_X1 U13338 ( .A1(n11414), .A2(n14430), .ZN(n11415) );
  NOR2_X1 U13339 ( .A1(n7610), .A2(n11415), .ZN(n11422) );
  INV_X1 U13340 ( .A(n14055), .ZN(n11427) );
  OAI22_X1 U13341 ( .A1(n14619), .A2(n11427), .B1(n11416), .B2(n14624), .ZN(
        n11417) );
  AOI21_X1 U13342 ( .B1(n14632), .B2(n11422), .A(n11417), .ZN(n11418) );
  OAI211_X1 U13343 ( .C1(n11420), .C2(n14602), .A(n11419), .B(n11418), .ZN(
        P2_U3258) );
  INV_X1 U13344 ( .A(n11420), .ZN(n11423) );
  AOI211_X1 U13345 ( .C1(n11423), .C2(n16558), .A(n11422), .B(n11421), .ZN(
        n11430) );
  INV_X1 U13346 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n11424) );
  OAI22_X1 U13347 ( .A1(n14768), .A2(n11427), .B1(n11936), .B2(n11424), .ZN(
        n11425) );
  INV_X1 U13348 ( .A(n11425), .ZN(n11426) );
  OAI21_X1 U13349 ( .B1(n11430), .B2(n16561), .A(n11426), .ZN(P2_U3451) );
  OAI22_X1 U13350 ( .A1(n14715), .A2(n11427), .B1(n16560), .B2(n10506), .ZN(
        n11428) );
  INV_X1 U13351 ( .A(n11428), .ZN(n11429) );
  OAI21_X1 U13352 ( .B1(n11430), .B2(n16559), .A(n11429), .ZN(P2_U3506) );
  NAND2_X1 U13353 ( .A1(n12998), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n11431) );
  OAI21_X1 U13354 ( .B1(n12574), .B2(n12998), .A(n11431), .ZN(P3_U3521) );
  NAND2_X1 U13355 ( .A1(n12998), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11432) );
  OAI21_X1 U13356 ( .B1(n13109), .B2(n12998), .A(n11432), .ZN(P3_U3520) );
  INV_X1 U13357 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n13383) );
  NAND2_X1 U13358 ( .A1(n9770), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n11435) );
  NAND2_X1 U13359 ( .A1(n11433), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n11434) );
  OAI211_X1 U13360 ( .C1(n11436), .C2(n13383), .A(n11435), .B(n11434), .ZN(
        n11437) );
  INV_X1 U13361 ( .A(n11437), .ZN(n11438) );
  NAND2_X1 U13362 ( .A1(n12998), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(n11440) );
  OAI21_X1 U13363 ( .B1(n13091), .B2(n12998), .A(n11440), .ZN(P3_U3522) );
  INV_X1 U13364 ( .A(n11441), .ZN(n11448) );
  NAND2_X1 U13365 ( .A1(n11442), .A2(n11443), .ZN(n11446) );
  OR2_X1 U13366 ( .A1(n11444), .A2(n11443), .ZN(n11445) );
  AND2_X1 U13367 ( .A1(n11446), .A2(n11445), .ZN(n11447) );
  NAND2_X1 U13368 ( .A1(n11448), .A2(n11447), .ZN(n11450) );
  INV_X1 U13369 ( .A(n11450), .ZN(n11449) );
  INV_X1 U13370 ( .A(n12733), .ZN(n11591) );
  NOR2_X1 U13371 ( .A1(n16593), .A2(n11591), .ZN(n16320) );
  NAND2_X2 U13372 ( .A1(n11449), .A2(n16320), .ZN(n13304) );
  INV_X1 U13373 ( .A(n16360), .ZN(n13291) );
  AOI21_X1 U13374 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n13291), .A(n11628), .ZN(
        n11451) );
  MUX2_X1 U13375 ( .A(n11452), .B(n11451), .S(n13310), .Z(n11453) );
  OAI21_X1 U13376 ( .B1(n11626), .B2(n13304), .A(n11453), .ZN(P3_U3233) );
  NAND2_X1 U13377 ( .A1(n11457), .A2(n11454), .ZN(n11455) );
  NAND2_X1 U13378 ( .A1(n11456), .A2(n11455), .ZN(n11461) );
  INV_X1 U13379 ( .A(n11457), .ZN(n11459) );
  NAND2_X1 U13380 ( .A1(n11459), .A2(n11458), .ZN(n11460) );
  NAND2_X1 U13381 ( .A1(n11461), .A2(n11460), .ZN(n11749) );
  NAND2_X1 U13382 ( .A1(n16465), .A2(n14917), .ZN(n11463) );
  NAND2_X1 U13383 ( .A1(n14916), .A2(n15323), .ZN(n11462) );
  NAND2_X1 U13384 ( .A1(n11463), .A2(n11462), .ZN(n11464) );
  XNOR2_X1 U13385 ( .A(n11464), .B(n14827), .ZN(n11750) );
  NAND2_X1 U13386 ( .A1(n16465), .A2(n14916), .ZN(n11465) );
  OAI21_X1 U13387 ( .B1(n11466), .B2(n14830), .A(n11465), .ZN(n11751) );
  XNOR2_X1 U13388 ( .A(n11750), .B(n11751), .ZN(n11748) );
  XNOR2_X1 U13389 ( .A(n11749), .B(n11748), .ZN(n11472) );
  OAI22_X1 U13390 ( .A1(n11467), .A2(n15293), .B1(n11768), .B2(n15016), .ZN(
        n11975) );
  NAND2_X1 U13391 ( .A1(n16614), .A2(n11975), .ZN(n11468) );
  OAI211_X1 U13392 ( .C1(n16619), .C2(n11979), .A(n11469), .B(n11468), .ZN(
        n11470) );
  AOI21_X1 U13393 ( .B1(n16610), .B2(n16465), .A(n11470), .ZN(n11471) );
  OAI21_X1 U13394 ( .B1(n11472), .B2(n15029), .A(n11471), .ZN(P1_U3239) );
  INV_X1 U13395 ( .A(n11473), .ZN(n11475) );
  INV_X1 U13396 ( .A(n15407), .ZN(n15927) );
  OAI222_X1 U13397 ( .A1(n15777), .A2(n11474), .B1(n15780), .B2(n11475), .C1(
        n15927), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U13398 ( .A(n15859), .ZN(n12340) );
  OAI222_X1 U13399 ( .A1(n14787), .A2(n11476), .B1(n14783), .B2(n11475), .C1(
        n12340), .C2(P2_U3088), .ZN(P2_U3311) );
  OAI211_X1 U13400 ( .C1(n16386), .C2(n11479), .A(n11478), .B(n11477), .ZN(
        n11485) );
  INV_X1 U13401 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n11480) );
  OAI22_X1 U13402 ( .A1(n14768), .A2(n11483), .B1(n11936), .B2(n11480), .ZN(
        n11481) );
  AOI21_X1 U13403 ( .B1(n11485), .B2(n11936), .A(n11481), .ZN(n11482) );
  INV_X1 U13404 ( .A(n11482), .ZN(P2_U3454) );
  OAI22_X1 U13405 ( .A1(n14715), .A2(n11483), .B1(n16560), .B2(n8694), .ZN(
        n11484) );
  AOI21_X1 U13406 ( .B1(n11485), .B2(n16560), .A(n11484), .ZN(n11486) );
  INV_X1 U13407 ( .A(n11486), .ZN(P2_U3507) );
  INV_X1 U13408 ( .A(n11487), .ZN(n11492) );
  XNOR2_X1 U13409 ( .A(n7502), .B(n15404), .ZN(n11490) );
  NOR2_X1 U13410 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n11490), .ZN(n15405) );
  AOI21_X1 U13411 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n11490), .A(n15405), 
        .ZN(n11504) );
  INV_X1 U13412 ( .A(n11491), .ZN(n11493) );
  OAI22_X1 U13413 ( .A1(n11495), .A2(n11494), .B1(n11493), .B2(n11492), .ZN(
        n15394) );
  XOR2_X1 U13414 ( .A(n11499), .B(n15394), .Z(n11496) );
  NOR2_X1 U13415 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n11496), .ZN(n15395) );
  AOI21_X1 U13416 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n11496), .A(n15395), 
        .ZN(n11497) );
  OR2_X1 U13417 ( .A1(n11497), .A2(n15925), .ZN(n11503) );
  NOR2_X1 U13418 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11498), .ZN(n11501) );
  NOR2_X1 U13419 ( .A1(n15928), .A2(n11499), .ZN(n11500) );
  AOI211_X1 U13420 ( .C1(n15892), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n11501), 
        .B(n11500), .ZN(n11502) );
  OAI211_X1 U13421 ( .C1(n11504), .C2(n16285), .A(n11503), .B(n11502), .ZN(
        P1_U3258) );
  OAI22_X1 U13422 ( .A1(n11368), .A2(n10481), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14624), .ZN(n11505) );
  AOI21_X1 U13423 ( .B1(n14628), .B2(n14027), .A(n11505), .ZN(n11506) );
  OAI21_X1 U13424 ( .B1(n14556), .B2(n11507), .A(n11506), .ZN(n11508) );
  AOI21_X1 U13425 ( .B1(n11509), .B2(n14630), .A(n11508), .ZN(n11510) );
  OAI21_X1 U13426 ( .B1(n14622), .B2(n11511), .A(n11510), .ZN(P2_U3262) );
  INV_X1 U13427 ( .A(n11512), .ZN(n11513) );
  XNOR2_X1 U13428 ( .A(n11703), .B(n12821), .ZN(n11618) );
  XNOR2_X1 U13429 ( .A(n11618), .B(n11926), .ZN(n11515) );
  AOI21_X1 U13430 ( .B1(n11516), .B2(n11515), .A(n11619), .ZN(n11522) );
  OAI22_X1 U13431 ( .A1(n12141), .A2(n11738), .B1(n12622), .B2(n12954), .ZN(
        n11517) );
  AOI211_X1 U13432 ( .C1(n11703), .C2(n12966), .A(n11518), .B(n11517), .ZN(
        n11521) );
  INV_X1 U13433 ( .A(n11965), .ZN(n11519) );
  NAND2_X1 U13434 ( .A1(n12978), .A2(n11519), .ZN(n11520) );
  OAI211_X1 U13435 ( .C1(n11522), .C2(n12969), .A(n11521), .B(n11520), .ZN(
        P3_U3167) );
  MUX2_X1 U13436 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13036), .Z(n11668) );
  XNOR2_X1 U13437 ( .A(n11668), .B(n11667), .ZN(n11669) );
  INV_X1 U13438 ( .A(n11523), .ZN(n11524) );
  XOR2_X1 U13439 ( .A(n11669), .B(n11670), .Z(n11545) );
  NAND2_X1 U13440 ( .A1(n11526), .A2(n11525), .ZN(n11528) );
  MUX2_X1 U13441 ( .A(P3_REG2_REG_8__SCAN_IN), .B(n11529), .S(n11667), .Z(
        n11530) );
  OAI21_X1 U13442 ( .B1(n11531), .B2(n11530), .A(n11659), .ZN(n11543) );
  INV_X1 U13443 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n13470) );
  NOR2_X1 U13444 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13470), .ZN(n12024) );
  AOI21_X1 U13445 ( .B1(n16259), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n12024), .ZN(
        n11532) );
  OAI21_X1 U13446 ( .B1(n16142), .B2(n11667), .A(n11532), .ZN(n11542) );
  NOR2_X1 U13447 ( .A1(n11534), .A2(n11533), .ZN(n11536) );
  MUX2_X1 U13448 ( .A(n11537), .B(P3_REG1_REG_8__SCAN_IN), .S(n11667), .Z(
        n11538) );
  NAND2_X1 U13449 ( .A1(n11539), .A2(n11538), .ZN(n11540) );
  AOI21_X1 U13450 ( .B1(n11663), .B2(n11540), .A(n16274), .ZN(n11541) );
  AOI211_X1 U13451 ( .C1(n16194), .C2(n11543), .A(n11542), .B(n11541), .ZN(
        n11544) );
  OAI21_X1 U13452 ( .B1(n11545), .B2(n16263), .A(n11544), .ZN(P3_U3190) );
  INV_X1 U13453 ( .A(n11546), .ZN(n11548) );
  INV_X1 U13454 ( .A(n15403), .ZN(n15904) );
  OAI222_X1 U13455 ( .A1(n15777), .A2(n11547), .B1(n15780), .B2(n11548), .C1(
        P1_U3086), .C2(n15904), .ZN(P1_U3338) );
  INV_X1 U13456 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11549) );
  INV_X1 U13457 ( .A(n12354), .ZN(n15868) );
  OAI222_X1 U13458 ( .A1(n14787), .A2(n11549), .B1(n14783), .B2(n11548), .C1(
        P2_U3088), .C2(n15868), .ZN(P2_U3310) );
  NAND2_X1 U13459 ( .A1(n11551), .A2(n11550), .ZN(n11552) );
  OAI211_X1 U13460 ( .C1(n13614), .C2(n13850), .A(n11552), .B(n12775), .ZN(
        P3_U3272) );
  AOI21_X1 U13461 ( .B1(n11554), .B2(P2_REG1_REG_13__SCAN_IN), .A(n11553), 
        .ZN(n11808) );
  XNOR2_X1 U13462 ( .A(n11555), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n11807) );
  XNOR2_X1 U13463 ( .A(n11808), .B(n11807), .ZN(n11566) );
  NAND2_X1 U13464 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n11892)
         );
  INV_X1 U13465 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11557) );
  NAND2_X1 U13466 ( .A1(n11555), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11803) );
  INV_X1 U13467 ( .A(n11803), .ZN(n11556) );
  AOI21_X1 U13468 ( .B1(n11557), .B2(n11806), .A(n11556), .ZN(n11561) );
  OAI21_X1 U13469 ( .B1(n11559), .B2(n12092), .A(n11558), .ZN(n11560) );
  NAND2_X1 U13470 ( .A1(n11561), .A2(n11560), .ZN(n11802) );
  OAI211_X1 U13471 ( .C1(n11561), .C2(n11560), .A(n15877), .B(n11802), .ZN(
        n11562) );
  NAND2_X1 U13472 ( .A1(n11892), .A2(n11562), .ZN(n11564) );
  NOR2_X1 U13473 ( .A1(n15842), .A2(n11806), .ZN(n11563) );
  AOI211_X1 U13474 ( .C1(n15875), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n11564), 
        .B(n11563), .ZN(n11565) );
  OAI21_X1 U13475 ( .B1(n11566), .B2(n15830), .A(n11565), .ZN(P2_U3228) );
  NOR2_X1 U13476 ( .A1(n11567), .A2(n15294), .ZN(n11569) );
  NAND2_X1 U13477 ( .A1(n11569), .A2(n11568), .ZN(n12781) );
  INV_X1 U13478 ( .A(n11570), .ZN(n11571) );
  NAND2_X2 U13479 ( .A1(n11572), .A2(n11571), .ZN(n16490) );
  AND2_X4 U13480 ( .A1(n12781), .A2(n16490), .ZN(n16522) );
  INV_X1 U13481 ( .A(n16522), .ZN(n15515) );
  AOI21_X1 U13482 ( .B1(n15217), .B2(n15515), .A(n16518), .ZN(n11584) );
  NAND2_X1 U13483 ( .A1(n11977), .A2(n11574), .ZN(n16302) );
  OR2_X1 U13484 ( .A1(n11575), .A2(n15417), .ZN(n15215) );
  NOR2_X1 U13485 ( .A1(n16522), .A2(n15215), .ZN(n16513) );
  NAND2_X1 U13486 ( .A1(n15327), .A2(n16327), .ZN(n15039) );
  NAND2_X1 U13487 ( .A1(n16331), .A2(n15039), .ZN(n16306) );
  NAND2_X1 U13488 ( .A1(n16370), .A2(n16479), .ZN(n11578) );
  AOI21_X1 U13489 ( .B1(n11578), .B2(n16306), .A(n11577), .ZN(n16303) );
  OAI22_X1 U13490 ( .A1(n16522), .A2(n16303), .B1(n11579), .B2(n16490), .ZN(
        n11582) );
  INV_X1 U13491 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n11580) );
  NOR2_X1 U13492 ( .A1(n15515), .A2(n11580), .ZN(n11581) );
  AOI211_X1 U13493 ( .C1(n16513), .C2(n16306), .A(n11582), .B(n11581), .ZN(
        n11583) );
  OAI21_X1 U13494 ( .B1(n11584), .B2(n16302), .A(n11583), .ZN(P1_U3293) );
  INV_X1 U13495 ( .A(n11585), .ZN(n11587) );
  INV_X1 U13496 ( .A(n14413), .ZN(n12345) );
  OAI222_X1 U13497 ( .A1(n14787), .A2(n11586), .B1(n14783), .B2(n11587), .C1(
        n12345), .C2(P2_U3088), .ZN(P2_U3309) );
  INV_X1 U13498 ( .A(n15410), .ZN(n15914) );
  OAI222_X1 U13499 ( .A1(n15777), .A2(n11588), .B1(n15780), .B2(n11587), .C1(
        n15914), .C2(P1_U3086), .ZN(P1_U3337) );
  NAND3_X1 U13500 ( .A1(n11731), .A2(n12608), .A3(n12738), .ZN(n11589) );
  AND2_X1 U13501 ( .A1(n11590), .A2(n11589), .ZN(n16415) );
  NAND2_X1 U13502 ( .A1(n12594), .A2(n11591), .ZN(n12123) );
  NAND2_X1 U13503 ( .A1(n16541), .A2(n12123), .ZN(n16367) );
  XNOR2_X1 U13504 ( .A(n11592), .B(n12610), .ZN(n11594) );
  OAI22_X1 U13505 ( .A1(n16351), .A2(n16350), .B1(n11926), .B2(n16352), .ZN(
        n11593) );
  AOI21_X1 U13506 ( .B1(n11594), .B2(n13299), .A(n11593), .ZN(n16418) );
  MUX2_X1 U13507 ( .A(n11595), .B(n16418), .S(n13310), .Z(n11599) );
  INV_X1 U13508 ( .A(n13304), .ZN(n13260) );
  AOI22_X1 U13509 ( .A1(n13260), .A2(n11597), .B1(n13291), .B2(n11596), .ZN(
        n11598) );
  OAI211_X1 U13510 ( .C1(n16415), .C2(n13313), .A(n11599), .B(n11598), .ZN(
        P3_U3229) );
  INV_X1 U13511 ( .A(n11600), .ZN(n11602) );
  OAI222_X1 U13512 ( .A1(n15777), .A2(n11601), .B1(n15780), .B2(n11602), .C1(
        P1_U3086), .C2(n15417), .ZN(P1_U3336) );
  INV_X1 U13513 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11603) );
  OAI222_X1 U13514 ( .A1(n14787), .A2(n11603), .B1(n14783), .B2(n11602), .C1(
        n14424), .C2(P2_U3088), .ZN(P2_U3308) );
  XNOR2_X1 U13515 ( .A(n11604), .B(n14297), .ZN(n14631) );
  AOI21_X1 U13516 ( .B1(n14629), .B2(n11605), .A(n7437), .ZN(n11606) );
  AND2_X1 U13517 ( .A1(n11606), .A2(n11639), .ZN(n14633) );
  OAI211_X1 U13518 ( .C1(n11608), .C2(n14297), .A(n11607), .B(n14606), .ZN(
        n11610) );
  NAND2_X1 U13519 ( .A1(n11610), .A2(n11609), .ZN(n14623) );
  AOI211_X1 U13520 ( .C1(n14717), .C2(n14631), .A(n14633), .B(n14623), .ZN(
        n11615) );
  INV_X1 U13521 ( .A(n14715), .ZN(n12239) );
  AOI22_X1 U13522 ( .A1(n14629), .A2(n12239), .B1(n16559), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11611) );
  OAI21_X1 U13523 ( .B1(n11615), .B2(n16559), .A(n11611), .ZN(P2_U3508) );
  INV_X1 U13524 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11612) );
  NOR2_X1 U13525 ( .A1(n11936), .A2(n11612), .ZN(n11613) );
  AOI21_X1 U13526 ( .B1(n14629), .B2(n9744), .A(n11613), .ZN(n11614) );
  OAI21_X1 U13527 ( .B1(n11615), .B2(n16561), .A(n11614), .ZN(P2_U3457) );
  INV_X1 U13528 ( .A(n11616), .ZN(n11706) );
  OAI222_X1 U13529 ( .A1(n15777), .A2(n11617), .B1(n15780), .B2(n11706), .C1(
        n15212), .C2(P1_U3086), .ZN(P1_U3335) );
  XNOR2_X1 U13530 ( .A(n12620), .B(n12821), .ZN(n11686) );
  XNOR2_X1 U13531 ( .A(n11686), .B(n12995), .ZN(n11620) );
  OAI211_X1 U13532 ( .C1(n11621), .C2(n11620), .A(n11688), .B(n7876), .ZN(
        n11625) );
  INV_X1 U13533 ( .A(n12620), .ZN(n16458) );
  NOR2_X1 U13534 ( .A1(n12981), .A2(n16458), .ZN(n11623) );
  OAI22_X1 U13535 ( .A1(n12141), .A2(n11926), .B1(n12022), .B2(n12954), .ZN(
        n11622) );
  AOI211_X1 U13536 ( .C1(P3_REG3_REG_6__SCAN_IN), .C2(P3_U3151), .A(n11623), 
        .B(n11622), .ZN(n11624) );
  OAI211_X1 U13537 ( .C1(n11920), .C2(n12955), .A(n11625), .B(n11624), .ZN(
        P3_U3179) );
  OAI22_X1 U13538 ( .A1(n13379), .A2(n11626), .B1(n16601), .B2(n10996), .ZN(
        n11627) );
  AOI21_X1 U13539 ( .B1(n11628), .B2(n16601), .A(n11627), .ZN(n11629) );
  INV_X1 U13540 ( .A(n11629), .ZN(P3_U3459) );
  XNOR2_X1 U13541 ( .A(n14073), .B(n14357), .ZN(n14296) );
  XOR2_X1 U13542 ( .A(n11630), .B(n14296), .Z(n16551) );
  XOR2_X1 U13543 ( .A(n14296), .B(n11631), .Z(n11634) );
  OAI22_X1 U13544 ( .A1(n11632), .A2(n13967), .B1(n11906), .B2(n13968), .ZN(
        n11633) );
  AOI21_X1 U13545 ( .B1(n11634), .B2(n14606), .A(n11633), .ZN(n11635) );
  OAI21_X1 U13546 ( .B1(n16551), .B2(n11636), .A(n11635), .ZN(n16555) );
  NAND2_X1 U13547 ( .A1(n16555), .A2(n11368), .ZN(n11644) );
  OAI22_X1 U13548 ( .A1(n11368), .A2(n11638), .B1(n11637), .B2(n14624), .ZN(
        n11642) );
  INV_X1 U13549 ( .A(n14073), .ZN(n16554) );
  INV_X1 U13550 ( .A(n11639), .ZN(n11640) );
  OAI211_X1 U13551 ( .C1(n16554), .C2(n11640), .A(n14430), .B(n11652), .ZN(
        n16552) );
  NOR2_X1 U13552 ( .A1(n16552), .A2(n14556), .ZN(n11641) );
  AOI211_X1 U13553 ( .C1(n14628), .C2(n14073), .A(n11642), .B(n11641), .ZN(
        n11643) );
  OAI211_X1 U13554 ( .C1(n16551), .C2(n14602), .A(n11644), .B(n11643), .ZN(
        P2_U3255) );
  XNOR2_X1 U13555 ( .A(n11645), .B(n14299), .ZN(n11935) );
  INV_X1 U13556 ( .A(n11935), .ZN(n11658) );
  XNOR2_X1 U13557 ( .A(n11647), .B(n11646), .ZN(n11650) );
  NAND2_X1 U13558 ( .A1(n14355), .A2(n14589), .ZN(n11649) );
  NAND2_X1 U13559 ( .A1(n14357), .A2(n14588), .ZN(n11648) );
  AND2_X1 U13560 ( .A1(n11649), .A2(n11648), .ZN(n11878) );
  OAI21_X1 U13561 ( .B1(n11650), .B2(n9148), .A(n11878), .ZN(n11933) );
  NAND2_X1 U13562 ( .A1(n11933), .A2(n11368), .ZN(n11657) );
  AOI211_X1 U13563 ( .C1(n14086), .C2(n11652), .A(n7437), .B(n11651), .ZN(
        n11934) );
  INV_X1 U13564 ( .A(n14086), .ZN(n11653) );
  NOR2_X1 U13565 ( .A1(n11653), .A2(n14619), .ZN(n11655) );
  OAI22_X1 U13566 ( .A1(n11368), .A2(n10707), .B1(n11875), .B2(n14624), .ZN(
        n11654) );
  AOI211_X1 U13567 ( .C1(n11934), .C2(n14632), .A(n11655), .B(n11654), .ZN(
        n11656) );
  OAI211_X1 U13568 ( .C1(n14580), .C2(n11658), .A(n11657), .B(n11656), .ZN(
        P2_U3254) );
  INV_X1 U13569 ( .A(n11667), .ZN(n11660) );
  OAI21_X1 U13570 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n11661), .A(n11832), .ZN(
        n11675) );
  INV_X1 U13571 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n16527) );
  NAND2_X1 U13572 ( .A1(n11667), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n11662) );
  XNOR2_X1 U13573 ( .A(n16527), .B(n11818), .ZN(n11664) );
  NAND2_X1 U13574 ( .A1(n11664), .A2(n16181), .ZN(n11666) );
  NOR2_X1 U13575 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13489), .ZN(n12143) );
  AOI21_X1 U13576 ( .B1(n16259), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n12143), .ZN(
        n11665) );
  OAI211_X1 U13577 ( .C1(n16142), .C2(n11831), .A(n11666), .B(n11665), .ZN(
        n11674) );
  MUX2_X1 U13578 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n13036), .Z(n11826) );
  XNOR2_X1 U13579 ( .A(n11826), .B(n11831), .ZN(n11672) );
  NOR2_X1 U13580 ( .A1(n11671), .A2(n11672), .ZN(n11825) );
  AOI211_X1 U13581 ( .C1(n11672), .C2(n11671), .A(n16263), .B(n11825), .ZN(
        n11673) );
  AOI211_X1 U13582 ( .C1(n16194), .C2(n11675), .A(n11674), .B(n11673), .ZN(
        n11676) );
  INV_X1 U13583 ( .A(n11676), .ZN(P3_U3191) );
  INV_X1 U13584 ( .A(n11677), .ZN(n11679) );
  OAI222_X1 U13585 ( .A1(n15777), .A2(n11678), .B1(n15780), .B2(n11679), .C1(
        P1_U3086), .C2(n15218), .ZN(P1_U3334) );
  OAI222_X1 U13586 ( .A1(n14787), .A2(n11680), .B1(n14783), .B2(n11679), .C1(
        n14276), .C2(P2_U3088), .ZN(P2_U3306) );
  INV_X1 U13587 ( .A(n11681), .ZN(n11685) );
  INV_X1 U13588 ( .A(n11682), .ZN(n11684) );
  OAI222_X1 U13589 ( .A1(P3_U3151), .A2(n11685), .B1(n13853), .B2(n11684), 
        .C1(n11683), .C2(n13850), .ZN(P3_U3271) );
  XNOR2_X1 U13590 ( .A(n11859), .B(n11080), .ZN(n12016) );
  XNOR2_X1 U13591 ( .A(n12016), .B(n12022), .ZN(n12017) );
  XNOR2_X1 U13592 ( .A(n12018), .B(n12017), .ZN(n11694) );
  INV_X1 U13593 ( .A(n11689), .ZN(n11852) );
  OAI21_X1 U13594 ( .B1(n12981), .B2(n11862), .A(n11690), .ZN(n11692) );
  OAI22_X1 U13595 ( .A1(n12141), .A2(n12622), .B1(n12140), .B2(n12954), .ZN(
        n11691) );
  AOI211_X1 U13596 ( .C1(n11852), .C2(n12978), .A(n11692), .B(n11691), .ZN(
        n11693) );
  OAI21_X1 U13597 ( .B1(n11694), .B2(n12969), .A(n11693), .ZN(P3_U3153) );
  OAI21_X1 U13598 ( .B1(n11695), .B2(n12746), .A(n11917), .ZN(n11970) );
  INV_X1 U13599 ( .A(n11696), .ZN(n11697) );
  AOI21_X1 U13600 ( .B1(n12746), .B2(n11698), .A(n11697), .ZN(n11699) );
  OAI222_X1 U13601 ( .A1(n16352), .A2(n12622), .B1(n16350), .B2(n11738), .C1(
        n16349), .C2(n11699), .ZN(n11967) );
  AOI21_X1 U13602 ( .B1(n16597), .B2(n11970), .A(n11967), .ZN(n11705) );
  INV_X1 U13603 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n11700) );
  OAI22_X1 U13604 ( .A1(n11966), .A2(n13837), .B1(n16602), .B2(n11700), .ZN(
        n11701) );
  INV_X1 U13605 ( .A(n11701), .ZN(n11702) );
  OAI21_X1 U13606 ( .B1(n11705), .B2(n16605), .A(n11702), .ZN(P3_U3405) );
  INV_X1 U13607 ( .A(n13379), .ZN(n13341) );
  AOI22_X1 U13608 ( .A1(n13341), .A2(n11703), .B1(n16599), .B2(
        P3_REG1_REG_5__SCAN_IN), .ZN(n11704) );
  OAI21_X1 U13609 ( .B1(n11705), .B2(n16599), .A(n11704), .ZN(P3_U3464) );
  OAI222_X1 U13610 ( .A1(n14787), .A2(n11707), .B1(P2_U3088), .B2(n14286), 
        .C1(n14783), .C2(n11706), .ZN(P2_U3307) );
  INV_X1 U13611 ( .A(n11708), .ZN(n11710) );
  XNOR2_X1 U13612 ( .A(n14086), .B(n10884), .ZN(n11712) );
  AND2_X1 U13613 ( .A1(n14356), .A2(n7437), .ZN(n11713) );
  NAND2_X1 U13614 ( .A1(n11712), .A2(n11713), .ZN(n11716) );
  INV_X1 U13615 ( .A(n11712), .ZN(n11907) );
  INV_X1 U13616 ( .A(n11713), .ZN(n11714) );
  NAND2_X1 U13617 ( .A1(n11907), .A2(n11714), .ZN(n11715) );
  NAND2_X1 U13618 ( .A1(n11716), .A2(n11715), .ZN(n11881) );
  XNOR2_X1 U13619 ( .A(n14094), .B(n10884), .ZN(n11717) );
  NAND2_X1 U13620 ( .A1(n14355), .A2(n7437), .ZN(n11718) );
  XNOR2_X1 U13621 ( .A(n11717), .B(n11718), .ZN(n11910) );
  INV_X1 U13622 ( .A(n11717), .ZN(n11724) );
  NAND2_X1 U13623 ( .A1(n11724), .A2(n11718), .ZN(n11719) );
  XNOR2_X1 U13624 ( .A(n14101), .B(n7433), .ZN(n11888) );
  NAND2_X1 U13625 ( .A1(n14354), .A2(n7437), .ZN(n11889) );
  INV_X1 U13626 ( .A(n11899), .ZN(n11728) );
  NOR2_X1 U13627 ( .A1(n13902), .A2(n14096), .ZN(n11723) );
  NAND2_X1 U13628 ( .A1(n13904), .A2(n14353), .ZN(n11721) );
  OAI211_X1 U13629 ( .C1(n13970), .C2(n12091), .A(n11721), .B(n11720), .ZN(
        n11722) );
  AOI211_X1 U13630 ( .C1(n7765), .C2(n13983), .A(n11723), .B(n11722), .ZN(
        n11727) );
  OAI22_X1 U13631 ( .A1(n11724), .A2(n13963), .B1(n14096), .B2(n13976), .ZN(
        n11725) );
  NAND3_X1 U13632 ( .A1(n11915), .A2(n8171), .A3(n11725), .ZN(n11726) );
  OAI211_X1 U13633 ( .C1(n11728), .C2(n13963), .A(n11727), .B(n11726), .ZN(
        P2_U3206) );
  INV_X1 U13634 ( .A(n12740), .ZN(n11729) );
  NAND3_X1 U13635 ( .A1(n16353), .A2(n12600), .A3(n11729), .ZN(n11730) );
  NAND2_X1 U13636 ( .A1(n11731), .A2(n11730), .ZN(n16393) );
  OAI22_X1 U13637 ( .A1(n13304), .A2(n16390), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n16360), .ZN(n11743) );
  INV_X1 U13638 ( .A(n11733), .ZN(n11734) );
  NAND2_X1 U13639 ( .A1(n11732), .A2(n11734), .ZN(n11735) );
  NAND2_X1 U13640 ( .A1(n11735), .A2(n12740), .ZN(n11737) );
  NAND3_X1 U13641 ( .A1(n11737), .A2(n13299), .A3(n11736), .ZN(n11741) );
  OAI22_X1 U13642 ( .A1(n16314), .A2(n16350), .B1(n11738), .B2(n16352), .ZN(
        n11739) );
  INV_X1 U13643 ( .A(n11739), .ZN(n11740) );
  NAND2_X1 U13644 ( .A1(n11741), .A2(n11740), .ZN(n16391) );
  MUX2_X1 U13645 ( .A(n16391), .B(P3_REG2_REG_3__SCAN_IN), .S(n16369), .Z(
        n11742) );
  AOI211_X1 U13646 ( .C1(n13266), .C2(n16393), .A(n11743), .B(n11742), .ZN(
        n11744) );
  INV_X1 U13647 ( .A(n11744), .ZN(P3_U3230) );
  NAND2_X1 U13648 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n15377) );
  NAND2_X1 U13649 ( .A1(n15008), .A2(n15321), .ZN(n11746) );
  NAND2_X1 U13650 ( .A1(n15006), .A2(n15323), .ZN(n11745) );
  NAND2_X1 U13651 ( .A1(n11746), .A2(n11745), .ZN(n16482) );
  NAND2_X1 U13652 ( .A1(n16614), .A2(n16482), .ZN(n11747) );
  OAI211_X1 U13653 ( .C1(n16619), .C2(n16489), .A(n15377), .B(n11747), .ZN(
        n11762) );
  NAND2_X1 U13654 ( .A1(n11749), .A2(n11748), .ZN(n11754) );
  INV_X1 U13655 ( .A(n11750), .ZN(n11752) );
  NAND2_X1 U13656 ( .A1(n11752), .A2(n11751), .ZN(n11753) );
  NAND2_X1 U13657 ( .A1(n11754), .A2(n11753), .ZN(n11785) );
  NAND2_X1 U13658 ( .A1(n15074), .A2(n14917), .ZN(n11757) );
  NAND2_X1 U13659 ( .A1(n14916), .A2(n15322), .ZN(n11756) );
  NAND2_X1 U13660 ( .A1(n11757), .A2(n11756), .ZN(n11758) );
  XNOR2_X1 U13661 ( .A(n11758), .B(n14919), .ZN(n11788) );
  NOR2_X1 U13662 ( .A1(n14830), .A2(n11768), .ZN(n11759) );
  AOI21_X1 U13663 ( .B1(n15074), .B2(n14916), .A(n11759), .ZN(n11786) );
  XNOR2_X1 U13664 ( .A(n11788), .B(n11786), .ZN(n11784) );
  XNOR2_X1 U13665 ( .A(n11785), .B(n11784), .ZN(n11760) );
  NOR2_X1 U13666 ( .A1(n11760), .A2(n15029), .ZN(n11761) );
  AOI211_X1 U13667 ( .C1(n16610), .C2(n15074), .A(n11762), .B(n11761), .ZN(
        n11763) );
  INV_X1 U13668 ( .A(n11763), .ZN(P1_U3213) );
  OAI21_X1 U13669 ( .B1(n11764), .B2(n11767), .A(n11765), .ZN(n16515) );
  AOI21_X1 U13670 ( .B1(n11766), .B2(n11767), .A(n16479), .ZN(n11771) );
  OAI22_X1 U13671 ( .A1(n11768), .A2(n15293), .B1(n12039), .B2(n15016), .ZN(
        n11796) );
  NOR2_X1 U13672 ( .A1(n16515), .A2(n16370), .ZN(n11769) );
  AOI211_X1 U13673 ( .C1(n11771), .C2(n11770), .A(n11796), .B(n11769), .ZN(
        n16521) );
  INV_X1 U13674 ( .A(n11772), .ZN(n16474) );
  INV_X1 U13675 ( .A(n12003), .ZN(n11773) );
  AOI211_X1 U13676 ( .C1(n15078), .C2(n16474), .A(n16437), .B(n11773), .ZN(
        n16519) );
  AOI21_X1 U13677 ( .B1(n16573), .B2(n15078), .A(n16519), .ZN(n11774) );
  OAI211_X1 U13678 ( .C1(n16468), .C2(n16515), .A(n16521), .B(n11774), .ZN(
        n11776) );
  NAND2_X1 U13679 ( .A1(n11776), .A2(n7435), .ZN(n11775) );
  OAI21_X1 U13680 ( .B1(n7435), .B2(n9354), .A(n11775), .ZN(P1_U3536) );
  INV_X1 U13681 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11778) );
  NAND2_X1 U13682 ( .A1(n11776), .A2(n16540), .ZN(n11777) );
  OAI21_X1 U13683 ( .B1(n16540), .B2(n11778), .A(n11777), .ZN(P1_U3483) );
  NAND2_X1 U13684 ( .A1(n15078), .A2(n14917), .ZN(n11780) );
  NAND2_X1 U13685 ( .A1(n14916), .A2(n15321), .ZN(n11779) );
  NAND2_X1 U13686 ( .A1(n11780), .A2(n11779), .ZN(n11781) );
  XNOR2_X1 U13687 ( .A(n11781), .B(n14827), .ZN(n12033) );
  NOR2_X1 U13688 ( .A1(n14830), .A2(n11782), .ZN(n11783) );
  AOI21_X1 U13689 ( .B1(n15078), .B2(n14916), .A(n11783), .ZN(n12032) );
  XNOR2_X1 U13690 ( .A(n12033), .B(n12032), .ZN(n11795) );
  NAND2_X1 U13691 ( .A1(n11785), .A2(n11784), .ZN(n11790) );
  INV_X1 U13692 ( .A(n11786), .ZN(n11787) );
  NAND2_X1 U13693 ( .A1(n11788), .A2(n11787), .ZN(n11789) );
  NAND2_X1 U13694 ( .A1(n11790), .A2(n11789), .ZN(n11794) );
  INV_X1 U13695 ( .A(n11795), .ZN(n11791) );
  INV_X1 U13696 ( .A(n12035), .ZN(n11793) );
  AOI21_X1 U13697 ( .B1(n11795), .B2(n11794), .A(n11793), .ZN(n11801) );
  NAND2_X1 U13698 ( .A1(n16614), .A2(n11796), .ZN(n11797) );
  OAI211_X1 U13699 ( .C1(n16619), .C2(n16507), .A(n11798), .B(n11797), .ZN(
        n11799) );
  AOI21_X1 U13700 ( .B1(n16610), .B2(n15078), .A(n11799), .ZN(n11800) );
  OAI21_X1 U13701 ( .B1(n11801), .B2(n15029), .A(n11800), .ZN(P1_U3221) );
  NAND2_X1 U13702 ( .A1(n11803), .A2(n11802), .ZN(n12336) );
  XNOR2_X1 U13703 ( .A(n12336), .B(n11815), .ZN(n11804) );
  NAND2_X1 U13704 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n11804), .ZN(n12337) );
  OAI211_X1 U13705 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n11804), .A(n15877), 
        .B(n12337), .ZN(n11811) );
  OAI22_X1 U13706 ( .A1(n11808), .A2(n11807), .B1(n11806), .B2(n11805), .ZN(
        n12348) );
  XNOR2_X1 U13707 ( .A(n11815), .B(n12348), .ZN(n11809) );
  NAND2_X1 U13708 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n11809), .ZN(n12350) );
  OAI211_X1 U13709 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n11809), .A(n15873), 
        .B(n12350), .ZN(n11810) );
  NAND2_X1 U13710 ( .A1(n11811), .A2(n11810), .ZN(n11813) );
  NAND2_X1 U13711 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n12388)
         );
  INV_X1 U13712 ( .A(n12388), .ZN(n11812) );
  AOI211_X1 U13713 ( .C1(n15875), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n11813), 
        .B(n11812), .ZN(n11814) );
  OAI21_X1 U13714 ( .B1(n11815), .B2(n15842), .A(n11814), .ZN(P2_U3229) );
  NOR2_X1 U13715 ( .A1(n11817), .A2(n11816), .ZN(n11819) );
  INV_X1 U13716 ( .A(n11834), .ZN(n13044) );
  NAND2_X1 U13717 ( .A1(n13044), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n13012) );
  INV_X1 U13718 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11820) );
  NAND2_X1 U13719 ( .A1(n11834), .A2(n11820), .ZN(n11821) );
  NAND2_X1 U13720 ( .A1(n13012), .A2(n11821), .ZN(n11823) );
  INV_X1 U13721 ( .A(n13013), .ZN(n11822) );
  AOI21_X1 U13722 ( .B1(n11824), .B2(n11823), .A(n11822), .ZN(n11844) );
  AOI21_X1 U13723 ( .B1(n11826), .B2(n11831), .A(n11825), .ZN(n11828) );
  MUX2_X1 U13724 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13036), .Z(n13026) );
  XNOR2_X1 U13725 ( .A(n13026), .B(n11834), .ZN(n11827) );
  NAND2_X1 U13726 ( .A1(n11828), .A2(n11827), .ZN(n13025) );
  OAI21_X1 U13727 ( .B1(n11828), .B2(n11827), .A(n13025), .ZN(n11829) );
  NAND2_X1 U13728 ( .A1(n11829), .A2(n16195), .ZN(n11843) );
  NAND2_X1 U13729 ( .A1(n11831), .A2(n11830), .ZN(n11833) );
  NAND2_X1 U13730 ( .A1(n11833), .A2(n11832), .ZN(n11838) );
  INV_X1 U13731 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11835) );
  MUX2_X1 U13732 ( .A(P3_REG2_REG_10__SCAN_IN), .B(n11835), .S(n11834), .Z(
        n11836) );
  INV_X1 U13733 ( .A(n11836), .ZN(n11837) );
  NAND2_X1 U13734 ( .A1(n11837), .A2(n11838), .ZN(n13045) );
  OAI21_X1 U13735 ( .B1(n11838), .B2(n11837), .A(n13045), .ZN(n11841) );
  NAND2_X1 U13736 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n12207)
         );
  NAND2_X1 U13737 ( .A1(n16259), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n11839) );
  OAI211_X1 U13738 ( .C1(n16142), .C2(n13044), .A(n12207), .B(n11839), .ZN(
        n11840) );
  AOI21_X1 U13739 ( .B1(n11841), .B2(n16194), .A(n11840), .ZN(n11842) );
  OAI211_X1 U13740 ( .C1(n11844), .C2(n16274), .A(n11843), .B(n11842), .ZN(
        P3_U3192) );
  OAI21_X1 U13741 ( .B1(n11846), .B2(n12624), .A(n11845), .ZN(n11858) );
  INV_X1 U13742 ( .A(n11858), .ZN(n11855) );
  XNOR2_X1 U13743 ( .A(n11847), .B(n12624), .ZN(n11850) );
  NAND2_X1 U13744 ( .A1(n12995), .A2(n12975), .ZN(n11848) );
  OAI21_X1 U13745 ( .B1(n12140), .B2(n16352), .A(n11848), .ZN(n11849) );
  AOI21_X1 U13746 ( .B1(n11850), .B2(n13299), .A(n11849), .ZN(n11856) );
  MUX2_X1 U13747 ( .A(n11856), .B(n11851), .S(n16369), .Z(n11854) );
  AOI22_X1 U13748 ( .A1(n13260), .A2(n11859), .B1(n13291), .B2(n11852), .ZN(
        n11853) );
  OAI211_X1 U13749 ( .C1(n11855), .C2(n13313), .A(n11854), .B(n11853), .ZN(
        P3_U3226) );
  INV_X1 U13750 ( .A(n11856), .ZN(n11857) );
  AOI21_X1 U13751 ( .B1(n16597), .B2(n11858), .A(n11857), .ZN(n11865) );
  AOI22_X1 U13752 ( .A1(n13341), .A2(n11859), .B1(n16599), .B2(
        P3_REG1_REG_7__SCAN_IN), .ZN(n11860) );
  OAI21_X1 U13753 ( .B1(n11865), .B2(n16599), .A(n11860), .ZN(P3_U3466) );
  INV_X1 U13754 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n11861) );
  OAI22_X1 U13755 ( .A1(n11862), .A2(n13837), .B1(n16602), .B2(n11861), .ZN(
        n11863) );
  INV_X1 U13756 ( .A(n11863), .ZN(n11864) );
  OAI21_X1 U13757 ( .B1(n11865), .B2(n16605), .A(n11864), .ZN(P3_U3411) );
  OAI21_X1 U13758 ( .B1(n11867), .B2(n12744), .A(n11866), .ZN(n11868) );
  AOI222_X1 U13759 ( .A1(n13299), .A2(n11868), .B1(n12992), .B2(n13251), .C1(
        n12994), .C2(n12975), .ZN(n16504) );
  OAI21_X1 U13760 ( .B1(n11870), .B2(n12629), .A(n11869), .ZN(n16502) );
  NOR2_X1 U13761 ( .A1(n13307), .A2(n11529), .ZN(n11873) );
  OAI22_X1 U13762 ( .A1(n13304), .A2(n11871), .B1(n12027), .B2(n16360), .ZN(
        n11872) );
  AOI211_X1 U13763 ( .C1(n16502), .C2(n13266), .A(n11873), .B(n11872), .ZN(
        n11874) );
  OAI21_X1 U13764 ( .B1(n16504), .B2(n16369), .A(n11874), .ZN(P3_U3225) );
  INV_X1 U13765 ( .A(n11875), .ZN(n11876) );
  AOI22_X1 U13766 ( .A1(n13985), .A2(n11876), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11877) );
  OAI21_X1 U13767 ( .B1(n13988), .B2(n11878), .A(n11877), .ZN(n11883) );
  INV_X1 U13768 ( .A(n11879), .ZN(n11909) );
  AOI211_X1 U13769 ( .C1(n11881), .C2(n11880), .A(n13963), .B(n11909), .ZN(
        n11882) );
  AOI211_X1 U13770 ( .C1(n14086), .C2(n13983), .A(n11883), .B(n11882), .ZN(
        n11884) );
  INV_X1 U13771 ( .A(n11884), .ZN(P2_U3208) );
  INV_X1 U13772 ( .A(n11885), .ZN(n11886) );
  OAI222_X1 U13773 ( .A1(P3_U3151), .A2(n11887), .B1(n13853), .B2(n11886), 
        .C1(n13610), .C2(n13850), .ZN(P3_U3270) );
  INV_X1 U13774 ( .A(n11888), .ZN(n11896) );
  INV_X1 U13775 ( .A(n11889), .ZN(n11890) );
  XNOR2_X1 U13776 ( .A(n14725), .B(n10884), .ZN(n12306) );
  NAND2_X1 U13777 ( .A1(n14353), .A2(n7437), .ZN(n12304) );
  XNOR2_X1 U13778 ( .A(n12306), .B(n12304), .ZN(n11897) );
  NOR2_X1 U13779 ( .A1(n13902), .A2(n11891), .ZN(n11895) );
  NAND2_X1 U13780 ( .A1(n13904), .A2(n14352), .ZN(n11893) );
  OAI211_X1 U13781 ( .C1(n13970), .C2(n12279), .A(n11893), .B(n11892), .ZN(
        n11894) );
  AOI211_X1 U13782 ( .C1(n14725), .C2(n13983), .A(n11895), .B(n11894), .ZN(
        n11901) );
  AOI22_X1 U13783 ( .A1(n11896), .A2(n13990), .B1(n13894), .B2(n14354), .ZN(
        n11898) );
  OR3_X1 U13784 ( .A1(n11899), .A2(n11898), .A3(n11897), .ZN(n11900) );
  OAI211_X1 U13785 ( .C1(n12305), .C2(n13963), .A(n11901), .B(n11900), .ZN(
        P2_U3187) );
  NAND2_X1 U13786 ( .A1(n14354), .A2(n14589), .ZN(n11903) );
  NAND2_X1 U13787 ( .A1(n14356), .A2(n14588), .ZN(n11902) );
  AND2_X1 U13788 ( .A1(n11903), .A2(n11902), .ZN(n11944) );
  INV_X1 U13789 ( .A(n11904), .ZN(n11948) );
  AOI22_X1 U13790 ( .A1(n13985), .A2(n11948), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11905) );
  OAI21_X1 U13791 ( .B1(n13988), .B2(n11944), .A(n11905), .ZN(n11913) );
  NOR3_X1 U13792 ( .A1(n11907), .A2(n11906), .A3(n13976), .ZN(n11908) );
  AOI21_X1 U13793 ( .B1(n11909), .B2(n13990), .A(n11908), .ZN(n11911) );
  NOR2_X1 U13794 ( .A1(n11911), .A2(n11910), .ZN(n11912) );
  AOI211_X1 U13795 ( .C1(n14094), .C2(n13983), .A(n11913), .B(n11912), .ZN(
        n11914) );
  OAI21_X1 U13796 ( .B1(n13963), .B2(n11915), .A(n11914), .ZN(P2_U3196) );
  INV_X1 U13797 ( .A(n12745), .ZN(n11916) );
  NAND3_X1 U13798 ( .A1(n11917), .A2(n11916), .A3(n12616), .ZN(n11918) );
  NAND2_X1 U13799 ( .A1(n11919), .A2(n11918), .ZN(n16461) );
  OAI22_X1 U13800 ( .A1(n13304), .A2(n16458), .B1(n11920), .B2(n16360), .ZN(
        n11931) );
  INV_X1 U13801 ( .A(n11921), .ZN(n11922) );
  NAND2_X1 U13802 ( .A1(n11696), .A2(n11922), .ZN(n11923) );
  NAND2_X1 U13803 ( .A1(n11923), .A2(n12745), .ZN(n11925) );
  NAND3_X1 U13804 ( .A1(n11925), .A2(n13299), .A3(n11924), .ZN(n11929) );
  OAI22_X1 U13805 ( .A1(n12022), .A2(n16352), .B1(n11926), .B2(n16350), .ZN(
        n11927) );
  INV_X1 U13806 ( .A(n11927), .ZN(n11928) );
  NAND2_X1 U13807 ( .A1(n11929), .A2(n11928), .ZN(n16459) );
  MUX2_X1 U13808 ( .A(n16459), .B(P3_REG2_REG_6__SCAN_IN), .S(n16369), .Z(
        n11930) );
  AOI211_X1 U13809 ( .C1(n13266), .C2(n16461), .A(n11931), .B(n11930), .ZN(
        n11932) );
  INV_X1 U13810 ( .A(n11932), .ZN(P3_U3227) );
  AOI211_X1 U13811 ( .C1(n14717), .C2(n11935), .A(n11934), .B(n11933), .ZN(
        n11940) );
  NOR2_X1 U13812 ( .A1(n11936), .A2(n8761), .ZN(n11937) );
  AOI21_X1 U13813 ( .B1(n14086), .B2(n9744), .A(n11937), .ZN(n11938) );
  OAI21_X1 U13814 ( .B1(n11940), .B2(n16561), .A(n11938), .ZN(P2_U3463) );
  AOI22_X1 U13815 ( .A1(n14086), .A2(n12239), .B1(n16559), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11939) );
  OAI21_X1 U13816 ( .B1(n11940), .B2(n16559), .A(n11939), .ZN(P2_U3510) );
  XOR2_X1 U13817 ( .A(n11941), .B(n14301), .Z(n12100) );
  INV_X1 U13818 ( .A(n12100), .ZN(n11953) );
  INV_X1 U13819 ( .A(n14301), .ZN(n11943) );
  OAI211_X1 U13820 ( .C1(n7606), .C2(n11943), .A(n11942), .B(n14606), .ZN(
        n11945) );
  NAND2_X1 U13821 ( .A1(n11945), .A2(n11944), .ZN(n12098) );
  INV_X1 U13822 ( .A(n12089), .ZN(n11946) );
  AOI211_X1 U13823 ( .C1(n14094), .C2(n11947), .A(n7437), .B(n11946), .ZN(
        n12099) );
  NAND2_X1 U13824 ( .A1(n12099), .A2(n14632), .ZN(n11950) );
  INV_X1 U13825 ( .A(n14624), .ZN(n14615) );
  AOI22_X1 U13826 ( .A1(n14622), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11948), 
        .B2(n14615), .ZN(n11949) );
  OAI211_X1 U13827 ( .C1(n9108), .C2(n14619), .A(n11950), .B(n11949), .ZN(
        n11951) );
  AOI21_X1 U13828 ( .B1(n11368), .B2(n12098), .A(n11951), .ZN(n11952) );
  OAI21_X1 U13829 ( .B1(n14580), .B2(n11953), .A(n11952), .ZN(P2_U3253) );
  OAI21_X1 U13830 ( .B1(n11955), .B2(n15245), .A(n11954), .ZN(n12075) );
  INV_X1 U13831 ( .A(n12075), .ZN(n11960) );
  NAND2_X1 U13832 ( .A1(n15008), .A2(n15318), .ZN(n12067) );
  NAND2_X1 U13833 ( .A1(n15006), .A2(n15320), .ZN(n12076) );
  NAND2_X1 U13834 ( .A1(n12067), .A2(n12076), .ZN(n12050) );
  INV_X1 U13835 ( .A(n12182), .ZN(n11956) );
  AOI211_X1 U13836 ( .C1(n15090), .C2(n7612), .A(n16437), .B(n11956), .ZN(
        n12068) );
  AOI211_X1 U13837 ( .C1(n16573), .C2(n15090), .A(n12050), .B(n12068), .ZN(
        n11959) );
  XNOR2_X1 U13838 ( .A(n11957), .B(n15245), .ZN(n11958) );
  NAND2_X1 U13839 ( .A1(n11958), .A2(n16536), .ZN(n12077) );
  OAI211_X1 U13840 ( .C1(n16576), .C2(n11960), .A(n11959), .B(n12077), .ZN(
        n11962) );
  NAND2_X1 U13841 ( .A1(n11962), .A2(n7435), .ZN(n11961) );
  OAI21_X1 U13842 ( .B1(n7435), .B2(n9387), .A(n11961), .ZN(P1_U3538) );
  INV_X1 U13843 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n11964) );
  NAND2_X1 U13844 ( .A1(n11962), .A2(n16540), .ZN(n11963) );
  OAI21_X1 U13845 ( .B1(n16540), .B2(n11964), .A(n11963), .ZN(P1_U3489) );
  OAI22_X1 U13846 ( .A1(n13304), .A2(n11966), .B1(n11965), .B2(n16360), .ZN(
        n11969) );
  MUX2_X1 U13847 ( .A(P3_REG2_REG_5__SCAN_IN), .B(n11967), .S(n13307), .Z(
        n11968) );
  AOI211_X1 U13848 ( .C1(n13266), .C2(n11970), .A(n11969), .B(n11968), .ZN(
        n11971) );
  INV_X1 U13849 ( .A(n11971), .ZN(P3_U3228) );
  INV_X1 U13850 ( .A(n16370), .ZN(n16483) );
  AOI21_X1 U13851 ( .B1(n16483), .B2(n15515), .A(n16513), .ZN(n15608) );
  XOR2_X1 U13852 ( .A(n11972), .B(n15238), .Z(n16469) );
  OAI21_X1 U13853 ( .B1(n11974), .B2(n9333), .A(n11973), .ZN(n11976) );
  AOI21_X1 U13854 ( .B1(n11976), .B2(n16536), .A(n11975), .ZN(n16467) );
  MUX2_X1 U13855 ( .A(n10571), .B(n16467), .S(n15515), .Z(n11982) );
  AOI211_X1 U13856 ( .C1(n16465), .C2(n16439), .A(n16437), .B(n16475), .ZN(
        n16464) );
  NAND2_X1 U13857 ( .A1(n11977), .A2(n15217), .ZN(n11978) );
  OAI22_X1 U13858 ( .A1(n16512), .A2(n7436), .B1(n16490), .B2(n11979), .ZN(
        n11980) );
  AOI21_X1 U13859 ( .B1(n16518), .B2(n16464), .A(n11980), .ZN(n11981) );
  OAI211_X1 U13860 ( .C1(n15608), .C2(n16469), .A(n11982), .B(n11981), .ZN(
        P1_U3287) );
  INV_X1 U13861 ( .A(n11983), .ZN(n11984) );
  OAI222_X1 U13862 ( .A1(n14787), .A2(n11985), .B1(n14783), .B2(n11984), .C1(
        n8539), .C2(P2_U3088), .ZN(P2_U3305) );
  OAI21_X1 U13863 ( .B1(n11988), .B2(n11987), .A(n11986), .ZN(n11990) );
  AOI21_X1 U13864 ( .B1(n11990), .B2(n16536), .A(n11989), .ZN(n16373) );
  NAND2_X1 U13865 ( .A1(n16522), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n11991) );
  OAI21_X1 U13866 ( .B1(n16490), .B2(n11992), .A(n11991), .ZN(n11995) );
  INV_X1 U13867 ( .A(n16518), .ZN(n15621) );
  NAND2_X1 U13868 ( .A1(n16329), .A2(n7812), .ZN(n11993) );
  NAND3_X1 U13869 ( .A1(n12107), .A2(n16473), .A3(n11993), .ZN(n16372) );
  NOR2_X1 U13870 ( .A1(n15621), .A2(n16372), .ZN(n11994) );
  AOI211_X1 U13871 ( .C1(n15619), .C2(n7812), .A(n11995), .B(n11994), .ZN(
        n11999) );
  INV_X1 U13872 ( .A(n15608), .ZN(n11997) );
  XNOR2_X1 U13873 ( .A(n11996), .B(n15234), .ZN(n16377) );
  NAND2_X1 U13874 ( .A1(n11997), .A2(n16377), .ZN(n11998) );
  OAI211_X1 U13875 ( .C1(n16522), .C2(n16373), .A(n11999), .B(n11998), .ZN(
        P1_U3291) );
  INV_X1 U13876 ( .A(n12001), .ZN(n12002) );
  AOI21_X1 U13877 ( .B1(n15241), .B2(n12000), .A(n12002), .ZN(n16534) );
  AOI21_X1 U13878 ( .B1(n16531), .B2(n12003), .A(n16437), .ZN(n12004) );
  NAND2_X1 U13879 ( .A1(n12004), .A2(n7612), .ZN(n16532) );
  INV_X1 U13880 ( .A(n16532), .ZN(n12012) );
  INV_X1 U13881 ( .A(n16531), .ZN(n12010) );
  NAND2_X1 U13882 ( .A1(n15008), .A2(n15319), .ZN(n12006) );
  NAND2_X1 U13883 ( .A1(n15006), .A2(n15321), .ZN(n12005) );
  NAND2_X1 U13884 ( .A1(n12006), .A2(n12005), .ZN(n16530) );
  INV_X1 U13885 ( .A(n16530), .ZN(n12007) );
  OAI22_X1 U13886 ( .A1(n16522), .A2(n12007), .B1(n12215), .B2(n16490), .ZN(
        n12008) );
  AOI21_X1 U13887 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n16522), .A(n12008), .ZN(
        n12009) );
  OAI21_X1 U13888 ( .B1(n12010), .B2(n16512), .A(n12009), .ZN(n12011) );
  AOI21_X1 U13889 ( .B1(n16518), .B2(n12012), .A(n12011), .ZN(n12015) );
  XOR2_X1 U13890 ( .A(n12013), .B(n15241), .Z(n16537) );
  NOR2_X1 U13891 ( .A1(n16522), .A2(n16479), .ZN(n15537) );
  NAND2_X1 U13892 ( .A1(n16537), .A2(n15537), .ZN(n12014) );
  OAI211_X1 U13893 ( .C1(n16534), .C2(n15608), .A(n12015), .B(n12014), .ZN(
        P1_U3284) );
  XNOR2_X1 U13894 ( .A(n16501), .B(n11080), .ZN(n12134) );
  XNOR2_X1 U13895 ( .A(n12140), .B(n12134), .ZN(n12135) );
  INV_X1 U13896 ( .A(n12016), .ZN(n12020) );
  OAI21_X1 U13897 ( .B1(n12022), .B2(n12020), .A(n12019), .ZN(n12136) );
  XOR2_X1 U13898 ( .A(n12135), .B(n12136), .Z(n12021) );
  NAND2_X1 U13899 ( .A1(n12021), .A2(n7876), .ZN(n12026) );
  OAI22_X1 U13900 ( .A1(n12141), .A2(n12022), .B1(n12133), .B2(n12954), .ZN(
        n12023) );
  AOI211_X1 U13901 ( .C1(n16501), .C2(n12966), .A(n12024), .B(n12023), .ZN(
        n12025) );
  OAI211_X1 U13902 ( .C1(n12027), .C2(n12955), .A(n12026), .B(n12025), .ZN(
        P3_U3161) );
  INV_X1 U13903 ( .A(n12028), .ZN(n12029) );
  OAI222_X1 U13904 ( .A1(n12031), .A2(P3_U3151), .B1(n13850), .B2(n12030), 
        .C1(n13853), .C2(n12029), .ZN(P3_U3269) );
  NAND2_X1 U13905 ( .A1(n12033), .A2(n12032), .ZN(n12034) );
  NAND2_X1 U13906 ( .A1(n16531), .A2(n14917), .ZN(n12037) );
  NAND2_X1 U13907 ( .A1(n14916), .A2(n15320), .ZN(n12036) );
  NAND2_X1 U13908 ( .A1(n12037), .A2(n12036), .ZN(n12038) );
  XNOR2_X1 U13909 ( .A(n12038), .B(n14827), .ZN(n12041) );
  NOR2_X1 U13910 ( .A1(n14830), .A2(n12039), .ZN(n12040) );
  AOI21_X1 U13911 ( .B1(n16531), .B2(n14916), .A(n12040), .ZN(n12042) );
  XNOR2_X1 U13912 ( .A(n12041), .B(n12042), .ZN(n12217) );
  INV_X1 U13913 ( .A(n12041), .ZN(n12044) );
  INV_X1 U13914 ( .A(n12042), .ZN(n12043) );
  NAND2_X1 U13915 ( .A1(n15090), .A2(n14917), .ZN(n12046) );
  NAND2_X1 U13916 ( .A1(n14916), .A2(n15319), .ZN(n12045) );
  NAND2_X1 U13917 ( .A1(n12046), .A2(n12045), .ZN(n12047) );
  XNOR2_X1 U13918 ( .A(n12047), .B(n14919), .ZN(n12250) );
  NOR2_X1 U13919 ( .A1(n14830), .A2(n12048), .ZN(n12049) );
  AOI21_X1 U13920 ( .B1(n15090), .B2(n14916), .A(n12049), .ZN(n12248) );
  XNOR2_X1 U13921 ( .A(n12250), .B(n12248), .ZN(n12251) );
  XNOR2_X1 U13922 ( .A(n12252), .B(n12251), .ZN(n12055) );
  NAND2_X1 U13923 ( .A1(n16614), .A2(n12050), .ZN(n12051) );
  OAI211_X1 U13924 ( .C1(n16619), .C2(n12071), .A(n12052), .B(n12051), .ZN(
        n12053) );
  AOI21_X1 U13925 ( .B1(n16610), .B2(n15090), .A(n12053), .ZN(n12054) );
  OAI21_X1 U13926 ( .B1(n12055), .B2(n15029), .A(n12054), .ZN(P1_U3217) );
  XNOR2_X1 U13927 ( .A(n12056), .B(n15236), .ZN(n16421) );
  INV_X1 U13928 ( .A(n12070), .ZN(n12057) );
  OAI211_X1 U13929 ( .C1(n12110), .C2(n15055), .A(n16473), .B(n16438), .ZN(
        n16426) );
  NOR2_X1 U13930 ( .A1(n15621), .A2(n16426), .ZN(n12063) );
  NOR2_X1 U13931 ( .A1(n16512), .A2(n15055), .ZN(n12062) );
  AND2_X1 U13932 ( .A1(n16522), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n12061) );
  INV_X1 U13933 ( .A(n16424), .ZN(n12059) );
  OAI22_X1 U13934 ( .A1(n16522), .A2(n12059), .B1(n12058), .B2(n16490), .ZN(
        n12060) );
  NOR4_X1 U13935 ( .A1(n12063), .A2(n12062), .A3(n12061), .A4(n12060), .ZN(
        n12066) );
  OR2_X1 U13936 ( .A1(n12064), .A2(n15236), .ZN(n16423) );
  NAND3_X1 U13937 ( .A1(n15537), .A2(n16422), .A3(n16423), .ZN(n12065) );
  OAI211_X1 U13938 ( .C1(n16421), .C2(n15592), .A(n12066), .B(n12065), .ZN(
        P1_U3289) );
  INV_X1 U13939 ( .A(n12067), .ZN(n12069) );
  AOI211_X1 U13940 ( .C1(n12075), .C2(n12070), .A(n12069), .B(n12068), .ZN(
        n12081) );
  NOR2_X1 U13941 ( .A1(n9626), .A2(n16512), .ZN(n12074) );
  OAI22_X1 U13942 ( .A1(n15515), .A2(n12072), .B1(n12071), .B2(n16490), .ZN(
        n12073) );
  AOI211_X1 U13943 ( .C1(n12075), .C2(n16513), .A(n12074), .B(n12073), .ZN(
        n12080) );
  AOI21_X1 U13944 ( .B1(n12077), .B2(n12076), .A(n16522), .ZN(n12078) );
  INV_X1 U13945 ( .A(n12078), .ZN(n12079) );
  OAI211_X1 U13946 ( .C1(n12081), .C2(n15621), .A(n12080), .B(n12079), .ZN(
        P1_U3283) );
  OAI21_X1 U13947 ( .B1(n12083), .B2(n14302), .A(n12082), .ZN(n12238) );
  INV_X1 U13948 ( .A(n12238), .ZN(n12097) );
  XNOR2_X1 U13949 ( .A(n12085), .B(n12084), .ZN(n12088) );
  OAI22_X1 U13950 ( .A1(n14096), .A2(n13967), .B1(n14107), .B2(n13968), .ZN(
        n12086) );
  AOI21_X1 U13951 ( .B1(n12238), .B2(n14591), .A(n12086), .ZN(n12087) );
  OAI21_X1 U13952 ( .B1(n9148), .B2(n12088), .A(n12087), .ZN(n12236) );
  NAND2_X1 U13953 ( .A1(n12236), .A2(n11368), .ZN(n12096) );
  AOI211_X1 U13954 ( .C1(n7765), .C2(n12089), .A(n7437), .B(n7969), .ZN(n12237) );
  NOR2_X1 U13955 ( .A1(n12090), .A2(n14619), .ZN(n12094) );
  OAI22_X1 U13956 ( .A1(n11368), .A2(n12092), .B1(n12091), .B2(n14624), .ZN(
        n12093) );
  AOI211_X1 U13957 ( .C1(n12237), .C2(n14632), .A(n12094), .B(n12093), .ZN(
        n12095) );
  OAI211_X1 U13958 ( .C1(n12097), .C2(n14602), .A(n12096), .B(n12095), .ZN(
        P2_U3252) );
  AOI211_X1 U13959 ( .C1(n14717), .C2(n12100), .A(n12099), .B(n12098), .ZN(
        n12103) );
  AOI22_X1 U13960 ( .A1(n14094), .A2(n12239), .B1(P2_REG1_REG_12__SCAN_IN), 
        .B2(n16559), .ZN(n12101) );
  OAI21_X1 U13961 ( .B1(n12103), .B2(n16559), .A(n12101), .ZN(P2_U3511) );
  AOI22_X1 U13962 ( .A1(n14094), .A2(n9744), .B1(P2_REG0_REG_12__SCAN_IN), 
        .B2(n16561), .ZN(n12102) );
  OAI21_X1 U13963 ( .B1(n12103), .B2(n16561), .A(n12102), .ZN(P2_U3466) );
  INV_X1 U13964 ( .A(n12104), .ZN(n12190) );
  AOI22_X1 U13965 ( .A1(n9704), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n15763), .ZN(n12105) );
  OAI21_X1 U13966 ( .B1(n12190), .B2(n15780), .A(n12105), .ZN(P1_U3331) );
  XNOR2_X1 U13967 ( .A(n15235), .B(n12106), .ZN(n16404) );
  NAND2_X1 U13968 ( .A1(n12107), .A2(n16396), .ZN(n12108) );
  NAND2_X1 U13969 ( .A1(n12108), .A2(n16473), .ZN(n12109) );
  NOR2_X1 U13970 ( .A1(n12110), .A2(n12109), .ZN(n16408) );
  OR2_X1 U13971 ( .A1(n15056), .A2(n15016), .ZN(n12112) );
  NAND2_X1 U13972 ( .A1(n15006), .A2(n9639), .ZN(n12111) );
  NAND2_X1 U13973 ( .A1(n12112), .A2(n12111), .ZN(n16406) );
  MUX2_X1 U13974 ( .A(n16406), .B(P1_REG2_REG_3__SCAN_IN), .S(n16522), .Z(
        n12114) );
  OAI22_X1 U13975 ( .A1(n16512), .A2(n9625), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n16490), .ZN(n12113) );
  AOI211_X1 U13976 ( .C1(n16408), .C2(n16518), .A(n12114), .B(n12113), .ZN(
        n12117) );
  XNOR2_X1 U13977 ( .A(n12115), .B(n15235), .ZN(n16405) );
  NAND2_X1 U13978 ( .A1(n15537), .A2(n16405), .ZN(n12116) );
  OAI211_X1 U13979 ( .C1(n16404), .C2(n15592), .A(n12117), .B(n12116), .ZN(
        P1_U3290) );
  INV_X1 U13980 ( .A(n12149), .ZN(n12120) );
  AOI21_X1 U13981 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n15763), .A(n12118), 
        .ZN(n12119) );
  OAI21_X1 U13982 ( .B1(n12120), .B2(n15780), .A(n12119), .ZN(P1_U3332) );
  INV_X1 U13983 ( .A(n12121), .ZN(n12636) );
  AND2_X1 U13984 ( .A1(n12636), .A2(n12635), .ZN(n12741) );
  XOR2_X1 U13985 ( .A(n12122), .B(n12741), .Z(n16524) );
  INV_X1 U13986 ( .A(n12123), .ZN(n12124) );
  AND2_X1 U13987 ( .A1(n13310), .A2(n12124), .ZN(n13197) );
  INV_X1 U13988 ( .A(n13197), .ZN(n12132) );
  XOR2_X1 U13989 ( .A(n12125), .B(n12741), .Z(n12127) );
  OAI22_X1 U13990 ( .A1(n12229), .A2(n16352), .B1(n12140), .B2(n16350), .ZN(
        n12126) );
  AOI21_X1 U13991 ( .B1(n12127), .B2(n13299), .A(n12126), .ZN(n12128) );
  OAI21_X1 U13992 ( .B1(n16524), .B2(n16541), .A(n12128), .ZN(n16526) );
  NAND2_X1 U13993 ( .A1(n16526), .A2(n13310), .ZN(n12131) );
  OAI22_X1 U13994 ( .A1(n13304), .A2(n16523), .B1(n12147), .B2(n16360), .ZN(
        n12129) );
  AOI21_X1 U13995 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n16369), .A(n12129), .ZN(
        n12130) );
  OAI211_X1 U13996 ( .C1(n16524), .C2(n12132), .A(n12131), .B(n12130), .ZN(
        P3_U3224) );
  XNOR2_X1 U13997 ( .A(n16523), .B(n12821), .ZN(n12199) );
  XNOR2_X1 U13998 ( .A(n12133), .B(n12199), .ZN(n12138) );
  OAI21_X1 U13999 ( .B1(n12138), .B2(n12137), .A(n12204), .ZN(n12139) );
  NAND2_X1 U14000 ( .A1(n12139), .A2(n7876), .ZN(n12146) );
  OAI22_X1 U14001 ( .A1(n12141), .A2(n12140), .B1(n12229), .B2(n12954), .ZN(
        n12142) );
  AOI211_X1 U14002 ( .C1(n12144), .C2(n12966), .A(n12143), .B(n12142), .ZN(
        n12145) );
  OAI211_X1 U14003 ( .C1(n12147), .C2(n12955), .A(n12146), .B(n12145), .ZN(
        P3_U3171) );
  NAND2_X1 U14004 ( .A1(n12149), .A2(n12148), .ZN(n12151) );
  AND2_X1 U14005 ( .A1(n12150), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14282) );
  INV_X1 U14006 ( .A(n14282), .ZN(n14327) );
  OAI211_X1 U14007 ( .C1(n12152), .C2(n14787), .A(n12151), .B(n14327), .ZN(
        P2_U3304) );
  OAI21_X1 U14008 ( .B1(n12154), .B2(n15246), .A(n12153), .ZN(n12325) );
  INV_X1 U14009 ( .A(n12325), .ZN(n12169) );
  NAND2_X1 U14010 ( .A1(n15101), .A2(n12183), .ZN(n12155) );
  NAND2_X1 U14011 ( .A1(n12155), .A2(n16473), .ZN(n12156) );
  OR2_X1 U14012 ( .A1(n12291), .A2(n12156), .ZN(n12327) );
  INV_X1 U14013 ( .A(n12327), .ZN(n12164) );
  INV_X1 U14014 ( .A(n15101), .ZN(n12162) );
  NAND2_X1 U14015 ( .A1(n15008), .A2(n15316), .ZN(n12158) );
  NAND2_X1 U14016 ( .A1(n15006), .A2(n15318), .ZN(n12157) );
  NAND2_X1 U14017 ( .A1(n12158), .A2(n12157), .ZN(n14940) );
  INV_X1 U14018 ( .A(n14940), .ZN(n12159) );
  OAI22_X1 U14019 ( .A1(n16522), .A2(n12159), .B1(n14942), .B2(n16490), .ZN(
        n12160) );
  AOI21_X1 U14020 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n16522), .A(n12160), 
        .ZN(n12161) );
  OAI21_X1 U14021 ( .B1(n12162), .B2(n16512), .A(n12161), .ZN(n12163) );
  AOI21_X1 U14022 ( .B1(n12164), .B2(n16518), .A(n12163), .ZN(n12168) );
  NAND2_X1 U14023 ( .A1(n12166), .A2(n15246), .ZN(n12326) );
  NAND3_X1 U14024 ( .A1(n12165), .A2(n12326), .A3(n15537), .ZN(n12167) );
  OAI211_X1 U14025 ( .C1(n12169), .C2(n15608), .A(n12168), .B(n12167), .ZN(
        P1_U3281) );
  INV_X1 U14026 ( .A(n12170), .ZN(n12172) );
  OAI222_X1 U14027 ( .A1(n13036), .A2(P3_U3151), .B1(n13853), .B2(n12172), 
        .C1(n12171), .C2(n13850), .ZN(P3_U3268) );
  XNOR2_X1 U14028 ( .A(n12173), .B(n12178), .ZN(n12176) );
  NAND2_X1 U14029 ( .A1(n15008), .A2(n15317), .ZN(n12175) );
  NAND2_X1 U14030 ( .A1(n15006), .A2(n15319), .ZN(n12174) );
  NAND2_X1 U14031 ( .A1(n12175), .A2(n12174), .ZN(n12260) );
  AOI21_X1 U14032 ( .B1(n12176), .B2(n16536), .A(n12260), .ZN(n16575) );
  OAI21_X1 U14033 ( .B1(n12179), .B2(n12178), .A(n12177), .ZN(n16577) );
  NAND2_X1 U14034 ( .A1(n16522), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n12180) );
  OAI21_X1 U14035 ( .B1(n16490), .B2(n12257), .A(n12180), .ZN(n12181) );
  AOI21_X1 U14036 ( .B1(n16572), .B2(n15619), .A(n12181), .ZN(n12186) );
  AOI21_X1 U14037 ( .B1(n16572), .B2(n12182), .A(n16437), .ZN(n12184) );
  AND2_X1 U14038 ( .A1(n12184), .A2(n12183), .ZN(n16571) );
  NAND2_X1 U14039 ( .A1(n16571), .A2(n16518), .ZN(n12185) );
  OAI211_X1 U14040 ( .C1(n16577), .C2(n15592), .A(n12186), .B(n12185), .ZN(
        n12187) );
  INV_X1 U14041 ( .A(n12187), .ZN(n12188) );
  OAI21_X1 U14042 ( .B1(n16522), .B2(n16575), .A(n12188), .ZN(P1_U3282) );
  OAI222_X1 U14043 ( .A1(n14787), .A2(n12191), .B1(n14783), .B2(n12190), .C1(
        P2_U3088), .C2(n12189), .ZN(P2_U3303) );
  XNOR2_X1 U14044 ( .A(n12192), .B(n12752), .ZN(n16546) );
  OAI211_X1 U14045 ( .C1(n8521), .C2(n12194), .A(n13299), .B(n12193), .ZN(
        n12195) );
  AOI22_X1 U14046 ( .A1(n12991), .A2(n13251), .B1(n12975), .B2(n12992), .ZN(
        n12208) );
  NAND2_X1 U14047 ( .A1(n12195), .A2(n12208), .ZN(n16542) );
  NAND2_X1 U14048 ( .A1(n16542), .A2(n13310), .ZN(n12198) );
  OAI22_X1 U14049 ( .A1(n13304), .A2(n12639), .B1(n12206), .B2(n16360), .ZN(
        n12196) );
  AOI21_X1 U14050 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n16369), .A(n12196), 
        .ZN(n12197) );
  OAI211_X1 U14051 ( .C1(n13313), .C2(n16546), .A(n12198), .B(n12197), .ZN(
        P3_U3223) );
  INV_X1 U14052 ( .A(n12204), .ZN(n12200) );
  NOR2_X1 U14053 ( .A1(n12199), .A2(n12992), .ZN(n12201) );
  XNOR2_X1 U14054 ( .A(n12639), .B(n12821), .ZN(n12264) );
  XNOR2_X1 U14055 ( .A(n12264), .B(n12640), .ZN(n12202) );
  OAI21_X1 U14056 ( .B1(n12200), .B2(n12201), .A(n12202), .ZN(n12205) );
  NOR2_X1 U14057 ( .A1(n12202), .A2(n12201), .ZN(n12203) );
  NAND3_X1 U14058 ( .A1(n12205), .A2(n7876), .A3(n12266), .ZN(n12212) );
  NOR2_X1 U14059 ( .A1(n12955), .A2(n12206), .ZN(n12210) );
  OAI21_X1 U14060 ( .B1(n12208), .B2(n12976), .A(n12207), .ZN(n12209) );
  AOI211_X1 U14061 ( .C1(n16543), .C2(n12966), .A(n12210), .B(n12209), .ZN(
        n12211) );
  NAND2_X1 U14062 ( .A1(n12212), .A2(n12211), .ZN(P3_U3157) );
  NAND2_X1 U14063 ( .A1(n16614), .A2(n16530), .ZN(n12213) );
  OAI211_X1 U14064 ( .C1(n16619), .C2(n12215), .A(n12214), .B(n12213), .ZN(
        n12219) );
  AOI211_X1 U14065 ( .C1(n12217), .C2(n12216), .A(n15029), .B(n7602), .ZN(
        n12218) );
  AOI211_X1 U14066 ( .C1(n16610), .C2(n16531), .A(n12219), .B(n12218), .ZN(
        n12220) );
  INV_X1 U14067 ( .A(n12220), .ZN(P1_U3231) );
  INV_X1 U14068 ( .A(n12221), .ZN(n12533) );
  OAI222_X1 U14069 ( .A1(n14787), .A2(n12223), .B1(n14783), .B2(n12533), .C1(
        n12222), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U14070 ( .A(n12193), .ZN(n12225) );
  OAI21_X1 U14071 ( .B1(n12225), .B2(n12224), .A(n12751), .ZN(n12227) );
  AOI21_X1 U14072 ( .B1(n12227), .B2(n12226), .A(n16349), .ZN(n12230) );
  OAI22_X1 U14073 ( .A1(n12229), .A2(n16350), .B1(n12228), .B2(n16352), .ZN(
        n12268) );
  NOR2_X1 U14074 ( .A1(n12230), .A2(n12268), .ZN(n16564) );
  OAI22_X1 U14075 ( .A1(n13307), .A2(n12231), .B1(n12270), .B2(n16360), .ZN(
        n12232) );
  AOI21_X1 U14076 ( .B1(n12272), .B2(n13260), .A(n12232), .ZN(n12235) );
  XNOR2_X1 U14077 ( .A(n12233), .B(n12751), .ZN(n16567) );
  NAND2_X1 U14078 ( .A1(n16567), .A2(n13266), .ZN(n12234) );
  OAI211_X1 U14079 ( .C1(n16564), .C2(n16369), .A(n12235), .B(n12234), .ZN(
        P3_U3222) );
  AOI211_X1 U14080 ( .C1(n16558), .C2(n12238), .A(n12237), .B(n12236), .ZN(
        n12242) );
  AOI22_X1 U14081 ( .A1(n7765), .A2(n12239), .B1(P2_REG1_REG_13__SCAN_IN), 
        .B2(n16559), .ZN(n12240) );
  OAI21_X1 U14082 ( .B1(n12242), .B2(n16559), .A(n12240), .ZN(P2_U3512) );
  AOI22_X1 U14083 ( .A1(n7765), .A2(n9744), .B1(P2_REG0_REG_13__SCAN_IN), .B2(
        n16561), .ZN(n12241) );
  OAI21_X1 U14084 ( .B1(n12242), .B2(n16561), .A(n12241), .ZN(P2_U3469) );
  INV_X1 U14085 ( .A(n16572), .ZN(n12263) );
  NAND2_X1 U14086 ( .A1(n16572), .A2(n14917), .ZN(n12244) );
  NAND2_X1 U14087 ( .A1(n14916), .A2(n15318), .ZN(n12243) );
  NAND2_X1 U14088 ( .A1(n12244), .A2(n12243), .ZN(n12245) );
  XNOR2_X1 U14089 ( .A(n12245), .B(n14919), .ZN(n12459) );
  NOR2_X1 U14090 ( .A1(n14830), .A2(n12246), .ZN(n12247) );
  AOI21_X1 U14091 ( .B1(n16572), .B2(n14916), .A(n12247), .ZN(n12460) );
  XNOR2_X1 U14092 ( .A(n12459), .B(n12460), .ZN(n12254) );
  INV_X1 U14093 ( .A(n12248), .ZN(n12249) );
  OAI21_X1 U14094 ( .B1(n12254), .B2(n12253), .A(n12463), .ZN(n12255) );
  NAND2_X1 U14095 ( .A1(n12255), .A2(n16612), .ZN(n12262) );
  INV_X1 U14096 ( .A(n12256), .ZN(n12259) );
  NOR2_X1 U14097 ( .A1(n16619), .A2(n12257), .ZN(n12258) );
  AOI211_X1 U14098 ( .C1(n16614), .C2(n12260), .A(n12259), .B(n12258), .ZN(
        n12261) );
  OAI211_X1 U14099 ( .C1(n12263), .C2(n15003), .A(n12262), .B(n12261), .ZN(
        P1_U3236) );
  NAND2_X1 U14100 ( .A1(n12264), .A2(n12640), .ZN(n12265) );
  XNOR2_X1 U14101 ( .A(n12272), .B(n11080), .ZN(n12398) );
  XNOR2_X1 U14102 ( .A(n12398), .B(n12267), .ZN(n12396) );
  XNOR2_X1 U14103 ( .A(n12397), .B(n12396), .ZN(n12274) );
  AOI22_X1 U14104 ( .A1(n12268), .A2(n12870), .B1(P3_REG3_REG_11__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12269) );
  OAI21_X1 U14105 ( .B1(n12270), .B2(n12955), .A(n12269), .ZN(n12271) );
  AOI21_X1 U14106 ( .B1(n12272), .B2(n12966), .A(n12271), .ZN(n12273) );
  OAI21_X1 U14107 ( .B1(n12274), .B2(n12969), .A(n12273), .ZN(P3_U3176) );
  XOR2_X1 U14108 ( .A(n12275), .B(n14303), .Z(n12276) );
  AOI222_X1 U14109 ( .A1(n14606), .A2(n12276), .B1(n14352), .B2(n14589), .C1(
        n14354), .C2(n14588), .ZN(n14727) );
  INV_X1 U14110 ( .A(n12376), .ZN(n12277) );
  AOI211_X1 U14111 ( .C1(n14725), .C2(n12278), .A(n7437), .B(n12277), .ZN(
        n14724) );
  INV_X1 U14112 ( .A(n12279), .ZN(n12280) );
  AOI22_X1 U14113 ( .A1(n14622), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n12280), 
        .B2(n14615), .ZN(n12281) );
  OAI21_X1 U14114 ( .B1(n7968), .B2(n14619), .A(n12281), .ZN(n12286) );
  OR2_X1 U14115 ( .A1(n12282), .A2(n14303), .ZN(n12283) );
  NAND2_X1 U14116 ( .A1(n12284), .A2(n12283), .ZN(n14728) );
  NOR2_X1 U14117 ( .A1(n14728), .A2(n14580), .ZN(n12285) );
  AOI211_X1 U14118 ( .C1(n14724), .C2(n14632), .A(n12286), .B(n12285), .ZN(
        n12287) );
  OAI21_X1 U14119 ( .B1(n14727), .B2(n14622), .A(n12287), .ZN(P2_U3251) );
  OAI21_X1 U14120 ( .B1(n12289), .B2(n15247), .A(n12288), .ZN(n12290) );
  INV_X1 U14121 ( .A(n12290), .ZN(n12446) );
  INV_X1 U14122 ( .A(n12291), .ZN(n12293) );
  INV_X1 U14123 ( .A(n12494), .ZN(n12292) );
  AOI211_X1 U14124 ( .C1(n15105), .C2(n12293), .A(n16437), .B(n12292), .ZN(
        n12443) );
  OAI22_X1 U14125 ( .A1(n12294), .A2(n16512), .B1(n10909), .B2(n15515), .ZN(
        n12295) );
  AOI21_X1 U14126 ( .B1(n12443), .B2(n16518), .A(n12295), .ZN(n12303) );
  OAI21_X1 U14127 ( .B1(n12298), .B2(n12297), .A(n12296), .ZN(n12299) );
  NAND2_X1 U14128 ( .A1(n12299), .A2(n16536), .ZN(n12444) );
  OAI22_X1 U14129 ( .A1(n12467), .A2(n15293), .B1(n14805), .B2(n15016), .ZN(
        n12479) );
  INV_X1 U14130 ( .A(n12479), .ZN(n12300) );
  OAI211_X1 U14131 ( .C1(n16490), .C2(n12482), .A(n12444), .B(n12300), .ZN(
        n12301) );
  NAND2_X1 U14132 ( .A1(n12301), .A2(n15515), .ZN(n12302) );
  OAI211_X1 U14133 ( .C1(n12446), .C2(n15592), .A(n12303), .B(n12302), .ZN(
        P1_U3280) );
  INV_X1 U14134 ( .A(n12304), .ZN(n12307) );
  XNOR2_X1 U14135 ( .A(n14716), .B(n10884), .ZN(n12310) );
  AND2_X1 U14136 ( .A1(n14352), .A2(n7437), .ZN(n12308) );
  NAND2_X1 U14137 ( .A1(n12310), .A2(n12308), .ZN(n12312) );
  OAI21_X1 U14138 ( .B1(n12310), .B2(n12308), .A(n12312), .ZN(n12391) );
  NOR2_X1 U14139 ( .A1(n13976), .A2(n12309), .ZN(n12311) );
  AOI22_X1 U14140 ( .A1(n12390), .A2(n13990), .B1(n12311), .B2(n12310), .ZN(
        n12324) );
  XNOR2_X1 U14141 ( .A(n14122), .B(n7433), .ZN(n12415) );
  NAND2_X1 U14142 ( .A1(n14351), .A2(n7437), .ZN(n12416) );
  XNOR2_X1 U14143 ( .A(n12415), .B(n12416), .ZN(n12313) );
  INV_X1 U14144 ( .A(n12313), .ZN(n12323) );
  INV_X1 U14145 ( .A(n12312), .ZN(n12314) );
  NAND2_X1 U14146 ( .A1(n14350), .A2(n14589), .ZN(n12316) );
  NAND2_X1 U14147 ( .A1(n14352), .A2(n14588), .ZN(n12315) );
  NAND2_X1 U14148 ( .A1(n12316), .A2(n12315), .ZN(n12431) );
  INV_X1 U14149 ( .A(n12317), .ZN(n12436) );
  OAI22_X1 U14150 ( .A1(n13970), .A2(n12436), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12318), .ZN(n12319) );
  AOI21_X1 U14151 ( .B1(n13972), .B2(n12431), .A(n12319), .ZN(n12320) );
  OAI21_X1 U14152 ( .B1(n14769), .B2(n13975), .A(n12320), .ZN(n12321) );
  AOI21_X1 U14153 ( .B1(n12427), .B2(n13990), .A(n12321), .ZN(n12322) );
  OAI21_X1 U14154 ( .B1(n12324), .B2(n12323), .A(n12322), .ZN(P2_U3198) );
  INV_X1 U14155 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n12332) );
  NAND2_X1 U14156 ( .A1(n12325), .A2(n16443), .ZN(n12330) );
  AOI21_X1 U14157 ( .B1(n15101), .B2(n16573), .A(n14940), .ZN(n12329) );
  NAND3_X1 U14158 ( .A1(n12165), .A2(n16536), .A3(n12326), .ZN(n12328) );
  NAND4_X1 U14159 ( .A1(n12330), .A2(n12329), .A3(n12328), .A4(n12327), .ZN(
        n12333) );
  NAND2_X1 U14160 ( .A1(n12333), .A2(n16540), .ZN(n12331) );
  OAI21_X1 U14161 ( .B1(n16540), .B2(n12332), .A(n12331), .ZN(P1_U3495) );
  NAND2_X1 U14162 ( .A1(n12333), .A2(n7435), .ZN(n12334) );
  OAI21_X1 U14163 ( .B1(n7435), .B2(n9419), .A(n12334), .ZN(P1_U3540) );
  NAND2_X1 U14164 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n12354), .ZN(n12341) );
  INV_X1 U14165 ( .A(n12341), .ZN(n12335) );
  AOI21_X1 U14166 ( .B1(n12518), .B2(n15868), .A(n12335), .ZN(n15878) );
  NAND2_X1 U14167 ( .A1(n12349), .A2(n12336), .ZN(n12338) );
  NAND2_X1 U14168 ( .A1(n12338), .A2(n12337), .ZN(n15863) );
  NOR2_X1 U14169 ( .A1(n12340), .A2(n12437), .ZN(n12339) );
  AOI21_X1 U14170 ( .B1(n12437), .B2(n12340), .A(n12339), .ZN(n15862) );
  NAND2_X1 U14171 ( .A1(n15863), .A2(n15862), .ZN(n15861) );
  OAI21_X1 U14172 ( .B1(n12437), .B2(n12340), .A(n15861), .ZN(n15879) );
  NAND2_X1 U14173 ( .A1(n15878), .A2(n15879), .ZN(n15876) );
  NAND2_X1 U14174 ( .A1(n12341), .A2(n15876), .ZN(n12342) );
  NOR2_X1 U14175 ( .A1(n12342), .A2(n14413), .ZN(n14418) );
  AOI21_X1 U14176 ( .B1(n12342), .B2(n14413), .A(n14418), .ZN(n12343) );
  INV_X1 U14177 ( .A(n12343), .ZN(n12344) );
  NOR2_X1 U14178 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n12344), .ZN(n14417) );
  AOI21_X1 U14179 ( .B1(n12344), .B2(P2_REG2_REG_18__SCAN_IN), .A(n14417), 
        .ZN(n12359) );
  NOR2_X1 U14180 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13969), .ZN(n12347) );
  NOR2_X1 U14181 ( .A1(n15842), .A2(n12345), .ZN(n12346) );
  AOI211_X1 U14182 ( .C1(n15875), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n12347), 
        .B(n12346), .ZN(n12358) );
  NAND2_X1 U14183 ( .A1(n12349), .A2(n12348), .ZN(n12351) );
  NAND2_X1 U14184 ( .A1(n12351), .A2(n12350), .ZN(n15856) );
  XNOR2_X1 U14185 ( .A(n15859), .B(n14713), .ZN(n15857) );
  NAND2_X1 U14186 ( .A1(n15856), .A2(n15857), .ZN(n12353) );
  NAND2_X1 U14187 ( .A1(n15859), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n12352) );
  NAND2_X1 U14188 ( .A1(n12353), .A2(n12352), .ZN(n15871) );
  INV_X1 U14189 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14706) );
  XNOR2_X1 U14190 ( .A(n12354), .B(n14706), .ZN(n15872) );
  AND2_X1 U14191 ( .A1(n12354), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n12355) );
  AOI21_X1 U14192 ( .B1(n15871), .B2(n15872), .A(n12355), .ZN(n14411) );
  XNOR2_X1 U14193 ( .A(n14411), .B(n14413), .ZN(n14414) );
  XOR2_X1 U14194 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14414), .Z(n12356) );
  NAND2_X1 U14195 ( .A1(n12356), .A2(n15873), .ZN(n12357) );
  OAI211_X1 U14196 ( .C1(n12359), .C2(n15848), .A(n12358), .B(n12357), .ZN(
        P2_U3232) );
  OAI21_X1 U14197 ( .B1(n12361), .B2(n12750), .A(n12360), .ZN(n16588) );
  INV_X1 U14198 ( .A(n16588), .ZN(n16585) );
  XNOR2_X1 U14199 ( .A(n12362), .B(n12750), .ZN(n12363) );
  AOI22_X1 U14200 ( .A1(n12991), .A2(n12975), .B1(n13251), .B2(n12990), .ZN(
        n12407) );
  OAI21_X1 U14201 ( .B1(n12363), .B2(n16349), .A(n12407), .ZN(n16587) );
  NAND2_X1 U14202 ( .A1(n16587), .A2(n13310), .ZN(n12366) );
  OAI22_X1 U14203 ( .A1(n13307), .A2(n13029), .B1(n12410), .B2(n16360), .ZN(
        n12364) );
  AOI21_X1 U14204 ( .B1(n12412), .B2(n13260), .A(n12364), .ZN(n12365) );
  OAI211_X1 U14205 ( .C1(n13313), .C2(n16585), .A(n12366), .B(n12365), .ZN(
        P3_U3221) );
  OAI21_X1 U14206 ( .B1(n12368), .B2(n14305), .A(n12367), .ZN(n12369) );
  NAND2_X1 U14207 ( .A1(n12369), .A2(n14606), .ZN(n12372) );
  NAND2_X1 U14208 ( .A1(n14353), .A2(n14588), .ZN(n12371) );
  NAND2_X1 U14209 ( .A1(n14351), .A2(n14589), .ZN(n12370) );
  AND2_X1 U14210 ( .A1(n12371), .A2(n12370), .ZN(n12389) );
  NAND2_X1 U14211 ( .A1(n12372), .A2(n12389), .ZN(n14723) );
  INV_X1 U14212 ( .A(n14723), .ZN(n12384) );
  NAND2_X1 U14213 ( .A1(n12373), .A2(n14305), .ZN(n12374) );
  NAND2_X1 U14214 ( .A1(n12375), .A2(n12374), .ZN(n14718) );
  NAND2_X1 U14215 ( .A1(n7757), .A2(n12376), .ZN(n12377) );
  NAND2_X1 U14216 ( .A1(n12377), .A2(n14430), .ZN(n12378) );
  OR2_X1 U14217 ( .A1(n12435), .A2(n12378), .ZN(n14719) );
  OAI22_X1 U14218 ( .A1(n11368), .A2(n12379), .B1(n12385), .B2(n14624), .ZN(
        n12380) );
  AOI21_X1 U14219 ( .B1(n7757), .B2(n14628), .A(n12380), .ZN(n12381) );
  OAI21_X1 U14220 ( .B1(n14719), .B2(n14556), .A(n12381), .ZN(n12382) );
  AOI21_X1 U14221 ( .B1(n14630), .B2(n14718), .A(n12382), .ZN(n12383) );
  OAI21_X1 U14222 ( .B1(n12384), .B2(n14622), .A(n12383), .ZN(P2_U3250) );
  INV_X1 U14223 ( .A(n12385), .ZN(n12386) );
  NAND2_X1 U14224 ( .A1(n13985), .A2(n12386), .ZN(n12387) );
  OAI211_X1 U14225 ( .C1(n13988), .C2(n12389), .A(n12388), .B(n12387), .ZN(
        n12394) );
  AOI211_X1 U14226 ( .C1(n12392), .C2(n12391), .A(n13963), .B(n12390), .ZN(
        n12393) );
  AOI211_X1 U14227 ( .C1(n7757), .C2(n13983), .A(n12394), .B(n12393), .ZN(
        n12395) );
  INV_X1 U14228 ( .A(n12395), .ZN(P2_U3213) );
  NAND2_X1 U14229 ( .A1(n12991), .A2(n12398), .ZN(n12399) );
  NAND2_X1 U14230 ( .A1(n12400), .A2(n12399), .ZN(n12795) );
  INV_X1 U14231 ( .A(n12653), .ZN(n12403) );
  INV_X1 U14232 ( .A(n12401), .ZN(n12402) );
  MUX2_X1 U14233 ( .A(n12403), .B(n12402), .S(n11080), .Z(n12794) );
  MUX2_X1 U14234 ( .A(n12404), .B(n12652), .S(n12821), .Z(n12793) );
  INV_X1 U14235 ( .A(n12793), .ZN(n12405) );
  NOR2_X1 U14236 ( .A1(n12794), .A2(n12405), .ZN(n12406) );
  XNOR2_X1 U14237 ( .A(n12795), .B(n12406), .ZN(n12414) );
  INV_X1 U14238 ( .A(n12407), .ZN(n12408) );
  AOI22_X1 U14239 ( .A1(n12408), .A2(n12870), .B1(P3_REG3_REG_12__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12409) );
  OAI21_X1 U14240 ( .B1(n12410), .B2(n12955), .A(n12409), .ZN(n12411) );
  AOI21_X1 U14241 ( .B1(n12412), .B2(n12966), .A(n12411), .ZN(n12413) );
  OAI21_X1 U14242 ( .B1(n12414), .B2(n12969), .A(n12413), .ZN(P3_U3164) );
  INV_X1 U14243 ( .A(n12415), .ZN(n12424) );
  INV_X1 U14244 ( .A(n12416), .ZN(n12417) );
  NOR2_X1 U14245 ( .A1(n12424), .A2(n12417), .ZN(n12418) );
  XNOR2_X1 U14246 ( .A(n14763), .B(n10884), .ZN(n12537) );
  NAND2_X1 U14247 ( .A1(n14350), .A2(n7437), .ZN(n12535) );
  XNOR2_X1 U14248 ( .A(n12537), .B(n12535), .ZN(n12425) );
  NAND2_X1 U14249 ( .A1(n14587), .A2(n14589), .ZN(n12420) );
  NAND2_X1 U14250 ( .A1(n14351), .A2(n14588), .ZN(n12419) );
  NAND2_X1 U14251 ( .A1(n12420), .A2(n12419), .ZN(n12515) );
  OAI22_X1 U14252 ( .A1(n13970), .A2(n12517), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12421), .ZN(n12423) );
  INV_X1 U14253 ( .A(n14763), .ZN(n14708) );
  NOR2_X1 U14254 ( .A1(n14708), .A2(n13975), .ZN(n12422) );
  AOI211_X1 U14255 ( .C1(n13972), .C2(n12515), .A(n12423), .B(n12422), .ZN(
        n12429) );
  AOI22_X1 U14256 ( .A1(n12424), .A2(n13990), .B1(n13894), .B2(n14351), .ZN(
        n12426) );
  OR3_X1 U14257 ( .A1(n12427), .A2(n12426), .A3(n12425), .ZN(n12428) );
  OAI211_X1 U14258 ( .C1(n12539), .C2(n13963), .A(n12429), .B(n12428), .ZN(
        P2_U3200) );
  XNOR2_X1 U14259 ( .A(n12430), .B(n14304), .ZN(n12432) );
  AOI21_X1 U14260 ( .B1(n12432), .B2(n14606), .A(n12431), .ZN(n14710) );
  OAI21_X1 U14261 ( .B1(n12434), .B2(n8856), .A(n12433), .ZN(n14711) );
  INV_X1 U14262 ( .A(n14711), .ZN(n12441) );
  OAI211_X1 U14263 ( .C1(n12435), .C2(n14769), .A(n14430), .B(n12519), .ZN(
        n14709) );
  OAI22_X1 U14264 ( .A1(n11368), .A2(n12437), .B1(n12436), .B2(n14624), .ZN(
        n12438) );
  AOI21_X1 U14265 ( .B1(n14122), .B2(n14628), .A(n12438), .ZN(n12439) );
  OAI21_X1 U14266 ( .B1(n14709), .B2(n14556), .A(n12439), .ZN(n12440) );
  AOI21_X1 U14267 ( .B1(n12441), .B2(n14630), .A(n12440), .ZN(n12442) );
  OAI21_X1 U14268 ( .B1(n14710), .B2(n14622), .A(n12442), .ZN(P2_U3249) );
  AOI211_X1 U14269 ( .C1(n16573), .C2(n15105), .A(n12479), .B(n12443), .ZN(
        n12445) );
  OAI211_X1 U14270 ( .C1(n16576), .C2(n12446), .A(n12445), .B(n12444), .ZN(
        n12448) );
  NAND2_X1 U14271 ( .A1(n12448), .A2(n16540), .ZN(n12447) );
  OAI21_X1 U14272 ( .B1(n16540), .B2(n9435), .A(n12447), .ZN(P1_U3498) );
  NAND2_X1 U14273 ( .A1(n12448), .A2(n7435), .ZN(n12449) );
  OAI21_X1 U14274 ( .B1(n7435), .B2(n9431), .A(n12449), .ZN(P1_U3541) );
  XNOR2_X1 U14275 ( .A(n12450), .B(n12796), .ZN(n16598) );
  INV_X1 U14276 ( .A(n16598), .ZN(n12458) );
  XNOR2_X1 U14277 ( .A(n12451), .B(n12796), .ZN(n12453) );
  AOI22_X1 U14278 ( .A1(n12452), .A2(n12975), .B1(n13251), .B2(n12989), .ZN(
        n12934) );
  OAI21_X1 U14279 ( .B1(n12453), .B2(n16349), .A(n12934), .ZN(n16595) );
  NOR2_X1 U14280 ( .A1(n16594), .A2(n13304), .ZN(n12456) );
  OAI22_X1 U14281 ( .A1(n13307), .A2(n12454), .B1(n12931), .B2(n16360), .ZN(
        n12455) );
  AOI211_X1 U14282 ( .C1(n16595), .C2(n13307), .A(n12456), .B(n12455), .ZN(
        n12457) );
  OAI21_X1 U14283 ( .B1(n13313), .B2(n12458), .A(n12457), .ZN(P3_U3220) );
  INV_X1 U14284 ( .A(n12459), .ZN(n12461) );
  NAND2_X1 U14285 ( .A1(n12461), .A2(n12460), .ZN(n12462) );
  NAND2_X1 U14286 ( .A1(n15101), .A2(n14917), .ZN(n12465) );
  NAND2_X1 U14287 ( .A1(n14916), .A2(n15317), .ZN(n12464) );
  NAND2_X1 U14288 ( .A1(n12465), .A2(n12464), .ZN(n12466) );
  XNOR2_X1 U14289 ( .A(n12466), .B(n14827), .ZN(n12470) );
  NOR2_X1 U14290 ( .A1(n14830), .A2(n12467), .ZN(n12468) );
  AOI21_X1 U14291 ( .B1(n15101), .B2(n14916), .A(n12468), .ZN(n12471) );
  XNOR2_X1 U14292 ( .A(n12470), .B(n12471), .ZN(n14946) );
  INV_X1 U14293 ( .A(n12470), .ZN(n12473) );
  INV_X1 U14294 ( .A(n12471), .ZN(n12472) );
  NAND2_X1 U14295 ( .A1(n12473), .A2(n12472), .ZN(n12474) );
  NAND2_X1 U14296 ( .A1(n14943), .A2(n12474), .ZN(n14797) );
  NAND2_X1 U14297 ( .A1(n15105), .A2(n14917), .ZN(n12476) );
  NAND2_X1 U14298 ( .A1(n14916), .A2(n15316), .ZN(n12475) );
  NAND2_X1 U14299 ( .A1(n12476), .A2(n12475), .ZN(n12477) );
  XNOR2_X1 U14300 ( .A(n12477), .B(n14919), .ZN(n14800) );
  NOR2_X1 U14301 ( .A1(n14830), .A2(n12488), .ZN(n12478) );
  AOI21_X1 U14302 ( .B1(n15105), .B2(n14916), .A(n12478), .ZN(n14798) );
  XNOR2_X1 U14303 ( .A(n14800), .B(n14798), .ZN(n14796) );
  XNOR2_X1 U14304 ( .A(n14797), .B(n14796), .ZN(n12485) );
  NAND2_X1 U14305 ( .A1(n16614), .A2(n12479), .ZN(n12480) );
  OAI211_X1 U14306 ( .C1(n16619), .C2(n12482), .A(n12481), .B(n12480), .ZN(
        n12483) );
  AOI21_X1 U14307 ( .B1(n15105), .B2(n16610), .A(n12483), .ZN(n12484) );
  OAI21_X1 U14308 ( .B1(n12485), .B2(n15029), .A(n12484), .ZN(P1_U3234) );
  XNOR2_X1 U14309 ( .A(n12486), .B(n15248), .ZN(n12489) );
  OAI22_X1 U14310 ( .A1(n12488), .A2(n15293), .B1(n12487), .B2(n15016), .ZN(
        n16615) );
  AOI21_X1 U14311 ( .B1(n12489), .B2(n16536), .A(n16615), .ZN(n15740) );
  OAI21_X1 U14312 ( .B1(n7446), .B2(n12491), .A(n12490), .ZN(n15741) );
  NAND2_X1 U14313 ( .A1(n16522), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n12492) );
  OAI21_X1 U14314 ( .B1(n16490), .B2(n16618), .A(n12492), .ZN(n12493) );
  AOI21_X1 U14315 ( .B1(n16611), .B2(n15619), .A(n12493), .ZN(n12497) );
  AOI21_X1 U14316 ( .B1(n16611), .B2(n12494), .A(n16437), .ZN(n12495) );
  AND2_X1 U14317 ( .A1(n12495), .A2(n12501), .ZN(n15738) );
  NAND2_X1 U14318 ( .A1(n15738), .A2(n16518), .ZN(n12496) );
  OAI211_X1 U14319 ( .C1(n15741), .C2(n15592), .A(n12497), .B(n12496), .ZN(
        n12498) );
  INV_X1 U14320 ( .A(n12498), .ZN(n12499) );
  OAI21_X1 U14321 ( .B1(n16522), .B2(n15740), .A(n12499), .ZN(P1_U3279) );
  XNOR2_X1 U14322 ( .A(n12500), .B(n12510), .ZN(n15737) );
  OAI21_X1 U14323 ( .B1(n8100), .B2(n8101), .A(n15631), .ZN(n15729) );
  INV_X1 U14324 ( .A(n15729), .ZN(n12508) );
  AND2_X1 U14325 ( .A1(n16518), .A2(n16473), .ZN(n15590) );
  NAND2_X1 U14326 ( .A1(n15008), .A2(n15313), .ZN(n12503) );
  NAND2_X1 U14327 ( .A1(n15006), .A2(n15315), .ZN(n12502) );
  NAND2_X1 U14328 ( .A1(n12503), .A2(n12502), .ZN(n15731) );
  INV_X1 U14329 ( .A(n15731), .ZN(n12504) );
  OAI22_X1 U14330 ( .A1(n16522), .A2(n12504), .B1(n15026), .B2(n16490), .ZN(
        n12505) );
  AOI21_X1 U14331 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n16522), .A(n12505), 
        .ZN(n12506) );
  OAI21_X1 U14332 ( .B1(n8100), .B2(n16512), .A(n12506), .ZN(n12507) );
  AOI21_X1 U14333 ( .B1(n12508), .B2(n15590), .A(n12507), .ZN(n12512) );
  NAND2_X1 U14334 ( .A1(n12509), .A2(n12510), .ZN(n15733) );
  NAND3_X1 U14335 ( .A1(n15734), .A2(n15733), .A3(n15537), .ZN(n12511) );
  OAI211_X1 U14336 ( .C1(n15737), .C2(n15592), .A(n12512), .B(n12511), .ZN(
        P1_U3278) );
  XNOR2_X1 U14337 ( .A(n12514), .B(n12513), .ZN(n12516) );
  AOI21_X1 U14338 ( .B1(n12516), .B2(n14606), .A(n12515), .ZN(n14703) );
  OAI22_X1 U14339 ( .A1(n11368), .A2(n12518), .B1(n12517), .B2(n14624), .ZN(
        n12523) );
  AOI21_X1 U14340 ( .B1(n12519), .B2(n14763), .A(n7437), .ZN(n12521) );
  INV_X1 U14341 ( .A(n12520), .ZN(n14613) );
  NAND2_X1 U14342 ( .A1(n12521), .A2(n14613), .ZN(n14702) );
  NOR2_X1 U14343 ( .A1(n14702), .A2(n14556), .ZN(n12522) );
  AOI211_X1 U14344 ( .C1(n14628), .C2(n14763), .A(n12523), .B(n12522), .ZN(
        n12526) );
  XNOR2_X1 U14345 ( .A(n12524), .B(n14307), .ZN(n14704) );
  OR2_X1 U14346 ( .A1(n14704), .A2(n14580), .ZN(n12525) );
  OAI211_X1 U14347 ( .C1(n14703), .C2(n14622), .A(n12526), .B(n12525), .ZN(
        P2_U3248) );
  INV_X1 U14348 ( .A(n12527), .ZN(n12528) );
  AND2_X1 U14349 ( .A1(n12530), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U14350 ( .A1(n12530), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U14351 ( .A1(n12530), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U14352 ( .A1(n12530), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U14353 ( .A1(n12530), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U14354 ( .A1(n12530), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U14355 ( .A1(n12530), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U14356 ( .A1(n12530), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U14357 ( .A1(n12530), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U14358 ( .A1(n12530), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U14359 ( .A1(n12530), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U14360 ( .A1(n12530), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U14361 ( .A1(n12530), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U14362 ( .A1(n12530), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U14363 ( .A1(n12530), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U14364 ( .A1(n12530), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U14365 ( .A1(n12530), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U14366 ( .A1(n12530), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U14367 ( .A1(n12530), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U14368 ( .A1(n12530), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U14369 ( .A1(n12530), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U14370 ( .A1(n12530), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U14371 ( .A1(n12530), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U14372 ( .A1(n12530), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U14373 ( .A1(n16301), .A2(n12529), .ZN(P1_U3085) );
  AND2_X1 U14374 ( .A1(n12530), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U14375 ( .A1(n12530), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U14376 ( .A1(n12530), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U14377 ( .A1(n12530), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U14378 ( .A1(n12530), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U14379 ( .A1(n12530), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  INV_X1 U14380 ( .A(n12531), .ZN(n12532) );
  OAI222_X1 U14381 ( .A1(P3_U3151), .A2(n7430), .B1(n13850), .B2(n13410), .C1(
        n13853), .C2(n12532), .ZN(P3_U3267) );
  OAI222_X1 U14382 ( .A1(n15777), .A2(n12534), .B1(n15780), .B2(n12533), .C1(
        P1_U3086), .C2(n9705), .ZN(P1_U3330) );
  XNOR2_X1 U14383 ( .A(n14596), .B(n10884), .ZN(n12542) );
  NAND2_X1 U14384 ( .A1(n14349), .A2(n7437), .ZN(n12543) );
  INV_X1 U14385 ( .A(n12535), .ZN(n12536) );
  XNOR2_X1 U14386 ( .A(n14698), .B(n10884), .ZN(n13895) );
  AND2_X1 U14387 ( .A1(n14587), .A2(n7437), .ZN(n12540) );
  NAND2_X1 U14388 ( .A1(n13895), .A2(n12540), .ZN(n12541) );
  OAI21_X1 U14389 ( .B1(n13895), .B2(n12540), .A(n12541), .ZN(n13964) );
  XNOR2_X1 U14390 ( .A(n12542), .B(n12543), .ZN(n13893) );
  XNOR2_X1 U14391 ( .A(n14688), .B(n10884), .ZN(n13953) );
  AND2_X1 U14392 ( .A1(n14590), .A2(n7437), .ZN(n12545) );
  NAND2_X1 U14393 ( .A1(n13953), .A2(n12545), .ZN(n13949) );
  XNOR2_X1 U14394 ( .A(n14551), .B(n10884), .ZN(n12546) );
  NOR2_X1 U14395 ( .A1(n14165), .A2(n14430), .ZN(n12547) );
  XNOR2_X1 U14396 ( .A(n12546), .B(n12547), .ZN(n13925) );
  INV_X1 U14397 ( .A(n12546), .ZN(n12548) );
  NAND2_X1 U14398 ( .A1(n12548), .A2(n12547), .ZN(n12549) );
  XNOR2_X1 U14399 ( .A(n14675), .B(n10884), .ZN(n13857) );
  AOI22_X1 U14400 ( .A1(n7603), .A2(n13990), .B1(n13894), .B2(n14347), .ZN(
        n12554) );
  OAI22_X1 U14401 ( .A1(n14177), .A2(n13968), .B1(n14165), .B2(n13967), .ZN(
        n14533) );
  OAI22_X1 U14402 ( .A1(n13970), .A2(n14540), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12550), .ZN(n12552) );
  INV_X1 U14403 ( .A(n14675), .ZN(n14173) );
  NOR2_X1 U14404 ( .A1(n14173), .A2(n13975), .ZN(n12551) );
  AOI211_X1 U14405 ( .C1(n13972), .C2(n14533), .A(n12552), .B(n12551), .ZN(
        n12553) );
  OAI21_X1 U14406 ( .B1(n13860), .B2(n12554), .A(n12553), .ZN(P2_U3207) );
  NAND2_X1 U14407 ( .A1(n15771), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12557) );
  XNOR2_X1 U14408 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n12565) );
  NAND2_X1 U14409 ( .A1(n12567), .A2(n12565), .ZN(n12559) );
  INV_X1 U14410 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15766) );
  NAND2_X1 U14411 ( .A1(n15766), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12558) );
  NAND2_X1 U14412 ( .A1(n12559), .A2(n12558), .ZN(n12561) );
  INV_X1 U14413 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n14231) );
  XNOR2_X1 U14414 ( .A(n14231), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n12560) );
  XNOR2_X1 U14415 ( .A(n12561), .B(n12560), .ZN(n13840) );
  NAND2_X1 U14416 ( .A1(n13840), .A2(n12568), .ZN(n12564) );
  NAND2_X1 U14417 ( .A1(n12562), .A2(SI_31_), .ZN(n12563) );
  NOR2_X1 U14418 ( .A1(n13380), .A2(n13091), .ZN(n12765) );
  INV_X1 U14419 ( .A(n12565), .ZN(n12566) );
  XNOR2_X1 U14420 ( .A(n12567), .B(n12566), .ZN(n12846) );
  NAND2_X1 U14421 ( .A1(n12846), .A2(n12568), .ZN(n12571) );
  INV_X1 U14422 ( .A(SI_30_), .ZN(n14226) );
  OR2_X1 U14423 ( .A1(n12569), .A2(n14226), .ZN(n12570) );
  NAND2_X1 U14424 ( .A1(n13384), .A2(n12574), .ZN(n12763) );
  NAND2_X1 U14425 ( .A1(n13384), .A2(n13091), .ZN(n12572) );
  INV_X1 U14426 ( .A(n13380), .ZN(n12575) );
  NOR2_X1 U14427 ( .A1(n12576), .A2(n12575), .ZN(n12577) );
  NOR2_X1 U14428 ( .A1(n12577), .A2(n12764), .ZN(n12578) );
  INV_X1 U14429 ( .A(n12580), .ZN(n12769) );
  NAND2_X1 U14430 ( .A1(n12581), .A2(n12731), .ZN(n12583) );
  INV_X1 U14431 ( .A(n13142), .ZN(n13145) );
  INV_X1 U14432 ( .A(n12586), .ZN(n12822) );
  NAND2_X1 U14433 ( .A1(n12587), .A2(n12822), .ZN(n12589) );
  NAND2_X1 U14434 ( .A1(n12589), .A2(n12588), .ZN(n12699) );
  NAND2_X1 U14435 ( .A1(n12591), .A2(n12595), .ZN(n12590) );
  NAND2_X1 U14436 ( .A1(n12590), .A2(n12597), .ZN(n12593) );
  INV_X1 U14437 ( .A(n12591), .ZN(n12592) );
  MUX2_X1 U14438 ( .A(n12593), .B(n12592), .S(n12731), .Z(n12606) );
  NAND2_X1 U14439 ( .A1(n12595), .A2(n12594), .ZN(n12596) );
  NAND4_X1 U14440 ( .A1(n12597), .A2(n16308), .A3(n12596), .A4(n12731), .ZN(
        n12598) );
  NAND2_X1 U14441 ( .A1(n10281), .A2(n12598), .ZN(n12605) );
  NAND2_X1 U14442 ( .A1(n12607), .A2(n12599), .ZN(n12602) );
  NAND2_X1 U14443 ( .A1(n12608), .A2(n12600), .ZN(n12601) );
  MUX2_X1 U14444 ( .A(n12602), .B(n12601), .S(n12731), .Z(n12603) );
  INV_X1 U14445 ( .A(n12603), .ZN(n12604) );
  OAI21_X1 U14446 ( .B1(n12606), .B2(n12605), .A(n12604), .ZN(n12611) );
  MUX2_X1 U14447 ( .A(n12608), .B(n12607), .S(n12731), .Z(n12609) );
  NAND3_X1 U14448 ( .A1(n12611), .A2(n12610), .A3(n12609), .ZN(n12615) );
  MUX2_X1 U14449 ( .A(n12613), .B(n12612), .S(n12731), .Z(n12614) );
  NAND3_X1 U14450 ( .A1(n12615), .A2(n12746), .A3(n12614), .ZN(n12619) );
  MUX2_X1 U14451 ( .A(n12617), .B(n12616), .S(n12728), .Z(n12618) );
  NAND3_X1 U14452 ( .A1(n12619), .A2(n12618), .A3(n12745), .ZN(n12625) );
  MUX2_X1 U14453 ( .A(n12995), .B(n12731), .S(n12620), .Z(n12621) );
  OAI21_X1 U14454 ( .B1(n12728), .B2(n12622), .A(n12621), .ZN(n12623) );
  NAND3_X1 U14455 ( .A1(n12625), .A2(n12624), .A3(n12623), .ZN(n12630) );
  MUX2_X1 U14456 ( .A(n12627), .B(n12626), .S(n12728), .Z(n12628) );
  NAND3_X1 U14457 ( .A1(n12630), .A2(n12629), .A3(n12628), .ZN(n12634) );
  MUX2_X1 U14458 ( .A(n12632), .B(n12631), .S(n12731), .Z(n12633) );
  NAND3_X1 U14459 ( .A1(n12634), .A2(n12741), .A3(n12633), .ZN(n12638) );
  MUX2_X1 U14460 ( .A(n12636), .B(n12635), .S(n12731), .Z(n12637) );
  NAND3_X1 U14461 ( .A1(n12638), .A2(n12752), .A3(n12637), .ZN(n12644) );
  NAND2_X1 U14462 ( .A1(n12640), .A2(n12639), .ZN(n12642) );
  MUX2_X1 U14463 ( .A(n12642), .B(n12641), .S(n12731), .Z(n12643) );
  NAND2_X1 U14464 ( .A1(n12644), .A2(n12643), .ZN(n12645) );
  NAND2_X1 U14465 ( .A1(n12645), .A2(n12751), .ZN(n12650) );
  NAND2_X1 U14466 ( .A1(n12653), .A2(n12646), .ZN(n12647) );
  NAND2_X1 U14467 ( .A1(n12647), .A2(n12728), .ZN(n12649) );
  INV_X1 U14468 ( .A(n12652), .ZN(n12648) );
  AOI21_X1 U14469 ( .B1(n12650), .B2(n12649), .A(n12648), .ZN(n12655) );
  INV_X1 U14470 ( .A(n12655), .ZN(n12657) );
  AOI21_X1 U14471 ( .B1(n12652), .B2(n12651), .A(n12728), .ZN(n12654) );
  OAI21_X1 U14472 ( .B1(n12655), .B2(n12654), .A(n12653), .ZN(n12656) );
  OAI21_X1 U14473 ( .B1(n12657), .B2(n12731), .A(n12656), .ZN(n12661) );
  MUX2_X1 U14474 ( .A(n12658), .B(n12799), .S(n12728), .Z(n12659) );
  NAND2_X1 U14475 ( .A1(n13297), .A2(n12659), .ZN(n12660) );
  AOI21_X1 U14476 ( .B1(n12661), .B2(n12796), .A(n12660), .ZN(n12667) );
  INV_X1 U14477 ( .A(n12662), .ZN(n12664) );
  MUX2_X1 U14478 ( .A(n12664), .B(n12663), .S(n12728), .Z(n12666) );
  OAI21_X1 U14479 ( .B1(n12667), .B2(n12666), .A(n10287), .ZN(n12672) );
  INV_X1 U14480 ( .A(n12668), .ZN(n12674) );
  NAND2_X1 U14481 ( .A1(n12673), .A2(n12674), .ZN(n13272) );
  INV_X1 U14482 ( .A(n13272), .ZN(n13270) );
  MUX2_X1 U14483 ( .A(n12670), .B(n12669), .S(n12731), .Z(n12671) );
  NAND3_X1 U14484 ( .A1(n12672), .A2(n13270), .A3(n12671), .ZN(n12676) );
  MUX2_X1 U14485 ( .A(n12674), .B(n12673), .S(n12728), .Z(n12675) );
  NAND2_X1 U14486 ( .A1(n12676), .A2(n12675), .ZN(n12691) );
  NAND2_X1 U14487 ( .A1(n12677), .A2(n13252), .ZN(n12678) );
  NAND2_X1 U14488 ( .A1(n12679), .A2(n12678), .ZN(n12685) );
  AND2_X1 U14489 ( .A1(n12685), .A2(n13250), .ZN(n12690) );
  INV_X1 U14490 ( .A(n12680), .ZN(n12681) );
  NAND2_X1 U14491 ( .A1(n10289), .A2(n12681), .ZN(n12682) );
  NAND3_X1 U14492 ( .A1(n12735), .A2(n12682), .A3(n13238), .ZN(n12688) );
  INV_X1 U14493 ( .A(n12683), .ZN(n12684) );
  NAND2_X1 U14494 ( .A1(n12685), .A2(n12684), .ZN(n12686) );
  NAND3_X1 U14495 ( .A1(n12736), .A2(n12686), .A3(n10289), .ZN(n12687) );
  MUX2_X1 U14496 ( .A(n12688), .B(n12687), .S(n12728), .Z(n12689) );
  AOI21_X1 U14497 ( .B1(n12691), .B2(n12690), .A(n12689), .ZN(n12694) );
  MUX2_X1 U14498 ( .A(n12735), .B(n12736), .S(n12731), .Z(n12692) );
  INV_X1 U14499 ( .A(n12692), .ZN(n12693) );
  OR3_X1 U14500 ( .A1(n12694), .A2(n12693), .A3(n13213), .ZN(n12702) );
  NAND2_X1 U14501 ( .A1(n12702), .A2(n12695), .ZN(n12697) );
  OR2_X1 U14502 ( .A1(n13185), .A2(n13201), .ZN(n12758) );
  INV_X1 U14503 ( .A(n12758), .ZN(n12701) );
  AOI21_X1 U14504 ( .B1(n12697), .B2(n12701), .A(n12699), .ZN(n12698) );
  MUX2_X1 U14505 ( .A(n12699), .B(n12698), .S(n12731), .Z(n12705) );
  NAND4_X1 U14506 ( .A1(n12702), .A2(n12728), .A3(n12701), .A4(n12700), .ZN(
        n12703) );
  INV_X1 U14507 ( .A(n13176), .ZN(n13170) );
  NAND2_X1 U14508 ( .A1(n12703), .A2(n13170), .ZN(n12704) );
  OR2_X1 U14509 ( .A1(n12705), .A2(n12704), .ZN(n12708) );
  MUX2_X1 U14510 ( .A(n12706), .B(n13158), .S(n12728), .Z(n12707) );
  NAND2_X1 U14511 ( .A1(n12708), .A2(n12707), .ZN(n12725) );
  INV_X1 U14512 ( .A(n12725), .ZN(n12720) );
  NAND2_X1 U14513 ( .A1(n12710), .A2(n12709), .ZN(n12712) );
  NAND2_X1 U14514 ( .A1(n12712), .A2(n12711), .ZN(n12713) );
  NAND2_X1 U14515 ( .A1(n12714), .A2(n12713), .ZN(n12715) );
  NAND3_X1 U14516 ( .A1(n12717), .A2(n12716), .A3(n12715), .ZN(n12719) );
  AND2_X1 U14517 ( .A1(n12719), .A2(n12718), .ZN(n12724) );
  OAI21_X1 U14518 ( .B1(n12760), .B2(n12720), .A(n12724), .ZN(n12721) );
  NAND2_X1 U14519 ( .A1(n12721), .A2(n13104), .ZN(n12723) );
  NAND2_X1 U14520 ( .A1(n12723), .A2(n12722), .ZN(n12730) );
  OAI211_X1 U14521 ( .C1(n12760), .C2(n12725), .A(n13104), .B(n12724), .ZN(
        n12727) );
  NAND2_X1 U14522 ( .A1(n12727), .A2(n12726), .ZN(n12729) );
  NAND2_X1 U14523 ( .A1(n12736), .A2(n12735), .ZN(n13224) );
  NOR2_X1 U14524 ( .A1(n12738), .A2(n12737), .ZN(n12742) );
  NAND4_X1 U14525 ( .A1(n12742), .A2(n12741), .A3(n12740), .A4(n16312), .ZN(
        n12749) );
  NOR2_X1 U14526 ( .A1(n12744), .A2(n12743), .ZN(n12747) );
  NAND4_X1 U14527 ( .A1(n12747), .A2(n12746), .A3(n10281), .A4(n12745), .ZN(
        n12748) );
  NOR2_X1 U14528 ( .A1(n12749), .A2(n12748), .ZN(n12753) );
  NAND4_X1 U14529 ( .A1(n12753), .A2(n12752), .A3(n12751), .A4(n12750), .ZN(
        n12754) );
  INV_X1 U14530 ( .A(n12796), .ZN(n12797) );
  NOR2_X1 U14531 ( .A1(n12754), .A2(n12797), .ZN(n12755) );
  NAND3_X1 U14532 ( .A1(n10287), .A2(n13297), .A3(n12755), .ZN(n12756) );
  OR4_X1 U14533 ( .A1(n13234), .A2(n13263), .A3(n12756), .A4(n13272), .ZN(
        n12757) );
  OR4_X1 U14534 ( .A1(n12758), .A2(n13213), .A3(n13224), .A4(n12757), .ZN(
        n12759) );
  INV_X1 U14535 ( .A(n13104), .ZN(n12761) );
  XNOR2_X1 U14536 ( .A(n12766), .B(n13086), .ZN(n12768) );
  NAND3_X1 U14537 ( .A1(n12771), .A2(n12770), .A3(n13036), .ZN(n12772) );
  OAI211_X1 U14538 ( .C1(n12773), .C2(n12775), .A(n12772), .B(P3_B_REG_SCAN_IN), .ZN(n12774) );
  OAI21_X1 U14539 ( .B1(n12776), .B2(n12775), .A(n12774), .ZN(P3_U3296) );
  NAND2_X1 U14540 ( .A1(n12778), .A2(n16518), .ZN(n12786) );
  OAI22_X1 U14541 ( .A1(n12781), .A2(n12780), .B1(n12779), .B2(n16490), .ZN(
        n12784) );
  NOR2_X1 U14542 ( .A1(n16522), .A2(n12782), .ZN(n12783) );
  AOI211_X1 U14543 ( .C1(n16522), .C2(P1_REG2_REG_29__SCAN_IN), .A(n12784), 
        .B(n12783), .ZN(n12785) );
  OAI211_X1 U14544 ( .C1(n15191), .C2(n16512), .A(n12786), .B(n12785), .ZN(
        n12787) );
  AOI21_X1 U14545 ( .B1(n12788), .B2(n15537), .A(n12787), .ZN(n12789) );
  OAI21_X1 U14546 ( .B1(n12777), .B2(n15592), .A(n12789), .ZN(P1_U3356) );
  INV_X1 U14547 ( .A(n12790), .ZN(n15770) );
  OAI222_X1 U14548 ( .A1(n14787), .A2(n12792), .B1(n14783), .B2(n15770), .C1(
        P2_U3088), .C2(n12791), .ZN(P2_U3298) );
  MUX2_X1 U14549 ( .A(n12797), .B(n12796), .S(n11080), .Z(n12938) );
  INV_X1 U14550 ( .A(n12938), .ZN(n12798) );
  MUX2_X1 U14551 ( .A(n12800), .B(n12799), .S(n12821), .Z(n12801) );
  XNOR2_X1 U14552 ( .A(n13836), .B(n12821), .ZN(n12803) );
  XNOR2_X1 U14553 ( .A(n12803), .B(n12989), .ZN(n12859) );
  INV_X1 U14554 ( .A(n12859), .ZN(n12802) );
  NAND2_X1 U14555 ( .A1(n12856), .A2(n12804), .ZN(n12971) );
  XNOR2_X1 U14556 ( .A(n13832), .B(n12821), .ZN(n12805) );
  XNOR2_X1 U14557 ( .A(n12805), .B(n12903), .ZN(n12970) );
  INV_X1 U14558 ( .A(n12805), .ZN(n12806) );
  XNOR2_X1 U14559 ( .A(n12897), .B(n12821), .ZN(n12807) );
  XNOR2_X1 U14560 ( .A(n12807), .B(n12988), .ZN(n12899) );
  INV_X1 U14561 ( .A(n12807), .ZN(n12808) );
  NAND2_X1 U14562 ( .A1(n12808), .A2(n12988), .ZN(n12809) );
  XNOR2_X1 U14563 ( .A(n13824), .B(n12821), .ZN(n12810) );
  XNOR2_X1 U14564 ( .A(n12810), .B(n13275), .ZN(n12907) );
  NAND2_X1 U14565 ( .A1(n12810), .A2(n12958), .ZN(n12811) );
  XNOR2_X1 U14566 ( .A(n13820), .B(n12821), .ZN(n12812) );
  XNOR2_X1 U14567 ( .A(n12812), .B(n13226), .ZN(n12952) );
  NAND2_X1 U14568 ( .A1(n12812), .A2(n13252), .ZN(n12813) );
  NAND2_X1 U14569 ( .A1(n12951), .A2(n12813), .ZN(n12878) );
  XNOR2_X1 U14570 ( .A(n12875), .B(n12821), .ZN(n12814) );
  XNOR2_X1 U14571 ( .A(n12814), .B(n12987), .ZN(n12877) );
  INV_X1 U14572 ( .A(n12814), .ZN(n12815) );
  NAND2_X1 U14573 ( .A1(n12815), .A2(n12987), .ZN(n12816) );
  XNOR2_X1 U14574 ( .A(n13216), .B(n12821), .ZN(n12818) );
  XNOR2_X1 U14575 ( .A(n12818), .B(n13227), .ZN(n12925) );
  INV_X1 U14576 ( .A(n12925), .ZN(n12817) );
  NAND2_X1 U14577 ( .A1(n12818), .A2(n13227), .ZN(n12819) );
  XOR2_X1 U14578 ( .A(n12821), .B(n13201), .Z(n12884) );
  INV_X1 U14579 ( .A(n12820), .ZN(n12823) );
  MUX2_X1 U14580 ( .A(n12823), .B(n12822), .S(n12821), .Z(n12824) );
  XNOR2_X1 U14581 ( .A(n13193), .B(n12821), .ZN(n12826) );
  NAND2_X1 U14582 ( .A1(n12943), .A2(n12867), .ZN(n12829) );
  INV_X1 U14583 ( .A(n12825), .ZN(n12827) );
  NAND2_X1 U14584 ( .A1(n12827), .A2(n12826), .ZN(n12828) );
  NAND2_X1 U14585 ( .A1(n12829), .A2(n12828), .ZN(n12830) );
  XNOR2_X1 U14586 ( .A(n13400), .B(n11080), .ZN(n12831) );
  XNOR2_X1 U14587 ( .A(n13164), .B(n12821), .ZN(n12833) );
  NAND2_X1 U14588 ( .A1(n12833), .A2(n12891), .ZN(n12834) );
  NAND2_X1 U14589 ( .A1(n12835), .A2(n12834), .ZN(n12889) );
  XNOR2_X1 U14590 ( .A(n13330), .B(n12821), .ZN(n12836) );
  NAND2_X1 U14591 ( .A1(n12889), .A2(n12890), .ZN(n12838) );
  NAND2_X1 U14592 ( .A1(n12836), .A2(n12915), .ZN(n12837) );
  XNOR2_X1 U14593 ( .A(n13326), .B(n12821), .ZN(n12839) );
  XNOR2_X1 U14594 ( .A(n10225), .B(n12821), .ZN(n12840) );
  XNOR2_X1 U14595 ( .A(n13104), .B(n12821), .ZN(n12841) );
  AOI22_X1 U14596 ( .A1(n13114), .A2(n12978), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12843) );
  NAND2_X1 U14597 ( .A1(n8270), .A2(n12959), .ZN(n12842) );
  OAI211_X1 U14598 ( .C1(n13109), .C2(n12954), .A(n12843), .B(n12842), .ZN(
        n12844) );
  AOI21_X1 U14599 ( .B1(n13113), .B2(n12966), .A(n12844), .ZN(n12845) );
  INV_X1 U14600 ( .A(n12846), .ZN(n12847) );
  OAI222_X1 U14601 ( .A1(P3_U3151), .A2(n7904), .B1(n13850), .B2(n14226), .C1(
        n13853), .C2(n12847), .ZN(P3_U3265) );
  INV_X1 U14602 ( .A(n12848), .ZN(n12849) );
  XNOR2_X1 U14603 ( .A(n12850), .B(n12849), .ZN(n12855) );
  AOI22_X1 U14604 ( .A1(n12983), .A2(n12959), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12852) );
  NAND2_X1 U14605 ( .A1(n13127), .A2(n12978), .ZN(n12851) );
  OAI211_X1 U14606 ( .C1(n13125), .C2(n12954), .A(n12852), .B(n12851), .ZN(
        n12853) );
  AOI21_X1 U14607 ( .B1(n10225), .B2(n12966), .A(n12853), .ZN(n12854) );
  OAI21_X1 U14608 ( .B1(n12855), .B2(n12969), .A(n12854), .ZN(P3_U3154) );
  INV_X1 U14609 ( .A(n12856), .ZN(n12857) );
  AOI21_X1 U14610 ( .B1(n12859), .B2(n12858), .A(n12857), .ZN(n12864) );
  INV_X1 U14611 ( .A(n13836), .ZN(n12862) );
  NOR2_X1 U14612 ( .A1(n12955), .A2(n13305), .ZN(n12861) );
  AOI22_X1 U14613 ( .A1(n12975), .A2(n12990), .B1(n12903), .B2(n13251), .ZN(
        n13302) );
  NAND2_X1 U14614 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n16207)
         );
  OAI21_X1 U14615 ( .B1(n13302), .B2(n12976), .A(n16207), .ZN(n12860) );
  AOI211_X1 U14616 ( .C1(n12862), .C2(n12966), .A(n12861), .B(n12860), .ZN(
        n12863) );
  OAI21_X1 U14617 ( .B1(n12864), .B2(n12969), .A(n12863), .ZN(P3_U3155) );
  XNOR2_X1 U14618 ( .A(n12865), .B(n12985), .ZN(n12874) );
  INV_X1 U14619 ( .A(n12866), .ZN(n13175) );
  OR2_X1 U14620 ( .A1(n12891), .A2(n16352), .ZN(n12869) );
  OR2_X1 U14621 ( .A1(n12867), .A2(n16350), .ZN(n12868) );
  NAND2_X1 U14622 ( .A1(n12869), .A2(n12868), .ZN(n13172) );
  AOI22_X1 U14623 ( .A1(n13172), .A2(n12870), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12871) );
  OAI21_X1 U14624 ( .B1(n13175), .B2(n12955), .A(n12871), .ZN(n12872) );
  AOI21_X1 U14625 ( .B1(n13400), .B2(n12966), .A(n12872), .ZN(n12873) );
  OAI21_X1 U14626 ( .B1(n12874), .B2(n12969), .A(n12873), .ZN(P3_U3156) );
  INV_X1 U14627 ( .A(n12875), .ZN(n13816) );
  OAI211_X1 U14628 ( .C1(n12878), .C2(n12877), .A(n12876), .B(n7876), .ZN(
        n12882) );
  NAND2_X1 U14629 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13083)
         );
  OAI21_X1 U14630 ( .B1(n12954), .B2(n13227), .A(n13083), .ZN(n12880) );
  NOR2_X1 U14631 ( .A1(n12955), .A2(n13228), .ZN(n12879) );
  AOI211_X1 U14632 ( .C1(n12959), .C2(n13252), .A(n12880), .B(n12879), .ZN(
        n12881) );
  OAI211_X1 U14633 ( .C1(n13816), .C2(n12981), .A(n12882), .B(n12881), .ZN(
        P3_U3159) );
  XOR2_X1 U14634 ( .A(n12884), .B(n12883), .Z(n12888) );
  AOI22_X1 U14635 ( .A1(n12944), .A2(n13251), .B1(n12975), .B2(n12986), .ZN(
        n13203) );
  OAI22_X1 U14636 ( .A1(n13203), .A2(n12976), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13666), .ZN(n12885) );
  AOI21_X1 U14637 ( .B1(n13205), .B2(n12978), .A(n12885), .ZN(n12887) );
  NAND2_X1 U14638 ( .A1(n13349), .A2(n12966), .ZN(n12886) );
  OAI211_X1 U14639 ( .C1(n12888), .C2(n12969), .A(n12887), .B(n12886), .ZN(
        P3_U3163) );
  XOR2_X1 U14640 ( .A(n12890), .B(n12889), .Z(n12896) );
  NOR2_X1 U14641 ( .A1(n12891), .A2(n16350), .ZN(n12892) );
  AOI21_X1 U14642 ( .B1(n12983), .B2(n13251), .A(n12892), .ZN(n13146) );
  AOI22_X1 U14643 ( .A1(n13148), .A2(n12978), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12893) );
  OAI21_X1 U14644 ( .B1(n13146), .B2(n12976), .A(n12893), .ZN(n12894) );
  AOI21_X1 U14645 ( .B1(n13330), .B2(n12966), .A(n12894), .ZN(n12895) );
  OAI21_X1 U14646 ( .B1(n12896), .B2(n12969), .A(n12895), .ZN(P3_U3165) );
  INV_X1 U14647 ( .A(n12897), .ZN(n13828) );
  OAI211_X1 U14648 ( .C1(n12900), .C2(n12899), .A(n12898), .B(n7876), .ZN(
        n12905) );
  NAND2_X1 U14649 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n16243)
         );
  OAI21_X1 U14650 ( .B1(n12954), .B2(n13275), .A(n16243), .ZN(n12902) );
  NOR2_X1 U14651 ( .A1(n12955), .A2(n13276), .ZN(n12901) );
  AOI211_X1 U14652 ( .C1(n12959), .C2(n12903), .A(n12902), .B(n12901), .ZN(
        n12904) );
  OAI211_X1 U14653 ( .C1(n13828), .C2(n12981), .A(n12905), .B(n12904), .ZN(
        P3_U3166) );
  OAI211_X1 U14654 ( .C1(n12908), .C2(n12907), .A(n12906), .B(n7876), .ZN(
        n12912) );
  NAND2_X1 U14655 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n16260)
         );
  OAI21_X1 U14656 ( .B1(n12954), .B2(n13226), .A(n16260), .ZN(n12910) );
  NOR2_X1 U14657 ( .A1(n12955), .A2(n13257), .ZN(n12909) );
  AOI211_X1 U14658 ( .C1(n12959), .C2(n12988), .A(n12910), .B(n12909), .ZN(
        n12911) );
  OAI211_X1 U14659 ( .C1(n12981), .C2(n13824), .A(n12912), .B(n12911), .ZN(
        P3_U3168) );
  XOR2_X1 U14660 ( .A(n12914), .B(n12913), .Z(n12921) );
  OR2_X1 U14661 ( .A1(n12915), .A2(n16352), .ZN(n12917) );
  NAND2_X1 U14662 ( .A1(n12985), .A2(n12975), .ZN(n12916) );
  AND2_X1 U14663 ( .A1(n12917), .A2(n12916), .ZN(n13154) );
  AOI22_X1 U14664 ( .A1(n13165), .A2(n12978), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12918) );
  OAI21_X1 U14665 ( .B1(n13154), .B2(n12976), .A(n12918), .ZN(n12919) );
  AOI21_X1 U14666 ( .B1(n13164), .B2(n12966), .A(n12919), .ZN(n12920) );
  OAI21_X1 U14667 ( .B1(n12921), .B2(n12969), .A(n12920), .ZN(P3_U3169) );
  INV_X1 U14668 ( .A(n12922), .ZN(n12923) );
  AOI21_X1 U14669 ( .B1(n12925), .B2(n12924), .A(n12923), .ZN(n12930) );
  AOI22_X1 U14670 ( .A1(n12945), .A2(n13251), .B1(n12987), .B2(n12975), .ZN(
        n13214) );
  INV_X1 U14671 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n12926) );
  OAI22_X1 U14672 ( .A1(n13214), .A2(n12976), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12926), .ZN(n12927) );
  AOI21_X1 U14673 ( .B1(n13217), .B2(n12978), .A(n12927), .ZN(n12929) );
  NAND2_X1 U14674 ( .A1(n13216), .A2(n12966), .ZN(n12928) );
  OAI211_X1 U14675 ( .C1(n12930), .C2(n12969), .A(n12929), .B(n12928), .ZN(
        P3_U3173) );
  INV_X1 U14676 ( .A(n16594), .ZN(n12941) );
  INV_X1 U14677 ( .A(n12931), .ZN(n12932) );
  NAND2_X1 U14678 ( .A1(n12978), .A2(n12932), .ZN(n12933) );
  NAND2_X1 U14679 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n16201)
         );
  OAI211_X1 U14680 ( .C1(n12934), .C2(n12976), .A(n12933), .B(n16201), .ZN(
        n12940) );
  INV_X1 U14681 ( .A(n12935), .ZN(n12936) );
  AOI211_X1 U14682 ( .C1(n12938), .C2(n12937), .A(n12969), .B(n12936), .ZN(
        n12939) );
  AOI211_X1 U14683 ( .C1(n12941), .C2(n12966), .A(n12940), .B(n12939), .ZN(
        n12942) );
  INV_X1 U14684 ( .A(n12942), .ZN(P3_U3174) );
  XNOR2_X1 U14685 ( .A(n12943), .B(n12944), .ZN(n12950) );
  AOI22_X1 U14686 ( .A1(n12945), .A2(n12959), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12947) );
  NAND2_X1 U14687 ( .A1(n12978), .A2(n13194), .ZN(n12946) );
  OAI211_X1 U14688 ( .C1(n13188), .C2(n12954), .A(n12947), .B(n12946), .ZN(
        n12948) );
  AOI21_X1 U14689 ( .B1(n13193), .B2(n12966), .A(n12948), .ZN(n12949) );
  OAI21_X1 U14690 ( .B1(n12950), .B2(n12969), .A(n12949), .ZN(P3_U3175) );
  OAI211_X1 U14691 ( .C1(n12953), .C2(n12952), .A(n12951), .B(n7876), .ZN(
        n12961) );
  NAND2_X1 U14692 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13064)
         );
  OAI21_X1 U14693 ( .B1(n12954), .B2(n13237), .A(n13064), .ZN(n12957) );
  NOR2_X1 U14694 ( .A1(n12955), .A2(n13243), .ZN(n12956) );
  AOI211_X1 U14695 ( .C1(n12959), .C2(n12958), .A(n12957), .B(n12956), .ZN(
        n12960) );
  OAI211_X1 U14696 ( .C1(n13820), .C2(n12981), .A(n12961), .B(n12960), .ZN(
        P3_U3178) );
  XOR2_X1 U14697 ( .A(n12963), .B(n12962), .Z(n12968) );
  AOI22_X1 U14698 ( .A1(n8270), .A2(n13251), .B1(n12975), .B2(n12984), .ZN(
        n13134) );
  AOI22_X1 U14699 ( .A1(n13136), .A2(n12978), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12964) );
  OAI21_X1 U14700 ( .B1(n13134), .B2(n12976), .A(n12964), .ZN(n12965) );
  AOI21_X1 U14701 ( .B1(n13326), .B2(n12966), .A(n12965), .ZN(n12967) );
  OAI21_X1 U14702 ( .B1(n12968), .B2(n12969), .A(n12967), .ZN(P3_U3180) );
  AOI21_X1 U14703 ( .B1(n12971), .B2(n12970), .A(n12969), .ZN(n12973) );
  NAND2_X1 U14704 ( .A1(n12973), .A2(n12972), .ZN(n12980) );
  INV_X1 U14705 ( .A(n12974), .ZN(n13290) );
  AOI22_X1 U14706 ( .A1(n12988), .A2(n13251), .B1(n12975), .B2(n12989), .ZN(
        n13288) );
  NAND2_X1 U14707 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n16225)
         );
  OAI21_X1 U14708 ( .B1(n13288), .B2(n12976), .A(n16225), .ZN(n12977) );
  AOI21_X1 U14709 ( .B1(n13290), .B2(n12978), .A(n12977), .ZN(n12979) );
  OAI211_X1 U14710 ( .C1(n12981), .C2(n13832), .A(n12980), .B(n12979), .ZN(
        P3_U3181) );
  MUX2_X1 U14711 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12982), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14712 ( .A(n8270), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12998), .Z(
        P3_U3518) );
  MUX2_X1 U14713 ( .A(n12983), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12998), .Z(
        P3_U3517) );
  MUX2_X1 U14714 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12984), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14715 ( .A(n12985), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12998), .Z(
        P3_U3514) );
  MUX2_X1 U14716 ( .A(n12986), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12998), .Z(
        P3_U3511) );
  MUX2_X1 U14717 ( .A(n12987), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12998), .Z(
        P3_U3510) );
  MUX2_X1 U14718 ( .A(n13252), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12998), .Z(
        P3_U3509) );
  MUX2_X1 U14719 ( .A(n12988), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12998), .Z(
        P3_U3507) );
  MUX2_X1 U14720 ( .A(n12989), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12998), .Z(
        P3_U3505) );
  MUX2_X1 U14721 ( .A(n12990), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12998), .Z(
        P3_U3504) );
  MUX2_X1 U14722 ( .A(n12991), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12998), .Z(
        P3_U3502) );
  MUX2_X1 U14723 ( .A(n12992), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12998), .Z(
        P3_U3500) );
  MUX2_X1 U14724 ( .A(n12993), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12998), .Z(
        P3_U3499) );
  MUX2_X1 U14725 ( .A(n12994), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12998), .Z(
        P3_U3498) );
  MUX2_X1 U14726 ( .A(n12995), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12998), .Z(
        P3_U3497) );
  MUX2_X1 U14727 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12996), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14728 ( .A(n9810), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12998), .Z(
        P3_U3494) );
  MUX2_X1 U14729 ( .A(n9794), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12998), .Z(
        P3_U3493) );
  MUX2_X1 U14730 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12997), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14731 ( .A(n12999), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12998), .Z(
        P3_U3491) );
  AND2_X1 U14732 ( .A1(n16274), .A2(n16263), .ZN(n13001) );
  NAND2_X1 U14733 ( .A1(n16277), .A2(n13001), .ZN(n13000) );
  AOI21_X1 U14734 ( .B1(n13000), .B2(n13002), .A(n16269), .ZN(n13007) );
  INV_X1 U14735 ( .A(n13001), .ZN(n13004) );
  INV_X1 U14736 ( .A(n13002), .ZN(n13003) );
  NAND2_X1 U14737 ( .A1(n13004), .A2(n13003), .ZN(n13006) );
  MUX2_X1 U14738 ( .A(n13007), .B(n13006), .S(n13005), .Z(n13011) );
  AOI22_X1 U14739 ( .A1(n16259), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n13010) );
  NAND2_X1 U14740 ( .A1(n16194), .A2(n13008), .ZN(n13009) );
  NAND3_X1 U14741 ( .A1(n13011), .A2(n13010), .A3(n13009), .ZN(P3_U3182) );
  INV_X1 U14742 ( .A(n13055), .ZN(n16232) );
  INV_X1 U14743 ( .A(n13052), .ZN(n16187) );
  INV_X1 U14744 ( .A(n13015), .ZN(n13014) );
  NOR2_X1 U14745 ( .A1(n16152), .A2(n13014), .ZN(n13016) );
  OR2_X1 U14746 ( .A1(n16166), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n13017) );
  NAND2_X1 U14747 ( .A1(n16166), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n13031) );
  NAND2_X1 U14748 ( .A1(n13017), .A2(n13031), .ZN(n13030) );
  OR2_X2 U14749 ( .A1(n16177), .A2(n13030), .ZN(n16178) );
  NOR2_X1 U14750 ( .A1(n16187), .A2(n7518), .ZN(n13018) );
  INV_X1 U14751 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n16600) );
  XNOR2_X1 U14752 ( .A(n16204), .B(P3_REG1_REG_14__SCAN_IN), .ZN(n16217) );
  OR2_X2 U14753 ( .A1(n16216), .A2(n16217), .ZN(n16214) );
  NAND2_X1 U14754 ( .A1(n16204), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13019) );
  INV_X1 U14755 ( .A(n13021), .ZN(n13020) );
  XNOR2_X1 U14756 ( .A(n16250), .B(n13370), .ZN(n16252) );
  AOI21_X1 U14757 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n13058), .A(n16251), 
        .ZN(n13023) );
  XNOR2_X1 U14758 ( .A(n16268), .B(n13023), .ZN(n16272) );
  NAND2_X1 U14759 ( .A1(n13065), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n13069) );
  OAI21_X1 U14760 ( .B1(n13065), .B2(P3_REG1_REG_18__SCAN_IN), .A(n13069), 
        .ZN(n13024) );
  AOI21_X1 U14761 ( .B1(n7576), .B2(n13024), .A(n13070), .ZN(n13068) );
  MUX2_X1 U14762 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13036), .Z(n13042) );
  MUX2_X1 U14763 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13036), .Z(n13040) );
  MUX2_X1 U14764 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n13036), .Z(n13038) );
  MUX2_X1 U14765 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n13036), .Z(n13034) );
  MUX2_X1 U14766 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13036), .Z(n13033) );
  OAI21_X1 U14767 ( .B1(n13026), .B2(n13044), .A(n13025), .ZN(n16154) );
  MUX2_X1 U14768 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13036), .Z(n13027) );
  XNOR2_X1 U14769 ( .A(n13027), .B(n16152), .ZN(n16153) );
  INV_X1 U14770 ( .A(n13027), .ZN(n13028) );
  AOI22_X1 U14771 ( .A1(n16154), .A2(n16153), .B1(n16152), .B2(n13028), .ZN(
        n16173) );
  XNOR2_X1 U14772 ( .A(n16166), .B(n13029), .ZN(n16169) );
  INV_X1 U14773 ( .A(n13030), .ZN(n16179) );
  MUX2_X1 U14774 ( .A(n16169), .B(n16179), .S(n13036), .Z(n16172) );
  NAND2_X1 U14775 ( .A1(n16173), .A2(n16172), .ZN(n16171) );
  NAND2_X1 U14776 ( .A1(n16166), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n13050) );
  MUX2_X1 U14777 ( .A(n13050), .B(n13031), .S(n13036), .Z(n13032) );
  XNOR2_X1 U14778 ( .A(n13033), .B(n16187), .ZN(n16189) );
  NAND2_X1 U14779 ( .A1(n16190), .A2(n16189), .ZN(n16188) );
  OAI21_X1 U14780 ( .B1(n13033), .B2(n13052), .A(n16188), .ZN(n16210) );
  XNOR2_X1 U14781 ( .A(n13034), .B(n16204), .ZN(n16211) );
  NOR2_X1 U14782 ( .A1(n16210), .A2(n16211), .ZN(n16209) );
  AOI21_X1 U14783 ( .B1(n13034), .B2(n16204), .A(n16209), .ZN(n13035) );
  INV_X1 U14784 ( .A(n13035), .ZN(n13037) );
  XNOR2_X1 U14785 ( .A(n13035), .B(n16232), .ZN(n16229) );
  MUX2_X1 U14786 ( .A(n16224), .B(n16234), .S(n13036), .Z(n16228) );
  NOR2_X1 U14787 ( .A1(n16229), .A2(n16228), .ZN(n16227) );
  XNOR2_X1 U14788 ( .A(n13038), .B(n13058), .ZN(n16246) );
  XNOR2_X1 U14789 ( .A(n13040), .B(n13039), .ZN(n16264) );
  AOI21_X1 U14790 ( .B1(n13040), .B2(n13039), .A(n16262), .ZN(n13078) );
  XNOR2_X1 U14791 ( .A(n13078), .B(n13077), .ZN(n13041) );
  NOR2_X1 U14792 ( .A1(n13041), .A2(n13042), .ZN(n13076) );
  AOI21_X1 U14793 ( .B1(n13042), .B2(n13041), .A(n13076), .ZN(n13043) );
  NOR2_X1 U14794 ( .A1(n13043), .A2(n16263), .ZN(n13067) );
  NAND2_X1 U14795 ( .A1(n13044), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n13046) );
  NAND2_X1 U14796 ( .A1(n13046), .A2(n13045), .ZN(n13048) );
  NAND2_X1 U14797 ( .A1(n13047), .A2(n13048), .ZN(n13049) );
  XNOR2_X1 U14798 ( .A(n13048), .B(n16152), .ZN(n16156) );
  NAND2_X1 U14799 ( .A1(P3_REG2_REG_11__SCAN_IN), .A2(n16156), .ZN(n16155) );
  NAND2_X1 U14800 ( .A1(n13052), .A2(n13051), .ZN(n13053) );
  INV_X1 U14801 ( .A(n16206), .ZN(n13054) );
  NOR2_X1 U14802 ( .A1(n16232), .A2(n13056), .ZN(n13057) );
  XOR2_X1 U14803 ( .A(n13056), .B(n13055), .Z(n16223) );
  NOR2_X1 U14804 ( .A1(n16224), .A2(n16223), .ZN(n16222) );
  AOI22_X1 U14805 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n16250), .B1(n13058), 
        .B2(n13277), .ZN(n16241) );
  NOR2_X1 U14806 ( .A1(n16242), .A2(n16241), .ZN(n16240) );
  NOR2_X1 U14807 ( .A1(n16268), .A2(n13059), .ZN(n13060) );
  XNOR2_X1 U14808 ( .A(n16268), .B(n13059), .ZN(n16258) );
  NOR2_X1 U14809 ( .A1(n13258), .A2(n16258), .ZN(n16257) );
  NAND2_X1 U14810 ( .A1(n13065), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n13071) );
  OAI21_X1 U14811 ( .B1(n13065), .B2(P3_REG2_REG_18__SCAN_IN), .A(n13071), 
        .ZN(n13061) );
  NAND2_X1 U14812 ( .A1(n16259), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n13063) );
  OAI211_X1 U14813 ( .C1(n16142), .C2(n13065), .A(n13064), .B(n13063), .ZN(
        n13066) );
  XNOR2_X1 U14814 ( .A(n13086), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13079) );
  INV_X1 U14815 ( .A(n13071), .ZN(n13072) );
  NOR2_X1 U14816 ( .A1(n13073), .A2(n13072), .ZN(n13075) );
  XNOR2_X1 U14817 ( .A(n13086), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13080) );
  INV_X1 U14818 ( .A(n13080), .ZN(n13074) );
  XNOR2_X1 U14819 ( .A(n13075), .B(n13074), .ZN(n13088) );
  AOI21_X1 U14820 ( .B1(n13078), .B2(n13077), .A(n13076), .ZN(n13082) );
  MUX2_X1 U14821 ( .A(n13080), .B(n13079), .S(n7432), .Z(n13081) );
  OAI21_X1 U14822 ( .B1(n16151), .B2(n13084), .A(n13083), .ZN(n13085) );
  AOI21_X1 U14823 ( .B1(n13086), .B2(n16269), .A(n13085), .ZN(n13087) );
  NOR2_X1 U14824 ( .A1(n13091), .A2(n13090), .ZN(n13381) );
  NOR2_X1 U14825 ( .A1(n13092), .A2(n16360), .ZN(n13097) );
  NOR3_X1 U14826 ( .A1(n13381), .A2(n13292), .A3(n13097), .ZN(n13095) );
  NOR2_X1 U14827 ( .A1(n13310), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13093) );
  OAI22_X1 U14828 ( .A1(n12575), .A2(n13304), .B1(n13095), .B2(n13093), .ZN(
        P3_U3202) );
  INV_X1 U14829 ( .A(n13384), .ZN(n13317) );
  NOR2_X1 U14830 ( .A1(n13310), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13094) );
  OAI22_X1 U14831 ( .A1(n13317), .A2(n13304), .B1(n13095), .B2(n13094), .ZN(
        P3_U3203) );
  INV_X1 U14832 ( .A(n13096), .ZN(n13103) );
  AOI21_X1 U14833 ( .B1(n16369), .B2(P3_REG2_REG_29__SCAN_IN), .A(n13097), 
        .ZN(n13098) );
  OAI21_X1 U14834 ( .B1(n13099), .B2(n13304), .A(n13098), .ZN(n13100) );
  AOI21_X1 U14835 ( .B1(n13101), .B2(n13310), .A(n13100), .ZN(n13102) );
  OAI21_X1 U14836 ( .B1(n13103), .B2(n13313), .A(n13102), .ZN(P3_U3204) );
  NAND2_X1 U14837 ( .A1(n13105), .A2(n13104), .ZN(n13106) );
  NAND2_X1 U14838 ( .A1(n13106), .A2(n13299), .ZN(n13107) );
  OAI22_X1 U14839 ( .A1(n13109), .A2(n16352), .B1(n13108), .B2(n16350), .ZN(
        n13110) );
  INV_X1 U14840 ( .A(n13110), .ZN(n13111) );
  INV_X1 U14841 ( .A(n13113), .ZN(n13390) );
  AOI22_X1 U14842 ( .A1(n13114), .A2(n13291), .B1(n16369), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13115) );
  OAI21_X1 U14843 ( .B1(n13390), .B2(n13304), .A(n13115), .ZN(n13116) );
  AOI21_X1 U14844 ( .B1(n13319), .B2(n13310), .A(n13116), .ZN(n13117) );
  OAI21_X1 U14845 ( .B1(n13318), .B2(n13313), .A(n13117), .ZN(P3_U3205) );
  INV_X1 U14846 ( .A(n13120), .ZN(n13121) );
  AOI21_X1 U14847 ( .B1(n13123), .B2(n13122), .A(n13121), .ZN(n13124) );
  OAI222_X1 U14848 ( .A1(n16350), .A2(n13126), .B1(n16352), .B2(n13125), .C1(
        n16349), .C2(n13124), .ZN(n13322) );
  AOI22_X1 U14849 ( .A1(n13127), .A2(n13291), .B1(n16369), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13128) );
  OAI21_X1 U14850 ( .B1(n8271), .B2(n13304), .A(n13128), .ZN(n13129) );
  AOI21_X1 U14851 ( .B1(n13322), .B2(n13310), .A(n13129), .ZN(n13130) );
  OAI21_X1 U14852 ( .B1(n13313), .B2(n13324), .A(n13130), .ZN(P3_U3206) );
  XOR2_X1 U14853 ( .A(n13131), .B(n13132), .Z(n13328) );
  XNOR2_X1 U14854 ( .A(n13133), .B(n13132), .ZN(n13135) );
  OAI21_X1 U14855 ( .B1(n13135), .B2(n16349), .A(n13134), .ZN(n13325) );
  INV_X1 U14856 ( .A(n13326), .ZN(n13138) );
  AOI22_X1 U14857 ( .A1(n13136), .A2(n13291), .B1(n13292), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13137) );
  OAI21_X1 U14858 ( .B1(n13138), .B2(n13304), .A(n13137), .ZN(n13139) );
  AOI21_X1 U14859 ( .B1(n13325), .B2(n13310), .A(n13139), .ZN(n13140) );
  OAI21_X1 U14860 ( .B1(n13328), .B2(n13313), .A(n13140), .ZN(P3_U3207) );
  OAI21_X1 U14861 ( .B1(n13143), .B2(n13142), .A(n13141), .ZN(n13332) );
  OAI211_X1 U14862 ( .C1(n7534), .C2(n13145), .A(n13299), .B(n13144), .ZN(
        n13147) );
  NAND2_X1 U14863 ( .A1(n13147), .A2(n13146), .ZN(n13329) );
  INV_X1 U14864 ( .A(n13330), .ZN(n13150) );
  AOI22_X1 U14865 ( .A1(n13148), .A2(n13291), .B1(n16369), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13149) );
  OAI21_X1 U14866 ( .B1(n13150), .B2(n13304), .A(n13149), .ZN(n13151) );
  AOI21_X1 U14867 ( .B1(n13329), .B2(n13310), .A(n13151), .ZN(n13152) );
  OAI21_X1 U14868 ( .B1(n13313), .B2(n13332), .A(n13152), .ZN(P3_U3208) );
  XNOR2_X1 U14869 ( .A(n13153), .B(n13162), .ZN(n13156) );
  INV_X1 U14870 ( .A(n13154), .ZN(n13155) );
  AOI21_X1 U14871 ( .B1(n13156), .B2(n13299), .A(n13155), .ZN(n13334) );
  OR2_X1 U14872 ( .A1(n13157), .A2(n13176), .ZN(n13178) );
  NAND2_X1 U14873 ( .A1(n13178), .A2(n13158), .ZN(n13163) );
  AND2_X1 U14874 ( .A1(n13160), .A2(n13159), .ZN(n13161) );
  OAI21_X1 U14875 ( .B1(n13163), .B2(n13162), .A(n13161), .ZN(n13333) );
  INV_X1 U14876 ( .A(n13333), .ZN(n13168) );
  INV_X1 U14877 ( .A(n13164), .ZN(n13397) );
  AOI22_X1 U14878 ( .A1(n13291), .A2(n13165), .B1(n16369), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n13166) );
  OAI21_X1 U14879 ( .B1(n13397), .B2(n13304), .A(n13166), .ZN(n13167) );
  AOI21_X1 U14880 ( .B1(n13168), .B2(n13266), .A(n13167), .ZN(n13169) );
  OAI21_X1 U14881 ( .B1(n16369), .B2(n13334), .A(n13169), .ZN(P3_U3209) );
  XNOR2_X1 U14882 ( .A(n13171), .B(n13170), .ZN(n13173) );
  AOI21_X1 U14883 ( .B1(n13173), .B2(n13299), .A(n13172), .ZN(n13338) );
  INV_X1 U14884 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n13174) );
  OAI22_X1 U14885 ( .A1(n13175), .A2(n16360), .B1(n13307), .B2(n13174), .ZN(
        n13180) );
  NAND2_X1 U14886 ( .A1(n13157), .A2(n13176), .ZN(n13177) );
  NAND2_X1 U14887 ( .A1(n13178), .A2(n13177), .ZN(n13339) );
  NOR2_X1 U14888 ( .A1(n13339), .A2(n13313), .ZN(n13179) );
  AOI211_X1 U14889 ( .C1(n13260), .C2(n13400), .A(n13180), .B(n13179), .ZN(
        n13181) );
  OAI21_X1 U14890 ( .B1(n13292), .B2(n13338), .A(n13181), .ZN(P3_U3210) );
  INV_X1 U14891 ( .A(n13182), .ZN(n13183) );
  AOI21_X1 U14892 ( .B1(n13185), .B2(n13184), .A(n13183), .ZN(n13192) );
  XNOR2_X1 U14893 ( .A(n13186), .B(n13185), .ZN(n13190) );
  OAI22_X1 U14894 ( .A1(n13188), .A2(n16352), .B1(n13187), .B2(n16350), .ZN(
        n13189) );
  AOI21_X1 U14895 ( .B1(n13190), .B2(n13299), .A(n13189), .ZN(n13191) );
  OAI21_X1 U14896 ( .B1(n13192), .B2(n16541), .A(n13191), .ZN(n13343) );
  INV_X1 U14897 ( .A(n13343), .ZN(n13199) );
  INV_X1 U14898 ( .A(n13192), .ZN(n13344) );
  INV_X1 U14899 ( .A(n13193), .ZN(n13406) );
  AOI22_X1 U14900 ( .A1(n13292), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n13291), 
        .B2(n13194), .ZN(n13195) );
  OAI21_X1 U14901 ( .B1(n13406), .B2(n13304), .A(n13195), .ZN(n13196) );
  AOI21_X1 U14902 ( .B1(n13344), .B2(n13197), .A(n13196), .ZN(n13198) );
  OAI21_X1 U14903 ( .B1(n13199), .B2(n13292), .A(n13198), .ZN(P3_U3211) );
  XOR2_X1 U14904 ( .A(n13201), .B(n13200), .Z(n13351) );
  XNOR2_X1 U14905 ( .A(n13202), .B(n13201), .ZN(n13204) );
  OAI21_X1 U14906 ( .B1(n13204), .B2(n16349), .A(n13203), .ZN(n13348) );
  INV_X1 U14907 ( .A(n13349), .ZN(n13207) );
  AOI22_X1 U14908 ( .A1(n16369), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n13291), 
        .B2(n13205), .ZN(n13206) );
  OAI21_X1 U14909 ( .B1(n13207), .B2(n13304), .A(n13206), .ZN(n13208) );
  AOI21_X1 U14910 ( .B1(n13348), .B2(n13310), .A(n13208), .ZN(n13209) );
  OAI21_X1 U14911 ( .B1(n13351), .B2(n13313), .A(n13209), .ZN(P3_U3212) );
  XNOR2_X1 U14912 ( .A(n13211), .B(n13210), .ZN(n13353) );
  INV_X1 U14913 ( .A(n13353), .ZN(n13221) );
  OAI211_X1 U14914 ( .C1(n8505), .C2(n13213), .A(n13299), .B(n13212), .ZN(
        n13215) );
  NAND2_X1 U14915 ( .A1(n13215), .A2(n13214), .ZN(n13352) );
  INV_X1 U14916 ( .A(n13216), .ZN(n13812) );
  AOI22_X1 U14917 ( .A1(n16369), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n13291), 
        .B2(n13217), .ZN(n13218) );
  OAI21_X1 U14918 ( .B1(n13812), .B2(n13304), .A(n13218), .ZN(n13219) );
  AOI21_X1 U14919 ( .B1(n13352), .B2(n13310), .A(n13219), .ZN(n13220) );
  OAI21_X1 U14920 ( .B1(n13221), .B2(n13313), .A(n13220), .ZN(P3_U3213) );
  NAND2_X1 U14921 ( .A1(n13241), .A2(n13238), .ZN(n13222) );
  XOR2_X1 U14922 ( .A(n13222), .B(n13224), .Z(n13357) );
  INV_X1 U14923 ( .A(n13357), .ZN(n13233) );
  XOR2_X1 U14924 ( .A(n13224), .B(n13223), .Z(n13225) );
  OAI222_X1 U14925 ( .A1(n16352), .A2(n13227), .B1(n16350), .B2(n13226), .C1(
        n16349), .C2(n13225), .ZN(n13356) );
  NOR2_X1 U14926 ( .A1(n13816), .A2(n13304), .ZN(n13231) );
  OAI22_X1 U14927 ( .A1(n13307), .A2(n13229), .B1(n13228), .B2(n16360), .ZN(
        n13230) );
  AOI211_X1 U14928 ( .C1(n13356), .C2(n13310), .A(n13231), .B(n13230), .ZN(
        n13232) );
  OAI21_X1 U14929 ( .B1(n13313), .B2(n13233), .A(n13232), .ZN(P3_U3214) );
  XNOR2_X1 U14930 ( .A(n13235), .B(n13234), .ZN(n13236) );
  OAI222_X1 U14931 ( .A1(n16352), .A2(n13237), .B1(n16350), .B2(n13275), .C1(
        n13236), .C2(n16349), .ZN(n13360) );
  INV_X1 U14932 ( .A(n13360), .ZN(n13248) );
  INV_X1 U14933 ( .A(n13238), .ZN(n13242) );
  OAI22_X1 U14934 ( .A1(n13242), .A2(n13241), .B1(n13240), .B2(n13239), .ZN(
        n13361) );
  NOR2_X1 U14935 ( .A1(n13820), .A2(n13304), .ZN(n13246) );
  INV_X1 U14936 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13244) );
  OAI22_X1 U14937 ( .A1(n13307), .A2(n13244), .B1(n13243), .B2(n16360), .ZN(
        n13245) );
  AOI211_X1 U14938 ( .C1(n13361), .C2(n13266), .A(n13246), .B(n13245), .ZN(
        n13247) );
  OAI21_X1 U14939 ( .B1(n13248), .B2(n16369), .A(n13247), .ZN(P3_U3215) );
  XNOR2_X1 U14940 ( .A(n13249), .B(n13250), .ZN(n13256) );
  NAND2_X1 U14941 ( .A1(n13252), .A2(n13251), .ZN(n13253) );
  OAI21_X1 U14942 ( .B1(n13254), .B2(n16350), .A(n13253), .ZN(n13255) );
  AOI21_X1 U14943 ( .B1(n13256), .B2(n13299), .A(n13255), .ZN(n13366) );
  INV_X1 U14944 ( .A(n13824), .ZN(n13261) );
  OAI22_X1 U14945 ( .A1(n13307), .A2(n13258), .B1(n13257), .B2(n16360), .ZN(
        n13259) );
  AOI21_X1 U14946 ( .B1(n13261), .B2(n13260), .A(n13259), .ZN(n13268) );
  INV_X1 U14947 ( .A(n13262), .ZN(n13264) );
  NAND2_X1 U14948 ( .A1(n13264), .A2(n13263), .ZN(n13364) );
  NAND3_X1 U14949 ( .A1(n13364), .A2(n13266), .A3(n13265), .ZN(n13267) );
  OAI211_X1 U14950 ( .C1(n13366), .C2(n13292), .A(n13268), .B(n13267), .ZN(
        P3_U3216) );
  XNOR2_X1 U14951 ( .A(n13269), .B(n13270), .ZN(n13369) );
  INV_X1 U14952 ( .A(n13369), .ZN(n13281) );
  XNOR2_X1 U14953 ( .A(n13271), .B(n13272), .ZN(n13273) );
  OAI222_X1 U14954 ( .A1(n16352), .A2(n13275), .B1(n16350), .B2(n13274), .C1(
        n13273), .C2(n16349), .ZN(n13368) );
  NOR2_X1 U14955 ( .A1(n13828), .A2(n13304), .ZN(n13279) );
  OAI22_X1 U14956 ( .A1(n13307), .A2(n13277), .B1(n13276), .B2(n16360), .ZN(
        n13278) );
  AOI211_X1 U14957 ( .C1(n13368), .C2(n13310), .A(n13279), .B(n13278), .ZN(
        n13280) );
  OAI21_X1 U14958 ( .B1(n13313), .B2(n13281), .A(n13280), .ZN(P3_U3217) );
  OAI21_X1 U14959 ( .B1(n13283), .B2(n10287), .A(n13282), .ZN(n13373) );
  INV_X1 U14960 ( .A(n13373), .ZN(n13296) );
  NAND3_X1 U14961 ( .A1(n13284), .A2(n10287), .A3(n13285), .ZN(n13286) );
  NAND3_X1 U14962 ( .A1(n13287), .A2(n13299), .A3(n13286), .ZN(n13289) );
  NAND2_X1 U14963 ( .A1(n13289), .A2(n13288), .ZN(n13372) );
  AOI22_X1 U14964 ( .A1(n13292), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n13291), 
        .B2(n13290), .ZN(n13293) );
  OAI21_X1 U14965 ( .B1(n13832), .B2(n13304), .A(n13293), .ZN(n13294) );
  AOI21_X1 U14966 ( .B1(n13372), .B2(n13310), .A(n13294), .ZN(n13295) );
  OAI21_X1 U14967 ( .B1(n13296), .B2(n13313), .A(n13295), .ZN(P3_U3218) );
  XNOR2_X1 U14968 ( .A(n13298), .B(n13297), .ZN(n13376) );
  INV_X1 U14969 ( .A(n13376), .ZN(n13312) );
  OAI211_X1 U14970 ( .C1(n13301), .C2(n13300), .A(n13284), .B(n13299), .ZN(
        n13303) );
  NAND2_X1 U14971 ( .A1(n13303), .A2(n13302), .ZN(n13375) );
  NOR2_X1 U14972 ( .A1(n13836), .A2(n13304), .ZN(n13309) );
  OAI22_X1 U14973 ( .A1(n13307), .A2(n13306), .B1(n13305), .B2(n16360), .ZN(
        n13308) );
  AOI211_X1 U14974 ( .C1(n13375), .C2(n13310), .A(n13309), .B(n13308), .ZN(
        n13311) );
  OAI21_X1 U14975 ( .B1(n13313), .B2(n13312), .A(n13311), .ZN(P3_U3219) );
  NAND2_X1 U14976 ( .A1(n13381), .A2(n16601), .ZN(n13315) );
  NAND2_X1 U14977 ( .A1(n16599), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13314) );
  OAI211_X1 U14978 ( .C1(n12575), .C2(n13379), .A(n13315), .B(n13314), .ZN(
        P3_U3490) );
  NAND2_X1 U14979 ( .A1(n16599), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13316) );
  OAI211_X1 U14980 ( .C1(n13317), .C2(n13379), .A(n13316), .B(n13315), .ZN(
        P3_U3489) );
  INV_X1 U14981 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13321) );
  AOI21_X1 U14982 ( .B1(n16544), .B2(n10225), .A(n13322), .ZN(n13323) );
  OAI21_X1 U14983 ( .B1(n16414), .B2(n13324), .A(n13323), .ZN(n13391) );
  MUX2_X1 U14984 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13391), .S(n16568), .Z(
        P3_U3486) );
  AOI21_X1 U14985 ( .B1(n16544), .B2(n13326), .A(n13325), .ZN(n13327) );
  OAI21_X1 U14986 ( .B1(n13328), .B2(n16414), .A(n13327), .ZN(n13392) );
  MUX2_X1 U14987 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n13392), .S(n16568), .Z(
        P3_U3485) );
  AOI21_X1 U14988 ( .B1(n16544), .B2(n13330), .A(n13329), .ZN(n13331) );
  OAI21_X1 U14989 ( .B1(n16414), .B2(n13332), .A(n13331), .ZN(n13393) );
  MUX2_X1 U14990 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13393), .S(n16601), .Z(
        P3_U3484) );
  OR2_X1 U14991 ( .A1(n13333), .A2(n16414), .ZN(n13335) );
  AND2_X1 U14992 ( .A1(n13335), .A2(n13334), .ZN(n13395) );
  INV_X1 U14993 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13336) );
  MUX2_X1 U14994 ( .A(n13395), .B(n13336), .S(n16599), .Z(n13337) );
  OAI21_X1 U14995 ( .B1(n13397), .B2(n13379), .A(n13337), .ZN(P3_U3483) );
  OAI21_X1 U14996 ( .B1(n13339), .B2(n16414), .A(n13338), .ZN(n13398) );
  MUX2_X1 U14997 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n13398), .S(n16601), .Z(
        n13340) );
  AOI21_X1 U14998 ( .B1(n13341), .B2(n13400), .A(n13340), .ZN(n13342) );
  INV_X1 U14999 ( .A(n13342), .ZN(P3_U3482) );
  INV_X1 U15000 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13346) );
  INV_X1 U15001 ( .A(n16584), .ZN(n13345) );
  AOI21_X1 U15002 ( .B1(n13345), .B2(n13344), .A(n13343), .ZN(n13403) );
  MUX2_X1 U15003 ( .A(n13346), .B(n13403), .S(n16601), .Z(n13347) );
  OAI21_X1 U15004 ( .B1(n13406), .B2(n13379), .A(n13347), .ZN(P3_U3481) );
  AOI21_X1 U15005 ( .B1(n16544), .B2(n13349), .A(n13348), .ZN(n13350) );
  OAI21_X1 U15006 ( .B1(n13351), .B2(n16414), .A(n13350), .ZN(n13806) );
  MUX2_X1 U15007 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n13806), .S(n16601), .Z(
        P3_U3480) );
  AOI21_X1 U15008 ( .B1(n13353), .B2(n16597), .A(n13352), .ZN(n13809) );
  MUX2_X1 U15009 ( .A(n13354), .B(n13809), .S(n16601), .Z(n13355) );
  OAI21_X1 U15010 ( .B1(n13812), .B2(n13379), .A(n13355), .ZN(P3_U3479) );
  AOI21_X1 U15011 ( .B1(n13357), .B2(n16597), .A(n13356), .ZN(n13813) );
  MUX2_X1 U15012 ( .A(n13358), .B(n13813), .S(n16601), .Z(n13359) );
  OAI21_X1 U15013 ( .B1(n13816), .B2(n13379), .A(n13359), .ZN(P3_U3478) );
  INV_X1 U15014 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13362) );
  AOI21_X1 U15015 ( .B1(n16597), .B2(n13361), .A(n13360), .ZN(n13817) );
  MUX2_X1 U15016 ( .A(n13362), .B(n13817), .S(n16601), .Z(n13363) );
  OAI21_X1 U15017 ( .B1(n13820), .B2(n13379), .A(n13363), .ZN(P3_U3477) );
  NAND3_X1 U15018 ( .A1(n13364), .A2(n13265), .A3(n16597), .ZN(n13365) );
  AND2_X1 U15019 ( .A1(n13366), .A2(n13365), .ZN(n13822) );
  MUX2_X1 U15020 ( .A(n16271), .B(n13822), .S(n16601), .Z(n13367) );
  OAI21_X1 U15021 ( .B1(n13379), .B2(n13824), .A(n13367), .ZN(P3_U3476) );
  AOI21_X1 U15022 ( .B1(n13369), .B2(n16597), .A(n13368), .ZN(n13825) );
  MUX2_X1 U15023 ( .A(n13370), .B(n13825), .S(n16601), .Z(n13371) );
  OAI21_X1 U15024 ( .B1(n13828), .B2(n13379), .A(n13371), .ZN(P3_U3475) );
  AOI21_X1 U15025 ( .B1(n13373), .B2(n16597), .A(n13372), .ZN(n13829) );
  MUX2_X1 U15026 ( .A(n16234), .B(n13829), .S(n16601), .Z(n13374) );
  OAI21_X1 U15027 ( .B1(n13379), .B2(n13832), .A(n13374), .ZN(P3_U3474) );
  INV_X1 U15028 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13377) );
  AOI21_X1 U15029 ( .B1(n13376), .B2(n16597), .A(n13375), .ZN(n13833) );
  MUX2_X1 U15030 ( .A(n13377), .B(n13833), .S(n16601), .Z(n13378) );
  OAI21_X1 U15031 ( .B1(n13379), .B2(n13836), .A(n13378), .ZN(P3_U3473) );
  INV_X1 U15032 ( .A(n13837), .ZN(n13401) );
  NAND2_X1 U15033 ( .A1(n13380), .A2(n13401), .ZN(n13382) );
  NAND2_X1 U15034 ( .A1(n13381), .A2(n16602), .ZN(n13385) );
  OAI211_X1 U15035 ( .C1(n16602), .C2(n13383), .A(n13382), .B(n13385), .ZN(
        P3_U3458) );
  NAND2_X1 U15036 ( .A1(n13384), .A2(n13401), .ZN(n13386) );
  OAI211_X1 U15037 ( .C1(n16602), .C2(n13387), .A(n13386), .B(n13385), .ZN(
        P3_U3457) );
  MUX2_X1 U15038 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n13391), .S(n16602), .Z(
        P3_U3454) );
  MUX2_X1 U15039 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n13392), .S(n16602), .Z(
        P3_U3453) );
  MUX2_X1 U15040 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n13393), .S(n16602), .Z(
        P3_U3452) );
  MUX2_X1 U15041 ( .A(n13395), .B(n13394), .S(n16605), .Z(n13396) );
  OAI21_X1 U15042 ( .B1(n13397), .B2(n13837), .A(n13396), .ZN(P3_U3451) );
  MUX2_X1 U15043 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n13398), .S(n16602), .Z(
        n13399) );
  AOI21_X1 U15044 ( .B1(n13401), .B2(n13400), .A(n13399), .ZN(n13402) );
  INV_X1 U15045 ( .A(n13402), .ZN(P3_U3450) );
  INV_X1 U15046 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13404) );
  MUX2_X1 U15047 ( .A(n13404), .B(n13403), .S(n16602), .Z(n13405) );
  OAI21_X1 U15048 ( .B1(n13406), .B2(n13837), .A(n13405), .ZN(P3_U3449) );
  XNOR2_X1 U15049 ( .A(P3_WR_REG_SCAN_IN), .B(keyinput_128), .ZN(n13409) );
  XNOR2_X1 U15050 ( .A(SI_31_), .B(keyinput_129), .ZN(n13408) );
  XNOR2_X1 U15051 ( .A(SI_30_), .B(keyinput_130), .ZN(n13407) );
  OAI21_X1 U15052 ( .B1(n13409), .B2(n13408), .A(n13407), .ZN(n13414) );
  XNOR2_X1 U15053 ( .A(n13410), .B(keyinput_132), .ZN(n13413) );
  XOR2_X1 U15054 ( .A(SI_27_), .B(keyinput_133), .Z(n13412) );
  XNOR2_X1 U15055 ( .A(n13851), .B(keyinput_131), .ZN(n13411) );
  NAND4_X1 U15056 ( .A1(n13414), .A2(n13413), .A3(n13412), .A4(n13411), .ZN(
        n13417) );
  XNOR2_X1 U15057 ( .A(SI_26_), .B(keyinput_134), .ZN(n13416) );
  XNOR2_X1 U15058 ( .A(n13610), .B(keyinput_135), .ZN(n13415) );
  AOI21_X1 U15059 ( .B1(n13417), .B2(n13416), .A(n13415), .ZN(n13420) );
  XOR2_X1 U15060 ( .A(SI_24_), .B(keyinput_136), .Z(n13419) );
  XNOR2_X1 U15061 ( .A(n13614), .B(keyinput_137), .ZN(n13418) );
  OAI21_X1 U15062 ( .B1(n13420), .B2(n13419), .A(n13418), .ZN(n13424) );
  XOR2_X1 U15063 ( .A(SI_22_), .B(keyinput_138), .Z(n13423) );
  XNOR2_X1 U15064 ( .A(SI_20_), .B(keyinput_140), .ZN(n13422) );
  XNOR2_X1 U15065 ( .A(SI_21_), .B(keyinput_139), .ZN(n13421) );
  NAND4_X1 U15066 ( .A1(n13424), .A2(n13423), .A3(n13422), .A4(n13421), .ZN(
        n13427) );
  XNOR2_X1 U15067 ( .A(SI_19_), .B(keyinput_141), .ZN(n13426) );
  XOR2_X1 U15068 ( .A(SI_18_), .B(keyinput_142), .Z(n13425) );
  AOI21_X1 U15069 ( .B1(n13427), .B2(n13426), .A(n13425), .ZN(n13432) );
  XNOR2_X1 U15070 ( .A(SI_17_), .B(keyinput_143), .ZN(n13431) );
  XNOR2_X1 U15071 ( .A(n13428), .B(keyinput_145), .ZN(n13430) );
  XNOR2_X1 U15072 ( .A(SI_16_), .B(keyinput_144), .ZN(n13429) );
  OAI211_X1 U15073 ( .C1(n13432), .C2(n13431), .A(n13430), .B(n13429), .ZN(
        n13435) );
  XNOR2_X1 U15074 ( .A(n13629), .B(keyinput_147), .ZN(n13434) );
  XNOR2_X1 U15075 ( .A(SI_14_), .B(keyinput_146), .ZN(n13433) );
  NAND3_X1 U15076 ( .A1(n13435), .A2(n13434), .A3(n13433), .ZN(n13447) );
  XNOR2_X1 U15077 ( .A(n13436), .B(keyinput_148), .ZN(n13446) );
  XOR2_X1 U15078 ( .A(SI_9_), .B(keyinput_151), .Z(n13441) );
  XNOR2_X1 U15079 ( .A(n13437), .B(keyinput_149), .ZN(n13440) );
  XNOR2_X1 U15080 ( .A(SI_7_), .B(keyinput_153), .ZN(n13439) );
  XNOR2_X1 U15081 ( .A(SI_6_), .B(keyinput_154), .ZN(n13438) );
  NOR4_X1 U15082 ( .A1(n13441), .A2(n13440), .A3(n13439), .A4(n13438), .ZN(
        n13444) );
  XOR2_X1 U15083 ( .A(SI_10_), .B(keyinput_150), .Z(n13443) );
  XOR2_X1 U15084 ( .A(SI_8_), .B(keyinput_152), .Z(n13442) );
  NAND3_X1 U15085 ( .A1(n13444), .A2(n13443), .A3(n13442), .ZN(n13445) );
  AOI21_X1 U15086 ( .B1(n13447), .B2(n13446), .A(n13445), .ZN(n13450) );
  XOR2_X1 U15087 ( .A(SI_5_), .B(keyinput_155), .Z(n13449) );
  XNOR2_X1 U15088 ( .A(SI_4_), .B(keyinput_156), .ZN(n13448) );
  NOR3_X1 U15089 ( .A1(n13450), .A2(n13449), .A3(n13448), .ZN(n13453) );
  XOR2_X1 U15090 ( .A(SI_3_), .B(keyinput_157), .Z(n13452) );
  XNOR2_X1 U15091 ( .A(SI_2_), .B(keyinput_158), .ZN(n13451) );
  NOR3_X1 U15092 ( .A1(n13453), .A2(n13452), .A3(n13451), .ZN(n13459) );
  XNOR2_X1 U15093 ( .A(n13650), .B(keyinput_159), .ZN(n13458) );
  XOR2_X1 U15094 ( .A(SI_0_), .B(keyinput_160), .Z(n13456) );
  XNOR2_X1 U15095 ( .A(P3_U3151), .B(keyinput_162), .ZN(n13455) );
  XNOR2_X1 U15096 ( .A(P3_RD_REG_SCAN_IN), .B(keyinput_161), .ZN(n13454) );
  NOR3_X1 U15097 ( .A1(n13456), .A2(n13455), .A3(n13454), .ZN(n13457) );
  OAI21_X1 U15098 ( .B1(n13459), .B2(n13458), .A(n13457), .ZN(n13465) );
  XNOR2_X1 U15099 ( .A(n13460), .B(keyinput_163), .ZN(n13464) );
  XOR2_X1 U15100 ( .A(P3_REG3_REG_14__SCAN_IN), .B(keyinput_165), .Z(n13463)
         );
  XNOR2_X1 U15101 ( .A(n13461), .B(keyinput_164), .ZN(n13462) );
  AOI211_X1 U15102 ( .C1(n13465), .C2(n13464), .A(n13463), .B(n13462), .ZN(
        n13468) );
  XOR2_X1 U15103 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_166), .Z(n13467)
         );
  XNOR2_X1 U15104 ( .A(P3_REG3_REG_10__SCAN_IN), .B(keyinput_167), .ZN(n13466)
         );
  OAI21_X1 U15105 ( .B1(n13468), .B2(n13467), .A(n13466), .ZN(n13482) );
  XNOR2_X1 U15106 ( .A(n13666), .B(keyinput_173), .ZN(n13474) );
  XOR2_X1 U15107 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput_170), .Z(n13473)
         );
  XNOR2_X1 U15108 ( .A(n13469), .B(keyinput_169), .ZN(n13472) );
  XOR2_X1 U15109 ( .A(n13470), .B(keyinput_171), .Z(n13471) );
  NAND4_X1 U15110 ( .A1(n13474), .A2(n13473), .A3(n13472), .A4(n13471), .ZN(
        n13479) );
  XOR2_X1 U15111 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_172), .Z(n13478) );
  XNOR2_X1 U15112 ( .A(n13475), .B(keyinput_168), .ZN(n13477) );
  XNOR2_X1 U15113 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput_174), .ZN(n13476)
         );
  NOR4_X1 U15114 ( .A1(n13479), .A2(n13478), .A3(n13477), .A4(n13476), .ZN(
        n13481) );
  XNOR2_X1 U15115 ( .A(P3_REG3_REG_25__SCAN_IN), .B(keyinput_175), .ZN(n13480)
         );
  AOI21_X1 U15116 ( .B1(n13482), .B2(n13481), .A(n13480), .ZN(n13485) );
  XOR2_X1 U15117 ( .A(P3_REG3_REG_16__SCAN_IN), .B(keyinput_176), .Z(n13484)
         );
  XNOR2_X1 U15118 ( .A(n13679), .B(keyinput_177), .ZN(n13483) );
  OAI21_X1 U15119 ( .B1(n13485), .B2(n13484), .A(n13483), .ZN(n13488) );
  XNOR2_X1 U15120 ( .A(n13680), .B(keyinput_178), .ZN(n13487) );
  XNOR2_X1 U15121 ( .A(P3_REG3_REG_24__SCAN_IN), .B(keyinput_179), .ZN(n13486)
         );
  AOI21_X1 U15122 ( .B1(n13488), .B2(n13487), .A(n13486), .ZN(n13492) );
  XNOR2_X1 U15123 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput_180), .ZN(n13491)
         );
  XNOR2_X1 U15124 ( .A(n13489), .B(keyinput_181), .ZN(n13490) );
  OAI21_X1 U15125 ( .B1(n13492), .B2(n13491), .A(n13490), .ZN(n13498) );
  XNOR2_X1 U15126 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_182), .ZN(n13497)
         );
  XOR2_X1 U15127 ( .A(P3_REG3_REG_20__SCAN_IN), .B(keyinput_183), .Z(n13495)
         );
  XNOR2_X1 U15128 ( .A(P3_REG3_REG_22__SCAN_IN), .B(keyinput_185), .ZN(n13494)
         );
  XNOR2_X1 U15129 ( .A(P3_REG3_REG_13__SCAN_IN), .B(keyinput_184), .ZN(n13493)
         );
  NAND3_X1 U15130 ( .A1(n13495), .A2(n13494), .A3(n13493), .ZN(n13496) );
  AOI21_X1 U15131 ( .B1(n13498), .B2(n13497), .A(n13496), .ZN(n13501) );
  XOR2_X1 U15132 ( .A(P3_REG3_REG_11__SCAN_IN), .B(keyinput_186), .Z(n13500)
         );
  XOR2_X1 U15133 ( .A(P3_REG3_REG_2__SCAN_IN), .B(keyinput_187), .Z(n13499) );
  OAI21_X1 U15134 ( .B1(n13501), .B2(n13500), .A(n13499), .ZN(n13505) );
  XNOR2_X1 U15135 ( .A(P3_REG3_REG_18__SCAN_IN), .B(keyinput_188), .ZN(n13504)
         );
  XOR2_X1 U15136 ( .A(P3_REG3_REG_26__SCAN_IN), .B(keyinput_190), .Z(n13503)
         );
  XNOR2_X1 U15137 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_189), .ZN(n13502)
         );
  AOI211_X1 U15138 ( .C1(n13505), .C2(n13504), .A(n13503), .B(n13502), .ZN(
        n13510) );
  XNOR2_X1 U15139 ( .A(P3_REG3_REG_15__SCAN_IN), .B(keyinput_191), .ZN(n13509)
         );
  XNOR2_X1 U15140 ( .A(n13506), .B(keyinput_192), .ZN(n13508) );
  XNOR2_X1 U15141 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(keyinput_193), .ZN(n13507) );
  OAI211_X1 U15142 ( .C1(n13510), .C2(n13509), .A(n13508), .B(n13507), .ZN(
        n13513) );
  XNOR2_X1 U15143 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(keyinput_194), .ZN(n13512) );
  XOR2_X1 U15144 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(keyinput_195), .Z(n13511)
         );
  AOI21_X1 U15145 ( .B1(n13513), .B2(n13512), .A(n13511), .ZN(n13516) );
  XNOR2_X1 U15146 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .ZN(n13515) );
  XNOR2_X1 U15147 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(keyinput_197), .ZN(n13514) );
  OAI21_X1 U15148 ( .B1(n13516), .B2(n13515), .A(n13514), .ZN(n13519) );
  XNOR2_X1 U15149 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(keyinput_199), .ZN(n13518) );
  XNOR2_X1 U15150 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(keyinput_198), .ZN(n13517) );
  NAND3_X1 U15151 ( .A1(n13519), .A2(n13518), .A3(n13517), .ZN(n13523) );
  XOR2_X1 U15152 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(keyinput_200), .Z(n13522)
         );
  XOR2_X1 U15153 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(keyinput_201), .Z(n13521)
         );
  XNOR2_X1 U15154 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(keyinput_202), .ZN(n13520) );
  AOI211_X1 U15155 ( .C1(n13523), .C2(n13522), .A(n13521), .B(n13520), .ZN(
        n13526) );
  XOR2_X1 U15156 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(keyinput_204), .Z(n13525)
         );
  XNOR2_X1 U15157 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(keyinput_203), .ZN(n13524) );
  NOR3_X1 U15158 ( .A1(n13526), .A2(n13525), .A3(n13524), .ZN(n13529) );
  XOR2_X1 U15159 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(keyinput_205), .Z(n13528)
         );
  XNOR2_X1 U15160 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .ZN(n13527) );
  NOR3_X1 U15161 ( .A1(n13529), .A2(n13528), .A3(n13527), .ZN(n13535) );
  XNOR2_X1 U15162 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(keyinput_207), .ZN(n13534) );
  XOR2_X1 U15163 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(keyinput_208), .Z(n13532)
         );
  XNOR2_X1 U15164 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(keyinput_210), .ZN(n13531) );
  XNOR2_X1 U15165 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(keyinput_209), .ZN(n13530) );
  NOR3_X1 U15166 ( .A1(n13532), .A2(n13531), .A3(n13530), .ZN(n13533) );
  OAI21_X1 U15167 ( .B1(n13535), .B2(n13534), .A(n13533), .ZN(n13539) );
  XOR2_X1 U15168 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(keyinput_213), .Z(n13538)
         );
  XOR2_X1 U15169 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(keyinput_212), .Z(n13537)
         );
  XNOR2_X1 U15170 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(keyinput_211), .ZN(n13536) );
  NAND4_X1 U15171 ( .A1(n13539), .A2(n13538), .A3(n13537), .A4(n13536), .ZN(
        n13542) );
  XOR2_X1 U15172 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(keyinput_215), .Z(n13541)
         );
  XOR2_X1 U15173 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .Z(n13540)
         );
  NAND3_X1 U15174 ( .A1(n13542), .A2(n13541), .A3(n13540), .ZN(n13545) );
  XOR2_X1 U15175 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(keyinput_216), .Z(n13544)
         );
  XNOR2_X1 U15176 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(keyinput_217), .ZN(n13543)
         );
  NAND3_X1 U15177 ( .A1(n13545), .A2(n13544), .A3(n13543), .ZN(n13548) );
  XOR2_X1 U15178 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(keyinput_218), .Z(n13547)
         );
  XOR2_X1 U15179 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(keyinput_219), .Z(n13546)
         );
  NAND3_X1 U15180 ( .A1(n13548), .A2(n13547), .A3(n13546), .ZN(n13552) );
  XOR2_X1 U15181 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(keyinput_222), .Z(n13551)
         );
  XNOR2_X1 U15182 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(keyinput_221), .ZN(n13550)
         );
  XNOR2_X1 U15183 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(keyinput_220), .ZN(n13549)
         );
  NAND4_X1 U15184 ( .A1(n13552), .A2(n13551), .A3(n13550), .A4(n13549), .ZN(
        n13555) );
  XNOR2_X1 U15185 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(keyinput_224), .ZN(n13554)
         );
  XNOR2_X1 U15186 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(keyinput_223), .ZN(n13553)
         );
  NAND3_X1 U15187 ( .A1(n13555), .A2(n13554), .A3(n13553), .ZN(n13558) );
  XOR2_X1 U15188 ( .A(P3_ADDR_REG_0__SCAN_IN), .B(keyinput_225), .Z(n13557) );
  XOR2_X1 U15189 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(keyinput_226), .Z(n13556) );
  AOI21_X1 U15190 ( .B1(n13558), .B2(n13557), .A(n13556), .ZN(n13561) );
  XNOR2_X1 U15191 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(keyinput_227), .ZN(n13560)
         );
  XNOR2_X1 U15192 ( .A(P3_ADDR_REG_3__SCAN_IN), .B(keyinput_228), .ZN(n13559)
         );
  OAI21_X1 U15193 ( .B1(n13561), .B2(n13560), .A(n13559), .ZN(n13564) );
  XNOR2_X1 U15194 ( .A(P3_ADDR_REG_4__SCAN_IN), .B(keyinput_229), .ZN(n13563)
         );
  XOR2_X1 U15195 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(keyinput_230), .Z(n13562) );
  AOI21_X1 U15196 ( .B1(n13564), .B2(n13563), .A(n13562), .ZN(n13567) );
  XOR2_X1 U15197 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(keyinput_231), .Z(n13566) );
  XNOR2_X1 U15198 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(keyinput_232), .ZN(n13565)
         );
  OAI21_X1 U15199 ( .B1(n13567), .B2(n13566), .A(n13565), .ZN(n13570) );
  XOR2_X1 U15200 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(keyinput_233), .Z(n13569) );
  XNOR2_X1 U15201 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(keyinput_234), .ZN(n13568)
         );
  NAND3_X1 U15202 ( .A1(n13570), .A2(n13569), .A3(n13568), .ZN(n13573) );
  XNOR2_X1 U15203 ( .A(n15887), .B(keyinput_235), .ZN(n13572) );
  XOR2_X1 U15204 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_236), .Z(n13571) );
  AOI21_X1 U15205 ( .B1(n13573), .B2(n13572), .A(n13571), .ZN(n13577) );
  XNOR2_X1 U15206 ( .A(n13770), .B(keyinput_237), .ZN(n13576) );
  XOR2_X1 U15207 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_239), .Z(n13575) );
  XNOR2_X1 U15208 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_238), .ZN(n13574) );
  NOR4_X1 U15209 ( .A1(n13577), .A2(n13576), .A3(n13575), .A4(n13574), .ZN(
        n13580) );
  XNOR2_X1 U15210 ( .A(n13775), .B(keyinput_240), .ZN(n13579) );
  XNOR2_X1 U15211 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_241), .ZN(n13578) );
  OAI21_X1 U15212 ( .B1(n13580), .B2(n13579), .A(n13578), .ZN(n13595) );
  XNOR2_X1 U15213 ( .A(n13581), .B(keyinput_243), .ZN(n13588) );
  XNOR2_X1 U15214 ( .A(n13582), .B(keyinput_242), .ZN(n13587) );
  XNOR2_X1 U15215 ( .A(n13583), .B(keyinput_244), .ZN(n13586) );
  XNOR2_X1 U15216 ( .A(n13584), .B(keyinput_245), .ZN(n13585) );
  NOR4_X1 U15217 ( .A1(n13588), .A2(n13587), .A3(n13586), .A4(n13585), .ZN(
        n13594) );
  XNOR2_X1 U15218 ( .A(n13589), .B(keyinput_246), .ZN(n13592) );
  XNOR2_X1 U15219 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_247), .ZN(n13591)
         );
  XNOR2_X1 U15220 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_248), .ZN(n13590)
         );
  NAND3_X1 U15221 ( .A1(n13592), .A2(n13591), .A3(n13590), .ZN(n13593) );
  AOI21_X1 U15222 ( .B1(n13595), .B2(n13594), .A(n13593), .ZN(n13599) );
  XNOR2_X1 U15223 ( .A(n13789), .B(keyinput_250), .ZN(n13598) );
  XOR2_X1 U15224 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_249), .Z(n13597) );
  XNOR2_X1 U15225 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_251), .ZN(n13596)
         );
  NOR4_X1 U15226 ( .A1(n13599), .A2(n13598), .A3(n13597), .A4(n13596), .ZN(
        n13602) );
  XOR2_X1 U15227 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_253), .Z(n13601) );
  XNOR2_X1 U15228 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_252), .ZN(n13600)
         );
  NOR3_X1 U15229 ( .A1(n13602), .A2(n13601), .A3(n13600), .ZN(n13805) );
  XNOR2_X1 U15230 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_254), .ZN(n13804)
         );
  XOR2_X1 U15231 ( .A(SI_31_), .B(keyinput_1), .Z(n13605) );
  XOR2_X1 U15232 ( .A(P3_WR_REG_SCAN_IN), .B(keyinput_0), .Z(n13604) );
  XOR2_X1 U15233 ( .A(SI_30_), .B(keyinput_2), .Z(n13603) );
  AOI21_X1 U15234 ( .B1(n13605), .B2(n13604), .A(n13603), .ZN(n13609) );
  XOR2_X1 U15235 ( .A(SI_27_), .B(keyinput_5), .Z(n13608) );
  XNOR2_X1 U15236 ( .A(SI_28_), .B(keyinput_4), .ZN(n13607) );
  XNOR2_X1 U15237 ( .A(SI_29_), .B(keyinput_3), .ZN(n13606) );
  NOR4_X1 U15238 ( .A1(n13609), .A2(n13608), .A3(n13607), .A4(n13606), .ZN(
        n13613) );
  XOR2_X1 U15239 ( .A(SI_26_), .B(keyinput_6), .Z(n13612) );
  XNOR2_X1 U15240 ( .A(n13610), .B(keyinput_7), .ZN(n13611) );
  OAI21_X1 U15241 ( .B1(n13613), .B2(n13612), .A(n13611), .ZN(n13617) );
  XNOR2_X1 U15242 ( .A(SI_24_), .B(keyinput_8), .ZN(n13616) );
  XNOR2_X1 U15243 ( .A(n13614), .B(keyinput_9), .ZN(n13615) );
  AOI21_X1 U15244 ( .B1(n13617), .B2(n13616), .A(n13615), .ZN(n13621) );
  XOR2_X1 U15245 ( .A(SI_21_), .B(keyinput_11), .Z(n13620) );
  XOR2_X1 U15246 ( .A(SI_20_), .B(keyinput_12), .Z(n13619) );
  XNOR2_X1 U15247 ( .A(SI_22_), .B(keyinput_10), .ZN(n13618) );
  NOR4_X1 U15248 ( .A1(n13621), .A2(n13620), .A3(n13619), .A4(n13618), .ZN(
        n13624) );
  XNOR2_X1 U15249 ( .A(SI_19_), .B(keyinput_13), .ZN(n13623) );
  XOR2_X1 U15250 ( .A(SI_18_), .B(keyinput_14), .Z(n13622) );
  OAI21_X1 U15251 ( .B1(n13624), .B2(n13623), .A(n13622), .ZN(n13628) );
  XNOR2_X1 U15252 ( .A(SI_17_), .B(keyinput_15), .ZN(n13627) );
  XNOR2_X1 U15253 ( .A(SI_15_), .B(keyinput_17), .ZN(n13626) );
  XNOR2_X1 U15254 ( .A(SI_16_), .B(keyinput_16), .ZN(n13625) );
  AOI211_X1 U15255 ( .C1(n13628), .C2(n13627), .A(n13626), .B(n13625), .ZN(
        n13632) );
  XNOR2_X1 U15256 ( .A(n13629), .B(keyinput_19), .ZN(n13631) );
  XNOR2_X1 U15257 ( .A(SI_14_), .B(keyinput_18), .ZN(n13630) );
  NOR3_X1 U15258 ( .A1(n13632), .A2(n13631), .A3(n13630), .ZN(n13643) );
  XNOR2_X1 U15259 ( .A(SI_12_), .B(keyinput_20), .ZN(n13642) );
  XOR2_X1 U15260 ( .A(SI_6_), .B(keyinput_26), .Z(n13634) );
  XOR2_X1 U15261 ( .A(SI_7_), .B(keyinput_25), .Z(n13633) );
  NAND2_X1 U15262 ( .A1(n13634), .A2(n13633), .ZN(n13640) );
  XNOR2_X1 U15263 ( .A(SI_10_), .B(keyinput_22), .ZN(n13636) );
  XNOR2_X1 U15264 ( .A(SI_11_), .B(keyinput_21), .ZN(n13635) );
  NAND2_X1 U15265 ( .A1(n13636), .A2(n13635), .ZN(n13639) );
  XNOR2_X1 U15266 ( .A(SI_8_), .B(keyinput_24), .ZN(n13638) );
  XNOR2_X1 U15267 ( .A(SI_9_), .B(keyinput_23), .ZN(n13637) );
  NOR4_X1 U15268 ( .A1(n13640), .A2(n13639), .A3(n13638), .A4(n13637), .ZN(
        n13641) );
  OAI21_X1 U15269 ( .B1(n13643), .B2(n13642), .A(n13641), .ZN(n13646) );
  XOR2_X1 U15270 ( .A(SI_5_), .B(keyinput_27), .Z(n13645) );
  XOR2_X1 U15271 ( .A(SI_4_), .B(keyinput_28), .Z(n13644) );
  NAND3_X1 U15272 ( .A1(n13646), .A2(n13645), .A3(n13644), .ZN(n13649) );
  XOR2_X1 U15273 ( .A(SI_3_), .B(keyinput_29), .Z(n13648) );
  XNOR2_X1 U15274 ( .A(SI_2_), .B(keyinput_30), .ZN(n13647) );
  NAND3_X1 U15275 ( .A1(n13649), .A2(n13648), .A3(n13647), .ZN(n13656) );
  XNOR2_X1 U15276 ( .A(n13650), .B(keyinput_31), .ZN(n13655) );
  XNOR2_X1 U15277 ( .A(P3_U3151), .B(keyinput_34), .ZN(n13653) );
  XNOR2_X1 U15278 ( .A(P3_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n13652) );
  XNOR2_X1 U15279 ( .A(SI_0_), .B(keyinput_32), .ZN(n13651) );
  NAND3_X1 U15280 ( .A1(n13653), .A2(n13652), .A3(n13651), .ZN(n13654) );
  AOI21_X1 U15281 ( .B1(n13656), .B2(n13655), .A(n13654), .ZN(n13660) );
  XNOR2_X1 U15282 ( .A(P3_REG3_REG_7__SCAN_IN), .B(keyinput_35), .ZN(n13659)
         );
  XNOR2_X1 U15283 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput_36), .ZN(n13658)
         );
  XNOR2_X1 U15284 ( .A(P3_REG3_REG_14__SCAN_IN), .B(keyinput_37), .ZN(n13657)
         );
  OAI211_X1 U15285 ( .C1(n13660), .C2(n13659), .A(n13658), .B(n13657), .ZN(
        n13663) );
  XOR2_X1 U15286 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_38), .Z(n13662) );
  XOR2_X1 U15287 ( .A(P3_REG3_REG_10__SCAN_IN), .B(keyinput_39), .Z(n13661) );
  AOI21_X1 U15288 ( .B1(n13663), .B2(n13662), .A(n13661), .ZN(n13674) );
  XNOR2_X1 U15289 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput_46), .ZN(n13673)
         );
  XNOR2_X1 U15290 ( .A(P3_REG3_REG_19__SCAN_IN), .B(keyinput_41), .ZN(n13665)
         );
  XNOR2_X1 U15291 ( .A(P3_REG3_REG_3__SCAN_IN), .B(keyinput_40), .ZN(n13664)
         );
  NAND2_X1 U15292 ( .A1(n13665), .A2(n13664), .ZN(n13672) );
  XOR2_X1 U15293 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput_42), .Z(n13670) );
  XOR2_X1 U15294 ( .A(P3_REG3_REG_8__SCAN_IN), .B(keyinput_43), .Z(n13669) );
  XNOR2_X1 U15295 ( .A(n13666), .B(keyinput_45), .ZN(n13668) );
  XNOR2_X1 U15296 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_44), .ZN(n13667)
         );
  NAND4_X1 U15297 ( .A1(n13670), .A2(n13669), .A3(n13668), .A4(n13667), .ZN(
        n13671) );
  NOR4_X1 U15298 ( .A1(n13674), .A2(n13673), .A3(n13672), .A4(n13671), .ZN(
        n13678) );
  XNOR2_X1 U15299 ( .A(n13675), .B(keyinput_47), .ZN(n13677) );
  XNOR2_X1 U15300 ( .A(P3_REG3_REG_16__SCAN_IN), .B(keyinput_48), .ZN(n13676)
         );
  OAI21_X1 U15301 ( .B1(n13678), .B2(n13677), .A(n13676), .ZN(n13683) );
  XNOR2_X1 U15302 ( .A(n13679), .B(keyinput_49), .ZN(n13682) );
  XNOR2_X1 U15303 ( .A(n13680), .B(keyinput_50), .ZN(n13681) );
  AOI21_X1 U15304 ( .B1(n13683), .B2(n13682), .A(n13681), .ZN(n13686) );
  XNOR2_X1 U15305 ( .A(P3_REG3_REG_24__SCAN_IN), .B(keyinput_51), .ZN(n13685)
         );
  XNOR2_X1 U15306 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput_52), .ZN(n13684)
         );
  OAI21_X1 U15307 ( .B1(n13686), .B2(n13685), .A(n13684), .ZN(n13689) );
  XNOR2_X1 U15308 ( .A(P3_REG3_REG_9__SCAN_IN), .B(keyinput_53), .ZN(n13688)
         );
  XNOR2_X1 U15309 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_54), .ZN(n13687)
         );
  AOI21_X1 U15310 ( .B1(n13689), .B2(n13688), .A(n13687), .ZN(n13694) );
  XOR2_X1 U15311 ( .A(P3_REG3_REG_22__SCAN_IN), .B(keyinput_57), .Z(n13693) );
  XOR2_X1 U15312 ( .A(P3_REG3_REG_20__SCAN_IN), .B(keyinput_55), .Z(n13692) );
  XNOR2_X1 U15313 ( .A(n13690), .B(keyinput_56), .ZN(n13691) );
  NOR4_X1 U15314 ( .A1(n13694), .A2(n13693), .A3(n13692), .A4(n13691), .ZN(
        n13697) );
  XNOR2_X1 U15315 ( .A(P3_REG3_REG_11__SCAN_IN), .B(keyinput_58), .ZN(n13696)
         );
  XNOR2_X1 U15316 ( .A(P3_REG3_REG_2__SCAN_IN), .B(keyinput_59), .ZN(n13695)
         );
  OAI21_X1 U15317 ( .B1(n13697), .B2(n13696), .A(n13695), .ZN(n13701) );
  XNOR2_X1 U15318 ( .A(P3_REG3_REG_18__SCAN_IN), .B(keyinput_60), .ZN(n13700)
         );
  XNOR2_X1 U15319 ( .A(P3_REG3_REG_26__SCAN_IN), .B(keyinput_62), .ZN(n13699)
         );
  XNOR2_X1 U15320 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_61), .ZN(n13698)
         );
  AOI211_X1 U15321 ( .C1(n13701), .C2(n13700), .A(n13699), .B(n13698), .ZN(
        n13706) );
  XNOR2_X1 U15322 ( .A(n13702), .B(keyinput_63), .ZN(n13705) );
  XOR2_X1 U15323 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .Z(n13704)
         );
  XNOR2_X1 U15324 ( .A(P3_B_REG_SCAN_IN), .B(keyinput_64), .ZN(n13703) );
  OAI211_X1 U15325 ( .C1(n13706), .C2(n13705), .A(n13704), .B(n13703), .ZN(
        n13709) );
  XNOR2_X1 U15326 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(keyinput_66), .ZN(n13708)
         );
  XOR2_X1 U15327 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .Z(n13707)
         );
  AOI21_X1 U15328 ( .B1(n13709), .B2(n13708), .A(n13707), .ZN(n13712) );
  XOR2_X1 U15329 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .Z(n13711)
         );
  XOR2_X1 U15330 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(keyinput_69), .Z(n13710)
         );
  OAI21_X1 U15331 ( .B1(n13712), .B2(n13711), .A(n13710), .ZN(n13715) );
  XNOR2_X1 U15332 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .ZN(n13714)
         );
  XNOR2_X1 U15333 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(keyinput_70), .ZN(n13713)
         );
  NAND3_X1 U15334 ( .A1(n13715), .A2(n13714), .A3(n13713), .ZN(n13719) );
  XOR2_X1 U15335 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .Z(n13718)
         );
  XOR2_X1 U15336 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .Z(n13717)
         );
  XNOR2_X1 U15337 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .ZN(n13716)
         );
  AOI211_X1 U15338 ( .C1(n13719), .C2(n13718), .A(n13717), .B(n13716), .ZN(
        n13725) );
  XOR2_X1 U15339 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .Z(n13721)
         );
  XNOR2_X1 U15340 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .ZN(n13720)
         );
  NAND2_X1 U15341 ( .A1(n13721), .A2(n13720), .ZN(n13724) );
  XOR2_X1 U15342 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .Z(n13723)
         );
  XNOR2_X1 U15343 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .ZN(n13722)
         );
  OAI211_X1 U15344 ( .C1(n13725), .C2(n13724), .A(n13723), .B(n13722), .ZN(
        n13731) );
  XOR2_X1 U15345 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .Z(n13730)
         );
  XOR2_X1 U15346 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .Z(n13728)
         );
  XOR2_X1 U15347 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(keyinput_80), .Z(n13727)
         );
  XNOR2_X1 U15348 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(keyinput_82), .ZN(n13726)
         );
  NAND3_X1 U15349 ( .A1(n13728), .A2(n13727), .A3(n13726), .ZN(n13729) );
  AOI21_X1 U15350 ( .B1(n13731), .B2(n13730), .A(n13729), .ZN(n13735) );
  XOR2_X1 U15351 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .Z(n13734)
         );
  XOR2_X1 U15352 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .Z(n13733)
         );
  XNOR2_X1 U15353 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(keyinput_84), .ZN(n13732)
         );
  NOR4_X1 U15354 ( .A1(n13735), .A2(n13734), .A3(n13733), .A4(n13732), .ZN(
        n13738) );
  XOR2_X1 U15355 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(keyinput_87), .Z(n13737) );
  XNOR2_X1 U15356 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .ZN(n13736)
         );
  NOR3_X1 U15357 ( .A1(n13738), .A2(n13737), .A3(n13736), .ZN(n13741) );
  XOR2_X1 U15358 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .Z(n13740) );
  XOR2_X1 U15359 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .Z(n13739) );
  NOR3_X1 U15360 ( .A1(n13741), .A2(n13740), .A3(n13739), .ZN(n13744) );
  XOR2_X1 U15361 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(keyinput_90), .Z(n13743) );
  XNOR2_X1 U15362 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(keyinput_91), .ZN(n13742)
         );
  NOR3_X1 U15363 ( .A1(n13744), .A2(n13743), .A3(n13742), .ZN(n13748) );
  XOR2_X1 U15364 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(keyinput_94), .Z(n13747) );
  XOR2_X1 U15365 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(keyinput_92), .Z(n13746) );
  XNOR2_X1 U15366 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(keyinput_93), .ZN(n13745)
         );
  NOR4_X1 U15367 ( .A1(n13748), .A2(n13747), .A3(n13746), .A4(n13745), .ZN(
        n13751) );
  XNOR2_X1 U15368 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(keyinput_96), .ZN(n13750)
         );
  XNOR2_X1 U15369 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(keyinput_95), .ZN(n13749)
         );
  NOR3_X1 U15370 ( .A1(n13751), .A2(n13750), .A3(n13749), .ZN(n13754) );
  XOR2_X1 U15371 ( .A(P3_ADDR_REG_0__SCAN_IN), .B(keyinput_97), .Z(n13753) );
  XNOR2_X1 U15372 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(keyinput_98), .ZN(n13752)
         );
  OAI21_X1 U15373 ( .B1(n13754), .B2(n13753), .A(n13752), .ZN(n13757) );
  XOR2_X1 U15374 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(keyinput_99), .Z(n13756) );
  XOR2_X1 U15375 ( .A(P3_ADDR_REG_3__SCAN_IN), .B(keyinput_100), .Z(n13755) );
  AOI21_X1 U15376 ( .B1(n13757), .B2(n13756), .A(n13755), .ZN(n13760) );
  XOR2_X1 U15377 ( .A(P3_ADDR_REG_4__SCAN_IN), .B(keyinput_101), .Z(n13759) );
  XOR2_X1 U15378 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(keyinput_102), .Z(n13758) );
  OAI21_X1 U15379 ( .B1(n13760), .B2(n13759), .A(n13758), .ZN(n13763) );
  XOR2_X1 U15380 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(keyinput_103), .Z(n13762) );
  XOR2_X1 U15381 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(keyinput_104), .Z(n13761) );
  AOI21_X1 U15382 ( .B1(n13763), .B2(n13762), .A(n13761), .ZN(n13766) );
  XNOR2_X1 U15383 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(keyinput_106), .ZN(n13765)
         );
  XNOR2_X1 U15384 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(keyinput_105), .ZN(n13764)
         );
  NOR3_X1 U15385 ( .A1(n13766), .A2(n13765), .A3(n13764), .ZN(n13769) );
  XNOR2_X1 U15386 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_107), .ZN(n13768) );
  XOR2_X1 U15387 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_108), .Z(n13767) );
  OAI21_X1 U15388 ( .B1(n13769), .B2(n13768), .A(n13767), .ZN(n13774) );
  XOR2_X1 U15389 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_111), .Z(n13773) );
  XOR2_X1 U15390 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_110), .Z(n13772) );
  XNOR2_X1 U15391 ( .A(n13770), .B(keyinput_109), .ZN(n13771) );
  NAND4_X1 U15392 ( .A1(n13774), .A2(n13773), .A3(n13772), .A4(n13771), .ZN(
        n13778) );
  XNOR2_X1 U15393 ( .A(n13775), .B(keyinput_112), .ZN(n13777) );
  XNOR2_X1 U15394 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_113), .ZN(n13776) );
  AOI21_X1 U15395 ( .B1(n13778), .B2(n13777), .A(n13776), .ZN(n13788) );
  XNOR2_X1 U15396 ( .A(n13582), .B(keyinput_114), .ZN(n13782) );
  XNOR2_X1 U15397 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_116), .ZN(n13781) );
  XNOR2_X1 U15398 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_115), .ZN(n13780) );
  XNOR2_X1 U15399 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_117), .ZN(n13779)
         );
  NAND4_X1 U15400 ( .A1(n13782), .A2(n13781), .A3(n13780), .A4(n13779), .ZN(
        n13787) );
  XNOR2_X1 U15401 ( .A(n9441), .B(keyinput_120), .ZN(n13786) );
  OAI22_X1 U15402 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput_118), .B1(
        P1_IR_REG_12__SCAN_IN), .B2(keyinput_119), .ZN(n13784) );
  AND2_X1 U15403 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput_119), .ZN(n13783)
         );
  AOI211_X1 U15404 ( .C1(P1_IR_REG_11__SCAN_IN), .C2(keyinput_118), .A(n13784), 
        .B(n13783), .ZN(n13785) );
  OAI211_X1 U15405 ( .C1(n13788), .C2(n13787), .A(n13786), .B(n13785), .ZN(
        n13797) );
  XOR2_X1 U15406 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_121), .Z(n13792) );
  XNOR2_X1 U15407 ( .A(n13789), .B(keyinput_122), .ZN(n13791) );
  XNOR2_X1 U15408 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_123), .ZN(n13790)
         );
  NOR3_X1 U15409 ( .A1(n13792), .A2(n13791), .A3(n13790), .ZN(n13796) );
  XNOR2_X1 U15410 ( .A(n13793), .B(keyinput_124), .ZN(n13795) );
  XNOR2_X1 U15411 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_125), .ZN(n13794)
         );
  AOI211_X1 U15412 ( .C1(n13797), .C2(n13796), .A(n13795), .B(n13794), .ZN(
        n13800) );
  XOR2_X1 U15413 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_126), .Z(n13799) );
  XOR2_X1 U15414 ( .A(keyinput_255), .B(keyinput_127), .Z(n13798) );
  OAI21_X1 U15415 ( .B1(n13800), .B2(n13799), .A(n13798), .ZN(n13803) );
  XNOR2_X1 U15416 ( .A(n13801), .B(keyinput_255), .ZN(n13802) );
  OAI211_X1 U15417 ( .C1(n13805), .C2(n13804), .A(n13803), .B(n13802), .ZN(
        n13808) );
  MUX2_X1 U15418 ( .A(P3_REG0_REG_21__SCAN_IN), .B(n13806), .S(n16602), .Z(
        n13807) );
  XNOR2_X1 U15419 ( .A(n13808), .B(n13807), .ZN(P3_U3448) );
  MUX2_X1 U15420 ( .A(n13810), .B(n13809), .S(n16602), .Z(n13811) );
  OAI21_X1 U15421 ( .B1(n13812), .B2(n13837), .A(n13811), .ZN(P3_U3447) );
  INV_X1 U15422 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13814) );
  MUX2_X1 U15423 ( .A(n13814), .B(n13813), .S(n16602), .Z(n13815) );
  OAI21_X1 U15424 ( .B1(n13816), .B2(n13837), .A(n13815), .ZN(P3_U3446) );
  INV_X1 U15425 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13818) );
  MUX2_X1 U15426 ( .A(n13818), .B(n13817), .S(n16602), .Z(n13819) );
  OAI21_X1 U15427 ( .B1(n13820), .B2(n13837), .A(n13819), .ZN(P3_U3444) );
  INV_X1 U15428 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13821) );
  MUX2_X1 U15429 ( .A(n13822), .B(n13821), .S(n16605), .Z(n13823) );
  OAI21_X1 U15430 ( .B1(n13837), .B2(n13824), .A(n13823), .ZN(P3_U3441) );
  INV_X1 U15431 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13826) );
  MUX2_X1 U15432 ( .A(n13826), .B(n13825), .S(n16602), .Z(n13827) );
  OAI21_X1 U15433 ( .B1(n13828), .B2(n13837), .A(n13827), .ZN(P3_U3438) );
  INV_X1 U15434 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13830) );
  MUX2_X1 U15435 ( .A(n13830), .B(n13829), .S(n16602), .Z(n13831) );
  OAI21_X1 U15436 ( .B1(n13837), .B2(n13832), .A(n13831), .ZN(P3_U3435) );
  INV_X1 U15437 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13834) );
  MUX2_X1 U15438 ( .A(n13834), .B(n13833), .S(n16602), .Z(n13835) );
  OAI21_X1 U15439 ( .B1(n13837), .B2(n13836), .A(n13835), .ZN(P3_U3432) );
  MUX2_X1 U15440 ( .A(n13839), .B(P3_D_REG_1__SCAN_IN), .S(n13838), .Z(
        P3_U3377) );
  INV_X1 U15441 ( .A(n13840), .ZN(n13848) );
  INV_X1 U15442 ( .A(n13841), .ZN(n13842) );
  NOR4_X1 U15443 ( .A1(n13842), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), 
        .A4(n13843), .ZN(n13845) );
  AOI21_X1 U15444 ( .B1(SI_31_), .B2(n13846), .A(n13845), .ZN(n13847) );
  OAI21_X1 U15445 ( .B1(n13848), .B2(n13853), .A(n13847), .ZN(P3_U3264) );
  INV_X1 U15446 ( .A(n13849), .ZN(n13852) );
  OAI222_X1 U15447 ( .A1(n13854), .A2(P3_U3151), .B1(n13853), .B2(n13852), 
        .C1(n13851), .C2(n13850), .ZN(P3_U3266) );
  MUX2_X1 U15448 ( .A(n13856), .B(n13855), .S(P3_STATE_REG_SCAN_IN), .Z(
        P3_U3294) );
  AND2_X1 U15449 ( .A1(n13858), .A2(n13857), .ZN(n13859) );
  XNOR2_X1 U15450 ( .A(n14671), .B(n10884), .ZN(n13861) );
  XNOR2_X1 U15451 ( .A(n14511), .B(n7433), .ZN(n13934) );
  NAND2_X1 U15452 ( .A1(n14345), .A2(n7437), .ZN(n13863) );
  NOR2_X1 U15453 ( .A1(n13934), .A2(n13863), .ZN(n13864) );
  AOI21_X1 U15454 ( .B1(n13934), .B2(n13863), .A(n13864), .ZN(n13942) );
  INV_X1 U15455 ( .A(n13864), .ZN(n13869) );
  XNOR2_X1 U15456 ( .A(n14497), .B(n10884), .ZN(n13865) );
  AND2_X1 U15457 ( .A1(n14344), .A2(n7437), .ZN(n13866) );
  NAND2_X1 U15458 ( .A1(n13865), .A2(n13866), .ZN(n13870) );
  INV_X1 U15459 ( .A(n13865), .ZN(n13978) );
  INV_X1 U15460 ( .A(n13866), .ZN(n13867) );
  NAND2_X1 U15461 ( .A1(n13978), .A2(n13867), .ZN(n13868) );
  NAND2_X1 U15462 ( .A1(n13870), .A2(n13868), .ZN(n13932) );
  XNOR2_X1 U15463 ( .A(n14482), .B(n7433), .ZN(n13873) );
  NAND2_X1 U15464 ( .A1(n14343), .A2(n7437), .ZN(n13872) );
  XNOR2_X1 U15465 ( .A(n13873), .B(n13872), .ZN(n13980) );
  INV_X1 U15466 ( .A(n13870), .ZN(n13871) );
  NAND2_X1 U15467 ( .A1(n13873), .A2(n13872), .ZN(n13874) );
  XNOR2_X1 U15468 ( .A(n14198), .B(n7433), .ZN(n13908) );
  NAND2_X1 U15469 ( .A1(n14342), .A2(n7437), .ZN(n13875) );
  NOR2_X1 U15470 ( .A1(n13908), .A2(n13875), .ZN(n13916) );
  AOI21_X1 U15471 ( .B1(n13908), .B2(n13875), .A(n13916), .ZN(n13876) );
  OAI211_X1 U15472 ( .C1(n13877), .C2(n13876), .A(n13918), .B(n13990), .ZN(
        n13884) );
  NAND2_X1 U15473 ( .A1(n14341), .A2(n14589), .ZN(n13879) );
  NAND2_X1 U15474 ( .A1(n14343), .A2(n14588), .ZN(n13878) );
  NAND2_X1 U15475 ( .A1(n13879), .A2(n13878), .ZN(n14470) );
  INV_X1 U15476 ( .A(n14467), .ZN(n13881) );
  OAI22_X1 U15477 ( .A1(n13881), .A2(n13970), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13880), .ZN(n13882) );
  AOI21_X1 U15478 ( .B1(n14470), .B2(n13972), .A(n13882), .ZN(n13883) );
  OAI211_X1 U15479 ( .C1(n14740), .C2(n13975), .A(n13884), .B(n13883), .ZN(
        P2_U3186) );
  INV_X1 U15480 ( .A(n13885), .ZN(n13892) );
  AOI22_X1 U15481 ( .A1(n13886), .A2(n13990), .B1(n13894), .B2(n14346), .ZN(
        n13891) );
  AND2_X1 U15482 ( .A1(n14347), .A2(n14588), .ZN(n13887) );
  AOI21_X1 U15483 ( .B1(n14345), .B2(n14589), .A(n13887), .ZN(n14522) );
  AOI22_X1 U15484 ( .A1(n13985), .A2(n14526), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13888) );
  OAI21_X1 U15485 ( .B1(n14522), .B2(n13988), .A(n13888), .ZN(n13889) );
  AOI21_X1 U15486 ( .B1(n14671), .B2(n13983), .A(n13889), .ZN(n13890) );
  OAI21_X1 U15487 ( .B1(n13892), .B2(n13891), .A(n13890), .ZN(P2_U3188) );
  INV_X1 U15488 ( .A(n14596), .ZN(n14759) );
  OAI21_X1 U15489 ( .B1(n7593), .B2(n13893), .A(n13990), .ZN(n13897) );
  NAND3_X1 U15490 ( .A1(n13895), .A2(n13894), .A3(n14587), .ZN(n13896) );
  NAND2_X1 U15491 ( .A1(n13897), .A2(n13896), .ZN(n13899) );
  NAND2_X1 U15492 ( .A1(n13899), .A2(n13898), .ZN(n13906) );
  NAND2_X1 U15493 ( .A1(n13985), .A2(n14597), .ZN(n13900) );
  NAND2_X1 U15494 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14422)
         );
  OAI211_X1 U15495 ( .C1(n13902), .C2(n13901), .A(n13900), .B(n14422), .ZN(
        n13903) );
  AOI21_X1 U15496 ( .B1(n13904), .B2(n14590), .A(n13903), .ZN(n13905) );
  OAI211_X1 U15497 ( .C1(n14759), .C2(n13975), .A(n13906), .B(n13905), .ZN(
        P2_U3191) );
  INV_X1 U15498 ( .A(n14342), .ZN(n13907) );
  NOR3_X1 U15499 ( .A1(n13908), .A2(n13907), .A3(n13976), .ZN(n13909) );
  AOI21_X1 U15500 ( .B1(n13910), .B2(n13990), .A(n13909), .ZN(n13922) );
  MUX2_X1 U15501 ( .A(n14193), .B(n14312), .S(n7437), .Z(n13911) );
  XNOR2_X1 U15502 ( .A(n13911), .B(n10884), .ZN(n13921) );
  INV_X1 U15503 ( .A(n13912), .ZN(n14455) );
  AOI22_X1 U15504 ( .A1(n14455), .A2(n13985), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13913) );
  OAI21_X1 U15505 ( .B1(n13914), .B2(n13988), .A(n13913), .ZN(n13915) );
  AOI21_X1 U15506 ( .B1(n14193), .B2(n13983), .A(n13915), .ZN(n13920) );
  INV_X1 U15507 ( .A(n13916), .ZN(n13917) );
  NAND4_X1 U15508 ( .A1(n13918), .A2(n13990), .A3(n13917), .A4(n13921), .ZN(
        n13919) );
  OAI211_X1 U15509 ( .C1(n13922), .C2(n13921), .A(n13920), .B(n13919), .ZN(
        P2_U3192) );
  OAI211_X1 U15510 ( .C1(n13923), .C2(n13925), .A(n13924), .B(n13990), .ZN(
        n13929) );
  OAI22_X1 U15511 ( .A1(n14172), .A2(n13968), .B1(n13958), .B2(n13967), .ZN(
        n14548) );
  OAI22_X1 U15512 ( .A1(n13970), .A2(n14552), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13926), .ZN(n13927) );
  AOI21_X1 U15513 ( .B1(n13972), .B2(n14548), .A(n13927), .ZN(n13928) );
  OAI211_X1 U15514 ( .C1(n14551), .C2(n13975), .A(n13929), .B(n13928), .ZN(
        P2_U3195) );
  NAND2_X1 U15515 ( .A1(n13931), .A2(n13932), .ZN(n13936) );
  NOR3_X1 U15516 ( .A1(n13934), .A2(n13933), .A3(n13976), .ZN(n13935) );
  AOI21_X1 U15517 ( .B1(n13936), .B2(n13990), .A(n13935), .ZN(n13941) );
  AND2_X1 U15518 ( .A1(n14345), .A2(n14588), .ZN(n13937) );
  AOI21_X1 U15519 ( .B1(n14343), .B2(n14589), .A(n13937), .ZN(n14493) );
  AOI22_X1 U15520 ( .A1(n13985), .A2(n14498), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13938) );
  OAI21_X1 U15521 ( .B1(n14493), .B2(n13988), .A(n13938), .ZN(n13939) );
  AOI21_X1 U15522 ( .B1(n14497), .B2(n13983), .A(n13939), .ZN(n13940) );
  OAI21_X1 U15523 ( .B1(n13930), .B2(n13941), .A(n13940), .ZN(P2_U3197) );
  OAI211_X1 U15524 ( .C1(n13943), .C2(n13942), .A(n13931), .B(n13990), .ZN(
        n13947) );
  NOR2_X1 U15525 ( .A1(n13970), .A2(n14512), .ZN(n13945) );
  AOI22_X1 U15526 ( .A1(n14344), .A2(n14589), .B1(n14588), .B2(n14346), .ZN(
        n14507) );
  NOR2_X1 U15527 ( .A1(n14507), .A2(n13988), .ZN(n13944) );
  AOI211_X1 U15528 ( .C1(P2_REG3_REG_24__SCAN_IN), .C2(P2_U3088), .A(n13945), 
        .B(n13944), .ZN(n13946) );
  OAI211_X1 U15529 ( .C1(n7963), .C2(n13975), .A(n13947), .B(n13946), .ZN(
        P2_U3201) );
  INV_X1 U15530 ( .A(n13923), .ZN(n13954) );
  INV_X1 U15531 ( .A(n13948), .ZN(n13950) );
  NAND2_X1 U15532 ( .A1(n13950), .A2(n13949), .ZN(n13952) );
  AOI22_X1 U15533 ( .A1(n13954), .A2(n13953), .B1(n13952), .B2(n13951), .ZN(
        n13962) );
  OAI22_X1 U15534 ( .A1(n14165), .A2(n13968), .B1(n14152), .B2(n13967), .ZN(
        n13955) );
  INV_X1 U15535 ( .A(n13955), .ZN(n14569) );
  INV_X1 U15536 ( .A(n13956), .ZN(n14574) );
  AOI22_X1 U15537 ( .A1(n13985), .A2(n14574), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13957) );
  OAI21_X1 U15538 ( .B1(n13988), .B2(n14569), .A(n13957), .ZN(n13960) );
  NOR3_X1 U15539 ( .A1(n13923), .A2(n13958), .A3(n13976), .ZN(n13959) );
  AOI211_X1 U15540 ( .C1(n14688), .C2(n13983), .A(n13960), .B(n13959), .ZN(
        n13961) );
  OAI21_X1 U15541 ( .B1(n13962), .B2(n13963), .A(n13961), .ZN(P2_U3205) );
  AOI211_X1 U15542 ( .C1(n13965), .C2(n13964), .A(n13963), .B(n7593), .ZN(
        n13966) );
  INV_X1 U15543 ( .A(n13966), .ZN(n13974) );
  OAI22_X1 U15544 ( .A1(n14152), .A2(n13968), .B1(n14133), .B2(n13967), .ZN(
        n14605) );
  OAI22_X1 U15545 ( .A1(n13970), .A2(n14614), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13969), .ZN(n13971) );
  AOI21_X1 U15546 ( .B1(n13972), .B2(n14605), .A(n13971), .ZN(n13973) );
  OAI211_X1 U15547 ( .C1(n9109), .C2(n13975), .A(n13974), .B(n13973), .ZN(
        P2_U3210) );
  NOR3_X1 U15548 ( .A1(n13978), .A2(n13977), .A3(n13976), .ZN(n13979) );
  AOI21_X1 U15549 ( .B1(n13930), .B2(n13990), .A(n13979), .ZN(n13993) );
  INV_X1 U15550 ( .A(n13980), .ZN(n13992) );
  AND2_X1 U15551 ( .A1(n14344), .A2(n14588), .ZN(n13982) );
  AOI21_X1 U15552 ( .B1(n14342), .B2(n14589), .A(n13982), .ZN(n14479) );
  NAND2_X1 U15553 ( .A1(n14482), .A2(n13983), .ZN(n13987) );
  INV_X1 U15554 ( .A(n13984), .ZN(n14483) );
  AOI22_X1 U15555 ( .A1(n14483), .A2(n13985), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13986) );
  OAI211_X1 U15556 ( .C1(n14479), .C2(n13988), .A(n13987), .B(n13986), .ZN(
        n13989) );
  OAI21_X1 U15557 ( .B1(n13993), .B2(n13992), .A(n13991), .ZN(P2_U3212) );
  NAND2_X1 U15558 ( .A1(n14332), .A2(n13996), .ZN(n13999) );
  NAND2_X1 U15559 ( .A1(n13994), .A2(n13999), .ZN(n13995) );
  NAND2_X1 U15560 ( .A1(n14000), .A2(n13995), .ZN(n13998) );
  INV_X1 U15561 ( .A(n13996), .ZN(n13997) );
  NAND2_X1 U15562 ( .A1(n13998), .A2(n14013), .ZN(n14003) );
  OAI211_X1 U15563 ( .C1(n14001), .C2(n14040), .A(n14000), .B(n13999), .ZN(
        n14002) );
  NAND2_X1 U15564 ( .A1(n14003), .A2(n14002), .ZN(n14009) );
  NAND2_X1 U15565 ( .A1(n14366), .A2(n14013), .ZN(n14005) );
  NAND2_X1 U15566 ( .A1(n14040), .A2(n14006), .ZN(n14004) );
  NAND2_X1 U15567 ( .A1(n14005), .A2(n14004), .ZN(n14008) );
  AOI22_X1 U15568 ( .A1(n14366), .A2(n14040), .B1(n14006), .B2(n14013), .ZN(
        n14007) );
  INV_X1 U15569 ( .A(n14017), .ZN(n14010) );
  NAND2_X1 U15570 ( .A1(n14010), .A2(n14020), .ZN(n14015) );
  NAND2_X1 U15571 ( .A1(n14365), .A2(n14031), .ZN(n14012) );
  NAND2_X1 U15572 ( .A1(n14012), .A2(n14011), .ZN(n14018) );
  AOI22_X1 U15573 ( .A1(n14365), .A2(n14013), .B1(n14235), .B2(n16381), .ZN(
        n14014) );
  AOI21_X1 U15574 ( .B1(n14015), .B2(n14018), .A(n14014), .ZN(n14016) );
  INV_X1 U15575 ( .A(n14016), .ZN(n14024) );
  INV_X1 U15576 ( .A(n14018), .ZN(n14019) );
  NAND2_X1 U15577 ( .A1(n14020), .A2(n14019), .ZN(n14021) );
  NOR2_X1 U15578 ( .A1(n14017), .A2(n14021), .ZN(n14022) );
  INV_X1 U15579 ( .A(n14022), .ZN(n14023) );
  NAND2_X1 U15580 ( .A1(n14027), .A2(n14031), .ZN(n14026) );
  NAND2_X1 U15581 ( .A1(n14364), .A2(n14013), .ZN(n14025) );
  NAND2_X1 U15582 ( .A1(n14027), .A2(n14256), .ZN(n14029) );
  INV_X1 U15583 ( .A(n14013), .ZN(n14031) );
  NAND2_X1 U15584 ( .A1(n14364), .A2(n14031), .ZN(n14028) );
  NAND2_X1 U15585 ( .A1(n14029), .A2(n14028), .ZN(n14030) );
  INV_X2 U15586 ( .A(n14235), .ZN(n14197) );
  NAND2_X1 U15587 ( .A1(n14034), .A2(n14197), .ZN(n14033) );
  NAND2_X1 U15588 ( .A1(n14363), .A2(n14031), .ZN(n14032) );
  NAND2_X1 U15589 ( .A1(n14033), .A2(n14032), .ZN(n14036) );
  AOI22_X1 U15590 ( .A1(n14034), .A2(n14031), .B1(n14363), .B2(n14197), .ZN(
        n14035) );
  NAND2_X1 U15591 ( .A1(n14041), .A2(n14031), .ZN(n14039) );
  NAND2_X1 U15592 ( .A1(n14362), .A2(n14197), .ZN(n14038) );
  NAND2_X1 U15593 ( .A1(n14041), .A2(n14197), .ZN(n14042) );
  OAI21_X1 U15594 ( .B1(n14043), .B2(n14256), .A(n14042), .ZN(n14044) );
  NAND2_X1 U15595 ( .A1(n14047), .A2(n14197), .ZN(n14046) );
  INV_X2 U15596 ( .A(n14013), .ZN(n14262) );
  NAND2_X1 U15597 ( .A1(n14361), .A2(n14262), .ZN(n14045) );
  NAND2_X1 U15598 ( .A1(n14046), .A2(n14045), .ZN(n14050) );
  AOI22_X1 U15599 ( .A1(n14047), .A2(n14262), .B1(n14361), .B2(n14197), .ZN(
        n14048) );
  AOI21_X1 U15600 ( .B1(n14051), .B2(n14050), .A(n14048), .ZN(n14049) );
  INV_X1 U15601 ( .A(n14049), .ZN(n14052) );
  NAND2_X1 U15602 ( .A1(n14055), .A2(n14262), .ZN(n14054) );
  NAND2_X1 U15603 ( .A1(n14360), .A2(n14197), .ZN(n14053) );
  NAND2_X1 U15604 ( .A1(n14055), .A2(n14197), .ZN(n14056) );
  OAI21_X1 U15605 ( .B1(n14057), .B2(n14256), .A(n14056), .ZN(n14058) );
  NAND2_X1 U15606 ( .A1(n14061), .A2(n14197), .ZN(n14060) );
  NAND2_X1 U15607 ( .A1(n14359), .A2(n14262), .ZN(n14059) );
  NAND2_X1 U15608 ( .A1(n14060), .A2(n14059), .ZN(n14063) );
  AOI22_X1 U15609 ( .A1(n14061), .A2(n14262), .B1(n14359), .B2(n14197), .ZN(
        n14062) );
  AOI21_X1 U15610 ( .B1(n14064), .B2(n14063), .A(n14062), .ZN(n14066) );
  NOR2_X1 U15611 ( .A1(n14064), .A2(n14063), .ZN(n14065) );
  NAND2_X1 U15612 ( .A1(n14629), .A2(n14262), .ZN(n14068) );
  NAND2_X1 U15613 ( .A1(n14358), .A2(n14197), .ZN(n14067) );
  NAND2_X1 U15614 ( .A1(n14068), .A2(n14067), .ZN(n14070) );
  AOI22_X1 U15615 ( .A1(n14629), .A2(n14197), .B1(n14262), .B2(n14358), .ZN(
        n14069) );
  NAND2_X1 U15616 ( .A1(n14073), .A2(n14197), .ZN(n14072) );
  NAND2_X1 U15617 ( .A1(n14357), .A2(n14262), .ZN(n14071) );
  NAND2_X1 U15618 ( .A1(n14072), .A2(n14071), .ZN(n14079) );
  NAND2_X1 U15619 ( .A1(n14078), .A2(n14079), .ZN(n14077) );
  NAND2_X1 U15620 ( .A1(n14073), .A2(n14262), .ZN(n14074) );
  OAI21_X1 U15621 ( .B1(n14075), .B2(n14235), .A(n14074), .ZN(n14076) );
  NAND2_X1 U15622 ( .A1(n14077), .A2(n14076), .ZN(n14083) );
  INV_X1 U15623 ( .A(n14078), .ZN(n14081) );
  NAND2_X1 U15624 ( .A1(n14081), .A2(n14080), .ZN(n14082) );
  NAND2_X1 U15625 ( .A1(n14083), .A2(n14082), .ZN(n14089) );
  NAND2_X1 U15626 ( .A1(n14086), .A2(n14262), .ZN(n14085) );
  NAND2_X1 U15627 ( .A1(n14356), .A2(n14197), .ZN(n14084) );
  NAND2_X1 U15628 ( .A1(n14085), .A2(n14084), .ZN(n14088) );
  AOI22_X1 U15629 ( .A1(n14086), .A2(n14197), .B1(n14262), .B2(n14356), .ZN(
        n14087) );
  AOI21_X1 U15630 ( .B1(n14089), .B2(n14088), .A(n14087), .ZN(n14091) );
  NOR2_X1 U15631 ( .A1(n14089), .A2(n14088), .ZN(n14090) );
  NAND2_X1 U15632 ( .A1(n14094), .A2(n14197), .ZN(n14093) );
  NAND2_X1 U15633 ( .A1(n14355), .A2(n14262), .ZN(n14092) );
  NAND2_X1 U15634 ( .A1(n14094), .A2(n14262), .ZN(n14095) );
  OAI21_X1 U15635 ( .B1(n14096), .B2(n14235), .A(n14095), .ZN(n14097) );
  NAND2_X1 U15636 ( .A1(n7765), .A2(n14262), .ZN(n14100) );
  NAND2_X1 U15637 ( .A1(n14354), .A2(n14197), .ZN(n14099) );
  NAND2_X1 U15638 ( .A1(n14100), .A2(n14099), .ZN(n14103) );
  AOI22_X1 U15639 ( .A1(n7765), .A2(n14197), .B1(n14262), .B2(n14354), .ZN(
        n14102) );
  NAND2_X1 U15640 ( .A1(n14725), .A2(n14197), .ZN(n14105) );
  NAND2_X1 U15641 ( .A1(n14353), .A2(n14262), .ZN(n14104) );
  NAND2_X1 U15642 ( .A1(n14105), .A2(n14104), .ZN(n14111) );
  NAND2_X1 U15643 ( .A1(n14110), .A2(n14111), .ZN(n14109) );
  NAND2_X1 U15644 ( .A1(n14725), .A2(n14262), .ZN(n14106) );
  OAI21_X1 U15645 ( .B1(n14107), .B2(n14235), .A(n14106), .ZN(n14108) );
  NAND2_X1 U15646 ( .A1(n14109), .A2(n14108), .ZN(n14115) );
  INV_X1 U15647 ( .A(n14110), .ZN(n14113) );
  INV_X1 U15648 ( .A(n14111), .ZN(n14112) );
  NAND2_X1 U15649 ( .A1(n14113), .A2(n14112), .ZN(n14114) );
  NAND2_X1 U15650 ( .A1(n7757), .A2(n14262), .ZN(n14117) );
  NAND2_X1 U15651 ( .A1(n14352), .A2(n14197), .ZN(n14116) );
  AOI22_X1 U15652 ( .A1(n7757), .A2(n14197), .B1(n14262), .B2(n14352), .ZN(
        n14118) );
  INV_X1 U15653 ( .A(n14118), .ZN(n14119) );
  NAND2_X1 U15654 ( .A1(n14122), .A2(n14256), .ZN(n14121) );
  NAND2_X1 U15655 ( .A1(n14351), .A2(n14262), .ZN(n14120) );
  NAND2_X1 U15656 ( .A1(n14121), .A2(n14120), .ZN(n14125) );
  AOI22_X1 U15657 ( .A1(n14122), .A2(n14262), .B1(n14351), .B2(n14256), .ZN(
        n14123) );
  AOI21_X1 U15658 ( .B1(n14126), .B2(n14125), .A(n14123), .ZN(n14124) );
  INV_X1 U15659 ( .A(n14124), .ZN(n14129) );
  NOR2_X1 U15660 ( .A1(n14126), .A2(n14125), .ZN(n14127) );
  INV_X1 U15661 ( .A(n14127), .ZN(n14128) );
  NAND2_X1 U15662 ( .A1(n14763), .A2(n14262), .ZN(n14131) );
  NAND2_X1 U15663 ( .A1(n14350), .A2(n14197), .ZN(n14130) );
  NAND2_X1 U15664 ( .A1(n14131), .A2(n14130), .ZN(n14137) );
  NAND2_X1 U15665 ( .A1(n14136), .A2(n14137), .ZN(n14135) );
  NAND2_X1 U15666 ( .A1(n14763), .A2(n14197), .ZN(n14132) );
  OAI21_X1 U15667 ( .B1(n14133), .B2(n14256), .A(n14132), .ZN(n14134) );
  NAND2_X1 U15668 ( .A1(n14135), .A2(n14134), .ZN(n14141) );
  INV_X1 U15669 ( .A(n14136), .ZN(n14139) );
  INV_X1 U15670 ( .A(n14137), .ZN(n14138) );
  NAND2_X1 U15671 ( .A1(n14139), .A2(n14138), .ZN(n14140) );
  NAND2_X1 U15672 ( .A1(n14698), .A2(n14256), .ZN(n14143) );
  NAND2_X1 U15673 ( .A1(n14587), .A2(n14262), .ZN(n14142) );
  NAND2_X1 U15674 ( .A1(n14143), .A2(n14142), .ZN(n14145) );
  AOI22_X1 U15675 ( .A1(n14698), .A2(n14262), .B1(n14587), .B2(n14197), .ZN(
        n14144) );
  AOI21_X1 U15676 ( .B1(n14146), .B2(n14145), .A(n14144), .ZN(n14148) );
  NOR2_X1 U15677 ( .A1(n14146), .A2(n14145), .ZN(n14147) );
  NAND2_X1 U15678 ( .A1(n14596), .A2(n14262), .ZN(n14150) );
  NAND2_X1 U15679 ( .A1(n14349), .A2(n14256), .ZN(n14149) );
  NAND2_X1 U15680 ( .A1(n14150), .A2(n14149), .ZN(n14156) );
  NAND2_X1 U15681 ( .A1(n14155), .A2(n14156), .ZN(n14154) );
  NAND2_X1 U15682 ( .A1(n14596), .A2(n14197), .ZN(n14151) );
  OAI21_X1 U15683 ( .B1(n14152), .B2(n14013), .A(n14151), .ZN(n14153) );
  NAND2_X1 U15684 ( .A1(n14154), .A2(n14153), .ZN(n14160) );
  INV_X1 U15685 ( .A(n14155), .ZN(n14158) );
  INV_X1 U15686 ( .A(n14156), .ZN(n14157) );
  NAND2_X1 U15687 ( .A1(n14158), .A2(n14157), .ZN(n14159) );
  NAND2_X1 U15688 ( .A1(n14688), .A2(n14197), .ZN(n14162) );
  NAND2_X1 U15689 ( .A1(n14590), .A2(n14031), .ZN(n14161) );
  AOI22_X1 U15690 ( .A1(n14688), .A2(n14262), .B1(n14590), .B2(n14256), .ZN(
        n14163) );
  INV_X1 U15691 ( .A(n14163), .ZN(n14164) );
  INV_X1 U15692 ( .A(n14168), .ZN(n14171) );
  OAI22_X1 U15693 ( .A1(n14551), .A2(n14256), .B1(n14165), .B2(n14235), .ZN(
        n14167) );
  INV_X1 U15694 ( .A(n14167), .ZN(n14170) );
  AOI22_X1 U15695 ( .A1(n14681), .A2(n14197), .B1(n14262), .B2(n14348), .ZN(
        n14166) );
  AOI21_X1 U15696 ( .B1(n14168), .B2(n14167), .A(n14166), .ZN(n14169) );
  AOI22_X1 U15697 ( .A1(n14675), .A2(n14197), .B1(n14031), .B2(n14347), .ZN(
        n14175) );
  OAI22_X1 U15698 ( .A1(n14173), .A2(n14013), .B1(n14172), .B2(n14235), .ZN(
        n14174) );
  OAI22_X1 U15699 ( .A1(n14529), .A2(n14013), .B1(n14177), .B2(n14235), .ZN(
        n14191) );
  AND2_X1 U15700 ( .A1(n14345), .A2(n14262), .ZN(n14178) );
  AOI21_X1 U15701 ( .B1(n14511), .B2(n14256), .A(n14178), .ZN(n14203) );
  NAND2_X1 U15702 ( .A1(n14511), .A2(n14262), .ZN(n14180) );
  NAND2_X1 U15703 ( .A1(n14345), .A2(n14256), .ZN(n14179) );
  NAND2_X1 U15704 ( .A1(n14180), .A2(n14179), .ZN(n14202) );
  AND2_X1 U15705 ( .A1(n14343), .A2(n14197), .ZN(n14181) );
  AOI21_X1 U15706 ( .B1(n14482), .B2(n14031), .A(n14181), .ZN(n14215) );
  NAND2_X1 U15707 ( .A1(n14482), .A2(n14256), .ZN(n14183) );
  NAND2_X1 U15708 ( .A1(n14343), .A2(n14262), .ZN(n14182) );
  NAND2_X1 U15709 ( .A1(n14183), .A2(n14182), .ZN(n14214) );
  NAND2_X1 U15710 ( .A1(n14215), .A2(n14214), .ZN(n14211) );
  AND2_X1 U15711 ( .A1(n14344), .A2(n14197), .ZN(n14184) );
  AOI21_X1 U15712 ( .B1(n14497), .B2(n14262), .A(n14184), .ZN(n14208) );
  NAND2_X1 U15713 ( .A1(n14497), .A2(n14197), .ZN(n14186) );
  NAND2_X1 U15714 ( .A1(n14344), .A2(n14031), .ZN(n14185) );
  NAND2_X1 U15715 ( .A1(n14186), .A2(n14185), .ZN(n14207) );
  NAND2_X1 U15716 ( .A1(n14208), .A2(n14207), .ZN(n14187) );
  AND2_X1 U15717 ( .A1(n14211), .A2(n14187), .ZN(n14201) );
  OAI21_X1 U15718 ( .B1(n14203), .B2(n14202), .A(n14201), .ZN(n14188) );
  INV_X1 U15719 ( .A(n14188), .ZN(n14189) );
  AOI22_X1 U15720 ( .A1(n14671), .A2(n14197), .B1(n14262), .B2(n14346), .ZN(
        n14190) );
  AND2_X1 U15721 ( .A1(n14341), .A2(n14262), .ZN(n14192) );
  AOI21_X1 U15722 ( .B1(n14193), .B2(n14197), .A(n14192), .ZN(n14242) );
  NAND2_X1 U15723 ( .A1(n14193), .A2(n14262), .ZN(n14195) );
  NAND2_X1 U15724 ( .A1(n14341), .A2(n14197), .ZN(n14194) );
  NAND2_X1 U15725 ( .A1(n14195), .A2(n14194), .ZN(n14241) );
  AND2_X1 U15726 ( .A1(n14342), .A2(n14262), .ZN(n14196) );
  AOI21_X1 U15727 ( .B1(n14198), .B2(n14197), .A(n14196), .ZN(n14240) );
  NAND2_X1 U15728 ( .A1(n14198), .A2(n14031), .ZN(n14200) );
  NAND2_X1 U15729 ( .A1(n14342), .A2(n14197), .ZN(n14199) );
  NAND2_X1 U15730 ( .A1(n14200), .A2(n14199), .ZN(n14239) );
  INV_X1 U15731 ( .A(n14201), .ZN(n14206) );
  INV_X1 U15732 ( .A(n14202), .ZN(n14205) );
  INV_X1 U15733 ( .A(n14203), .ZN(n14204) );
  OR3_X1 U15734 ( .A1(n14206), .A2(n14205), .A3(n14204), .ZN(n14213) );
  INV_X1 U15735 ( .A(n14207), .ZN(n14210) );
  INV_X1 U15736 ( .A(n14208), .ZN(n14209) );
  NAND3_X1 U15737 ( .A1(n14211), .A2(n14210), .A3(n14209), .ZN(n14212) );
  OAI211_X1 U15738 ( .C1(n14215), .C2(n14214), .A(n14213), .B(n14212), .ZN(
        n14216) );
  INV_X1 U15739 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n14639) );
  OR2_X1 U15740 ( .A1(n8851), .A2(n14639), .ZN(n14222) );
  INV_X1 U15741 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14730) );
  OR2_X1 U15742 ( .A1(n14219), .A2(n14730), .ZN(n14220) );
  AND3_X1 U15743 ( .A1(n14222), .A2(n14221), .A3(n14220), .ZN(n14434) );
  INV_X1 U15744 ( .A(n14434), .ZN(n14338) );
  INV_X1 U15745 ( .A(n14225), .ZN(n14227) );
  XNOR2_X1 U15746 ( .A(n14228), .B(SI_31_), .ZN(n14229) );
  NAND2_X1 U15747 ( .A1(n15207), .A2(n8612), .ZN(n14233) );
  OR2_X1 U15748 ( .A1(n14253), .A2(n14231), .ZN(n14232) );
  AOI22_X1 U15749 ( .A1(n14234), .A2(n14256), .B1(n14031), .B2(n14340), .ZN(
        n14264) );
  INV_X1 U15750 ( .A(n14264), .ZN(n14238) );
  OAI22_X1 U15751 ( .A1(n14447), .A2(n14013), .B1(n14236), .B2(n14235), .ZN(
        n14263) );
  NAND2_X1 U15752 ( .A1(n14238), .A2(n14237), .ZN(n14247) );
  NOR2_X1 U15753 ( .A1(n14240), .A2(n14239), .ZN(n14245) );
  INV_X1 U15754 ( .A(n14241), .ZN(n14244) );
  INV_X1 U15755 ( .A(n14242), .ZN(n14243) );
  AOI22_X1 U15756 ( .A1(n8515), .A2(n14245), .B1(n14244), .B2(n14243), .ZN(
        n14246) );
  NAND3_X1 U15757 ( .A1(n14250), .A2(n14249), .A3(n14248), .ZN(n14268) );
  MUX2_X1 U15758 ( .A(n14434), .B(n14256), .S(n14435), .Z(n14251) );
  AOI21_X1 U15759 ( .B1(n14262), .B2(n14338), .A(n14251), .ZN(n14266) );
  NAND2_X1 U15760 ( .A1(n15200), .A2(n8612), .ZN(n14255) );
  INV_X1 U15761 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n14777) );
  OR2_X1 U15762 ( .A1(n14253), .A2(n14777), .ZN(n14254) );
  NAND2_X1 U15763 ( .A1(n14338), .A2(n14256), .ZN(n14272) );
  INV_X1 U15764 ( .A(n14257), .ZN(n14258) );
  NAND2_X1 U15765 ( .A1(n14258), .A2(n14286), .ZN(n14277) );
  NAND3_X1 U15766 ( .A1(n14272), .A2(n14259), .A3(n14277), .ZN(n14260) );
  AOI22_X1 U15767 ( .A1(n14429), .A2(n14031), .B1(n14339), .B2(n14260), .ZN(
        n14261) );
  INV_X1 U15768 ( .A(n14261), .ZN(n14270) );
  AOI22_X1 U15769 ( .A1(n14429), .A2(n14197), .B1(n14262), .B2(n14339), .ZN(
        n14269) );
  AOI22_X1 U15770 ( .A1(n14270), .A2(n14269), .B1(n14264), .B2(n14263), .ZN(
        n14265) );
  NAND2_X1 U15771 ( .A1(n14268), .A2(n14267), .ZN(n14271) );
  NAND2_X1 U15772 ( .A1(n14271), .A2(n8508), .ZN(n14275) );
  MUX2_X1 U15773 ( .A(n14338), .B(n14013), .S(n14435), .Z(n14273) );
  NAND2_X1 U15774 ( .A1(n14273), .A2(n14272), .ZN(n14274) );
  NAND2_X1 U15775 ( .A1(n14275), .A2(n14274), .ZN(n14330) );
  AOI21_X1 U15776 ( .B1(n14323), .B2(n14276), .A(n7431), .ZN(n14283) );
  OAI21_X1 U15777 ( .B1(n14278), .B2(n14424), .A(n14277), .ZN(n14279) );
  NAND2_X1 U15778 ( .A1(n14330), .A2(n14280), .ZN(n14281) );
  OAI211_X1 U15779 ( .C1(n14330), .C2(n14283), .A(n14282), .B(n14281), .ZN(
        n14337) );
  XOR2_X1 U15780 ( .A(n14339), .B(n14429), .Z(n14317) );
  XOR2_X1 U15781 ( .A(n14346), .B(n14671), .Z(n14520) );
  NOR4_X1 U15782 ( .A1(n14287), .A2(n14286), .A3(n14285), .A4(n14284), .ZN(
        n14291) );
  NAND4_X1 U15783 ( .A1(n14291), .A2(n14290), .A3(n14289), .A4(n14288), .ZN(
        n14292) );
  NOR4_X1 U15784 ( .A1(n14295), .A2(n14294), .A3(n14293), .A4(n14292), .ZN(
        n14298) );
  NAND4_X1 U15785 ( .A1(n14299), .A2(n14298), .A3(n14297), .A4(n14296), .ZN(
        n14300) );
  NOR4_X1 U15786 ( .A1(n14303), .A2(n14302), .A3(n14301), .A4(n14300), .ZN(
        n14306) );
  NAND4_X1 U15787 ( .A1(n14567), .A2(n14306), .A3(n14305), .A4(n14304), .ZN(
        n14308) );
  NOR4_X1 U15788 ( .A1(n14308), .A2(n14586), .A3(n14609), .A4(n14307), .ZN(
        n14309) );
  NAND4_X1 U15789 ( .A1(n14310), .A2(n14309), .A3(n14541), .A4(n14558), .ZN(
        n14311) );
  NOR4_X1 U15790 ( .A1(n14312), .A2(n14505), .A3(n14520), .A4(n14311), .ZN(
        n14315) );
  NAND4_X1 U15791 ( .A1(n14315), .A2(n14314), .A3(n14462), .A4(n14313), .ZN(
        n14316) );
  NOR3_X1 U15792 ( .A1(n14318), .A2(n14317), .A3(n14316), .ZN(n14319) );
  XNOR2_X1 U15793 ( .A(n14319), .B(n7431), .ZN(n14321) );
  NOR3_X1 U15794 ( .A1(n14321), .A2(n14320), .A3(n14327), .ZN(n14322) );
  OAI21_X1 U15795 ( .B1(n14330), .B2(n14323), .A(n14322), .ZN(n14336) );
  NAND3_X1 U15796 ( .A1(n14588), .A2(n14325), .A3(n14324), .ZN(n14329) );
  NOR2_X1 U15797 ( .A1(n14327), .A2(n14326), .ZN(n14331) );
  INV_X1 U15798 ( .A(n14331), .ZN(n14328) );
  OAI211_X1 U15799 ( .C1(n15822), .C2(n14329), .A(P2_B_REG_SCAN_IN), .B(n14328), .ZN(n14335) );
  INV_X1 U15800 ( .A(n14330), .ZN(n14333) );
  NAND3_X1 U15801 ( .A1(n14333), .A2(n14332), .A3(n14331), .ZN(n14334) );
  NAND4_X1 U15802 ( .A1(n14337), .A2(n14336), .A3(n14335), .A4(n14334), .ZN(
        P2_U3328) );
  MUX2_X1 U15803 ( .A(n14338), .B(P2_DATAO_REG_31__SCAN_IN), .S(n14367), .Z(
        P2_U3562) );
  MUX2_X1 U15804 ( .A(n14339), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14367), .Z(
        P2_U3561) );
  MUX2_X1 U15805 ( .A(n14340), .B(P2_DATAO_REG_29__SCAN_IN), .S(n14367), .Z(
        P2_U3560) );
  MUX2_X1 U15806 ( .A(n14341), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14367), .Z(
        P2_U3559) );
  MUX2_X1 U15807 ( .A(n14342), .B(P2_DATAO_REG_27__SCAN_IN), .S(n14367), .Z(
        P2_U3558) );
  MUX2_X1 U15808 ( .A(n14343), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14367), .Z(
        P2_U3557) );
  MUX2_X1 U15809 ( .A(n14344), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14367), .Z(
        P2_U3556) );
  MUX2_X1 U15810 ( .A(n14345), .B(P2_DATAO_REG_24__SCAN_IN), .S(n14367), .Z(
        P2_U3555) );
  MUX2_X1 U15811 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n14346), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15812 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n14347), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U15813 ( .A(n14348), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14367), .Z(
        P2_U3552) );
  MUX2_X1 U15814 ( .A(n14590), .B(P2_DATAO_REG_20__SCAN_IN), .S(n14367), .Z(
        P2_U3551) );
  MUX2_X1 U15815 ( .A(n14349), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14367), .Z(
        P2_U3550) );
  MUX2_X1 U15816 ( .A(n14587), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14367), .Z(
        P2_U3549) );
  MUX2_X1 U15817 ( .A(n14350), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14367), .Z(
        P2_U3548) );
  MUX2_X1 U15818 ( .A(n14351), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14367), .Z(
        P2_U3547) );
  MUX2_X1 U15819 ( .A(n14352), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14367), .Z(
        P2_U3546) );
  MUX2_X1 U15820 ( .A(n14353), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14367), .Z(
        P2_U3545) );
  MUX2_X1 U15821 ( .A(n14354), .B(P2_DATAO_REG_13__SCAN_IN), .S(n14367), .Z(
        P2_U3544) );
  MUX2_X1 U15822 ( .A(n14355), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14367), .Z(
        P2_U3543) );
  MUX2_X1 U15823 ( .A(n14356), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14367), .Z(
        P2_U3542) );
  MUX2_X1 U15824 ( .A(n14357), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14367), .Z(
        P2_U3541) );
  MUX2_X1 U15825 ( .A(n14358), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14367), .Z(
        P2_U3540) );
  MUX2_X1 U15826 ( .A(n14359), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14367), .Z(
        P2_U3539) );
  MUX2_X1 U15827 ( .A(n14360), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14367), .Z(
        P2_U3538) );
  MUX2_X1 U15828 ( .A(n14361), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14367), .Z(
        P2_U3537) );
  MUX2_X1 U15829 ( .A(n14362), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14367), .Z(
        P2_U3536) );
  MUX2_X1 U15830 ( .A(n14363), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14367), .Z(
        P2_U3535) );
  MUX2_X1 U15831 ( .A(n14364), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14367), .Z(
        P2_U3534) );
  MUX2_X1 U15832 ( .A(n14365), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14367), .Z(
        P2_U3533) );
  MUX2_X1 U15833 ( .A(n14366), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14367), .Z(
        P2_U3532) );
  MUX2_X1 U15834 ( .A(n13994), .B(P2_DATAO_REG_0__SCAN_IN), .S(n14367), .Z(
        P2_U3531) );
  INV_X1 U15835 ( .A(n15842), .ZN(n15860) );
  INV_X1 U15836 ( .A(n14381), .ZN(n14368) );
  AOI211_X1 U15837 ( .C1(n14370), .C2(n14369), .A(n14368), .B(n15848), .ZN(
        n14371) );
  AOI21_X1 U15838 ( .B1(n15860), .B2(n14372), .A(n14371), .ZN(n14378) );
  AOI22_X1 U15839 ( .A1(n15875), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n14377) );
  OAI21_X1 U15840 ( .B1(n10534), .B2(n14374), .A(n14373), .ZN(n14375) );
  NAND3_X1 U15841 ( .A1(n15873), .A2(n14389), .A3(n14375), .ZN(n14376) );
  NAND3_X1 U15842 ( .A1(n14378), .A2(n14377), .A3(n14376), .ZN(P2_U3215) );
  AND3_X1 U15843 ( .A1(n14381), .A2(n14380), .A3(n14379), .ZN(n14382) );
  NOR3_X1 U15844 ( .A1(n15848), .A2(n14383), .A3(n14382), .ZN(n14384) );
  AOI21_X1 U15845 ( .B1(n15860), .B2(n14385), .A(n14384), .ZN(n14394) );
  AOI22_X1 U15846 ( .A1(n15875), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14393) );
  INV_X1 U15847 ( .A(n14386), .ZN(n14391) );
  NAND3_X1 U15848 ( .A1(n14389), .A2(n14388), .A3(n14387), .ZN(n14390) );
  NAND3_X1 U15849 ( .A1(n15873), .A2(n14391), .A3(n14390), .ZN(n14392) );
  NAND3_X1 U15850 ( .A1(n14394), .A2(n14393), .A3(n14392), .ZN(P2_U3216) );
  INV_X1 U15851 ( .A(n14395), .ZN(n14399) );
  NOR3_X1 U15852 ( .A1(n15826), .A2(n14397), .A3(n14396), .ZN(n14398) );
  NOR3_X1 U15853 ( .A1(n15848), .A2(n14399), .A3(n14398), .ZN(n14400) );
  AOI21_X1 U15854 ( .B1(n15860), .B2(n14401), .A(n14400), .ZN(n14410) );
  MUX2_X1 U15855 ( .A(n10501), .B(P2_REG1_REG_4__SCAN_IN), .S(n14401), .Z(
        n14404) );
  INV_X1 U15856 ( .A(n14402), .ZN(n14403) );
  NAND2_X1 U15857 ( .A1(n14404), .A2(n14403), .ZN(n14406) );
  OAI211_X1 U15858 ( .C1(n15831), .C2(n14406), .A(n15873), .B(n14405), .ZN(
        n14408) );
  NAND2_X1 U15859 ( .A1(n15875), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n14407) );
  NAND4_X1 U15860 ( .A1(n14410), .A2(n14409), .A3(n14408), .A4(n14407), .ZN(
        P2_U3218) );
  INV_X1 U15861 ( .A(n14411), .ZN(n14412) );
  AOI22_X1 U15862 ( .A1(n14414), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n14413), 
        .B2(n14412), .ZN(n14416) );
  XNOR2_X1 U15863 ( .A(n7431), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n14415) );
  XNOR2_X1 U15864 ( .A(n14416), .B(n14415), .ZN(n14428) );
  NOR2_X1 U15865 ( .A1(n14418), .A2(n14417), .ZN(n14421) );
  INV_X1 U15866 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14419) );
  MUX2_X1 U15867 ( .A(n14419), .B(P2_REG2_REG_19__SCAN_IN), .S(n7431), .Z(
        n14420) );
  XNOR2_X1 U15868 ( .A(n14421), .B(n14420), .ZN(n14426) );
  NAND2_X1 U15869 ( .A1(n15875), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n14423) );
  OAI211_X1 U15870 ( .C1(n15842), .C2(n14424), .A(n14423), .B(n14422), .ZN(
        n14425) );
  AOI21_X1 U15871 ( .B1(n14426), .B2(n15877), .A(n14425), .ZN(n14427) );
  OAI21_X1 U15872 ( .B1(n14428), .B2(n15830), .A(n14427), .ZN(P2_U3233) );
  NAND2_X1 U15873 ( .A1(n14736), .A2(n14439), .ZN(n14438) );
  INV_X1 U15874 ( .A(n14432), .ZN(n14433) );
  OR2_X1 U15875 ( .A1(n14434), .A2(n14433), .ZN(n14641) );
  NOR2_X1 U15876 ( .A1(n14622), .A2(n14641), .ZN(n14441) );
  INV_X1 U15877 ( .A(n14435), .ZN(n14732) );
  NOR2_X1 U15878 ( .A1(n14732), .A2(n14619), .ZN(n14436) );
  AOI211_X1 U15879 ( .C1(P2_REG2_REG_31__SCAN_IN), .C2(n14622), .A(n14441), 
        .B(n14436), .ZN(n14437) );
  OAI21_X1 U15880 ( .B1(n14556), .B2(n14638), .A(n14437), .ZN(P2_U3234) );
  OAI211_X1 U15881 ( .C1(n14736), .C2(n14439), .A(n14430), .B(n14438), .ZN(
        n14642) );
  NOR2_X1 U15882 ( .A1(n14736), .A2(n14619), .ZN(n14440) );
  AOI211_X1 U15883 ( .C1(n14622), .C2(P2_REG2_REG_30__SCAN_IN), .A(n14441), 
        .B(n14440), .ZN(n14442) );
  OAI21_X1 U15884 ( .B1(n14556), .B2(n14642), .A(n14442), .ZN(P2_U3235) );
  INV_X1 U15885 ( .A(n14443), .ZN(n14453) );
  INV_X1 U15886 ( .A(n14444), .ZN(n14445) );
  AOI22_X1 U15887 ( .A1(n14445), .A2(n14615), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14622), .ZN(n14446) );
  OAI21_X1 U15888 ( .B1(n14447), .B2(n14619), .A(n14446), .ZN(n14448) );
  AOI21_X1 U15889 ( .B1(n14449), .B2(n14632), .A(n14448), .ZN(n14452) );
  NAND2_X1 U15890 ( .A1(n14450), .A2(n14630), .ZN(n14451) );
  OAI211_X1 U15891 ( .C1(n14453), .C2(n14622), .A(n14452), .B(n14451), .ZN(
        P2_U3236) );
  NAND2_X1 U15892 ( .A1(n14454), .A2(n14632), .ZN(n14460) );
  AOI22_X1 U15893 ( .A1(n14455), .A2(n14615), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n14622), .ZN(n14456) );
  OAI21_X1 U15894 ( .B1(n14648), .B2(n14619), .A(n14456), .ZN(n14457) );
  AOI21_X1 U15895 ( .B1(n14458), .B2(n11368), .A(n14457), .ZN(n14459) );
  OAI211_X1 U15896 ( .C1(n14461), .C2(n14602), .A(n14460), .B(n14459), .ZN(
        P2_U3237) );
  NAND2_X1 U15897 ( .A1(n14463), .A2(n14462), .ZN(n14464) );
  NAND2_X1 U15898 ( .A1(n14465), .A2(n14464), .ZN(n14649) );
  OAI211_X1 U15899 ( .C1(n14481), .C2(n14740), .A(n14430), .B(n14466), .ZN(
        n14650) );
  INV_X1 U15900 ( .A(n14650), .ZN(n14474) );
  AOI22_X1 U15901 ( .A1(n14467), .A2(n14615), .B1(n14622), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n14468) );
  OAI21_X1 U15902 ( .B1(n14740), .B2(n14619), .A(n14468), .ZN(n14473) );
  XNOR2_X1 U15903 ( .A(n14469), .B(n9065), .ZN(n14471) );
  AOI21_X1 U15904 ( .B1(n14471), .B2(n14606), .A(n14470), .ZN(n14651) );
  NOR2_X1 U15905 ( .A1(n14651), .A2(n14622), .ZN(n14472) );
  AOI211_X1 U15906 ( .C1(n14474), .C2(n14632), .A(n14473), .B(n14472), .ZN(
        n14475) );
  OAI21_X1 U15907 ( .B1(n14580), .B2(n14649), .A(n14475), .ZN(P2_U3238) );
  OAI21_X1 U15908 ( .B1(n14477), .B2(n14478), .A(n14476), .ZN(n14656) );
  INV_X1 U15909 ( .A(n14656), .ZN(n14488) );
  OAI21_X1 U15910 ( .B1(n14480), .B2(n9148), .A(n14479), .ZN(n14654) );
  INV_X1 U15911 ( .A(n14482), .ZN(n14744) );
  AOI211_X1 U15912 ( .C1(n14482), .C2(n14495), .A(n7437), .B(n14481), .ZN(
        n14655) );
  NAND2_X1 U15913 ( .A1(n14655), .A2(n14632), .ZN(n14485) );
  AOI22_X1 U15914 ( .A1(n14622), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n14483), 
        .B2(n14615), .ZN(n14484) );
  OAI211_X1 U15915 ( .C1(n14744), .C2(n14619), .A(n14485), .B(n14484), .ZN(
        n14486) );
  AOI21_X1 U15916 ( .B1(n14654), .B2(n11368), .A(n14486), .ZN(n14487) );
  OAI21_X1 U15917 ( .B1(n14488), .B2(n14580), .A(n14487), .ZN(P2_U3239) );
  OAI21_X1 U15918 ( .B1(n14490), .B2(n14491), .A(n14489), .ZN(n14661) );
  INV_X1 U15919 ( .A(n14661), .ZN(n14503) );
  XNOR2_X1 U15920 ( .A(n14492), .B(n14491), .ZN(n14494) );
  OAI21_X1 U15921 ( .B1(n14494), .B2(n9148), .A(n14493), .ZN(n14659) );
  INV_X1 U15922 ( .A(n14497), .ZN(n14748) );
  INV_X1 U15923 ( .A(n14495), .ZN(n14496) );
  AOI211_X1 U15924 ( .C1(n14497), .C2(n14509), .A(n7437), .B(n14496), .ZN(
        n14660) );
  NAND2_X1 U15925 ( .A1(n14660), .A2(n14632), .ZN(n14500) );
  AOI22_X1 U15926 ( .A1(n14622), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n14498), 
        .B2(n14615), .ZN(n14499) );
  OAI211_X1 U15927 ( .C1(n14748), .C2(n14619), .A(n14500), .B(n14499), .ZN(
        n14501) );
  AOI21_X1 U15928 ( .B1(n14659), .B2(n11368), .A(n14501), .ZN(n14502) );
  OAI21_X1 U15929 ( .B1(n14503), .B2(n14580), .A(n14502), .ZN(P2_U3240) );
  OAI21_X1 U15930 ( .B1(n8219), .B2(n14505), .A(n14504), .ZN(n14666) );
  INV_X1 U15931 ( .A(n14666), .ZN(n14518) );
  XNOR2_X1 U15932 ( .A(n14506), .B(n14505), .ZN(n14508) );
  OAI21_X1 U15933 ( .B1(n14508), .B2(n9148), .A(n14507), .ZN(n14664) );
  INV_X1 U15934 ( .A(n14509), .ZN(n14510) );
  AOI211_X1 U15935 ( .C1(n14511), .C2(n14524), .A(n7437), .B(n14510), .ZN(
        n14665) );
  NAND2_X1 U15936 ( .A1(n14665), .A2(n14632), .ZN(n14515) );
  INV_X1 U15937 ( .A(n14512), .ZN(n14513) );
  AOI22_X1 U15938 ( .A1(n14622), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n14513), 
        .B2(n14615), .ZN(n14514) );
  OAI211_X1 U15939 ( .C1(n7963), .C2(n14619), .A(n14515), .B(n14514), .ZN(
        n14516) );
  AOI21_X1 U15940 ( .B1(n14664), .B2(n11368), .A(n14516), .ZN(n14517) );
  OAI21_X1 U15941 ( .B1(n14518), .B2(n14580), .A(n14517), .ZN(P2_U3241) );
  XNOR2_X1 U15942 ( .A(n14519), .B(n14520), .ZN(n14673) );
  XNOR2_X1 U15943 ( .A(n14521), .B(n14520), .ZN(n14523) );
  OAI21_X1 U15944 ( .B1(n14523), .B2(n9148), .A(n14522), .ZN(n14669) );
  INV_X1 U15945 ( .A(n14524), .ZN(n14525) );
  AOI211_X1 U15946 ( .C1(n14671), .C2(n7967), .A(n7437), .B(n14525), .ZN(
        n14670) );
  NAND2_X1 U15947 ( .A1(n14670), .A2(n14632), .ZN(n14528) );
  AOI22_X1 U15948 ( .A1(n14622), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n14526), 
        .B2(n14615), .ZN(n14527) );
  OAI211_X1 U15949 ( .C1(n14529), .C2(n14619), .A(n14528), .B(n14527), .ZN(
        n14530) );
  AOI21_X1 U15950 ( .B1(n14669), .B2(n11368), .A(n14530), .ZN(n14531) );
  OAI21_X1 U15951 ( .B1(n14580), .B2(n14673), .A(n14531), .ZN(P2_U3242) );
  XNOR2_X1 U15952 ( .A(n14532), .B(n14541), .ZN(n14534) );
  AOI21_X1 U15953 ( .B1(n14534), .B2(n14606), .A(n14533), .ZN(n14677) );
  NAND2_X1 U15954 ( .A1(n14550), .A2(n14675), .ZN(n14535) );
  NAND2_X1 U15955 ( .A1(n14535), .A2(n14430), .ZN(n14536) );
  NOR2_X1 U15956 ( .A1(n14537), .A2(n14536), .ZN(n14674) );
  NAND2_X1 U15957 ( .A1(n14675), .A2(n14628), .ZN(n14539) );
  NAND2_X1 U15958 ( .A1(n14622), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n14538) );
  OAI211_X1 U15959 ( .C1(n14624), .C2(n14540), .A(n14539), .B(n14538), .ZN(
        n14545) );
  OAI21_X1 U15960 ( .B1(n14543), .B2(n8965), .A(n14542), .ZN(n14678) );
  NOR2_X1 U15961 ( .A1(n14678), .A2(n14580), .ZN(n14544) );
  AOI211_X1 U15962 ( .C1(n14674), .C2(n14632), .A(n14545), .B(n14544), .ZN(
        n14546) );
  OAI21_X1 U15963 ( .B1(n14622), .B2(n14677), .A(n14546), .ZN(P2_U3243) );
  OAI21_X1 U15964 ( .B1(n7513), .B2(n14558), .A(n14547), .ZN(n14549) );
  AOI21_X1 U15965 ( .B1(n14549), .B2(n14606), .A(n14548), .ZN(n14685) );
  OAI211_X1 U15966 ( .C1(n14572), .C2(n14551), .A(n14430), .B(n14550), .ZN(
        n14682) );
  INV_X1 U15967 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n14553) );
  OAI22_X1 U15968 ( .A1(n11368), .A2(n14553), .B1(n14552), .B2(n14624), .ZN(
        n14554) );
  AOI21_X1 U15969 ( .B1(n14681), .B2(n14628), .A(n14554), .ZN(n14555) );
  OAI21_X1 U15970 ( .B1(n14682), .B2(n14556), .A(n14555), .ZN(n14557) );
  INV_X1 U15971 ( .A(n14557), .ZN(n14561) );
  NAND2_X1 U15972 ( .A1(n14559), .A2(n14558), .ZN(n14679) );
  NAND3_X1 U15973 ( .A1(n14680), .A2(n14679), .A3(n14630), .ZN(n14560) );
  OAI211_X1 U15974 ( .C1(n14685), .C2(n14622), .A(n14561), .B(n14560), .ZN(
        P2_U3244) );
  OAI21_X1 U15975 ( .B1(n14564), .B2(n14563), .A(n14562), .ZN(n14565) );
  INV_X1 U15976 ( .A(n14565), .ZN(n14690) );
  NAND2_X1 U15977 ( .A1(n14566), .A2(n14606), .ZN(n14571) );
  AOI21_X1 U15978 ( .B1(n14583), .B2(n14568), .A(n14567), .ZN(n14570) );
  OAI21_X1 U15979 ( .B1(n14571), .B2(n14570), .A(n14569), .ZN(n14686) );
  INV_X1 U15980 ( .A(n14595), .ZN(n14573) );
  AOI211_X1 U15981 ( .C1(n14688), .C2(n14573), .A(n7437), .B(n14572), .ZN(
        n14687) );
  NAND2_X1 U15982 ( .A1(n14687), .A2(n14632), .ZN(n14576) );
  AOI22_X1 U15983 ( .A1(n14622), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14574), 
        .B2(n14615), .ZN(n14575) );
  OAI211_X1 U15984 ( .C1(n14577), .C2(n14619), .A(n14576), .B(n14575), .ZN(
        n14578) );
  AOI21_X1 U15985 ( .B1(n14686), .B2(n11368), .A(n14578), .ZN(n14579) );
  OAI21_X1 U15986 ( .B1(n14580), .B2(n14690), .A(n14579), .ZN(P2_U3245) );
  OAI21_X1 U15987 ( .B1(n14582), .B2(n14586), .A(n14581), .ZN(n14693) );
  INV_X1 U15988 ( .A(n14693), .ZN(n14603) );
  INV_X1 U15989 ( .A(n14583), .ZN(n14584) );
  AOI21_X1 U15990 ( .B1(n14586), .B2(n14585), .A(n14584), .ZN(n14594) );
  AOI22_X1 U15991 ( .A1(n14590), .A2(n14589), .B1(n14588), .B2(n14587), .ZN(
        n14593) );
  NAND2_X1 U15992 ( .A1(n14693), .A2(n14591), .ZN(n14592) );
  OAI211_X1 U15993 ( .C1(n14594), .C2(n9148), .A(n14593), .B(n14592), .ZN(
        n14691) );
  NAND2_X1 U15994 ( .A1(n14691), .A2(n11368), .ZN(n14601) );
  AOI211_X1 U15995 ( .C1(n14596), .C2(n14611), .A(n7437), .B(n14595), .ZN(
        n14692) );
  AOI22_X1 U15996 ( .A1(n14622), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14597), 
        .B2(n14615), .ZN(n14598) );
  OAI21_X1 U15997 ( .B1(n14759), .B2(n14619), .A(n14598), .ZN(n14599) );
  AOI21_X1 U15998 ( .B1(n14692), .B2(n14632), .A(n14599), .ZN(n14600) );
  OAI211_X1 U15999 ( .C1(n14603), .C2(n14602), .A(n14601), .B(n14600), .ZN(
        P2_U3246) );
  XOR2_X1 U16000 ( .A(n14609), .B(n14604), .Z(n14607) );
  AOI21_X1 U16001 ( .B1(n14607), .B2(n14606), .A(n14605), .ZN(n14700) );
  OAI21_X1 U16002 ( .B1(n14610), .B2(n14609), .A(n14608), .ZN(n14696) );
  INV_X1 U16003 ( .A(n14611), .ZN(n14612) );
  AOI211_X1 U16004 ( .C1(n14698), .C2(n14613), .A(n7437), .B(n14612), .ZN(
        n14697) );
  NAND2_X1 U16005 ( .A1(n14697), .A2(n14632), .ZN(n14618) );
  INV_X1 U16006 ( .A(n14614), .ZN(n14616) );
  AOI22_X1 U16007 ( .A1(n14622), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14616), 
        .B2(n14615), .ZN(n14617) );
  OAI211_X1 U16008 ( .C1(n9109), .C2(n14619), .A(n14618), .B(n14617), .ZN(
        n14620) );
  AOI21_X1 U16009 ( .B1(n14630), .B2(n14696), .A(n14620), .ZN(n14621) );
  OAI21_X1 U16010 ( .B1(n14622), .B2(n14700), .A(n14621), .ZN(P2_U3247) );
  NAND2_X1 U16011 ( .A1(n14623), .A2(n11368), .ZN(n14637) );
  OAI22_X1 U16012 ( .A1(n11368), .A2(n14626), .B1(n14625), .B2(n14624), .ZN(
        n14627) );
  AOI21_X1 U16013 ( .B1(n14629), .B2(n14628), .A(n14627), .ZN(n14636) );
  NAND2_X1 U16014 ( .A1(n14631), .A2(n14630), .ZN(n14635) );
  NAND2_X1 U16015 ( .A1(n14633), .A2(n14632), .ZN(n14634) );
  NAND4_X1 U16016 ( .A1(n14637), .A2(n14636), .A3(n14635), .A4(n14634), .ZN(
        P2_U3256) );
  MUX2_X1 U16017 ( .A(n14639), .B(n14729), .S(n16560), .Z(n14640) );
  OAI21_X1 U16018 ( .B1(n14732), .B2(n14715), .A(n14640), .ZN(P2_U3530) );
  INV_X1 U16019 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14643) );
  AND2_X1 U16020 ( .A1(n14642), .A2(n14641), .ZN(n14733) );
  MUX2_X1 U16021 ( .A(n14643), .B(n14733), .S(n16560), .Z(n14644) );
  OAI21_X1 U16022 ( .B1(n14736), .B2(n14715), .A(n14644), .ZN(P2_U3529) );
  INV_X1 U16023 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n14645) );
  NAND2_X1 U16024 ( .A1(n16559), .A2(n14645), .ZN(n14646) );
  AND2_X1 U16025 ( .A1(n14651), .A2(n14650), .ZN(n14652) );
  INV_X1 U16026 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n14657) );
  MUX2_X1 U16027 ( .A(n14657), .B(n14741), .S(n16560), .Z(n14658) );
  OAI21_X1 U16028 ( .B1(n14744), .B2(n14715), .A(n14658), .ZN(P2_U3525) );
  INV_X1 U16029 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14662) );
  AOI211_X1 U16030 ( .C1(n14717), .C2(n14661), .A(n14660), .B(n14659), .ZN(
        n14745) );
  MUX2_X1 U16031 ( .A(n14662), .B(n14745), .S(n16560), .Z(n14663) );
  OAI21_X1 U16032 ( .B1(n14748), .B2(n14715), .A(n14663), .ZN(P2_U3524) );
  INV_X1 U16033 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n14667) );
  AOI211_X1 U16034 ( .C1(n14717), .C2(n14666), .A(n14665), .B(n14664), .ZN(
        n14749) );
  MUX2_X1 U16035 ( .A(n14667), .B(n14749), .S(n16560), .Z(n14668) );
  OAI21_X1 U16036 ( .B1(n7963), .B2(n14715), .A(n14668), .ZN(P2_U3523) );
  AOI211_X1 U16037 ( .C1(n16382), .C2(n14671), .A(n14670), .B(n14669), .ZN(
        n14672) );
  OAI21_X1 U16038 ( .B1(n16386), .B2(n14673), .A(n14672), .ZN(n14752) );
  MUX2_X1 U16039 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14752), .S(n16560), .Z(
        P2_U3522) );
  AOI21_X1 U16040 ( .B1(n16382), .B2(n14675), .A(n14674), .ZN(n14676) );
  OAI211_X1 U16041 ( .C1(n14678), .C2(n16386), .A(n14677), .B(n14676), .ZN(
        n14753) );
  MUX2_X1 U16042 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14753), .S(n16560), .Z(
        P2_U3521) );
  NAND3_X1 U16043 ( .A1(n14680), .A2(n14679), .A3(n14717), .ZN(n14684) );
  NAND2_X1 U16044 ( .A1(n14681), .A2(n16382), .ZN(n14683) );
  NAND4_X1 U16045 ( .A1(n14685), .A2(n14684), .A3(n14683), .A4(n14682), .ZN(
        n14754) );
  MUX2_X1 U16046 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14754), .S(n16560), .Z(
        P2_U3520) );
  AOI211_X1 U16047 ( .C1(n16382), .C2(n14688), .A(n14687), .B(n14686), .ZN(
        n14689) );
  OAI21_X1 U16048 ( .B1(n16386), .B2(n14690), .A(n14689), .ZN(n14755) );
  MUX2_X1 U16049 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14755), .S(n16560), .Z(
        P2_U3519) );
  INV_X1 U16050 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14694) );
  AOI211_X1 U16051 ( .C1(n16558), .C2(n14693), .A(n14692), .B(n14691), .ZN(
        n14756) );
  MUX2_X1 U16052 ( .A(n14694), .B(n14756), .S(n16560), .Z(n14695) );
  OAI21_X1 U16053 ( .B1(n14759), .B2(n14715), .A(n14695), .ZN(P2_U3518) );
  INV_X1 U16054 ( .A(n14696), .ZN(n14701) );
  AOI21_X1 U16055 ( .B1(n16382), .B2(n14698), .A(n14697), .ZN(n14699) );
  OAI211_X1 U16056 ( .C1(n16386), .C2(n14701), .A(n14700), .B(n14699), .ZN(
        n14760) );
  MUX2_X1 U16057 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14760), .S(n16560), .Z(
        P2_U3517) );
  OAI211_X1 U16058 ( .C1(n16386), .C2(n14704), .A(n14703), .B(n14702), .ZN(
        n14761) );
  INV_X1 U16059 ( .A(n14761), .ZN(n14705) );
  MUX2_X1 U16060 ( .A(n14706), .B(n14705), .S(n16560), .Z(n14707) );
  OAI21_X1 U16061 ( .B1(n14708), .B2(n14715), .A(n14707), .ZN(P2_U3516) );
  OAI211_X1 U16062 ( .C1(n16386), .C2(n14711), .A(n14710), .B(n14709), .ZN(
        n14712) );
  INV_X1 U16063 ( .A(n14712), .ZN(n14765) );
  MUX2_X1 U16064 ( .A(n14713), .B(n14765), .S(n16560), .Z(n14714) );
  OAI21_X1 U16065 ( .B1(n14769), .B2(n14715), .A(n14714), .ZN(P2_U3515) );
  INV_X1 U16066 ( .A(n7757), .ZN(n14721) );
  NAND2_X1 U16067 ( .A1(n14718), .A2(n14717), .ZN(n14720) );
  OAI211_X1 U16068 ( .C1(n14721), .C2(n16553), .A(n14720), .B(n14719), .ZN(
        n14722) );
  OR2_X1 U16069 ( .A1(n14723), .A2(n14722), .ZN(n14770) );
  MUX2_X1 U16070 ( .A(n14770), .B(P2_REG1_REG_15__SCAN_IN), .S(n16559), .Z(
        P2_U3514) );
  AOI21_X1 U16071 ( .B1(n16382), .B2(n14725), .A(n14724), .ZN(n14726) );
  OAI211_X1 U16072 ( .C1(n16386), .C2(n14728), .A(n14727), .B(n14726), .ZN(
        n14771) );
  MUX2_X1 U16073 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14771), .S(n16560), .Z(
        P2_U3513) );
  MUX2_X1 U16074 ( .A(n14730), .B(n14729), .S(n11936), .Z(n14731) );
  OAI21_X1 U16075 ( .B1(n14732), .B2(n14768), .A(n14731), .ZN(P2_U3498) );
  MUX2_X1 U16076 ( .A(n14734), .B(n14733), .S(n11936), .Z(n14735) );
  OAI21_X1 U16077 ( .B1(n14736), .B2(n14768), .A(n14735), .ZN(P2_U3497) );
  INV_X1 U16078 ( .A(n14737), .ZN(n14738) );
  MUX2_X1 U16079 ( .A(n14742), .B(n14741), .S(n11936), .Z(n14743) );
  OAI21_X1 U16080 ( .B1(n14744), .B2(n14768), .A(n14743), .ZN(P2_U3493) );
  MUX2_X1 U16081 ( .A(n14746), .B(n14745), .S(n11936), .Z(n14747) );
  OAI21_X1 U16082 ( .B1(n14748), .B2(n14768), .A(n14747), .ZN(P2_U3492) );
  MUX2_X1 U16083 ( .A(n14750), .B(n14749), .S(n11936), .Z(n14751) );
  OAI21_X1 U16084 ( .B1(n7963), .B2(n14768), .A(n14751), .ZN(P2_U3491) );
  MUX2_X1 U16085 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14752), .S(n11936), .Z(
        P2_U3490) );
  MUX2_X1 U16086 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14753), .S(n11936), .Z(
        P2_U3489) );
  MUX2_X1 U16087 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14754), .S(n11936), .Z(
        P2_U3488) );
  MUX2_X1 U16088 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14755), .S(n11936), .Z(
        P2_U3487) );
  INV_X1 U16089 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14757) );
  MUX2_X1 U16090 ( .A(n14757), .B(n14756), .S(n11936), .Z(n14758) );
  OAI21_X1 U16091 ( .B1(n14759), .B2(n14768), .A(n14758), .ZN(P2_U3486) );
  MUX2_X1 U16092 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14760), .S(n11936), .Z(
        P2_U3484) );
  MUX2_X1 U16093 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14761), .S(n11936), .Z(
        n14762) );
  AOI21_X1 U16094 ( .B1(n9744), .B2(n14763), .A(n14762), .ZN(n14764) );
  INV_X1 U16095 ( .A(n14764), .ZN(P2_U3481) );
  MUX2_X1 U16096 ( .A(n14766), .B(n14765), .S(n11936), .Z(n14767) );
  OAI21_X1 U16097 ( .B1(n14769), .B2(n14768), .A(n14767), .ZN(P2_U3478) );
  MUX2_X1 U16098 ( .A(n14770), .B(P2_REG0_REG_15__SCAN_IN), .S(n16561), .Z(
        P2_U3475) );
  MUX2_X1 U16099 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n14771), .S(n11936), .Z(
        P2_U3472) );
  INV_X1 U16100 ( .A(n15207), .ZN(n15765) );
  NOR4_X1 U16101 ( .A1(n14773), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14772), .A4(
        P2_U3088), .ZN(n14774) );
  AOI21_X1 U16102 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n7626), .A(n14774), 
        .ZN(n14775) );
  OAI21_X1 U16103 ( .B1(n15765), .B2(n14783), .A(n14775), .ZN(P2_U3296) );
  INV_X1 U16104 ( .A(n15200), .ZN(n15768) );
  OAI222_X1 U16105 ( .A1(n14783), .A2(n15768), .B1(P2_U3088), .B2(n14776), 
        .C1(n14777), .C2(n14787), .ZN(P2_U3297) );
  INV_X1 U16106 ( .A(n14778), .ZN(n15773) );
  AOI21_X1 U16107 ( .B1(n7626), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14779), 
        .ZN(n14780) );
  OAI21_X1 U16108 ( .B1(n15773), .B2(n14783), .A(n14780), .ZN(P2_U3299) );
  INV_X1 U16109 ( .A(n14781), .ZN(n15775) );
  OAI222_X1 U16110 ( .A1(n14787), .A2(n14784), .B1(n14783), .B2(n15775), .C1(
        n14782), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U16111 ( .A(n14785), .ZN(n14789) );
  INV_X1 U16112 ( .A(n14786), .ZN(n15779) );
  OAI222_X1 U16113 ( .A1(P2_U3088), .A2(n14789), .B1(n14783), .B2(n15779), 
        .C1(n14788), .C2(n14787), .ZN(P2_U3301) );
  INV_X1 U16114 ( .A(n14791), .ZN(n14792) );
  MUX2_X1 U16115 ( .A(n14792), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U16116 ( .A1(n15659), .A2(n14917), .ZN(n14794) );
  NAND2_X1 U16117 ( .A1(n14916), .A2(n15302), .ZN(n14793) );
  NAND2_X1 U16118 ( .A1(n14794), .A2(n14793), .ZN(n14795) );
  XNOR2_X1 U16119 ( .A(n14795), .B(n14919), .ZN(n14911) );
  AOI22_X1 U16120 ( .A1(n15659), .A2(n14916), .B1(n14918), .B2(n15302), .ZN(
        n14912) );
  XNOR2_X1 U16121 ( .A(n14911), .B(n14912), .ZN(n14914) );
  INV_X1 U16122 ( .A(n14798), .ZN(n14799) );
  NAND2_X1 U16123 ( .A1(n14800), .A2(n14799), .ZN(n14801) );
  NAND2_X1 U16124 ( .A1(n16611), .A2(n14917), .ZN(n14803) );
  NAND2_X1 U16125 ( .A1(n14916), .A2(n15315), .ZN(n14802) );
  NAND2_X1 U16126 ( .A1(n14803), .A2(n14802), .ZN(n14804) );
  XNOR2_X1 U16127 ( .A(n14804), .B(n14827), .ZN(n14807) );
  NOR2_X1 U16128 ( .A1(n14830), .A2(n14805), .ZN(n14806) );
  AOI21_X1 U16129 ( .B1(n16611), .B2(n14916), .A(n14806), .ZN(n14808) );
  NAND2_X1 U16130 ( .A1(n14807), .A2(n14808), .ZN(n14812) );
  INV_X1 U16131 ( .A(n14807), .ZN(n14810) );
  INV_X1 U16132 ( .A(n14808), .ZN(n14809) );
  NAND2_X1 U16133 ( .A1(n14810), .A2(n14809), .ZN(n14811) );
  NAND2_X1 U16134 ( .A1(n14812), .A2(n14811), .ZN(n16606) );
  AOI22_X1 U16135 ( .A1(n15732), .A2(n14917), .B1(n14916), .B2(n15314), .ZN(
        n14813) );
  XNOR2_X1 U16136 ( .A(n14813), .B(n14919), .ZN(n14815) );
  AOI22_X1 U16137 ( .A1(n15732), .A2(n14916), .B1(n14918), .B2(n15314), .ZN(
        n15023) );
  NAND2_X1 U16138 ( .A1(n15725), .A2(n14917), .ZN(n14817) );
  NAND2_X1 U16139 ( .A1(n14916), .A2(n15313), .ZN(n14816) );
  NAND2_X1 U16140 ( .A1(n14817), .A2(n14816), .ZN(n14818) );
  XNOR2_X1 U16141 ( .A(n14818), .B(n14827), .ZN(n14822) );
  NOR2_X1 U16142 ( .A1(n14830), .A2(n14819), .ZN(n14820) );
  AOI21_X1 U16143 ( .B1(n15725), .B2(n14916), .A(n14820), .ZN(n14821) );
  NAND2_X1 U16144 ( .A1(n14822), .A2(n14821), .ZN(n14823) );
  OAI21_X1 U16145 ( .B1(n14822), .B2(n14821), .A(n14823), .ZN(n14959) );
  INV_X1 U16146 ( .A(n14823), .ZN(n14824) );
  NAND2_X1 U16147 ( .A1(n15715), .A2(n14917), .ZN(n14826) );
  NAND2_X1 U16148 ( .A1(n14916), .A2(n15312), .ZN(n14825) );
  NAND2_X1 U16149 ( .A1(n14826), .A2(n14825), .ZN(n14828) );
  XNOR2_X1 U16150 ( .A(n14828), .B(n14827), .ZN(n14833) );
  NOR2_X1 U16151 ( .A1(n14830), .A2(n14829), .ZN(n14831) );
  AOI21_X1 U16152 ( .B1(n15715), .B2(n14916), .A(n14831), .ZN(n14832) );
  NOR2_X1 U16153 ( .A1(n14833), .A2(n14832), .ZN(n14968) );
  NAND2_X1 U16154 ( .A1(n14833), .A2(n14832), .ZN(n14966) );
  NAND2_X1 U16155 ( .A1(n15710), .A2(n14917), .ZN(n14835) );
  NAND2_X1 U16156 ( .A1(n15311), .A2(n14916), .ZN(n14834) );
  NAND2_X1 U16157 ( .A1(n14835), .A2(n14834), .ZN(n14836) );
  XNOR2_X1 U16158 ( .A(n14836), .B(n14919), .ZN(n14837) );
  AOI22_X1 U16159 ( .A1(n15710), .A2(n14916), .B1(n14918), .B2(n15311), .ZN(
        n14838) );
  XNOR2_X1 U16160 ( .A(n14837), .B(n14838), .ZN(n15005) );
  INV_X1 U16161 ( .A(n14837), .ZN(n14839) );
  AOI22_X1 U16162 ( .A1(n15703), .A2(n14916), .B1(n14918), .B2(n15310), .ZN(
        n14843) );
  NAND2_X1 U16163 ( .A1(n15703), .A2(n14917), .ZN(n14841) );
  NAND2_X1 U16164 ( .A1(n15310), .A2(n14916), .ZN(n14840) );
  NAND2_X1 U16165 ( .A1(n14841), .A2(n14840), .ZN(n14842) );
  XNOR2_X1 U16166 ( .A(n14842), .B(n14919), .ZN(n14845) );
  XOR2_X1 U16167 ( .A(n14843), .B(n14845), .Z(n14905) );
  INV_X1 U16168 ( .A(n14843), .ZN(n14844) );
  OR2_X1 U16169 ( .A1(n14845), .A2(n14844), .ZN(n14846) );
  OAI21_X2 U16170 ( .B1(n14904), .B2(n14905), .A(n14846), .ZN(n14988) );
  AND2_X1 U16171 ( .A1(n15309), .A2(n14918), .ZN(n14847) );
  AOI21_X1 U16172 ( .B1(n15699), .B2(n14916), .A(n14847), .ZN(n14851) );
  NAND2_X1 U16173 ( .A1(n15699), .A2(n14917), .ZN(n14849) );
  NAND2_X1 U16174 ( .A1(n15309), .A2(n14916), .ZN(n14848) );
  NAND2_X1 U16175 ( .A1(n14849), .A2(n14848), .ZN(n14850) );
  XNOR2_X1 U16176 ( .A(n14850), .B(n14919), .ZN(n14853) );
  XOR2_X1 U16177 ( .A(n14851), .B(n14853), .Z(n14989) );
  INV_X1 U16178 ( .A(n14851), .ZN(n14852) );
  AND2_X1 U16179 ( .A1(n14853), .A2(n14852), .ZN(n14854) );
  NAND2_X1 U16180 ( .A1(n15694), .A2(n14917), .ZN(n14856) );
  NAND2_X1 U16181 ( .A1(n15308), .A2(n14916), .ZN(n14855) );
  NAND2_X1 U16182 ( .A1(n14856), .A2(n14855), .ZN(n14857) );
  XNOR2_X1 U16183 ( .A(n14857), .B(n14919), .ZN(n14860) );
  AOI22_X1 U16184 ( .A1(n15694), .A2(n14916), .B1(n14918), .B2(n15308), .ZN(
        n14858) );
  XNOR2_X1 U16185 ( .A(n14860), .B(n14858), .ZN(n14933) );
  INV_X1 U16186 ( .A(n14858), .ZN(n14859) );
  OR2_X1 U16187 ( .A1(n15688), .A2(n14863), .ZN(n14862) );
  INV_X1 U16188 ( .A(n15146), .ZN(n15307) );
  NAND2_X1 U16189 ( .A1(n15307), .A2(n14918), .ZN(n14861) );
  NAND2_X1 U16190 ( .A1(n14862), .A2(n14861), .ZN(n14865) );
  OAI22_X1 U16191 ( .A1(n15688), .A2(n11208), .B1(n15146), .B2(n14863), .ZN(
        n14864) );
  XNOR2_X1 U16192 ( .A(n14864), .B(n14919), .ZN(n14866) );
  XOR2_X1 U16193 ( .A(n14865), .B(n14866), .Z(n14995) );
  OR2_X1 U16194 ( .A1(n14866), .A2(n14865), .ZN(n14867) );
  NAND2_X1 U16195 ( .A1(n15681), .A2(n14917), .ZN(n14869) );
  NAND2_X1 U16196 ( .A1(n14916), .A2(n15306), .ZN(n14868) );
  NAND2_X1 U16197 ( .A1(n14869), .A2(n14868), .ZN(n14870) );
  XNOR2_X1 U16198 ( .A(n14870), .B(n14919), .ZN(n14871) );
  AOI22_X1 U16199 ( .A1(n15681), .A2(n14916), .B1(n14918), .B2(n15306), .ZN(
        n14872) );
  XNOR2_X1 U16200 ( .A(n14871), .B(n14872), .ZN(n14899) );
  INV_X1 U16201 ( .A(n14871), .ZN(n14873) );
  AOI22_X1 U16202 ( .A1(n15675), .A2(n14916), .B1(n14918), .B2(n15305), .ZN(
        n14877) );
  NAND2_X1 U16203 ( .A1(n15675), .A2(n14917), .ZN(n14875) );
  NAND2_X1 U16204 ( .A1(n14916), .A2(n15305), .ZN(n14874) );
  NAND2_X1 U16205 ( .A1(n14875), .A2(n14874), .ZN(n14876) );
  XNOR2_X1 U16206 ( .A(n14876), .B(n14919), .ZN(n14879) );
  XOR2_X1 U16207 ( .A(n14877), .B(n14879), .Z(n14977) );
  INV_X1 U16208 ( .A(n14877), .ZN(n14878) );
  NAND2_X1 U16209 ( .A1(n15668), .A2(n14917), .ZN(n14881) );
  NAND2_X1 U16210 ( .A1(n14916), .A2(n15304), .ZN(n14880) );
  NAND2_X1 U16211 ( .A1(n14881), .A2(n14880), .ZN(n14882) );
  XNOR2_X1 U16212 ( .A(n14882), .B(n14919), .ZN(n14883) );
  AOI22_X1 U16213 ( .A1(n15668), .A2(n14916), .B1(n14918), .B2(n15304), .ZN(
        n14884) );
  XNOR2_X1 U16214 ( .A(n14883), .B(n14884), .ZN(n14951) );
  INV_X1 U16215 ( .A(n14883), .ZN(n14885) );
  AOI22_X1 U16216 ( .A1(n15664), .A2(n14916), .B1(n14918), .B2(n15303), .ZN(
        n14889) );
  NAND2_X1 U16217 ( .A1(n15664), .A2(n14917), .ZN(n14887) );
  NAND2_X1 U16218 ( .A1(n14916), .A2(n15303), .ZN(n14886) );
  NAND2_X1 U16219 ( .A1(n14887), .A2(n14886), .ZN(n14888) );
  XNOR2_X1 U16220 ( .A(n14888), .B(n14919), .ZN(n14891) );
  XOR2_X1 U16221 ( .A(n14889), .B(n14891), .Z(n15015) );
  INV_X1 U16222 ( .A(n14889), .ZN(n14890) );
  XOR2_X1 U16223 ( .A(n14914), .B(n14915), .Z(n14897) );
  NAND2_X1 U16224 ( .A1(n15008), .A2(n15301), .ZN(n14893) );
  NAND2_X1 U16225 ( .A1(n15006), .A2(n15303), .ZN(n14892) );
  NAND2_X1 U16226 ( .A1(n14893), .A2(n14892), .ZN(n15658) );
  AOI22_X1 U16227 ( .A1(n16614), .A2(n15658), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14894) );
  OAI21_X1 U16228 ( .B1(n15455), .B2(n16619), .A(n14894), .ZN(n14895) );
  AOI21_X1 U16229 ( .B1(n15659), .B2(n16610), .A(n14895), .ZN(n14896) );
  OAI21_X1 U16230 ( .B1(n14897), .B2(n15029), .A(n14896), .ZN(P1_U3214) );
  XOR2_X1 U16231 ( .A(n14899), .B(n14898), .Z(n14903) );
  OAI22_X1 U16232 ( .A1(n15146), .A2(n15293), .B1(n14953), .B2(n15016), .ZN(
        n15680) );
  AOI22_X1 U16233 ( .A1(n15680), .A2(n16614), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14900) );
  OAI21_X1 U16234 ( .B1(n15513), .B2(n16619), .A(n14900), .ZN(n14901) );
  AOI21_X1 U16235 ( .B1(n15681), .B2(n16610), .A(n14901), .ZN(n14902) );
  OAI21_X1 U16236 ( .B1(n14903), .B2(n15029), .A(n14902), .ZN(P1_U3216) );
  XOR2_X1 U16237 ( .A(n14905), .B(n14904), .Z(n14910) );
  NOR2_X1 U16238 ( .A1(n16619), .A2(n15576), .ZN(n14908) );
  AND2_X1 U16239 ( .A1(n15311), .A2(n15006), .ZN(n14906) );
  AOI21_X1 U16240 ( .B1(n15309), .B2(n15008), .A(n14906), .ZN(n15585) );
  NAND2_X1 U16241 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15419)
         );
  OAI21_X1 U16242 ( .B1(n15009), .B2(n15585), .A(n15419), .ZN(n14907) );
  AOI211_X1 U16243 ( .C1(n15703), .C2(n16610), .A(n14908), .B(n14907), .ZN(
        n14909) );
  OAI21_X1 U16244 ( .B1(n14910), .B2(n15029), .A(n14909), .ZN(P1_U3219) );
  INV_X1 U16245 ( .A(n14911), .ZN(n14913) );
  AOI22_X1 U16246 ( .A1(n15651), .A2(n14917), .B1(n14916), .B2(n15301), .ZN(
        n14922) );
  AOI22_X1 U16247 ( .A1(n15651), .A2(n14916), .B1(n14918), .B2(n15301), .ZN(
        n14920) );
  XNOR2_X1 U16248 ( .A(n14920), .B(n14919), .ZN(n14921) );
  XOR2_X1 U16249 ( .A(n14922), .B(n14921), .Z(n14923) );
  XNOR2_X1 U16250 ( .A(n14924), .B(n14923), .ZN(n14930) );
  OR2_X1 U16251 ( .A1(n15192), .A2(n15016), .ZN(n14926) );
  NAND2_X1 U16252 ( .A1(n15006), .A2(n15302), .ZN(n14925) );
  NAND2_X1 U16253 ( .A1(n14926), .A2(n14925), .ZN(n15650) );
  AOI22_X1 U16254 ( .A1(n16614), .A2(n15650), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14927) );
  OAI21_X1 U16255 ( .B1(n15440), .B2(n16619), .A(n14927), .ZN(n14928) );
  AOI21_X1 U16256 ( .B1(n15651), .B2(n16610), .A(n14928), .ZN(n14929) );
  OAI21_X1 U16257 ( .B1(n14930), .B2(n15029), .A(n14929), .ZN(P1_U3220) );
  OAI21_X1 U16258 ( .B1(n14933), .B2(n14932), .A(n14931), .ZN(n14938) );
  NAND2_X1 U16259 ( .A1(n15694), .A2(n16610), .ZN(n14936) );
  OAI22_X1 U16260 ( .A1(n15146), .A2(n15016), .B1(n14934), .B2(n15293), .ZN(
        n15539) );
  AOI22_X1 U16261 ( .A1(n15539), .A2(n16614), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14935) );
  OAI211_X1 U16262 ( .C1(n16619), .C2(n15547), .A(n14936), .B(n14935), .ZN(
        n14937) );
  AOI21_X1 U16263 ( .B1(n14938), .B2(n16612), .A(n14937), .ZN(n14939) );
  INV_X1 U16264 ( .A(n14939), .ZN(P1_U3223) );
  AOI22_X1 U16265 ( .A1(n16614), .A2(n14940), .B1(P1_REG3_REG_12__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14941) );
  OAI21_X1 U16266 ( .B1(n14942), .B2(n16619), .A(n14941), .ZN(n14948) );
  INV_X1 U16267 ( .A(n14943), .ZN(n14944) );
  AOI211_X1 U16268 ( .C1(n14946), .C2(n14945), .A(n15029), .B(n14944), .ZN(
        n14947) );
  AOI211_X1 U16269 ( .C1(n16610), .C2(n15101), .A(n14948), .B(n14947), .ZN(
        n14949) );
  INV_X1 U16270 ( .A(n14949), .ZN(P1_U3224) );
  XOR2_X1 U16271 ( .A(n14951), .B(n14950), .Z(n14957) );
  OAI22_X1 U16272 ( .A1(n14953), .A2(n15293), .B1(n14952), .B2(n15016), .ZN(
        n15480) );
  AOI22_X1 U16273 ( .A1(n16614), .A2(n15480), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14954) );
  OAI21_X1 U16274 ( .B1(n15487), .B2(n16619), .A(n14954), .ZN(n14955) );
  AOI21_X1 U16275 ( .B1(n15668), .B2(n16610), .A(n14955), .ZN(n14956) );
  OAI21_X1 U16276 ( .B1(n14957), .B2(n15029), .A(n14956), .ZN(P1_U3225) );
  AOI21_X1 U16277 ( .B1(n14959), .B2(n14958), .A(n7609), .ZN(n14965) );
  NAND2_X1 U16278 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n15930)
         );
  NAND2_X1 U16279 ( .A1(n15312), .A2(n15008), .ZN(n14961) );
  NAND2_X1 U16280 ( .A1(n15006), .A2(n15314), .ZN(n14960) );
  NAND2_X1 U16281 ( .A1(n14961), .A2(n14960), .ZN(n15724) );
  NAND2_X1 U16282 ( .A1(n16614), .A2(n15724), .ZN(n14962) );
  OAI211_X1 U16283 ( .C1(n16619), .C2(n15634), .A(n15930), .B(n14962), .ZN(
        n14963) );
  AOI21_X1 U16284 ( .B1(n15725), .B2(n16610), .A(n14963), .ZN(n14964) );
  OAI21_X1 U16285 ( .B1(n14965), .B2(n15029), .A(n14964), .ZN(P1_U3226) );
  INV_X1 U16286 ( .A(n14966), .ZN(n14967) );
  NOR2_X1 U16287 ( .A1(n14968), .A2(n14967), .ZN(n14969) );
  XNOR2_X1 U16288 ( .A(n14970), .B(n14969), .ZN(n14975) );
  NOR2_X1 U16289 ( .A1(n16619), .A2(n15616), .ZN(n14973) );
  AND2_X1 U16290 ( .A1(n15313), .A2(n15006), .ZN(n14971) );
  AOI21_X1 U16291 ( .B1(n15311), .B2(n15008), .A(n14971), .ZN(n15716) );
  NAND2_X1 U16292 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n15906)
         );
  OAI21_X1 U16293 ( .B1(n15009), .B2(n15716), .A(n15906), .ZN(n14972) );
  AOI211_X1 U16294 ( .C1(n15715), .C2(n16610), .A(n14973), .B(n14972), .ZN(
        n14974) );
  OAI21_X1 U16295 ( .B1(n14975), .B2(n15029), .A(n14974), .ZN(P1_U3228) );
  XOR2_X1 U16296 ( .A(n14977), .B(n14976), .Z(n14983) );
  NAND2_X1 U16297 ( .A1(n15008), .A2(n15304), .ZN(n14979) );
  NAND2_X1 U16298 ( .A1(n15006), .A2(n15306), .ZN(n14978) );
  NAND2_X1 U16299 ( .A1(n14979), .A2(n14978), .ZN(n15495) );
  AOI22_X1 U16300 ( .A1(n16614), .A2(n15495), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14980) );
  OAI21_X1 U16301 ( .B1(n15502), .B2(n16619), .A(n14980), .ZN(n14981) );
  AOI21_X1 U16302 ( .B1(n15675), .B2(n16610), .A(n14981), .ZN(n14982) );
  OAI21_X1 U16303 ( .B1(n14983), .B2(n15029), .A(n14982), .ZN(P1_U3229) );
  NAND2_X1 U16304 ( .A1(n15308), .A2(n15008), .ZN(n14985) );
  NAND2_X1 U16305 ( .A1(n15310), .A2(n15006), .ZN(n14984) );
  NAND2_X1 U16306 ( .A1(n14985), .A2(n14984), .ZN(n15556) );
  AOI22_X1 U16307 ( .A1(n16614), .A2(n15556), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14986) );
  OAI21_X1 U16308 ( .B1(n15563), .B2(n16619), .A(n14986), .ZN(n14991) );
  AOI211_X1 U16309 ( .C1(n14989), .C2(n14988), .A(n15029), .B(n14987), .ZN(
        n14990) );
  AOI211_X1 U16310 ( .C1(n16610), .C2(n15699), .A(n14991), .B(n14990), .ZN(
        n14992) );
  INV_X1 U16311 ( .A(n14992), .ZN(P1_U3233) );
  OAI21_X1 U16312 ( .B1(n14995), .B2(n14994), .A(n14993), .ZN(n14996) );
  NAND2_X1 U16313 ( .A1(n14996), .A2(n16612), .ZN(n15002) );
  INV_X1 U16314 ( .A(n16619), .ZN(n14999) );
  AOI22_X1 U16315 ( .A1(n15308), .A2(n15006), .B1(n15008), .B2(n15306), .ZN(
        n15686) );
  INV_X1 U16316 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14997) );
  OAI22_X1 U16317 ( .A1(n15009), .A2(n15686), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14997), .ZN(n14998) );
  AOI21_X1 U16318 ( .B1(n15000), .B2(n14999), .A(n14998), .ZN(n15001) );
  OAI211_X1 U16319 ( .C1(n15003), .C2(n15688), .A(n15002), .B(n15001), .ZN(
        P1_U3235) );
  XOR2_X1 U16320 ( .A(n15004), .B(n15005), .Z(n15013) );
  NOR2_X1 U16321 ( .A1(n16619), .A2(n15594), .ZN(n15011) );
  AND2_X1 U16322 ( .A1(n15312), .A2(n15006), .ZN(n15007) );
  AOI21_X1 U16323 ( .B1(n15310), .B2(n15008), .A(n15007), .ZN(n15604) );
  NAND2_X1 U16324 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15916)
         );
  OAI21_X1 U16325 ( .B1(n15009), .B2(n15604), .A(n15916), .ZN(n15010) );
  AOI211_X1 U16326 ( .C1(n15710), .C2(n16610), .A(n15011), .B(n15010), .ZN(
        n15012) );
  OAI21_X1 U16327 ( .B1(n15013), .B2(n15029), .A(n15012), .ZN(P1_U3238) );
  XOR2_X1 U16328 ( .A(n15015), .B(n15014), .Z(n15022) );
  INV_X1 U16329 ( .A(n15302), .ZN(n15017) );
  OAI22_X1 U16330 ( .A1(n15018), .A2(n15293), .B1(n15017), .B2(n15016), .ZN(
        n15465) );
  AOI22_X1 U16331 ( .A1(n16614), .A2(n15465), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15019) );
  OAI21_X1 U16332 ( .B1(n15467), .B2(n16619), .A(n15019), .ZN(n15020) );
  AOI21_X1 U16333 ( .B1(n15664), .B2(n16610), .A(n15020), .ZN(n15021) );
  OAI21_X1 U16334 ( .B1(n15022), .B2(n15029), .A(n15021), .ZN(P1_U3240) );
  XNOR2_X1 U16335 ( .A(n15024), .B(n15023), .ZN(n15030) );
  AOI22_X1 U16336 ( .A1(n16614), .A2(n15731), .B1(P1_REG3_REG_15__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15025) );
  OAI21_X1 U16337 ( .B1(n15026), .B2(n16619), .A(n15025), .ZN(n15027) );
  AOI21_X1 U16338 ( .B1(n15732), .B2(n16610), .A(n15027), .ZN(n15028) );
  OAI21_X1 U16339 ( .B1(n15030), .B2(n15029), .A(n15028), .ZN(P1_U3241) );
  NAND2_X1 U16340 ( .A1(n15213), .A2(n15417), .ZN(n15031) );
  NAND2_X1 U16341 ( .A1(n15034), .A2(n15031), .ZN(n15032) );
  NAND2_X1 U16342 ( .A1(n15032), .A2(n15212), .ZN(n15037) );
  OAI21_X1 U16343 ( .B1(n15218), .B2(n15417), .A(n15033), .ZN(n15035) );
  NAND2_X1 U16344 ( .A1(n15035), .A2(n15034), .ZN(n15036) );
  NAND2_X4 U16345 ( .A1(n15037), .A2(n15036), .ZN(n15211) );
  AOI21_X1 U16346 ( .B1(n15211), .B2(n15326), .A(n16396), .ZN(n15053) );
  AND2_X1 U16347 ( .A1(n15039), .A2(n15038), .ZN(n15040) );
  OAI211_X1 U16348 ( .C1(n15041), .C2(n15040), .A(n15049), .B(n15044), .ZN(
        n15043) );
  NAND4_X1 U16349 ( .A1(n15043), .A2(n15046), .A3(n15042), .A4(n15211), .ZN(
        n15052) );
  INV_X1 U16350 ( .A(n15044), .ZN(n15047) );
  OAI211_X1 U16351 ( .C1(n15047), .C2(n16331), .A(n15046), .B(n15045), .ZN(
        n15050) );
  NAND4_X1 U16352 ( .A1(n15050), .A2(n15065), .A3(n15049), .A4(n15048), .ZN(
        n15051) );
  OAI211_X1 U16353 ( .C1(n15054), .C2(n15053), .A(n15052), .B(n15051), .ZN(
        n15059) );
  MUX2_X1 U16354 ( .A(n15056), .B(n15055), .S(n15211), .Z(n15058) );
  MUX2_X1 U16355 ( .A(n16425), .B(n15325), .S(n15211), .Z(n15057) );
  NAND2_X1 U16356 ( .A1(n15059), .A2(n15058), .ZN(n15060) );
  MUX2_X1 U16357 ( .A(n15324), .B(n16448), .S(n15065), .Z(n15063) );
  MUX2_X1 U16358 ( .A(n15324), .B(n16448), .S(n15211), .Z(n15062) );
  MUX2_X1 U16359 ( .A(n15323), .B(n16465), .S(n15211), .Z(n15069) );
  NAND2_X1 U16360 ( .A1(n15068), .A2(n15069), .ZN(n15067) );
  MUX2_X1 U16361 ( .A(n15323), .B(n16465), .S(n15065), .Z(n15066) );
  NAND2_X1 U16362 ( .A1(n15067), .A2(n15066), .ZN(n15073) );
  INV_X1 U16363 ( .A(n15068), .ZN(n15071) );
  INV_X1 U16364 ( .A(n15069), .ZN(n15070) );
  NAND2_X1 U16365 ( .A1(n15071), .A2(n15070), .ZN(n15072) );
  MUX2_X1 U16366 ( .A(n15322), .B(n15074), .S(n15065), .Z(n15076) );
  MUX2_X1 U16367 ( .A(n15322), .B(n15074), .S(n15211), .Z(n15075) );
  INV_X1 U16368 ( .A(n15076), .ZN(n15077) );
  MUX2_X1 U16369 ( .A(n15321), .B(n15078), .S(n15211), .Z(n15082) );
  NAND2_X1 U16370 ( .A1(n15081), .A2(n15082), .ZN(n15080) );
  MUX2_X1 U16371 ( .A(n15321), .B(n15078), .S(n15065), .Z(n15079) );
  NAND2_X1 U16372 ( .A1(n15080), .A2(n15079), .ZN(n15086) );
  INV_X1 U16373 ( .A(n15081), .ZN(n15084) );
  INV_X1 U16374 ( .A(n15082), .ZN(n15083) );
  NAND2_X1 U16375 ( .A1(n15084), .A2(n15083), .ZN(n15085) );
  MUX2_X1 U16376 ( .A(n15320), .B(n16531), .S(n15065), .Z(n15088) );
  MUX2_X1 U16377 ( .A(n15320), .B(n16531), .S(n15211), .Z(n15087) );
  INV_X1 U16378 ( .A(n15088), .ZN(n15089) );
  MUX2_X1 U16379 ( .A(n15319), .B(n15090), .S(n15211), .Z(n15093) );
  MUX2_X1 U16380 ( .A(n15319), .B(n15090), .S(n15065), .Z(n15091) );
  MUX2_X1 U16381 ( .A(n15318), .B(n16572), .S(n15065), .Z(n15097) );
  MUX2_X1 U16382 ( .A(n15318), .B(n16572), .S(n15211), .Z(n15094) );
  NAND2_X1 U16383 ( .A1(n15095), .A2(n15094), .ZN(n15100) );
  INV_X1 U16384 ( .A(n15096), .ZN(n15098) );
  NAND2_X1 U16385 ( .A1(n15098), .A2(n8469), .ZN(n15099) );
  MUX2_X1 U16386 ( .A(n15317), .B(n15101), .S(n15211), .Z(n15103) );
  MUX2_X1 U16387 ( .A(n15317), .B(n15101), .S(n15065), .Z(n15102) );
  INV_X1 U16388 ( .A(n15103), .ZN(n15104) );
  MUX2_X1 U16389 ( .A(n15316), .B(n15105), .S(n15065), .Z(n15107) );
  MUX2_X1 U16390 ( .A(n15316), .B(n15105), .S(n15211), .Z(n15106) );
  INV_X1 U16391 ( .A(n15107), .ZN(n15108) );
  MUX2_X1 U16392 ( .A(n15315), .B(n16611), .S(n15211), .Z(n15112) );
  NAND2_X1 U16393 ( .A1(n15111), .A2(n15112), .ZN(n15110) );
  MUX2_X1 U16394 ( .A(n15315), .B(n16611), .S(n15065), .Z(n15109) );
  NAND2_X1 U16395 ( .A1(n15110), .A2(n15109), .ZN(n15116) );
  INV_X1 U16396 ( .A(n15111), .ZN(n15114) );
  INV_X1 U16397 ( .A(n15112), .ZN(n15113) );
  NAND2_X1 U16398 ( .A1(n15114), .A2(n15113), .ZN(n15115) );
  MUX2_X1 U16399 ( .A(n15314), .B(n15732), .S(n15065), .Z(n15118) );
  MUX2_X1 U16400 ( .A(n15314), .B(n15732), .S(n15211), .Z(n15117) );
  INV_X1 U16401 ( .A(n15118), .ZN(n15119) );
  MUX2_X1 U16402 ( .A(n15313), .B(n15725), .S(n15211), .Z(n15122) );
  MUX2_X1 U16403 ( .A(n15313), .B(n15725), .S(n15065), .Z(n15120) );
  INV_X1 U16404 ( .A(n15122), .ZN(n15123) );
  MUX2_X1 U16405 ( .A(n15312), .B(n15715), .S(n15065), .Z(n15127) );
  MUX2_X1 U16406 ( .A(n15312), .B(n15715), .S(n15211), .Z(n15124) );
  NAND2_X1 U16407 ( .A1(n15125), .A2(n15124), .ZN(n15130) );
  INV_X1 U16408 ( .A(n15126), .ZN(n15128) );
  NAND2_X1 U16409 ( .A1(n15128), .A2(n8464), .ZN(n15129) );
  NAND2_X1 U16410 ( .A1(n15130), .A2(n15129), .ZN(n15132) );
  MUX2_X1 U16411 ( .A(n15311), .B(n15710), .S(n15211), .Z(n15133) );
  MUX2_X1 U16412 ( .A(n15311), .B(n15710), .S(n15065), .Z(n15131) );
  INV_X1 U16413 ( .A(n15133), .ZN(n15134) );
  MUX2_X1 U16414 ( .A(n15310), .B(n15703), .S(n15065), .Z(n15136) );
  MUX2_X1 U16415 ( .A(n15310), .B(n15703), .S(n15211), .Z(n15135) );
  INV_X1 U16416 ( .A(n15136), .ZN(n15137) );
  MUX2_X1 U16417 ( .A(n15309), .B(n15699), .S(n15211), .Z(n15141) );
  NAND2_X1 U16418 ( .A1(n15140), .A2(n15141), .ZN(n15139) );
  MUX2_X1 U16419 ( .A(n15309), .B(n15699), .S(n15065), .Z(n15138) );
  INV_X1 U16420 ( .A(n15140), .ZN(n15143) );
  INV_X1 U16421 ( .A(n15141), .ZN(n15142) );
  MUX2_X1 U16422 ( .A(n15308), .B(n15694), .S(n15065), .Z(n15160) );
  AOI21_X1 U16423 ( .B1(n15160), .B2(n15307), .A(n8506), .ZN(n15150) );
  NAND2_X1 U16424 ( .A1(n15307), .A2(n15211), .ZN(n15154) );
  OR2_X1 U16425 ( .A1(n15694), .A2(n15154), .ZN(n15145) );
  NAND2_X1 U16426 ( .A1(n8506), .A2(n15146), .ZN(n15144) );
  AND2_X1 U16427 ( .A1(n15145), .A2(n15144), .ZN(n15156) );
  NAND2_X1 U16428 ( .A1(n15160), .A2(n15146), .ZN(n15147) );
  OR2_X1 U16429 ( .A1(n15694), .A2(n15065), .ZN(n15152) );
  NAND2_X1 U16430 ( .A1(n15147), .A2(n15152), .ZN(n15148) );
  NAND2_X1 U16431 ( .A1(n15688), .A2(n15148), .ZN(n15149) );
  OAI211_X1 U16432 ( .C1(n15150), .C2(n15688), .A(n15156), .B(n15149), .ZN(
        n15151) );
  INV_X1 U16433 ( .A(n15152), .ZN(n15153) );
  NAND2_X1 U16434 ( .A1(n15160), .A2(n15153), .ZN(n15155) );
  NAND2_X1 U16435 ( .A1(n15155), .A2(n15154), .ZN(n15158) );
  INV_X1 U16436 ( .A(n15156), .ZN(n15157) );
  AOI22_X1 U16437 ( .A1(n15688), .A2(n15158), .B1(n15160), .B2(n15157), .ZN(
        n15162) );
  NOR2_X1 U16438 ( .A1(n15307), .A2(n15211), .ZN(n15159) );
  AOI21_X1 U16439 ( .B1(n15160), .B2(n8506), .A(n15159), .ZN(n15161) );
  MUX2_X1 U16440 ( .A(n15306), .B(n15681), .S(n15065), .Z(n15166) );
  MUX2_X1 U16441 ( .A(n15306), .B(n15681), .S(n15211), .Z(n15164) );
  INV_X1 U16442 ( .A(n15166), .ZN(n15167) );
  MUX2_X1 U16443 ( .A(n15305), .B(n15675), .S(n15211), .Z(n15171) );
  MUX2_X1 U16444 ( .A(n15305), .B(n15675), .S(n15065), .Z(n15168) );
  NAND2_X1 U16445 ( .A1(n15169), .A2(n15168), .ZN(n15175) );
  INV_X1 U16446 ( .A(n15170), .ZN(n15173) );
  INV_X1 U16447 ( .A(n15171), .ZN(n15172) );
  NAND2_X1 U16448 ( .A1(n15173), .A2(n15172), .ZN(n15174) );
  MUX2_X1 U16449 ( .A(n15304), .B(n15668), .S(n15065), .Z(n15177) );
  MUX2_X1 U16450 ( .A(n15304), .B(n15668), .S(n15211), .Z(n15176) );
  MUX2_X1 U16451 ( .A(n15303), .B(n15664), .S(n15211), .Z(n15181) );
  MUX2_X1 U16452 ( .A(n15303), .B(n15664), .S(n15065), .Z(n15179) );
  MUX2_X1 U16453 ( .A(n15302), .B(n15659), .S(n15065), .Z(n15183) );
  MUX2_X1 U16454 ( .A(n15302), .B(n15659), .S(n15211), .Z(n15182) );
  INV_X1 U16455 ( .A(n15183), .ZN(n15184) );
  MUX2_X1 U16456 ( .A(n15301), .B(n15651), .S(n15211), .Z(n15186) );
  NAND2_X1 U16457 ( .A1(n15185), .A2(n15186), .ZN(n15190) );
  MUX2_X1 U16458 ( .A(n15651), .B(n15301), .S(n15211), .Z(n15189) );
  INV_X1 U16459 ( .A(n15185), .ZN(n15188) );
  INV_X1 U16460 ( .A(n15186), .ZN(n15187) );
  MUX2_X1 U16461 ( .A(n15192), .B(n15191), .S(n15211), .Z(n15220) );
  INV_X1 U16462 ( .A(n15192), .ZN(n15300) );
  MUX2_X1 U16463 ( .A(n15300), .B(n15193), .S(n15065), .Z(n15219) );
  INV_X1 U16464 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n15194) );
  NOR2_X1 U16465 ( .A1(n7778), .A2(n15194), .ZN(n15199) );
  INV_X1 U16466 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n15423) );
  NOR2_X1 U16467 ( .A1(n9477), .A2(n15423), .ZN(n15198) );
  INV_X1 U16468 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n15196) );
  NOR2_X1 U16469 ( .A1(n9634), .A2(n15196), .ZN(n15197) );
  OR3_X1 U16470 ( .A1(n15199), .A2(n15198), .A3(n15197), .ZN(n15424) );
  OAI21_X1 U16471 ( .B1(n15424), .B2(n15212), .A(n15299), .ZN(n15203) );
  NAND2_X1 U16472 ( .A1(n15200), .A2(n15206), .ZN(n15202) );
  NAND2_X1 U16473 ( .A1(n7460), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n15201) );
  MUX2_X1 U16474 ( .A(n15203), .B(n15648), .S(n15065), .Z(n15224) );
  OAI21_X1 U16475 ( .B1(n15424), .B2(n15218), .A(n15299), .ZN(n15204) );
  INV_X1 U16476 ( .A(n15204), .ZN(n15205) );
  MUX2_X1 U16477 ( .A(n15205), .B(n15232), .S(n15211), .Z(n15223) );
  NAND2_X1 U16478 ( .A1(n15224), .A2(n15223), .ZN(n15283) );
  OAI21_X1 U16479 ( .B1(n15220), .B2(n15219), .A(n15283), .ZN(n15230) );
  NAND2_X1 U16480 ( .A1(n15207), .A2(n15206), .ZN(n15209) );
  NAND2_X1 U16481 ( .A1(n7459), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n15208) );
  INV_X1 U16482 ( .A(n15424), .ZN(n15210) );
  NOR2_X1 U16483 ( .A1(n15065), .A2(n15210), .ZN(n15267) );
  NAND2_X1 U16484 ( .A1(n15645), .A2(n15267), .ZN(n15263) );
  NOR2_X1 U16485 ( .A1(n15211), .A2(n15424), .ZN(n15271) );
  NAND2_X1 U16486 ( .A1(n15427), .A2(n15271), .ZN(n15262) );
  NAND2_X1 U16487 ( .A1(n15213), .A2(n15212), .ZN(n15214) );
  NAND2_X1 U16488 ( .A1(n15033), .A2(n15214), .ZN(n15216) );
  NAND2_X1 U16489 ( .A1(n15216), .A2(n15215), .ZN(n15272) );
  NAND2_X1 U16490 ( .A1(n15218), .A2(n15217), .ZN(n15280) );
  NAND4_X1 U16491 ( .A1(n15263), .A2(n15262), .A3(n15272), .A4(n15280), .ZN(
        n15282) );
  NOR3_X1 U16492 ( .A1(n15229), .A2(n15230), .A3(n15282), .ZN(n15292) );
  INV_X1 U16493 ( .A(n15219), .ZN(n15222) );
  INV_X1 U16494 ( .A(n15220), .ZN(n15221) );
  NOR2_X1 U16495 ( .A1(n15222), .A2(n15221), .ZN(n15284) );
  INV_X1 U16496 ( .A(n15284), .ZN(n15228) );
  INV_X1 U16497 ( .A(n15272), .ZN(n15270) );
  INV_X1 U16498 ( .A(n15223), .ZN(n15226) );
  INV_X1 U16499 ( .A(n15224), .ZN(n15225) );
  NAND2_X1 U16500 ( .A1(n15226), .A2(n15225), .ZN(n15264) );
  NAND3_X1 U16501 ( .A1(n15231), .A2(n15270), .A3(n15264), .ZN(n15288) );
  INV_X1 U16502 ( .A(n15288), .ZN(n15227) );
  INV_X1 U16503 ( .A(n15230), .ZN(n15289) );
  NOR3_X1 U16504 ( .A1(n15234), .A2(n15233), .A3(n16306), .ZN(n15237) );
  NAND3_X1 U16505 ( .A1(n15237), .A2(n15236), .A3(n15235), .ZN(n15239) );
  NOR4_X1 U16506 ( .A1(n16477), .A2(n16434), .A3(n15239), .A4(n15238), .ZN(
        n15242) );
  NAND4_X1 U16507 ( .A1(n15243), .A2(n15242), .A3(n15241), .A4(n15240), .ZN(
        n15244) );
  NOR4_X1 U16508 ( .A1(n15247), .A2(n15246), .A3(n15245), .A4(n15244), .ZN(
        n15250) );
  NAND4_X1 U16509 ( .A1(n15625), .A2(n15250), .A3(n15249), .A4(n15248), .ZN(
        n15251) );
  NOR4_X1 U16510 ( .A1(n15580), .A2(n15601), .A3(n15611), .A4(n15251), .ZN(
        n15253) );
  NAND4_X1 U16511 ( .A1(n15524), .A2(n15253), .A3(n15252), .A4(n15559), .ZN(
        n15254) );
  NOR4_X1 U16512 ( .A1(n15483), .A2(n15498), .A3(n15255), .A4(n15254), .ZN(
        n15257) );
  NAND4_X1 U16513 ( .A1(n15258), .A2(n15257), .A3(n15256), .A4(n15463), .ZN(
        n15259) );
  XNOR2_X1 U16514 ( .A(n15261), .B(n15417), .ZN(n15281) );
  INV_X1 U16515 ( .A(n15262), .ZN(n15266) );
  INV_X1 U16516 ( .A(n15263), .ZN(n15265) );
  NOR4_X1 U16517 ( .A1(n15266), .A2(n15265), .A3(n15264), .A4(n15270), .ZN(
        n15279) );
  NAND2_X1 U16518 ( .A1(n15424), .A2(n15272), .ZN(n15269) );
  INV_X1 U16519 ( .A(n15267), .ZN(n15268) );
  MUX2_X1 U16520 ( .A(n15272), .B(n15269), .S(n15268), .Z(n15277) );
  NOR3_X1 U16521 ( .A1(n15271), .A2(n15270), .A3(n15424), .ZN(n15275) );
  INV_X1 U16522 ( .A(n15271), .ZN(n15273) );
  NOR2_X1 U16523 ( .A1(n15273), .A2(n15272), .ZN(n15274) );
  OAI21_X1 U16524 ( .B1(n15275), .B2(n15274), .A(n15427), .ZN(n15276) );
  OAI211_X1 U16525 ( .C1(n15277), .C2(n15427), .A(n15276), .B(n15280), .ZN(
        n15278) );
  OAI22_X1 U16526 ( .A1(n15281), .A2(n15280), .B1(n15279), .B2(n15278), .ZN(
        n15287) );
  INV_X1 U16527 ( .A(n15282), .ZN(n15285) );
  NAND3_X1 U16528 ( .A1(n15285), .A2(n15284), .A3(n15283), .ZN(n15286) );
  OAI211_X1 U16529 ( .C1(n15289), .C2(n15288), .A(n15287), .B(n15286), .ZN(
        n15290) );
  NOR3_X1 U16530 ( .A1(n15292), .A2(n15291), .A3(n15290), .ZN(n15298) );
  NOR3_X1 U16531 ( .A1(n15294), .A2(n15885), .A3(n15293), .ZN(n15296) );
  OAI21_X1 U16532 ( .B1(n15297), .B2(n15783), .A(P1_B_REG_SCAN_IN), .ZN(n15295) );
  OAI22_X1 U16533 ( .A1(n15298), .A2(n15297), .B1(n15296), .B2(n15295), .ZN(
        P1_U3242) );
  MUX2_X1 U16534 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n15424), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16535 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n15299), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16536 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n15300), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16537 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n15301), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16538 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n15302), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16539 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n15303), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16540 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n15304), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16541 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n15305), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16542 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n15306), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16543 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n15307), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16544 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n15308), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16545 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n15309), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16546 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n15310), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16547 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15311), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16548 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n15312), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16549 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n15313), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16550 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n15314), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16551 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n15315), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16552 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n15316), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16553 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n15317), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16554 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n15318), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16555 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n15319), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16556 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n15320), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16557 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n15321), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16558 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n15322), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16559 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n15323), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16560 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n15324), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16561 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n15325), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16562 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n15326), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16563 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9639), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16564 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9636), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16565 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n15327), .S(P1_U4016), .Z(
        P1_U3560) );
  NAND2_X1 U16566 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n15343) );
  INV_X1 U16567 ( .A(n15343), .ZN(n15331) );
  MUX2_X1 U16568 ( .A(n9255), .B(P1_REG2_REG_1__SCAN_IN), .S(n15336), .Z(
        n15330) );
  INV_X1 U16569 ( .A(n15328), .ZN(n15329) );
  OAI211_X1 U16570 ( .C1(n15331), .C2(n15330), .A(n15415), .B(n15329), .ZN(
        n15342) );
  INV_X1 U16571 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n15333) );
  OAI22_X1 U16572 ( .A1(n16301), .A2(n15333), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15332), .ZN(n15334) );
  AOI21_X1 U16573 ( .B1(n16287), .B2(n15335), .A(n15334), .ZN(n15341) );
  MUX2_X1 U16574 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10587), .S(n15336), .Z(
        n15337) );
  OAI21_X1 U16575 ( .B1(n9246), .B2(n15887), .A(n15337), .ZN(n15338) );
  NAND3_X1 U16576 ( .A1(n16294), .A2(n15339), .A3(n15338), .ZN(n15340) );
  NAND3_X1 U16577 ( .A1(n15342), .A2(n15341), .A3(n15340), .ZN(P1_U3244) );
  MUX2_X1 U16578 ( .A(n15344), .B(n15343), .S(n15345), .Z(n15349) );
  NAND2_X1 U16579 ( .A1(n15345), .A2(n11580), .ZN(n15346) );
  NAND2_X1 U16580 ( .A1(n15347), .A2(n15346), .ZN(n15884) );
  NAND2_X1 U16581 ( .A1(n15884), .A2(n15887), .ZN(n15890) );
  AND2_X1 U16582 ( .A1(P1_U4016), .A2(n15890), .ZN(n15348) );
  OAI21_X1 U16583 ( .B1(n15349), .B2(n15772), .A(n15348), .ZN(n16297) );
  OAI22_X1 U16584 ( .A1(n16301), .A2(n15950), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11992), .ZN(n15350) );
  AOI21_X1 U16585 ( .B1(n16287), .B2(n15351), .A(n15350), .ZN(n15361) );
  OAI211_X1 U16586 ( .C1(n15353), .C2(n15352), .A(n16294), .B(n15366), .ZN(
        n15360) );
  MUX2_X1 U16587 ( .A(n15355), .B(P1_REG2_REG_2__SCAN_IN), .S(n15354), .Z(
        n15358) );
  INV_X1 U16588 ( .A(n15356), .ZN(n15357) );
  OAI211_X1 U16589 ( .C1(n15358), .C2(n15357), .A(n15415), .B(n15371), .ZN(
        n15359) );
  NAND4_X1 U16590 ( .A1(n16297), .A2(n15361), .A3(n15360), .A4(n15359), .ZN(
        P1_U3245) );
  AND2_X1 U16591 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n16397) );
  NOR2_X1 U16592 ( .A1(n15928), .A2(n15362), .ZN(n15363) );
  AOI211_X1 U16593 ( .C1(n15892), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n16397), .B(
        n15363), .ZN(n15376) );
  MUX2_X1 U16594 ( .A(n10592), .B(P1_REG1_REG_3__SCAN_IN), .S(n15364), .Z(
        n15367) );
  NAND3_X1 U16595 ( .A1(n15367), .A2(n15366), .A3(n15365), .ZN(n15368) );
  NAND3_X1 U16596 ( .A1(n16294), .A2(n16291), .A3(n15368), .ZN(n15375) );
  INV_X1 U16597 ( .A(n16282), .ZN(n15373) );
  NAND3_X1 U16598 ( .A1(n15371), .A2(n15370), .A3(n15369), .ZN(n15372) );
  NAND3_X1 U16599 ( .A1(n15415), .A2(n15373), .A3(n15372), .ZN(n15374) );
  NAND3_X1 U16600 ( .A1(n15376), .A2(n15375), .A3(n15374), .ZN(P1_U3246) );
  INV_X1 U16601 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n15996) );
  OAI21_X1 U16602 ( .B1(n16301), .B2(n15996), .A(n15377), .ZN(n15378) );
  AOI21_X1 U16603 ( .B1(n16287), .B2(n15385), .A(n15378), .ZN(n15393) );
  INV_X1 U16604 ( .A(n15379), .ZN(n15384) );
  NAND3_X1 U16605 ( .A1(n15382), .A2(n15381), .A3(n15380), .ZN(n15383) );
  NAND3_X1 U16606 ( .A1(n15415), .A2(n15384), .A3(n15383), .ZN(n15392) );
  MUX2_X1 U16607 ( .A(n10602), .B(P1_REG1_REG_7__SCAN_IN), .S(n15385), .Z(
        n15386) );
  NAND3_X1 U16608 ( .A1(n15388), .A2(n15387), .A3(n15386), .ZN(n15389) );
  NAND3_X1 U16609 ( .A1(n16294), .A2(n15390), .A3(n15389), .ZN(n15391) );
  NAND3_X1 U16610 ( .A1(n15393), .A2(n15392), .A3(n15391), .ZN(P1_U3250) );
  AOI22_X1 U16611 ( .A1(n15403), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n15398), 
        .B2(n15904), .ZN(n15901) );
  AOI22_X1 U16612 ( .A1(n15407), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n15397), 
        .B2(n15927), .ZN(n15923) );
  NOR2_X1 U16613 ( .A1(n15404), .A2(n15394), .ZN(n15396) );
  NOR2_X1 U16614 ( .A1(n15396), .A2(n15395), .ZN(n15922) );
  NAND2_X1 U16615 ( .A1(n15923), .A2(n15922), .ZN(n15921) );
  OAI21_X1 U16616 ( .B1(n15397), .B2(n15927), .A(n15921), .ZN(n15900) );
  NAND2_X1 U16617 ( .A1(n15901), .A2(n15900), .ZN(n15899) );
  OAI21_X1 U16618 ( .B1(n15398), .B2(n15904), .A(n15899), .ZN(n15399) );
  XNOR2_X1 U16619 ( .A(n15914), .B(n15399), .ZN(n15911) );
  NAND2_X1 U16620 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n15911), .ZN(n15910) );
  NAND2_X1 U16621 ( .A1(n15410), .A2(n15399), .ZN(n15400) );
  NAND2_X1 U16622 ( .A1(n15910), .A2(n15400), .ZN(n15402) );
  XNOR2_X1 U16623 ( .A(n15402), .B(n15401), .ZN(n15416) );
  INV_X1 U16624 ( .A(n15416), .ZN(n15413) );
  AOI22_X1 U16625 ( .A1(n15403), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n15615), 
        .B2(n15904), .ZN(n15898) );
  NAND2_X1 U16626 ( .A1(n15407), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n15408) );
  NOR2_X1 U16627 ( .A1(n15404), .A2(n7502), .ZN(n15406) );
  AOI22_X1 U16628 ( .A1(n15407), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9476), 
        .B2(n15927), .ZN(n15919) );
  NAND2_X1 U16629 ( .A1(n15920), .A2(n15919), .ZN(n15918) );
  NAND2_X1 U16630 ( .A1(n15408), .A2(n15918), .ZN(n15897) );
  NAND2_X1 U16631 ( .A1(n15898), .A2(n15897), .ZN(n15896) );
  OAI21_X1 U16632 ( .B1(n15615), .B2(n15904), .A(n15896), .ZN(n15409) );
  XNOR2_X1 U16633 ( .A(n15914), .B(n15409), .ZN(n15909) );
  NAND2_X1 U16634 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n15909), .ZN(n15908) );
  NAND2_X1 U16635 ( .A1(n15410), .A2(n15409), .ZN(n15411) );
  NOR2_X1 U16636 ( .A1(n15414), .A2(n16285), .ZN(n15412) );
  AOI22_X1 U16637 ( .A1(n15416), .A2(n16294), .B1(n15415), .B2(n15414), .ZN(
        n15418) );
  OAI211_X1 U16638 ( .C1(n15421), .C2(n16301), .A(n15420), .B(n15419), .ZN(
        P1_U3262) );
  XNOR2_X1 U16639 ( .A(n15645), .B(n15429), .ZN(n15422) );
  NAND2_X1 U16640 ( .A1(n15422), .A2(n16473), .ZN(n15644) );
  NOR2_X1 U16641 ( .A1(n15515), .A2(n15423), .ZN(n15426) );
  NAND2_X1 U16642 ( .A1(n15425), .A2(n15424), .ZN(n15646) );
  NOR2_X1 U16643 ( .A1(n16522), .A2(n15646), .ZN(n15431) );
  AOI211_X1 U16644 ( .C1(n15427), .C2(n15619), .A(n15426), .B(n15431), .ZN(
        n15428) );
  OAI21_X1 U16645 ( .B1(n15644), .B2(n15621), .A(n15428), .ZN(P1_U3263) );
  OAI211_X1 U16646 ( .C1(n15648), .C2(n15430), .A(n16473), .B(n15429), .ZN(
        n15647) );
  NAND2_X1 U16647 ( .A1(n16522), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n15433) );
  INV_X1 U16648 ( .A(n15431), .ZN(n15432) );
  OAI211_X1 U16649 ( .C1(n15648), .C2(n16512), .A(n15433), .B(n15432), .ZN(
        n15434) );
  INV_X1 U16650 ( .A(n15434), .ZN(n15435) );
  OAI21_X1 U16651 ( .B1(n15647), .B2(n15621), .A(n15435), .ZN(P1_U3264) );
  XNOR2_X1 U16652 ( .A(n15436), .B(n15445), .ZN(n15655) );
  INV_X1 U16653 ( .A(n15537), .ZN(n15643) );
  NAND2_X1 U16654 ( .A1(n15453), .A2(n15651), .ZN(n15437) );
  NAND2_X1 U16655 ( .A1(n15437), .A2(n16473), .ZN(n15438) );
  NOR2_X1 U16656 ( .A1(n15439), .A2(n15438), .ZN(n15649) );
  INV_X1 U16657 ( .A(n15650), .ZN(n15441) );
  OAI22_X1 U16658 ( .A1(n16522), .A2(n15441), .B1(n15440), .B2(n16490), .ZN(
        n15442) );
  AOI21_X1 U16659 ( .B1(P1_REG2_REG_28__SCAN_IN), .B2(n16522), .A(n15442), 
        .ZN(n15443) );
  OAI21_X1 U16660 ( .B1(n8114), .B2(n16512), .A(n15443), .ZN(n15444) );
  AOI21_X1 U16661 ( .B1(n15649), .B2(n16518), .A(n15444), .ZN(n15449) );
  INV_X1 U16662 ( .A(n15592), .ZN(n15641) );
  NAND3_X1 U16663 ( .A1(n15652), .A2(n15641), .A3(n15447), .ZN(n15448) );
  OAI211_X1 U16664 ( .C1(n15655), .C2(n15643), .A(n15449), .B(n15448), .ZN(
        P1_U3265) );
  XNOR2_X1 U16665 ( .A(n15450), .B(n15451), .ZN(n15662) );
  XNOR2_X1 U16666 ( .A(n15452), .B(n15451), .ZN(n15656) );
  INV_X1 U16667 ( .A(n15453), .ZN(n15454) );
  AOI211_X1 U16668 ( .C1(n15659), .C2(n15470), .A(n16437), .B(n15454), .ZN(
        n15657) );
  NAND2_X1 U16669 ( .A1(n15657), .A2(n16518), .ZN(n15459) );
  INV_X1 U16670 ( .A(n15658), .ZN(n15456) );
  OAI22_X1 U16671 ( .A1(n16522), .A2(n15456), .B1(n15455), .B2(n16490), .ZN(
        n15457) );
  AOI21_X1 U16672 ( .B1(P1_REG2_REG_27__SCAN_IN), .B2(n16522), .A(n15457), 
        .ZN(n15458) );
  OAI211_X1 U16673 ( .C1(n15460), .C2(n16512), .A(n15459), .B(n15458), .ZN(
        n15461) );
  AOI21_X1 U16674 ( .B1(n15656), .B2(n15537), .A(n15461), .ZN(n15462) );
  OAI21_X1 U16675 ( .B1(n15662), .B2(n15608), .A(n15462), .ZN(P1_U3266) );
  XNOR2_X1 U16676 ( .A(n15464), .B(n15463), .ZN(n15466) );
  OAI21_X1 U16677 ( .B1(n15467), .B2(n16490), .A(n15666), .ZN(n15475) );
  OAI21_X1 U16678 ( .B1(n15469), .B2(n8413), .A(n15468), .ZN(n15667) );
  AOI22_X1 U16679 ( .A1(n15664), .A2(n15619), .B1(n16522), .B2(
        P1_REG2_REG_26__SCAN_IN), .ZN(n15473) );
  AOI21_X1 U16680 ( .B1(n15482), .B2(n15664), .A(n16437), .ZN(n15471) );
  NAND2_X1 U16681 ( .A1(n15663), .A2(n16518), .ZN(n15472) );
  OAI211_X1 U16682 ( .C1(n15667), .C2(n15592), .A(n15473), .B(n15472), .ZN(
        n15474) );
  AOI21_X1 U16683 ( .B1(n15475), .B2(n15515), .A(n15474), .ZN(n15476) );
  INV_X1 U16684 ( .A(n15476), .ZN(P1_U3267) );
  OAI21_X1 U16685 ( .B1(n15479), .B2(n15478), .A(n15477), .ZN(n15481) );
  AOI21_X1 U16686 ( .B1(n15481), .B2(n16536), .A(n15480), .ZN(n15673) );
  OAI211_X1 U16687 ( .C1(n7491), .C2(n8102), .A(n16473), .B(n15482), .ZN(
        n15670) );
  OR2_X1 U16688 ( .A1(n15484), .A2(n15483), .ZN(n15669) );
  NAND3_X1 U16689 ( .A1(n15669), .A2(n15641), .A3(n15485), .ZN(n15490) );
  NAND2_X1 U16690 ( .A1(n16522), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n15486) );
  OAI21_X1 U16691 ( .B1(n16490), .B2(n15487), .A(n15486), .ZN(n15488) );
  AOI21_X1 U16692 ( .B1(n15668), .B2(n15619), .A(n15488), .ZN(n15489) );
  OAI211_X1 U16693 ( .C1(n15670), .C2(n15621), .A(n15490), .B(n15489), .ZN(
        n15491) );
  INV_X1 U16694 ( .A(n15491), .ZN(n15492) );
  OAI21_X1 U16695 ( .B1(n15673), .B2(n16522), .A(n15492), .ZN(P1_U3268) );
  AOI211_X1 U16696 ( .C1(n15498), .C2(n15494), .A(n16479), .B(n15493), .ZN(
        n15496) );
  NOR2_X1 U16697 ( .A1(n15496), .A2(n15495), .ZN(n15677) );
  OAI21_X1 U16698 ( .B1(n15499), .B2(n15498), .A(n15497), .ZN(n15500) );
  INV_X1 U16699 ( .A(n15500), .ZN(n15678) );
  NAND2_X1 U16700 ( .A1(n16522), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n15501) );
  OAI21_X1 U16701 ( .B1(n16490), .B2(n15502), .A(n15501), .ZN(n15503) );
  AOI21_X1 U16702 ( .B1(n15675), .B2(n15619), .A(n15503), .ZN(n15507) );
  NAND2_X1 U16703 ( .A1(n15511), .A2(n15675), .ZN(n15504) );
  NAND2_X1 U16704 ( .A1(n15504), .A2(n16473), .ZN(n15505) );
  NOR2_X1 U16705 ( .A1(n7491), .A2(n15505), .ZN(n15674) );
  NAND2_X1 U16706 ( .A1(n15674), .A2(n16518), .ZN(n15506) );
  OAI211_X1 U16707 ( .C1(n15678), .C2(n15608), .A(n15507), .B(n15506), .ZN(
        n15508) );
  INV_X1 U16708 ( .A(n15508), .ZN(n15509) );
  OAI21_X1 U16709 ( .B1(n15677), .B2(n16522), .A(n15509), .ZN(P1_U3269) );
  XNOR2_X1 U16710 ( .A(n15510), .B(n8442), .ZN(n15685) );
  AOI21_X1 U16711 ( .B1(n15681), .B2(n15530), .A(n16437), .ZN(n15512) );
  AND2_X1 U16712 ( .A1(n15512), .A2(n15511), .ZN(n15679) );
  NAND2_X1 U16713 ( .A1(n15681), .A2(n15619), .ZN(n15518) );
  NOR2_X1 U16714 ( .A1(n16490), .A2(n15513), .ZN(n15514) );
  AOI21_X1 U16715 ( .B1(n15680), .B2(n15515), .A(n15514), .ZN(n15517) );
  NAND2_X1 U16716 ( .A1(n16522), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n15516) );
  NAND3_X1 U16717 ( .A1(n15518), .A2(n15517), .A3(n15516), .ZN(n15519) );
  AOI21_X1 U16718 ( .B1(n15679), .B2(n16518), .A(n15519), .ZN(n15523) );
  NAND2_X1 U16719 ( .A1(n15521), .A2(n8442), .ZN(n15682) );
  NAND3_X1 U16720 ( .A1(n15520), .A2(n15682), .A3(n15641), .ZN(n15522) );
  OAI211_X1 U16721 ( .C1(n15685), .C2(n15643), .A(n15523), .B(n15522), .ZN(
        P1_U3270) );
  XNOR2_X1 U16722 ( .A(n15525), .B(n15524), .ZN(n15692) );
  AOI21_X1 U16723 ( .B1(n15528), .B2(n15527), .A(n7781), .ZN(n15529) );
  INV_X1 U16724 ( .A(n15529), .ZN(n15690) );
  OAI211_X1 U16725 ( .C1(n15531), .C2(n15688), .A(n15530), .B(n16473), .ZN(
        n15687) );
  OAI22_X1 U16726 ( .A1(n15686), .A2(n16522), .B1(n15532), .B2(n16490), .ZN(
        n15534) );
  NOR2_X1 U16727 ( .A1(n15688), .A2(n16512), .ZN(n15533) );
  AOI211_X1 U16728 ( .C1(n16522), .C2(P1_REG2_REG_22__SCAN_IN), .A(n15534), 
        .B(n15533), .ZN(n15535) );
  OAI21_X1 U16729 ( .B1(n15621), .B2(n15687), .A(n15535), .ZN(n15536) );
  AOI21_X1 U16730 ( .B1(n15690), .B2(n15537), .A(n15536), .ZN(n15538) );
  OAI21_X1 U16731 ( .B1(n15592), .B2(n15692), .A(n15538), .ZN(P1_U3271) );
  AOI21_X1 U16732 ( .B1(n7524), .B2(n15543), .A(n16479), .ZN(n15541) );
  AOI21_X1 U16733 ( .B1(n15541), .B2(n15540), .A(n15539), .ZN(n15696) );
  OAI21_X1 U16734 ( .B1(n15544), .B2(n15543), .A(n15542), .ZN(n15545) );
  INV_X1 U16735 ( .A(n15545), .ZN(n15697) );
  NAND2_X1 U16736 ( .A1(n16522), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n15546) );
  OAI21_X1 U16737 ( .B1(n16490), .B2(n15547), .A(n15546), .ZN(n15548) );
  AOI21_X1 U16738 ( .B1(n15694), .B2(n15619), .A(n15548), .ZN(n15552) );
  INV_X1 U16739 ( .A(n15694), .ZN(n15549) );
  XNOR2_X1 U16740 ( .A(n15565), .B(n15549), .ZN(n15550) );
  AND2_X1 U16741 ( .A1(n15550), .A2(n16473), .ZN(n15693) );
  NAND2_X1 U16742 ( .A1(n15693), .A2(n16518), .ZN(n15551) );
  OAI211_X1 U16743 ( .C1(n15697), .C2(n15592), .A(n15552), .B(n15551), .ZN(
        n15553) );
  INV_X1 U16744 ( .A(n15553), .ZN(n15554) );
  OAI21_X1 U16745 ( .B1(n16522), .B2(n15696), .A(n15554), .ZN(P1_U3272) );
  OAI211_X1 U16746 ( .C1(n7574), .C2(n15559), .A(n15555), .B(n16536), .ZN(
        n15558) );
  INV_X1 U16747 ( .A(n15556), .ZN(n15557) );
  AND2_X1 U16748 ( .A1(n15558), .A2(n15557), .ZN(n15701) );
  OAI21_X1 U16749 ( .B1(n15561), .B2(n9667), .A(n15560), .ZN(n15702) );
  NAND2_X1 U16750 ( .A1(n16522), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n15562) );
  OAI21_X1 U16751 ( .B1(n16490), .B2(n15563), .A(n15562), .ZN(n15564) );
  AOI21_X1 U16752 ( .B1(n15699), .B2(n15619), .A(n15564), .ZN(n15568) );
  AOI21_X1 U16753 ( .B1(n15573), .B2(n15699), .A(n16437), .ZN(n15566) );
  AND2_X1 U16754 ( .A1(n15566), .A2(n15565), .ZN(n15698) );
  NAND2_X1 U16755 ( .A1(n15698), .A2(n16518), .ZN(n15567) );
  OAI211_X1 U16756 ( .C1(n15702), .C2(n15592), .A(n15568), .B(n15567), .ZN(
        n15569) );
  INV_X1 U16757 ( .A(n15569), .ZN(n15570) );
  OAI21_X1 U16758 ( .B1(n16522), .B2(n15701), .A(n15570), .ZN(P1_U3273) );
  XOR2_X1 U16759 ( .A(n15571), .B(n15580), .Z(n15707) );
  INV_X1 U16760 ( .A(n15572), .ZN(n15575) );
  INV_X1 U16761 ( .A(n15573), .ZN(n15574) );
  AOI21_X1 U16762 ( .B1(n15703), .B2(n15575), .A(n15574), .ZN(n15704) );
  INV_X1 U16763 ( .A(n15576), .ZN(n15577) );
  AOI22_X1 U16764 ( .A1(n16522), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n15577), 
        .B2(n16508), .ZN(n15578) );
  OAI21_X1 U16765 ( .B1(n15579), .B2(n16512), .A(n15578), .ZN(n15589) );
  INV_X1 U16766 ( .A(n15602), .ZN(n15582) );
  OAI21_X1 U16767 ( .B1(n15582), .B2(n15581), .A(n15580), .ZN(n15584) );
  AOI21_X1 U16768 ( .B1(n15584), .B2(n15583), .A(n16479), .ZN(n15587) );
  INV_X1 U16769 ( .A(n15585), .ZN(n15586) );
  NOR2_X1 U16770 ( .A1(n15587), .A2(n15586), .ZN(n15706) );
  NOR2_X1 U16771 ( .A1(n15706), .A2(n16522), .ZN(n15588) );
  AOI211_X1 U16772 ( .C1(n15704), .C2(n15590), .A(n15589), .B(n15588), .ZN(
        n15591) );
  OAI21_X1 U16773 ( .B1(n15707), .B2(n15592), .A(n15591), .ZN(P1_U3274) );
  XOR2_X1 U16774 ( .A(n15593), .B(n15601), .Z(n15708) );
  INV_X1 U16775 ( .A(n15708), .ZN(n15609) );
  INV_X1 U16776 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15595) );
  OAI22_X1 U16777 ( .A1(n15515), .A2(n15595), .B1(n15594), .B2(n16490), .ZN(
        n15599) );
  INV_X1 U16778 ( .A(n15710), .ZN(n15596) );
  XNOR2_X1 U16779 ( .A(n15613), .B(n15596), .ZN(n15597) );
  NAND2_X1 U16780 ( .A1(n15597), .A2(n16473), .ZN(n15711) );
  NOR2_X1 U16781 ( .A1(n15711), .A2(n15621), .ZN(n15598) );
  AOI211_X1 U16782 ( .C1(n15619), .C2(n15710), .A(n15599), .B(n15598), .ZN(
        n15607) );
  AOI21_X1 U16783 ( .B1(n15600), .B2(n15601), .A(n16479), .ZN(n15603) );
  NAND2_X1 U16784 ( .A1(n15603), .A2(n15602), .ZN(n15712) );
  INV_X1 U16785 ( .A(n15712), .ZN(n15605) );
  INV_X1 U16786 ( .A(n15604), .ZN(n15709) );
  OAI21_X1 U16787 ( .B1(n15605), .B2(n15709), .A(n15515), .ZN(n15606) );
  OAI211_X1 U16788 ( .C1(n15609), .C2(n15608), .A(n15607), .B(n15606), .ZN(
        P1_U3275) );
  XNOR2_X1 U16789 ( .A(n15610), .B(n15611), .ZN(n15721) );
  XNOR2_X1 U16790 ( .A(n15612), .B(n15611), .ZN(n15719) );
  AOI21_X1 U16791 ( .B1(n15632), .B2(n15715), .A(n16437), .ZN(n15614) );
  NAND2_X1 U16792 ( .A1(n15614), .A2(n15613), .ZN(n15717) );
  NOR2_X1 U16793 ( .A1(n15515), .A2(n15615), .ZN(n15618) );
  OAI22_X1 U16794 ( .A1(n16522), .A2(n15716), .B1(n15616), .B2(n16490), .ZN(
        n15617) );
  AOI211_X1 U16795 ( .C1(n15715), .C2(n15619), .A(n15618), .B(n15617), .ZN(
        n15620) );
  OAI21_X1 U16796 ( .B1(n15717), .B2(n15621), .A(n15620), .ZN(n15622) );
  AOI21_X1 U16797 ( .B1(n15719), .B2(n15641), .A(n15622), .ZN(n15623) );
  OAI21_X1 U16798 ( .B1(n15721), .B2(n15643), .A(n15623), .ZN(P1_U3276) );
  OAI21_X1 U16799 ( .B1(n15626), .B2(n15625), .A(n15624), .ZN(n15627) );
  INV_X1 U16800 ( .A(n15627), .ZN(n15728) );
  OAI21_X1 U16801 ( .B1(n15630), .B2(n15629), .A(n15628), .ZN(n15722) );
  INV_X1 U16802 ( .A(n15725), .ZN(n15639) );
  AOI21_X1 U16803 ( .B1(n15631), .B2(n15725), .A(n16437), .ZN(n15633) );
  AND2_X1 U16804 ( .A1(n15633), .A2(n15632), .ZN(n15723) );
  NAND2_X1 U16805 ( .A1(n15723), .A2(n16518), .ZN(n15638) );
  INV_X1 U16806 ( .A(n15724), .ZN(n15635) );
  OAI22_X1 U16807 ( .A1(n16522), .A2(n15635), .B1(n15634), .B2(n16490), .ZN(
        n15636) );
  AOI21_X1 U16808 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n16522), .A(n15636), 
        .ZN(n15637) );
  OAI211_X1 U16809 ( .C1(n15639), .C2(n16512), .A(n15638), .B(n15637), .ZN(
        n15640) );
  AOI21_X1 U16810 ( .B1(n15722), .B2(n15641), .A(n15640), .ZN(n15642) );
  OAI21_X1 U16811 ( .B1(n15728), .B2(n15643), .A(n15642), .ZN(P1_U3277) );
  OAI211_X1 U16812 ( .C1(n15645), .C2(n16476), .A(n15644), .B(n15646), .ZN(
        n15742) );
  MUX2_X1 U16813 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15742), .S(n7435), .Z(
        P1_U3559) );
  OAI211_X1 U16814 ( .C1(n15648), .C2(n16476), .A(n15647), .B(n15646), .ZN(
        n15743) );
  MUX2_X1 U16815 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15743), .S(n7435), .Z(
        P1_U3558) );
  AOI211_X1 U16816 ( .C1(n16573), .C2(n15651), .A(n15650), .B(n15649), .ZN(
        n15654) );
  NAND3_X1 U16817 ( .A1(n15652), .A2(n16443), .A3(n15447), .ZN(n15653) );
  OAI211_X1 U16818 ( .C1(n15655), .C2(n16479), .A(n15654), .B(n15653), .ZN(
        n15744) );
  MUX2_X1 U16819 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15744), .S(n7435), .Z(
        P1_U3556) );
  NAND2_X1 U16820 ( .A1(n15656), .A2(n16536), .ZN(n15661) );
  AOI211_X1 U16821 ( .C1(n16573), .C2(n15659), .A(n15658), .B(n15657), .ZN(
        n15660) );
  OAI211_X1 U16822 ( .C1(n16576), .C2(n15662), .A(n15661), .B(n15660), .ZN(
        n15745) );
  MUX2_X1 U16823 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15745), .S(n7435), .Z(
        P1_U3555) );
  AOI21_X1 U16824 ( .B1(n16573), .B2(n15664), .A(n15663), .ZN(n15665) );
  OAI211_X1 U16825 ( .C1(n16576), .C2(n15667), .A(n15666), .B(n15665), .ZN(
        n15746) );
  MUX2_X1 U16826 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15746), .S(n7435), .Z(
        P1_U3554) );
  NAND2_X1 U16827 ( .A1(n15668), .A2(n16573), .ZN(n15672) );
  NAND3_X1 U16828 ( .A1(n15669), .A2(n16443), .A3(n15485), .ZN(n15671) );
  NAND4_X1 U16829 ( .A1(n15673), .A2(n15672), .A3(n15671), .A4(n15670), .ZN(
        n15747) );
  MUX2_X1 U16830 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15747), .S(n7435), .Z(
        P1_U3553) );
  AOI21_X1 U16831 ( .B1(n16573), .B2(n15675), .A(n15674), .ZN(n15676) );
  OAI211_X1 U16832 ( .C1(n16576), .C2(n15678), .A(n15677), .B(n15676), .ZN(
        n15748) );
  MUX2_X1 U16833 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15748), .S(n7435), .Z(
        P1_U3552) );
  AOI211_X1 U16834 ( .C1(n16573), .C2(n15681), .A(n15680), .B(n15679), .ZN(
        n15684) );
  NAND3_X1 U16835 ( .A1(n15520), .A2(n16443), .A3(n15682), .ZN(n15683) );
  OAI211_X1 U16836 ( .C1(n15685), .C2(n16479), .A(n15684), .B(n15683), .ZN(
        n15749) );
  MUX2_X1 U16837 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15749), .S(n7435), .Z(
        P1_U3551) );
  OAI211_X1 U16838 ( .C1(n16476), .C2(n15688), .A(n15687), .B(n15686), .ZN(
        n15689) );
  AOI21_X1 U16839 ( .B1(n15690), .B2(n16536), .A(n15689), .ZN(n15691) );
  OAI21_X1 U16840 ( .B1(n16576), .B2(n15692), .A(n15691), .ZN(n15750) );
  MUX2_X1 U16841 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15750), .S(n7435), .Z(
        P1_U3550) );
  AOI21_X1 U16842 ( .B1(n16573), .B2(n15694), .A(n15693), .ZN(n15695) );
  OAI211_X1 U16843 ( .C1(n15697), .C2(n16576), .A(n15696), .B(n15695), .ZN(
        n15751) );
  MUX2_X1 U16844 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15751), .S(n7435), .Z(
        P1_U3549) );
  AOI21_X1 U16845 ( .B1(n16573), .B2(n15699), .A(n15698), .ZN(n15700) );
  OAI211_X1 U16846 ( .C1(n15702), .C2(n16576), .A(n15701), .B(n15700), .ZN(
        n15752) );
  MUX2_X1 U16847 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15752), .S(n7435), .Z(
        P1_U3548) );
  AOI22_X1 U16848 ( .A1(n15704), .A2(n16473), .B1(n16573), .B2(n15703), .ZN(
        n15705) );
  OAI211_X1 U16849 ( .C1(n15707), .C2(n16576), .A(n15706), .B(n15705), .ZN(
        n15753) );
  MUX2_X1 U16850 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15753), .S(n7435), .Z(
        P1_U3547) );
  NAND2_X1 U16851 ( .A1(n15708), .A2(n16443), .ZN(n15714) );
  AOI21_X1 U16852 ( .B1(n15710), .B2(n16573), .A(n15709), .ZN(n15713) );
  NAND4_X1 U16853 ( .A1(n15714), .A2(n15713), .A3(n15712), .A4(n15711), .ZN(
        n15754) );
  MUX2_X1 U16854 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15754), .S(n7435), .Z(
        P1_U3546) );
  OAI211_X1 U16855 ( .C1(n8098), .C2(n16476), .A(n15717), .B(n15716), .ZN(
        n15718) );
  AOI21_X1 U16856 ( .B1(n15719), .B2(n16443), .A(n15718), .ZN(n15720) );
  OAI21_X1 U16857 ( .B1(n16479), .B2(n15721), .A(n15720), .ZN(n15755) );
  MUX2_X1 U16858 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15755), .S(n7435), .Z(
        P1_U3545) );
  NAND2_X1 U16859 ( .A1(n15722), .A2(n16443), .ZN(n15727) );
  AOI211_X1 U16860 ( .C1(n16573), .C2(n15725), .A(n15724), .B(n15723), .ZN(
        n15726) );
  OAI211_X1 U16861 ( .C1(n15728), .C2(n16479), .A(n15727), .B(n15726), .ZN(
        n15756) );
  MUX2_X1 U16862 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15756), .S(n7435), .Z(
        P1_U3544) );
  NOR2_X1 U16863 ( .A1(n15729), .A2(n16437), .ZN(n15730) );
  AOI211_X1 U16864 ( .C1(n16573), .C2(n15732), .A(n15731), .B(n15730), .ZN(
        n15736) );
  NAND3_X1 U16865 ( .A1(n15734), .A2(n16536), .A3(n15733), .ZN(n15735) );
  OAI211_X1 U16866 ( .C1(n15737), .C2(n16576), .A(n15736), .B(n15735), .ZN(
        n15757) );
  MUX2_X1 U16867 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15757), .S(n7435), .Z(
        P1_U3543) );
  AOI21_X1 U16868 ( .B1(n16573), .B2(n16611), .A(n15738), .ZN(n15739) );
  OAI211_X1 U16869 ( .C1(n15741), .C2(n16576), .A(n15740), .B(n15739), .ZN(
        n15758) );
  MUX2_X1 U16870 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15758), .S(n7435), .Z(
        P1_U3542) );
  MUX2_X1 U16871 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15742), .S(n16540), .Z(
        P1_U3527) );
  MUX2_X1 U16872 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15743), .S(n16540), .Z(
        P1_U3526) );
  MUX2_X1 U16873 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15744), .S(n16540), .Z(
        P1_U3524) );
  MUX2_X1 U16874 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15745), .S(n16540), .Z(
        P1_U3523) );
  MUX2_X1 U16875 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15746), .S(n16540), .Z(
        P1_U3522) );
  MUX2_X1 U16876 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15747), .S(n16540), .Z(
        P1_U3521) );
  MUX2_X1 U16877 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15748), .S(n16540), .Z(
        P1_U3520) );
  MUX2_X1 U16878 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15749), .S(n16540), .Z(
        P1_U3519) );
  MUX2_X1 U16879 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15750), .S(n16540), .Z(
        P1_U3518) );
  MUX2_X1 U16880 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15751), .S(n16540), .Z(
        P1_U3517) );
  MUX2_X1 U16881 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15752), .S(n16540), .Z(
        P1_U3516) );
  MUX2_X1 U16882 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15753), .S(n16540), .Z(
        P1_U3515) );
  MUX2_X1 U16883 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15754), .S(n16540), .Z(
        P1_U3513) );
  MUX2_X1 U16884 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15755), .S(n16540), .Z(
        P1_U3510) );
  MUX2_X1 U16885 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15756), .S(n16540), .Z(
        P1_U3507) );
  MUX2_X1 U16886 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15757), .S(n16540), .Z(
        P1_U3504) );
  MUX2_X1 U16887 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15758), .S(n16540), .Z(
        P1_U3501) );
  MUX2_X1 U16888 ( .A(P1_D_REG_0__SCAN_IN), .B(n15759), .S(n15816), .Z(
        P1_U3445) );
  NOR4_X1 U16889 ( .A1(n15761), .A2(P1_IR_REG_30__SCAN_IN), .A3(n15760), .A4(
        P1_U3086), .ZN(n15762) );
  AOI21_X1 U16890 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n15763), .A(n15762), 
        .ZN(n15764) );
  OAI21_X1 U16891 ( .B1(n15765), .B2(n15780), .A(n15764), .ZN(P1_U3324) );
  OAI222_X1 U16892 ( .A1(n15777), .A2(n15771), .B1(n15780), .B2(n15770), .C1(
        P1_U3086), .C2(n15769), .ZN(P1_U3326) );
  OAI222_X1 U16893 ( .A1(n15777), .A2(n15774), .B1(n15780), .B2(n15773), .C1(
        P1_U3086), .C2(n15772), .ZN(P1_U3327) );
  OAI222_X1 U16894 ( .A1(n15777), .A2(n15776), .B1(n15780), .B2(n15775), .C1(
        P1_U3086), .C2(n15885), .ZN(P1_U3328) );
  OAI222_X1 U16895 ( .A1(P1_U3086), .A2(n15781), .B1(n15780), .B2(n15779), 
        .C1(n15778), .C2(n15777), .ZN(P1_U3329) );
  MUX2_X1 U16896 ( .A(n15783), .B(n15782), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16897 ( .A(n15784), .ZN(n15785) );
  MUX2_X1 U16898 ( .A(n15785), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16899 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15786) );
  NOR2_X1 U16900 ( .A1(n15816), .A2(n15786), .ZN(P1_U3323) );
  INV_X1 U16901 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n15787) );
  NOR2_X1 U16902 ( .A1(n15816), .A2(n15787), .ZN(P1_U3322) );
  INV_X1 U16903 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15788) );
  NOR2_X1 U16904 ( .A1(n15816), .A2(n15788), .ZN(P1_U3321) );
  INV_X1 U16905 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15789) );
  NOR2_X1 U16906 ( .A1(n15816), .A2(n15789), .ZN(P1_U3320) );
  INV_X1 U16907 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n15790) );
  NOR2_X1 U16908 ( .A1(n15816), .A2(n15790), .ZN(P1_U3319) );
  INV_X1 U16909 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15791) );
  NOR2_X1 U16910 ( .A1(n15816), .A2(n15791), .ZN(P1_U3318) );
  INV_X1 U16911 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15792) );
  NOR2_X1 U16912 ( .A1(n15816), .A2(n15792), .ZN(P1_U3317) );
  INV_X1 U16913 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15793) );
  NOR2_X1 U16914 ( .A1(n15816), .A2(n15793), .ZN(P1_U3316) );
  INV_X1 U16915 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15794) );
  NOR2_X1 U16916 ( .A1(n15816), .A2(n15794), .ZN(P1_U3315) );
  INV_X1 U16917 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15795) );
  NOR2_X1 U16918 ( .A1(n15816), .A2(n15795), .ZN(P1_U3314) );
  INV_X1 U16919 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n15796) );
  NOR2_X1 U16920 ( .A1(n15816), .A2(n15796), .ZN(P1_U3313) );
  INV_X1 U16921 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15797) );
  NOR2_X1 U16922 ( .A1(n15816), .A2(n15797), .ZN(P1_U3312) );
  INV_X1 U16923 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15798) );
  NOR2_X1 U16924 ( .A1(n15816), .A2(n15798), .ZN(P1_U3311) );
  INV_X1 U16925 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15799) );
  NOR2_X1 U16926 ( .A1(n15816), .A2(n15799), .ZN(P1_U3310) );
  INV_X1 U16927 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15800) );
  NOR2_X1 U16928 ( .A1(n15816), .A2(n15800), .ZN(P1_U3309) );
  INV_X1 U16929 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15801) );
  NOR2_X1 U16930 ( .A1(n15816), .A2(n15801), .ZN(P1_U3308) );
  INV_X1 U16931 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15802) );
  NOR2_X1 U16932 ( .A1(n15816), .A2(n15802), .ZN(P1_U3307) );
  INV_X1 U16933 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15803) );
  NOR2_X1 U16934 ( .A1(n15816), .A2(n15803), .ZN(P1_U3306) );
  INV_X1 U16935 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15804) );
  NOR2_X1 U16936 ( .A1(n15816), .A2(n15804), .ZN(P1_U3305) );
  INV_X1 U16937 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15805) );
  NOR2_X1 U16938 ( .A1(n15816), .A2(n15805), .ZN(P1_U3304) );
  INV_X1 U16939 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n15806) );
  NOR2_X1 U16940 ( .A1(n15816), .A2(n15806), .ZN(P1_U3303) );
  INV_X1 U16941 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15807) );
  NOR2_X1 U16942 ( .A1(n15816), .A2(n15807), .ZN(P1_U3302) );
  INV_X1 U16943 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15808) );
  NOR2_X1 U16944 ( .A1(n15816), .A2(n15808), .ZN(P1_U3301) );
  INV_X1 U16945 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15809) );
  NOR2_X1 U16946 ( .A1(n15816), .A2(n15809), .ZN(P1_U3300) );
  INV_X1 U16947 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n15810) );
  NOR2_X1 U16948 ( .A1(n15816), .A2(n15810), .ZN(P1_U3299) );
  INV_X1 U16949 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n15811) );
  NOR2_X1 U16950 ( .A1(n15816), .A2(n15811), .ZN(P1_U3298) );
  INV_X1 U16951 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15812) );
  NOR2_X1 U16952 ( .A1(n15816), .A2(n15812), .ZN(P1_U3297) );
  INV_X1 U16953 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15813) );
  NOR2_X1 U16954 ( .A1(n15816), .A2(n15813), .ZN(P1_U3296) );
  INV_X1 U16955 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15814) );
  NOR2_X1 U16956 ( .A1(n15816), .A2(n15814), .ZN(P1_U3295) );
  INV_X1 U16957 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15815) );
  NOR2_X1 U16958 ( .A1(n15816), .A2(n15815), .ZN(P1_U3294) );
  AOI21_X1 U16959 ( .B1(n15818), .B2(n15822), .A(n15817), .ZN(P2_U3417) );
  AND2_X1 U16960 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15820), .ZN(P2_U3295) );
  AND2_X1 U16961 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15820), .ZN(P2_U3294) );
  AND2_X1 U16962 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15820), .ZN(P2_U3293) );
  AND2_X1 U16963 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15820), .ZN(P2_U3292) );
  AND2_X1 U16964 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15820), .ZN(P2_U3291) );
  AND2_X1 U16965 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15820), .ZN(P2_U3290) );
  AND2_X1 U16966 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15820), .ZN(P2_U3289) );
  AND2_X1 U16967 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15820), .ZN(P2_U3288) );
  AND2_X1 U16968 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15820), .ZN(P2_U3287) );
  AND2_X1 U16969 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15820), .ZN(P2_U3286) );
  AND2_X1 U16970 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15820), .ZN(P2_U3285) );
  AND2_X1 U16971 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15820), .ZN(P2_U3284) );
  AND2_X1 U16972 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15820), .ZN(P2_U3283) );
  AND2_X1 U16973 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15820), .ZN(P2_U3282) );
  AND2_X1 U16974 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15820), .ZN(P2_U3281) );
  AND2_X1 U16975 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15820), .ZN(P2_U3280) );
  AND2_X1 U16976 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15820), .ZN(P2_U3279) );
  AND2_X1 U16977 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15820), .ZN(P2_U3278) );
  AND2_X1 U16978 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15820), .ZN(P2_U3277) );
  AND2_X1 U16979 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15820), .ZN(P2_U3276) );
  AND2_X1 U16980 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15820), .ZN(P2_U3275) );
  AND2_X1 U16981 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15820), .ZN(P2_U3274) );
  AND2_X1 U16982 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15820), .ZN(P2_U3273) );
  AND2_X1 U16983 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15820), .ZN(P2_U3272) );
  AND2_X1 U16984 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15820), .ZN(P2_U3271) );
  AND2_X1 U16985 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15820), .ZN(P2_U3270) );
  AND2_X1 U16986 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15820), .ZN(P2_U3269) );
  AND2_X1 U16987 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15820), .ZN(P2_U3268) );
  AND2_X1 U16988 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15820), .ZN(P2_U3267) );
  AND2_X1 U16989 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15820), .ZN(P2_U3266) );
  NOR2_X1 U16990 ( .A1(n15875), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U16991 ( .A1(P3_U3897), .A2(n16259), .ZN(P3_U3150) );
  AOI21_X1 U16992 ( .B1(n15823), .B2(n15822), .A(n15821), .ZN(P2_U3416) );
  OAI21_X1 U16993 ( .B1(n15869), .B2(n15824), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15825) );
  OAI21_X1 U16994 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15825), .ZN(n15838) );
  AOI211_X1 U16995 ( .C1(n15828), .C2(n15827), .A(n15826), .B(n15848), .ZN(
        n15829) );
  INV_X1 U16996 ( .A(n15829), .ZN(n15837) );
  AOI211_X1 U16997 ( .C1(n15833), .C2(n15832), .A(n15831), .B(n15830), .ZN(
        n15834) );
  INV_X1 U16998 ( .A(n15834), .ZN(n15836) );
  NAND2_X1 U16999 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(n15875), .ZN(n15835) );
  NAND4_X1 U17000 ( .A1(n15838), .A2(n15837), .A3(n15836), .A4(n15835), .ZN(
        P2_U3217) );
  NAND2_X1 U17001 ( .A1(n15875), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n15839) );
  OAI211_X1 U17002 ( .C1(n15842), .C2(n15841), .A(n15840), .B(n15839), .ZN(
        n15843) );
  INV_X1 U17003 ( .A(n15843), .ZN(n15855) );
  NAND2_X1 U17004 ( .A1(n15845), .A2(n15844), .ZN(n15846) );
  NAND3_X1 U17005 ( .A1(n15873), .A2(n15847), .A3(n15846), .ZN(n15854) );
  AOI211_X1 U17006 ( .C1(n15851), .C2(n15850), .A(n15849), .B(n15848), .ZN(
        n15852) );
  INV_X1 U17007 ( .A(n15852), .ZN(n15853) );
  NAND3_X1 U17008 ( .A1(n15855), .A2(n15854), .A3(n15853), .ZN(P2_U3220) );
  AOI22_X1 U17009 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .B1(
        P2_ADDR_REG_16__SCAN_IN), .B2(n15875), .ZN(n15867) );
  XOR2_X1 U17010 ( .A(n15857), .B(n15856), .Z(n15858) );
  NAND2_X1 U17011 ( .A1(n15858), .A2(n15873), .ZN(n15866) );
  NAND2_X1 U17012 ( .A1(n15860), .A2(n15859), .ZN(n15865) );
  OAI211_X1 U17013 ( .C1(n15863), .C2(n15862), .A(n15861), .B(n15877), .ZN(
        n15864) );
  NAND4_X1 U17014 ( .A1(n15867), .A2(n15866), .A3(n15865), .A4(n15864), .ZN(
        P2_U3230) );
  OAI21_X1 U17015 ( .B1(n15869), .B2(n15868), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15870) );
  OAI21_X1 U17016 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15870), .ZN(n15883) );
  XOR2_X1 U17017 ( .A(n15872), .B(n15871), .Z(n15874) );
  NAND2_X1 U17018 ( .A1(n15874), .A2(n15873), .ZN(n15882) );
  NAND2_X1 U17019 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n15875), .ZN(n15881) );
  OAI211_X1 U17020 ( .C1(n15879), .C2(n15878), .A(n15877), .B(n15876), .ZN(
        n15880) );
  NAND4_X1 U17021 ( .A1(n15883), .A2(n15882), .A3(n15881), .A4(n15880), .ZN(
        P2_U3231) );
  INV_X1 U17022 ( .A(n15884), .ZN(n15886) );
  NAND2_X1 U17023 ( .A1(n15885), .A2(n9246), .ZN(n15888) );
  NAND2_X1 U17024 ( .A1(n15886), .A2(n15888), .ZN(n15889) );
  MUX2_X1 U17025 ( .A(n15889), .B(n15888), .S(n15887), .Z(n15891) );
  NAND2_X1 U17026 ( .A1(n15891), .A2(n15890), .ZN(n15894) );
  AOI22_X1 U17027 ( .A1(n15892), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15893) );
  OAI21_X1 U17028 ( .B1(n15895), .B2(n15894), .A(n15893), .ZN(P1_U3243) );
  INV_X1 U17029 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n16088) );
  OAI21_X1 U17030 ( .B1(n15898), .B2(n15897), .A(n15896), .ZN(n15903) );
  OAI21_X1 U17031 ( .B1(n15901), .B2(n15900), .A(n15899), .ZN(n15902) );
  OAI222_X1 U17032 ( .A1(n15928), .A2(n15904), .B1(n16285), .B2(n15903), .C1(
        n15925), .C2(n15902), .ZN(n15905) );
  INV_X1 U17033 ( .A(n15905), .ZN(n15907) );
  OAI211_X1 U17034 ( .C1(n16088), .C2(n16301), .A(n15907), .B(n15906), .ZN(
        P1_U3260) );
  INV_X1 U17035 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n16101) );
  OAI21_X1 U17036 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n15909), .A(n15908), 
        .ZN(n15913) );
  OAI21_X1 U17037 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n15911), .A(n15910), 
        .ZN(n15912) );
  OAI222_X1 U17038 ( .A1(n15928), .A2(n15914), .B1(n16285), .B2(n15913), .C1(
        n15925), .C2(n15912), .ZN(n15915) );
  INV_X1 U17039 ( .A(n15915), .ZN(n15917) );
  OAI211_X1 U17040 ( .C1(n16101), .C2(n16301), .A(n15917), .B(n15916), .ZN(
        P1_U3261) );
  INV_X1 U17041 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n16078) );
  OAI21_X1 U17042 ( .B1(n15920), .B2(n15919), .A(n15918), .ZN(n15926) );
  OAI21_X1 U17043 ( .B1(n15923), .B2(n15922), .A(n15921), .ZN(n15924) );
  OAI222_X1 U17044 ( .A1(n15928), .A2(n15927), .B1(n16285), .B2(n15926), .C1(
        n15925), .C2(n15924), .ZN(n15929) );
  INV_X1 U17045 ( .A(n15929), .ZN(n15931) );
  OAI211_X1 U17046 ( .C1(n16078), .C2(n16301), .A(n15931), .B(n15930), .ZN(
        P1_U3259) );
  INV_X1 U17047 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n15932) );
  AOI22_X1 U17048 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .B1(n15932), .B2(n15933), .ZN(n15934) );
  XOR2_X1 U17049 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15934), .Z(SUB_1596_U53) );
  INV_X1 U17050 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15946) );
  XOR2_X1 U17051 ( .A(n15938), .B(n15937), .Z(n16112) );
  NAND2_X1 U17052 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15934), .ZN(n16111) );
  NAND2_X1 U17053 ( .A1(n16112), .A2(n16111), .ZN(n15935) );
  NOR2_X1 U17054 ( .A1(n16112), .A2(n16111), .ZN(n16110) );
  AOI21_X1 U17055 ( .B1(P2_ADDR_REG_1__SCAN_IN), .B2(n15935), .A(n16110), .ZN(
        n15936) );
  INV_X1 U17056 ( .A(n15936), .ZN(n15943) );
  INV_X1 U17057 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n15941) );
  XNOR2_X1 U17058 ( .A(n15950), .B(n15951), .ZN(n15942) );
  NAND2_X1 U17059 ( .A1(n15943), .A2(n15942), .ZN(n15945) );
  NOR2_X1 U17060 ( .A1(n15943), .A2(n15942), .ZN(n15944) );
  INV_X1 U17061 ( .A(n15944), .ZN(n15948) );
  NAND2_X1 U17062 ( .A1(n15946), .A2(n15945), .ZN(n15947) );
  OAI222_X1 U17063 ( .A1(n15946), .A2(n15945), .B1(n15946), .B2(n15948), .C1(
        n15944), .C2(n15947), .ZN(SUB_1596_U61) );
  NAND2_X1 U17064 ( .A1(n15948), .A2(n15947), .ZN(n15961) );
  INV_X1 U17065 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n16130) );
  NAND2_X1 U17066 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n15949), .ZN(n15952) );
  XNOR2_X1 U17067 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n15957), .ZN(n15962) );
  XOR2_X1 U17068 ( .A(n15961), .B(n15962), .Z(n15954) );
  INV_X1 U17069 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15953) );
  NAND2_X1 U17070 ( .A1(n15954), .A2(n15953), .ZN(n15963) );
  OAI21_X1 U17071 ( .B1(n15954), .B2(n15953), .A(n15963), .ZN(SUB_1596_U60) );
  NAND2_X1 U17072 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n15955), .ZN(n15959) );
  INV_X1 U17073 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15956) );
  NAND2_X1 U17074 ( .A1(n15957), .A2(n15956), .ZN(n15958) );
  NAND2_X1 U17075 ( .A1(n15962), .A2(n15961), .ZN(n15964) );
  NAND2_X1 U17076 ( .A1(n15964), .A2(n15963), .ZN(n15965) );
  NOR2_X1 U17077 ( .A1(n15966), .A2(n15965), .ZN(n15973) );
  AOI21_X1 U17078 ( .B1(n15966), .B2(n15965), .A(n15973), .ZN(SUB_1596_U59) );
  NAND2_X1 U17079 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n15967), .ZN(n15970) );
  INV_X1 U17080 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n16300) );
  NAND2_X1 U17081 ( .A1(n15968), .A2(n16300), .ZN(n15969) );
  INV_X1 U17082 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15976) );
  NOR2_X1 U17083 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n15976), .ZN(n15977) );
  AOI21_X1 U17084 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(n15976), .A(n15977), .ZN(
        n15971) );
  XOR2_X1 U17085 ( .A(n15978), .B(n15971), .Z(n15982) );
  AND2_X1 U17086 ( .A1(n15972), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n15974) );
  NAND2_X1 U17087 ( .A1(n15983), .A2(n15982), .ZN(n15984) );
  OAI21_X1 U17088 ( .B1(n15982), .B2(n15983), .A(n15984), .ZN(n15975) );
  XNOR2_X1 U17089 ( .A(n15975), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  NAND2_X1 U17090 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n15976), .ZN(n15979) );
  INV_X1 U17091 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n16150) );
  NAND2_X1 U17092 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n16150), .ZN(n15980) );
  OAI21_X1 U17093 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n16150), .A(n15980), .ZN(
        n15981) );
  XOR2_X1 U17094 ( .A(n15987), .B(n15981), .Z(n16108) );
  NAND2_X1 U17095 ( .A1(n16108), .A2(n16107), .ZN(n15985) );
  OR2_X1 U17096 ( .A1(n16150), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n15986) );
  XNOR2_X1 U17097 ( .A(n15988), .B(n15995), .ZN(n15997) );
  XNOR2_X1 U17098 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n15997), .ZN(n15989) );
  OAI21_X1 U17099 ( .B1(n15990), .B2(n15989), .A(n15993), .ZN(SUB_1596_U56) );
  INV_X1 U17100 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n15991) );
  NAND2_X1 U17101 ( .A1(n15992), .A2(n15991), .ZN(n15994) );
  NAND2_X1 U17102 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n15995), .ZN(n15999) );
  NAND2_X1 U17103 ( .A1(n15997), .A2(n15996), .ZN(n15998) );
  XOR2_X1 U17104 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n16006), .Z(n16007) );
  XNOR2_X1 U17105 ( .A(n16007), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n16003) );
  INV_X1 U17106 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n16000) );
  OAI21_X1 U17107 ( .B1(n16001), .B2(n16000), .A(n16004), .ZN(SUB_1596_U55) );
  NAND2_X1 U17108 ( .A1(n16003), .A2(n16002), .ZN(n16005) );
  INV_X1 U17109 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n16012) );
  NOR2_X1 U17110 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n16012), .ZN(n16013) );
  AOI21_X1 U17111 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n16012), .A(n16013), .ZN(
        n16010) );
  NOR2_X1 U17112 ( .A1(P3_ADDR_REG_8__SCAN_IN), .A2(n16006), .ZN(n16009) );
  XOR2_X1 U17113 ( .A(n16010), .B(n16015), .Z(n16017) );
  OAI21_X1 U17114 ( .B1(n16016), .B2(n16017), .A(n16018), .ZN(n16011) );
  XNOR2_X1 U17115 ( .A(n16011), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  NAND2_X1 U17116 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n16012), .ZN(n16014) );
  XOR2_X1 U17117 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n16024) );
  XOR2_X1 U17118 ( .A(n16025), .B(n16024), .Z(n16021) );
  AOI21_X1 U17119 ( .B1(n16021), .B2(n16020), .A(n16022), .ZN(n16019) );
  XOR2_X1 U17120 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n16019), .Z(SUB_1596_U70)
         );
  NAND2_X1 U17121 ( .A1(n16021), .A2(n16020), .ZN(n16023) );
  XNOR2_X1 U17122 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n16030) );
  INV_X1 U17123 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n16027) );
  XNOR2_X1 U17124 ( .A(n16030), .B(n16029), .ZN(n16033) );
  AOI21_X1 U17125 ( .B1(n16034), .B2(n16033), .A(n16035), .ZN(n16028) );
  XOR2_X1 U17126 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n16028), .Z(SUB_1596_U69)
         );
  NAND2_X1 U17127 ( .A1(n16030), .A2(n16029), .ZN(n16031) );
  XOR2_X1 U17128 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .Z(n16037) );
  XOR2_X1 U17129 ( .A(n16038), .B(n16037), .Z(n16043) );
  AOI21_X1 U17130 ( .B1(n16043), .B2(n16042), .A(n16044), .ZN(n16036) );
  XOR2_X1 U17131 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n16036), .Z(SUB_1596_U68)
         );
  XNOR2_X1 U17132 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n16041) );
  XNOR2_X1 U17133 ( .A(n16041), .B(n16053), .ZN(n16047) );
  INV_X1 U17134 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n16045) );
  OAI21_X1 U17135 ( .B1(n16046), .B2(n16045), .A(n16049), .ZN(SUB_1596_U67) );
  NAND2_X1 U17136 ( .A1(n16048), .A2(n16047), .ZN(n16050) );
  INV_X1 U17137 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n16054) );
  NOR2_X1 U17138 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n16051), .ZN(n16052) );
  OAI22_X1 U17139 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n16054), .B1(n16053), 
        .B2(n16052), .ZN(n16059) );
  XNOR2_X1 U17140 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n16060) );
  XOR2_X1 U17141 ( .A(n16059), .B(n16060), .Z(n16057) );
  OAI21_X1 U17142 ( .B1(n16056), .B2(n16057), .A(n16058), .ZN(n16055) );
  XNOR2_X1 U17143 ( .A(n16055), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  INV_X1 U17144 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n16066) );
  INV_X1 U17145 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n16062) );
  NAND2_X1 U17146 ( .A1(n16060), .A2(n16059), .ZN(n16061) );
  INV_X1 U17147 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n16072) );
  XNOR2_X1 U17148 ( .A(n16072), .B(P1_ADDR_REG_15__SCAN_IN), .ZN(n16069) );
  XOR2_X1 U17149 ( .A(n16070), .B(n16069), .Z(n16063) );
  NAND2_X1 U17150 ( .A1(n7499), .A2(n16063), .ZN(n16065) );
  OAI222_X1 U17151 ( .A1(n16066), .A2(n16065), .B1(n16066), .B2(n16068), .C1(
        n16064), .C2(n16067), .ZN(SUB_1596_U65) );
  INV_X1 U17152 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n16077) );
  NOR2_X1 U17153 ( .A1(n16070), .A2(n16069), .ZN(n16071) );
  AOI21_X1 U17154 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n16072), .A(n16071), 
        .ZN(n16079) );
  XNOR2_X1 U17155 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n16079), .ZN(n16080) );
  XNOR2_X1 U17156 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n16080), .ZN(n16074) );
  INV_X1 U17157 ( .A(n16075), .ZN(n16084) );
  OAI222_X1 U17158 ( .A1(n16077), .A2(n16076), .B1(n16077), .B2(n16084), .C1(
        n16075), .C2(n16083), .ZN(SUB_1596_U64) );
  NAND2_X1 U17159 ( .A1(n16079), .A2(n16078), .ZN(n16082) );
  NAND2_X1 U17160 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n16080), .ZN(n16081) );
  NAND2_X1 U17161 ( .A1(n16082), .A2(n16081), .ZN(n16087) );
  XNOR2_X1 U17162 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n16087), .ZN(n16089) );
  XNOR2_X1 U17163 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n16089), .ZN(n16093) );
  XNOR2_X1 U17164 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n16093), .ZN(n16086) );
  NAND2_X1 U17165 ( .A1(n16084), .A2(n16083), .ZN(n16085) );
  AOI21_X1 U17166 ( .B1(n16086), .B2(n16085), .A(n16094), .ZN(SUB_1596_U63) );
  XNOR2_X1 U17167 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n16092) );
  NAND2_X1 U17168 ( .A1(n16088), .A2(n16087), .ZN(n16091) );
  NAND2_X1 U17169 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n16089), .ZN(n16090) );
  NAND2_X1 U17170 ( .A1(n16091), .A2(n16090), .ZN(n16102) );
  XOR2_X1 U17171 ( .A(n16092), .B(n16102), .Z(n16097) );
  AND2_X1 U17172 ( .A1(n16093), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n16095) );
  NAND2_X1 U17173 ( .A1(n16098), .A2(n16097), .ZN(n16099) );
  OAI21_X1 U17174 ( .B1(n16097), .B2(n16098), .A(n16099), .ZN(n16096) );
  XNOR2_X1 U17175 ( .A(n16096), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NOR2_X1 U17176 ( .A1(n16098), .A2(n16097), .ZN(n16100) );
  AND2_X1 U17177 ( .A1(n16101), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n16103) );
  OAI22_X1 U17178 ( .A1(n16103), .A2(n16102), .B1(P3_ADDR_REG_18__SCAN_IN), 
        .B2(n16101), .ZN(n16104) );
  XNOR2_X1 U17179 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n16105) );
  AOI21_X1 U17180 ( .B1(n16108), .B2(n16107), .A(n16106), .ZN(n16109) );
  XOR2_X1 U17181 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n16109), .Z(SUB_1596_U57) );
  AOI21_X1 U17182 ( .B1(n16112), .B2(n16111), .A(n16110), .ZN(n16113) );
  XOR2_X1 U17183 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n16113), .Z(SUB_1596_U5) );
  XNOR2_X1 U17184 ( .A(n16115), .B(n16114), .ZN(n16119) );
  AOI21_X1 U17185 ( .B1(n11003), .B2(n16117), .A(n16116), .ZN(n16118) );
  OAI22_X1 U17186 ( .A1(n16277), .A2(n16119), .B1(n16118), .B2(n16274), .ZN(
        n16127) );
  INV_X1 U17187 ( .A(n16120), .ZN(n16125) );
  NAND3_X1 U17188 ( .A1(n16123), .A2(n16122), .A3(n16121), .ZN(n16124) );
  AOI21_X1 U17189 ( .B1(n16125), .B2(n16124), .A(n16263), .ZN(n16126) );
  AOI211_X1 U17190 ( .C1(n16269), .C2(n7767), .A(n16127), .B(n16126), .ZN(
        n16129) );
  NAND2_X1 U17191 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_U3151), .ZN(n16128) );
  OAI211_X1 U17192 ( .C1(n16151), .C2(n16130), .A(n16129), .B(n16128), .ZN(
        P3_U3185) );
  MUX2_X1 U17193 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n16131), .S(n16143), .Z(
        n16134) );
  NAND2_X1 U17194 ( .A1(n16133), .A2(n16134), .ZN(n16132) );
  OAI21_X1 U17195 ( .B1(n16134), .B2(n16133), .A(n16132), .ZN(n16147) );
  NAND2_X1 U17196 ( .A1(n16136), .A2(n16135), .ZN(n16137) );
  AOI21_X1 U17197 ( .B1(n16138), .B2(n16137), .A(n16274), .ZN(n16146) );
  NAND2_X1 U17198 ( .A1(n7622), .A2(n16139), .ZN(n16140) );
  XNOR2_X1 U17199 ( .A(n16141), .B(n16140), .ZN(n16144) );
  OAI22_X1 U17200 ( .A1(n16144), .A2(n16263), .B1(n16143), .B2(n16142), .ZN(
        n16145) );
  AOI211_X1 U17201 ( .C1(n16194), .C2(n16147), .A(n16146), .B(n16145), .ZN(
        n16149) );
  NAND2_X1 U17202 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n16148) );
  OAI211_X1 U17203 ( .C1(n16151), .C2(n16150), .A(n16149), .B(n16148), .ZN(
        P3_U3188) );
  AOI22_X1 U17204 ( .A1(n16269), .A2(n16152), .B1(n16259), .B2(
        P3_ADDR_REG_11__SCAN_IN), .ZN(n16165) );
  XNOR2_X1 U17205 ( .A(n16154), .B(n16153), .ZN(n16158) );
  OAI21_X1 U17206 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n16156), .A(n16155), 
        .ZN(n16157) );
  AOI22_X1 U17207 ( .A1(n16158), .A2(n16195), .B1(n16194), .B2(n16157), .ZN(
        n16164) );
  NAND2_X1 U17208 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(P3_U3151), .ZN(n16163)
         );
  AOI21_X1 U17209 ( .B1(n16160), .B2(n9944), .A(n16159), .ZN(n16161) );
  OR2_X1 U17210 ( .A1(n16161), .A2(n16274), .ZN(n16162) );
  NAND4_X1 U17211 ( .A1(n16165), .A2(n16164), .A3(n16163), .A4(n16162), .ZN(
        P3_U3193) );
  INV_X1 U17212 ( .A(n16166), .ZN(n16167) );
  AOI22_X1 U17213 ( .A1(n16269), .A2(n16167), .B1(n16259), .B2(
        P3_ADDR_REG_12__SCAN_IN), .ZN(n16186) );
  OAI21_X1 U17214 ( .B1(n16170), .B2(n16169), .A(n16168), .ZN(n16176) );
  OAI211_X1 U17215 ( .C1(n16173), .C2(n16172), .A(n16171), .B(n16195), .ZN(
        n16174) );
  INV_X1 U17216 ( .A(n16174), .ZN(n16175) );
  AOI21_X1 U17217 ( .B1(n16194), .B2(n16176), .A(n16175), .ZN(n16185) );
  NAND2_X1 U17218 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_U3151), .ZN(n16184)
         );
  INV_X1 U17219 ( .A(n16177), .ZN(n16180) );
  OAI21_X1 U17220 ( .B1(n16180), .B2(n16179), .A(n16178), .ZN(n16182) );
  NAND2_X1 U17221 ( .A1(n16182), .A2(n16181), .ZN(n16183) );
  NAND4_X1 U17222 ( .A1(n16186), .A2(n16185), .A3(n16184), .A4(n16183), .ZN(
        P3_U3194) );
  AOI22_X1 U17223 ( .A1(n16269), .A2(n16187), .B1(n16259), .B2(
        P3_ADDR_REG_13__SCAN_IN), .ZN(n16203) );
  OAI21_X1 U17224 ( .B1(n16190), .B2(n16189), .A(n16188), .ZN(n16196) );
  OAI21_X1 U17225 ( .B1(P3_REG2_REG_13__SCAN_IN), .B2(n16192), .A(n16191), 
        .ZN(n16193) );
  AOI22_X1 U17226 ( .A1(n16196), .A2(n16195), .B1(n16194), .B2(n16193), .ZN(
        n16202) );
  AOI21_X1 U17227 ( .B1(n16198), .B2(n16600), .A(n16197), .ZN(n16199) );
  OR2_X1 U17228 ( .A1(n16199), .A2(n16274), .ZN(n16200) );
  NAND4_X1 U17229 ( .A1(n16203), .A2(n16202), .A3(n16201), .A4(n16200), .ZN(
        P3_U3195) );
  XNOR2_X1 U17230 ( .A(n7787), .B(n13306), .ZN(n16205) );
  XNOR2_X1 U17231 ( .A(n16206), .B(n16205), .ZN(n16221) );
  NAND2_X1 U17232 ( .A1(n16259), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n16208) );
  NAND2_X1 U17233 ( .A1(n16208), .A2(n16207), .ZN(n16213) );
  AOI211_X1 U17234 ( .C1(n16211), .C2(n16210), .A(n16263), .B(n16209), .ZN(
        n16212) );
  AOI211_X1 U17235 ( .C1(n16269), .C2(n7787), .A(n16213), .B(n16212), .ZN(
        n16220) );
  INV_X1 U17236 ( .A(n16214), .ZN(n16215) );
  AOI21_X1 U17237 ( .B1(n16217), .B2(n16216), .A(n16215), .ZN(n16218) );
  OR2_X1 U17238 ( .A1(n16218), .A2(n16274), .ZN(n16219) );
  OAI211_X1 U17239 ( .C1(n16277), .C2(n16221), .A(n16220), .B(n16219), .ZN(
        P3_U3196) );
  AOI21_X1 U17240 ( .B1(n16224), .B2(n16223), .A(n16222), .ZN(n16239) );
  NAND2_X1 U17241 ( .A1(n16259), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n16226) );
  NAND2_X1 U17242 ( .A1(n16226), .A2(n16225), .ZN(n16231) );
  AOI211_X1 U17243 ( .C1(n16229), .C2(n16228), .A(n16263), .B(n16227), .ZN(
        n16230) );
  AOI211_X1 U17244 ( .C1(n16269), .C2(n16232), .A(n16231), .B(n16230), .ZN(
        n16238) );
  AOI21_X1 U17245 ( .B1(n16235), .B2(n16234), .A(n16233), .ZN(n16236) );
  OR2_X1 U17246 ( .A1(n16236), .A2(n16274), .ZN(n16237) );
  OAI211_X1 U17247 ( .C1(n16239), .C2(n16277), .A(n16238), .B(n16237), .ZN(
        P3_U3197) );
  AOI21_X1 U17248 ( .B1(n16242), .B2(n16241), .A(n16240), .ZN(n16256) );
  NAND2_X1 U17249 ( .A1(n16259), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n16244) );
  NAND2_X1 U17250 ( .A1(n16244), .A2(n16243), .ZN(n16249) );
  AOI211_X1 U17251 ( .C1(n16247), .C2(n16246), .A(n16263), .B(n16245), .ZN(
        n16248) );
  AOI211_X1 U17252 ( .C1(n16269), .C2(n16250), .A(n16249), .B(n16248), .ZN(
        n16255) );
  AOI21_X1 U17253 ( .B1(n7512), .B2(n16252), .A(n16251), .ZN(n16253) );
  OR2_X1 U17254 ( .A1(n16253), .A2(n16274), .ZN(n16254) );
  OAI211_X1 U17255 ( .C1(n16256), .C2(n16277), .A(n16255), .B(n16254), .ZN(
        P3_U3198) );
  AOI21_X1 U17256 ( .B1(n13258), .B2(n16258), .A(n16257), .ZN(n16278) );
  NAND2_X1 U17257 ( .A1(n16259), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n16261) );
  NAND2_X1 U17258 ( .A1(n16261), .A2(n16260), .ZN(n16267) );
  AOI211_X1 U17259 ( .C1(n16265), .C2(n16264), .A(n16263), .B(n16262), .ZN(
        n16266) );
  AOI211_X1 U17260 ( .C1(n16269), .C2(n16268), .A(n16267), .B(n16266), .ZN(
        n16276) );
  AOI21_X1 U17261 ( .B1(n16272), .B2(n16271), .A(n16270), .ZN(n16273) );
  OR2_X1 U17262 ( .A1(n16274), .A2(n16273), .ZN(n16275) );
  OAI211_X1 U17263 ( .C1(n16278), .C2(n16277), .A(n16276), .B(n16275), .ZN(
        P3_U3199) );
  INV_X1 U17264 ( .A(n16279), .ZN(n16284) );
  NOR3_X1 U17265 ( .A1(n16282), .A2(n16281), .A3(n16280), .ZN(n16283) );
  NOR3_X1 U17266 ( .A1(n16285), .A2(n16284), .A3(n16283), .ZN(n16286) );
  AOI21_X1 U17267 ( .B1(n16287), .B2(n16288), .A(n16286), .ZN(n16296) );
  MUX2_X1 U17268 ( .A(n10595), .B(P1_REG1_REG_4__SCAN_IN), .S(n16288), .Z(
        n16289) );
  NAND3_X1 U17269 ( .A1(n16291), .A2(n16290), .A3(n16289), .ZN(n16292) );
  NAND3_X1 U17270 ( .A1(n16294), .A2(n16293), .A3(n16292), .ZN(n16295) );
  AND3_X1 U17271 ( .A1(n16297), .A2(n16296), .A3(n16295), .ZN(n16299) );
  OAI211_X1 U17272 ( .C1(n16301), .C2(n16300), .A(n16299), .B(n16298), .ZN(
        P1_U3247) );
  INV_X1 U17273 ( .A(n16302), .ZN(n16305) );
  INV_X1 U17274 ( .A(n16303), .ZN(n16304) );
  AOI211_X1 U17275 ( .C1(n16486), .C2(n16306), .A(n16305), .B(n16304), .ZN(
        n16307) );
  AOI22_X1 U17276 ( .A1(n7435), .A2(n16307), .B1(n9246), .B2(n16579), .ZN(
        P1_U3528) );
  AOI22_X1 U17277 ( .A1(n16540), .A2(n16307), .B1(n9247), .B2(n16580), .ZN(
        P1_U3459) );
  XNOR2_X1 U17278 ( .A(n16312), .B(n16308), .ZN(n16319) );
  NOR2_X1 U17279 ( .A1(n16319), .A2(n16414), .ZN(n16315) );
  INV_X1 U17280 ( .A(n16309), .ZN(n16310) );
  AOI21_X1 U17281 ( .B1(n16312), .B2(n16311), .A(n16310), .ZN(n16313) );
  OAI222_X1 U17282 ( .A1(n16350), .A2(n10278), .B1(n16352), .B2(n16314), .C1(
        n16349), .C2(n16313), .ZN(n16322) );
  AOI211_X1 U17283 ( .C1(n16544), .C2(n16316), .A(n16315), .B(n16322), .ZN(
        n16317) );
  AOI22_X1 U17284 ( .A1(n16601), .A2(n16317), .B1(n10991), .B2(n16599), .ZN(
        P3_U3460) );
  INV_X1 U17285 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n16318) );
  AOI22_X1 U17286 ( .A1(n16605), .A2(n16318), .B1(n16317), .B2(n16602), .ZN(
        P3_U3393) );
  INV_X1 U17287 ( .A(n16319), .ZN(n16324) );
  INV_X1 U17288 ( .A(n16320), .ZN(n16362) );
  OAI22_X1 U17289 ( .A1(n8116), .A2(n16362), .B1(n16321), .B2(n16360), .ZN(
        n16323) );
  AOI211_X1 U17290 ( .C1(n16367), .C2(n16324), .A(n16323), .B(n16322), .ZN(
        n16325) );
  AOI22_X1 U17291 ( .A1(n16369), .A2(n10992), .B1(n16325), .B2(n13310), .ZN(
        P3_U3232) );
  XNOR2_X1 U17292 ( .A(n15233), .B(n16326), .ZN(n16341) );
  OR2_X1 U17293 ( .A1(n16327), .A2(n16339), .ZN(n16328) );
  AND3_X1 U17294 ( .A1(n16473), .A2(n16329), .A3(n16328), .ZN(n16342) );
  INV_X1 U17295 ( .A(n16342), .ZN(n16330) );
  OAI21_X1 U17296 ( .B1(n16339), .B2(n16476), .A(n16330), .ZN(n16336) );
  XOR2_X1 U17297 ( .A(n16331), .B(n15233), .Z(n16332) );
  NOR2_X1 U17298 ( .A1(n16332), .A2(n16479), .ZN(n16333) );
  AOI211_X1 U17299 ( .C1(n16483), .C2(n16341), .A(n16334), .B(n16333), .ZN(
        n16345) );
  INV_X1 U17300 ( .A(n16345), .ZN(n16335) );
  AOI211_X1 U17301 ( .C1(n16486), .C2(n16341), .A(n16336), .B(n16335), .ZN(
        n16337) );
  AOI22_X1 U17302 ( .A1(n7435), .A2(n16337), .B1(n10587), .B2(n16579), .ZN(
        P1_U3529) );
  AOI22_X1 U17303 ( .A1(n16540), .A2(n16337), .B1(n9256), .B2(n16580), .ZN(
        P1_U3462) );
  AOI22_X1 U17304 ( .A1(n16522), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n16508), .ZN(n16338) );
  OAI21_X1 U17305 ( .B1(n16512), .B2(n16339), .A(n16338), .ZN(n16340) );
  INV_X1 U17306 ( .A(n16340), .ZN(n16344) );
  AOI22_X1 U17307 ( .A1(n16518), .A2(n16342), .B1(n16513), .B2(n16341), .ZN(
        n16343) );
  OAI211_X1 U17308 ( .C1(n16522), .C2(n16345), .A(n16344), .B(n16343), .ZN(
        P1_U3292) );
  NAND3_X1 U17309 ( .A1(n16309), .A2(n10281), .A3(n16346), .ZN(n16347) );
  AND2_X1 U17310 ( .A1(n11732), .A2(n16347), .ZN(n16348) );
  OAI222_X1 U17311 ( .A1(n16352), .A2(n16351), .B1(n16350), .B2(n9780), .C1(
        n16349), .C2(n16348), .ZN(n16364) );
  INV_X1 U17312 ( .A(n16353), .ZN(n16354) );
  AOI21_X1 U17313 ( .B1(n10277), .B2(n16355), .A(n16354), .ZN(n16359) );
  OAI22_X1 U17314 ( .A1(n16359), .A2(n16414), .B1(n16593), .B2(n16363), .ZN(
        n16356) );
  NOR2_X1 U17315 ( .A1(n16364), .A2(n16356), .ZN(n16357) );
  AOI22_X1 U17316 ( .A1(n16568), .A2(n16357), .B1(n10998), .B2(n16599), .ZN(
        P3_U3461) );
  INV_X1 U17317 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n16358) );
  AOI22_X1 U17318 ( .A1(n16605), .A2(n16358), .B1(n16357), .B2(n16602), .ZN(
        P3_U3396) );
  INV_X1 U17319 ( .A(n16359), .ZN(n16366) );
  OAI22_X1 U17320 ( .A1(n16363), .A2(n16362), .B1(n16361), .B2(n16360), .ZN(
        n16365) );
  AOI211_X1 U17321 ( .C1(n16367), .C2(n16366), .A(n16365), .B(n16364), .ZN(
        n16368) );
  AOI22_X1 U17322 ( .A1(n16369), .A2(n10999), .B1(n16368), .B2(n13310), .ZN(
        P3_U3231) );
  INV_X1 U17323 ( .A(n16377), .ZN(n16371) );
  NOR2_X1 U17324 ( .A1(n16371), .A2(n16370), .ZN(n16376) );
  OAI211_X1 U17325 ( .C1(n16374), .C2(n16476), .A(n16373), .B(n16372), .ZN(
        n16375) );
  AOI211_X1 U17326 ( .C1(n16486), .C2(n16377), .A(n16376), .B(n16375), .ZN(
        n16379) );
  AOI22_X1 U17327 ( .A1(n7435), .A2(n16379), .B1(n10591), .B2(n16579), .ZN(
        P1_U3530) );
  INV_X1 U17328 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n16378) );
  AOI22_X1 U17329 ( .A1(n16540), .A2(n16379), .B1(n16378), .B2(n16580), .ZN(
        P1_U3465) );
  AOI21_X1 U17330 ( .B1(n16382), .B2(n16381), .A(n16380), .ZN(n16383) );
  OAI211_X1 U17331 ( .C1(n16386), .C2(n16385), .A(n16384), .B(n16383), .ZN(
        n16387) );
  INV_X1 U17332 ( .A(n16387), .ZN(n16389) );
  AOI22_X1 U17333 ( .A1(n16560), .A2(n16389), .B1(n8576), .B2(n16559), .ZN(
        P2_U3501) );
  INV_X1 U17334 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n16388) );
  AOI22_X1 U17335 ( .A1(n11936), .A2(n16389), .B1(n16388), .B2(n16561), .ZN(
        P2_U3436) );
  NOR2_X1 U17336 ( .A1(n16390), .A2(n16593), .ZN(n16392) );
  AOI211_X1 U17337 ( .C1(n16597), .C2(n16393), .A(n16392), .B(n16391), .ZN(
        n16394) );
  AOI22_X1 U17338 ( .A1(n16568), .A2(n16394), .B1(n11003), .B2(n16599), .ZN(
        P3_U3462) );
  INV_X1 U17339 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n16395) );
  AOI22_X1 U17340 ( .A1(n16605), .A2(n16395), .B1(n16394), .B2(n16602), .ZN(
        P3_U3399) );
  AND2_X1 U17341 ( .A1(n16396), .A2(n16573), .ZN(n16407) );
  AOI21_X1 U17342 ( .B1(n16398), .B2(n16407), .A(n16397), .ZN(n16403) );
  XOR2_X1 U17343 ( .A(n16400), .B(n16399), .Z(n16401) );
  AOI22_X1 U17344 ( .A1(n16401), .A2(n16612), .B1(n16614), .B2(n16406), .ZN(
        n16402) );
  OAI211_X1 U17345 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n16619), .A(n16403), .B(
        n16402), .ZN(P1_U3218) );
  INV_X1 U17346 ( .A(n16404), .ZN(n16411) );
  AND2_X1 U17347 ( .A1(n16405), .A2(n16536), .ZN(n16409) );
  OR4_X1 U17348 ( .A1(n16409), .A2(n16408), .A3(n16407), .A4(n16406), .ZN(
        n16410) );
  AOI21_X1 U17349 ( .B1(n16411), .B2(n16443), .A(n16410), .ZN(n16412) );
  AOI22_X1 U17350 ( .A1(n7435), .A2(n16412), .B1(n10592), .B2(n16579), .ZN(
        P1_U3531) );
  AOI22_X1 U17351 ( .A1(n16540), .A2(n16412), .B1(n9281), .B2(n16580), .ZN(
        P1_U3468) );
  OAI22_X1 U17352 ( .A1(n16415), .A2(n16414), .B1(n16593), .B2(n16413), .ZN(
        n16416) );
  INV_X1 U17353 ( .A(n16416), .ZN(n16417) );
  AND2_X1 U17354 ( .A1(n16418), .A2(n16417), .ZN(n16419) );
  AOI22_X1 U17355 ( .A1(n16568), .A2(n16419), .B1(n11008), .B2(n16599), .ZN(
        P3_U3463) );
  INV_X1 U17356 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n16420) );
  AOI22_X1 U17357 ( .A1(n16605), .A2(n16420), .B1(n16419), .B2(n16602), .ZN(
        P3_U3402) );
  INV_X1 U17358 ( .A(n16421), .ZN(n16430) );
  NAND3_X1 U17359 ( .A1(n16423), .A2(n16422), .A3(n16536), .ZN(n16428) );
  AOI21_X1 U17360 ( .B1(n16573), .B2(n16425), .A(n16424), .ZN(n16427) );
  NAND3_X1 U17361 ( .A1(n16428), .A2(n16427), .A3(n16426), .ZN(n16429) );
  AOI21_X1 U17362 ( .B1(n16430), .B2(n16443), .A(n16429), .ZN(n16432) );
  AOI22_X1 U17363 ( .A1(n7435), .A2(n16432), .B1(n10595), .B2(n16579), .ZN(
        P1_U3532) );
  INV_X1 U17364 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n16431) );
  AOI22_X1 U17365 ( .A1(n16540), .A2(n16432), .B1(n16431), .B2(n16580), .ZN(
        P1_U3471) );
  XNOR2_X1 U17366 ( .A(n16433), .B(n16434), .ZN(n16453) );
  XOR2_X1 U17367 ( .A(n16435), .B(n16434), .Z(n16436) );
  NOR2_X1 U17368 ( .A1(n16436), .A2(n16479), .ZN(n16446) );
  AOI21_X1 U17369 ( .B1(n16438), .B2(n16448), .A(n16437), .ZN(n16440) );
  AND2_X1 U17370 ( .A1(n16440), .A2(n16439), .ZN(n16454) );
  OR4_X1 U17371 ( .A1(n16446), .A2(n16441), .A3(n16454), .A4(n16447), .ZN(
        n16442) );
  AOI21_X1 U17372 ( .B1(n16453), .B2(n16443), .A(n16442), .ZN(n16445) );
  AOI22_X1 U17373 ( .A1(n7435), .A2(n16445), .B1(n9312), .B2(n16579), .ZN(
        P1_U3533) );
  INV_X1 U17374 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n16444) );
  AOI22_X1 U17375 ( .A1(n16540), .A2(n16445), .B1(n16444), .B2(n16580), .ZN(
        P1_U3474) );
  AOI211_X1 U17376 ( .C1(n16483), .C2(n16453), .A(n16447), .B(n16446), .ZN(
        n16457) );
  NOR2_X1 U17377 ( .A1(n16490), .A2(n16449), .ZN(n16450) );
  AOI21_X1 U17378 ( .B1(n16522), .B2(P1_REG2_REG_5__SCAN_IN), .A(n16450), .ZN(
        n16451) );
  OAI21_X1 U17379 ( .B1(n16512), .B2(n8096), .A(n16451), .ZN(n16452) );
  INV_X1 U17380 ( .A(n16452), .ZN(n16456) );
  AOI22_X1 U17381 ( .A1(n16518), .A2(n16454), .B1(n16513), .B2(n16453), .ZN(
        n16455) );
  OAI211_X1 U17382 ( .C1(n16522), .C2(n16457), .A(n16456), .B(n16455), .ZN(
        P1_U3288) );
  NOR2_X1 U17383 ( .A1(n16458), .A2(n16593), .ZN(n16460) );
  AOI211_X1 U17384 ( .C1(n16597), .C2(n16461), .A(n16460), .B(n16459), .ZN(
        n16462) );
  AOI22_X1 U17385 ( .A1(n16568), .A2(n16462), .B1(n11253), .B2(n16599), .ZN(
        P3_U3465) );
  INV_X1 U17386 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n16463) );
  AOI22_X1 U17387 ( .A1(n16605), .A2(n16463), .B1(n16462), .B2(n16602), .ZN(
        P3_U3408) );
  INV_X1 U17388 ( .A(n16469), .ZN(n16471) );
  AOI21_X1 U17389 ( .B1(n16573), .B2(n16465), .A(n16464), .ZN(n16466) );
  OAI211_X1 U17390 ( .C1(n16469), .C2(n16468), .A(n16467), .B(n16466), .ZN(
        n16470) );
  AOI21_X1 U17391 ( .B1(n16483), .B2(n16471), .A(n16470), .ZN(n16472) );
  AOI22_X1 U17392 ( .A1(n7435), .A2(n16472), .B1(n9323), .B2(n16579), .ZN(
        P1_U3534) );
  AOI22_X1 U17393 ( .A1(n16540), .A2(n16472), .B1(n9327), .B2(n16580), .ZN(
        P1_U3477) );
  OAI21_X1 U17394 ( .B1(n7613), .B2(n16477), .A(n8293), .ZN(n16497) );
  OAI211_X1 U17395 ( .C1(n16493), .C2(n16475), .A(n16474), .B(n16473), .ZN(
        n16495) );
  OAI21_X1 U17396 ( .B1(n16493), .B2(n16476), .A(n16495), .ZN(n16485) );
  XNOR2_X1 U17397 ( .A(n16478), .B(n16477), .ZN(n16480) );
  NOR2_X1 U17398 ( .A1(n16480), .A2(n16479), .ZN(n16481) );
  AOI211_X1 U17399 ( .C1(n16483), .C2(n16497), .A(n16482), .B(n16481), .ZN(
        n16500) );
  INV_X1 U17400 ( .A(n16500), .ZN(n16484) );
  AOI211_X1 U17401 ( .C1(n16486), .C2(n16497), .A(n16485), .B(n16484), .ZN(
        n16488) );
  AOI22_X1 U17402 ( .A1(n7435), .A2(n16488), .B1(n10602), .B2(n16579), .ZN(
        P1_U3535) );
  INV_X1 U17403 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n16487) );
  AOI22_X1 U17404 ( .A1(n16540), .A2(n16488), .B1(n16487), .B2(n16580), .ZN(
        P1_U3480) );
  NOR2_X1 U17405 ( .A1(n16490), .A2(n16489), .ZN(n16491) );
  AOI21_X1 U17406 ( .B1(n16522), .B2(P1_REG2_REG_7__SCAN_IN), .A(n16491), .ZN(
        n16492) );
  OAI21_X1 U17407 ( .B1(n16512), .B2(n16493), .A(n16492), .ZN(n16494) );
  INV_X1 U17408 ( .A(n16494), .ZN(n16499) );
  INV_X1 U17409 ( .A(n16495), .ZN(n16496) );
  AOI22_X1 U17410 ( .A1(n16497), .A2(n16513), .B1(n16518), .B2(n16496), .ZN(
        n16498) );
  OAI211_X1 U17411 ( .C1(n16522), .C2(n16500), .A(n16499), .B(n16498), .ZN(
        P1_U3286) );
  AOI22_X1 U17412 ( .A1(n16502), .A2(n16597), .B1(n16544), .B2(n16501), .ZN(
        n16503) );
  AND2_X1 U17413 ( .A1(n16504), .A2(n16503), .ZN(n16505) );
  AOI22_X1 U17414 ( .A1(n16568), .A2(n16505), .B1(n11537), .B2(n16599), .ZN(
        P3_U3467) );
  INV_X1 U17415 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n16506) );
  AOI22_X1 U17416 ( .A1(n16605), .A2(n16506), .B1(n16505), .B2(n16602), .ZN(
        P3_U3414) );
  INV_X1 U17417 ( .A(n16507), .ZN(n16509) );
  AOI22_X1 U17418 ( .A1(n16522), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n16509), 
        .B2(n16508), .ZN(n16510) );
  OAI21_X1 U17419 ( .B1(n16512), .B2(n16511), .A(n16510), .ZN(n16517) );
  INV_X1 U17420 ( .A(n16513), .ZN(n16514) );
  NOR2_X1 U17421 ( .A1(n16515), .A2(n16514), .ZN(n16516) );
  AOI211_X1 U17422 ( .C1(n16519), .C2(n16518), .A(n16517), .B(n16516), .ZN(
        n16520) );
  OAI21_X1 U17423 ( .B1(n16522), .B2(n16521), .A(n16520), .ZN(P1_U3285) );
  OAI22_X1 U17424 ( .A1(n16524), .A2(n16584), .B1(n16593), .B2(n16523), .ZN(
        n16525) );
  NOR2_X1 U17425 ( .A1(n16526), .A2(n16525), .ZN(n16528) );
  AOI22_X1 U17426 ( .A1(n16568), .A2(n16528), .B1(n16527), .B2(n16599), .ZN(
        P3_U3468) );
  INV_X1 U17427 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n16529) );
  AOI22_X1 U17428 ( .A1(n16605), .A2(n16529), .B1(n16528), .B2(n16602), .ZN(
        P3_U3417) );
  AOI21_X1 U17429 ( .B1(n16531), .B2(n16573), .A(n16530), .ZN(n16533) );
  OAI211_X1 U17430 ( .C1(n16534), .C2(n16576), .A(n16533), .B(n16532), .ZN(
        n16535) );
  AOI21_X1 U17431 ( .B1(n16537), .B2(n16536), .A(n16535), .ZN(n16539) );
  AOI22_X1 U17432 ( .A1(n7435), .A2(n16539), .B1(n9373), .B2(n16579), .ZN(
        P1_U3537) );
  INV_X1 U17433 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n16538) );
  AOI22_X1 U17434 ( .A1(n16540), .A2(n16539), .B1(n16538), .B2(n16580), .ZN(
        P1_U3486) );
  INV_X1 U17435 ( .A(n16541), .ZN(n16589) );
  INV_X1 U17436 ( .A(n16546), .ZN(n16548) );
  AOI21_X1 U17437 ( .B1(n16544), .B2(n16543), .A(n16542), .ZN(n16545) );
  OAI21_X1 U17438 ( .B1(n16546), .B2(n16584), .A(n16545), .ZN(n16547) );
  AOI21_X1 U17439 ( .B1(n16589), .B2(n16548), .A(n16547), .ZN(n16549) );
  AOI22_X1 U17440 ( .A1(n16568), .A2(n16549), .B1(n11820), .B2(n16599), .ZN(
        P3_U3469) );
  INV_X1 U17441 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n16550) );
  AOI22_X1 U17442 ( .A1(n16605), .A2(n16550), .B1(n16549), .B2(n16602), .ZN(
        P3_U3420) );
  INV_X1 U17443 ( .A(n16551), .ZN(n16557) );
  OAI21_X1 U17444 ( .B1(n16554), .B2(n16553), .A(n16552), .ZN(n16556) );
  AOI211_X1 U17445 ( .C1(n16558), .C2(n16557), .A(n16556), .B(n16555), .ZN(
        n16563) );
  AOI22_X1 U17446 ( .A1(n16560), .A2(n16563), .B1(n8733), .B2(n16559), .ZN(
        P2_U3509) );
  INV_X1 U17447 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n16562) );
  AOI22_X1 U17448 ( .A1(n11936), .A2(n16563), .B1(n16562), .B2(n16561), .ZN(
        P2_U3460) );
  OAI21_X1 U17449 ( .B1(n16593), .B2(n16565), .A(n16564), .ZN(n16566) );
  AOI21_X1 U17450 ( .B1(n16567), .B2(n16597), .A(n16566), .ZN(n16569) );
  AOI22_X1 U17451 ( .A1(n16568), .A2(n16569), .B1(n9944), .B2(n16599), .ZN(
        P3_U3470) );
  INV_X1 U17452 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n16570) );
  AOI22_X1 U17453 ( .A1(n16605), .A2(n16570), .B1(n16569), .B2(n16602), .ZN(
        P3_U3423) );
  AOI21_X1 U17454 ( .B1(n16573), .B2(n16572), .A(n16571), .ZN(n16574) );
  OAI211_X1 U17455 ( .C1(n16577), .C2(n16576), .A(n16575), .B(n16574), .ZN(
        n16578) );
  INV_X1 U17456 ( .A(n16578), .ZN(n16582) );
  AOI22_X1 U17457 ( .A1(n7435), .A2(n16582), .B1(n9403), .B2(n16579), .ZN(
        P1_U3539) );
  INV_X1 U17458 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n16581) );
  AOI22_X1 U17459 ( .A1(n16540), .A2(n16582), .B1(n16581), .B2(n16580), .ZN(
        P1_U3492) );
  OAI22_X1 U17460 ( .A1(n16585), .A2(n16584), .B1(n16593), .B2(n16583), .ZN(
        n16586) );
  AOI211_X1 U17461 ( .C1(n16589), .C2(n16588), .A(n16587), .B(n16586), .ZN(
        n16591) );
  AOI22_X1 U17462 ( .A1(n16601), .A2(n16591), .B1(n16590), .B2(n16599), .ZN(
        P3_U3471) );
  INV_X1 U17463 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n16592) );
  AOI22_X1 U17464 ( .A1(n16605), .A2(n16592), .B1(n16591), .B2(n16602), .ZN(
        P3_U3426) );
  NOR2_X1 U17465 ( .A1(n16594), .A2(n16593), .ZN(n16596) );
  AOI211_X1 U17466 ( .C1(n16598), .C2(n16597), .A(n16596), .B(n16595), .ZN(
        n16603) );
  AOI22_X1 U17467 ( .A1(n16601), .A2(n16603), .B1(n16600), .B2(n16599), .ZN(
        P3_U3472) );
  INV_X1 U17468 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n16604) );
  AOI22_X1 U17469 ( .A1(n16605), .A2(n16604), .B1(n16603), .B2(n16602), .ZN(
        P3_U3429) );
  NAND2_X1 U17470 ( .A1(n16607), .A2(n16606), .ZN(n16608) );
  NAND2_X1 U17471 ( .A1(n16609), .A2(n16608), .ZN(n16613) );
  AOI222_X1 U17472 ( .A1(n16615), .A2(n16614), .B1(n16613), .B2(n16612), .C1(
        n16611), .C2(n16610), .ZN(n16617) );
  OAI211_X1 U17473 ( .C1(n16619), .C2(n16618), .A(n16617), .B(n16616), .ZN(
        P1_U3215) );
  AOI21_X1 U17474 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16620) );
  OAI21_X1 U17475 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16620), 
        .ZN(U28) );
  NAND2_X1 U7558 ( .A1(n16422), .A2(n9300), .ZN(n16435) );
  CLKBUF_X1 U7547 ( .A(n15526), .Z(n7781) );
endmodule

