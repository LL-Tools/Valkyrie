

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, 
        keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, 
        keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, 
        keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, 
        keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, 
        keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, 
        keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, 
        keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, 
        keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, 
        keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, 
        keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597;

  AND2_X1 U2250 ( .A1(n2115), .A2(n2114), .ZN(n3642) );
  OR2_X1 U2251 ( .A1(n3496), .A2(n3490), .ZN(n3497) );
  BUF_X2 U2252 ( .A(n3435), .Z(n3321) );
  NAND2_X1 U2253 ( .A1(n2170), .A2(n3743), .ZN(n2553) );
  NAND3_X1 U2254 ( .A1(n2258), .A2(n2257), .A3(n2256), .ZN(n3543) );
  INV_X2 U2255 ( .A(n3544), .ZN(n2742) );
  CLKBUF_X1 U2256 ( .A(n4253), .Z(n2008) );
  AND2_X1 U2257 ( .A1(n2767), .A2(n2771), .ZN(n2820) );
  INV_X2 U2258 ( .A(n2820), .ZN(n3410) );
  OAI22_X1 U2259 ( .A1(n4300), .A2(n4302), .B1(REG2_REG_13__SCAN_IN), .B2(
        n3897), .ZN(n3898) );
  BUF_X1 U2260 ( .A(n2011), .Z(n3666) );
  OAI22_X1 U2261 ( .A1(n2971), .A2(n2314), .B1(n2973), .B2(n3828), .ZN(n2890)
         );
  INV_X1 U2262 ( .A(n3834), .ZN(n2730) );
  NAND2_X1 U2263 ( .A1(n2630), .A2(IR_REG_31__SCAN_IN), .ZN(n2239) );
  XNOR2_X1 U2264 ( .A(n2239), .B(IR_REG_30__SCAN_IN), .ZN(n4240) );
  AND2_X1 U2265 ( .A1(n2532), .A2(n2458), .ZN(n4247) );
  NAND2_X2 U2266 ( .A1(n3291), .A2(n2423), .ZN(n3356) );
  NAND2_X1 U2267 ( .A1(n2542), .A2(n2551), .ZN(n2767) );
  XNOR2_X1 U2268 ( .A(n2168), .B(IR_REG_1__SCAN_IN), .ZN(n4253) );
  BUF_X4 U2269 ( .A(n2438), .Z(n2012) );
  AND2_X1 U2270 ( .A1(n3320), .A2(n3319), .ZN(n3331) );
  AND2_X1 U2271 ( .A1(n2049), .A2(n2048), .ZN(n4141) );
  NOR2_X1 U2272 ( .A1(n4309), .A2(n2082), .ZN(n3900) );
  NAND2_X1 U2273 ( .A1(n2185), .A2(n2184), .ZN(n3089) );
  INV_X4 U2274 ( .A(n3451), .ZN(n2903) );
  INV_X2 U2275 ( .A(n2551), .ZN(n2583) );
  INV_X1 U2276 ( .A(n3832), .ZN(n3020) );
  NAND4_X2 U2277 ( .A1(n2249), .A2(n2250), .A3(n2248), .A4(n2251), .ZN(n3834)
         );
  NAND4_X1 U2278 ( .A1(n2277), .A2(n2276), .A3(n2275), .A4(n2274), .ZN(n3831)
         );
  CLKBUF_X2 U2279 ( .A(n2285), .Z(n2013) );
  CLKBUF_X2 U2280 ( .A(n2285), .Z(n2014) );
  AND2_X1 U2281 ( .A1(n4240), .A2(n4241), .ZN(n2438) );
  NOR2_X1 U2282 ( .A1(n2101), .A2(n2100), .ZN(n3463) );
  NAND2_X1 U2283 ( .A1(n2129), .A2(n3249), .ZN(n3316) );
  AOI21_X1 U2284 ( .B1(n2176), .B2(n2174), .A(n2173), .ZN(n2466) );
  INV_X1 U2285 ( .A(n2049), .ZN(n4132) );
  NAND2_X1 U2286 ( .A1(n4321), .A2(n3296), .ZN(n4320) );
  XNOR2_X1 U2287 ( .A(n3900), .B(n2421), .ZN(n4321) );
  NAND2_X1 U2288 ( .A1(n3233), .A2(n2400), .ZN(n3343) );
  NAND2_X1 U2289 ( .A1(n3234), .A2(n3711), .ZN(n3233) );
  NAND2_X1 U2290 ( .A1(n4291), .A2(REG2_REG_12__SCAN_IN), .ZN(n4290) );
  AOI21_X1 U2291 ( .B1(n2124), .B2(n2991), .A(n2121), .ZN(n2120) );
  INV_X2 U2292 ( .A(n4263), .ZN(n2009) );
  CLKBUF_X1 U2293 ( .A(n2820), .Z(n3435) );
  AND2_X2 U2294 ( .A1(n2614), .A2(n2542), .ZN(n4421) );
  AND2_X2 U2295 ( .A1(n2767), .A2(n2813), .ZN(n3451) );
  NOR2_X1 U2296 ( .A1(n2849), .A2(n2848), .ZN(n3025) );
  INV_X1 U2297 ( .A(n4247), .ZN(n3908) );
  NAND2_X1 U2298 ( .A1(n2532), .A2(IR_REG_31__SCAN_IN), .ZN(n2534) );
  NAND4_X1 U2299 ( .A1(n2264), .A2(n2263), .A3(n2262), .A4(n2261), .ZN(n3832)
         );
  NAND2_X1 U2300 ( .A1(n2269), .A2(n2268), .ZN(n2848) );
  NAND2_X1 U2301 ( .A1(n2285), .A2(REG1_REG_1__SCAN_IN), .ZN(n2251) );
  INV_X2 U2302 ( .A(n2255), .ZN(n2011) );
  OR2_X1 U2303 ( .A1(n2260), .A2(n2247), .ZN(n2249) );
  CLKBUF_X1 U2304 ( .A(n2260), .Z(n3670) );
  XNOR2_X1 U2305 ( .A(n2588), .B(IR_REG_24__SCAN_IN), .ZN(n4244) );
  NAND2_X1 U2306 ( .A1(n2242), .A2(n2241), .ZN(n2255) );
  OR2_X1 U2307 ( .A1(n2655), .A2(n2231), .ZN(n2095) );
  NAND2_X1 U2308 ( .A1(n2050), .A2(IR_REG_31__SCAN_IN), .ZN(n2655) );
  NOR2_X1 U2309 ( .A1(n2228), .A2(n2227), .ZN(n2015) );
  AND2_X1 U2310 ( .A1(n2350), .A2(n2219), .ZN(n2370) );
  AND2_X1 U2311 ( .A1(n2218), .A2(n2349), .ZN(n2219) );
  AND2_X1 U2312 ( .A1(n2214), .A2(n2301), .ZN(n2172) );
  AND3_X1 U2313 ( .A1(n2044), .A2(n2322), .A3(n2043), .ZN(n2350) );
  AND3_X1 U2314 ( .A1(n2229), .A2(n2594), .A3(n2592), .ZN(n2230) );
  INV_X1 U2315 ( .A(IR_REG_15__SCAN_IN), .ZN(n2430) );
  INV_X1 U2316 ( .A(IR_REG_19__SCAN_IN), .ZN(n4518) );
  INV_X1 U2317 ( .A(IR_REG_23__SCAN_IN), .ZN(n2594) );
  INV_X1 U2318 ( .A(IR_REG_16__SCAN_IN), .ZN(n2428) );
  INV_X1 U2319 ( .A(IR_REG_17__SCAN_IN), .ZN(n2444) );
  NOR2_X1 U2320 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_21__SCAN_IN), .ZN(n2225)
         );
  INV_X1 U2321 ( .A(IR_REG_14__SCAN_IN), .ZN(n2429) );
  NOR2_X1 U2322 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2214)
         );
  AOI21_X2 U2323 ( .B1(n3993), .B2(n2491), .A(n2490), .ZN(n3974) );
  OAI21_X2 U2324 ( .B1(n3089), .B2(n2362), .A(n2361), .ZN(n3181) );
  OAI21_X2 U2325 ( .B1(n3181), .B2(n2210), .A(n2208), .ZN(n3263) );
  INV_X1 U2326 ( .A(n2255), .ZN(n2010) );
  NAND2_X2 U2327 ( .A1(n3555), .A2(n3613), .ZN(n3612) );
  OAI21_X4 U2328 ( .B1(n3633), .B2(n3409), .A(n3408), .ZN(n3555) );
  NOR3_X4 U2329 ( .A1(n3522), .A2(n3438), .A3(n3437), .ZN(n3601) );
  OAI21_X2 U2330 ( .B1(n3522), .B2(n3438), .A(n3437), .ZN(n3602) );
  NAND2_X4 U2331 ( .A1(n2093), .A2(n2232), .ZN(n2265) );
  XNOR2_X2 U2332 ( .A(n2538), .B(n2537), .ZN(n2551) );
  AND2_X1 U2333 ( .A1(n4241), .A2(n2241), .ZN(n2285) );
  XNOR2_X2 U2334 ( .A(n2534), .B(n2533), .ZN(n2542) );
  INV_X1 U2335 ( .A(IR_REG_10__SCAN_IN), .ZN(n2218) );
  INV_X1 U2336 ( .A(IR_REG_27__SCAN_IN), .ZN(n2231) );
  OR2_X1 U2337 ( .A1(n3927), .A2(n3465), .ZN(n3913) );
  OAI21_X1 U2338 ( .B1(n2177), .B2(n2175), .A(n2033), .ZN(n2173) );
  OR2_X1 U2339 ( .A1(n2113), .A2(n2112), .ZN(n2109) );
  AND2_X1 U2340 ( .A1(n3640), .A2(n2114), .ZN(n2113) );
  NOR2_X1 U2341 ( .A1(n2112), .A2(n2111), .ZN(n2110) );
  AND2_X1 U2342 ( .A1(n2769), .A2(n2768), .ZN(n2817) );
  NAND2_X1 U2343 ( .A1(n2035), .A2(n2684), .ZN(n2686) );
  NAND2_X1 U2344 ( .A1(n2682), .A2(REG1_REG_3__SCAN_IN), .ZN(n2035) );
  XNOR2_X1 U2345 ( .A(n2686), .B(n4251), .ZN(n3862) );
  NAND2_X1 U2346 ( .A1(n2041), .A2(n2040), .ZN(n2158) );
  INV_X1 U2347 ( .A(n4275), .ZN(n2040) );
  AOI21_X1 U2348 ( .B1(n2200), .B2(n2198), .A(n2197), .ZN(n2196) );
  INV_X1 U2349 ( .A(n2201), .ZN(n2198) );
  NAND2_X1 U2350 ( .A1(n3820), .A2(n3583), .ZN(n2423) );
  AND4_X1 U2351 ( .A1(n2223), .A2(n2025), .A3(n2015), .A4(n2369), .ZN(n2238)
         );
  NOR2_X1 U2352 ( .A1(n3249), .A2(n2133), .ZN(n2132) );
  INV_X1 U2353 ( .A(n4053), .ZN(n2175) );
  INV_X1 U2354 ( .A(n2076), .ZN(n2071) );
  INV_X1 U2355 ( .A(n3651), .ZN(n2145) );
  AOI21_X1 U2356 ( .B1(n2120), .B2(n2123), .A(n2119), .ZN(n2118) );
  INV_X1 U2357 ( .A(n3059), .ZN(n2119) );
  OR2_X1 U2358 ( .A1(n3197), .A2(n3198), .ZN(n2138) );
  INV_X1 U2359 ( .A(n4241), .ZN(n2242) );
  INV_X1 U2360 ( .A(IR_REG_1__SCAN_IN), .ZN(n2171) );
  AND2_X1 U2361 ( .A1(n4314), .A2(REG2_REG_15__SCAN_IN), .ZN(n2082) );
  AOI21_X1 U2362 ( .B1(n4037), .B2(n3795), .A(n3687), .ZN(n3977) );
  NOR2_X1 U2363 ( .A1(n2179), .A2(n2175), .ZN(n2174) );
  NAND2_X1 U2364 ( .A1(n2080), .A2(n3719), .ZN(n2078) );
  NOR2_X1 U2365 ( .A1(n3787), .A2(n2081), .ZN(n2080) );
  AOI21_X1 U2366 ( .B1(n2181), .B2(n2178), .A(n2024), .ZN(n2177) );
  INV_X1 U2367 ( .A(n2435), .ZN(n2178) );
  INV_X1 U2368 ( .A(n2181), .ZN(n2179) );
  NAND2_X1 U2369 ( .A1(n2211), .A2(n2386), .ZN(n2210) );
  INV_X1 U2370 ( .A(n3765), .ZN(n2088) );
  INV_X1 U2371 ( .A(n3760), .ZN(n2085) );
  AND2_X1 U2372 ( .A1(n2551), .A2(n4245), .ZN(n2642) );
  NAND2_X1 U2373 ( .A1(n3344), .A2(n2045), .ZN(n3293) );
  AND2_X1 U2374 ( .A1(n3657), .A2(n2422), .ZN(n2045) );
  NOR2_X1 U2375 ( .A1(n3552), .A2(n2154), .ZN(n2153) );
  OAI21_X1 U2376 ( .B1(n2109), .B2(n2106), .A(n2031), .ZN(n2105) );
  INV_X1 U2377 ( .A(n3513), .ZN(n2106) );
  NAND2_X1 U2378 ( .A1(n2107), .A2(n2116), .ZN(n2103) );
  AND2_X1 U2379 ( .A1(n3368), .A2(n2145), .ZN(n2144) );
  AND2_X1 U2380 ( .A1(n3579), .A2(n2142), .ZN(n2141) );
  NAND2_X1 U2381 ( .A1(n3383), .A2(n2145), .ZN(n2142) );
  AOI21_X1 U2382 ( .B1(n3458), .B2(n2774), .A(n2773), .ZN(n2775) );
  NAND2_X1 U2383 ( .A1(n2817), .A2(n2772), .ZN(n2778) );
  NAND2_X1 U2384 ( .A1(n2447), .A2(REG3_REG_19__SCAN_IN), .ZN(n2469) );
  AND2_X1 U2385 ( .A1(n3209), .A2(n3208), .ZN(n3250) );
  NAND2_X1 U2386 ( .A1(n3197), .A2(n3198), .ZN(n2136) );
  NOR2_X1 U2387 ( .A1(n3623), .A2(n2151), .ZN(n2150) );
  INV_X1 U2388 ( .A(n3553), .ZN(n2151) );
  NAND2_X1 U2389 ( .A1(n2095), .A2(n2094), .ZN(n2093) );
  INV_X1 U2390 ( .A(n3568), .ZN(n2114) );
  NAND3_X1 U2391 ( .A1(n4244), .A2(n4243), .A3(n2627), .ZN(n2771) );
  AND2_X1 U2392 ( .A1(n2012), .A2(REG3_REG_0__SCAN_IN), .ZN(n2254) );
  INV_X1 U2393 ( .A(IR_REG_3__SCAN_IN), .ZN(n2279) );
  NAND2_X1 U2394 ( .A1(n2055), .A2(n2693), .ZN(n2694) );
  NAND2_X1 U2395 ( .A1(n2690), .A2(REG2_REG_3__SCAN_IN), .ZN(n2055) );
  XNOR2_X1 U2396 ( .A(n2694), .B(n2054), .ZN(n2695) );
  INV_X1 U2397 ( .A(n4251), .ZN(n2054) );
  OAI21_X1 U2398 ( .B1(n2748), .B2(n2747), .A(n2749), .ZN(n2801) );
  OR2_X1 U2399 ( .A1(n4264), .A2(n3875), .ZN(n2041) );
  NOR2_X1 U2400 ( .A1(n3877), .A2(n4285), .ZN(n4296) );
  INV_X1 U2401 ( .A(n2156), .ZN(n3876) );
  OR2_X1 U2402 ( .A1(n4296), .A2(n4295), .ZN(n2037) );
  NAND2_X1 U2403 ( .A1(n4280), .A2(n3893), .ZN(n3895) );
  NOR2_X1 U2404 ( .A1(n4306), .A2(n2167), .ZN(n3882) );
  AND2_X1 U2405 ( .A1(n4314), .A2(REG1_REG_15__SCAN_IN), .ZN(n2167) );
  OR2_X1 U2406 ( .A1(n2163), .A2(n4342), .ZN(n2039) );
  NOR2_X1 U2407 ( .A1(n2199), .A2(n2194), .ZN(n2193) );
  INV_X1 U2408 ( .A(n2504), .ZN(n2194) );
  INV_X1 U2409 ( .A(n2200), .ZN(n2199) );
  NOR2_X1 U2410 ( .A1(n2523), .A2(n2202), .ZN(n2201) );
  INV_X1 U2411 ( .A(n2514), .ZN(n2202) );
  AOI21_X1 U2412 ( .B1(n2201), .B2(n2515), .A(n2203), .ZN(n2200) );
  NOR2_X1 U2413 ( .A1(n3644), .A2(n3515), .ZN(n2203) );
  INV_X1 U2414 ( .A(n3728), .ZN(n3478) );
  INV_X1 U2415 ( .A(n3481), .ZN(n3966) );
  NAND2_X1 U2416 ( .A1(n2492), .A2(REG3_REG_24__SCAN_IN), .ZN(n2498) );
  NOR2_X1 U2417 ( .A1(n4069), .A2(n4045), .ZN(n2053) );
  AND2_X1 U2418 ( .A1(n4055), .A2(n4039), .ZN(n2476) );
  AND2_X1 U2419 ( .A1(n4108), .A2(n3596), .ZN(n2434) );
  AND2_X1 U2420 ( .A1(n4111), .A2(n2182), .ZN(n2181) );
  INV_X1 U2421 ( .A(n2434), .ZN(n2182) );
  NAND2_X1 U2422 ( .A1(n3356), .A2(n2435), .ZN(n2183) );
  AND2_X1 U2423 ( .A1(n3581), .A2(n3657), .ZN(n2190) );
  NAND2_X1 U2424 ( .A1(n2063), .A2(n2061), .ZN(n3682) );
  AND2_X1 U2425 ( .A1(n2062), .A2(n3779), .ZN(n2061) );
  NAND2_X1 U2426 ( .A1(n2065), .A2(n2068), .ZN(n2062) );
  NOR2_X1 U2427 ( .A1(n2388), .A2(n2191), .ZN(n3234) );
  AND2_X1 U2428 ( .A1(n3268), .A2(n3822), .ZN(n2191) );
  AOI21_X1 U2429 ( .B1(n3336), .B2(n3276), .A(n3263), .ZN(n2388) );
  NAND2_X1 U2430 ( .A1(n2064), .A2(n3781), .ZN(n3266) );
  NAND2_X1 U2431 ( .A1(n3179), .A2(n3775), .ZN(n2064) );
  NAND2_X1 U2432 ( .A1(n2563), .A2(n3766), .ZN(n3085) );
  OR2_X1 U2433 ( .A1(n3047), .A2(n3772), .ZN(n2563) );
  AOI21_X1 U2434 ( .B1(n2016), .B2(n2189), .A(n2023), .ZN(n2184) );
  AND2_X1 U2435 ( .A1(n2560), .A2(n3760), .ZN(n3757) );
  AND2_X1 U2436 ( .A1(n2205), .A2(n2304), .ZN(n2204) );
  AOI21_X1 U2437 ( .B1(n2738), .B2(n2553), .A(n2215), .ZN(n2839) );
  NAND2_X1 U2438 ( .A1(n4092), .A2(n4067), .ZN(n4069) );
  AND2_X1 U2439 ( .A1(n3274), .A2(n3235), .ZN(n3344) );
  NOR2_X2 U2440 ( .A1(n3153), .A2(n3268), .ZN(n3274) );
  AND2_X1 U2441 ( .A1(n2771), .A2(n4374), .ZN(n2787) );
  NOR2_X1 U2442 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2220)
         );
  INV_X1 U2443 ( .A(n3824), .ZN(n3212) );
  INV_X1 U2444 ( .A(n3360), .ZN(n3596) );
  INV_X1 U2445 ( .A(n3182), .ZN(n3189) );
  OR2_X1 U2446 ( .A1(n2265), .A2(n2267), .ZN(n2269) );
  NAND2_X1 U2447 ( .A1(n2265), .A2(DATAI_2_), .ZN(n2268) );
  INV_X1 U2448 ( .A(n3373), .ZN(n3657) );
  NAND2_X1 U2449 ( .A1(n2531), .A2(n2530), .ZN(n3927) );
  OAI21_X1 U2450 ( .B1(n3862), .B2(n2685), .A(n2687), .ZN(n2710) );
  XNOR2_X1 U2451 ( .A(n2715), .B(n2057), .ZN(n2714) );
  XNOR2_X1 U2452 ( .A(n3895), .B(n4384), .ZN(n4291) );
  NOR2_X1 U2453 ( .A1(n4286), .A2(n4287), .ZN(n4285) );
  XNOR2_X1 U2454 ( .A(n3882), .B(n2421), .ZN(n4324) );
  NAND2_X1 U2455 ( .A1(n4324), .A2(n4323), .ZN(n4322) );
  NAND2_X1 U2456 ( .A1(n4334), .A2(n4335), .ZN(n4333) );
  INV_X1 U2457 ( .A(n2039), .ZN(n4341) );
  INV_X1 U2458 ( .A(n2162), .ZN(n2161) );
  AOI21_X1 U2459 ( .B1(n2163), .B2(n4342), .A(n4433), .ZN(n2162) );
  AOI21_X1 U2460 ( .B1(n4442), .B2(ADDR_REG_18__SCAN_IN), .A(n4343), .ZN(n2160) );
  AND2_X1 U2461 ( .A1(n2672), .A2(n2665), .ZN(n4348) );
  NAND2_X1 U2462 ( .A1(n2186), .A2(n2187), .ZN(n3046) );
  OR2_X1 U2463 ( .A1(n2889), .A2(n2189), .ZN(n2186) );
  INV_X1 U2464 ( .A(n3754), .ZN(n2074) );
  INV_X1 U2465 ( .A(n3762), .ZN(n2070) );
  INV_X1 U2466 ( .A(n2032), .ZN(n2112) );
  NOR2_X1 U2467 ( .A1(n2132), .A2(n2128), .ZN(n2127) );
  INV_X1 U2468 ( .A(n2138), .ZN(n2128) );
  OR2_X1 U2469 ( .A1(n2132), .A2(n2134), .ZN(n2126) );
  NOR2_X1 U2470 ( .A1(n3250), .A2(n2135), .ZN(n2134) );
  NAND2_X1 U2471 ( .A1(n2136), .A2(n3317), .ZN(n2135) );
  OR2_X1 U2472 ( .A1(n2498), .A2(n3571), .ZN(n2506) );
  INV_X1 U2473 ( .A(n3781), .ZN(n2068) );
  AND2_X1 U2474 ( .A1(n3776), .A2(n2066), .ZN(n2065) );
  NAND2_X1 U2475 ( .A1(n3781), .A2(n2067), .ZN(n2066) );
  INV_X1 U2476 ( .A(n3775), .ZN(n2067) );
  OAI21_X1 U2477 ( .B1(n3016), .B2(n2072), .A(n2069), .ZN(n2972) );
  INV_X1 U2478 ( .A(n2073), .ZN(n2072) );
  AOI21_X1 U2479 ( .B1(n2071), .B2(n2073), .A(n2070), .ZN(n2069) );
  NOR2_X1 U2480 ( .A1(n2933), .A2(n2074), .ZN(n2073) );
  NOR2_X1 U2481 ( .A1(n2557), .A2(n2077), .ZN(n2076) );
  INV_X1 U2482 ( .A(n3750), .ZN(n2077) );
  INV_X1 U2483 ( .A(n2848), .ZN(n2270) );
  NAND2_X1 U2484 ( .A1(n3020), .A2(n2848), .ZN(n3745) );
  NOR2_X1 U2485 ( .A1(n3968), .A2(n3943), .ZN(n3471) );
  OR2_X1 U2486 ( .A1(n3188), .A2(n3214), .ZN(n3153) );
  NAND2_X1 U2487 ( .A1(n2052), .A2(n3048), .ZN(n3052) );
  INV_X1 U2488 ( .A(n3003), .ZN(n2884) );
  INV_X1 U2489 ( .A(n3018), .ZN(n3024) );
  INV_X1 U2490 ( .A(n2635), .ZN(n2760) );
  INV_X1 U2491 ( .A(IR_REG_6__SCAN_IN), .ZN(n2349) );
  INV_X1 U2492 ( .A(IR_REG_9__SCAN_IN), .ZN(n2044) );
  NOR2_X1 U2493 ( .A1(n2957), .A2(n2122), .ZN(n2121) );
  NAND2_X1 U2494 ( .A1(n3124), .A2(n3123), .ZN(n2099) );
  AND2_X1 U2495 ( .A1(n3396), .A2(n3395), .ZN(n3534) );
  OR2_X1 U2496 ( .A1(n2315), .A2(n4576), .ZN(n2329) );
  INV_X1 U2497 ( .A(n3822), .ZN(n3336) );
  OAI21_X1 U2498 ( .B1(n2265), .B2(n4504), .A(n2259), .ZN(n2774) );
  NAND2_X1 U2499 ( .A1(n3612), .A2(n2153), .ZN(n2152) );
  NAND2_X1 U2500 ( .A1(n2353), .A2(REG3_REG_10__SCAN_IN), .ZN(n2363) );
  INV_X1 U2501 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4484) );
  INV_X1 U2502 ( .A(n2831), .ZN(n2098) );
  INV_X1 U2503 ( .A(n2833), .ZN(n2097) );
  NOR2_X1 U2504 ( .A1(n2413), .A2(n2412), .ZN(n2436) );
  NAND2_X1 U2505 ( .A1(n2307), .A2(REG3_REG_6__SCAN_IN), .ZN(n2315) );
  NAND2_X1 U2506 ( .A1(n3369), .A2(n2030), .ZN(n3649) );
  OR2_X1 U2507 ( .A1(n2401), .A2(n3656), .ZN(n2413) );
  AND2_X1 U2508 ( .A1(n2522), .A2(n2521), .ZN(n3644) );
  XNOR2_X1 U2509 ( .A(n2692), .B(n2678), .ZN(n2690) );
  OR2_X1 U2510 ( .A1(n2703), .A2(n2702), .ZN(n2060) );
  NAND2_X1 U2511 ( .A1(n2060), .A2(n2059), .ZN(n2058) );
  NAND2_X1 U2512 ( .A1(n4250), .A2(REG2_REG_5__SCAN_IN), .ZN(n2059) );
  AOI21_X1 U2513 ( .B1(n2721), .B2(REG2_REG_6__SCAN_IN), .A(n2056), .ZN(n2723)
         );
  AND2_X1 U2514 ( .A1(n2058), .A2(n2720), .ZN(n2056) );
  OR2_X1 U2515 ( .A1(n2807), .A2(n2806), .ZN(n2166) );
  INV_X1 U2516 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2800) );
  AND2_X1 U2517 ( .A1(n2166), .A2(n2165), .ZN(n3874) );
  NAND2_X1 U2518 ( .A1(n3873), .A2(REG1_REG_9__SCAN_IN), .ZN(n2165) );
  NAND2_X1 U2519 ( .A1(n2158), .A2(n2157), .ZN(n2156) );
  NAND2_X1 U2520 ( .A1(n3888), .A2(REG1_REG_11__SCAN_IN), .ZN(n2157) );
  XNOR2_X1 U2521 ( .A(n3879), .B(n4444), .ZN(n4435) );
  AND2_X1 U2522 ( .A1(n2037), .A2(n2036), .ZN(n3879) );
  NAND2_X1 U2523 ( .A1(n3897), .A2(REG1_REG_13__SCAN_IN), .ZN(n2036) );
  NOR2_X1 U2524 ( .A1(n4435), .A2(n4436), .ZN(n4434) );
  NAND2_X1 U2525 ( .A1(n4320), .A2(n3901), .ZN(n4331) );
  NAND2_X1 U2526 ( .A1(n4333), .A2(n2164), .ZN(n2163) );
  NAND2_X1 U2527 ( .A1(n4378), .A2(n4186), .ZN(n2164) );
  NAND2_X1 U2528 ( .A1(n3472), .A2(n2047), .ZN(n2049) );
  NOR2_X1 U2529 ( .A1(n3934), .A2(n3926), .ZN(n2047) );
  OR2_X1 U2530 ( .A1(n2524), .A2(n3464), .ZN(n2546) );
  NAND2_X1 U2531 ( .A1(n3476), .A2(n3674), .ZN(n3916) );
  NAND2_X1 U2532 ( .A1(n3945), .A2(n4109), .ZN(n2090) );
  NOR2_X1 U2533 ( .A1(n2485), .A2(n3526), .ZN(n2492) );
  INV_X1 U2534 ( .A(n3986), .ZN(n3981) );
  OR2_X1 U2535 ( .A1(n4040), .A2(n4030), .ZN(n2484) );
  OR2_X1 U2536 ( .A1(n2469), .A2(n2468), .ZN(n2478) );
  OR2_X1 U2537 ( .A1(n2478), .A2(n4485), .ZN(n2485) );
  AND2_X1 U2538 ( .A1(n4042), .A2(n3731), .ZN(n2464) );
  INV_X1 U2539 ( .A(n4002), .ZN(n4040) );
  INV_X1 U2540 ( .A(n2080), .ZN(n2079) );
  NAND2_X1 U2541 ( .A1(n3298), .A2(n2080), .ZN(n4057) );
  OAI21_X1 U2542 ( .B1(n3356), .B2(n2179), .A(n2177), .ZN(n4075) );
  NAND2_X1 U2543 ( .A1(n3298), .A2(n3683), .ZN(n4079) );
  NAND2_X1 U2544 ( .A1(n3300), .A2(n3299), .ZN(n3298) );
  OR2_X1 U2545 ( .A1(n3349), .A2(n3716), .ZN(n3347) );
  NAND2_X1 U2546 ( .A1(n2399), .A2(n3235), .ZN(n2400) );
  INV_X1 U2547 ( .A(n2209), .ZN(n2208) );
  OAI21_X1 U2548 ( .B1(n2210), .B2(n2372), .A(n2387), .ZN(n2209) );
  OR2_X1 U2549 ( .A1(n3214), .A2(n3823), .ZN(n2387) );
  AND2_X1 U2550 ( .A1(n2376), .A2(REG3_REG_13__SCAN_IN), .ZN(n2389) );
  INV_X1 U2551 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2373) );
  NAND2_X1 U2552 ( .A1(n2564), .A2(n3771), .ZN(n3179) );
  AOI21_X1 U2553 ( .B1(n2338), .B2(n2188), .A(n2018), .ZN(n2187) );
  INV_X1 U2554 ( .A(n2327), .ZN(n2188) );
  AOI21_X1 U2555 ( .B1(n2087), .B2(n2085), .A(n2084), .ZN(n2083) );
  INV_X1 U2556 ( .A(n2087), .ZN(n2086) );
  INV_X1 U2557 ( .A(n3759), .ZN(n2084) );
  INV_X1 U2558 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2704) );
  NAND2_X1 U2559 ( .A1(n2075), .A2(n3754), .ZN(n2935) );
  NAND2_X1 U2560 ( .A1(n3016), .A2(n2076), .ZN(n2075) );
  INV_X1 U2561 ( .A(n3830), .ZN(n2937) );
  NAND2_X1 U2562 ( .A1(n3025), .A2(n3024), .ZN(n3496) );
  NAND2_X1 U2563 ( .A1(n3016), .A2(n3750), .ZN(n3489) );
  NAND2_X1 U2564 ( .A1(n2169), .A2(n2842), .ZN(n2843) );
  INV_X1 U2565 ( .A(n2555), .ZN(n2169) );
  OR2_X1 U2566 ( .A1(n2553), .A2(n3741), .ZN(n2841) );
  AND2_X1 U2567 ( .A1(n2780), .A2(n2787), .ZN(n2881) );
  INV_X1 U2568 ( .A(n4025), .ZN(n4101) );
  NAND2_X1 U2569 ( .A1(n3472), .A2(n3465), .ZN(n3933) );
  OR2_X1 U2570 ( .A1(n3985), .A2(n2503), .ZN(n3968) );
  NAND2_X1 U2571 ( .A1(n4007), .A2(n3986), .ZN(n3985) );
  NOR2_X1 U2572 ( .A1(n4164), .A2(n4006), .ZN(n4007) );
  INV_X1 U2573 ( .A(n3527), .ZN(n4006) );
  INV_X1 U2574 ( .A(n2053), .ZN(n4047) );
  NOR2_X2 U2575 ( .A1(n2046), .A2(n2034), .ZN(n4092) );
  NAND2_X1 U2576 ( .A1(n3190), .A2(n3189), .ZN(n3188) );
  INV_X1 U2577 ( .A(n2052), .ZN(n3053) );
  INV_X1 U2578 ( .A(n4410), .ZN(n4416) );
  NAND2_X1 U2579 ( .A1(n2792), .A2(n2742), .ZN(n2849) );
  INV_X1 U2580 ( .A(IR_REG_28__SCAN_IN), .ZN(n2544) );
  INV_X1 U2581 ( .A(IR_REG_26__SCAN_IN), .ZN(n2051) );
  NOR2_X1 U2582 ( .A1(n2539), .A2(IR_REG_22__SCAN_IN), .ZN(n2586) );
  INV_X1 U2583 ( .A(IR_REG_20__SCAN_IN), .ZN(n2533) );
  NOR2_X1 U2584 ( .A1(n2346), .A2(n2585), .ZN(n2321) );
  OAI21_X1 U2585 ( .B1(n2958), .B2(n2123), .A(n2120), .ZN(n3060) );
  INV_X1 U2586 ( .A(n3480), .ZN(n3515) );
  NAND2_X1 U2587 ( .A1(n2104), .A2(n2109), .ZN(n3514) );
  NAND2_X1 U2588 ( .A1(n3566), .A2(n2110), .ZN(n2104) );
  NOR2_X1 U2589 ( .A1(n2155), .A2(n2149), .ZN(n2148) );
  NOR2_X1 U2590 ( .A1(n2155), .A2(n2150), .ZN(n2147) );
  INV_X1 U2591 ( .A(n2153), .ZN(n2149) );
  INV_X1 U2592 ( .A(n3400), .ZN(n4090) );
  INV_X1 U2593 ( .A(n2105), .ZN(n2102) );
  INV_X1 U2594 ( .A(n2562), .ZN(n3081) );
  INV_X1 U2595 ( .A(n4039), .ZN(n4045) );
  NAND2_X1 U2596 ( .A1(n2137), .A2(n2136), .ZN(n3251) );
  INV_X1 U2597 ( .A(n2558), .ZN(n2941) );
  AOI21_X1 U2598 ( .B1(n2141), .B2(n2143), .A(n3384), .ZN(n2139) );
  INV_X1 U2599 ( .A(n2141), .ZN(n2140) );
  NOR2_X1 U2600 ( .A1(n2030), .A2(n2144), .ZN(n2143) );
  INV_X1 U2601 ( .A(n2774), .ZN(n2792) );
  NAND2_X1 U2602 ( .A1(n2265), .A2(DATAI_20_), .ZN(n4067) );
  NAND2_X1 U2603 ( .A1(n2137), .A2(n2130), .ZN(n2129) );
  NOR2_X1 U2604 ( .A1(n3250), .A2(n2131), .ZN(n2130) );
  INV_X1 U2605 ( .A(n2136), .ZN(n2131) );
  NAND2_X1 U2606 ( .A1(n2152), .A2(n3553), .ZN(n3622) );
  NAND2_X1 U2607 ( .A1(n2958), .A2(n2957), .ZN(n2993) );
  NAND2_X1 U2608 ( .A1(n3566), .A2(n3567), .ZN(n2115) );
  NAND3_X1 U2609 ( .A1(n2857), .A2(n2856), .A3(n3818), .ZN(n3661) );
  INV_X1 U2610 ( .A(n3644), .ZN(n3945) );
  OAI21_X1 U2611 ( .B1(n3643), .B2(n2513), .A(n2512), .ZN(n3481) );
  OAI211_X1 U2612 ( .C1(n3987), .C2(n2513), .A(n2495), .B(n2494), .ZN(n4001)
         );
  NAND4_X1 U2613 ( .A1(n2453), .A2(n2452), .A3(n2451), .A4(n2450), .ZN(n4063)
         );
  NAND2_X1 U2614 ( .A1(n2438), .A2(REG3_REG_1__SCAN_IN), .ZN(n2250) );
  NOR2_X1 U2615 ( .A1(n2254), .A2(n2253), .ZN(n2258) );
  NAND2_X1 U2616 ( .A1(n3835), .A2(n3843), .ZN(n3853) );
  XNOR2_X1 U2617 ( .A(n2683), .B(n2678), .ZN(n2682) );
  AND2_X1 U2618 ( .A1(n2291), .A2(n2281), .ZN(n2691) );
  INV_X1 U2619 ( .A(n2695), .ZN(n3860) );
  INV_X1 U2620 ( .A(n2060), .ZN(n2701) );
  XNOR2_X1 U2621 ( .A(n2058), .B(n2057), .ZN(n2721) );
  NAND2_X1 U2622 ( .A1(n2042), .A2(n2716), .ZN(n2748) );
  NAND2_X1 U2623 ( .A1(n2714), .A2(REG1_REG_6__SCAN_IN), .ZN(n2042) );
  INV_X1 U2624 ( .A(n2166), .ZN(n3872) );
  XNOR2_X1 U2625 ( .A(n3874), .B(n4273), .ZN(n4265) );
  INV_X1 U2626 ( .A(n2041), .ZN(n4276) );
  INV_X1 U2627 ( .A(n2158), .ZN(n4274) );
  XNOR2_X1 U2628 ( .A(n2156), .B(n3894), .ZN(n4286) );
  INV_X1 U2629 ( .A(n2037), .ZN(n4294) );
  NAND2_X1 U2630 ( .A1(n4290), .A2(n3896), .ZN(n4302) );
  AND2_X1 U2631 ( .A1(n2410), .A2(n2419), .ZN(n4314) );
  NAND2_X1 U2632 ( .A1(n4322), .A2(n3883), .ZN(n4334) );
  AND2_X1 U2633 ( .A1(n2672), .A2(n3844), .ZN(n4337) );
  INV_X1 U2634 ( .A(n4337), .ZN(n4433) );
  AND2_X1 U2635 ( .A1(n2039), .A2(n2038), .ZN(n3885) );
  NAND2_X1 U2636 ( .A1(n3903), .A2(REG1_REG_18__SCAN_IN), .ZN(n2038) );
  NAND2_X1 U2637 ( .A1(n2192), .A2(n2196), .ZN(n3929) );
  NAND2_X1 U2638 ( .A1(n2195), .A2(n2200), .ZN(n3925) );
  NAND2_X1 U2639 ( .A1(n3938), .A2(n2201), .ZN(n2195) );
  AOI21_X1 U2640 ( .B1(n2092), .B2(n4032), .A(n2089), .ZN(n3505) );
  NAND2_X1 U2641 ( .A1(n2091), .A2(n2090), .ZN(n2089) );
  XNOR2_X1 U2642 ( .A(n3916), .B(n2197), .ZN(n2092) );
  INV_X1 U2643 ( .A(n2582), .ZN(n2091) );
  OAI21_X1 U2644 ( .B1(n3938), .B2(n2515), .A(n2514), .ZN(n3470) );
  NAND2_X1 U2645 ( .A1(n2053), .A2(n4030), .ZN(n4164) );
  NAND2_X1 U2646 ( .A1(n2183), .A2(n2181), .ZN(n4110) );
  NOR2_X1 U2647 ( .A1(n2180), .A2(n2434), .ZN(n4112) );
  INV_X1 U2648 ( .A(n2183), .ZN(n2180) );
  NAND2_X1 U2649 ( .A1(n3344), .A2(n3657), .ZN(n3294) );
  NAND2_X1 U2650 ( .A1(n3180), .A2(n2372), .ZN(n3152) );
  INV_X1 U2651 ( .A(n3757), .ZN(n2325) );
  AND2_X1 U2652 ( .A1(n4263), .A2(n3908), .ZN(n4116) );
  NAND2_X1 U2653 ( .A1(n3486), .A2(n2293), .ZN(n2934) );
  AND2_X1 U2654 ( .A1(n4116), .A2(n4421), .ZN(n4358) );
  INV_X1 U2655 ( .A(n4358), .ZN(n4095) );
  NAND2_X1 U2656 ( .A1(n4402), .A2(n2788), .ZN(n4352) );
  OR2_X1 U2657 ( .A1(n2616), .A2(n2880), .ZN(n4430) );
  INV_X2 U2658 ( .A(n4422), .ZN(n4423) );
  NOR2_X1 U2659 ( .A1(IR_REG_29__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .ZN(n2237)
         );
  NAND2_X1 U2660 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .ZN(n2234) );
  XNOR2_X1 U2661 ( .A(n2590), .B(IR_REG_26__SCAN_IN), .ZN(n4243) );
  AND2_X1 U2662 ( .A1(n2644), .A2(STATE_REG_SCAN_IN), .ZN(n4374) );
  INV_X1 U2663 ( .A(n2552), .ZN(n4245) );
  INV_X1 U2664 ( .A(IR_REG_21__SCAN_IN), .ZN(n2537) );
  INV_X1 U2665 ( .A(n3897), .ZN(n4383) );
  XNOR2_X1 U2666 ( .A(n2292), .B(IR_REG_4__SCAN_IN), .ZN(n4251) );
  OAI21_X1 U2667 ( .B1(IR_REG_1__SCAN_IN), .B2(IR_REG_0__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2266) );
  NAND2_X1 U2668 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2168)
         );
  INV_X1 U2669 ( .A(n2159), .ZN(n4350) );
  OAI21_X1 U2670 ( .B1(n4341), .B2(n2161), .A(n2160), .ZN(n2159) );
  AOI21_X1 U2671 ( .B1(n3369), .B2(n3368), .A(n3383), .ZN(n3578) );
  AND2_X1 U2672 ( .A1(n2187), .A2(n2020), .ZN(n2016) );
  AND2_X1 U2673 ( .A1(n3751), .A2(n3754), .ZN(n2017) );
  INV_X1 U2674 ( .A(n2992), .ZN(n2122) );
  INV_X1 U2675 ( .A(n3924), .ZN(n2197) );
  AND2_X1 U2676 ( .A1(n3827), .A2(n3081), .ZN(n2018) );
  AND2_X1 U2677 ( .A1(n2152), .A2(n2150), .ZN(n2019) );
  NAND2_X1 U2678 ( .A1(n2222), .A2(n2214), .ZN(n2300) );
  NAND2_X1 U2679 ( .A1(n3826), .A2(n3118), .ZN(n2020) );
  AND2_X1 U2680 ( .A1(n3136), .A2(n3128), .ZN(n2021) );
  NOR2_X1 U2681 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2022)
         );
  AND2_X1 U2682 ( .A1(n3138), .A2(n3048), .ZN(n2023) );
  NOR2_X1 U2683 ( .A1(n4087), .A2(n4113), .ZN(n2024) );
  AOI21_X1 U2684 ( .B1(n3612), .B2(n2148), .A(n2147), .ZN(n2146) );
  XNOR2_X1 U2685 ( .A(n2814), .B(n2903), .ZN(n2863) );
  AND2_X1 U2686 ( .A1(n2026), .A2(n2022), .ZN(n2025) );
  AND2_X1 U2687 ( .A1(n2230), .A2(n2207), .ZN(n2026) );
  AND2_X1 U2688 ( .A1(n3685), .A2(n2078), .ZN(n2027) );
  AND2_X1 U2689 ( .A1(n2804), .A2(n4248), .ZN(n2028) );
  AND2_X1 U2690 ( .A1(n2369), .A2(n2051), .ZN(n2029) );
  INV_X1 U2691 ( .A(n2108), .ZN(n2107) );
  NAND2_X1 U2692 ( .A1(n2110), .A2(n3513), .ZN(n2108) );
  CLKBUF_X3 U2693 ( .A(n3459), .Z(n3203) );
  CLKBUF_X3 U2694 ( .A(n2824), .Z(n3459) );
  INV_X1 U2695 ( .A(n2720), .ZN(n2057) );
  INV_X1 U2696 ( .A(n3317), .ZN(n2133) );
  AND2_X1 U2697 ( .A1(n3383), .A2(n3368), .ZN(n2030) );
  INV_X1 U2698 ( .A(n3683), .ZN(n2081) );
  INV_X1 U2699 ( .A(IR_REG_8__SCAN_IN), .ZN(n2043) );
  INV_X1 U2700 ( .A(IR_REG_22__SCAN_IN), .ZN(n2207) );
  INV_X1 U2701 ( .A(n3567), .ZN(n2111) );
  NAND2_X1 U2702 ( .A1(n2223), .A2(n2369), .ZN(n2396) );
  NAND2_X1 U2703 ( .A1(n3455), .A2(n3456), .ZN(n2031) );
  OR2_X1 U2704 ( .A1(n3293), .A2(n3596), .ZN(n2046) );
  INV_X1 U2705 ( .A(n2212), .ZN(n3180) );
  NAND2_X1 U2706 ( .A1(n3450), .A2(n3449), .ZN(n2032) );
  INV_X1 U2707 ( .A(n3604), .ZN(n2116) );
  NAND2_X1 U2708 ( .A1(n4102), .A2(n4090), .ZN(n2033) );
  NOR2_X1 U2709 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2345)
         );
  OR2_X1 U2710 ( .A1(n3400), .A2(n4113), .ZN(n2034) );
  OR2_X1 U2711 ( .A1(n4421), .A2(n3410), .ZN(n3424) );
  INV_X1 U2712 ( .A(n3894), .ZN(n4384) );
  AND2_X1 U2713 ( .A1(n2583), .A2(n2552), .ZN(n2614) );
  OR2_X1 U2714 ( .A1(n3487), .A2(n2017), .ZN(n3486) );
  NAND2_X1 U2715 ( .A1(n2099), .A2(n2021), .ZN(n3168) );
  NAND2_X1 U2716 ( .A1(n2099), .A2(n3128), .ZN(n3134) );
  OR2_X1 U2717 ( .A1(n2238), .A2(n2585), .ZN(n2543) );
  AND2_X1 U2718 ( .A1(n2581), .A2(n2580), .ZN(n4104) );
  INV_X1 U2719 ( .A(n4104), .ZN(n4032) );
  NAND2_X1 U2720 ( .A1(n2265), .A2(DATAI_22_), .ZN(n4030) );
  INV_X1 U2721 ( .A(IR_REG_2__SCAN_IN), .ZN(n2221) );
  INV_X1 U2722 ( .A(IR_REG_29__SCAN_IN), .ZN(n2235) );
  INV_X1 U2723 ( .A(IR_REG_31__SCAN_IN), .ZN(n2585) );
  NOR2_X1 U2724 ( .A1(n2803), .A2(n2028), .ZN(n2807) );
  INV_X1 U2725 ( .A(n2046), .ZN(n4114) );
  NAND2_X1 U2726 ( .A1(n3933), .A2(n3934), .ZN(n2048) );
  AND2_X2 U2727 ( .A1(n3471), .A2(n3515), .ZN(n3472) );
  NAND4_X1 U2728 ( .A1(n2026), .A2(n2015), .A3(n2223), .A4(n2369), .ZN(n2589)
         );
  NAND4_X1 U2729 ( .A1(n2029), .A2(n2026), .A3(n2223), .A4(n2015), .ZN(n2050)
         );
  NAND3_X1 U2730 ( .A1(n2015), .A2(n2369), .A3(n2223), .ZN(n2539) );
  NOR2_X2 U2731 ( .A1(n3052), .A2(n3140), .ZN(n3190) );
  NOR2_X2 U2732 ( .A1(n3038), .A2(n3081), .ZN(n2052) );
  NAND2_X1 U2733 ( .A1(n3179), .A2(n2065), .ZN(n2063) );
  OAI21_X1 U2734 ( .B1(n3300), .B2(n2079), .A(n2027), .ZN(n2574) );
  OAI21_X1 U2735 ( .B1(n2876), .B2(n2086), .A(n2083), .ZN(n3047) );
  OAI21_X1 U2736 ( .B1(n2876), .B2(n2561), .A(n3760), .ZN(n3032) );
  AOI21_X1 U2737 ( .B1(n2561), .B2(n3760), .A(n2088), .ZN(n2087) );
  NAND2_X1 U2738 ( .A1(n2574), .A2(n3790), .ZN(n4037) );
  AOI21_X1 U2739 ( .B1(n3958), .B2(n3796), .A(n3802), .ZN(n3477) );
  NOR2_X1 U2740 ( .A1(n3977), .A2(n3798), .ZN(n3958) );
  NAND2_X1 U2741 ( .A1(n2559), .A2(n3756), .ZN(n2876) );
  AOI21_X1 U2742 ( .B1(n3903), .B2(REG2_REG_18__SCAN_IN), .A(n4344), .ZN(n3905) );
  NOR2_X1 U2743 ( .A1(n3899), .A2(n4438), .ZN(n4311) );
  OAI21_X1 U2744 ( .B1(n3055), .B2(n3890), .A(n3889), .ZN(n3891) );
  NAND2_X1 U2745 ( .A1(n2555), .A2(n3721), .ZN(n2844) );
  NAND2_X1 U2746 ( .A1(n2010), .A2(REG0_REG_1__SCAN_IN), .ZN(n2248) );
  NAND2_X1 U2747 ( .A1(n2568), .A2(n3677), .ZN(n3349) );
  AND2_X2 U2748 ( .A1(n2370), .A2(n2220), .ZN(n2223) );
  MUX2_X1 U2749 ( .A(n2008), .B(DATAI_1_), .S(n2265), .Z(n3544) );
  NAND2_X1 U2750 ( .A1(n2655), .A2(n2544), .ZN(n2094) );
  OAI21_X1 U2751 ( .B1(n2831), .B2(n2833), .A(n2867), .ZN(n2096) );
  NAND2_X1 U2752 ( .A1(n2096), .A2(n2894), .ZN(n2900) );
  NAND2_X1 U2753 ( .A1(n2868), .A2(n2867), .ZN(n2895) );
  NAND2_X1 U2754 ( .A1(n2098), .A2(n2097), .ZN(n2868) );
  OAI21_X1 U2755 ( .B1(n3601), .B2(n3604), .A(n3602), .ZN(n3566) );
  NOR2_X1 U2756 ( .A1(n3602), .A2(n2108), .ZN(n2100) );
  OAI21_X1 U2757 ( .B1(n3601), .B2(n2103), .A(n2102), .ZN(n2101) );
  NAND2_X1 U2758 ( .A1(n2958), .A2(n2120), .ZN(n2117) );
  NAND2_X1 U2759 ( .A1(n2118), .A2(n2117), .ZN(n3065) );
  NOR2_X1 U2760 ( .A1(n2991), .A2(n2992), .ZN(n2123) );
  NAND2_X1 U2761 ( .A1(n2957), .A2(n2122), .ZN(n2124) );
  NAND2_X1 U2762 ( .A1(n3199), .A2(n2138), .ZN(n2137) );
  NAND2_X1 U2763 ( .A1(n2125), .A2(n2126), .ZN(n3315) );
  NAND2_X1 U2764 ( .A1(n3199), .A2(n2127), .ZN(n2125) );
  OAI21_X2 U2765 ( .B1(n3369), .B2(n2140), .A(n2139), .ZN(n3592) );
  INV_X1 U2766 ( .A(n2146), .ZN(n3522) );
  NAND2_X1 U2767 ( .A1(n3612), .A2(n3615), .ZN(n3559) );
  INV_X1 U2768 ( .A(n3615), .ZN(n2154) );
  OR2_X1 U2769 ( .A1(n3523), .A2(n3524), .ZN(n2155) );
  XNOR2_X2 U2770 ( .A(n2236), .B(n2235), .ZN(n4241) );
  NAND2_X1 U2771 ( .A1(n2730), .A2(n3544), .ZN(n2170) );
  NAND3_X1 U2772 ( .A1(n3746), .A2(n3745), .A3(n2170), .ZN(n3749) );
  NAND2_X1 U2773 ( .A1(n2841), .A2(n2170), .ZN(n2555) );
  NAND3_X1 U2774 ( .A1(n4504), .A2(n2171), .A3(n2221), .ZN(n2278) );
  NAND2_X1 U2775 ( .A1(n3834), .A2(n3458), .ZN(n2822) );
  AND2_X4 U2776 ( .A1(n2222), .A2(n2172), .ZN(n2369) );
  INV_X1 U2777 ( .A(n3356), .ZN(n2176) );
  NAND2_X1 U2778 ( .A1(n2889), .A2(n2016), .ZN(n2185) );
  NAND2_X1 U2779 ( .A1(n2889), .A2(n2327), .ZN(n3031) );
  INV_X1 U2780 ( .A(n2338), .ZN(n2189) );
  AOI21_X2 U2781 ( .B1(n3343), .B2(n2411), .A(n2190), .ZN(n3292) );
  NAND2_X1 U2782 ( .A1(n2505), .A2(n2504), .ZN(n3938) );
  NAND2_X1 U2783 ( .A1(n2505), .A2(n2193), .ZN(n2192) );
  NAND2_X1 U2784 ( .A1(n2206), .A2(n2204), .ZN(n2306) );
  NAND2_X1 U2785 ( .A1(n2017), .A2(n2293), .ZN(n2205) );
  NAND2_X1 U2786 ( .A1(n3487), .A2(n2293), .ZN(n2206) );
  NAND2_X1 U2787 ( .A1(n3720), .A2(n2372), .ZN(n2211) );
  NOR2_X1 U2788 ( .A1(n3181), .A2(n3720), .ZN(n2212) );
  MUX2_X2 U2789 ( .A(REG0_REG_28__SCAN_IN), .B(n2617), .S(n4423), .Z(n2618) );
  MUX2_X2 U2790 ( .A(REG1_REG_28__SCAN_IN), .B(n2617), .S(n4432), .Z(n2613) );
  AND2_X1 U2791 ( .A1(n2369), .A2(n2349), .ZN(n2346) );
  INV_X1 U2792 ( .A(n3820), .ZN(n3653) );
  OAI211_X1 U2793 ( .C1(n3570), .C2(n2513), .A(n2502), .B(n2501), .ZN(n3944)
         );
  OR2_X1 U2794 ( .A1(n3944), .A2(n2503), .ZN(n2213) );
  INV_X1 U2795 ( .A(n3338), .ZN(n3235) );
  AND2_X1 U2796 ( .A1(n3834), .A2(n3544), .ZN(n2215) );
  INV_X1 U2797 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2412) );
  OR2_X1 U2798 ( .A1(n3508), .A2(n4236), .ZN(n2216) );
  OR2_X1 U2799 ( .A1(n3508), .A2(n4188), .ZN(n2217) );
  NAND2_X1 U2800 ( .A1(n3168), .A2(n3167), .ZN(n3199) );
  NAND4_X1 U2801 ( .A1(n2381), .A2(n2380), .A3(n2379), .A4(n2378), .ZN(n3823)
         );
  INV_X1 U2802 ( .A(n2771), .ZN(n2854) );
  INV_X1 U2803 ( .A(IR_REG_13__SCAN_IN), .ZN(n2226) );
  AND2_X1 U2804 ( .A1(n3729), .A2(n3939), .ZN(n3796) );
  AND2_X1 U2805 ( .A1(n3264), .A2(n2565), .ZN(n3776) );
  INV_X1 U2806 ( .A(IR_REG_24__SCAN_IN), .ZN(n2229) );
  INV_X1 U2807 ( .A(n2767), .ZN(n2766) );
  AND2_X1 U2808 ( .A1(n3407), .A2(n3532), .ZN(n3408) );
  INV_X1 U2809 ( .A(n3135), .ZN(n3136) );
  CLKBUF_X3 U2810 ( .A(n3458), .Z(n3444) );
  INV_X1 U2811 ( .A(n3572), .ZN(n2503) );
  NAND2_X1 U2812 ( .A1(n3823), .A2(n3214), .ZN(n2386) );
  INV_X1 U2813 ( .A(n2842), .ZN(n3721) );
  NAND2_X1 U2814 ( .A1(n2265), .A2(DATAI_0_), .ZN(n2259) );
  INV_X1 U2815 ( .A(IR_REG_18__SCAN_IN), .ZN(n2455) );
  INV_X1 U2816 ( .A(n2949), .ZN(n2907) );
  NOR2_X1 U2817 ( .A1(n2506), .A2(n4479), .ZN(n2516) );
  NAND2_X1 U2818 ( .A1(n3927), .A2(n3926), .ZN(n3928) );
  NAND2_X1 U2819 ( .A1(n3944), .A2(n2503), .ZN(n2504) );
  AND2_X1 U2820 ( .A1(n4026), .A2(n4006), .ZN(n2490) );
  INV_X1 U2821 ( .A(n3352), .ZN(n2399) );
  NAND2_X1 U2822 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2294) );
  INV_X1 U2823 ( .A(n3276), .ZN(n3268) );
  INV_X1 U2824 ( .A(n2973), .ZN(n2980) );
  INV_X1 U2825 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4576) );
  NAND2_X1 U2826 ( .A1(n2389), .A2(REG3_REG_14__SCAN_IN), .ZN(n2401) );
  INV_X1 U2827 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2328) );
  NOR2_X1 U2828 ( .A1(n2374), .A2(n2373), .ZN(n2376) );
  NOR2_X1 U2829 ( .A1(n2339), .A2(n2800), .ZN(n2353) );
  OR2_X1 U2830 ( .A1(n2363), .A2(n4484), .ZN(n2374) );
  AND2_X1 U2831 ( .A1(n2436), .A2(n4589), .ZN(n2447) );
  OR2_X1 U2832 ( .A1(n2507), .A2(n2516), .ZN(n3643) );
  NOR2_X1 U2833 ( .A1(n2750), .A2(n4453), .ZN(n2803) );
  AND2_X1 U2834 ( .A1(n2614), .A2(n4246), .ZN(n4127) );
  INV_X1 U2835 ( .A(n3930), .ZN(n3931) );
  INV_X1 U2836 ( .A(n4030), .ZN(n4017) );
  INV_X1 U2837 ( .A(n4063), .ZN(n4102) );
  INV_X1 U2838 ( .A(n3821), .ZN(n3581) );
  AND2_X1 U2839 ( .A1(n3781), .A2(n3775), .ZN(n3720) );
  NOR2_X1 U2840 ( .A1(n2294), .A2(n2704), .ZN(n2307) );
  INV_X1 U2841 ( .A(n4127), .ZN(n4134) );
  INV_X1 U2842 ( .A(IR_REG_25__SCAN_IN), .ZN(n2592) );
  OR2_X1 U2843 ( .A1(n2371), .A2(n2585), .ZN(n2383) );
  AND2_X1 U2844 ( .A1(n2524), .A2(n2517), .ZN(n3519) );
  AND2_X1 U2845 ( .A1(n2546), .A2(n2525), .ZN(n3506) );
  OR2_X1 U2846 ( .A1(n2329), .A2(n2328), .ZN(n2339) );
  INV_X1 U2847 ( .A(n3149), .ZN(n3214) );
  INV_X1 U2848 ( .A(n3658), .ZN(n3636) );
  NAND4_X1 U2849 ( .A1(n2395), .A2(n2394), .A3(n2393), .A4(n2392), .ZN(n3352)
         );
  AND2_X1 U2850 ( .A1(n2352), .A2(n2359), .ZN(n3873) );
  AND2_X1 U2851 ( .A1(n2672), .A2(n2791), .ZN(n4315) );
  INV_X1 U2852 ( .A(n2546), .ZN(n3923) );
  AND2_X1 U2853 ( .A1(n4254), .A2(n2642), .ZN(n4109) );
  AND2_X1 U2854 ( .A1(n4263), .A2(n2891), .ZN(n4121) );
  INV_X1 U2855 ( .A(n4352), .ZN(n4367) );
  AND2_X1 U2856 ( .A1(n4363), .A2(n2552), .ZN(n4402) );
  INV_X1 U2857 ( .A(n2691), .ZN(n2678) );
  AND2_X1 U2858 ( .A1(n2647), .A2(n2659), .ZN(n4442) );
  OR2_X1 U2859 ( .A1(n2790), .A2(n2765), .ZN(n3664) );
  AOI21_X1 U2860 ( .B1(n3923), .B2(n2012), .A(n2550), .ZN(n3699) );
  NAND4_X1 U2861 ( .A1(n2463), .A2(n2462), .A3(n2461), .A4(n2460), .ZN(n4042)
         );
  NAND4_X1 U2862 ( .A1(n2246), .A2(n2245), .A3(n2244), .A4(n2243), .ZN(n3822)
         );
  INV_X1 U2863 ( .A(n4315), .ZN(n4445) );
  INV_X1 U2864 ( .A(n4121), .ZN(n4098) );
  NAND2_X1 U2865 ( .A1(n4432), .A2(n4421), .ZN(n4188) );
  INV_X2 U2866 ( .A(n4430), .ZN(n4432) );
  NAND2_X1 U2867 ( .A1(n4423), .A2(n4421), .ZN(n4236) );
  OR2_X1 U2868 ( .A1(n2616), .A2(n2761), .ZN(n4422) );
  INV_X1 U2869 ( .A(n3902), .ZN(n4378) );
  AND2_X1 U2870 ( .A1(n2324), .A2(n2335), .ZN(n4249) );
  INV_X1 U2871 ( .A(n3833), .ZN(U4043) );
  INV_X1 U2872 ( .A(n2278), .ZN(n2222) );
  NAND2_X1 U2873 ( .A1(n2396), .A2(IR_REG_31__SCAN_IN), .ZN(n2224) );
  XNOR2_X1 U2874 ( .A(n2224), .B(IR_REG_13__SCAN_IN), .ZN(n3897) );
  INV_X1 U2875 ( .A(DATAI_13_), .ZN(n2233) );
  NAND4_X1 U2876 ( .A1(n2225), .A2(n4518), .A3(n2429), .A4(n2455), .ZN(n2228)
         );
  NAND4_X1 U2877 ( .A1(n2430), .A2(n2226), .A3(n2444), .A4(n2428), .ZN(n2227)
         );
  NAND2_X1 U2878 ( .A1(n2544), .A2(IR_REG_27__SCAN_IN), .ZN(n2232) );
  MUX2_X1 U2879 ( .A(n4383), .B(n2233), .S(n2265), .Z(n3276) );
  NAND2_X1 U2880 ( .A1(n2543), .A2(n2234), .ZN(n2236) );
  NAND2_X1 U2881 ( .A1(n2238), .A2(n2237), .ZN(n2630) );
  INV_X1 U2882 ( .A(n4240), .ZN(n2241) );
  NAND2_X1 U2883 ( .A1(n2013), .A2(REG1_REG_13__SCAN_IN), .ZN(n2246) );
  NOR2_X1 U2884 ( .A1(n2376), .A2(REG3_REG_13__SCAN_IN), .ZN(n2240) );
  OR2_X1 U2885 ( .A1(n2389), .A2(n2240), .ZN(n3278) );
  INV_X1 U2886 ( .A(n3278), .ZN(n3260) );
  NAND2_X1 U2887 ( .A1(n2012), .A2(n3260), .ZN(n2245) );
  NAND2_X1 U2888 ( .A1(n2011), .A2(REG0_REG_13__SCAN_IN), .ZN(n2244) );
  NAND2_X2 U2889 ( .A1(n2242), .A2(n4240), .ZN(n2260) );
  INV_X1 U2890 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3279) );
  OR2_X1 U2891 ( .A1(n2260), .A2(n3279), .ZN(n2243) );
  INV_X1 U2892 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2247) );
  NAND2_X1 U2893 ( .A1(n3834), .A2(n2742), .ZN(n3743) );
  INV_X1 U2894 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2252) );
  NOR2_X1 U2895 ( .A1(n2260), .A2(n2252), .ZN(n2253) );
  NAND2_X1 U2896 ( .A1(n2014), .A2(REG1_REG_0__SCAN_IN), .ZN(n2257) );
  NAND2_X1 U2897 ( .A1(n2011), .A2(REG0_REG_0__SCAN_IN), .ZN(n2256) );
  AND2_X1 U2898 ( .A1(n3543), .A2(n2774), .ZN(n2738) );
  NAND2_X1 U2899 ( .A1(n2012), .A2(REG3_REG_2__SCAN_IN), .ZN(n2264) );
  NAND2_X1 U2900 ( .A1(n2011), .A2(REG0_REG_2__SCAN_IN), .ZN(n2263) );
  NAND2_X1 U2901 ( .A1(n2013), .A2(REG1_REG_2__SCAN_IN), .ZN(n2262) );
  INV_X1 U2902 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2928) );
  OR2_X1 U2903 ( .A1(n2260), .A2(n2928), .ZN(n2261) );
  XNOR2_X2 U2904 ( .A(n2266), .B(IR_REG_2__SCAN_IN), .ZN(n4252) );
  INV_X1 U2905 ( .A(n4252), .ZN(n2267) );
  NAND2_X1 U2906 ( .A1(n3832), .A2(n2270), .ZN(n3748) );
  NAND2_X1 U2907 ( .A1(n3748), .A2(n3745), .ZN(n2842) );
  NAND2_X1 U2908 ( .A1(n2839), .A2(n2842), .ZN(n2838) );
  NAND2_X1 U2909 ( .A1(n3020), .A2(n2270), .ZN(n2271) );
  NAND2_X1 U2910 ( .A1(n2838), .A2(n2271), .ZN(n3015) );
  NAND2_X1 U2911 ( .A1(n2013), .A2(REG1_REG_3__SCAN_IN), .ZN(n2277) );
  INV_X1 U2912 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2272) );
  NAND2_X1 U2913 ( .A1(n2012), .A2(n2272), .ZN(n2276) );
  NAND2_X1 U2914 ( .A1(n2011), .A2(REG0_REG_3__SCAN_IN), .ZN(n2275) );
  INV_X1 U2915 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2273) );
  OR2_X1 U2916 ( .A1(n2260), .A2(n2273), .ZN(n2274) );
  NAND2_X1 U2917 ( .A1(n2278), .A2(IR_REG_31__SCAN_IN), .ZN(n2280) );
  NAND2_X1 U2918 ( .A1(n2280), .A2(n2279), .ZN(n2291) );
  OR2_X1 U2919 ( .A1(n2280), .A2(n2279), .ZN(n2281) );
  MUX2_X1 U2920 ( .A(n2691), .B(DATAI_3_), .S(n2265), .Z(n3018) );
  NAND2_X1 U2921 ( .A1(n3831), .A2(n3018), .ZN(n2282) );
  NAND2_X1 U2922 ( .A1(n3015), .A2(n2282), .ZN(n2284) );
  INV_X1 U2923 ( .A(n3831), .ZN(n2556) );
  NAND2_X1 U2924 ( .A1(n2556), .A2(n3024), .ZN(n2283) );
  NAND2_X1 U2925 ( .A1(n2284), .A2(n2283), .ZN(n3487) );
  NAND2_X1 U2926 ( .A1(n2014), .A2(REG1_REG_4__SCAN_IN), .ZN(n2290) );
  OAI21_X1 U2927 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2294), .ZN(n3500) );
  INV_X1 U2928 ( .A(n3500), .ZN(n2952) );
  NAND2_X1 U2929 ( .A1(n2012), .A2(n2952), .ZN(n2289) );
  NAND2_X1 U2930 ( .A1(n2011), .A2(REG0_REG_4__SCAN_IN), .ZN(n2288) );
  INV_X1 U2931 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2286) );
  OR2_X1 U2932 ( .A1(n2260), .A2(n2286), .ZN(n2287) );
  NAND4_X1 U2933 ( .A1(n2290), .A2(n2289), .A3(n2288), .A4(n2287), .ZN(n3830)
         );
  NAND2_X1 U2934 ( .A1(n2291), .A2(IR_REG_31__SCAN_IN), .ZN(n2292) );
  MUX2_X1 U2935 ( .A(n4251), .B(DATAI_4_), .S(n2265), .Z(n3490) );
  NAND2_X1 U2936 ( .A1(n2937), .A2(n3490), .ZN(n3751) );
  INV_X1 U2937 ( .A(n3490), .ZN(n3498) );
  NAND2_X1 U2938 ( .A1(n3830), .A2(n3498), .ZN(n3754) );
  NAND2_X1 U2939 ( .A1(n3830), .A2(n3490), .ZN(n2293) );
  NAND2_X1 U2940 ( .A1(n2014), .A2(REG1_REG_5__SCAN_IN), .ZN(n2299) );
  AND2_X1 U2941 ( .A1(n2294), .A2(n2704), .ZN(n2295) );
  NOR2_X1 U2942 ( .A1(n2307), .A2(n2295), .ZN(n2942) );
  NAND2_X1 U2943 ( .A1(n2012), .A2(n2942), .ZN(n2298) );
  NAND2_X1 U2944 ( .A1(n3666), .A2(REG0_REG_5__SCAN_IN), .ZN(n2297) );
  INV_X1 U2945 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2940) );
  OR2_X1 U2946 ( .A1(n2260), .A2(n2940), .ZN(n2296) );
  NAND4_X1 U2947 ( .A1(n2299), .A2(n2298), .A3(n2297), .A4(n2296), .ZN(n3829)
         );
  INV_X1 U2948 ( .A(n3829), .ZN(n2965) );
  NAND2_X1 U2949 ( .A1(n2300), .A2(IR_REG_31__SCAN_IN), .ZN(n2302) );
  INV_X1 U2950 ( .A(IR_REG_5__SCAN_IN), .ZN(n2301) );
  XNOR2_X1 U2951 ( .A(n2302), .B(n2301), .ZN(n2706) );
  INV_X1 U2952 ( .A(DATAI_5_), .ZN(n2303) );
  MUX2_X1 U2953 ( .A(n2706), .B(n2303), .S(n2265), .Z(n2558) );
  NAND2_X1 U2954 ( .A1(n2965), .A2(n2558), .ZN(n2304) );
  NAND2_X1 U2955 ( .A1(n3829), .A2(n2941), .ZN(n2305) );
  NAND2_X1 U2956 ( .A1(n2306), .A2(n2305), .ZN(n2971) );
  NAND2_X1 U2957 ( .A1(n2014), .A2(REG1_REG_6__SCAN_IN), .ZN(n2312) );
  OR2_X1 U2958 ( .A1(n2307), .A2(REG3_REG_6__SCAN_IN), .ZN(n2308) );
  AND2_X1 U2959 ( .A1(n2315), .A2(n2308), .ZN(n4351) );
  NAND2_X1 U2960 ( .A1(n2012), .A2(n4351), .ZN(n2311) );
  NAND2_X1 U2961 ( .A1(n2011), .A2(REG0_REG_6__SCAN_IN), .ZN(n2310) );
  INV_X1 U2962 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4354) );
  OR2_X1 U2963 ( .A1(n3670), .A2(n4354), .ZN(n2309) );
  NAND4_X1 U2964 ( .A1(n2312), .A2(n2311), .A3(n2310), .A4(n2309), .ZN(n3828)
         );
  OR2_X1 U2965 ( .A1(n2369), .A2(n2585), .ZN(n2313) );
  XNOR2_X1 U2966 ( .A(n2313), .B(IR_REG_6__SCAN_IN), .ZN(n2720) );
  MUX2_X1 U2967 ( .A(n2720), .B(DATAI_6_), .S(n2265), .Z(n2973) );
  AND2_X1 U2968 ( .A1(n3828), .A2(n2973), .ZN(n2314) );
  INV_X1 U2969 ( .A(n2890), .ZN(n2326) );
  NAND2_X1 U2970 ( .A1(n2014), .A2(REG1_REG_7__SCAN_IN), .ZN(n2320) );
  NAND2_X1 U2971 ( .A1(n2315), .A2(n4576), .ZN(n2316) );
  AND2_X1 U2972 ( .A1(n2329), .A2(n2316), .ZN(n3004) );
  NAND2_X1 U2973 ( .A1(n2012), .A2(n3004), .ZN(n2319) );
  NAND2_X1 U2974 ( .A1(n2011), .A2(REG0_REG_7__SCAN_IN), .ZN(n2318) );
  OR2_X1 U2975 ( .A1(n2260), .A2(n2886), .ZN(n2317) );
  NAND4_X1 U2976 ( .A1(n2320), .A2(n2319), .A3(n2318), .A4(n2317), .ZN(n2997)
         );
  INV_X1 U2977 ( .A(n2997), .ZN(n3078) );
  NAND2_X1 U2978 ( .A1(n2321), .A2(IR_REG_7__SCAN_IN), .ZN(n2324) );
  INV_X1 U2979 ( .A(n2321), .ZN(n2323) );
  INV_X1 U2980 ( .A(IR_REG_7__SCAN_IN), .ZN(n2322) );
  NAND2_X1 U2981 ( .A1(n2323), .A2(n2322), .ZN(n2335) );
  MUX2_X1 U2982 ( .A(n4249), .B(DATAI_7_), .S(n2265), .Z(n3003) );
  NAND2_X1 U2983 ( .A1(n3078), .A2(n3003), .ZN(n2560) );
  NAND2_X1 U2984 ( .A1(n2997), .A2(n2884), .ZN(n3760) );
  NAND2_X1 U2985 ( .A1(n2326), .A2(n2325), .ZN(n2889) );
  NAND2_X1 U2986 ( .A1(n2997), .A2(n3003), .ZN(n2327) );
  NAND2_X1 U2987 ( .A1(n2013), .A2(REG1_REG_8__SCAN_IN), .ZN(n2334) );
  NAND2_X1 U2988 ( .A1(n2329), .A2(n2328), .ZN(n2330) );
  NAND2_X1 U2989 ( .A1(n2339), .A2(n2330), .ZN(n3084) );
  INV_X1 U2990 ( .A(n3084), .ZN(n3040) );
  NAND2_X1 U2991 ( .A1(n2012), .A2(n3040), .ZN(n2333) );
  NAND2_X1 U2992 ( .A1(n2011), .A2(REG0_REG_8__SCAN_IN), .ZN(n2332) );
  INV_X1 U2993 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2796) );
  OR2_X1 U2994 ( .A1(n2260), .A2(n2796), .ZN(n2331) );
  NAND4_X1 U2995 ( .A1(n2334), .A2(n2333), .A3(n2332), .A4(n2331), .ZN(n3827)
         );
  INV_X1 U2996 ( .A(n3827), .ZN(n3115) );
  NAND2_X1 U2997 ( .A1(n2335), .A2(IR_REG_31__SCAN_IN), .ZN(n2336) );
  XNOR2_X1 U2998 ( .A(n2336), .B(n2043), .ZN(n2802) );
  INV_X1 U2999 ( .A(DATAI_8_), .ZN(n2337) );
  MUX2_X1 U3000 ( .A(n2802), .B(n2337), .S(n2265), .Z(n2562) );
  NAND2_X1 U3001 ( .A1(n3115), .A2(n2562), .ZN(n2338) );
  NAND2_X1 U3002 ( .A1(n2014), .A2(REG1_REG_9__SCAN_IN), .ZN(n2344) );
  AND2_X1 U3003 ( .A1(n2339), .A2(n2800), .ZN(n2340) );
  NOR2_X1 U3004 ( .A1(n2353), .A2(n2340), .ZN(n3119) );
  NAND2_X1 U3005 ( .A1(n2012), .A2(n3119), .ZN(n2343) );
  NAND2_X1 U3006 ( .A1(n2011), .A2(REG0_REG_9__SCAN_IN), .ZN(n2342) );
  INV_X1 U3007 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3055) );
  OR2_X1 U3008 ( .A1(n2260), .A2(n3055), .ZN(n2341) );
  NAND4_X1 U3009 ( .A1(n2344), .A2(n2343), .A3(n2342), .A4(n2341), .ZN(n3826)
         );
  NAND2_X1 U3010 ( .A1(n2346), .A2(n2345), .ZN(n2347) );
  NAND2_X1 U3011 ( .A1(n2347), .A2(IR_REG_31__SCAN_IN), .ZN(n2348) );
  MUX2_X1 U3012 ( .A(IR_REG_31__SCAN_IN), .B(n2348), .S(IR_REG_9__SCAN_IN), 
        .Z(n2352) );
  AND2_X1 U3013 ( .A1(n2350), .A2(n2349), .ZN(n2351) );
  NAND2_X1 U3014 ( .A1(n2369), .A2(n2351), .ZN(n2359) );
  MUX2_X1 U3015 ( .A(n3873), .B(DATAI_9_), .S(n2265), .Z(n3118) );
  INV_X1 U3016 ( .A(n3826), .ZN(n3138) );
  INV_X1 U3017 ( .A(n3118), .ZN(n3048) );
  NAND2_X1 U3018 ( .A1(n2014), .A2(REG1_REG_10__SCAN_IN), .ZN(n2358) );
  OR2_X1 U3019 ( .A1(n2353), .A2(REG3_REG_10__SCAN_IN), .ZN(n2354) );
  AND2_X1 U3020 ( .A1(n2354), .A2(n2363), .ZN(n3093) );
  NAND2_X1 U3021 ( .A1(n2012), .A2(n3093), .ZN(n2357) );
  NAND2_X1 U3022 ( .A1(n2011), .A2(REG0_REG_10__SCAN_IN), .ZN(n2356) );
  INV_X1 U3023 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3094) );
  OR2_X1 U3024 ( .A1(n2260), .A2(n3094), .ZN(n2355) );
  NAND4_X1 U3025 ( .A1(n2358), .A2(n2357), .A3(n2356), .A4(n2355), .ZN(n3825)
         );
  NAND2_X1 U3026 ( .A1(n2359), .A2(IR_REG_31__SCAN_IN), .ZN(n2360) );
  XNOR2_X1 U3027 ( .A(n2360), .B(IR_REG_10__SCAN_IN), .ZN(n4386) );
  MUX2_X1 U3028 ( .A(n4386), .B(DATAI_10_), .S(n2265), .Z(n3140) );
  NOR2_X1 U3029 ( .A1(n3825), .A2(n3140), .ZN(n2362) );
  NAND2_X1 U3030 ( .A1(n3825), .A2(n3140), .ZN(n2361) );
  NAND2_X1 U3031 ( .A1(n2013), .A2(REG1_REG_11__SCAN_IN), .ZN(n2368) );
  NAND2_X1 U3032 ( .A1(n2363), .A2(n4484), .ZN(n2364) );
  AND2_X1 U3033 ( .A1(n2374), .A2(n2364), .ZN(n3191) );
  NAND2_X1 U3034 ( .A1(n2012), .A2(n3191), .ZN(n2367) );
  NAND2_X1 U3035 ( .A1(n2011), .A2(REG0_REG_11__SCAN_IN), .ZN(n2366) );
  INV_X1 U3036 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3193) );
  OR2_X1 U3037 ( .A1(n2260), .A2(n3193), .ZN(n2365) );
  NAND4_X1 U3038 ( .A1(n2368), .A2(n2367), .A3(n2366), .A4(n2365), .ZN(n3824)
         );
  AND2_X1 U3039 ( .A1(n2370), .A2(n2369), .ZN(n2371) );
  XNOR2_X1 U3040 ( .A(n2383), .B(IR_REG_11__SCAN_IN), .ZN(n3888) );
  MUX2_X1 U3041 ( .A(n3888), .B(DATAI_11_), .S(n2265), .Z(n3182) );
  NAND2_X1 U3042 ( .A1(n3212), .A2(n3182), .ZN(n3781) );
  NAND2_X1 U3043 ( .A1(n3824), .A2(n3189), .ZN(n3775) );
  NAND2_X1 U3044 ( .A1(n3212), .A2(n3189), .ZN(n2372) );
  NAND2_X1 U3045 ( .A1(n2014), .A2(REG1_REG_12__SCAN_IN), .ZN(n2381) );
  AND2_X1 U3046 ( .A1(n2374), .A2(n2373), .ZN(n2375) );
  NOR2_X1 U3047 ( .A1(n2376), .A2(n2375), .ZN(n3215) );
  NAND2_X1 U3048 ( .A1(n2012), .A2(n3215), .ZN(n2380) );
  NAND2_X1 U3049 ( .A1(n2011), .A2(REG0_REG_12__SCAN_IN), .ZN(n2379) );
  INV_X1 U3050 ( .A(REG2_REG_12__SCAN_IN), .ZN(n2377) );
  OR2_X1 U3051 ( .A1(n2260), .A2(n2377), .ZN(n2378) );
  INV_X1 U3052 ( .A(n3823), .ZN(n3270) );
  INV_X1 U3053 ( .A(IR_REG_11__SCAN_IN), .ZN(n2382) );
  NAND2_X1 U3054 ( .A1(n2383), .A2(n2382), .ZN(n2384) );
  NAND2_X1 U3055 ( .A1(n2384), .A2(IR_REG_31__SCAN_IN), .ZN(n2385) );
  XNOR2_X1 U3056 ( .A(n2385), .B(IR_REG_12__SCAN_IN), .ZN(n3894) );
  INV_X1 U3057 ( .A(DATAI_12_), .ZN(n4577) );
  MUX2_X1 U3058 ( .A(n4384), .B(n4577), .S(n2265), .Z(n3149) );
  NAND2_X1 U3059 ( .A1(n2014), .A2(REG1_REG_14__SCAN_IN), .ZN(n2395) );
  OR2_X1 U3060 ( .A1(n2389), .A2(REG3_REG_14__SCAN_IN), .ZN(n2390) );
  AND2_X1 U3061 ( .A1(n2401), .A2(n2390), .ZN(n3339) );
  NAND2_X1 U3062 ( .A1(n2012), .A2(n3339), .ZN(n2394) );
  NAND2_X1 U3063 ( .A1(n2011), .A2(REG0_REG_14__SCAN_IN), .ZN(n2393) );
  INV_X1 U3064 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2391) );
  OR2_X1 U3065 ( .A1(n2260), .A2(n2391), .ZN(n2392) );
  INV_X1 U3066 ( .A(n2396), .ZN(n2397) );
  NAND2_X1 U3067 ( .A1(n2397), .A2(n2226), .ZN(n2432) );
  NAND2_X1 U3068 ( .A1(n2432), .A2(IR_REG_31__SCAN_IN), .ZN(n2398) );
  XNOR2_X1 U3069 ( .A(n2398), .B(IR_REG_14__SCAN_IN), .ZN(n4381) );
  MUX2_X1 U3070 ( .A(n4381), .B(DATAI_14_), .S(n2265), .Z(n3338) );
  NAND2_X1 U3071 ( .A1(n2399), .A2(n3338), .ZN(n3677) );
  NAND2_X1 U3072 ( .A1(n3352), .A2(n3235), .ZN(n3678) );
  NAND2_X1 U3073 ( .A1(n3677), .A2(n3678), .ZN(n3711) );
  NAND2_X1 U3074 ( .A1(n2014), .A2(REG1_REG_15__SCAN_IN), .ZN(n2406) );
  INV_X1 U3075 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3656) );
  NAND2_X1 U3076 ( .A1(n2401), .A2(n3656), .ZN(n2402) );
  AND2_X1 U3077 ( .A1(n2413), .A2(n2402), .ZN(n3662) );
  NAND2_X1 U3078 ( .A1(n2012), .A2(n3662), .ZN(n2405) );
  NAND2_X1 U3079 ( .A1(n2011), .A2(REG0_REG_15__SCAN_IN), .ZN(n2404) );
  INV_X1 U3080 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3346) );
  OR2_X1 U3081 ( .A1(n2260), .A2(n3346), .ZN(n2403) );
  NAND4_X1 U3082 ( .A1(n2406), .A2(n2405), .A3(n2404), .A4(n2403), .ZN(n3821)
         );
  OR2_X1 U3083 ( .A1(n2432), .A2(IR_REG_14__SCAN_IN), .ZN(n2407) );
  NAND2_X1 U3084 ( .A1(n2407), .A2(IR_REG_31__SCAN_IN), .ZN(n2409) );
  INV_X1 U3085 ( .A(n2409), .ZN(n2408) );
  NAND2_X1 U3086 ( .A1(n2408), .A2(IR_REG_15__SCAN_IN), .ZN(n2410) );
  NAND2_X1 U3087 ( .A1(n2409), .A2(n2430), .ZN(n2419) );
  MUX2_X1 U3088 ( .A(n4314), .B(DATAI_15_), .S(n2265), .Z(n3373) );
  NAND2_X1 U3089 ( .A1(n3821), .A2(n3373), .ZN(n2411) );
  NAND2_X1 U3090 ( .A1(n2013), .A2(REG1_REG_16__SCAN_IN), .ZN(n2418) );
  AND2_X1 U3091 ( .A1(n2413), .A2(n2412), .ZN(n2414) );
  NOR2_X1 U3092 ( .A1(n2436), .A2(n2414), .ZN(n3584) );
  NAND2_X1 U3093 ( .A1(n2012), .A2(n3584), .ZN(n2417) );
  NAND2_X1 U3094 ( .A1(n3666), .A2(REG0_REG_16__SCAN_IN), .ZN(n2416) );
  INV_X1 U3095 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3296) );
  OR2_X1 U3096 ( .A1(n3670), .A2(n3296), .ZN(n2415) );
  NAND4_X1 U3097 ( .A1(n2418), .A2(n2417), .A3(n2416), .A4(n2415), .ZN(n3820)
         );
  NAND2_X1 U3098 ( .A1(n2419), .A2(IR_REG_31__SCAN_IN), .ZN(n2420) );
  XNOR2_X1 U3099 ( .A(n2420), .B(n2428), .ZN(n4379) );
  INV_X1 U3100 ( .A(n4379), .ZN(n2421) );
  MUX2_X1 U3101 ( .A(n2421), .B(DATAI_16_), .S(n2265), .Z(n3583) );
  NAND2_X1 U3102 ( .A1(n3653), .A2(n3583), .ZN(n3788) );
  INV_X1 U3103 ( .A(n3583), .ZN(n2422) );
  NAND2_X1 U3104 ( .A1(n3820), .A2(n2422), .ZN(n3683) );
  NAND2_X1 U3105 ( .A1(n3788), .A2(n3683), .ZN(n3719) );
  NAND2_X1 U3106 ( .A1(n3292), .A2(n3719), .ZN(n3291) );
  NAND2_X1 U3107 ( .A1(n2014), .A2(REG1_REG_17__SCAN_IN), .ZN(n2427) );
  INV_X1 U3108 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3593) );
  XNOR2_X1 U3109 ( .A(n2436), .B(n3593), .ZN(n3597) );
  NAND2_X1 U3110 ( .A1(n2012), .A2(n3597), .ZN(n2426) );
  NAND2_X1 U3111 ( .A1(n3666), .A2(REG0_REG_17__SCAN_IN), .ZN(n2425) );
  INV_X1 U3112 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3363) );
  OR2_X1 U3113 ( .A1(n3670), .A2(n3363), .ZN(n2424) );
  NAND4_X1 U3114 ( .A1(n2427), .A2(n2426), .A3(n2425), .A4(n2424), .ZN(n4108)
         );
  INV_X1 U3115 ( .A(n4108), .ZN(n3634) );
  NAND3_X1 U3116 ( .A1(n2430), .A2(n2429), .A3(n2428), .ZN(n2431) );
  NOR2_X2 U3117 ( .A1(n2432), .A2(n2431), .ZN(n2445) );
  OR2_X1 U3118 ( .A1(n2445), .A2(n2585), .ZN(n2433) );
  XNOR2_X1 U3119 ( .A(n2433), .B(IR_REG_17__SCAN_IN), .ZN(n3902) );
  INV_X1 U3120 ( .A(DATAI_17_), .ZN(n4377) );
  MUX2_X1 U3121 ( .A(n4378), .B(n4377), .S(n2265), .Z(n3360) );
  NAND2_X1 U3122 ( .A1(n3634), .A2(n3360), .ZN(n2435) );
  NAND2_X1 U3123 ( .A1(n2014), .A2(REG1_REG_18__SCAN_IN), .ZN(n2443) );
  AND2_X1 U3124 ( .A1(REG3_REG_18__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .ZN(
        n4589) );
  AOI21_X1 U3125 ( .B1(n2436), .B2(REG3_REG_17__SCAN_IN), .A(
        REG3_REG_18__SCAN_IN), .ZN(n2437) );
  NOR2_X1 U3126 ( .A1(n2447), .A2(n2437), .ZN(n4117) );
  NAND2_X1 U3127 ( .A1(n2012), .A2(n4117), .ZN(n2442) );
  NAND2_X1 U3128 ( .A1(n3666), .A2(REG0_REG_18__SCAN_IN), .ZN(n2441) );
  INV_X1 U3129 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2439) );
  OR2_X1 U3130 ( .A1(n2260), .A2(n2439), .ZN(n2440) );
  NAND4_X1 U3131 ( .A1(n2443), .A2(n2442), .A3(n2441), .A4(n2440), .ZN(n4087)
         );
  INV_X1 U3132 ( .A(n4087), .ZN(n3594) );
  NAND2_X1 U3133 ( .A1(n2445), .A2(n2444), .ZN(n2454) );
  NAND2_X1 U3134 ( .A1(n2454), .A2(IR_REG_31__SCAN_IN), .ZN(n2446) );
  XNOR2_X1 U3135 ( .A(n2446), .B(IR_REG_18__SCAN_IN), .ZN(n3903) );
  MUX2_X1 U3136 ( .A(n3903), .B(DATAI_18_), .S(n2265), .Z(n4113) );
  NAND2_X1 U3137 ( .A1(n3594), .A2(n4113), .ZN(n4080) );
  INV_X1 U3138 ( .A(n4113), .ZN(n4100) );
  NAND2_X1 U3139 ( .A1(n4087), .A2(n4100), .ZN(n4081) );
  NAND2_X1 U3140 ( .A1(n4080), .A2(n4081), .ZN(n4111) );
  NAND2_X1 U3141 ( .A1(n2013), .A2(REG1_REG_19__SCAN_IN), .ZN(n2453) );
  OR2_X1 U3142 ( .A1(n2447), .A2(REG3_REG_19__SCAN_IN), .ZN(n2448) );
  AND2_X1 U3143 ( .A1(n2469), .A2(n2448), .ZN(n4093) );
  NAND2_X1 U3144 ( .A1(n2012), .A2(n4093), .ZN(n2452) );
  NAND2_X1 U3145 ( .A1(n3666), .A2(REG0_REG_19__SCAN_IN), .ZN(n2451) );
  INV_X1 U3146 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2449) );
  OR2_X1 U3147 ( .A1(n3670), .A2(n2449), .ZN(n2450) );
  INV_X1 U31480 ( .A(n2454), .ZN(n2456) );
  NAND2_X1 U31490 ( .A1(n2456), .A2(n2455), .ZN(n2457) );
  NAND2_X2 U3150 ( .A1(n2457), .A2(IR_REG_31__SCAN_IN), .ZN(n2536) );
  NAND2_X1 U3151 ( .A1(n2536), .A2(n4518), .ZN(n2532) );
  OR2_X1 U3152 ( .A1(n2536), .A2(n4518), .ZN(n2458) );
  MUX2_X1 U3153 ( .A(n4247), .B(DATAI_19_), .S(n2265), .Z(n3400) );
  NAND2_X1 U3154 ( .A1(n4063), .A2(n3400), .ZN(n4053) );
  NAND2_X1 U3155 ( .A1(n2014), .A2(REG1_REG_20__SCAN_IN), .ZN(n2463) );
  XNOR2_X1 U3156 ( .A(n2469), .B(REG3_REG_20__SCAN_IN), .ZN(n4070) );
  NAND2_X1 U3157 ( .A1(n2012), .A2(n4070), .ZN(n2462) );
  NAND2_X1 U3158 ( .A1(n3666), .A2(REG0_REG_20__SCAN_IN), .ZN(n2461) );
  INV_X1 U3159 ( .A(REG2_REG_20__SCAN_IN), .ZN(n2459) );
  OR2_X1 U3160 ( .A1(n2260), .A2(n2459), .ZN(n2460) );
  INV_X1 U3161 ( .A(n4042), .ZN(n4085) );
  NAND2_X1 U3162 ( .A1(n4085), .A2(n4067), .ZN(n2465) );
  INV_X1 U3163 ( .A(n4067), .ZN(n3731) );
  AOI21_X1 U3164 ( .B1(n2466), .B2(n2465), .A(n2464), .ZN(n4036) );
  NAND2_X1 U3165 ( .A1(n2014), .A2(REG1_REG_21__SCAN_IN), .ZN(n2475) );
  INV_X1 U3166 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3617) );
  INV_X1 U3167 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2467) );
  OAI21_X1 U3168 ( .B1(n2469), .B2(n3617), .A(n2467), .ZN(n2470) );
  NAND2_X1 U3169 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2468) );
  AND2_X1 U3170 ( .A1(n2470), .A2(n2478), .ZN(n4048) );
  NAND2_X1 U3171 ( .A1(n2012), .A2(n4048), .ZN(n2474) );
  NAND2_X1 U3172 ( .A1(n3666), .A2(REG0_REG_21__SCAN_IN), .ZN(n2473) );
  INV_X1 U3173 ( .A(REG2_REG_21__SCAN_IN), .ZN(n2471) );
  OR2_X1 U3174 ( .A1(n3670), .A2(n2471), .ZN(n2472) );
  NAND4_X1 U3175 ( .A1(n2475), .A2(n2474), .A3(n2473), .A4(n2472), .ZN(n4027)
         );
  NAND2_X1 U3176 ( .A1(n2265), .A2(DATAI_21_), .ZN(n4039) );
  NAND2_X1 U3177 ( .A1(n4027), .A2(n4045), .ZN(n2477) );
  INV_X1 U3178 ( .A(n4027), .ZN(n4055) );
  AOI21_X1 U3179 ( .B1(n4036), .B2(n2477), .A(n2476), .ZN(n4016) );
  INV_X1 U3180 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4485) );
  NAND2_X1 U3181 ( .A1(n2478), .A2(n4485), .ZN(n2479) );
  NAND2_X1 U3182 ( .A1(n2485), .A2(n2479), .ZN(n4018) );
  INV_X1 U3183 ( .A(n4018), .ZN(n3627) );
  NAND2_X1 U3184 ( .A1(n3627), .A2(n2012), .ZN(n2483) );
  NAND2_X1 U3185 ( .A1(n2013), .A2(REG1_REG_22__SCAN_IN), .ZN(n2482) );
  INV_X1 U3186 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4019) );
  OR2_X1 U3187 ( .A1(n3670), .A2(n4019), .ZN(n2481) );
  NAND2_X1 U3188 ( .A1(n3666), .A2(REG0_REG_22__SCAN_IN), .ZN(n2480) );
  NAND4_X1 U3189 ( .A1(n2483), .A2(n2482), .A3(n2481), .A4(n2480), .ZN(n4002)
         );
  NAND2_X1 U3190 ( .A1(n4040), .A2(n4017), .ZN(n3998) );
  NAND2_X1 U3191 ( .A1(n4002), .A2(n4030), .ZN(n2576) );
  NAND2_X1 U3192 ( .A1(n3998), .A2(n2576), .ZN(n4015) );
  NAND2_X1 U3193 ( .A1(n4016), .A2(n4015), .ZN(n4014) );
  NAND2_X1 U3194 ( .A1(n4014), .A2(n2484), .ZN(n3993) );
  INV_X1 U3195 ( .A(REG2_REG_23__SCAN_IN), .ZN(n2489) );
  INV_X1 U3196 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3526) );
  AND2_X1 U3197 ( .A1(n2485), .A2(n3526), .ZN(n2486) );
  NOR2_X1 U3198 ( .A1(n2492), .A2(n2486), .ZN(n4009) );
  NAND2_X1 U3199 ( .A1(n4009), .A2(n2012), .ZN(n2488) );
  AOI22_X1 U3200 ( .A1(n2014), .A2(REG1_REG_23__SCAN_IN), .B1(n2011), .B2(
        REG0_REG_23__SCAN_IN), .ZN(n2487) );
  OAI211_X1 U3201 ( .C1(n3670), .C2(n2489), .A(n2488), .B(n2487), .ZN(n4026)
         );
  INV_X1 U3202 ( .A(n4026), .ZN(n3624) );
  NAND2_X1 U3203 ( .A1(n2265), .A2(DATAI_23_), .ZN(n3527) );
  NAND2_X1 U3204 ( .A1(n3624), .A2(n3527), .ZN(n2491) );
  OR2_X1 U3205 ( .A1(n2492), .A2(REG3_REG_24__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U3206 ( .A1(n2498), .A2(n2493), .ZN(n3987) );
  INV_X1 U3207 ( .A(n2012), .ZN(n2513) );
  INV_X1 U3208 ( .A(n2260), .ZN(n2500) );
  AOI22_X1 U3209 ( .A1(n2500), .A2(REG2_REG_24__SCAN_IN), .B1(n2013), .B2(
        REG1_REG_24__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U32100 ( .A1(n3666), .A2(REG0_REG_24__SCAN_IN), .ZN(n2494) );
  NAND2_X1 U32110 ( .A1(n2265), .A2(DATAI_24_), .ZN(n3986) );
  NAND2_X1 U32120 ( .A1(n4001), .A2(n3981), .ZN(n2497) );
  NOR2_X1 U32130 ( .A1(n4001), .A2(n3981), .ZN(n2496) );
  AOI21_X1 U32140 ( .B1(n3974), .B2(n2497), .A(n2496), .ZN(n3957) );
  INV_X1 U32150 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3571) );
  NAND2_X1 U32160 ( .A1(n2498), .A2(n3571), .ZN(n2499) );
  NAND2_X1 U32170 ( .A1(n2506), .A2(n2499), .ZN(n3570) );
  AOI22_X1 U32180 ( .A1(n2500), .A2(REG2_REG_25__SCAN_IN), .B1(n2014), .B2(
        REG1_REG_25__SCAN_IN), .ZN(n2502) );
  NAND2_X1 U32190 ( .A1(n3666), .A2(REG0_REG_25__SCAN_IN), .ZN(n2501) );
  NAND2_X1 U32200 ( .A1(n2265), .A2(DATAI_25_), .ZN(n3572) );
  NAND2_X1 U32210 ( .A1(n3957), .A2(n2213), .ZN(n2505) );
  INV_X1 U32220 ( .A(n3944), .ZN(n3984) );
  INV_X1 U32230 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4479) );
  AND2_X1 U32240 ( .A1(n2506), .A2(n4479), .ZN(n2507) );
  INV_X1 U32250 ( .A(REG2_REG_26__SCAN_IN), .ZN(n2510) );
  NAND2_X1 U32260 ( .A1(n3666), .A2(REG0_REG_26__SCAN_IN), .ZN(n2509) );
  NAND2_X1 U32270 ( .A1(n2014), .A2(REG1_REG_26__SCAN_IN), .ZN(n2508) );
  OAI211_X1 U32280 ( .C1(n3670), .C2(n2510), .A(n2509), .B(n2508), .ZN(n2511)
         );
  INV_X1 U32290 ( .A(n2511), .ZN(n2512) );
  NAND2_X1 U32300 ( .A1(n2265), .A2(DATAI_26_), .ZN(n3950) );
  NOR2_X1 U32310 ( .A1(n3966), .A2(n3950), .ZN(n2515) );
  NAND2_X1 U32320 ( .A1(n3966), .A2(n3950), .ZN(n2514) );
  NAND2_X1 U32330 ( .A1(n2516), .A2(REG3_REG_27__SCAN_IN), .ZN(n2524) );
  OR2_X1 U32340 ( .A1(n2516), .A2(REG3_REG_27__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U32350 ( .A1(n3519), .A2(n2012), .ZN(n2522) );
  INV_X1 U32360 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3473) );
  NAND2_X1 U32370 ( .A1(n2013), .A2(REG1_REG_27__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U32380 ( .A1(n3666), .A2(REG0_REG_27__SCAN_IN), .ZN(n2518) );
  OAI211_X1 U32390 ( .C1(n3473), .C2(n3670), .A(n2519), .B(n2518), .ZN(n2520)
         );
  INV_X1 U32400 ( .A(n2520), .ZN(n2521) );
  AND2_X1 U32410 ( .A1(n2265), .A2(DATAI_27_), .ZN(n3480) );
  NOR2_X1 U32420 ( .A1(n3945), .A2(n3480), .ZN(n2523) );
  INV_X1 U32430 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3464) );
  NAND2_X1 U32440 ( .A1(n2524), .A2(n3464), .ZN(n2525) );
  NAND2_X1 U32450 ( .A1(n3506), .A2(n2012), .ZN(n2531) );
  INV_X1 U32460 ( .A(REG2_REG_28__SCAN_IN), .ZN(n2528) );
  NAND2_X1 U32470 ( .A1(n2014), .A2(REG1_REG_28__SCAN_IN), .ZN(n2527) );
  NAND2_X1 U32480 ( .A1(n3666), .A2(REG0_REG_28__SCAN_IN), .ZN(n2526) );
  OAI211_X1 U32490 ( .C1(n2528), .C2(n3670), .A(n2527), .B(n2526), .ZN(n2529)
         );
  INV_X1 U32500 ( .A(n2529), .ZN(n2530) );
  NAND2_X1 U32510 ( .A1(n2265), .A2(DATAI_28_), .ZN(n3465) );
  NAND2_X1 U32520 ( .A1(n3927), .A2(n3465), .ZN(n3915) );
  NAND2_X1 U32530 ( .A1(n3913), .A2(n3915), .ZN(n3924) );
  XNOR2_X1 U32540 ( .A(n3925), .B(n3924), .ZN(n3512) );
  OAI21_X1 U32550 ( .B1(IR_REG_20__SCAN_IN), .B2(IR_REG_19__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2535) );
  NAND2_X1 U32560 ( .A1(n2536), .A2(n2535), .ZN(n2538) );
  NAND2_X1 U32570 ( .A1(n2539), .A2(IR_REG_31__SCAN_IN), .ZN(n2540) );
  XNOR2_X1 U32580 ( .A(n2540), .B(n2207), .ZN(n2552) );
  XNOR2_X1 U32590 ( .A(n2767), .B(n4245), .ZN(n2541) );
  NAND2_X1 U32600 ( .A1(n2541), .A2(n3908), .ZN(n4065) );
  AND2_X1 U32610 ( .A1(n2542), .A2(n4247), .ZN(n4363) );
  INV_X1 U32620 ( .A(n4402), .ZN(n4394) );
  NAND2_X1 U32630 ( .A1(n4065), .A2(n4394), .ZN(n4410) );
  INV_X1 U32640 ( .A(n2543), .ZN(n2545) );
  MUX2_X1 U32650 ( .A(n2543), .B(n2545), .S(n2544), .Z(n4254) );
  INV_X1 U32660 ( .A(REG2_REG_29__SCAN_IN), .ZN(n2549) );
  NAND2_X1 U32670 ( .A1(n3666), .A2(REG0_REG_29__SCAN_IN), .ZN(n2548) );
  NAND2_X1 U32680 ( .A1(n2014), .A2(REG1_REG_29__SCAN_IN), .ZN(n2547) );
  OAI211_X1 U32690 ( .C1(n3670), .C2(n2549), .A(n2548), .B(n2547), .ZN(n2550)
         );
  INV_X1 U32700 ( .A(n2642), .ZN(n2763) );
  NOR2_X2 U32710 ( .A1(n4254), .A2(n2763), .ZN(n4025) );
  INV_X1 U32720 ( .A(n2542), .ZN(n4246) );
  OAI22_X1 U32730 ( .A1(n3699), .A2(n4101), .B1(n3465), .B2(n4134), .ZN(n2582)
         );
  INV_X1 U32740 ( .A(n3543), .ZN(n2554) );
  NAND2_X1 U32750 ( .A1(n2554), .A2(n2774), .ZN(n3741) );
  NAND2_X1 U32760 ( .A1(n2844), .A2(n3745), .ZN(n3017) );
  NAND2_X1 U32770 ( .A1(n2556), .A2(n3018), .ZN(n3750) );
  NAND2_X1 U32780 ( .A1(n3831), .A2(n3024), .ZN(n3747) );
  AND2_X1 U32790 ( .A1(n3750), .A2(n3747), .ZN(n3714) );
  NAND2_X1 U32800 ( .A1(n3017), .A2(n3714), .ZN(n3016) );
  INV_X1 U32810 ( .A(n3751), .ZN(n2557) );
  AND2_X1 U32820 ( .A1(n3829), .A2(n2558), .ZN(n2933) );
  NAND2_X1 U32830 ( .A1(n2965), .A2(n2941), .ZN(n3762) );
  NAND2_X1 U32840 ( .A1(n3828), .A2(n2980), .ZN(n3761) );
  NAND2_X1 U32850 ( .A1(n2972), .A2(n3761), .ZN(n2559) );
  INV_X1 U32860 ( .A(n3828), .ZN(n3000) );
  NAND2_X1 U32870 ( .A1(n3000), .A2(n2973), .ZN(n3756) );
  INV_X1 U32880 ( .A(n2560), .ZN(n2561) );
  NAND2_X1 U32890 ( .A1(n3115), .A2(n3081), .ZN(n3765) );
  NAND2_X1 U32900 ( .A1(n3827), .A2(n2562), .ZN(n3759) );
  AND2_X1 U32910 ( .A1(n3826), .A2(n3048), .ZN(n3772) );
  NAND2_X1 U32920 ( .A1(n3138), .A2(n3118), .ZN(n3766) );
  INV_X1 U32930 ( .A(n3140), .ZN(n3091) );
  NAND2_X1 U32940 ( .A1(n3825), .A2(n3091), .ZN(n3774) );
  NAND2_X1 U32950 ( .A1(n3085), .A2(n3774), .ZN(n2564) );
  INV_X1 U32960 ( .A(n3825), .ZN(n3114) );
  NAND2_X1 U32970 ( .A1(n3114), .A2(n3140), .ZN(n3771) );
  NAND2_X1 U32980 ( .A1(n3823), .A2(n3149), .ZN(n3264) );
  NAND2_X1 U32990 ( .A1(n3822), .A2(n3276), .ZN(n2565) );
  NOR2_X1 U33000 ( .A1(n3823), .A2(n3149), .ZN(n3265) );
  NOR2_X1 U33010 ( .A1(n3822), .A2(n3276), .ZN(n2566) );
  AOI21_X1 U33020 ( .B1(n3776), .B2(n3265), .A(n2566), .ZN(n3779) );
  INV_X1 U33030 ( .A(n3711), .ZN(n2567) );
  NAND2_X1 U33040 ( .A1(n3682), .A2(n2567), .ZN(n2568) );
  NAND2_X1 U33050 ( .A1(n3581), .A2(n3373), .ZN(n3681) );
  NAND2_X1 U33060 ( .A1(n3821), .A2(n3657), .ZN(n3679) );
  NAND2_X1 U33070 ( .A1(n3681), .A2(n3679), .ZN(n3716) );
  NAND2_X1 U33080 ( .A1(n3347), .A2(n3679), .ZN(n3300) );
  INV_X1 U33090 ( .A(n3719), .ZN(n3299) );
  NAND2_X1 U33100 ( .A1(n4063), .A2(n4090), .ZN(n2569) );
  AND2_X1 U33110 ( .A1(n4081), .A2(n2569), .ZN(n2571) );
  NAND2_X1 U33120 ( .A1(n4108), .A2(n3360), .ZN(n4076) );
  NAND2_X1 U33130 ( .A1(n2571), .A2(n4076), .ZN(n3787) );
  NAND2_X1 U33140 ( .A1(n3634), .A2(n3596), .ZN(n4077) );
  NAND2_X1 U33150 ( .A1(n4080), .A2(n4077), .ZN(n2572) );
  NOR2_X1 U33160 ( .A1(n4063), .A2(n4090), .ZN(n2570) );
  AOI21_X1 U33170 ( .B1(n2572), .B2(n2571), .A(n2570), .ZN(n4056) );
  NAND2_X1 U33180 ( .A1(n4085), .A2(n3731), .ZN(n2573) );
  AND2_X1 U33190 ( .A1(n4056), .A2(n2573), .ZN(n3685) );
  NAND2_X1 U33200 ( .A1(n4042), .A2(n4067), .ZN(n3790) );
  INV_X1 U33210 ( .A(n3998), .ZN(n2575) );
  NOR2_X1 U33220 ( .A1(n4027), .A2(n4039), .ZN(n3995) );
  NOR2_X1 U33230 ( .A1(n2575), .A2(n3995), .ZN(n3795) );
  NAND2_X1 U33240 ( .A1(n4026), .A2(n3527), .ZN(n3705) );
  AND2_X1 U33250 ( .A1(n3705), .A2(n2576), .ZN(n3800) );
  AND2_X1 U33260 ( .A1(n4027), .A2(n4039), .ZN(n3994) );
  NAND2_X1 U33270 ( .A1(n3998), .A2(n3994), .ZN(n2577) );
  NAND2_X1 U33280 ( .A1(n3800), .A2(n2577), .ZN(n3687) );
  OR2_X1 U33290 ( .A1(n4001), .A2(n3986), .ZN(n3702) );
  OR2_X1 U33300 ( .A1(n4026), .A2(n3527), .ZN(n3975) );
  NAND2_X1 U33310 ( .A1(n3702), .A2(n3975), .ZN(n3798) );
  OR2_X1 U33320 ( .A1(n3481), .A2(n3950), .ZN(n3729) );
  OR2_X1 U33330 ( .A1(n3944), .A2(n3572), .ZN(n3939) );
  NAND2_X1 U33340 ( .A1(n3944), .A2(n3572), .ZN(n3701) );
  NAND2_X1 U33350 ( .A1(n4001), .A2(n3986), .ZN(n3959) );
  AND2_X1 U33360 ( .A1(n3701), .A2(n3959), .ZN(n3689) );
  INV_X1 U33370 ( .A(n3689), .ZN(n3940) );
  NAND2_X1 U33380 ( .A1(n3796), .A2(n3940), .ZN(n2578) );
  AND2_X1 U33390 ( .A1(n3481), .A2(n3950), .ZN(n3673) );
  INV_X1 U33400 ( .A(n3673), .ZN(n3730) );
  NAND2_X1 U33410 ( .A1(n2578), .A2(n3730), .ZN(n3802) );
  NOR2_X1 U33420 ( .A1(n3644), .A2(n3480), .ZN(n3804) );
  INV_X1 U33430 ( .A(n3804), .ZN(n2579) );
  NAND2_X1 U33440 ( .A1(n3644), .A2(n3480), .ZN(n3674) );
  NAND2_X1 U33450 ( .A1(n2579), .A2(n3674), .ZN(n3728) );
  NAND2_X1 U33460 ( .A1(n3477), .A2(n3478), .ZN(n3476) );
  NAND2_X1 U33470 ( .A1(n4246), .A2(n2551), .ZN(n2581) );
  NAND2_X1 U33480 ( .A1(n4247), .A2(n4245), .ZN(n2580) );
  OAI21_X1 U33490 ( .B1(n3512), .B2(n4416), .A(n3505), .ZN(n2617) );
  NAND2_X1 U33500 ( .A1(n4402), .A2(n2583), .ZN(n2610) );
  NAND2_X1 U33510 ( .A1(n2542), .A2(n3908), .ZN(n2584) );
  NAND2_X1 U33520 ( .A1(n2584), .A2(n2642), .ZN(n2780) );
  OR2_X1 U3353 ( .A1(n2586), .A2(n2585), .ZN(n2595) );
  NAND2_X1 U33540 ( .A1(n2595), .A2(n2594), .ZN(n2587) );
  NAND2_X1 U3355 ( .A1(n2587), .A2(IR_REG_31__SCAN_IN), .ZN(n2588) );
  NAND2_X1 U3356 ( .A1(n2589), .A2(IR_REG_31__SCAN_IN), .ZN(n2590) );
  OAI21_X1 U3357 ( .B1(IR_REG_23__SCAN_IN), .B2(IR_REG_24__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2591) );
  NAND2_X1 U3358 ( .A1(n2595), .A2(n2591), .ZN(n2593) );
  XNOR2_X1 U3359 ( .A(n2593), .B(n2592), .ZN(n2627) );
  XNOR2_X1 U3360 ( .A(n2595), .B(n2594), .ZN(n2644) );
  INV_X1 U3361 ( .A(n2627), .ZN(n2598) );
  NAND2_X1 U3362 ( .A1(n2598), .A2(B_REG_SCAN_IN), .ZN(n2596) );
  MUX2_X1 U3363 ( .A(n2596), .B(B_REG_SCAN_IN), .S(n4244), .Z(n2597) );
  NAND2_X1 U3364 ( .A1(n2597), .A2(n4243), .ZN(n2635) );
  INV_X1 U3365 ( .A(n4243), .ZN(n2638) );
  NAND2_X1 U3366 ( .A1(n2598), .A2(n2638), .ZN(n2636) );
  OAI21_X1 U3367 ( .B1(n2635), .B2(D_REG_1__SCAN_IN), .A(n2636), .ZN(n2609) );
  NOR4_X1 U3368 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n4559) );
  NOR2_X1 U3369 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .ZN(n2601)
         );
  NOR4_X1 U3370 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2600) );
  NOR4_X1 U3371 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_31__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2599) );
  AND4_X1 U3372 ( .A1(n4559), .A2(n2601), .A3(n2600), .A4(n2599), .ZN(n2607)
         );
  NOR4_X1 U3373 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2605) );
  NOR4_X1 U3374 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2604) );
  NOR4_X1 U3375 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2603) );
  NOR4_X1 U3376 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2602) );
  AND4_X1 U3377 ( .A1(n2605), .A2(n2604), .A3(n2603), .A4(n2602), .ZN(n2606)
         );
  NAND2_X1 U3378 ( .A1(n2607), .A2(n2606), .ZN(n2756) );
  NAND2_X1 U3379 ( .A1(n2760), .A2(n2756), .ZN(n2608) );
  NAND4_X1 U3380 ( .A1(n2610), .A2(n2881), .A3(n2609), .A4(n2608), .ZN(n2616)
         );
  INV_X1 U3381 ( .A(D_REG_0__SCAN_IN), .ZN(n2641) );
  NAND2_X1 U3382 ( .A1(n2760), .A2(n2641), .ZN(n2612) );
  INV_X1 U3383 ( .A(n4244), .ZN(n2639) );
  NAND2_X1 U3384 ( .A1(n2639), .A2(n2638), .ZN(n2611) );
  NAND2_X1 U3385 ( .A1(n2612), .A2(n2611), .ZN(n2880) );
  INV_X1 U3386 ( .A(n2613), .ZN(n2615) );
  NOR2_X2 U3387 ( .A1(n3497), .A2(n2941), .ZN(n2981) );
  AND2_X2 U3388 ( .A1(n2981), .A2(n2980), .ZN(n2983) );
  NAND2_X2 U3389 ( .A1(n2983), .A2(n2884), .ZN(n3038) );
  INV_X1 U3390 ( .A(n3950), .ZN(n3943) );
  OAI21_X1 U3391 ( .B1(n3472), .B2(n3465), .A(n3933), .ZN(n3508) );
  NAND2_X1 U3392 ( .A1(n2615), .A2(n2217), .ZN(U3546) );
  INV_X1 U3393 ( .A(n2880), .ZN(n2761) );
  INV_X1 U3394 ( .A(n2618), .ZN(n2619) );
  NAND2_X1 U3395 ( .A1(n2619), .A2(n2216), .ZN(U3514) );
  INV_X1 U3396 ( .A(n4374), .ZN(n2620) );
  OR2_X2 U3397 ( .A1(n2771), .A2(n2620), .ZN(n3833) );
  INV_X2 U3398 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3399 ( .A(DATAI_3_), .ZN(n2621) );
  MUX2_X1 U3400 ( .A(n2678), .B(n2621), .S(U3149), .Z(n2622) );
  INV_X1 U3401 ( .A(n2622), .ZN(U3349) );
  INV_X1 U3402 ( .A(DATAI_6_), .ZN(n2623) );
  MUX2_X1 U3403 ( .A(n2057), .B(n2623), .S(U3149), .Z(n2624) );
  INV_X1 U3404 ( .A(n2624), .ZN(U3346) );
  INV_X1 U3405 ( .A(n3873), .ZN(n3890) );
  INV_X1 U3406 ( .A(DATAI_9_), .ZN(n2625) );
  MUX2_X1 U3407 ( .A(n3890), .B(n2625), .S(U3149), .Z(n2626) );
  INV_X1 U3408 ( .A(n2626), .ZN(U3343) );
  INV_X1 U3409 ( .A(DATAI_25_), .ZN(n2629) );
  NAND2_X1 U3410 ( .A1(n2627), .A2(STATE_REG_SCAN_IN), .ZN(n2628) );
  OAI21_X1 U3411 ( .B1(STATE_REG_SCAN_IN), .B2(n2629), .A(n2628), .ZN(U3327)
         );
  INV_X1 U3412 ( .A(DATAI_31_), .ZN(n2632) );
  OR4_X1 U3413 ( .A1(n2630), .A2(IR_REG_30__SCAN_IN), .A3(n2585), .A4(U3149), 
        .ZN(n2631) );
  OAI21_X1 U3414 ( .B1(STATE_REG_SCAN_IN), .B2(n2632), .A(n2631), .ZN(U3321)
         );
  INV_X1 U3415 ( .A(DATAI_21_), .ZN(n2634) );
  NAND2_X1 U3416 ( .A1(n2551), .A2(STATE_REG_SCAN_IN), .ZN(n2633) );
  OAI21_X1 U3417 ( .B1(STATE_REG_SCAN_IN), .B2(n2634), .A(n2633), .ZN(U3331)
         );
  NAND2_X1 U3418 ( .A1(n2635), .A2(n2787), .ZN(n4373) );
  INV_X1 U3419 ( .A(D_REG_1__SCAN_IN), .ZN(n2637) );
  INV_X1 U3420 ( .A(n2636), .ZN(n2758) );
  AOI22_X1 U3421 ( .A1(n4373), .A2(n2637), .B1(n2758), .B2(n4374), .ZN(U3459)
         );
  AND2_X1 U3422 ( .A1(n2638), .A2(n4374), .ZN(n2640) );
  AOI22_X1 U3423 ( .A1(n4373), .A2(n2641), .B1(n2640), .B2(n2639), .ZN(U3458)
         );
  NAND2_X1 U3424 ( .A1(n2642), .A2(n2644), .ZN(n2643) );
  AND2_X1 U3425 ( .A1(n2643), .A2(n2265), .ZN(n2660) );
  INV_X1 U3426 ( .A(n2660), .ZN(n2647) );
  INV_X1 U3427 ( .A(n2644), .ZN(n2645) );
  NAND2_X1 U3428 ( .A1(n2645), .A2(STATE_REG_SCAN_IN), .ZN(n3818) );
  INV_X1 U3429 ( .A(n3818), .ZN(n2646) );
  OR2_X1 U3430 ( .A1(n2787), .A2(n2646), .ZN(n2659) );
  NOR2_X1 U3431 ( .A1(n4442), .A2(U4043), .ZN(U3148) );
  INV_X1 U3432 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n4469) );
  NAND2_X1 U3433 ( .A1(n2997), .A2(U4043), .ZN(n2648) );
  OAI21_X1 U3434 ( .B1(U4043), .B2(n4469), .A(n2648), .ZN(U3557) );
  INV_X1 U3435 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n4468) );
  NAND2_X1 U3436 ( .A1(n3352), .A2(U4043), .ZN(n2649) );
  OAI21_X1 U3437 ( .B1(U4043), .B2(n4468), .A(n2649), .ZN(U3564) );
  INV_X1 U3438 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4478) );
  INV_X1 U3439 ( .A(REG2_REG_31__SCAN_IN), .ZN(n2652) );
  NAND2_X1 U3440 ( .A1(n2014), .A2(REG1_REG_31__SCAN_IN), .ZN(n2651) );
  NAND2_X1 U3441 ( .A1(n3666), .A2(REG0_REG_31__SCAN_IN), .ZN(n2650) );
  OAI211_X1 U3442 ( .C1(n3670), .C2(n2652), .A(n2651), .B(n2650), .ZN(n4123)
         );
  NAND2_X1 U3443 ( .A1(n4123), .A2(U4043), .ZN(n2653) );
  OAI21_X1 U3444 ( .B1(U4043), .B2(n4478), .A(n2653), .ZN(U3581) );
  INV_X1 U3445 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4466) );
  NAND2_X1 U3446 ( .A1(n3543), .A2(U4043), .ZN(n2654) );
  OAI21_X1 U3447 ( .B1(U4043), .B2(n4466), .A(n2654), .ZN(U3550) );
  INV_X1 U3448 ( .A(n4442), .ZN(n4318) );
  INV_X1 U3449 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n2664) );
  XNOR2_X1 U3450 ( .A(n2655), .B(IR_REG_27__SCAN_IN), .ZN(n4242) );
  NAND2_X1 U3451 ( .A1(n4242), .A2(n2252), .ZN(n2656) );
  AND2_X1 U3452 ( .A1(n4254), .A2(n2656), .ZN(n3848) );
  OAI21_X1 U3453 ( .B1(n4242), .B2(REG1_REG_0__SCAN_IN), .A(n4504), .ZN(n2658)
         );
  INV_X1 U3454 ( .A(IR_REG_0__SCAN_IN), .ZN(n4504) );
  NOR2_X1 U3455 ( .A1(n3848), .A2(IR_REG_0__SCAN_IN), .ZN(n2657) );
  AOI21_X1 U3456 ( .B1(n3848), .B2(n2658), .A(n2657), .ZN(n2661) );
  AND2_X1 U3457 ( .A1(n2660), .A2(n2659), .ZN(n2672) );
  AOI22_X1 U34580 ( .A1(n2661), .A2(n2672), .B1(REG3_REG_0__SCAN_IN), .B2(
        U3149), .ZN(n2663) );
  INV_X1 U34590 ( .A(n4242), .ZN(n3844) );
  INV_X1 U3460 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2770) );
  NAND3_X1 U3461 ( .A1(n4337), .A2(n2770), .A3(IR_REG_0__SCAN_IN), .ZN(n2662)
         );
  OAI211_X1 U3462 ( .C1(n4318), .C2(n2664), .A(n2663), .B(n2662), .ZN(U3240)
         );
  NOR2_X1 U3463 ( .A1(STATE_REG_SCAN_IN), .A2(n2272), .ZN(n2871) );
  INV_X1 U3464 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n4464) );
  NAND2_X1 U3465 ( .A1(n4254), .A2(n4242), .ZN(n3814) );
  INV_X1 U3466 ( .A(n3814), .ZN(n2665) );
  MUX2_X1 U34670 ( .A(REG2_REG_2__SCAN_IN), .B(n2928), .S(n4252), .Z(n2667) );
  MUX2_X1 U3468 ( .A(REG2_REG_1__SCAN_IN), .B(n2247), .S(n4253), .Z(n3835) );
  AND2_X1 U34690 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3843) );
  NAND2_X1 U3470 ( .A1(n2008), .A2(REG2_REG_1__SCAN_IN), .ZN(n3852) );
  NAND2_X1 U34710 ( .A1(n3853), .A2(n3852), .ZN(n2666) );
  NAND2_X1 U3472 ( .A1(n2667), .A2(n2666), .ZN(n3856) );
  NAND2_X1 U34730 ( .A1(n4252), .A2(REG2_REG_2__SCAN_IN), .ZN(n2668) );
  NAND2_X1 U3474 ( .A1(n3856), .A2(n2668), .ZN(n2692) );
  XOR2_X1 U34750 ( .A(REG2_REG_3__SCAN_IN), .B(n2690), .Z(n2669) );
  NAND2_X1 U3476 ( .A1(n4348), .A2(n2669), .ZN(n2670) );
  OAI21_X1 U34770 ( .B1(n4464), .B2(n4318), .A(n2670), .ZN(n2671) );
  NOR2_X1 U3478 ( .A1(n2871), .A2(n2671), .ZN(n2681) );
  INV_X1 U34790 ( .A(n4254), .ZN(n2791) );
  XNOR2_X1 U3480 ( .A(n4252), .B(REG1_REG_2__SCAN_IN), .ZN(n3850) );
  INV_X1 U34810 ( .A(n3850), .ZN(n2675) );
  INV_X1 U3482 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2673) );
  XNOR2_X1 U34830 ( .A(n2008), .B(n2673), .ZN(n3838) );
  AND2_X1 U3484 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3837)
         );
  NAND2_X1 U34850 ( .A1(n3838), .A2(n3837), .ZN(n3836) );
  NAND2_X1 U3486 ( .A1(n2008), .A2(REG1_REG_1__SCAN_IN), .ZN(n2674) );
  NAND2_X1 U34870 ( .A1(n3836), .A2(n2674), .ZN(n3849) );
  NAND2_X1 U3488 ( .A1(n2675), .A2(n3849), .ZN(n2677) );
  NAND2_X1 U34890 ( .A1(n4252), .A2(REG1_REG_2__SCAN_IN), .ZN(n2676) );
  NAND2_X1 U3490 ( .A1(n2677), .A2(n2676), .ZN(n2683) );
  XOR2_X1 U34910 ( .A(REG1_REG_3__SCAN_IN), .B(n2682), .Z(n2679) );
  AOI22_X1 U3492 ( .A1(n2691), .A2(n4315), .B1(n4337), .B2(n2679), .ZN(n2680)
         );
  NAND2_X1 U34930 ( .A1(n2681), .A2(n2680), .ZN(U3243) );
  NAND2_X1 U3494 ( .A1(n2683), .A2(n2691), .ZN(n2684) );
  INV_X1 U34950 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2685) );
  NAND2_X1 U3496 ( .A1(n2686), .A2(n4251), .ZN(n2687) );
  INV_X1 U34970 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2688) );
  MUX2_X1 U3498 ( .A(n2688), .B(REG1_REG_5__SCAN_IN), .S(n2706), .Z(n2711) );
  NAND2_X1 U34990 ( .A1(n2710), .A2(n2711), .ZN(n2709) );
  OR2_X1 U3500 ( .A1(n2706), .A2(n2688), .ZN(n2689) );
  NAND2_X1 U35010 ( .A1(n2709), .A2(n2689), .ZN(n2715) );
  XNOR2_X1 U3502 ( .A(n2714), .B(REG1_REG_6__SCAN_IN), .ZN(n2700) );
  INV_X1 U35030 ( .A(n2706), .ZN(n4250) );
  NAND2_X1 U3504 ( .A1(n2692), .A2(n2691), .ZN(n2693) );
  AOI22_X1 U35050 ( .A1(n2695), .A2(REG2_REG_4__SCAN_IN), .B1(n4251), .B2(
        n2694), .ZN(n2703) );
  MUX2_X1 U35060 ( .A(REG2_REG_5__SCAN_IN), .B(n2940), .S(n2706), .Z(n2702) );
  XOR2_X1 U35070 ( .A(REG2_REG_6__SCAN_IN), .B(n2721), .Z(n2698) );
  INV_X1 U35080 ( .A(REG3_REG_6__SCAN_IN), .ZN(n4481) );
  NOR2_X1 U35090 ( .A1(STATE_REG_SCAN_IN), .A2(n4481), .ZN(n2967) );
  AOI21_X1 U35100 ( .B1(n4442), .B2(ADDR_REG_6__SCAN_IN), .A(n2967), .ZN(n2696) );
  OAI21_X1 U35110 ( .B1(n4445), .B2(n2057), .A(n2696), .ZN(n2697) );
  AOI21_X1 U35120 ( .B1(n4348), .B2(n2698), .A(n2697), .ZN(n2699) );
  OAI21_X1 U35130 ( .B1(n2700), .B2(n4433), .A(n2699), .ZN(U3246) );
  INV_X1 U35140 ( .A(n4348), .ZN(n4437) );
  AOI211_X1 U35150 ( .C1(n2703), .C2(n2702), .A(n2701), .B(n4437), .ZN(n2708)
         );
  NOR2_X1 U35160 ( .A1(n2704), .A2(STATE_REG_SCAN_IN), .ZN(n2920) );
  AOI21_X1 U35170 ( .B1(n4442), .B2(ADDR_REG_5__SCAN_IN), .A(n2920), .ZN(n2705) );
  OAI21_X1 U35180 ( .B1(n4445), .B2(n2706), .A(n2705), .ZN(n2707) );
  NOR2_X1 U35190 ( .A1(n2708), .A2(n2707), .ZN(n2713) );
  OAI211_X1 U35200 ( .C1(n2711), .C2(n2710), .A(n4337), .B(n2709), .ZN(n2712)
         );
  NAND2_X1 U35210 ( .A1(n2713), .A2(n2712), .ZN(U3245) );
  NAND2_X1 U35220 ( .A1(n2715), .A2(n2720), .ZN(n2716) );
  INV_X1 U35230 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4428) );
  XNOR2_X1 U35240 ( .A(n4249), .B(n4428), .ZN(n2717) );
  XNOR2_X1 U35250 ( .A(n2748), .B(n2717), .ZN(n2727) );
  INV_X1 U35260 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n2719) );
  NOR2_X1 U35270 ( .A1(STATE_REG_SCAN_IN), .A2(n4576), .ZN(n3002) );
  INV_X1 U35280 ( .A(n3002), .ZN(n2718) );
  OAI21_X1 U35290 ( .B1(n4318), .B2(n2719), .A(n2718), .ZN(n2725) );
  INV_X1 U35300 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2886) );
  MUX2_X1 U35310 ( .A(n2886), .B(REG2_REG_7__SCAN_IN), .S(n4249), .Z(n2722) );
  NOR2_X1 U35320 ( .A1(n2723), .A2(n2722), .ZN(n2746) );
  AOI211_X1 U35330 ( .C1(n2723), .C2(n2722), .A(n4437), .B(n2746), .ZN(n2724)
         );
  AOI211_X1 U35340 ( .C1(n4315), .C2(n4249), .A(n2725), .B(n2724), .ZN(n2726)
         );
  OAI21_X1 U35350 ( .B1(n4433), .B2(n2727), .A(n2726), .ZN(U3247) );
  INV_X1 U35360 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4476) );
  NAND2_X1 U35370 ( .A1(n4002), .A2(U4043), .ZN(n2728) );
  OAI21_X1 U35380 ( .B1(U4043), .B2(n4476), .A(n2728), .ZN(U3572) );
  NAND2_X1 U35390 ( .A1(n3543), .A2(n2792), .ZN(n3742) );
  AND2_X1 U35400 ( .A1(n3741), .A2(n3742), .ZN(n3733) );
  INV_X1 U35410 ( .A(n3733), .ZN(n4369) );
  INV_X1 U35420 ( .A(n2614), .ZN(n2729) );
  NOR2_X1 U35430 ( .A1(n2792), .A2(n2729), .ZN(n4366) );
  INV_X1 U35440 ( .A(n4065), .ZN(n2978) );
  NOR2_X1 U35450 ( .A1(n2978), .A2(n4032), .ZN(n2731) );
  OAI22_X1 U35460 ( .A1(n3733), .A2(n2731), .B1(n2730), .B2(n4101), .ZN(n4364)
         );
  AOI211_X1 U35470 ( .C1(n4402), .C2(n4369), .A(n4366), .B(n4364), .ZN(n4389)
         );
  NAND2_X1 U35480 ( .A1(n4430), .A2(REG1_REG_0__SCAN_IN), .ZN(n2732) );
  OAI21_X1 U35490 ( .B1(n4389), .B2(n4430), .A(n2732), .ZN(U3518) );
  NAND2_X1 U35500 ( .A1(n2553), .A2(n3741), .ZN(n2733) );
  NAND2_X1 U35510 ( .A1(n2841), .A2(n2733), .ZN(n2737) );
  NAND2_X1 U35520 ( .A1(n3543), .A2(n4109), .ZN(n2735) );
  NAND2_X1 U35530 ( .A1(n3832), .A2(n4025), .ZN(n2734) );
  OAI211_X1 U35540 ( .C1(n4134), .C2(n2742), .A(n2735), .B(n2734), .ZN(n2736)
         );
  AOI21_X1 U35550 ( .B1(n2737), .B2(n4032), .A(n2736), .ZN(n2741) );
  INV_X1 U35560 ( .A(n2738), .ZN(n2739) );
  XNOR2_X1 U35570 ( .A(n2553), .B(n2739), .ZN(n3013) );
  NAND2_X1 U35580 ( .A1(n3013), .A2(n2978), .ZN(n2740) );
  NAND2_X1 U35590 ( .A1(n2741), .A2(n2740), .ZN(n3010) );
  INV_X1 U35600 ( .A(n3013), .ZN(n2743) );
  INV_X1 U35610 ( .A(n4421), .ZN(n4393) );
  OAI21_X1 U35620 ( .B1(n2792), .B2(n2742), .A(n2849), .ZN(n3009) );
  OAI22_X1 U35630 ( .A1(n2743), .A2(n4394), .B1(n4393), .B2(n3009), .ZN(n2744)
         );
  NOR2_X1 U35640 ( .A1(n3010), .A2(n2744), .ZN(n4391) );
  NAND2_X1 U35650 ( .A1(n4430), .A2(REG1_REG_1__SCAN_IN), .ZN(n2745) );
  OAI21_X1 U35660 ( .B1(n4391), .B2(n4430), .A(n2745), .ZN(U3519) );
  AOI21_X1 U35670 ( .B1(n4249), .B2(REG2_REG_7__SCAN_IN), .A(n2746), .ZN(n2795) );
  XNOR2_X1 U35680 ( .A(n2795), .B(n2802), .ZN(n2797) );
  XNOR2_X1 U35690 ( .A(n2797), .B(REG2_REG_8__SCAN_IN), .ZN(n2754) );
  INV_X1 U35700 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4453) );
  AND2_X1 U35710 ( .A1(n4249), .A2(REG1_REG_7__SCAN_IN), .ZN(n2747) );
  OR2_X1 U35720 ( .A1(n4249), .A2(REG1_REG_7__SCAN_IN), .ZN(n2749) );
  XNOR2_X1 U35730 ( .A(n2801), .B(n2802), .ZN(n2750) );
  AOI211_X1 U35740 ( .C1(n4453), .C2(n2750), .A(n4433), .B(n2803), .ZN(n2753)
         );
  AND2_X1 U35750 ( .A1(U3149), .A2(REG3_REG_8__SCAN_IN), .ZN(n3080) );
  AOI21_X1 U35760 ( .B1(n4442), .B2(ADDR_REG_8__SCAN_IN), .A(n3080), .ZN(n2751) );
  OAI21_X1 U35770 ( .B1(n4445), .B2(n2802), .A(n2751), .ZN(n2752) );
  AOI211_X1 U35780 ( .C1(n2754), .C2(n4348), .A(n2753), .B(n2752), .ZN(n2755)
         );
  INV_X1 U35790 ( .A(n2755), .ZN(U3248) );
  INV_X1 U35800 ( .A(n2756), .ZN(n2757) );
  NAND2_X1 U35810 ( .A1(n2757), .A2(D_REG_1__SCAN_IN), .ZN(n2759) );
  AOI21_X1 U3582 ( .B1(n2760), .B2(n2759), .A(n2758), .ZN(n2882) );
  NAND2_X1 U3583 ( .A1(n2882), .A2(n2761), .ZN(n2790) );
  NAND2_X1 U3584 ( .A1(n2614), .A2(n4247), .ZN(n2762) );
  NAND2_X1 U3585 ( .A1(n2763), .A2(n2762), .ZN(n2764) );
  NOR2_X1 U3586 ( .A1(n2764), .A2(n4127), .ZN(n2779) );
  NAND2_X1 U3587 ( .A1(n2779), .A2(n2787), .ZN(n2765) );
  AND2_X4 U3588 ( .A1(n2766), .A2(n2771), .ZN(n3458) );
  NAND2_X1 U3589 ( .A1(n3543), .A2(n3458), .ZN(n2769) );
  NAND2_X1 U3590 ( .A1(n2774), .A2(n2820), .ZN(n2768) );
  OR2_X1 U3591 ( .A1(n2771), .A2(n2770), .ZN(n2772) );
  INV_X1 U3592 ( .A(n3424), .ZN(n2824) );
  NAND2_X1 U3593 ( .A1(n3543), .A2(n2824), .ZN(n2776) );
  AND2_X1 U3594 ( .A1(n2854), .A2(IR_REG_0__SCAN_IN), .ZN(n2773) );
  NAND2_X1 U3595 ( .A1(n2776), .A2(n2775), .ZN(n2777) );
  NAND2_X1 U3596 ( .A1(n2778), .A2(n2777), .ZN(n2819) );
  OAI21_X1 U3597 ( .B1(n2778), .B2(n2777), .A(n2819), .ZN(n3846) );
  OAI21_X1 U3598 ( .B1(n4127), .B2(n2779), .A(n2790), .ZN(n2781) );
  NAND2_X1 U3599 ( .A1(n2781), .A2(n2780), .ZN(n2855) );
  INV_X1 U3600 ( .A(n2855), .ZN(n2785) );
  NAND2_X1 U3601 ( .A1(n3908), .A2(n4245), .ZN(n2813) );
  INV_X1 U3602 ( .A(n2813), .ZN(n2782) );
  AND2_X1 U3603 ( .A1(n2782), .A2(n4374), .ZN(n2783) );
  NAND2_X1 U3604 ( .A1(n3444), .A2(n2783), .ZN(n3815) );
  INV_X1 U3605 ( .A(n3815), .ZN(n2784) );
  NAND2_X1 U3606 ( .A1(n2790), .A2(n2784), .ZN(n2856) );
  NAND3_X1 U3607 ( .A1(n2785), .A2(n2787), .A3(n2856), .ZN(n3548) );
  INV_X1 U3608 ( .A(n2787), .ZN(n2786) );
  NOR3_X1 U3609 ( .A1(n2790), .A2(n4134), .A3(n2786), .ZN(n2789) );
  AND2_X1 U3610 ( .A1(n2787), .A2(n2583), .ZN(n2788) );
  NOR2_X2 U3611 ( .A1(n2789), .A2(n4367), .ZN(n3658) );
  NOR2_X1 U3612 ( .A1(n2790), .A2(n3815), .ZN(n2834) );
  NAND2_X1 U3613 ( .A1(n2834), .A2(n2791), .ZN(n3654) );
  OAI22_X1 U3614 ( .A1(n3658), .A2(n2792), .B1(n2730), .B2(n3654), .ZN(n2793)
         );
  AOI21_X1 U3615 ( .B1(REG3_REG_0__SCAN_IN), .B2(n3548), .A(n2793), .ZN(n2794)
         );
  OAI21_X1 U3616 ( .B1(n3664), .B2(n3846), .A(n2794), .ZN(U3229) );
  OAI22_X1 U3617 ( .A1(n2797), .A2(n2796), .B1(n2795), .B2(n2802), .ZN(n2799)
         );
  MUX2_X1 U3618 ( .A(REG2_REG_9__SCAN_IN), .B(n3055), .S(n3873), .Z(n2798) );
  NAND2_X1 U3619 ( .A1(n2799), .A2(n2798), .ZN(n3889) );
  OAI211_X1 U3620 ( .C1(n2799), .C2(n2798), .A(n3889), .B(n4348), .ZN(n2810)
         );
  NOR2_X1 U3621 ( .A1(STATE_REG_SCAN_IN), .A2(n2800), .ZN(n3117) );
  INV_X1 U3622 ( .A(n2801), .ZN(n2804) );
  INV_X1 U3623 ( .A(n2802), .ZN(n4248) );
  INV_X1 U3624 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2805) );
  MUX2_X1 U3625 ( .A(n2805), .B(REG1_REG_9__SCAN_IN), .S(n3873), .Z(n2806) );
  AOI211_X1 U3626 ( .C1(n2807), .C2(n2806), .A(n3872), .B(n4433), .ZN(n2808)
         );
  AOI211_X1 U3627 ( .C1(n4442), .C2(ADDR_REG_9__SCAN_IN), .A(n3117), .B(n2808), 
        .ZN(n2809) );
  OAI211_X1 U3628 ( .C1(n4445), .C2(n3890), .A(n2810), .B(n2809), .ZN(U3249)
         );
  NAND2_X1 U3629 ( .A1(n3832), .A2(n3458), .ZN(n2812) );
  NAND2_X1 U3630 ( .A1(n2848), .A2(n3435), .ZN(n2811) );
  NAND2_X1 U3631 ( .A1(n2812), .A2(n2811), .ZN(n2814) );
  NAND2_X1 U3632 ( .A1(n3832), .A2(n3459), .ZN(n2816) );
  NAND2_X1 U3633 ( .A1(n3458), .A2(n2848), .ZN(n2815) );
  NAND2_X1 U3634 ( .A1(n2816), .A2(n2815), .ZN(n2864) );
  XNOR2_X1 U3635 ( .A(n2863), .B(n2864), .ZN(n2833) );
  NAND2_X1 U3636 ( .A1(n2817), .A2(n3451), .ZN(n2818) );
  NAND2_X1 U3637 ( .A1(n2819), .A2(n2818), .ZN(n3546) );
  NAND2_X1 U3638 ( .A1(n3544), .A2(n3435), .ZN(n2821) );
  NAND2_X1 U3639 ( .A1(n2822), .A2(n2821), .ZN(n2823) );
  XNOR2_X1 U3640 ( .A(n2823), .B(n3451), .ZN(n2827) );
  NAND2_X1 U3641 ( .A1(n3834), .A2(n2824), .ZN(n2826) );
  NAND2_X1 U3642 ( .A1(n3544), .A2(n3458), .ZN(n2825) );
  NAND2_X1 U3643 ( .A1(n2826), .A2(n2825), .ZN(n2828) );
  XNOR2_X1 U3644 ( .A(n2827), .B(n2828), .ZN(n3547) );
  NAND2_X1 U3645 ( .A1(n3546), .A2(n3547), .ZN(n3545) );
  INV_X1 U3646 ( .A(n2827), .ZN(n2829) );
  NAND2_X1 U3647 ( .A1(n2829), .A2(n2828), .ZN(n2830) );
  NAND2_X1 U3648 ( .A1(n3545), .A2(n2830), .ZN(n2831) );
  INV_X1 U3649 ( .A(n2868), .ZN(n2832) );
  AOI21_X1 U3650 ( .B1(n2833), .B2(n2831), .A(n2832), .ZN(n2837) );
  NAND2_X1 U3651 ( .A1(n2834), .A2(n4254), .ZN(n3655) );
  INV_X1 U3652 ( .A(n3655), .ZN(n3561) );
  AOI22_X1 U3653 ( .A1(n3636), .A2(n2848), .B1(n3561), .B2(n3834), .ZN(n2836)
         );
  INV_X1 U3654 ( .A(n3654), .ZN(n3560) );
  AOI22_X1 U3655 ( .A1(n3548), .A2(REG3_REG_2__SCAN_IN), .B1(n3560), .B2(n3831), .ZN(n2835) );
  OAI211_X1 U3656 ( .C1(n2837), .C2(n3664), .A(n2836), .B(n2835), .ZN(U3234)
         );
  OAI21_X1 U3657 ( .B1(n2839), .B2(n2842), .A(n2838), .ZN(n2924) );
  INV_X1 U3658 ( .A(n4109), .ZN(n3303) );
  AOI22_X1 U3659 ( .A1(n3831), .A2(n4025), .B1(n2848), .B2(n4127), .ZN(n2840)
         );
  OAI21_X1 U3660 ( .B1(n2730), .B2(n3303), .A(n2840), .ZN(n2846) );
  AOI21_X1 U3661 ( .B1(n2844), .B2(n2843), .A(n4104), .ZN(n2845) );
  AOI211_X1 U3662 ( .C1(n2978), .C2(n2924), .A(n2846), .B(n2845), .ZN(n2927)
         );
  INV_X1 U3663 ( .A(n2927), .ZN(n2847) );
  AOI21_X1 U3664 ( .B1(n4402), .B2(n2924), .A(n2847), .ZN(n2853) );
  INV_X1 U3665 ( .A(n4188), .ZN(n3223) );
  AND2_X1 U3666 ( .A1(n2849), .A2(n2848), .ZN(n2850) );
  NOR2_X1 U3667 ( .A1(n3025), .A2(n2850), .ZN(n2929) );
  AOI22_X1 U3668 ( .A1(n3223), .A2(n2929), .B1(REG1_REG_2__SCAN_IN), .B2(n4430), .ZN(n2851) );
  OAI21_X1 U3669 ( .B1(n2853), .B2(n4430), .A(n2851), .ZN(U3520) );
  INV_X1 U3670 ( .A(n4236), .ZN(n3227) );
  AOI22_X1 U3671 ( .A1(n3227), .A2(n2929), .B1(n4422), .B2(REG0_REG_2__SCAN_IN), .ZN(n2852) );
  OAI21_X1 U3672 ( .B1(n2853), .B2(n4422), .A(n2852), .ZN(U3471) );
  OAI21_X1 U3673 ( .B1(n2855), .B2(n2854), .A(STATE_REG_SCAN_IN), .ZN(n2857)
         );
  INV_X1 U3674 ( .A(n3661), .ZN(n3144) );
  NAND2_X1 U3675 ( .A1(n3831), .A2(n3458), .ZN(n2859) );
  NAND2_X1 U3676 ( .A1(n3018), .A2(n3321), .ZN(n2858) );
  NAND2_X1 U3677 ( .A1(n2859), .A2(n2858), .ZN(n2860) );
  XNOR2_X1 U3678 ( .A(n2860), .B(n3451), .ZN(n2898) );
  NAND2_X1 U3679 ( .A1(n3831), .A2(n3459), .ZN(n2862) );
  NAND2_X1 U3680 ( .A1(n3444), .A2(n3018), .ZN(n2861) );
  NAND2_X1 U3681 ( .A1(n2862), .A2(n2861), .ZN(n2896) );
  XNOR2_X1 U3682 ( .A(n2898), .B(n2896), .ZN(n2894) );
  INV_X1 U3683 ( .A(n2863), .ZN(n2866) );
  INV_X1 U3684 ( .A(n2864), .ZN(n2865) );
  NAND2_X1 U3685 ( .A1(n2866), .A2(n2865), .ZN(n2867) );
  XNOR2_X1 U3686 ( .A(n2894), .B(n2895), .ZN(n2869) );
  INV_X1 U3687 ( .A(n3664), .ZN(n3557) );
  NAND2_X1 U3688 ( .A1(n2869), .A2(n3557), .ZN(n2873) );
  OAI22_X1 U3689 ( .A1(n3020), .A2(n3655), .B1(n3654), .B2(n2937), .ZN(n2870)
         );
  AOI211_X1 U3690 ( .C1(n3018), .C2(n3636), .A(n2871), .B(n2870), .ZN(n2872)
         );
  OAI211_X1 U3691 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3144), .A(n2873), .B(n2872), 
        .ZN(U3215) );
  NAND2_X1 U3692 ( .A1(n3833), .A2(DATAO_REG_29__SCAN_IN), .ZN(n2874) );
  OAI21_X1 U3693 ( .B1(n3699), .B2(n3833), .A(n2874), .ZN(U3579) );
  INV_X1 U3694 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4475) );
  NAND2_X1 U3695 ( .A1(n3481), .A2(U4043), .ZN(n2875) );
  OAI21_X1 U3696 ( .B1(U4043), .B2(n4475), .A(n2875), .ZN(U3576) );
  XNOR2_X1 U3697 ( .A(n2876), .B(n3757), .ZN(n2879) );
  AOI22_X1 U3698 ( .A1(n3827), .A2(n4025), .B1(n4127), .B2(n3003), .ZN(n2877)
         );
  OAI21_X1 U3699 ( .B1(n3000), .B2(n3303), .A(n2877), .ZN(n2878) );
  AOI21_X1 U3700 ( .B1(n2879), .B2(n4032), .A(n2878), .ZN(n4414) );
  NAND3_X1 U3701 ( .A1(n2882), .A2(n2881), .A3(n2880), .ZN(n2883) );
  NAND2_X2 U3702 ( .A1(n2883), .A2(n4352), .ZN(n4263) );
  OAI211_X1 U3703 ( .C1(n2983), .C2(n2884), .A(n4421), .B(n3038), .ZN(n4413)
         );
  INV_X1 U3704 ( .A(n4413), .ZN(n2888) );
  INV_X1 U3705 ( .A(n3004), .ZN(n2885) );
  OAI22_X1 U3706 ( .A1(n4263), .A2(n2886), .B1(n2885), .B2(n4352), .ZN(n2887)
         );
  AOI21_X1 U3707 ( .B1(n2888), .B2(n4116), .A(n2887), .ZN(n2893) );
  NAND2_X1 U3708 ( .A1(n2890), .A2(n3757), .ZN(n4411) );
  OR2_X1 U3709 ( .A1(n2767), .A2(n3908), .ZN(n2925) );
  NAND2_X1 U3710 ( .A1(n4065), .A2(n2925), .ZN(n2891) );
  NAND3_X1 U3711 ( .A1(n2889), .A2(n4411), .A3(n4121), .ZN(n2892) );
  OAI211_X1 U3712 ( .C1(n4414), .C2(n2009), .A(n2893), .B(n2892), .ZN(U3283)
         );
  INV_X1 U3713 ( .A(n2942), .ZN(n2923) );
  INV_X1 U3714 ( .A(n2896), .ZN(n2897) );
  NAND2_X1 U3715 ( .A1(n2898), .A2(n2897), .ZN(n2899) );
  NAND2_X1 U3716 ( .A1(n2900), .A2(n2899), .ZN(n2948) );
  INV_X1 U3717 ( .A(n2948), .ZN(n2908) );
  NAND2_X1 U3718 ( .A1(n3830), .A2(n3458), .ZN(n2902) );
  NAND2_X1 U3719 ( .A1(n3490), .A2(n3321), .ZN(n2901) );
  NAND2_X1 U3720 ( .A1(n2902), .A2(n2901), .ZN(n2904) );
  XNOR2_X1 U3721 ( .A(n2904), .B(n2903), .ZN(n2910) );
  NAND2_X1 U3722 ( .A1(n3830), .A2(n3203), .ZN(n2906) );
  NAND2_X1 U3723 ( .A1(n3444), .A2(n3490), .ZN(n2905) );
  NAND2_X1 U3724 ( .A1(n2906), .A2(n2905), .ZN(n2909) );
  XNOR2_X1 U3725 ( .A(n2910), .B(n2909), .ZN(n2949) );
  NAND2_X1 U3726 ( .A1(n2908), .A2(n2907), .ZN(n2946) );
  NAND2_X1 U3727 ( .A1(n2910), .A2(n2909), .ZN(n2911) );
  NAND2_X1 U3728 ( .A1(n2946), .A2(n2911), .ZN(n2918) );
  NAND2_X1 U3729 ( .A1(n3829), .A2(n3458), .ZN(n2913) );
  NAND2_X1 U3730 ( .A1(n2941), .A2(n3321), .ZN(n2912) );
  NAND2_X1 U3731 ( .A1(n2913), .A2(n2912), .ZN(n2914) );
  XNOR2_X1 U3732 ( .A(n2914), .B(n3451), .ZN(n2954) );
  NAND2_X1 U3733 ( .A1(n3829), .A2(n3203), .ZN(n2916) );
  NAND2_X1 U3734 ( .A1(n2941), .A2(n3458), .ZN(n2915) );
  NAND2_X1 U3735 ( .A1(n2916), .A2(n2915), .ZN(n2955) );
  XNOR2_X1 U3736 ( .A(n2954), .B(n2955), .ZN(n2917) );
  NAND2_X1 U3737 ( .A1(n2918), .A2(n2917), .ZN(n2958) );
  OAI211_X1 U3738 ( .C1(n2918), .C2(n2917), .A(n2958), .B(n3557), .ZN(n2922)
         );
  OAI22_X1 U3739 ( .A1(n2937), .A2(n3655), .B1(n3654), .B2(n3000), .ZN(n2919)
         );
  AOI211_X1 U3740 ( .C1(n2941), .C2(n3636), .A(n2920), .B(n2919), .ZN(n2921)
         );
  OAI211_X1 U3741 ( .C1(n3144), .C2(n2923), .A(n2922), .B(n2921), .ZN(U3224)
         );
  INV_X1 U3742 ( .A(n2924), .ZN(n2932) );
  INV_X1 U3743 ( .A(n2925), .ZN(n2926) );
  AND2_X1 U3744 ( .A1(n4263), .A2(n2926), .ZN(n4368) );
  INV_X1 U3745 ( .A(n4368), .ZN(n3504) );
  MUX2_X1 U3746 ( .A(n2928), .B(n2927), .S(n4263), .Z(n2931) );
  AOI22_X1 U3747 ( .A1(n4358), .A2(n2929), .B1(REG3_REG_2__SCAN_IN), .B2(n4367), .ZN(n2930) );
  OAI211_X1 U3748 ( .C1(n2932), .C2(n3504), .A(n2931), .B(n2930), .ZN(U3288)
         );
  INV_X1 U3749 ( .A(n2933), .ZN(n3753) );
  NAND2_X1 U3750 ( .A1(n3753), .A2(n3762), .ZN(n3712) );
  XNOR2_X1 U3751 ( .A(n2934), .B(n3712), .ZN(n4404) );
  XNOR2_X1 U3752 ( .A(n2935), .B(n3712), .ZN(n2939) );
  AOI22_X1 U3753 ( .A1(n3828), .A2(n4025), .B1(n2941), .B2(n4127), .ZN(n2936)
         );
  OAI21_X1 U3754 ( .B1(n2937), .B2(n3303), .A(n2936), .ZN(n2938) );
  AOI21_X1 U3755 ( .B1(n2939), .B2(n4032), .A(n2938), .ZN(n4405) );
  MUX2_X1 U3756 ( .A(n4405), .B(n2940), .S(n2009), .Z(n2944) );
  AOI21_X1 U3757 ( .B1(n2941), .B2(n3497), .A(n2981), .ZN(n4408) );
  AOI22_X1 U3758 ( .A1(n4408), .A2(n4358), .B1(n2942), .B2(n4367), .ZN(n2943)
         );
  OAI211_X1 U3759 ( .C1(n4098), .C2(n4404), .A(n2944), .B(n2943), .ZN(U3285)
         );
  AOI22_X1 U3760 ( .A1(n3560), .A2(n3829), .B1(n3561), .B2(n3831), .ZN(n2945)
         );
  NAND2_X1 U3761 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3864) );
  OAI211_X1 U3762 ( .C1(n3658), .C2(n3498), .A(n2945), .B(n3864), .ZN(n2951)
         );
  INV_X1 U3763 ( .A(n2946), .ZN(n2947) );
  AOI211_X1 U3764 ( .C1(n2949), .C2(n2948), .A(n3664), .B(n2947), .ZN(n2950)
         );
  AOI211_X1 U3765 ( .C1(n2952), .C2(n3661), .A(n2951), .B(n2950), .ZN(n2953)
         );
  INV_X1 U3766 ( .A(n2953), .ZN(U3227) );
  INV_X1 U3767 ( .A(n2954), .ZN(n2956) );
  NAND2_X1 U3768 ( .A1(n2956), .A2(n2955), .ZN(n2957) );
  NAND2_X1 U3769 ( .A1(n3828), .A2(n3203), .ZN(n2960) );
  NAND2_X1 U3770 ( .A1(n3444), .A2(n2973), .ZN(n2959) );
  NAND2_X1 U3771 ( .A1(n2960), .A2(n2959), .ZN(n2992) );
  NAND2_X1 U3772 ( .A1(n3828), .A2(n3458), .ZN(n2962) );
  NAND2_X1 U3773 ( .A1(n2973), .A2(n3321), .ZN(n2961) );
  NAND2_X1 U3774 ( .A1(n2962), .A2(n2961), .ZN(n2963) );
  XNOR2_X1 U3775 ( .A(n2963), .B(n2903), .ZN(n2991) );
  XOR2_X1 U3776 ( .A(n2992), .B(n2991), .Z(n2964) );
  XNOR2_X1 U3777 ( .A(n2993), .B(n2964), .ZN(n2970) );
  OAI22_X1 U3778 ( .A1(n3078), .A2(n3654), .B1(n3655), .B2(n2965), .ZN(n2966)
         );
  AOI211_X1 U3779 ( .C1(n2973), .C2(n3636), .A(n2967), .B(n2966), .ZN(n2969)
         );
  NAND2_X1 U3780 ( .A1(n3661), .A2(n4351), .ZN(n2968) );
  OAI211_X1 U3781 ( .C1(n2970), .C2(n3664), .A(n2969), .B(n2968), .ZN(U3236)
         );
  NAND2_X1 U3782 ( .A1(n3756), .A2(n3761), .ZN(n3718) );
  XOR2_X1 U3783 ( .A(n2971), .B(n3718), .Z(n4359) );
  INV_X1 U3784 ( .A(n4359), .ZN(n2979) );
  XNOR2_X1 U3785 ( .A(n2972), .B(n3718), .ZN(n2976) );
  AOI22_X1 U3786 ( .A1(n2997), .A2(n4025), .B1(n2973), .B2(n4127), .ZN(n2975)
         );
  NAND2_X1 U3787 ( .A1(n3829), .A2(n4109), .ZN(n2974) );
  OAI211_X1 U3788 ( .C1(n2976), .C2(n4104), .A(n2975), .B(n2974), .ZN(n2977)
         );
  AOI21_X1 U3789 ( .B1(n2978), .B2(n4359), .A(n2977), .ZN(n4362) );
  OAI21_X1 U3790 ( .B1(n4394), .B2(n2979), .A(n4362), .ZN(n2989) );
  NOR2_X1 U3791 ( .A1(n2981), .A2(n2980), .ZN(n2982) );
  OR2_X1 U3792 ( .A1(n2983), .A2(n2982), .ZN(n4356) );
  INV_X1 U3793 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2984) );
  OAI22_X1 U3794 ( .A1(n4356), .A2(n4188), .B1(n4432), .B2(n2984), .ZN(n2985)
         );
  AOI21_X1 U3795 ( .B1(n2989), .B2(n4432), .A(n2985), .ZN(n2986) );
  INV_X1 U3796 ( .A(n2986), .ZN(U3524) );
  INV_X1 U3797 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2987) );
  OAI22_X1 U3798 ( .A1(n4356), .A2(n4236), .B1(n4423), .B2(n2987), .ZN(n2988)
         );
  AOI21_X1 U3799 ( .B1(n2989), .B2(n4423), .A(n2988), .ZN(n2990) );
  INV_X1 U3800 ( .A(n2990), .ZN(U3479) );
  NAND2_X1 U3801 ( .A1(n2997), .A2(n3458), .ZN(n2995) );
  NAND2_X1 U3802 ( .A1(n3003), .A2(n3321), .ZN(n2994) );
  NAND2_X1 U3803 ( .A1(n2995), .A2(n2994), .ZN(n2996) );
  XNOR2_X1 U3804 ( .A(n2996), .B(n3451), .ZN(n3061) );
  NAND2_X1 U3805 ( .A1(n2997), .A2(n3203), .ZN(n2999) );
  NAND2_X1 U3806 ( .A1(n3444), .A2(n3003), .ZN(n2998) );
  NAND2_X1 U3807 ( .A1(n2999), .A2(n2998), .ZN(n3062) );
  XNOR2_X1 U3808 ( .A(n3061), .B(n3062), .ZN(n3059) );
  XNOR2_X1 U3809 ( .A(n3060), .B(n3059), .ZN(n3007) );
  OAI22_X1 U3810 ( .A1(n3000), .A2(n3655), .B1(n3654), .B2(n3115), .ZN(n3001)
         );
  AOI211_X1 U3811 ( .C1(n3003), .C2(n3636), .A(n3002), .B(n3001), .ZN(n3006)
         );
  NAND2_X1 U3812 ( .A1(n3661), .A2(n3004), .ZN(n3005) );
  OAI211_X1 U3813 ( .C1(n3007), .C2(n3664), .A(n3006), .B(n3005), .ZN(U3210)
         );
  INV_X1 U3814 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3008) );
  OAI22_X1 U3815 ( .A1(n4095), .A2(n3009), .B1(n3008), .B2(n4352), .ZN(n3012)
         );
  MUX2_X1 U3816 ( .A(n3010), .B(REG2_REG_1__SCAN_IN), .S(n2009), .Z(n3011) );
  AOI211_X1 U3817 ( .C1(n4368), .C2(n3013), .A(n3012), .B(n3011), .ZN(n3014)
         );
  INV_X1 U3818 ( .A(n3014), .ZN(U3289) );
  XNOR2_X1 U3819 ( .A(n3015), .B(n3714), .ZN(n4395) );
  OAI21_X1 U3820 ( .B1(n3714), .B2(n3017), .A(n3016), .ZN(n3022) );
  AOI22_X1 U3821 ( .A1(n3830), .A2(n4025), .B1(n4127), .B2(n3018), .ZN(n3019)
         );
  OAI21_X1 U3822 ( .B1(n3020), .B2(n3303), .A(n3019), .ZN(n3021) );
  AOI21_X1 U3823 ( .B1(n3022), .B2(n4032), .A(n3021), .ZN(n3023) );
  OAI21_X1 U3824 ( .B1(n4395), .B2(n4065), .A(n3023), .ZN(n4397) );
  INV_X1 U3825 ( .A(n4397), .ZN(n3030) );
  INV_X1 U3826 ( .A(n4395), .ZN(n3028) );
  OAI21_X1 U3827 ( .B1(n3025), .B2(n3024), .A(n3496), .ZN(n4392) );
  AOI22_X1 U3828 ( .A1(n2009), .A2(REG2_REG_3__SCAN_IN), .B1(n4367), .B2(n2272), .ZN(n3026) );
  OAI21_X1 U3829 ( .B1(n4095), .B2(n4392), .A(n3026), .ZN(n3027) );
  AOI21_X1 U3830 ( .B1(n3028), .B2(n4368), .A(n3027), .ZN(n3029) );
  OAI21_X1 U3831 ( .B1(n3030), .B2(n2009), .A(n3029), .ZN(U3287) );
  AND2_X1 U3832 ( .A1(n3765), .A2(n3759), .ZN(n3707) );
  XOR2_X1 U3833 ( .A(n3707), .B(n3031), .Z(n3037) );
  XOR2_X1 U3834 ( .A(n3707), .B(n3032), .Z(n3035) );
  AOI22_X1 U3835 ( .A1(n3826), .A2(n4025), .B1(n3081), .B2(n4127), .ZN(n3033)
         );
  OAI21_X1 U3836 ( .B1(n3078), .B2(n3303), .A(n3033), .ZN(n3034) );
  AOI21_X1 U3837 ( .B1(n3035), .B2(n4032), .A(n3034), .ZN(n3036) );
  OAI21_X1 U3838 ( .B1(n3037), .B2(n4065), .A(n3036), .ZN(n3099) );
  INV_X1 U3839 ( .A(n3099), .ZN(n3044) );
  INV_X1 U3840 ( .A(n3037), .ZN(n3100) );
  NAND2_X1 U3841 ( .A1(n3038), .A2(n3081), .ZN(n3039) );
  NAND2_X1 U3842 ( .A1(n3053), .A2(n3039), .ZN(n3105) );
  AOI22_X1 U3843 ( .A1(n2009), .A2(REG2_REG_8__SCAN_IN), .B1(n3040), .B2(n4367), .ZN(n3041) );
  OAI21_X1 U3844 ( .B1(n3105), .B2(n4095), .A(n3041), .ZN(n3042) );
  AOI21_X1 U3845 ( .B1(n3100), .B2(n4368), .A(n3042), .ZN(n3043) );
  OAI21_X1 U3846 ( .B1(n3044), .B2(n2009), .A(n3043), .ZN(U3282) );
  INV_X1 U3847 ( .A(n3772), .ZN(n3045) );
  NAND2_X1 U3848 ( .A1(n3045), .A2(n3766), .ZN(n3713) );
  XNOR2_X1 U3849 ( .A(n3046), .B(n3713), .ZN(n4417) );
  XOR2_X1 U3850 ( .A(n3713), .B(n3047), .Z(n3051) );
  OAI22_X1 U3851 ( .A1(n3114), .A2(n4101), .B1(n4134), .B2(n3048), .ZN(n3049)
         );
  AOI21_X1 U3852 ( .B1(n4109), .B2(n3827), .A(n3049), .ZN(n3050) );
  OAI21_X1 U3853 ( .B1(n3051), .B2(n4104), .A(n3050), .ZN(n4418) );
  NAND2_X1 U3854 ( .A1(n4418), .A2(n4263), .ZN(n3058) );
  INV_X1 U3855 ( .A(n3052), .ZN(n3092) );
  AOI21_X1 U3856 ( .B1(n3118), .B2(n3053), .A(n3092), .ZN(n4420) );
  INV_X1 U3857 ( .A(n3119), .ZN(n3054) );
  OAI22_X1 U3858 ( .A1(n4263), .A2(n3055), .B1(n3054), .B2(n4352), .ZN(n3056)
         );
  AOI21_X1 U3859 ( .B1(n4420), .B2(n4358), .A(n3056), .ZN(n3057) );
  OAI211_X1 U3860 ( .C1(n4417), .C2(n4098), .A(n3058), .B(n3057), .ZN(U3281)
         );
  INV_X1 U3861 ( .A(n3061), .ZN(n3063) );
  NAND2_X1 U3862 ( .A1(n3063), .A2(n3062), .ZN(n3064) );
  NAND2_X1 U3863 ( .A1(n3065), .A2(n3064), .ZN(n3108) );
  NAND2_X1 U3864 ( .A1(n3827), .A2(n3458), .ZN(n3067) );
  NAND2_X1 U3865 ( .A1(n3081), .A2(n3321), .ZN(n3066) );
  NAND2_X1 U3866 ( .A1(n3067), .A2(n3066), .ZN(n3068) );
  XNOR2_X1 U3867 ( .A(n3068), .B(n2903), .ZN(n3071) );
  NAND2_X1 U3868 ( .A1(n3827), .A2(n3203), .ZN(n3070) );
  NAND2_X1 U3869 ( .A1(n3081), .A2(n3458), .ZN(n3069) );
  NAND2_X1 U3870 ( .A1(n3070), .A2(n3069), .ZN(n3072) );
  AND2_X1 U3871 ( .A1(n3071), .A2(n3072), .ZN(n3107) );
  INV_X1 U3872 ( .A(n3107), .ZN(n3075) );
  INV_X1 U3873 ( .A(n3071), .ZN(n3074) );
  INV_X1 U3874 ( .A(n3072), .ZN(n3073) );
  NAND2_X1 U3875 ( .A1(n3074), .A2(n3073), .ZN(n3106) );
  NAND2_X1 U3876 ( .A1(n3075), .A2(n3106), .ZN(n3076) );
  XNOR2_X1 U3877 ( .A(n3108), .B(n3076), .ZN(n3077) );
  NAND2_X1 U3878 ( .A1(n3077), .A2(n3557), .ZN(n3083) );
  OAI22_X1 U3879 ( .A1(n3138), .A2(n3654), .B1(n3655), .B2(n3078), .ZN(n3079)
         );
  AOI211_X1 U3880 ( .C1(n3081), .C2(n3636), .A(n3080), .B(n3079), .ZN(n3082)
         );
  OAI211_X1 U3881 ( .C1(n3144), .C2(n3084), .A(n3083), .B(n3082), .ZN(U3218)
         );
  AND2_X1 U3882 ( .A1(n3771), .A2(n3774), .ZN(n3708) );
  XOR2_X1 U3883 ( .A(n3708), .B(n3085), .Z(n3088) );
  OAI22_X1 U3884 ( .A1(n3212), .A2(n4101), .B1(n4134), .B2(n3091), .ZN(n3086)
         );
  AOI21_X1 U3885 ( .B1(n4109), .B2(n3826), .A(n3086), .ZN(n3087) );
  OAI21_X1 U3886 ( .B1(n3088), .B2(n4104), .A(n3087), .ZN(n3158) );
  INV_X1 U3887 ( .A(n3158), .ZN(n3098) );
  XOR2_X1 U3888 ( .A(n3708), .B(n3089), .Z(n3159) );
  INV_X1 U3889 ( .A(n3190), .ZN(n3090) );
  OAI21_X1 U3890 ( .B1(n3092), .B2(n3091), .A(n3090), .ZN(n3164) );
  NOR2_X1 U3891 ( .A1(n3164), .A2(n4095), .ZN(n3096) );
  INV_X1 U3892 ( .A(n3093), .ZN(n3143) );
  OAI22_X1 U3893 ( .A1(n4263), .A2(n3094), .B1(n3143), .B2(n4352), .ZN(n3095)
         );
  AOI211_X1 U3894 ( .C1(n3159), .C2(n4121), .A(n3096), .B(n3095), .ZN(n3097)
         );
  OAI21_X1 U3895 ( .B1(n3098), .B2(n2009), .A(n3097), .ZN(U3280) );
  INV_X1 U3896 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3101) );
  AOI21_X1 U3897 ( .B1(n4402), .B2(n3100), .A(n3099), .ZN(n3103) );
  MUX2_X1 U3898 ( .A(n3101), .B(n3103), .S(n4423), .Z(n3102) );
  OAI21_X1 U3899 ( .B1(n3105), .B2(n4236), .A(n3102), .ZN(U3483) );
  MUX2_X1 U3900 ( .A(n4453), .B(n3103), .S(n4432), .Z(n3104) );
  OAI21_X1 U3901 ( .B1(n3105), .B2(n4188), .A(n3104), .ZN(U3526) );
  OAI21_X1 U3902 ( .B1(n3108), .B2(n3107), .A(n3106), .ZN(n3124) );
  NAND2_X1 U3903 ( .A1(n3826), .A2(n3444), .ZN(n3110) );
  NAND2_X1 U3904 ( .A1(n3118), .A2(n3321), .ZN(n3109) );
  NAND2_X1 U3905 ( .A1(n3110), .A2(n3109), .ZN(n3111) );
  XNOR2_X1 U3906 ( .A(n3111), .B(n3451), .ZN(n3127) );
  NAND2_X1 U3907 ( .A1(n3826), .A2(n3203), .ZN(n3113) );
  NAND2_X1 U3908 ( .A1(n3444), .A2(n3118), .ZN(n3112) );
  NAND2_X1 U3909 ( .A1(n3113), .A2(n3112), .ZN(n3125) );
  XNOR2_X1 U3910 ( .A(n3127), .B(n3125), .ZN(n3123) );
  XOR2_X1 U3911 ( .A(n3124), .B(n3123), .Z(n3122) );
  OAI22_X1 U3912 ( .A1(n3115), .A2(n3655), .B1(n3654), .B2(n3114), .ZN(n3116)
         );
  AOI211_X1 U3913 ( .C1(n3118), .C2(n3636), .A(n3117), .B(n3116), .ZN(n3121)
         );
  NAND2_X1 U3914 ( .A1(n3661), .A2(n3119), .ZN(n3120) );
  OAI211_X1 U3915 ( .C1(n3122), .C2(n3664), .A(n3121), .B(n3120), .ZN(U3228)
         );
  INV_X1 U3916 ( .A(n3125), .ZN(n3126) );
  NAND2_X1 U3917 ( .A1(n3127), .A2(n3126), .ZN(n3128) );
  NAND2_X1 U3918 ( .A1(n3825), .A2(n3444), .ZN(n3130) );
  NAND2_X1 U3919 ( .A1(n3140), .A2(n3321), .ZN(n3129) );
  NAND2_X1 U3920 ( .A1(n3130), .A2(n3129), .ZN(n3131) );
  XNOR2_X1 U3921 ( .A(n3131), .B(n2903), .ZN(n3166) );
  NAND2_X1 U3922 ( .A1(n3825), .A2(n3203), .ZN(n3133) );
  NAND2_X1 U3923 ( .A1(n3444), .A2(n3140), .ZN(n3132) );
  NAND2_X1 U3924 ( .A1(n3133), .A2(n3132), .ZN(n3165) );
  XNOR2_X1 U3925 ( .A(n3166), .B(n3165), .ZN(n3135) );
  AOI21_X1 U3926 ( .B1(n3134), .B2(n3135), .A(n3664), .ZN(n3137) );
  NAND2_X1 U3927 ( .A1(n3137), .A2(n3168), .ZN(n3142) );
  AND2_X1 U3928 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n4268) );
  OAI22_X1 U3929 ( .A1(n3138), .A2(n3655), .B1(n3654), .B2(n3212), .ZN(n3139)
         );
  AOI211_X1 U3930 ( .C1(n3140), .C2(n3636), .A(n4268), .B(n3139), .ZN(n3141)
         );
  OAI211_X1 U3931 ( .C1(n3144), .C2(n3143), .A(n3142), .B(n3141), .ZN(U3214)
         );
  INV_X1 U3932 ( .A(n3264), .ZN(n3145) );
  OR2_X1 U3933 ( .A1(n3145), .A2(n3265), .ZN(n3706) );
  INV_X1 U3934 ( .A(n3706), .ZN(n3146) );
  XNOR2_X1 U3935 ( .A(n3266), .B(n3146), .ZN(n3151) );
  NAND2_X1 U3936 ( .A1(n3824), .A2(n4109), .ZN(n3148) );
  NAND2_X1 U3937 ( .A1(n3822), .A2(n4025), .ZN(n3147) );
  OAI211_X1 U3938 ( .C1(n4134), .C2(n3149), .A(n3148), .B(n3147), .ZN(n3150)
         );
  AOI21_X1 U3939 ( .B1(n3151), .B2(n4032), .A(n3150), .ZN(n3220) );
  XNOR2_X1 U3940 ( .A(n3152), .B(n3706), .ZN(n3219) );
  INV_X1 U3941 ( .A(n3153), .ZN(n3277) );
  AOI21_X1 U3942 ( .B1(n3214), .B2(n3188), .A(n3277), .ZN(n3228) );
  INV_X1 U3943 ( .A(n3228), .ZN(n3155) );
  AOI22_X1 U3944 ( .A1(n2009), .A2(REG2_REG_12__SCAN_IN), .B1(n3215), .B2(
        n4367), .ZN(n3154) );
  OAI21_X1 U3945 ( .B1(n3155), .B2(n4095), .A(n3154), .ZN(n3156) );
  AOI21_X1 U3946 ( .B1(n3219), .B2(n4121), .A(n3156), .ZN(n3157) );
  OAI21_X1 U3947 ( .B1(n2009), .B2(n3220), .A(n3157), .ZN(U3278) );
  INV_X1 U3948 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4266) );
  AOI21_X1 U3949 ( .B1(n4410), .B2(n3159), .A(n3158), .ZN(n3161) );
  MUX2_X1 U3950 ( .A(n4266), .B(n3161), .S(n4432), .Z(n3160) );
  OAI21_X1 U3951 ( .B1(n3164), .B2(n4188), .A(n3160), .ZN(U3528) );
  INV_X1 U3952 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3162) );
  MUX2_X1 U3953 ( .A(n3162), .B(n3161), .S(n4423), .Z(n3163) );
  OAI21_X1 U3954 ( .B1(n3164), .B2(n4236), .A(n3163), .ZN(U3487) );
  NAND2_X1 U3955 ( .A1(n3166), .A2(n3165), .ZN(n3167) );
  NAND2_X1 U3956 ( .A1(n3824), .A2(n3203), .ZN(n3170) );
  NAND2_X1 U3957 ( .A1(n3444), .A2(n3182), .ZN(n3169) );
  NAND2_X1 U3958 ( .A1(n3170), .A2(n3169), .ZN(n3198) );
  NAND2_X1 U3959 ( .A1(n3824), .A2(n3444), .ZN(n3172) );
  NAND2_X1 U3960 ( .A1(n3182), .A2(n3321), .ZN(n3171) );
  NAND2_X1 U3961 ( .A1(n3172), .A2(n3171), .ZN(n3173) );
  XNOR2_X1 U3962 ( .A(n3173), .B(n2903), .ZN(n3197) );
  XOR2_X1 U3963 ( .A(n3198), .B(n3197), .Z(n3174) );
  XNOR2_X1 U3964 ( .A(n3199), .B(n3174), .ZN(n3178) );
  AOI22_X1 U3965 ( .A1(n3561), .A2(n3825), .B1(n3560), .B2(n3823), .ZN(n3175)
         );
  NAND2_X1 U3966 ( .A1(REG3_REG_11__SCAN_IN), .A2(U3149), .ZN(n4277) );
  OAI211_X1 U3967 ( .C1(n3658), .C2(n3189), .A(n3175), .B(n4277), .ZN(n3176)
         );
  AOI21_X1 U3968 ( .B1(n3191), .B2(n3661), .A(n3176), .ZN(n3177) );
  OAI21_X1 U3969 ( .B1(n3178), .B2(n3664), .A(n3177), .ZN(U3233) );
  XNOR2_X1 U3970 ( .A(n3179), .B(n3720), .ZN(n3186) );
  AOI21_X1 U3971 ( .B1(n3720), .B2(n3181), .A(n2212), .ZN(n3187) );
  AOI22_X1 U3972 ( .A1(n3823), .A2(n4025), .B1(n4127), .B2(n3182), .ZN(n3184)
         );
  NAND2_X1 U3973 ( .A1(n3825), .A2(n4109), .ZN(n3183) );
  OAI211_X1 U3974 ( .C1(n3187), .C2(n4065), .A(n3184), .B(n3183), .ZN(n3185)
         );
  AOI21_X1 U3975 ( .B1(n3186), .B2(n4032), .A(n3185), .ZN(n3241) );
  INV_X1 U3976 ( .A(n3187), .ZN(n3243) );
  OAI21_X1 U3977 ( .B1(n3190), .B2(n3189), .A(n3188), .ZN(n3248) );
  NOR2_X1 U3978 ( .A1(n3248), .A2(n4095), .ZN(n3195) );
  INV_X1 U3979 ( .A(n3191), .ZN(n3192) );
  OAI22_X1 U3980 ( .A1(n4263), .A2(n3193), .B1(n3192), .B2(n4352), .ZN(n3194)
         );
  AOI211_X1 U3981 ( .C1(n3243), .C2(n4368), .A(n3195), .B(n3194), .ZN(n3196)
         );
  OAI21_X1 U3982 ( .B1(n3241), .B2(n2009), .A(n3196), .ZN(U3279) );
  NAND2_X1 U3983 ( .A1(n3823), .A2(n3444), .ZN(n3201) );
  NAND2_X1 U3984 ( .A1(n3214), .A2(n3321), .ZN(n3200) );
  NAND2_X1 U3985 ( .A1(n3201), .A2(n3200), .ZN(n3202) );
  XNOR2_X1 U3986 ( .A(n3202), .B(n2903), .ZN(n3209) );
  INV_X1 U3987 ( .A(n3209), .ZN(n3207) );
  NAND2_X1 U3988 ( .A1(n3823), .A2(n3203), .ZN(n3205) );
  NAND2_X1 U3989 ( .A1(n3214), .A2(n3444), .ZN(n3204) );
  NAND2_X1 U3990 ( .A1(n3205), .A2(n3204), .ZN(n3208) );
  INV_X1 U3991 ( .A(n3208), .ZN(n3206) );
  NAND2_X1 U3992 ( .A1(n3207), .A2(n3206), .ZN(n3249) );
  INV_X1 U3993 ( .A(n3249), .ZN(n3210) );
  NOR2_X1 U3994 ( .A1(n3210), .A2(n3250), .ZN(n3211) );
  XNOR2_X1 U3995 ( .A(n3251), .B(n3211), .ZN(n3218) );
  AND2_X1 U3996 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n4288) );
  OAI22_X1 U3997 ( .A1(n3212), .A2(n3655), .B1(n3654), .B2(n3336), .ZN(n3213)
         );
  AOI211_X1 U3998 ( .C1(n3214), .C2(n3636), .A(n4288), .B(n3213), .ZN(n3217)
         );
  NAND2_X1 U3999 ( .A1(n3661), .A2(n3215), .ZN(n3216) );
  OAI211_X1 U4000 ( .C1(n3218), .C2(n3664), .A(n3217), .B(n3216), .ZN(U3221)
         );
  NAND2_X1 U4001 ( .A1(n3219), .A2(n4410), .ZN(n3221) );
  NAND2_X1 U4002 ( .A1(n3221), .A2(n3220), .ZN(n3225) );
  MUX2_X1 U4003 ( .A(REG1_REG_12__SCAN_IN), .B(n3225), .S(n4432), .Z(n3222) );
  AOI21_X1 U4004 ( .B1(n3223), .B2(n3228), .A(n3222), .ZN(n3224) );
  INV_X1 U4005 ( .A(n3224), .ZN(U3530) );
  MUX2_X1 U4006 ( .A(REG0_REG_12__SCAN_IN), .B(n3225), .S(n4423), .Z(n3226) );
  AOI21_X1 U4007 ( .B1(n3228), .B2(n3227), .A(n3226), .ZN(n3229) );
  INV_X1 U4008 ( .A(n3229), .ZN(U3491) );
  XNOR2_X1 U4009 ( .A(n3682), .B(n3711), .ZN(n3232) );
  OAI22_X1 U4010 ( .A1(n3581), .A2(n4101), .B1(n4134), .B2(n3235), .ZN(n3230)
         );
  AOI21_X1 U4011 ( .B1(n4109), .B2(n3822), .A(n3230), .ZN(n3231) );
  OAI21_X1 U4012 ( .B1(n3232), .B2(n4104), .A(n3231), .ZN(n3284) );
  INV_X1 U4013 ( .A(n3284), .ZN(n3240) );
  OAI21_X1 U4014 ( .B1(n3234), .B2(n3711), .A(n3233), .ZN(n3285) );
  NOR2_X1 U4015 ( .A1(n3274), .A2(n3235), .ZN(n3236) );
  OR2_X1 U4016 ( .A1(n3344), .A2(n3236), .ZN(n3290) );
  AOI22_X1 U4017 ( .A1(n2009), .A2(REG2_REG_14__SCAN_IN), .B1(n3339), .B2(
        n4367), .ZN(n3237) );
  OAI21_X1 U4018 ( .B1(n3290), .B2(n4095), .A(n3237), .ZN(n3238) );
  AOI21_X1 U4019 ( .B1(n3285), .B2(n4121), .A(n3238), .ZN(n3239) );
  OAI21_X1 U4020 ( .B1(n2009), .B2(n3240), .A(n3239), .ZN(U3276) );
  INV_X1 U4021 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4548) );
  INV_X1 U4022 ( .A(n3241), .ZN(n3242) );
  AOI21_X1 U4023 ( .B1(n4402), .B2(n3243), .A(n3242), .ZN(n3245) );
  MUX2_X1 U4024 ( .A(n4548), .B(n3245), .S(n4432), .Z(n3244) );
  OAI21_X1 U4025 ( .B1(n4188), .B2(n3248), .A(n3244), .ZN(U3529) );
  INV_X1 U4026 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3246) );
  MUX2_X1 U4027 ( .A(n3246), .B(n3245), .S(n4423), .Z(n3247) );
  OAI21_X1 U4028 ( .B1(n3248), .B2(n4236), .A(n3247), .ZN(U3489) );
  NAND2_X1 U4029 ( .A1(n3822), .A2(n3203), .ZN(n3253) );
  NAND2_X1 U4030 ( .A1(n3268), .A2(n3458), .ZN(n3252) );
  NAND2_X1 U4031 ( .A1(n3253), .A2(n3252), .ZN(n3314) );
  NAND2_X1 U4032 ( .A1(n3822), .A2(n3444), .ZN(n3255) );
  NAND2_X1 U4033 ( .A1(n3268), .A2(n3321), .ZN(n3254) );
  NAND2_X1 U4034 ( .A1(n3255), .A2(n3254), .ZN(n3256) );
  XNOR2_X1 U4035 ( .A(n3256), .B(n3451), .ZN(n3317) );
  XOR2_X1 U4036 ( .A(n3314), .B(n3317), .Z(n3257) );
  XNOR2_X1 U4037 ( .A(n3316), .B(n3257), .ZN(n3262) );
  AOI22_X1 U4038 ( .A1(n3561), .A2(n3823), .B1(n3560), .B2(n3352), .ZN(n3258)
         );
  NAND2_X1 U4039 ( .A1(REG3_REG_13__SCAN_IN), .A2(U3149), .ZN(n4297) );
  OAI211_X1 U4040 ( .C1(n3658), .C2(n3276), .A(n3258), .B(n4297), .ZN(n3259)
         );
  AOI21_X1 U4041 ( .B1(n3260), .B2(n3661), .A(n3259), .ZN(n3261) );
  OAI21_X1 U4042 ( .B1(n3262), .B2(n3664), .A(n3261), .ZN(U3231) );
  XNOR2_X1 U40430 ( .A(n3822), .B(n3276), .ZN(n3735) );
  XOR2_X1 U4044 ( .A(n3735), .B(n3263), .Z(n3306) );
  OAI21_X1 U4045 ( .B1(n3266), .B2(n3265), .A(n3264), .ZN(n3267) );
  XNOR2_X1 U4046 ( .A(n3267), .B(n3735), .ZN(n3272) );
  AOI22_X1 U4047 ( .A1(n3352), .A2(n4025), .B1(n3268), .B2(n4127), .ZN(n3269)
         );
  OAI21_X1 U4048 ( .B1(n3270), .B2(n3303), .A(n3269), .ZN(n3271) );
  AOI21_X1 U4049 ( .B1(n3272), .B2(n4032), .A(n3271), .ZN(n3273) );
  OAI21_X1 U4050 ( .B1(n3306), .B2(n4065), .A(n3273), .ZN(n3307) );
  NAND2_X1 U4051 ( .A1(n3307), .A2(n4263), .ZN(n3283) );
  INV_X1 U4052 ( .A(n3274), .ZN(n3275) );
  OAI21_X1 U4053 ( .B1(n3277), .B2(n3276), .A(n3275), .ZN(n3313) );
  INV_X1 U4054 ( .A(n3313), .ZN(n3281) );
  OAI22_X1 U4055 ( .A1(n4263), .A2(n3279), .B1(n3278), .B2(n4352), .ZN(n3280)
         );
  AOI21_X1 U4056 ( .B1(n3281), .B2(n4358), .A(n3280), .ZN(n3282) );
  OAI211_X1 U4057 ( .C1(n3306), .C2(n3504), .A(n3283), .B(n3282), .ZN(U3277)
         );
  INV_X1 U4058 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3286) );
  AOI21_X1 U4059 ( .B1(n3285), .B2(n4410), .A(n3284), .ZN(n3288) );
  MUX2_X1 U4060 ( .A(n3286), .B(n3288), .S(n4423), .Z(n3287) );
  OAI21_X1 U4061 ( .B1(n3290), .B2(n4236), .A(n3287), .ZN(U3495) );
  INV_X1 U4062 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4436) );
  MUX2_X1 U4063 ( .A(n4436), .B(n3288), .S(n4432), .Z(n3289) );
  OAI21_X1 U4064 ( .B1(n4188), .B2(n3290), .A(n3289), .ZN(U3532) );
  OAI21_X1 U4065 ( .B1(n3292), .B2(n3719), .A(n3291), .ZN(n4192) );
  INV_X1 U4066 ( .A(n3293), .ZN(n3361) );
  AOI21_X1 U4067 ( .B1(n3583), .B2(n3294), .A(n3361), .ZN(n4190) );
  INV_X1 U4068 ( .A(n3584), .ZN(n3295) );
  OAI22_X1 U4069 ( .A1(n4263), .A2(n3296), .B1(n3295), .B2(n4352), .ZN(n3297)
         );
  AOI21_X1 U4070 ( .B1(n4190), .B2(n4358), .A(n3297), .ZN(n3305) );
  OAI211_X1 U4071 ( .C1(n3300), .C2(n3299), .A(n3298), .B(n4032), .ZN(n3302)
         );
  AOI22_X1 U4072 ( .A1(n4108), .A2(n4025), .B1(n4127), .B2(n3583), .ZN(n3301)
         );
  OAI211_X1 U4073 ( .C1(n3581), .C2(n3303), .A(n3302), .B(n3301), .ZN(n4189)
         );
  NAND2_X1 U4074 ( .A1(n4189), .A2(n4263), .ZN(n3304) );
  OAI211_X1 U4075 ( .C1(n4192), .C2(n4098), .A(n3305), .B(n3304), .ZN(U3274)
         );
  INV_X1 U4076 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3878) );
  INV_X1 U4077 ( .A(n3306), .ZN(n3308) );
  AOI21_X1 U4078 ( .B1(n4402), .B2(n3308), .A(n3307), .ZN(n3310) );
  MUX2_X1 U4079 ( .A(n3878), .B(n3310), .S(n4432), .Z(n3309) );
  OAI21_X1 U4080 ( .B1(n4188), .B2(n3313), .A(n3309), .ZN(U3531) );
  INV_X1 U4081 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3311) );
  MUX2_X1 U4082 ( .A(n3311), .B(n3310), .S(n4423), .Z(n3312) );
  OAI21_X1 U4083 ( .B1(n3313), .B2(n4236), .A(n3312), .ZN(U3493) );
  NAND2_X1 U4084 ( .A1(n3315), .A2(n3314), .ZN(n3320) );
  INV_X1 U4085 ( .A(n3316), .ZN(n3318) );
  NAND2_X1 U4086 ( .A1(n3318), .A2(n2133), .ZN(n3319) );
  NAND2_X1 U4087 ( .A1(n3352), .A2(n3444), .ZN(n3323) );
  NAND2_X1 U4088 ( .A1(n3338), .A2(n3321), .ZN(n3322) );
  NAND2_X1 U4089 ( .A1(n3323), .A2(n3322), .ZN(n3324) );
  XNOR2_X1 U4090 ( .A(n3324), .B(n2903), .ZN(n3327) );
  NAND2_X1 U4091 ( .A1(n3352), .A2(n3203), .ZN(n3326) );
  NAND2_X1 U4092 ( .A1(n3444), .A2(n3338), .ZN(n3325) );
  NAND2_X1 U4093 ( .A1(n3326), .A2(n3325), .ZN(n3328) );
  NAND2_X1 U4094 ( .A1(n3327), .A2(n3328), .ZN(n3332) );
  NAND2_X1 U4095 ( .A1(n3331), .A2(n3332), .ZN(n3369) );
  INV_X1 U4096 ( .A(n3369), .ZN(n3334) );
  INV_X1 U4097 ( .A(n3327), .ZN(n3330) );
  INV_X1 U4098 ( .A(n3328), .ZN(n3329) );
  NAND2_X1 U4099 ( .A1(n3330), .A2(n3329), .ZN(n3368) );
  AOI21_X1 U4100 ( .B1(n3368), .B2(n3332), .A(n3331), .ZN(n3333) );
  AOI21_X1 U4101 ( .B1(n3334), .B2(n3368), .A(n3333), .ZN(n3342) );
  INV_X1 U4102 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3335) );
  NOR2_X1 U4103 ( .A1(STATE_REG_SCAN_IN), .A2(n3335), .ZN(n4441) );
  OAI22_X1 U4104 ( .A1(n3336), .A2(n3655), .B1(n3654), .B2(n3581), .ZN(n3337)
         );
  AOI211_X1 U4105 ( .C1(n3338), .C2(n3636), .A(n4441), .B(n3337), .ZN(n3341)
         );
  NAND2_X1 U4106 ( .A1(n3661), .A2(n3339), .ZN(n3340) );
  OAI211_X1 U4107 ( .C1(n3342), .C2(n3664), .A(n3341), .B(n3340), .ZN(U3212)
         );
  XOR2_X1 U4108 ( .A(n3716), .B(n3343), .Z(n4196) );
  XNOR2_X1 U4109 ( .A(n3344), .B(n3373), .ZN(n4193) );
  INV_X1 U4110 ( .A(n3662), .ZN(n3345) );
  OAI22_X1 U4111 ( .A1(n4263), .A2(n3346), .B1(n3345), .B2(n4352), .ZN(n3354)
         );
  OAI22_X1 U4112 ( .A1(n3653), .A2(n4101), .B1(n4134), .B2(n3657), .ZN(n3351)
         );
  INV_X1 U4113 ( .A(n3347), .ZN(n3348) );
  AOI211_X1 U4114 ( .C1(n3349), .C2(n3716), .A(n4104), .B(n3348), .ZN(n3350)
         );
  AOI211_X1 U4115 ( .C1(n4109), .C2(n3352), .A(n3351), .B(n3350), .ZN(n4195)
         );
  NOR2_X1 U4116 ( .A1(n4195), .A2(n2009), .ZN(n3353) );
  AOI211_X1 U4117 ( .C1(n4358), .C2(n4193), .A(n3354), .B(n3353), .ZN(n3355)
         );
  OAI21_X1 U4118 ( .B1(n4196), .B2(n4098), .A(n3355), .ZN(U3275) );
  NAND2_X1 U4119 ( .A1(n4077), .A2(n4076), .ZN(n3715) );
  XOR2_X1 U4120 ( .A(n3715), .B(n3356), .Z(n4185) );
  INV_X1 U4121 ( .A(n4185), .ZN(n3367) );
  XOR2_X1 U4122 ( .A(n3715), .B(n4079), .Z(n3359) );
  OAI22_X1 U4123 ( .A1(n3594), .A2(n4101), .B1(n3360), .B2(n4134), .ZN(n3357)
         );
  AOI21_X1 U4124 ( .B1(n4109), .B2(n3820), .A(n3357), .ZN(n3358) );
  OAI21_X1 U4125 ( .B1(n3359), .B2(n4104), .A(n3358), .ZN(n4184) );
  OAI21_X1 U4126 ( .B1(n3361), .B2(n3360), .A(n2046), .ZN(n4237) );
  NOR2_X1 U4127 ( .A1(n4237), .A2(n4095), .ZN(n3365) );
  INV_X1 U4128 ( .A(n3597), .ZN(n3362) );
  OAI22_X1 U4129 ( .A1(n4263), .A2(n3363), .B1(n3362), .B2(n4352), .ZN(n3364)
         );
  AOI211_X1 U4130 ( .C1(n4184), .C2(n4263), .A(n3365), .B(n3364), .ZN(n3366)
         );
  OAI21_X1 U4131 ( .B1(n3367), .B2(n4098), .A(n3366), .ZN(U3273) );
  NAND2_X1 U4132 ( .A1(n3821), .A2(n3444), .ZN(n3371) );
  NAND2_X1 U4133 ( .A1(n3373), .A2(n3321), .ZN(n3370) );
  NAND2_X1 U4134 ( .A1(n3371), .A2(n3370), .ZN(n3372) );
  XNOR2_X1 U4135 ( .A(n3372), .B(n2903), .ZN(n3383) );
  NAND2_X1 U4136 ( .A1(n3821), .A2(n3203), .ZN(n3375) );
  NAND2_X1 U4137 ( .A1(n3444), .A2(n3373), .ZN(n3374) );
  AND2_X1 U4138 ( .A1(n3375), .A2(n3374), .ZN(n3651) );
  NAND2_X1 U4139 ( .A1(n3820), .A2(n3444), .ZN(n3377) );
  NAND2_X1 U4140 ( .A1(n3583), .A2(n3435), .ZN(n3376) );
  NAND2_X1 U4141 ( .A1(n3377), .A2(n3376), .ZN(n3378) );
  XNOR2_X1 U4142 ( .A(n3378), .B(n2903), .ZN(n3382) );
  NAND2_X1 U4143 ( .A1(n3820), .A2(n3203), .ZN(n3380) );
  NAND2_X1 U4144 ( .A1(n3444), .A2(n3583), .ZN(n3379) );
  NAND2_X1 U4145 ( .A1(n3380), .A2(n3379), .ZN(n3381) );
  NOR2_X1 U4146 ( .A1(n3382), .A2(n3381), .ZN(n3384) );
  AOI21_X1 U4147 ( .B1(n3382), .B2(n3381), .A(n3384), .ZN(n3579) );
  NAND2_X1 U4148 ( .A1(n4108), .A2(n3444), .ZN(n3386) );
  NAND2_X1 U4149 ( .A1(n3596), .A2(n3321), .ZN(n3385) );
  NAND2_X1 U4150 ( .A1(n3386), .A2(n3385), .ZN(n3387) );
  XNOR2_X1 U4151 ( .A(n3387), .B(n2903), .ZN(n3391) );
  NAND2_X1 U4152 ( .A1(n4108), .A2(n3203), .ZN(n3389) );
  NAND2_X1 U4153 ( .A1(n3596), .A2(n3444), .ZN(n3388) );
  NAND2_X1 U4154 ( .A1(n3389), .A2(n3388), .ZN(n3390) );
  NAND2_X1 U4155 ( .A1(n3391), .A2(n3390), .ZN(n3589) );
  NOR2_X1 U4156 ( .A1(n3391), .A2(n3390), .ZN(n3588) );
  AOI21_X2 U4157 ( .B1(n3592), .B2(n3589), .A(n3588), .ZN(n3633) );
  NAND2_X1 U4158 ( .A1(n4087), .A2(n3458), .ZN(n3393) );
  NAND2_X1 U4159 ( .A1(n4113), .A2(n3321), .ZN(n3392) );
  NAND2_X1 U4160 ( .A1(n3393), .A2(n3392), .ZN(n3394) );
  XNOR2_X1 U4161 ( .A(n3394), .B(n3451), .ZN(n3631) );
  NAND2_X1 U4162 ( .A1(n4087), .A2(n3459), .ZN(n3396) );
  NAND2_X1 U4163 ( .A1(n3458), .A2(n4113), .ZN(n3395) );
  NAND2_X1 U4164 ( .A1(n4063), .A2(n3444), .ZN(n3398) );
  NAND2_X1 U4165 ( .A1(n3400), .A2(n3321), .ZN(n3397) );
  NAND2_X1 U4166 ( .A1(n3398), .A2(n3397), .ZN(n3399) );
  XNOR2_X1 U4167 ( .A(n3399), .B(n2903), .ZN(n3403) );
  NAND2_X1 U4168 ( .A1(n4063), .A2(n3203), .ZN(n3402) );
  NAND2_X1 U4169 ( .A1(n3444), .A2(n3400), .ZN(n3401) );
  NAND2_X1 U4170 ( .A1(n3402), .A2(n3401), .ZN(n3404) );
  NAND2_X1 U4171 ( .A1(n3403), .A2(n3404), .ZN(n3533) );
  OAI21_X1 U4172 ( .B1(n3631), .B2(n3534), .A(n3533), .ZN(n3409) );
  NAND3_X1 U4173 ( .A1(n3533), .A2(n3534), .A3(n3631), .ZN(n3407) );
  INV_X1 U4174 ( .A(n3403), .ZN(n3406) );
  INV_X1 U4175 ( .A(n3404), .ZN(n3405) );
  NAND2_X1 U4176 ( .A1(n3406), .A2(n3405), .ZN(n3532) );
  NAND2_X1 U4177 ( .A1(n4042), .A2(n3444), .ZN(n3412) );
  OR2_X1 U4178 ( .A1(n3410), .A2(n4067), .ZN(n3411) );
  NAND2_X1 U4179 ( .A1(n3412), .A2(n3411), .ZN(n3413) );
  XNOR2_X1 U4180 ( .A(n3413), .B(n3451), .ZN(n3416) );
  INV_X1 U4181 ( .A(n3458), .ZN(n3453) );
  NOR2_X1 U4182 ( .A1(n3453), .A2(n4067), .ZN(n3414) );
  AOI21_X1 U4183 ( .B1(n4042), .B2(n3459), .A(n3414), .ZN(n3415) );
  OR2_X1 U4184 ( .A1(n3416), .A2(n3415), .ZN(n3613) );
  NAND2_X1 U4185 ( .A1(n3416), .A2(n3415), .ZN(n3615) );
  NAND2_X1 U4186 ( .A1(n4027), .A2(n3444), .ZN(n3418) );
  OR2_X1 U4187 ( .A1(n3410), .A2(n4039), .ZN(n3417) );
  NAND2_X1 U4188 ( .A1(n3418), .A2(n3417), .ZN(n3419) );
  XNOR2_X1 U4189 ( .A(n3419), .B(n3451), .ZN(n3422) );
  NOR2_X1 U4190 ( .A1(n3453), .A2(n4039), .ZN(n3420) );
  AOI21_X1 U4191 ( .B1(n4027), .B2(n3459), .A(n3420), .ZN(n3421) );
  AND2_X1 U4192 ( .A1(n3422), .A2(n3421), .ZN(n3552) );
  OR2_X1 U4193 ( .A1(n3422), .A2(n3421), .ZN(n3553) );
  OAI22_X1 U4194 ( .A1(n4040), .A2(n3453), .B1(n3410), .B2(n4030), .ZN(n3423)
         );
  XNOR2_X1 U4195 ( .A(n3423), .B(n2903), .ZN(n3426) );
  OAI22_X1 U4196 ( .A1(n4040), .A2(n3424), .B1(n3453), .B2(n4030), .ZN(n3425)
         );
  XNOR2_X1 U4197 ( .A(n3426), .B(n3425), .ZN(n3623) );
  NOR2_X1 U4198 ( .A1(n3426), .A2(n3425), .ZN(n3524) );
  NAND2_X1 U4199 ( .A1(n4026), .A2(n3444), .ZN(n3428) );
  OR2_X1 U4200 ( .A1(n3410), .A2(n3527), .ZN(n3427) );
  NAND2_X1 U4201 ( .A1(n3428), .A2(n3427), .ZN(n3429) );
  XNOR2_X1 U4202 ( .A(n3429), .B(n3451), .ZN(n3432) );
  NOR2_X1 U4203 ( .A1(n3453), .A2(n3527), .ZN(n3430) );
  AOI21_X1 U4204 ( .B1(n4026), .B2(n3459), .A(n3430), .ZN(n3431) );
  XNOR2_X1 U4205 ( .A(n3432), .B(n3431), .ZN(n3523) );
  NOR2_X1 U4206 ( .A1(n3432), .A2(n3431), .ZN(n3438) );
  NAND2_X1 U4207 ( .A1(n4001), .A2(n3459), .ZN(n3434) );
  NAND2_X1 U4208 ( .A1(n3444), .A2(n3981), .ZN(n3433) );
  NAND2_X1 U4209 ( .A1(n3434), .A2(n3433), .ZN(n3437) );
  AOI22_X1 U4210 ( .A1(n4001), .A2(n3444), .B1(n3435), .B2(n3981), .ZN(n3436)
         );
  XNOR2_X1 U4211 ( .A(n3436), .B(n2903), .ZN(n3604) );
  NOR2_X1 U4212 ( .A1(n3410), .A2(n3572), .ZN(n3439) );
  AOI21_X1 U4213 ( .B1(n3944), .B2(n3444), .A(n3439), .ZN(n3440) );
  XNOR2_X1 U4214 ( .A(n3440), .B(n2903), .ZN(n3443) );
  NOR2_X1 U4215 ( .A1(n3453), .A2(n3572), .ZN(n3441) );
  AOI21_X1 U4216 ( .B1(n3944), .B2(n3459), .A(n3441), .ZN(n3442) );
  NAND2_X1 U4217 ( .A1(n3443), .A2(n3442), .ZN(n3567) );
  NOR2_X1 U4218 ( .A1(n3443), .A2(n3442), .ZN(n3568) );
  NAND2_X1 U4219 ( .A1(n3481), .A2(n3444), .ZN(n3446) );
  OR2_X1 U4220 ( .A1(n3410), .A2(n3950), .ZN(n3445) );
  NAND2_X1 U4221 ( .A1(n3446), .A2(n3445), .ZN(n3447) );
  XNOR2_X1 U4222 ( .A(n3447), .B(n3451), .ZN(n3450) );
  NOR2_X1 U4223 ( .A1(n3453), .A2(n3950), .ZN(n3448) );
  AOI21_X1 U4224 ( .B1(n3481), .B2(n3459), .A(n3448), .ZN(n3449) );
  OR2_X1 U4225 ( .A1(n3450), .A2(n3449), .ZN(n3640) );
  OAI22_X1 U4226 ( .A1(n3644), .A2(n3453), .B1(n3515), .B2(n3410), .ZN(n3452)
         );
  XNOR2_X1 U4227 ( .A(n3452), .B(n3451), .ZN(n3454) );
  OAI22_X1 U4228 ( .A1(n3644), .A2(n3424), .B1(n3515), .B2(n3453), .ZN(n3456)
         );
  XNOR2_X1 U4229 ( .A(n3454), .B(n3456), .ZN(n3513) );
  INV_X1 U4230 ( .A(n3454), .ZN(n3455) );
  INV_X1 U4231 ( .A(n3465), .ZN(n3926) );
  AOI22_X1 U4232 ( .A1(n3927), .A2(n3444), .B1(n3321), .B2(n3926), .ZN(n3457)
         );
  XNOR2_X1 U4233 ( .A(n3457), .B(n2903), .ZN(n3461) );
  AOI22_X1 U4234 ( .A1(n3927), .A2(n3459), .B1(n3458), .B2(n3926), .ZN(n3460)
         );
  XNOR2_X1 U4235 ( .A(n3461), .B(n3460), .ZN(n3462) );
  XNOR2_X1 U4236 ( .A(n3463), .B(n3462), .ZN(n3469) );
  OAI22_X1 U4237 ( .A1(n3658), .A2(n3465), .B1(STATE_REG_SCAN_IN), .B2(n3464), 
        .ZN(n3467) );
  OAI22_X1 U4238 ( .A1(n3699), .A2(n3654), .B1(n3644), .B2(n3655), .ZN(n3466)
         );
  AOI211_X1 U4239 ( .C1(n3506), .C2(n3661), .A(n3467), .B(n3466), .ZN(n3468)
         );
  OAI21_X1 U4240 ( .B1(n3469), .B2(n3664), .A(n3468), .ZN(U3217) );
  XNOR2_X1 U4241 ( .A(n3470), .B(n3478), .ZN(n4147) );
  INV_X1 U4242 ( .A(n3471), .ZN(n3949) );
  AOI21_X1 U4243 ( .B1(n3480), .B2(n3949), .A(n3472), .ZN(n4145) );
  INV_X1 U4244 ( .A(n3519), .ZN(n3474) );
  OAI22_X1 U4245 ( .A1(n3474), .A2(n4352), .B1(n3473), .B2(n4263), .ZN(n3475)
         );
  AOI21_X1 U4246 ( .B1(n4145), .B2(n4358), .A(n3475), .ZN(n3485) );
  INV_X1 U4247 ( .A(n3927), .ZN(n3516) );
  OAI21_X1 U4248 ( .B1(n3478), .B2(n3477), .A(n3476), .ZN(n3479) );
  NAND2_X1 U4249 ( .A1(n3479), .A2(n4032), .ZN(n3483) );
  AOI22_X1 U4250 ( .A1(n3481), .A2(n4109), .B1(n3480), .B2(n4127), .ZN(n3482)
         );
  OAI211_X1 U4251 ( .C1(n3516), .C2(n4101), .A(n3483), .B(n3482), .ZN(n4144)
         );
  NAND2_X1 U4252 ( .A1(n4144), .A2(n4263), .ZN(n3484) );
  OAI211_X1 U4253 ( .C1(n4147), .C2(n4098), .A(n3485), .B(n3484), .ZN(U3263)
         );
  NAND2_X1 U4254 ( .A1(n3487), .A2(n2017), .ZN(n3488) );
  NAND2_X1 U4255 ( .A1(n3486), .A2(n3488), .ZN(n4398) );
  XNOR2_X1 U4256 ( .A(n2017), .B(n3489), .ZN(n3494) );
  AOI22_X1 U4257 ( .A1(n3831), .A2(n4109), .B1(n3490), .B2(n4127), .ZN(n3492)
         );
  NAND2_X1 U4258 ( .A1(n3829), .A2(n4025), .ZN(n3491) );
  OAI211_X1 U4259 ( .C1(n4398), .C2(n4065), .A(n3492), .B(n3491), .ZN(n3493)
         );
  AOI21_X1 U4260 ( .B1(n3494), .B2(n4032), .A(n3493), .ZN(n3495) );
  INV_X1 U4261 ( .A(n3495), .ZN(n4400) );
  INV_X1 U4262 ( .A(n3496), .ZN(n3499) );
  OAI211_X1 U4263 ( .C1(n3499), .C2(n3498), .A(n4421), .B(n3497), .ZN(n4399)
         );
  OAI22_X1 U4264 ( .A1(n4399), .A2(n4247), .B1(n4352), .B2(n3500), .ZN(n3501)
         );
  OAI21_X1 U4265 ( .B1(n4400), .B2(n3501), .A(n4263), .ZN(n3503) );
  NAND2_X1 U4266 ( .A1(n2009), .A2(REG2_REG_4__SCAN_IN), .ZN(n3502) );
  OAI211_X1 U4267 ( .C1(n4398), .C2(n3504), .A(n3503), .B(n3502), .ZN(U3286)
         );
  INV_X1 U4268 ( .A(n3505), .ZN(n3510) );
  AOI22_X1 U4269 ( .A1(n3506), .A2(n4367), .B1(REG2_REG_28__SCAN_IN), .B2(
        n2009), .ZN(n3507) );
  OAI21_X1 U4270 ( .B1(n3508), .B2(n4095), .A(n3507), .ZN(n3509) );
  AOI21_X1 U4271 ( .B1(n3510), .B2(n4263), .A(n3509), .ZN(n3511) );
  OAI21_X1 U4272 ( .B1(n3512), .B2(n4098), .A(n3511), .ZN(U3262) );
  XNOR2_X1 U4273 ( .A(n3514), .B(n3513), .ZN(n3521) );
  INV_X1 U4274 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4496) );
  OAI22_X1 U4275 ( .A1(n3658), .A2(n3515), .B1(STATE_REG_SCAN_IN), .B2(n4496), 
        .ZN(n3518) );
  OAI22_X1 U4276 ( .A1(n3516), .A2(n3654), .B1(n3966), .B2(n3655), .ZN(n3517)
         );
  AOI211_X1 U4277 ( .C1(n3519), .C2(n3661), .A(n3518), .B(n3517), .ZN(n3520)
         );
  OAI21_X1 U4278 ( .B1(n3521), .B2(n3664), .A(n3520), .ZN(U3211) );
  OAI21_X1 U4279 ( .B1(n2019), .B2(n3524), .A(n3523), .ZN(n3525) );
  NAND3_X1 U4280 ( .A1(n2146), .A2(n3557), .A3(n3525), .ZN(n3531) );
  INV_X1 U4281 ( .A(n4001), .ZN(n3573) );
  OAI22_X1 U4282 ( .A1(n3573), .A2(n3654), .B1(n3655), .B2(n4040), .ZN(n3529)
         );
  OAI22_X1 U4283 ( .A1(n3658), .A2(n3527), .B1(STATE_REG_SCAN_IN), .B2(n3526), 
        .ZN(n3528) );
  AOI211_X1 U4284 ( .C1(n4009), .C2(n3661), .A(n3529), .B(n3528), .ZN(n3530)
         );
  NAND2_X1 U4285 ( .A1(n3531), .A2(n3530), .ZN(U3213) );
  NAND2_X1 U4286 ( .A1(n3533), .A2(n3532), .ZN(n3538) );
  INV_X1 U4287 ( .A(n3534), .ZN(n3630) );
  NOR2_X1 U4288 ( .A1(n3633), .A2(n3630), .ZN(n3536) );
  INV_X1 U4289 ( .A(n3633), .ZN(n3535) );
  OAI22_X1 U4290 ( .A1(n3536), .A2(n3631), .B1(n3535), .B2(n3534), .ZN(n3537)
         );
  XOR2_X1 U4291 ( .A(n3538), .B(n3537), .Z(n3542) );
  AOI22_X1 U4292 ( .A1(n3561), .A2(n4087), .B1(n3560), .B2(n4042), .ZN(n3539)
         );
  NAND2_X1 U4293 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3907) );
  OAI211_X1 U4294 ( .C1(n3658), .C2(n4090), .A(n3539), .B(n3907), .ZN(n3540)
         );
  AOI21_X1 U4295 ( .B1(n4093), .B2(n3661), .A(n3540), .ZN(n3541) );
  OAI21_X1 U4296 ( .B1(n3542), .B2(n3664), .A(n3541), .ZN(U3216) );
  AOI22_X1 U4297 ( .A1(n3636), .A2(n3544), .B1(n3561), .B2(n3543), .ZN(n3551)
         );
  OAI211_X1 U4298 ( .C1(n3547), .C2(n3546), .A(n3545), .B(n3557), .ZN(n3550)
         );
  AOI22_X1 U4299 ( .A1(n3548), .A2(REG3_REG_1__SCAN_IN), .B1(n3560), .B2(n3832), .ZN(n3549) );
  NAND3_X1 U4300 ( .A1(n3551), .A2(n3550), .A3(n3549), .ZN(U3219) );
  INV_X1 U4301 ( .A(n3552), .ZN(n3554) );
  NAND2_X1 U4302 ( .A1(n3554), .A2(n3553), .ZN(n3558) );
  OAI211_X1 U4303 ( .C1(n3555), .C2(n2154), .A(n3613), .B(n3558), .ZN(n3556)
         );
  OAI211_X1 U4304 ( .C1(n3559), .C2(n3558), .A(n3557), .B(n3556), .ZN(n3565)
         );
  AOI22_X1 U4305 ( .A1(n3636), .A2(n4045), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3564) );
  AOI22_X1 U4306 ( .A1(n3561), .A2(n4042), .B1(n3560), .B2(n4002), .ZN(n3563)
         );
  NAND2_X1 U4307 ( .A1(n3661), .A2(n4048), .ZN(n3562) );
  NAND4_X1 U4308 ( .A1(n3565), .A2(n3564), .A3(n3563), .A4(n3562), .ZN(U3220)
         );
  NOR2_X1 U4309 ( .A1(n3568), .A2(n2111), .ZN(n3569) );
  XNOR2_X1 U4310 ( .A(n3566), .B(n3569), .ZN(n3577) );
  INV_X1 U4311 ( .A(n3570), .ZN(n3969) );
  OAI22_X1 U4312 ( .A1(n3658), .A2(n3572), .B1(STATE_REG_SCAN_IN), .B2(n3571), 
        .ZN(n3575) );
  OAI22_X1 U4313 ( .A1(n3966), .A2(n3654), .B1(n3573), .B2(n3655), .ZN(n3574)
         );
  AOI211_X1 U4314 ( .C1(n3969), .C2(n3661), .A(n3575), .B(n3574), .ZN(n3576)
         );
  OAI21_X1 U4315 ( .B1(n3577), .B2(n3664), .A(n3576), .ZN(U3222) );
  AOI21_X1 U4316 ( .B1(n3651), .B2(n3649), .A(n3578), .ZN(n3580) );
  XNOR2_X1 U4317 ( .A(n3580), .B(n3579), .ZN(n3587) );
  NOR2_X1 U4318 ( .A1(STATE_REG_SCAN_IN), .A2(n2412), .ZN(n4319) );
  OAI22_X1 U4319 ( .A1(n3581), .A2(n3655), .B1(n3654), .B2(n3634), .ZN(n3582)
         );
  AOI211_X1 U4320 ( .C1(n3583), .C2(n3636), .A(n4319), .B(n3582), .ZN(n3586)
         );
  NAND2_X1 U4321 ( .A1(n3661), .A2(n3584), .ZN(n3585) );
  OAI211_X1 U4322 ( .C1(n3587), .C2(n3664), .A(n3586), .B(n3585), .ZN(U3223)
         );
  INV_X1 U4323 ( .A(n3588), .ZN(n3590) );
  NAND2_X1 U4324 ( .A1(n3590), .A2(n3589), .ZN(n3591) );
  XNOR2_X1 U4325 ( .A(n3592), .B(n3591), .ZN(n3600) );
  NOR2_X1 U4326 ( .A1(STATE_REG_SCAN_IN), .A2(n3593), .ZN(n4329) );
  OAI22_X1 U4327 ( .A1(n3594), .A2(n3654), .B1(n3655), .B2(n3653), .ZN(n3595)
         );
  AOI211_X1 U4328 ( .C1(n3596), .C2(n3636), .A(n4329), .B(n3595), .ZN(n3599)
         );
  NAND2_X1 U4329 ( .A1(n3661), .A2(n3597), .ZN(n3598) );
  OAI211_X1 U4330 ( .C1(n3600), .C2(n3664), .A(n3599), .B(n3598), .ZN(U3225)
         );
  INV_X1 U4331 ( .A(n3601), .ZN(n3603) );
  NAND2_X1 U4332 ( .A1(n3603), .A2(n3602), .ZN(n3605) );
  XNOR2_X1 U4333 ( .A(n3605), .B(n3604), .ZN(n3611) );
  INV_X1 U4334 ( .A(n3987), .ZN(n3609) );
  OAI22_X1 U4335 ( .A1(n3984), .A2(n3654), .B1(n3655), .B2(n3624), .ZN(n3608)
         );
  INV_X1 U4336 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3606) );
  OAI22_X1 U4337 ( .A1(n3658), .A2(n3986), .B1(STATE_REG_SCAN_IN), .B2(n3606), 
        .ZN(n3607) );
  AOI211_X1 U4338 ( .C1(n3609), .C2(n3661), .A(n3608), .B(n3607), .ZN(n3610)
         );
  OAI21_X1 U4339 ( .B1(n3611), .B2(n3664), .A(n3610), .ZN(U3226) );
  INV_X1 U4340 ( .A(n3612), .ZN(n3616) );
  AOI21_X1 U4341 ( .B1(n3613), .B2(n3615), .A(n3555), .ZN(n3614) );
  AOI21_X1 U4342 ( .B1(n3616), .B2(n3615), .A(n3614), .ZN(n3621) );
  OAI22_X1 U4343 ( .A1(n4102), .A2(n3655), .B1(n3654), .B2(n4055), .ZN(n3619)
         );
  OAI22_X1 U4344 ( .A1(n3658), .A2(n4067), .B1(STATE_REG_SCAN_IN), .B2(n3617), 
        .ZN(n3618) );
  AOI211_X1 U4345 ( .C1(n4070), .C2(n3661), .A(n3619), .B(n3618), .ZN(n3620)
         );
  OAI21_X1 U4346 ( .B1(n3621), .B2(n3664), .A(n3620), .ZN(U3230) );
  AOI21_X1 U4347 ( .B1(n3623), .B2(n3622), .A(n2019), .ZN(n3629) );
  OAI22_X1 U4348 ( .A1(n3624), .A2(n3654), .B1(n3655), .B2(n4055), .ZN(n3626)
         );
  OAI22_X1 U4349 ( .A1(n3658), .A2(n4030), .B1(STATE_REG_SCAN_IN), .B2(n4485), 
        .ZN(n3625) );
  AOI211_X1 U4350 ( .C1(n3627), .C2(n3661), .A(n3626), .B(n3625), .ZN(n3628)
         );
  OAI21_X1 U4351 ( .B1(n3629), .B2(n3664), .A(n3628), .ZN(U3232) );
  XNOR2_X1 U4352 ( .A(n3631), .B(n3630), .ZN(n3632) );
  XNOR2_X1 U4353 ( .A(n3633), .B(n3632), .ZN(n3639) );
  INV_X1 U4354 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4482) );
  NOR2_X1 U4355 ( .A1(STATE_REG_SCAN_IN), .A2(n4482), .ZN(n4343) );
  OAI22_X1 U4356 ( .A1(n4102), .A2(n3654), .B1(n3655), .B2(n3634), .ZN(n3635)
         );
  AOI211_X1 U4357 ( .C1(n4113), .C2(n3636), .A(n4343), .B(n3635), .ZN(n3638)
         );
  NAND2_X1 U4358 ( .A1(n3661), .A2(n4117), .ZN(n3637) );
  OAI211_X1 U4359 ( .C1(n3639), .C2(n3664), .A(n3638), .B(n3637), .ZN(U3235)
         );
  NAND2_X1 U4360 ( .A1(n2032), .A2(n3640), .ZN(n3641) );
  XNOR2_X1 U4361 ( .A(n3642), .B(n3641), .ZN(n3648) );
  INV_X1 U4362 ( .A(n3643), .ZN(n3952) );
  OAI22_X1 U4363 ( .A1(n3658), .A2(n3950), .B1(STATE_REG_SCAN_IN), .B2(n4479), 
        .ZN(n3646) );
  OAI22_X1 U4364 ( .A1(n3644), .A2(n3654), .B1(n3984), .B2(n3655), .ZN(n3645)
         );
  AOI211_X1 U4365 ( .C1(n3952), .C2(n3661), .A(n3646), .B(n3645), .ZN(n3647)
         );
  OAI21_X1 U4366 ( .B1(n3648), .B2(n3664), .A(n3647), .ZN(U3237) );
  INV_X1 U4367 ( .A(n3578), .ZN(n3650) );
  NAND2_X1 U4368 ( .A1(n3650), .A2(n3649), .ZN(n3652) );
  XNOR2_X1 U4369 ( .A(n3652), .B(n3651), .ZN(n3665) );
  OAI22_X1 U4370 ( .A1(n2399), .A2(n3655), .B1(n3654), .B2(n3653), .ZN(n3660)
         );
  OAI22_X1 U4371 ( .A1(n3658), .A2(n3657), .B1(STATE_REG_SCAN_IN), .B2(n3656), 
        .ZN(n3659) );
  AOI211_X1 U4372 ( .C1(n3662), .C2(n3661), .A(n3660), .B(n3659), .ZN(n3663)
         );
  OAI21_X1 U4373 ( .B1(n3665), .B2(n3664), .A(n3663), .ZN(U3238) );
  INV_X1 U4374 ( .A(REG2_REG_30__SCAN_IN), .ZN(n3669) );
  NAND2_X1 U4375 ( .A1(n2013), .A2(REG1_REG_30__SCAN_IN), .ZN(n3668) );
  NAND2_X1 U4376 ( .A1(n3666), .A2(REG0_REG_30__SCAN_IN), .ZN(n3667) );
  OAI211_X1 U4377 ( .C1(n3670), .C2(n3669), .A(n3668), .B(n3667), .ZN(n3919)
         );
  NAND2_X1 U4378 ( .A1(n2265), .A2(DATAI_30_), .ZN(n4135) );
  NAND2_X1 U4379 ( .A1(n3919), .A2(n4135), .ZN(n3704) );
  AND2_X1 U4380 ( .A1(n3704), .A2(n4123), .ZN(n3698) );
  NAND2_X1 U4381 ( .A1(n2265), .A2(DATAI_31_), .ZN(n4125) );
  INV_X1 U4382 ( .A(n3699), .ZN(n3671) );
  NAND2_X1 U4383 ( .A1(n2265), .A2(DATAI_29_), .ZN(n3700) );
  NAND2_X1 U4384 ( .A1(n3671), .A2(n3700), .ZN(n3672) );
  NAND2_X1 U4385 ( .A1(n3672), .A2(n3915), .ZN(n3801) );
  NOR3_X1 U4386 ( .A1(n3673), .A2(n3728), .A3(n3801), .ZN(n3695) );
  NAND2_X1 U4387 ( .A1(n3913), .A2(n3674), .ZN(n3694) );
  INV_X1 U4388 ( .A(n3694), .ZN(n3676) );
  NAND2_X1 U4389 ( .A1(n4123), .A2(n4125), .ZN(n3805) );
  OR2_X1 U4390 ( .A1(n3919), .A2(n4135), .ZN(n3675) );
  AND2_X1 U4391 ( .A1(n3805), .A2(n3675), .ZN(n3732) );
  INV_X1 U4392 ( .A(n3700), .ZN(n3934) );
  NAND2_X1 U4393 ( .A1(n3699), .A2(n3934), .ZN(n3692) );
  OAI211_X1 U4394 ( .C1(n3676), .C2(n3801), .A(n3732), .B(n3692), .ZN(n3809)
         );
  NAND2_X1 U4395 ( .A1(n3677), .A2(n3681), .ZN(n3777) );
  NAND2_X1 U4396 ( .A1(n3679), .A2(n3678), .ZN(n3680) );
  NAND2_X1 U4397 ( .A1(n3681), .A2(n3680), .ZN(n3783) );
  OAI21_X1 U4398 ( .B1(n3682), .B2(n3777), .A(n3783), .ZN(n3684) );
  AOI211_X1 U4399 ( .C1(n3684), .C2(n3788), .A(n2081), .B(n3787), .ZN(n3686)
         );
  INV_X1 U4400 ( .A(n3685), .ZN(n3792) );
  OAI21_X1 U4401 ( .B1(n3686), .B2(n3792), .A(n3790), .ZN(n3688) );
  AOI21_X1 U4402 ( .B1(n3795), .B2(n3688), .A(n3687), .ZN(n3690) );
  OAI21_X1 U4403 ( .B1(n3690), .B2(n3798), .A(n3689), .ZN(n3691) );
  NAND4_X1 U4404 ( .A1(n3796), .A2(n3732), .A3(n3692), .A4(n3691), .ZN(n3693)
         );
  OAI22_X1 U4405 ( .A1(n3695), .A2(n3809), .B1(n3694), .B2(n3693), .ZN(n3696)
         );
  OAI21_X1 U4406 ( .B1(n4123), .B2(n4135), .A(n3696), .ZN(n3697) );
  OAI21_X1 U4407 ( .B1(n3698), .B2(n4125), .A(n3697), .ZN(n3740) );
  XOR2_X1 U4408 ( .A(n3700), .B(n3699), .Z(n3930) );
  NAND2_X1 U4409 ( .A1(n3939), .A2(n3701), .ZN(n3961) );
  NAND2_X1 U4410 ( .A1(n3702), .A2(n3959), .ZN(n3978) );
  OR2_X1 U4411 ( .A1(n4123), .A2(n4125), .ZN(n3703) );
  NAND2_X1 U4412 ( .A1(n3704), .A2(n3703), .ZN(n3806) );
  NOR3_X1 U4413 ( .A1(n3961), .A2(n3978), .A3(n3806), .ZN(n3710) );
  NAND2_X1 U4414 ( .A1(n3975), .A2(n3705), .ZN(n3999) );
  NOR2_X1 U4415 ( .A1(n3999), .A2(n3706), .ZN(n3709) );
  NAND4_X1 U4416 ( .A1(n3710), .A2(n3709), .A3(n3708), .A4(n3707), .ZN(n3727)
         );
  NOR4_X1 U4417 ( .A1(n3713), .A2(n3712), .A3(n4111), .A4(n3711), .ZN(n3725)
         );
  INV_X1 U4418 ( .A(n3714), .ZN(n3717) );
  OR2_X1 U4419 ( .A1(n3994), .A2(n3995), .ZN(n4038) );
  NOR4_X1 U4420 ( .A1(n3717), .A2(n3716), .A3(n4038), .A4(n3715), .ZN(n3724)
         );
  NOR4_X1 U4421 ( .A1(n4015), .A2(n3719), .A3(n2553), .A4(n3718), .ZN(n3723)
         );
  AND4_X1 U4422 ( .A1(n3721), .A2(n2017), .A3(n3720), .A4(n3757), .ZN(n3722)
         );
  NAND4_X1 U4423 ( .A1(n3725), .A2(n3724), .A3(n3723), .A4(n3722), .ZN(n3726)
         );
  NOR4_X1 U4424 ( .A1(n3930), .A2(n3728), .A3(n3727), .A4(n3726), .ZN(n3738)
         );
  NAND2_X1 U4425 ( .A1(n3730), .A2(n3729), .ZN(n3941) );
  INV_X1 U4426 ( .A(n3941), .ZN(n3734) );
  XNOR2_X1 U4427 ( .A(n4042), .B(n3731), .ZN(n4059) );
  NAND4_X1 U4428 ( .A1(n3734), .A2(n4059), .A3(n3733), .A4(n3732), .ZN(n3736)
         );
  XNOR2_X1 U4429 ( .A(n4063), .B(n4090), .ZN(n4084) );
  NOR4_X1 U4430 ( .A1(n3736), .A2(n3924), .A3(n4084), .A4(n3735), .ZN(n3737)
         );
  NAND2_X1 U4431 ( .A1(n3738), .A2(n3737), .ZN(n3739) );
  MUX2_X1 U4432 ( .A(n3740), .B(n3739), .S(n2583), .Z(n3812) );
  INV_X1 U4433 ( .A(n3741), .ZN(n3744) );
  OAI211_X1 U4434 ( .C1(n3744), .C2(n2551), .A(n3743), .B(n3742), .ZN(n3746)
         );
  NAND3_X1 U4435 ( .A1(n3749), .A2(n3748), .A3(n3747), .ZN(n3752) );
  NAND3_X1 U4436 ( .A1(n3752), .A2(n3751), .A3(n3750), .ZN(n3755) );
  NAND4_X1 U4437 ( .A1(n3755), .A2(n3754), .A3(n3753), .A4(n3761), .ZN(n3758)
         );
  NAND3_X1 U4438 ( .A1(n3758), .A2(n3757), .A3(n3756), .ZN(n3770) );
  NAND2_X1 U4439 ( .A1(n3760), .A2(n3759), .ZN(n3763) );
  INV_X1 U4440 ( .A(n3763), .ZN(n3769) );
  INV_X1 U4441 ( .A(n3761), .ZN(n3764) );
  NOR3_X1 U4442 ( .A1(n3764), .A2(n3763), .A3(n3762), .ZN(n3768) );
  NAND2_X1 U4443 ( .A1(n3766), .A2(n3765), .ZN(n3767) );
  AOI211_X1 U4444 ( .C1(n3770), .C2(n3769), .A(n3768), .B(n3767), .ZN(n3773)
         );
  OAI21_X1 U4445 ( .B1(n3773), .B2(n3772), .A(n3771), .ZN(n3785) );
  AND4_X1 U4446 ( .A1(n3783), .A2(n3776), .A3(n3775), .A4(n3774), .ZN(n3784)
         );
  INV_X1 U4447 ( .A(n3776), .ZN(n3780) );
  INV_X1 U4448 ( .A(n3777), .ZN(n3778) );
  OAI211_X1 U4449 ( .C1(n3781), .C2(n3780), .A(n3779), .B(n3778), .ZN(n3782)
         );
  AOI22_X1 U4450 ( .A1(n3785), .A2(n3784), .B1(n3783), .B2(n3782), .ZN(n3786)
         );
  OR2_X1 U4451 ( .A1(n3786), .A2(n2081), .ZN(n3789) );
  AOI21_X1 U4452 ( .B1(n3789), .B2(n3788), .A(n3787), .ZN(n3793) );
  INV_X1 U4453 ( .A(n3994), .ZN(n3791) );
  OAI211_X1 U4454 ( .C1(n3793), .C2(n3792), .A(n3791), .B(n3790), .ZN(n3794)
         );
  NAND2_X1 U4455 ( .A1(n3795), .A2(n3794), .ZN(n3799) );
  INV_X1 U4456 ( .A(n3796), .ZN(n3797) );
  AOI211_X1 U4457 ( .C1(n3800), .C2(n3799), .A(n3798), .B(n3797), .ZN(n3803)
         );
  NOR4_X1 U4458 ( .A1(n3804), .A2(n3803), .A3(n3802), .A4(n3801), .ZN(n3810)
         );
  INV_X1 U4459 ( .A(n3805), .ZN(n3808) );
  INV_X1 U4460 ( .A(n3806), .ZN(n3807) );
  OAI22_X1 U4461 ( .A1(n3810), .A2(n3809), .B1(n3808), .B2(n3807), .ZN(n3811)
         );
  MUX2_X1 U4462 ( .A(n3812), .B(n3811), .S(n2542), .Z(n3813) );
  XNOR2_X1 U4463 ( .A(n3813), .B(n3908), .ZN(n3819) );
  NOR2_X1 U4464 ( .A1(n3815), .A2(n3814), .ZN(n3817) );
  OAI21_X1 U4465 ( .B1(n3818), .B2(n4245), .A(B_REG_SCAN_IN), .ZN(n3816) );
  OAI22_X1 U4466 ( .A1(n3819), .A2(n3818), .B1(n3817), .B2(n3816), .ZN(U3239)
         );
  MUX2_X1 U4467 ( .A(DATAO_REG_30__SCAN_IN), .B(n3919), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4468 ( .A(n3927), .B(DATAO_REG_28__SCAN_IN), .S(n3833), .Z(U3578)
         );
  MUX2_X1 U4469 ( .A(n3945), .B(DATAO_REG_27__SCAN_IN), .S(n3833), .Z(U3577)
         );
  MUX2_X1 U4470 ( .A(n3944), .B(DATAO_REG_25__SCAN_IN), .S(n3833), .Z(U3575)
         );
  MUX2_X1 U4471 ( .A(n4001), .B(DATAO_REG_24__SCAN_IN), .S(n3833), .Z(U3574)
         );
  MUX2_X1 U4472 ( .A(n4026), .B(DATAO_REG_23__SCAN_IN), .S(n3833), .Z(U3573)
         );
  MUX2_X1 U4473 ( .A(n4027), .B(DATAO_REG_21__SCAN_IN), .S(n3833), .Z(U3571)
         );
  MUX2_X1 U4474 ( .A(n4042), .B(DATAO_REG_20__SCAN_IN), .S(n3833), .Z(U3570)
         );
  MUX2_X1 U4475 ( .A(n4063), .B(DATAO_REG_19__SCAN_IN), .S(n3833), .Z(U3569)
         );
  MUX2_X1 U4476 ( .A(n4087), .B(DATAO_REG_18__SCAN_IN), .S(n3833), .Z(U3568)
         );
  MUX2_X1 U4477 ( .A(n4108), .B(DATAO_REG_17__SCAN_IN), .S(n3833), .Z(U3567)
         );
  MUX2_X1 U4478 ( .A(n3820), .B(DATAO_REG_16__SCAN_IN), .S(n3833), .Z(U3566)
         );
  MUX2_X1 U4479 ( .A(n3821), .B(DATAO_REG_15__SCAN_IN), .S(n3833), .Z(U3565)
         );
  MUX2_X1 U4480 ( .A(n3822), .B(DATAO_REG_13__SCAN_IN), .S(n3833), .Z(U3563)
         );
  MUX2_X1 U4481 ( .A(n3823), .B(DATAO_REG_12__SCAN_IN), .S(n3833), .Z(U3562)
         );
  MUX2_X1 U4482 ( .A(n3824), .B(DATAO_REG_11__SCAN_IN), .S(n3833), .Z(U3561)
         );
  MUX2_X1 U4483 ( .A(n3825), .B(DATAO_REG_10__SCAN_IN), .S(n3833), .Z(U3560)
         );
  MUX2_X1 U4484 ( .A(n3826), .B(DATAO_REG_9__SCAN_IN), .S(n3833), .Z(U3559) );
  MUX2_X1 U4485 ( .A(n3827), .B(DATAO_REG_8__SCAN_IN), .S(n3833), .Z(U3558) );
  MUX2_X1 U4486 ( .A(n3828), .B(DATAO_REG_6__SCAN_IN), .S(n3833), .Z(U3556) );
  MUX2_X1 U4487 ( .A(n3829), .B(DATAO_REG_5__SCAN_IN), .S(n3833), .Z(U3555) );
  MUX2_X1 U4488 ( .A(n3830), .B(DATAO_REG_4__SCAN_IN), .S(n3833), .Z(U3554) );
  MUX2_X1 U4489 ( .A(n3831), .B(DATAO_REG_3__SCAN_IN), .S(n3833), .Z(U3553) );
  MUX2_X1 U4490 ( .A(n3832), .B(DATAO_REG_2__SCAN_IN), .S(n3833), .Z(U3552) );
  MUX2_X1 U4491 ( .A(n3834), .B(DATAO_REG_1__SCAN_IN), .S(n3833), .Z(U3551) );
  AOI22_X1 U4492 ( .A1(n4442), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3842) );
  OAI211_X1 U4493 ( .C1(n3843), .C2(n3835), .A(n4348), .B(n3853), .ZN(n3841)
         );
  OAI211_X1 U4494 ( .C1(n3838), .C2(n3837), .A(n4337), .B(n3836), .ZN(n3840)
         );
  NAND2_X1 U4495 ( .A1(n4315), .A2(n2008), .ZN(n3839) );
  NAND4_X1 U4496 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(U3241)
         );
  OR2_X1 U4497 ( .A1(n3844), .A2(n3843), .ZN(n3845) );
  OAI211_X1 U4498 ( .C1(n3846), .C2(n4242), .A(n4254), .B(n3845), .ZN(n3847)
         );
  OAI211_X1 U4499 ( .C1(IR_REG_0__SCAN_IN), .C2(n3848), .A(n3847), .B(U4043), 
        .ZN(n3870) );
  AOI22_X1 U4500 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4442), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3859) );
  XNOR2_X1 U4501 ( .A(n3850), .B(n3849), .ZN(n3851) );
  AOI22_X1 U4502 ( .A1(n4252), .A2(n4315), .B1(n4337), .B2(n3851), .ZN(n3858)
         );
  MUX2_X1 U4503 ( .A(n2928), .B(REG2_REG_2__SCAN_IN), .S(n4252), .Z(n3854) );
  NAND3_X1 U4504 ( .A1(n3854), .A2(n3853), .A3(n3852), .ZN(n3855) );
  NAND3_X1 U4505 ( .A1(n4348), .A2(n3856), .A3(n3855), .ZN(n3857) );
  NAND4_X1 U4506 ( .A1(n3870), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(U3242)
         );
  NAND2_X1 U4507 ( .A1(n4442), .A2(ADDR_REG_4__SCAN_IN), .ZN(n3869) );
  XNOR2_X1 U4508 ( .A(n3860), .B(REG2_REG_4__SCAN_IN), .ZN(n3861) );
  NAND2_X1 U4509 ( .A1(n4348), .A2(n3861), .ZN(n3867) );
  XNOR2_X1 U4510 ( .A(n3862), .B(REG1_REG_4__SCAN_IN), .ZN(n3863) );
  NAND2_X1 U4511 ( .A1(n4337), .A2(n3863), .ZN(n3866) );
  NAND2_X1 U4512 ( .A1(n4315), .A2(n4251), .ZN(n3865) );
  AND4_X1 U4513 ( .A1(n3867), .A2(n3866), .A3(n3865), .A4(n3864), .ZN(n3868)
         );
  NAND3_X1 U4514 ( .A1(n3870), .A2(n3869), .A3(n3868), .ZN(U3244) );
  INV_X1 U4515 ( .A(n3903), .ZN(n4376) );
  INV_X1 U4516 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4517 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4376), .B1(n3903), .B2(
        n3871), .ZN(n4342) );
  INV_X1 U4518 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4186) );
  AOI22_X1 U4519 ( .A1(n3902), .A2(REG1_REG_17__SCAN_IN), .B1(n4186), .B2(
        n4378), .ZN(n4335) );
  INV_X1 U4520 ( .A(n4386), .ZN(n4273) );
  NOR2_X1 U4521 ( .A1(n3874), .A2(n4273), .ZN(n3875) );
  NOR2_X1 U4522 ( .A1(n4266), .A2(n4265), .ZN(n4264) );
  INV_X1 U4523 ( .A(n3888), .ZN(n4385) );
  AOI22_X1 U4524 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4385), .B1(n3888), .B2(
        n4548), .ZN(n4275) );
  NOR2_X1 U4525 ( .A1(n3876), .A2(n4384), .ZN(n3877) );
  INV_X1 U4526 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4287) );
  AOI22_X1 U4527 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4383), .B1(n3897), .B2(
        n3878), .ZN(n4295) );
  INV_X1 U4528 ( .A(n4381), .ZN(n4444) );
  NOR2_X1 U4529 ( .A1(n3879), .A2(n4444), .ZN(n3880) );
  NOR2_X1 U4530 ( .A1(n3880), .A2(n4434), .ZN(n4308) );
  INV_X1 U4531 ( .A(n4314), .ZN(n4380) );
  INV_X1 U4532 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4533 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4380), .B1(n4314), .B2(
        n3881), .ZN(n4307) );
  NOR2_X1 U4534 ( .A1(n4308), .A2(n4307), .ZN(n4306) );
  NAND2_X1 U4535 ( .A1(n3882), .A2(n4379), .ZN(n3883) );
  INV_X1 U4536 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4323) );
  XNOR2_X1 U4537 ( .A(n4247), .B(REG1_REG_19__SCAN_IN), .ZN(n3884) );
  XNOR2_X1 U4538 ( .A(n3885), .B(n3884), .ZN(n3912) );
  NAND2_X1 U4539 ( .A1(REG2_REG_18__SCAN_IN), .A2(n3903), .ZN(n3886) );
  OAI21_X1 U4540 ( .B1(REG2_REG_18__SCAN_IN), .B2(n3903), .A(n3886), .ZN(n4346) );
  NOR2_X1 U4541 ( .A1(n3902), .A2(REG2_REG_17__SCAN_IN), .ZN(n3887) );
  AOI21_X1 U4542 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3902), .A(n3887), .ZN(n4332) );
  NOR2_X1 U4543 ( .A1(n3279), .A2(n4383), .ZN(n4300) );
  NAND2_X1 U4544 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3888), .ZN(n3893) );
  AOI22_X1 U4545 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3888), .B1(n4385), .B2(
        n3193), .ZN(n4282) );
  NAND2_X1 U4546 ( .A1(n4386), .A2(n3891), .ZN(n3892) );
  XNOR2_X1 U4547 ( .A(n4273), .B(n3891), .ZN(n4270) );
  NAND2_X1 U4548 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4270), .ZN(n4269) );
  NAND2_X1 U4549 ( .A1(n3892), .A2(n4269), .ZN(n4281) );
  NAND2_X1 U4550 ( .A1(n4282), .A2(n4281), .ZN(n4280) );
  NAND2_X1 U4551 ( .A1(n3894), .A2(n3895), .ZN(n3896) );
  NOR2_X1 U4552 ( .A1(n4444), .A2(n3898), .ZN(n3899) );
  XOR2_X1 U4553 ( .A(n4381), .B(n3898), .Z(n4439) );
  NOR2_X1 U4554 ( .A1(n2391), .A2(n4439), .ZN(n4438) );
  AOI22_X1 U4555 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4380), .B1(n4314), .B2(
        n3346), .ZN(n4310) );
  NOR2_X1 U4556 ( .A1(n4311), .A2(n4310), .ZN(n4309) );
  NAND2_X1 U4557 ( .A1(n3900), .A2(n4379), .ZN(n3901) );
  NAND2_X1 U4558 ( .A1(n4332), .A2(n4331), .ZN(n4330) );
  OAI21_X1 U4559 ( .B1(n3902), .B2(REG2_REG_17__SCAN_IN), .A(n4330), .ZN(n4345) );
  NOR2_X1 U4560 ( .A1(n4346), .A2(n4345), .ZN(n4344) );
  MUX2_X1 U4561 ( .A(REG2_REG_19__SCAN_IN), .B(n2449), .S(n4247), .Z(n3904) );
  XNOR2_X1 U4562 ( .A(n3905), .B(n3904), .ZN(n3910) );
  NAND2_X1 U4563 ( .A1(n4442), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3906) );
  OAI211_X1 U4564 ( .C1(n4445), .C2(n3908), .A(n3907), .B(n3906), .ZN(n3909)
         );
  AOI21_X1 U4565 ( .B1(n3910), .B2(n4348), .A(n3909), .ZN(n3911) );
  OAI21_X1 U4566 ( .B1(n3912), .B2(n4433), .A(n3911), .ZN(U3259) );
  INV_X1 U4567 ( .A(n3913), .ZN(n3914) );
  AOI21_X1 U4568 ( .B1(n3916), .B2(n3915), .A(n3914), .ZN(n3917) );
  XNOR2_X1 U4569 ( .A(n3917), .B(n3931), .ZN(n3922) );
  NAND2_X1 U4570 ( .A1(n4242), .A2(B_REG_SCAN_IN), .ZN(n3918) );
  AND2_X1 U4571 ( .A1(n4025), .A2(n3918), .ZN(n4124) );
  AOI22_X1 U4572 ( .A1(n4124), .A2(n3919), .B1(n4127), .B2(n3934), .ZN(n3921)
         );
  NAND2_X1 U4573 ( .A1(n3927), .A2(n4109), .ZN(n3920) );
  OAI211_X1 U4574 ( .C1(n3922), .C2(n4104), .A(n3921), .B(n3920), .ZN(n4140)
         );
  AOI21_X1 U4575 ( .B1(n3923), .B2(n4367), .A(n4140), .ZN(n3937) );
  NAND2_X1 U4576 ( .A1(n3929), .A2(n3928), .ZN(n3932) );
  XNOR2_X1 U4577 ( .A(n3932), .B(n3931), .ZN(n4139) );
  NAND2_X1 U4578 ( .A1(n4139), .A2(n4121), .ZN(n3936) );
  AOI22_X1 U4579 ( .A1(n4141), .A2(n4358), .B1(REG2_REG_29__SCAN_IN), .B2(
        n2009), .ZN(n3935) );
  OAI211_X1 U4580 ( .C1(n2009), .C2(n3937), .A(n3936), .B(n3935), .ZN(U3354)
         );
  XOR2_X1 U4581 ( .A(n3941), .B(n3938), .Z(n4149) );
  INV_X1 U4582 ( .A(n4149), .ZN(n3956) );
  OAI21_X1 U4583 ( .B1(n3958), .B2(n3940), .A(n3939), .ZN(n3942) );
  XNOR2_X1 U4584 ( .A(n3942), .B(n3941), .ZN(n3948) );
  AOI22_X1 U4585 ( .A1(n3944), .A2(n4109), .B1(n3943), .B2(n4127), .ZN(n3947)
         );
  NAND2_X1 U4586 ( .A1(n3945), .A2(n4025), .ZN(n3946) );
  OAI211_X1 U4587 ( .C1(n3948), .C2(n4104), .A(n3947), .B(n3946), .ZN(n4148)
         );
  INV_X1 U4588 ( .A(n3968), .ZN(n3951) );
  OAI21_X1 U4589 ( .B1(n3951), .B2(n3950), .A(n3949), .ZN(n4208) );
  AOI22_X1 U4590 ( .A1(n3952), .A2(n4367), .B1(REG2_REG_26__SCAN_IN), .B2(
        n2009), .ZN(n3953) );
  OAI21_X1 U4591 ( .B1(n4208), .B2(n4095), .A(n3953), .ZN(n3954) );
  AOI21_X1 U4592 ( .B1(n4148), .B2(n4263), .A(n3954), .ZN(n3955) );
  OAI21_X1 U4593 ( .B1(n3956), .B2(n4098), .A(n3955), .ZN(U3264) );
  XOR2_X1 U4594 ( .A(n3961), .B(n3957), .Z(n4153) );
  INV_X1 U4595 ( .A(n4153), .ZN(n3973) );
  INV_X1 U4596 ( .A(n3958), .ZN(n3960) );
  NAND2_X1 U4597 ( .A1(n3960), .A2(n3959), .ZN(n3962) );
  XNOR2_X1 U4598 ( .A(n3962), .B(n3961), .ZN(n3963) );
  NAND2_X1 U4599 ( .A1(n3963), .A2(n4032), .ZN(n3965) );
  AOI22_X1 U4600 ( .A1(n4001), .A2(n4109), .B1(n2503), .B2(n4127), .ZN(n3964)
         );
  OAI211_X1 U4601 ( .C1(n3966), .C2(n4101), .A(n3965), .B(n3964), .ZN(n4152)
         );
  NAND2_X1 U4602 ( .A1(n3985), .A2(n2503), .ZN(n3967) );
  NAND2_X1 U4603 ( .A1(n3968), .A2(n3967), .ZN(n4211) );
  AOI22_X1 U4604 ( .A1(n2009), .A2(REG2_REG_25__SCAN_IN), .B1(n3969), .B2(
        n4367), .ZN(n3970) );
  OAI21_X1 U4605 ( .B1(n4211), .B2(n4095), .A(n3970), .ZN(n3971) );
  AOI21_X1 U4606 ( .B1(n4152), .B2(n4263), .A(n3971), .ZN(n3972) );
  OAI21_X1 U4607 ( .B1(n3973), .B2(n4098), .A(n3972), .ZN(U3265) );
  XNOR2_X1 U4608 ( .A(n3974), .B(n3978), .ZN(n4156) );
  INV_X1 U4609 ( .A(n4156), .ZN(n3992) );
  INV_X1 U4610 ( .A(n3975), .ZN(n3976) );
  NOR2_X1 U4611 ( .A1(n3977), .A2(n3976), .ZN(n3979) );
  XNOR2_X1 U4612 ( .A(n3979), .B(n3978), .ZN(n3980) );
  NAND2_X1 U4613 ( .A1(n3980), .A2(n4032), .ZN(n3983) );
  AOI22_X1 U4614 ( .A1(n4026), .A2(n4109), .B1(n4127), .B2(n3981), .ZN(n3982)
         );
  OAI211_X1 U4615 ( .C1(n3984), .C2(n4101), .A(n3983), .B(n3982), .ZN(n4155)
         );
  OAI21_X1 U4616 ( .B1(n4007), .B2(n3986), .A(n3985), .ZN(n4214) );
  NOR2_X1 U4617 ( .A1(n4214), .A2(n4095), .ZN(n3990) );
  INV_X1 U4618 ( .A(REG2_REG_24__SCAN_IN), .ZN(n3988) );
  OAI22_X1 U4619 ( .A1(n4263), .A2(n3988), .B1(n3987), .B2(n4352), .ZN(n3989)
         );
  AOI211_X1 U4620 ( .C1(n4155), .C2(n4263), .A(n3990), .B(n3989), .ZN(n3991)
         );
  OAI21_X1 U4621 ( .B1(n3992), .B2(n4098), .A(n3991), .ZN(U3266) );
  XOR2_X1 U4622 ( .A(n3999), .B(n3993), .Z(n4160) );
  INV_X1 U4623 ( .A(n4160), .ZN(n4013) );
  OR2_X1 U4624 ( .A1(n4037), .A2(n3994), .ZN(n3997) );
  INV_X1 U4625 ( .A(n3995), .ZN(n3996) );
  NAND2_X1 U4626 ( .A1(n3997), .A2(n3996), .ZN(n4023) );
  INV_X1 U4627 ( .A(n4015), .ZN(n4024) );
  NAND2_X1 U4628 ( .A1(n4023), .A2(n4024), .ZN(n4022) );
  NAND2_X1 U4629 ( .A1(n4022), .A2(n3998), .ZN(n4000) );
  XNOR2_X1 U4630 ( .A(n4000), .B(n3999), .ZN(n4005) );
  AOI22_X1 U4631 ( .A1(n4001), .A2(n4025), .B1(n4006), .B2(n4127), .ZN(n4004)
         );
  NAND2_X1 U4632 ( .A1(n4002), .A2(n4109), .ZN(n4003) );
  OAI211_X1 U4633 ( .C1(n4005), .C2(n4104), .A(n4004), .B(n4003), .ZN(n4159)
         );
  AND2_X1 U4634 ( .A1(n4164), .A2(n4006), .ZN(n4008) );
  OR2_X1 U4635 ( .A1(n4008), .A2(n4007), .ZN(n4218) );
  AOI22_X1 U4636 ( .A1(n2009), .A2(REG2_REG_23__SCAN_IN), .B1(n4009), .B2(
        n4367), .ZN(n4010) );
  OAI21_X1 U4637 ( .B1(n4218), .B2(n4095), .A(n4010), .ZN(n4011) );
  AOI21_X1 U4638 ( .B1(n4159), .B2(n4263), .A(n4011), .ZN(n4012) );
  OAI21_X1 U4639 ( .B1(n4013), .B2(n4098), .A(n4012), .ZN(U3267) );
  OAI21_X1 U4640 ( .B1(n4016), .B2(n4015), .A(n4014), .ZN(n4167) );
  NAND2_X1 U4641 ( .A1(n4047), .A2(n4017), .ZN(n4163) );
  AND2_X1 U4642 ( .A1(n4163), .A2(n4358), .ZN(n4021) );
  OAI22_X1 U4643 ( .A1(n4263), .A2(n4019), .B1(n4018), .B2(n4352), .ZN(n4020)
         );
  AOI21_X1 U4644 ( .B1(n4021), .B2(n4164), .A(n4020), .ZN(n4035) );
  OAI21_X1 U4645 ( .B1(n4024), .B2(n4023), .A(n4022), .ZN(n4033) );
  NAND2_X1 U4646 ( .A1(n4026), .A2(n4025), .ZN(n4029) );
  NAND2_X1 U4647 ( .A1(n4027), .A2(n4109), .ZN(n4028) );
  OAI211_X1 U4648 ( .C1(n4134), .C2(n4030), .A(n4029), .B(n4028), .ZN(n4031)
         );
  AOI21_X1 U4649 ( .B1(n4033), .B2(n4032), .A(n4031), .ZN(n4166) );
  OR2_X1 U4650 ( .A1(n4166), .A2(n2009), .ZN(n4034) );
  OAI211_X1 U4651 ( .C1(n4167), .C2(n4098), .A(n4035), .B(n4034), .ZN(U3268)
         );
  XNOR2_X1 U4652 ( .A(n4036), .B(n4038), .ZN(n4169) );
  INV_X1 U4653 ( .A(n4169), .ZN(n4052) );
  XOR2_X1 U4654 ( .A(n4038), .B(n4037), .Z(n4044) );
  OAI22_X1 U4655 ( .A1(n4040), .A2(n4101), .B1(n4134), .B2(n4039), .ZN(n4041)
         );
  AOI21_X1 U4656 ( .B1(n4109), .B2(n4042), .A(n4041), .ZN(n4043) );
  OAI21_X1 U4657 ( .B1(n4044), .B2(n4104), .A(n4043), .ZN(n4168) );
  NAND2_X1 U4658 ( .A1(n4069), .A2(n4045), .ZN(n4046) );
  NAND2_X1 U4659 ( .A1(n4047), .A2(n4046), .ZN(n4223) );
  AOI22_X1 U4660 ( .A1(n2009), .A2(REG2_REG_21__SCAN_IN), .B1(n4048), .B2(
        n4367), .ZN(n4049) );
  OAI21_X1 U4661 ( .B1(n4223), .B2(n4095), .A(n4049), .ZN(n4050) );
  AOI21_X1 U4662 ( .B1(n4168), .B2(n4263), .A(n4050), .ZN(n4051) );
  OAI21_X1 U4663 ( .B1(n4052), .B2(n4098), .A(n4051), .ZN(U3269) );
  AOI22_X1 U4664 ( .A1(n4075), .A2(n4053), .B1(n4102), .B2(n4090), .ZN(n4054)
         );
  XOR2_X1 U4665 ( .A(n4059), .B(n4054), .Z(n4066) );
  OAI22_X1 U4666 ( .A1(n4055), .A2(n4101), .B1(n4134), .B2(n4067), .ZN(n4062)
         );
  NAND2_X1 U4667 ( .A1(n4057), .A2(n4056), .ZN(n4058) );
  XOR2_X1 U4668 ( .A(n4059), .B(n4058), .Z(n4060) );
  NOR2_X1 U4669 ( .A1(n4060), .A2(n4104), .ZN(n4061) );
  AOI211_X1 U4670 ( .C1(n4109), .C2(n4063), .A(n4062), .B(n4061), .ZN(n4064)
         );
  OAI21_X1 U4671 ( .B1(n4066), .B2(n4065), .A(n4064), .ZN(n4172) );
  INV_X1 U4672 ( .A(n4172), .ZN(n4074) );
  INV_X1 U4673 ( .A(n4066), .ZN(n4173) );
  OR2_X1 U4674 ( .A1(n4092), .A2(n4067), .ZN(n4068) );
  NAND2_X1 U4675 ( .A1(n4069), .A2(n4068), .ZN(n4227) );
  AOI22_X1 U4676 ( .A1(n2009), .A2(REG2_REG_20__SCAN_IN), .B1(n4070), .B2(
        n4367), .ZN(n4071) );
  OAI21_X1 U4677 ( .B1(n4227), .B2(n4095), .A(n4071), .ZN(n4072) );
  AOI21_X1 U4678 ( .B1(n4173), .B2(n4368), .A(n4072), .ZN(n4073) );
  OAI21_X1 U4679 ( .B1(n4074), .B2(n2009), .A(n4073), .ZN(U3270) );
  XNOR2_X1 U4680 ( .A(n4075), .B(n4084), .ZN(n4177) );
  INV_X1 U4681 ( .A(n4177), .ZN(n4099) );
  INV_X1 U4682 ( .A(n4076), .ZN(n4078) );
  OAI21_X1 U4683 ( .B1(n4079), .B2(n4078), .A(n4077), .ZN(n4103) );
  INV_X1 U4684 ( .A(n4080), .ZN(n4082) );
  OAI21_X1 U4685 ( .B1(n4103), .B2(n4082), .A(n4081), .ZN(n4083) );
  XOR2_X1 U4686 ( .A(n4084), .B(n4083), .Z(n4089) );
  OAI22_X1 U4687 ( .A1(n4085), .A2(n4101), .B1(n4134), .B2(n4090), .ZN(n4086)
         );
  AOI21_X1 U4688 ( .B1(n4109), .B2(n4087), .A(n4086), .ZN(n4088) );
  OAI21_X1 U4689 ( .B1(n4089), .B2(n4104), .A(n4088), .ZN(n4176) );
  AOI21_X1 U4690 ( .B1(n4114), .B2(n4100), .A(n4090), .ZN(n4091) );
  OR2_X1 U4691 ( .A1(n4092), .A2(n4091), .ZN(n4231) );
  AOI22_X1 U4692 ( .A1(n2009), .A2(REG2_REG_19__SCAN_IN), .B1(n4093), .B2(
        n4367), .ZN(n4094) );
  OAI21_X1 U4693 ( .B1(n4231), .B2(n4095), .A(n4094), .ZN(n4096) );
  AOI21_X1 U4694 ( .B1(n4176), .B2(n4263), .A(n4096), .ZN(n4097) );
  OAI21_X1 U4695 ( .B1(n4099), .B2(n4098), .A(n4097), .ZN(U3271) );
  OAI22_X1 U4696 ( .A1(n4102), .A2(n4101), .B1(n4134), .B2(n4100), .ZN(n4107)
         );
  XNOR2_X1 U4697 ( .A(n4103), .B(n4111), .ZN(n4105) );
  NOR2_X1 U4698 ( .A1(n4105), .A2(n4104), .ZN(n4106) );
  AOI211_X1 U4699 ( .C1(n4109), .C2(n4108), .A(n4107), .B(n4106), .ZN(n4182)
         );
  OAI21_X1 U4700 ( .B1(n4112), .B2(n4111), .A(n4110), .ZN(n4180) );
  XNOR2_X1 U4701 ( .A(n4114), .B(n4113), .ZN(n4115) );
  NAND2_X1 U4702 ( .A1(n4115), .A2(n4421), .ZN(n4181) );
  INV_X1 U4703 ( .A(n4116), .ZN(n4119) );
  AOI22_X1 U4704 ( .A1(n2009), .A2(REG2_REG_18__SCAN_IN), .B1(n4117), .B2(
        n4367), .ZN(n4118) );
  OAI21_X1 U4705 ( .B1(n4181), .B2(n4119), .A(n4118), .ZN(n4120) );
  AOI21_X1 U4706 ( .B1(n4180), .B2(n4121), .A(n4120), .ZN(n4122) );
  OAI21_X1 U4707 ( .B1(n2009), .B2(n4182), .A(n4122), .ZN(U3272) );
  NAND2_X1 U4708 ( .A1(n4132), .A2(n4135), .ZN(n4131) );
  XNOR2_X1 U4709 ( .A(n4131), .B(n4125), .ZN(n4256) );
  INV_X1 U4710 ( .A(n4256), .ZN(n4199) );
  NAND2_X1 U4711 ( .A1(n4124), .A2(n4123), .ZN(n4133) );
  INV_X1 U4712 ( .A(n4125), .ZN(n4126) );
  NAND2_X1 U4713 ( .A1(n4127), .A2(n4126), .ZN(n4128) );
  AND2_X1 U4714 ( .A1(n4133), .A2(n4128), .ZN(n4258) );
  INV_X1 U4715 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4129) );
  MUX2_X1 U4716 ( .A(n4258), .B(n4129), .S(n4430), .Z(n4130) );
  OAI21_X1 U4717 ( .B1(n4199), .B2(n4188), .A(n4130), .ZN(U3549) );
  OAI21_X1 U4718 ( .B1(n4132), .B2(n4135), .A(n4131), .ZN(n4259) );
  OAI21_X1 U4719 ( .B1(n4135), .B2(n4134), .A(n4133), .ZN(n4260) );
  INV_X1 U4720 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4136) );
  NOR2_X1 U4721 ( .A1(n4432), .A2(n4136), .ZN(n4137) );
  AOI21_X1 U4722 ( .B1(n4432), .B2(n4260), .A(n4137), .ZN(n4138) );
  OAI21_X1 U4723 ( .B1(n4259), .B2(n4188), .A(n4138), .ZN(U3548) );
  NAND2_X1 U4724 ( .A1(n4139), .A2(n4410), .ZN(n4143) );
  AOI21_X1 U4725 ( .B1(n4421), .B2(n4141), .A(n4140), .ZN(n4142) );
  NAND2_X1 U4726 ( .A1(n4143), .A2(n4142), .ZN(n4203) );
  MUX2_X1 U4727 ( .A(REG1_REG_29__SCAN_IN), .B(n4203), .S(n4432), .Z(U3547) );
  AOI21_X1 U4728 ( .B1(n4421), .B2(n4145), .A(n4144), .ZN(n4146) );
  OAI21_X1 U4729 ( .B1(n4147), .B2(n4416), .A(n4146), .ZN(n4204) );
  MUX2_X1 U4730 ( .A(REG1_REG_27__SCAN_IN), .B(n4204), .S(n4432), .Z(U3545) );
  INV_X1 U4731 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4150) );
  AOI21_X1 U4732 ( .B1(n4149), .B2(n4410), .A(n4148), .ZN(n4205) );
  MUX2_X1 U4733 ( .A(n4150), .B(n4205), .S(n4432), .Z(n4151) );
  OAI21_X1 U4734 ( .B1(n4188), .B2(n4208), .A(n4151), .ZN(U3544) );
  INV_X1 U4735 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4561) );
  AOI21_X1 U4736 ( .B1(n4153), .B2(n4410), .A(n4152), .ZN(n4209) );
  MUX2_X1 U4737 ( .A(n4561), .B(n4209), .S(n4432), .Z(n4154) );
  OAI21_X1 U4738 ( .B1(n4188), .B2(n4211), .A(n4154), .ZN(U3543) );
  INV_X1 U4739 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4157) );
  AOI21_X1 U4740 ( .B1(n4156), .B2(n4410), .A(n4155), .ZN(n4212) );
  MUX2_X1 U4741 ( .A(n4157), .B(n4212), .S(n4432), .Z(n4158) );
  OAI21_X1 U4742 ( .B1(n4188), .B2(n4214), .A(n4158), .ZN(U3542) );
  INV_X1 U4743 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4161) );
  AOI21_X1 U4744 ( .B1(n4160), .B2(n4410), .A(n4159), .ZN(n4215) );
  MUX2_X1 U4745 ( .A(n4161), .B(n4215), .S(n4432), .Z(n4162) );
  OAI21_X1 U4746 ( .B1(n4188), .B2(n4218), .A(n4162), .ZN(U3541) );
  NAND3_X1 U4747 ( .A1(n4164), .A2(n4421), .A3(n4163), .ZN(n4165) );
  OAI211_X1 U4748 ( .C1(n4167), .C2(n4416), .A(n4166), .B(n4165), .ZN(n4219)
         );
  MUX2_X1 U4749 ( .A(REG1_REG_22__SCAN_IN), .B(n4219), .S(n4432), .Z(U3540) );
  INV_X1 U4750 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4170) );
  AOI21_X1 U4751 ( .B1(n4169), .B2(n4410), .A(n4168), .ZN(n4220) );
  MUX2_X1 U4752 ( .A(n4170), .B(n4220), .S(n4432), .Z(n4171) );
  OAI21_X1 U4753 ( .B1(n4188), .B2(n4223), .A(n4171), .ZN(U3539) );
  INV_X1 U4754 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4174) );
  AOI21_X1 U4755 ( .B1(n4402), .B2(n4173), .A(n4172), .ZN(n4224) );
  MUX2_X1 U4756 ( .A(n4174), .B(n4224), .S(n4432), .Z(n4175) );
  OAI21_X1 U4757 ( .B1(n4188), .B2(n4227), .A(n4175), .ZN(U3538) );
  INV_X1 U4758 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4178) );
  AOI21_X1 U4759 ( .B1(n4177), .B2(n4410), .A(n4176), .ZN(n4228) );
  MUX2_X1 U4760 ( .A(n4178), .B(n4228), .S(n4432), .Z(n4179) );
  OAI21_X1 U4761 ( .B1(n4188), .B2(n4231), .A(n4179), .ZN(U3537) );
  INV_X1 U4762 ( .A(n4180), .ZN(n4183) );
  OAI211_X1 U4763 ( .C1(n4183), .C2(n4416), .A(n4182), .B(n4181), .ZN(n4232)
         );
  MUX2_X1 U4764 ( .A(REG1_REG_18__SCAN_IN), .B(n4232), .S(n4432), .Z(U3536) );
  AOI21_X1 U4765 ( .B1(n4185), .B2(n4410), .A(n4184), .ZN(n4233) );
  MUX2_X1 U4766 ( .A(n4186), .B(n4233), .S(n4432), .Z(n4187) );
  OAI21_X1 U4767 ( .B1(n4188), .B2(n4237), .A(n4187), .ZN(U3535) );
  AOI21_X1 U4768 ( .B1(n4421), .B2(n4190), .A(n4189), .ZN(n4191) );
  OAI21_X1 U4769 ( .B1(n4192), .B2(n4416), .A(n4191), .ZN(n4238) );
  MUX2_X1 U4770 ( .A(REG1_REG_16__SCAN_IN), .B(n4238), .S(n4432), .Z(U3534) );
  NAND2_X1 U4771 ( .A1(n4193), .A2(n4421), .ZN(n4194) );
  OAI211_X1 U4772 ( .C1(n4196), .C2(n4416), .A(n4195), .B(n4194), .ZN(n4239)
         );
  MUX2_X1 U4773 ( .A(REG1_REG_15__SCAN_IN), .B(n4239), .S(n4432), .Z(U3533) );
  INV_X1 U4774 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4197) );
  MUX2_X1 U4775 ( .A(n4258), .B(n4197), .S(n4422), .Z(n4198) );
  OAI21_X1 U4776 ( .B1(n4199), .B2(n4236), .A(n4198), .ZN(U3517) );
  INV_X1 U4777 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4200) );
  NOR2_X1 U4778 ( .A1(n4423), .A2(n4200), .ZN(n4201) );
  AOI21_X1 U4779 ( .B1(n4423), .B2(n4260), .A(n4201), .ZN(n4202) );
  OAI21_X1 U4780 ( .B1(n4259), .B2(n4236), .A(n4202), .ZN(U3516) );
  MUX2_X1 U4781 ( .A(REG0_REG_29__SCAN_IN), .B(n4203), .S(n4423), .Z(U3515) );
  MUX2_X1 U4782 ( .A(REG0_REG_27__SCAN_IN), .B(n4204), .S(n4423), .Z(U3513) );
  INV_X1 U4783 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4206) );
  MUX2_X1 U4784 ( .A(n4206), .B(n4205), .S(n4423), .Z(n4207) );
  OAI21_X1 U4785 ( .B1(n4208), .B2(n4236), .A(n4207), .ZN(U3512) );
  INV_X1 U4786 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4451) );
  MUX2_X1 U4787 ( .A(n4451), .B(n4209), .S(n4423), .Z(n4210) );
  OAI21_X1 U4788 ( .B1(n4211), .B2(n4236), .A(n4210), .ZN(U3511) );
  INV_X1 U4789 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4565) );
  MUX2_X1 U4790 ( .A(n4565), .B(n4212), .S(n4423), .Z(n4213) );
  OAI21_X1 U4791 ( .B1(n4214), .B2(n4236), .A(n4213), .ZN(U3510) );
  INV_X1 U4792 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4216) );
  MUX2_X1 U4793 ( .A(n4216), .B(n4215), .S(n4423), .Z(n4217) );
  OAI21_X1 U4794 ( .B1(n4218), .B2(n4236), .A(n4217), .ZN(U3509) );
  MUX2_X1 U4795 ( .A(REG0_REG_22__SCAN_IN), .B(n4219), .S(n4423), .Z(U3508) );
  INV_X1 U4796 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4221) );
  MUX2_X1 U4797 ( .A(n4221), .B(n4220), .S(n4423), .Z(n4222) );
  OAI21_X1 U4798 ( .B1(n4223), .B2(n4236), .A(n4222), .ZN(U3507) );
  INV_X1 U4799 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4225) );
  MUX2_X1 U4800 ( .A(n4225), .B(n4224), .S(n4423), .Z(n4226) );
  OAI21_X1 U4801 ( .B1(n4227), .B2(n4236), .A(n4226), .ZN(U3506) );
  INV_X1 U4802 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4229) );
  MUX2_X1 U4803 ( .A(n4229), .B(n4228), .S(n4423), .Z(n4230) );
  OAI21_X1 U4804 ( .B1(n4231), .B2(n4236), .A(n4230), .ZN(U3505) );
  MUX2_X1 U4805 ( .A(REG0_REG_18__SCAN_IN), .B(n4232), .S(n4423), .Z(U3503) );
  INV_X1 U4806 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4234) );
  MUX2_X1 U4807 ( .A(n4234), .B(n4233), .S(n4423), .Z(n4235) );
  OAI21_X1 U4808 ( .B1(n4237), .B2(n4236), .A(n4235), .ZN(U3501) );
  MUX2_X1 U4809 ( .A(REG0_REG_16__SCAN_IN), .B(n4238), .S(n4423), .Z(U3499) );
  MUX2_X1 U4810 ( .A(REG0_REG_15__SCAN_IN), .B(n4239), .S(n4423), .Z(U3497) );
  MUX2_X1 U4811 ( .A(DATAI_30_), .B(n4240), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4812 ( .A(DATAI_29_), .B(n4241), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U4813 ( .A(n4242), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U4814 ( .A(n4243), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4815 ( .A(n4244), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U4816 ( .A(n4245), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U4817 ( .A(DATAI_20_), .B(n4246), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4818 ( .A(n4247), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4819 ( .A(DATAI_8_), .B(n4248), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U4820 ( .A(n4249), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4821 ( .A(n4250), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4822 ( .A(DATAI_4_), .B(n4251), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4823 ( .A(n4252), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4824 ( .A(n2008), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  OAI22_X1 U4825 ( .A1(U3149), .A2(n4254), .B1(DATAI_28_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4255) );
  INV_X1 U4826 ( .A(n4255), .ZN(U3324) );
  AOI22_X1 U4827 ( .A1(n4256), .A2(n4358), .B1(n2009), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4257) );
  OAI21_X1 U4828 ( .B1(n2009), .B2(n4258), .A(n4257), .ZN(U3260) );
  INV_X1 U4829 ( .A(n4259), .ZN(n4261) );
  AOI22_X1 U4830 ( .A1(n4261), .A2(n4358), .B1(n4263), .B2(n4260), .ZN(n4262)
         );
  OAI21_X1 U4831 ( .B1(n3669), .B2(n4263), .A(n4262), .ZN(U3261) );
  AOI211_X1 U4832 ( .C1(n4266), .C2(n4265), .A(n4264), .B(n4433), .ZN(n4267)
         );
  AOI211_X1 U4833 ( .C1(n4442), .C2(ADDR_REG_10__SCAN_IN), .A(n4268), .B(n4267), .ZN(n4272) );
  OAI211_X1 U4834 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4270), .A(n4348), .B(n4269), .ZN(n4271) );
  OAI211_X1 U4835 ( .C1(n4445), .C2(n4273), .A(n4272), .B(n4271), .ZN(U3250)
         );
  AOI211_X1 U4836 ( .C1(n4276), .C2(n4275), .A(n4274), .B(n4433), .ZN(n4279)
         );
  INV_X1 U4837 ( .A(n4277), .ZN(n4278) );
  AOI211_X1 U4838 ( .C1(n4442), .C2(ADDR_REG_11__SCAN_IN), .A(n4279), .B(n4278), .ZN(n4284) );
  OAI211_X1 U4839 ( .C1(n4282), .C2(n4281), .A(n4348), .B(n4280), .ZN(n4283)
         );
  OAI211_X1 U4840 ( .C1(n4445), .C2(n4385), .A(n4284), .B(n4283), .ZN(U3251)
         );
  AOI211_X1 U4841 ( .C1(n4287), .C2(n4286), .A(n4285), .B(n4433), .ZN(n4289)
         );
  AOI211_X1 U4842 ( .C1(n4442), .C2(ADDR_REG_12__SCAN_IN), .A(n4289), .B(n4288), .ZN(n4293) );
  OAI211_X1 U4843 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4291), .A(n4348), .B(n4290), .ZN(n4292) );
  OAI211_X1 U4844 ( .C1(n4445), .C2(n4384), .A(n4293), .B(n4292), .ZN(U3252)
         );
  AOI211_X1 U4845 ( .C1(n4296), .C2(n4295), .A(n4294), .B(n4433), .ZN(n4299)
         );
  INV_X1 U4846 ( .A(n4297), .ZN(n4298) );
  AOI211_X1 U4847 ( .C1(n4442), .C2(ADDR_REG_13__SCAN_IN), .A(n4299), .B(n4298), .ZN(n4305) );
  AOI21_X1 U4848 ( .B1(n3279), .B2(n4383), .A(n4300), .ZN(n4303) );
  AOI21_X1 U4849 ( .B1(n4303), .B2(n4302), .A(n4437), .ZN(n4301) );
  OAI21_X1 U4850 ( .B1(n4303), .B2(n4302), .A(n4301), .ZN(n4304) );
  OAI211_X1 U4851 ( .C1(n4445), .C2(n4383), .A(n4305), .B(n4304), .ZN(U3253)
         );
  INV_X1 U4852 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4462) );
  AOI211_X1 U4853 ( .C1(n4308), .C2(n4307), .A(n4306), .B(n4433), .ZN(n4313)
         );
  AOI211_X1 U4854 ( .C1(n4311), .C2(n4310), .A(n4309), .B(n4437), .ZN(n4312)
         );
  AOI211_X1 U4855 ( .C1(n4315), .C2(n4314), .A(n4313), .B(n4312), .ZN(n4317)
         );
  NAND2_X1 U4856 ( .A1(REG3_REG_15__SCAN_IN), .A2(U3149), .ZN(n4316) );
  OAI211_X1 U4857 ( .C1(n4318), .C2(n4462), .A(n4317), .B(n4316), .ZN(U3255)
         );
  AOI21_X1 U4858 ( .B1(n4442), .B2(ADDR_REG_16__SCAN_IN), .A(n4319), .ZN(n4328) );
  OAI21_X1 U4859 ( .B1(n4321), .B2(n3296), .A(n4320), .ZN(n4326) );
  OAI21_X1 U4860 ( .B1(n4324), .B2(n4323), .A(n4322), .ZN(n4325) );
  AOI22_X1 U4861 ( .A1(n4348), .A2(n4326), .B1(n4337), .B2(n4325), .ZN(n4327)
         );
  OAI211_X1 U4862 ( .C1(n4379), .C2(n4445), .A(n4328), .B(n4327), .ZN(U3256)
         );
  AOI21_X1 U4863 ( .B1(n4442), .B2(ADDR_REG_17__SCAN_IN), .A(n4329), .ZN(n4340) );
  OAI21_X1 U4864 ( .B1(n4332), .B2(n4331), .A(n4330), .ZN(n4338) );
  OAI21_X1 U4865 ( .B1(n4335), .B2(n4334), .A(n4333), .ZN(n4336) );
  AOI22_X1 U4866 ( .A1(n4348), .A2(n4338), .B1(n4337), .B2(n4336), .ZN(n4339)
         );
  OAI211_X1 U4867 ( .C1(n4378), .C2(n4445), .A(n4340), .B(n4339), .ZN(U3257)
         );
  AOI21_X1 U4868 ( .B1(n4346), .B2(n4345), .A(n4344), .ZN(n4347) );
  NAND2_X1 U4869 ( .A1(n4348), .A2(n4347), .ZN(n4349) );
  OAI211_X1 U4870 ( .C1(n4445), .C2(n4376), .A(n4350), .B(n4349), .ZN(U3258)
         );
  INV_X1 U4871 ( .A(n4351), .ZN(n4353) );
  OAI22_X1 U4872 ( .A1(n4263), .A2(n4354), .B1(n4353), .B2(n4352), .ZN(n4355)
         );
  INV_X1 U4873 ( .A(n4355), .ZN(n4361) );
  INV_X1 U4874 ( .A(n4356), .ZN(n4357) );
  AOI22_X1 U4875 ( .A1(n4359), .A2(n4368), .B1(n4358), .B2(n4357), .ZN(n4360)
         );
  OAI211_X1 U4876 ( .C1(n2009), .C2(n4362), .A(n4361), .B(n4360), .ZN(U3284)
         );
  INV_X1 U4877 ( .A(n4363), .ZN(n4365) );
  AOI21_X1 U4878 ( .B1(n4366), .B2(n4365), .A(n4364), .ZN(n4371) );
  AOI22_X1 U4879 ( .A1(n4369), .A2(n4368), .B1(REG3_REG_0__SCAN_IN), .B2(n4367), .ZN(n4370) );
  OAI221_X1 U4880 ( .B1(n2009), .B2(n4371), .C1(n4263), .C2(n2252), .A(n4370), 
        .ZN(U3290) );
  INV_X1 U4881 ( .A(n4373), .ZN(n4372) );
  INV_X1 U4882 ( .A(D_REG_31__SCAN_IN), .ZN(n4532) );
  NOR2_X1 U4883 ( .A1(n4372), .A2(n4532), .ZN(U3291) );
  AND2_X1 U4884 ( .A1(D_REG_30__SCAN_IN), .A2(n4373), .ZN(U3292) );
  AND2_X1 U4885 ( .A1(D_REG_29__SCAN_IN), .A2(n4373), .ZN(U3293) );
  INV_X1 U4886 ( .A(D_REG_28__SCAN_IN), .ZN(n4533) );
  NOR2_X1 U4887 ( .A1(n4372), .A2(n4533), .ZN(U3294) );
  AND2_X1 U4888 ( .A1(D_REG_27__SCAN_IN), .A2(n4373), .ZN(U3295) );
  INV_X1 U4889 ( .A(D_REG_26__SCAN_IN), .ZN(n4529) );
  NOR2_X1 U4890 ( .A1(n4372), .A2(n4529), .ZN(U3296) );
  AND2_X1 U4891 ( .A1(D_REG_25__SCAN_IN), .A2(n4373), .ZN(U3297) );
  AND2_X1 U4892 ( .A1(D_REG_24__SCAN_IN), .A2(n4373), .ZN(U3298) );
  AND2_X1 U4893 ( .A1(D_REG_23__SCAN_IN), .A2(n4373), .ZN(U3299) );
  INV_X1 U4894 ( .A(D_REG_22__SCAN_IN), .ZN(n4530) );
  NOR2_X1 U4895 ( .A1(n4372), .A2(n4530), .ZN(U3300) );
  AND2_X1 U4896 ( .A1(D_REG_21__SCAN_IN), .A2(n4373), .ZN(U3301) );
  AND2_X1 U4897 ( .A1(D_REG_20__SCAN_IN), .A2(n4373), .ZN(U3302) );
  AND2_X1 U4898 ( .A1(D_REG_19__SCAN_IN), .A2(n4373), .ZN(U3303) );
  AND2_X1 U4899 ( .A1(D_REG_18__SCAN_IN), .A2(n4373), .ZN(U3304) );
  AND2_X1 U4900 ( .A1(D_REG_17__SCAN_IN), .A2(n4373), .ZN(U3305) );
  AND2_X1 U4901 ( .A1(D_REG_16__SCAN_IN), .A2(n4373), .ZN(U3306) );
  INV_X1 U4902 ( .A(D_REG_15__SCAN_IN), .ZN(n4526) );
  NOR2_X1 U4903 ( .A1(n4372), .A2(n4526), .ZN(U3307) );
  INV_X1 U4904 ( .A(D_REG_14__SCAN_IN), .ZN(n4527) );
  NOR2_X1 U4905 ( .A1(n4372), .A2(n4527), .ZN(U3308) );
  AND2_X1 U4906 ( .A1(D_REG_13__SCAN_IN), .A2(n4373), .ZN(U3309) );
  AND2_X1 U4907 ( .A1(D_REG_12__SCAN_IN), .A2(n4373), .ZN(U3310) );
  AND2_X1 U4908 ( .A1(D_REG_11__SCAN_IN), .A2(n4373), .ZN(U3311) );
  INV_X1 U4909 ( .A(D_REG_10__SCAN_IN), .ZN(n4513) );
  NOR2_X1 U4910 ( .A1(n4372), .A2(n4513), .ZN(U3312) );
  AND2_X1 U4911 ( .A1(D_REG_9__SCAN_IN), .A2(n4373), .ZN(U3313) );
  AND2_X1 U4912 ( .A1(D_REG_8__SCAN_IN), .A2(n4373), .ZN(U3314) );
  AND2_X1 U4913 ( .A1(D_REG_7__SCAN_IN), .A2(n4373), .ZN(U3315) );
  AND2_X1 U4914 ( .A1(D_REG_6__SCAN_IN), .A2(n4373), .ZN(U3316) );
  AND2_X1 U4915 ( .A1(D_REG_5__SCAN_IN), .A2(n4373), .ZN(U3317) );
  INV_X1 U4916 ( .A(D_REG_4__SCAN_IN), .ZN(n4514) );
  NOR2_X1 U4917 ( .A1(n4372), .A2(n4514), .ZN(U3318) );
  AND2_X1 U4918 ( .A1(D_REG_3__SCAN_IN), .A2(n4373), .ZN(U3319) );
  AND2_X1 U4919 ( .A1(D_REG_2__SCAN_IN), .A2(n4373), .ZN(U3320) );
  INV_X1 U4920 ( .A(DATAI_23_), .ZN(n4375) );
  AOI21_X1 U4921 ( .B1(U3149), .B2(n4375), .A(n4374), .ZN(U3329) );
  INV_X1 U4922 ( .A(DATAI_18_), .ZN(n4491) );
  AOI22_X1 U4923 ( .A1(STATE_REG_SCAN_IN), .A2(n4376), .B1(n4491), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U4924 ( .A1(STATE_REG_SCAN_IN), .A2(n4378), .B1(n4377), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U4925 ( .A(DATAI_16_), .ZN(n4493) );
  AOI22_X1 U4926 ( .A1(STATE_REG_SCAN_IN), .A2(n4379), .B1(n4493), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U4927 ( .A(DATAI_15_), .ZN(n4575) );
  AOI22_X1 U4928 ( .A1(STATE_REG_SCAN_IN), .A2(n4380), .B1(n4575), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U4929 ( .A1(U3149), .A2(n4381), .B1(DATAI_14_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4382) );
  INV_X1 U4930 ( .A(n4382), .ZN(U3338) );
  AOI22_X1 U4931 ( .A1(STATE_REG_SCAN_IN), .A2(n4383), .B1(n2233), .B2(U3149), 
        .ZN(U3339) );
  AOI22_X1 U4932 ( .A1(STATE_REG_SCAN_IN), .A2(n4384), .B1(n4577), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U4933 ( .A(DATAI_11_), .ZN(n4579) );
  AOI22_X1 U4934 ( .A1(STATE_REG_SCAN_IN), .A2(n4385), .B1(n4579), .B2(U3149), 
        .ZN(U3341) );
  OAI22_X1 U4935 ( .A1(U3149), .A2(n4386), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4387) );
  INV_X1 U4936 ( .A(n4387), .ZN(U3342) );
  OAI22_X1 U4937 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4388) );
  INV_X1 U4938 ( .A(n4388), .ZN(U3352) );
  INV_X1 U4939 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4578) );
  AOI22_X1 U4940 ( .A1(n4423), .A2(n4389), .B1(n4578), .B2(n4422), .ZN(U3467)
         );
  INV_X1 U4941 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4390) );
  AOI22_X1 U4942 ( .A1(n4423), .A2(n4391), .B1(n4390), .B2(n4422), .ZN(U3469)
         );
  OAI22_X1 U4943 ( .A1(n4395), .A2(n4394), .B1(n4393), .B2(n4392), .ZN(n4396)
         );
  NOR2_X1 U4944 ( .A1(n4397), .A2(n4396), .ZN(n4425) );
  INV_X1 U4945 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4535) );
  AOI22_X1 U4946 ( .A1(n4423), .A2(n4425), .B1(n4535), .B2(n4422), .ZN(U3473)
         );
  INV_X1 U4947 ( .A(n4398), .ZN(n4403) );
  INV_X1 U4948 ( .A(n4399), .ZN(n4401) );
  AOI211_X1 U4949 ( .C1(n4403), .C2(n4402), .A(n4401), .B(n4400), .ZN(n4426)
         );
  INV_X1 U4950 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4449) );
  AOI22_X1 U4951 ( .A1(n4423), .A2(n4426), .B1(n4449), .B2(n4422), .ZN(U3475)
         );
  NOR2_X1 U4952 ( .A1(n4404), .A2(n4416), .ZN(n4407) );
  INV_X1 U4953 ( .A(n4405), .ZN(n4406) );
  AOI211_X1 U4954 ( .C1(n4421), .C2(n4408), .A(n4407), .B(n4406), .ZN(n4427)
         );
  INV_X1 U4955 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4409) );
  AOI22_X1 U4956 ( .A1(n4423), .A2(n4427), .B1(n4409), .B2(n4422), .ZN(U3477)
         );
  NAND3_X1 U4957 ( .A1(n2889), .A2(n4411), .A3(n4410), .ZN(n4412) );
  AND3_X1 U4958 ( .A1(n4414), .A2(n4413), .A3(n4412), .ZN(n4429) );
  INV_X1 U4959 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4415) );
  AOI22_X1 U4960 ( .A1(n4423), .A2(n4429), .B1(n4415), .B2(n4422), .ZN(U3481)
         );
  NOR2_X1 U4961 ( .A1(n4417), .A2(n4416), .ZN(n4419) );
  AOI211_X1 U4962 ( .C1(n4421), .C2(n4420), .A(n4419), .B(n4418), .ZN(n4431)
         );
  INV_X1 U4963 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4562) );
  AOI22_X1 U4964 ( .A1(n4423), .A2(n4431), .B1(n4562), .B2(n4422), .ZN(U3485)
         );
  INV_X1 U4965 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4424) );
  AOI22_X1 U4966 ( .A1(n4432), .A2(n4425), .B1(n4424), .B2(n4430), .ZN(U3521)
         );
  AOI22_X1 U4967 ( .A1(n4432), .A2(n4426), .B1(n2685), .B2(n4430), .ZN(U3522)
         );
  AOI22_X1 U4968 ( .A1(n4432), .A2(n4427), .B1(n2688), .B2(n4430), .ZN(U3523)
         );
  AOI22_X1 U4969 ( .A1(n4432), .A2(n4429), .B1(n4428), .B2(n4430), .ZN(U3525)
         );
  AOI22_X1 U4970 ( .A1(n4432), .A2(n4431), .B1(n2805), .B2(n4430), .ZN(U3527)
         );
  AOI211_X1 U4971 ( .C1(n4436), .C2(n4435), .A(n4434), .B(n4433), .ZN(n4447)
         );
  AOI211_X1 U4972 ( .C1(n2391), .C2(n4439), .A(n4438), .B(n4437), .ZN(n4440)
         );
  AOI211_X1 U4973 ( .C1(n4442), .C2(ADDR_REG_14__SCAN_IN), .A(n4441), .B(n4440), .ZN(n4443) );
  OAI21_X1 U4974 ( .B1(n4445), .B2(n4444), .A(n4443), .ZN(n4446) );
  NOR2_X1 U4975 ( .A1(n4447), .A2(n4446), .ZN(n4597) );
  AOI22_X1 U4976 ( .A1(n4449), .A2(keyinput59), .B1(n4562), .B2(keyinput6), 
        .ZN(n4448) );
  OAI221_X1 U4977 ( .B1(n4449), .B2(keyinput59), .C1(n4562), .C2(keyinput6), 
        .A(n4448), .ZN(n4459) );
  AOI22_X1 U4978 ( .A1(n4565), .A2(keyinput35), .B1(n4451), .B2(keyinput31), 
        .ZN(n4450) );
  OAI221_X1 U4979 ( .B1(n4565), .B2(keyinput35), .C1(n4451), .C2(keyinput31), 
        .A(n4450), .ZN(n4458) );
  INV_X1 U4980 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4563) );
  INV_X1 U4981 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4564) );
  AOI22_X1 U4982 ( .A1(n4563), .A2(keyinput46), .B1(n4564), .B2(keyinput42), 
        .ZN(n4452) );
  OAI221_X1 U4983 ( .B1(n4563), .B2(keyinput46), .C1(n4564), .C2(keyinput42), 
        .A(n4452), .ZN(n4457) );
  XOR2_X1 U4984 ( .A(n4453), .B(keyinput11), .Z(n4455) );
  XNOR2_X1 U4985 ( .A(REG1_REG_2__SCAN_IN), .B(keyinput27), .ZN(n4454) );
  NAND2_X1 U4986 ( .A1(n4455), .A2(n4454), .ZN(n4456) );
  NOR4_X1 U4987 ( .A1(n4459), .A2(n4458), .A3(n4457), .A4(n4456), .ZN(n4558)
         );
  INV_X1 U4988 ( .A(ADDR_REG_10__SCAN_IN), .ZN(n4461) );
  OAI22_X1 U4989 ( .A1(n4462), .A2(keyinput7), .B1(n4461), .B2(keyinput38), 
        .ZN(n4460) );
  AOI221_X1 U4990 ( .B1(n4462), .B2(keyinput7), .C1(keyinput38), .C2(n4461), 
        .A(n4460), .ZN(n4473) );
  OAI22_X1 U4991 ( .A1(keyinput15), .A2(n2719), .B1(n4464), .B2(keyinput5), 
        .ZN(n4463) );
  AOI221_X1 U4992 ( .B1(n2719), .B2(keyinput15), .C1(n4464), .C2(keyinput5), 
        .A(n4463), .ZN(n4472) );
  OAI22_X1 U4993 ( .A1(n2664), .A2(keyinput50), .B1(n4466), .B2(keyinput55), 
        .ZN(n4465) );
  AOI221_X1 U4994 ( .B1(n2664), .B2(keyinput50), .C1(keyinput55), .C2(n4466), 
        .A(n4465), .ZN(n4471) );
  OAI22_X1 U4995 ( .A1(n4469), .A2(keyinput48), .B1(n4468), .B2(keyinput14), 
        .ZN(n4467) );
  AOI221_X1 U4996 ( .B1(n4469), .B2(keyinput48), .C1(keyinput14), .C2(n4468), 
        .A(n4467), .ZN(n4470) );
  NAND4_X1 U4997 ( .A1(n4473), .A2(n4472), .A3(n4471), .A4(n4470), .ZN(n4546)
         );
  OAI22_X1 U4998 ( .A1(n4476), .A2(keyinput45), .B1(n4475), .B2(keyinput39), 
        .ZN(n4474) );
  AOI221_X1 U4999 ( .B1(n4476), .B2(keyinput45), .C1(keyinput39), .C2(n4475), 
        .A(n4474), .ZN(n4489) );
  OAI22_X1 U5000 ( .A1(n4479), .A2(keyinput17), .B1(n4478), .B2(keyinput12), 
        .ZN(n4477) );
  AOI221_X1 U5001 ( .B1(n4479), .B2(keyinput17), .C1(keyinput12), .C2(n4478), 
        .A(n4477), .ZN(n4488) );
  OAI22_X1 U5002 ( .A1(n4482), .A2(keyinput44), .B1(n4481), .B2(keyinput54), 
        .ZN(n4480) );
  AOI221_X1 U5003 ( .B1(n4482), .B2(keyinput44), .C1(keyinput54), .C2(n4481), 
        .A(n4480), .ZN(n4487) );
  OAI22_X1 U5004 ( .A1(n4485), .A2(keyinput13), .B1(n4484), .B2(keyinput10), 
        .ZN(n4483) );
  AOI221_X1 U5005 ( .B1(n4485), .B2(keyinput13), .C1(keyinput10), .C2(n4484), 
        .A(n4483), .ZN(n4486) );
  NAND4_X1 U5006 ( .A1(n4489), .A2(n4488), .A3(n4487), .A4(n4486), .ZN(n4545)
         );
  INV_X1 U5007 ( .A(DATAI_26_), .ZN(n4574) );
  AOI22_X1 U5008 ( .A1(n4574), .A2(keyinput18), .B1(n4491), .B2(keyinput25), 
        .ZN(n4490) );
  OAI221_X1 U5009 ( .B1(n4574), .B2(keyinput18), .C1(n4491), .C2(keyinput25), 
        .A(n4490), .ZN(n4500) );
  AOI22_X1 U5010 ( .A1(n4575), .A2(keyinput43), .B1(n4493), .B2(keyinput29), 
        .ZN(n4492) );
  OAI221_X1 U5011 ( .B1(n4575), .B2(keyinput43), .C1(n4493), .C2(keyinput29), 
        .A(n4492), .ZN(n4499) );
  AOI22_X1 U5012 ( .A1(n4577), .A2(keyinput56), .B1(keyinput26), .B2(n4579), 
        .ZN(n4494) );
  OAI221_X1 U5013 ( .B1(n4577), .B2(keyinput56), .C1(n4579), .C2(keyinput26), 
        .A(n4494), .ZN(n4498) );
  AOI22_X1 U5014 ( .A1(n4576), .A2(keyinput36), .B1(n4496), .B2(keyinput9), 
        .ZN(n4495) );
  OAI221_X1 U5015 ( .B1(n4576), .B2(keyinput36), .C1(n4496), .C2(keyinput9), 
        .A(n4495), .ZN(n4497) );
  NOR4_X1 U5016 ( .A1(n4500), .A2(n4499), .A3(n4498), .A4(n4497), .ZN(n4543)
         );
  AOI22_X1 U5017 ( .A1(n2467), .A2(keyinput16), .B1(keyinput23), .B2(n2412), 
        .ZN(n4501) );
  OAI221_X1 U5018 ( .B1(n2467), .B2(keyinput16), .C1(n2412), .C2(keyinput23), 
        .A(n4501), .ZN(n4511) );
  INV_X1 U5019 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4503) );
  AOI22_X1 U5020 ( .A1(n4504), .A2(keyinput51), .B1(keyinput34), .B2(n4503), 
        .ZN(n4502) );
  OAI221_X1 U5021 ( .B1(n4504), .B2(keyinput51), .C1(n4503), .C2(keyinput34), 
        .A(n4502), .ZN(n4510) );
  XOR2_X1 U5022 ( .A(n2221), .B(keyinput33), .Z(n4508) );
  XNOR2_X1 U5023 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput32), .ZN(n4507) );
  XNOR2_X1 U5024 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput30), .ZN(n4506) );
  XNOR2_X1 U5025 ( .A(IR_REG_6__SCAN_IN), .B(keyinput0), .ZN(n4505) );
  NAND4_X1 U5026 ( .A1(n4508), .A2(n4507), .A3(n4506), .A4(n4505), .ZN(n4509)
         );
  NOR3_X1 U5027 ( .A1(n4511), .A2(n4510), .A3(n4509), .ZN(n4542) );
  AOI22_X1 U5028 ( .A1(n4514), .A2(keyinput22), .B1(keyinput21), .B2(n4513), 
        .ZN(n4512) );
  OAI221_X1 U5029 ( .B1(n4514), .B2(keyinput22), .C1(n4513), .C2(keyinput21), 
        .A(n4512), .ZN(n4524) );
  INV_X1 U5030 ( .A(IR_REG_12__SCAN_IN), .ZN(n4516) );
  AOI22_X1 U5031 ( .A1(n2382), .A2(keyinput4), .B1(keyinput57), .B2(n4516), 
        .ZN(n4515) );
  OAI221_X1 U5032 ( .B1(n2382), .B2(keyinput4), .C1(n4516), .C2(keyinput57), 
        .A(n4515), .ZN(n4523) );
  AOI22_X1 U5033 ( .A1(n4518), .A2(keyinput49), .B1(n2226), .B2(keyinput41), 
        .ZN(n4517) );
  OAI221_X1 U5034 ( .B1(n4518), .B2(keyinput49), .C1(n2226), .C2(keyinput41), 
        .A(n4517), .ZN(n4522) );
  XOR2_X1 U5035 ( .A(n2235), .B(keyinput53), .Z(n4520) );
  XNOR2_X1 U5036 ( .A(IR_REG_24__SCAN_IN), .B(keyinput47), .ZN(n4519) );
  NAND2_X1 U5037 ( .A1(n4520), .A2(n4519), .ZN(n4521) );
  NOR4_X1 U5038 ( .A1(n4524), .A2(n4523), .A3(n4522), .A4(n4521), .ZN(n4541)
         );
  AOI22_X1 U5039 ( .A1(n4527), .A2(keyinput61), .B1(keyinput24), .B2(n4526), 
        .ZN(n4525) );
  OAI221_X1 U5040 ( .B1(n4527), .B2(keyinput61), .C1(n4526), .C2(keyinput24), 
        .A(n4525), .ZN(n4539) );
  AOI22_X1 U5041 ( .A1(n4530), .A2(keyinput3), .B1(n4529), .B2(keyinput8), 
        .ZN(n4528) );
  OAI221_X1 U5042 ( .B1(n4530), .B2(keyinput3), .C1(n4529), .C2(keyinput8), 
        .A(n4528), .ZN(n4538) );
  AOI22_X1 U5043 ( .A1(n4533), .A2(keyinput28), .B1(keyinput2), .B2(n4532), 
        .ZN(n4531) );
  OAI221_X1 U5044 ( .B1(n4533), .B2(keyinput28), .C1(n4532), .C2(keyinput2), 
        .A(n4531), .ZN(n4537) );
  AOI22_X1 U5045 ( .A1(n4578), .A2(keyinput37), .B1(n4535), .B2(keyinput52), 
        .ZN(n4534) );
  OAI221_X1 U5046 ( .B1(n4578), .B2(keyinput37), .C1(n4535), .C2(keyinput52), 
        .A(n4534), .ZN(n4536) );
  NOR4_X1 U5047 ( .A1(n4539), .A2(n4538), .A3(n4537), .A4(n4536), .ZN(n4540)
         );
  NAND4_X1 U5048 ( .A1(n4543), .A2(n4542), .A3(n4541), .A4(n4540), .ZN(n4544)
         );
  NOR3_X1 U5049 ( .A1(n4546), .A2(n4545), .A3(n4544), .ZN(n4557) );
  AOI22_X1 U5050 ( .A1(n4548), .A2(keyinput1), .B1(n4561), .B2(keyinput40), 
        .ZN(n4547) );
  OAI221_X1 U5051 ( .B1(n4548), .B2(keyinput1), .C1(n4561), .C2(keyinput40), 
        .A(n4547), .ZN(n4555) );
  INV_X1 U5052 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4560) );
  AOI22_X1 U5053 ( .A1(n2273), .A2(keyinput20), .B1(n4560), .B2(keyinput60), 
        .ZN(n4549) );
  OAI221_X1 U5054 ( .B1(n2273), .B2(keyinput20), .C1(n4560), .C2(keyinput60), 
        .A(n4549), .ZN(n4554) );
  AOI22_X1 U5055 ( .A1(n2489), .A2(keyinput63), .B1(keyinput62), .B2(n3296), 
        .ZN(n4550) );
  OAI221_X1 U5056 ( .B1(n2489), .B2(keyinput63), .C1(n3296), .C2(keyinput62), 
        .A(n4550), .ZN(n4553) );
  AOI22_X1 U5057 ( .A1(n2528), .A2(keyinput19), .B1(keyinput58), .B2(n3669), 
        .ZN(n4551) );
  OAI221_X1 U5058 ( .B1(n2528), .B2(keyinput19), .C1(n3669), .C2(keyinput58), 
        .A(n4551), .ZN(n4552) );
  NOR4_X1 U5059 ( .A1(n4555), .A2(n4554), .A3(n4553), .A4(n4552), .ZN(n4556)
         );
  NAND3_X1 U5060 ( .A1(n4558), .A2(n4557), .A3(n4556), .ZN(n4595) );
  INV_X1 U5061 ( .A(n4559), .ZN(n4593) );
  NOR4_X1 U5062 ( .A1(REG1_REG_8__SCAN_IN), .A2(REG2_REG_3__SCAN_IN), .A3(
        n4561), .A4(n4560), .ZN(n4587) );
  NAND4_X1 U5063 ( .A1(REG2_REG_23__SCAN_IN), .A2(n2528), .A3(n3296), .A4(
        n3669), .ZN(n4568) );
  NAND4_X1 U5064 ( .A1(REG0_REG_4__SCAN_IN), .A2(n4564), .A3(n4563), .A4(n4562), .ZN(n4567) );
  NAND3_X1 U5065 ( .A1(REG0_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .A3(
        n4565), .ZN(n4566) );
  NOR4_X1 U5066 ( .A1(DATAO_REG_31__SCAN_IN), .A2(n4568), .A3(n4567), .A4(
        n4566), .ZN(n4586) );
  NAND3_X1 U5067 ( .A1(ADDR_REG_15__SCAN_IN), .A2(DATAO_REG_7__SCAN_IN), .A3(
        DATAO_REG_14__SCAN_IN), .ZN(n4573) );
  NAND4_X1 U5068 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_5__SCAN_IN), .A3(
        DATAO_REG_0__SCAN_IN), .A4(n2412), .ZN(n4572) );
  NOR3_X1 U5069 ( .A1(REG3_REG_11__SCAN_IN), .A2(DATAO_REG_22__SCAN_IN), .A3(
        DATAO_REG_26__SCAN_IN), .ZN(n4570) );
  NOR3_X1 U5070 ( .A1(REG3_REG_6__SCAN_IN), .A2(ADDR_REG_7__SCAN_IN), .A3(
        ADDR_REG_3__SCAN_IN), .ZN(n4569) );
  NAND4_X1 U5071 ( .A1(REG3_REG_22__SCAN_IN), .A2(ADDR_REG_10__SCAN_IN), .A3(
        n4570), .A4(n4569), .ZN(n4571) );
  NOR4_X1 U5072 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4573), .A3(n4572), .A4(n4571), 
        .ZN(n4585) );
  NAND4_X1 U5073 ( .A1(DATAI_16_), .A2(REG3_REG_13__SCAN_IN), .A3(n4575), .A4(
        n4574), .ZN(n4583) );
  NAND4_X1 U5074 ( .A1(REG3_REG_27__SCAN_IN), .A2(DATAI_18_), .A3(n4577), .A4(
        n4576), .ZN(n4582) );
  NAND4_X1 U5075 ( .A1(D_REG_22__SCAN_IN), .A2(REG0_REG_3__SCAN_IN), .A3(n4579), .A4(n4578), .ZN(n4581) );
  NAND4_X1 U5076 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_31__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(IR_REG_29__SCAN_IN), .ZN(n4580) );
  NOR4_X1 U5077 ( .A1(n4583), .A2(n4582), .A3(n4581), .A4(n4580), .ZN(n4584)
         );
  NAND4_X1 U5078 ( .A1(n4587), .A2(n4586), .A3(n4585), .A4(n4584), .ZN(n4592)
         );
  NAND4_X1 U5079 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .A3(
        REG1_REG_11__SCAN_IN), .A4(REG1_REG_2__SCAN_IN), .ZN(n4588) );
  OR4_X1 U5080 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .A3(
        IR_REG_12__SCAN_IN), .A4(n4588), .ZN(n4591) );
  NAND4_X1 U5081 ( .A1(n4589), .A2(IR_REG_2__SCAN_IN), .A3(IR_REG_13__SCAN_IN), 
        .A4(IR_REG_0__SCAN_IN), .ZN(n4590) );
  NOR4_X1 U5082 ( .A1(n4593), .A2(n4592), .A3(n4591), .A4(n4590), .ZN(n4594)
         );
  XNOR2_X1 U5083 ( .A(n4595), .B(n4594), .ZN(n4596) );
  XNOR2_X1 U5084 ( .A(n4597), .B(n4596), .ZN(U3254) );
endmodule

