

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9694, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
         n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
         n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
         n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
         n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
         n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036,
         n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
         n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
         n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
         n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
         n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
         n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
         n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
         n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
         n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156,
         n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
         n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
         n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
         n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
         n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
         n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204,
         n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
         n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220,
         n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228,
         n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
         n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
         n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252,
         n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260,
         n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268,
         n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
         n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
         n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292,
         n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300,
         n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308,
         n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
         n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324,
         n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332,
         n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340,
         n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348,
         n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356,
         n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364,
         n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372,
         n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380,
         n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388,
         n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396,
         n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404,
         n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412,
         n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420,
         n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428,
         n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436,
         n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444,
         n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452,
         n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460,
         n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468,
         n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476,
         n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484,
         n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492,
         n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500,
         n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508,
         n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516,
         n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524,
         n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532,
         n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540,
         n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548,
         n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556,
         n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564,
         n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572,
         n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580,
         n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588,
         n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596,
         n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
         n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612,
         n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620,
         n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
         n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636,
         n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644,
         n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652,
         n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660,
         n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668,
         n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
         n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684,
         n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692,
         n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700,
         n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708,
         n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716,
         n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724,
         n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732,
         n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740,
         n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748,
         n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756,
         n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764,
         n21765, n21766, n21767, n21768, n21769, n21770;

  INV_X1 U11127 ( .A(n21089), .ZN(n21040) );
  INV_X1 U11128 ( .A(n21086), .ZN(n21041) );
  NOR2_X1 U11129 ( .A1(n17565), .A2(n10299), .ZN(n17551) );
  INV_X1 U11130 ( .A(n15899), .ZN(n15889) );
  AND2_X1 U11131 ( .A1(n17109), .A2(n11086), .ZN(n10203) );
  OAI21_X2 U11132 ( .B1(n17140), .B2(n17141), .A(n10226), .ZN(n17132) );
  OAI21_X1 U11133 ( .B1(n9687), .B2(n10215), .A(n10214), .ZN(n17080) );
  NAND2_X1 U11134 ( .A1(n10415), .A2(n9722), .ZN(n16753) );
  NAND4_X2 U11135 ( .A1(n10200), .A2(n9925), .A3(n9924), .A4(n10841), .ZN(
        n11084) );
  CLKBUF_X1 U11136 ( .A(n12214), .Z(n17446) );
  NAND2_X1 U11137 ( .A1(n15187), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15191) );
  NAND2_X1 U11138 ( .A1(n12227), .A2(n12226), .ZN(n12229) );
  NOR2_X2 U11139 ( .A1(n10048), .A2(n14582), .ZN(n10792) );
  INV_X1 U11140 ( .A(n10781), .ZN(n17183) );
  NAND4_X1 U11141 ( .A1(n10871), .A2(n10870), .A3(n10869), .A4(n10868), .ZN(
        n11477) );
  BUF_X2 U11142 ( .A(n11207), .Z(n11473) );
  CLKBUF_X2 U11143 ( .A(n12611), .Z(n9705) );
  CLKBUF_X2 U11144 ( .A(n12610), .Z(n15355) );
  CLKBUF_X2 U11145 ( .A(n12605), .Z(n15197) );
  CLKBUF_X2 U11146 ( .A(n12589), .Z(n15360) );
  AND2_X1 U11147 ( .A1(n15772), .A2(n13126), .ZN(n10087) );
  CLKBUF_X2 U11148 ( .A(n15302), .Z(n9694) );
  INV_X1 U11149 ( .A(n9756), .ZN(n18551) );
  OR2_X1 U11150 ( .A1(n12635), .A2(n12634), .ZN(n13766) );
  INV_X1 U11151 ( .A(n14449), .ZN(n15394) );
  INV_X4 U11152 ( .A(n18464), .ZN(n18472) );
  CLKBUF_X2 U11153 ( .A(n17765), .Z(n18545) );
  NAND2_X1 U11154 ( .A1(n20964), .A2(n20968), .ZN(n15442) );
  OR2_X1 U11155 ( .A1(n12576), .A2(n12575), .ZN(n14464) );
  CLKBUF_X1 U11156 ( .A(n12626), .Z(n14460) );
  INV_X1 U11157 ( .A(n12012), .ZN(n17682) );
  CLKBUF_X1 U11160 ( .A(n13345), .Z(n18517) );
  AND4_X1 U11161 ( .A1(n12557), .A2(n12556), .A3(n12555), .A4(n12554), .ZN(
        n12564) );
  INV_X1 U11162 ( .A(n9746), .ZN(n18477) );
  INV_X1 U11163 ( .A(n10712), .ZN(n9921) );
  AND2_X2 U11164 ( .A1(n14287), .A2(n12518), .ZN(n9704) );
  AND2_X1 U11165 ( .A1(n12520), .A2(n12519), .ZN(n12589) );
  AND2_X2 U11166 ( .A1(n12517), .A2(n14290), .ZN(n12536) );
  NAND2_X2 U11167 ( .A1(n13529), .A2(n11672), .ZN(n9756) );
  CLKBUF_X1 U11168 ( .A(n19606), .Z(n9683) );
  NOR2_X1 U11169 ( .A1(n19864), .A2(n19589), .ZN(n19606) );
  CLKBUF_X1 U11170 ( .A(n19849), .Z(n9684) );
  NOR2_X1 U11171 ( .A1(n19864), .A2(n19735), .ZN(n19849) );
  INV_X1 U11172 ( .A(n15442), .ZN(n9692) );
  AND2_X2 U11173 ( .A1(n14287), .A2(n12518), .ZN(n12581) );
  OR2_X1 U11174 ( .A1(n14464), .A2(n21641), .ZN(n15329) );
  AND2_X1 U11175 ( .A1(n14290), .A2(n12518), .ZN(n12687) );
  AND4_X1 U11176 ( .A1(n12515), .A2(n12514), .A3(n12513), .A4(n12512), .ZN(
        n12526) );
  NOR2_X1 U11177 ( .A1(n10770), .A2(n17183), .ZN(n10812) );
  INV_X2 U11178 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14353) );
  INV_X1 U11179 ( .A(n9756), .ZN(n17784) );
  NAND2_X1 U11181 ( .A1(n12594), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12602) );
  INV_X1 U11182 ( .A(n15329), .ZN(n15379) );
  INV_X1 U11184 ( .A(n11361), .ZN(n11512) );
  NOR2_X1 U11185 ( .A1(n15434), .A2(n11482), .ZN(n11484) );
  INV_X1 U11186 ( .A(n11091), .ZN(n11558) );
  INV_X1 U11187 ( .A(n11477), .ZN(n11482) );
  NAND2_X1 U11188 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13537) );
  AND4_X1 U11189 ( .A1(n12621), .A2(n12620), .A3(n12619), .A4(n12618), .ZN(
        n12622) );
  NAND2_X1 U11190 ( .A1(n15626), .A2(n10039), .ZN(n15595) );
  NAND2_X1 U11191 ( .A1(n15823), .A2(n12695), .ZN(n12588) );
  XNOR2_X1 U11193 ( .A(n11484), .B(n11483), .ZN(n11485) );
  AOI211_X1 U11194 ( .C1(n14919), .C2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14918), .B(n14917), .ZN(n14920) );
  INV_X1 U11195 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n17491) );
  INV_X1 U11196 ( .A(n18432), .ZN(n18408) );
  INV_X1 U11197 ( .A(n19443), .ZN(n13546) );
  NAND2_X1 U11198 ( .A1(n18032), .A2(n20046), .ZN(n14235) );
  NOR2_X1 U11199 ( .A1(n18987), .A2(n18973), .ZN(n18968) );
  INV_X1 U11200 ( .A(n15775), .ZN(n21036) );
  NAND2_X1 U11201 ( .A1(n15479), .A2(n15465), .ZN(n15447) );
  NOR2_X1 U11202 ( .A1(n10187), .A2(n14862), .ZN(n16966) );
  OAI21_X1 U11203 ( .B1(n20540), .B2(n20539), .A(n20538), .ZN(n20558) );
  INV_X1 U11204 ( .A(n20031), .ZN(n19420) );
  NAND2_X1 U11205 ( .A1(n13546), .A2(n19440), .ZN(n13433) );
  NAND2_X1 U11206 ( .A1(n19289), .A2(n19306), .ZN(n19318) );
  OR2_X1 U11207 ( .A1(n15453), .A2(n15451), .ZN(n15775) );
  INV_X1 U11208 ( .A(n20346), .ZN(n20355) );
  NAND2_X1 U11209 ( .A1(n19870), .A2(n20038), .ZN(n18041) );
  AOI211_X1 U11210 ( .C1(n18087), .C2(n18453), .A(n18078), .B(n18077), .ZN(
        n18079) );
  AND2_X1 U11211 ( .A1(n13912), .A2(n9809), .ZN(n9685) );
  AND2_X2 U11212 ( .A1(n14287), .A2(n12520), .ZN(n12611) );
  AND2_X1 U11214 ( .A1(n12518), .A2(n10275), .ZN(n9686) );
  AND2_X4 U11215 ( .A1(n12518), .A2(n10275), .ZN(n12594) );
  AND2_X1 U11216 ( .A1(n12517), .A2(n12519), .ZN(n9699) );
  NAND2_X2 U11217 ( .A1(n13687), .A2(n13686), .ZN(n13688) );
  OAI21_X1 U11218 ( .B1(n16691), .B2(n12435), .A(n12434), .ZN(n12457) );
  NAND2_X2 U11220 ( .A1(n11415), .A2(n12192), .ZN(n14828) );
  XNOR2_X2 U11221 ( .A(n13519), .B(n12795), .ZN(n13583) );
  INV_X2 U11222 ( .A(n11084), .ZN(n9942) );
  AND2_X4 U11223 ( .A1(n11683), .A2(n10249), .ZN(n13472) );
  BUF_X2 U11224 ( .A(n11077), .Z(n9687) );
  NAND2_X2 U11225 ( .A1(n14442), .A2(n12729), .ZN(n12732) );
  XNOR2_X2 U11226 ( .A(n13118), .B(n13117), .ZN(n15388) );
  NAND2_X1 U11227 ( .A1(n12867), .A2(n12866), .ZN(n9688) );
  NAND2_X1 U11228 ( .A1(n12867), .A2(n12866), .ZN(n9689) );
  NAND2_X4 U11229 ( .A1(n12867), .A2(n12866), .ZN(n12890) );
  INV_X4 U11230 ( .A(n12890), .ZN(n16103) );
  OAI211_X2 U11231 ( .C1(n19052), .C2(n9981), .A(n9978), .B(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19043) );
  NAND2_X2 U11232 ( .A1(n12788), .A2(n12787), .ZN(n13519) );
  XNOR2_X1 U11233 ( .A(n12090), .B(n12089), .ZN(n12092) );
  OAI21_X2 U11234 ( .B1(n16710), .B2(n12365), .A(n12364), .ZN(n16705) );
  NAND2_X2 U11235 ( .A1(n16759), .A2(n10121), .ZN(n16710) );
  NOR2_X2 U11236 ( .A1(n18258), .A2(n13721), .ZN(n13890) );
  NOR2_X2 U11237 ( .A1(n14574), .A2(n18954), .ZN(n18971) );
  AOI211_X2 U11238 ( .C1(n11202), .C2(n11389), .A(n11201), .B(n11200), .ZN(
        n11203) );
  NAND2_X2 U11239 ( .A1(n10020), .A2(n10201), .ZN(n17032) );
  NAND2_X1 U11240 ( .A1(n9902), .A2(n10463), .ZN(n16675) );
  OAI21_X1 U11241 ( .B1(n11422), .B2(n10223), .A(n10222), .ZN(n16957) );
  AND2_X1 U11242 ( .A1(n17550), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10297) );
  XNOR2_X1 U11244 ( .A(n11084), .B(n11085), .ZN(n11077) );
  NAND2_X1 U11245 ( .A1(n18816), .A2(n18966), .ZN(n18821) );
  OR2_X1 U11246 ( .A1(n17370), .A2(n11562), .ZN(n17253) );
  NOR2_X1 U11247 ( .A1(n21581), .A2(n21451), .ZN(n21632) );
  NAND2_X1 U11248 ( .A1(n12802), .A2(n12811), .ZN(n21743) );
  NAND2_X1 U11249 ( .A1(n17383), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17370) );
  NOR2_X1 U11250 ( .A1(n17433), .A2(n11407), .ZN(n17406) );
  AND2_X1 U11251 ( .A1(n10285), .A2(n10284), .ZN(n18124) );
  NAND2_X1 U11252 ( .A1(n12112), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18951) );
  NAND2_X4 U11253 ( .A1(n14828), .A2(n11399), .ZN(n10181) );
  INV_X1 U11254 ( .A(n21082), .ZN(n21068) );
  INV_X2 U11255 ( .A(n17455), .ZN(n10780) );
  NAND2_X1 U11256 ( .A1(n10762), .A2(n10763), .ZN(n10782) );
  INV_X1 U11257 ( .A(n10044), .ZN(n10042) );
  AND2_X1 U11258 ( .A1(n14235), .A2(n9808), .ZN(n13373) );
  CLKBUF_X1 U11259 ( .A(n11195), .Z(n14404) );
  INV_X1 U11260 ( .A(n12940), .ZN(n12948) );
  INV_X4 U11261 ( .A(n13223), .ZN(n16694) );
  INV_X1 U11262 ( .A(n18681), .ZN(n10081) );
  AND3_X1 U11263 ( .A1(n9990), .A2(n9989), .A3(n9726), .ZN(n11390) );
  NAND3_X1 U11264 ( .A1(n12004), .A2(n12002), .A3(n12003), .ZN(n19448) );
  NAND2_X1 U11265 ( .A1(n9920), .A2(n9919), .ZN(n11382) );
  NAND2_X1 U11266 ( .A1(n10494), .A2(n10495), .ZN(n11219) );
  AND4_X1 U11267 ( .A1(n12604), .A2(n12603), .A3(n12602), .A4(n12601), .ZN(
        n12625) );
  INV_X8 U11268 ( .A(n17799), .ZN(n17774) );
  INV_X1 U11269 ( .A(n18539), .ZN(n11716) );
  INV_X8 U11270 ( .A(n17769), .ZN(n18552) );
  BUF_X2 U11271 ( .A(n12665), .Z(n15254) );
  CLKBUF_X2 U11272 ( .A(n12536), .Z(n15202) );
  CLKBUF_X2 U11274 ( .A(n12717), .Z(n15361) );
  CLKBUF_X2 U11275 ( .A(n12696), .Z(n15341) );
  INV_X4 U11276 ( .A(n18541), .ZN(n18524) );
  INV_X4 U11277 ( .A(n17767), .ZN(n9690) );
  INV_X1 U11278 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13539) );
  NAND2_X1 U11279 ( .A1(n10127), .A2(n10210), .ZN(n10209) );
  XNOR2_X1 U11280 ( .A(n10151), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17622) );
  NOR2_X1 U11281 ( .A1(n16675), .A2(n16650), .ZN(n16672) );
  NAND2_X1 U11282 ( .A1(n10367), .A2(n10365), .ZN(n15418) );
  OR2_X1 U11283 ( .A1(n15447), .A2(n10369), .ZN(n10365) );
  XNOR2_X1 U11284 ( .A(n10280), .B(n15920), .ZN(n16154) );
  OR2_X1 U11285 ( .A1(n17551), .A2(n17550), .ZN(n10151) );
  NAND2_X1 U11286 ( .A1(n10464), .A2(n10465), .ZN(n10463) );
  OAI21_X1 U11287 ( .B1(n10282), .B2(n9761), .A(n10281), .ZN(n10280) );
  AOI21_X1 U11288 ( .B1(n10038), .B2(n15567), .A(n10034), .ZN(n10033) );
  NAND2_X1 U11289 ( .A1(n10282), .A2(n15919), .ZN(n10281) );
  AND2_X1 U11290 ( .A1(n15270), .A2(n9817), .ZN(n15479) );
  OR2_X1 U11291 ( .A1(n10297), .A2(n10073), .ZN(n10072) );
  OR2_X1 U11292 ( .A1(n16084), .A2(n16083), .ZN(n16081) );
  INV_X1 U11293 ( .A(n15967), .ZN(n15956) );
  NAND2_X1 U11294 ( .A1(n9800), .A2(n15741), .ZN(n21011) );
  NAND2_X1 U11295 ( .A1(n9747), .A2(n15698), .ZN(n15699) );
  AND2_X1 U11296 ( .A1(n12889), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9884) );
  AOI21_X1 U11297 ( .B1(n15975), .B2(n12885), .A(n12884), .ZN(n12888) );
  CLKBUF_X1 U11298 ( .A(n15918), .Z(n15967) );
  AND2_X1 U11299 ( .A1(n16144), .A2(n16143), .ZN(n9997) );
  NOR2_X1 U11300 ( .A1(n9769), .A2(n11478), .ZN(n11479) );
  NOR2_X1 U11301 ( .A1(n10301), .A2(n10300), .ZN(n17582) );
  AND2_X1 U11302 ( .A1(n17046), .A2(n9804), .ZN(n10544) );
  AND2_X1 U11303 ( .A1(n10512), .A2(n10140), .ZN(n10229) );
  AND2_X1 U11304 ( .A1(n10006), .A2(n10162), .ZN(n9880) );
  NOR2_X1 U11305 ( .A1(n15468), .A2(n13114), .ZN(n13115) );
  INV_X1 U11306 ( .A(n14646), .ZN(n10358) );
  AND2_X1 U11307 ( .A1(n11466), .A2(n11465), .ZN(n16429) );
  OAI221_X1 U11308 ( .B1(n10557), .B2(n21530), .C1(n10557), .C2(n21339), .A(
        n21529), .ZN(n21358) );
  OAI22_X1 U11309 ( .A1(n21535), .A2(n21534), .B1(n21533), .B2(n21532), .ZN(
        n21565) );
  OAI211_X1 U11310 ( .C1(n10556), .C2(n21530), .A(n21529), .B(n21528), .ZN(
        n21566) );
  INV_X1 U11311 ( .A(n10279), .ZN(n10095) );
  NAND3_X1 U11312 ( .A1(n10842), .A2(n10449), .A3(n11073), .ZN(n17177) );
  INV_X1 U11313 ( .A(n20592), .ZN(n20584) );
  NAND2_X1 U11314 ( .A1(n10200), .A2(n10841), .ZN(n11073) );
  OAI211_X1 U11315 ( .C1(n21401), .C2(n21400), .A(n21463), .B(n21399), .ZN(
        n21419) );
  INV_X2 U11316 ( .A(n17509), .ZN(n20821) );
  AND2_X1 U11317 ( .A1(n19031), .A2(n10157), .ZN(n18847) );
  NAND2_X1 U11318 ( .A1(n10517), .A2(n10516), .ZN(n10515) );
  NAND2_X1 U11319 ( .A1(n10839), .A2(n10840), .ZN(n10842) );
  INV_X2 U11320 ( .A(n17507), .ZN(n20747) );
  NOR2_X1 U11321 ( .A1(n17863), .A2(n10228), .ZN(n10227) );
  AOI211_X1 U11322 ( .C1(n18111), .C2(n18108), .A(n18107), .B(n18106), .ZN(
        n18109) );
  CLKBUF_X1 U11323 ( .A(n11464), .Z(n11481) );
  NOR2_X1 U11324 ( .A1(n16141), .A2(n10266), .ZN(n16130) );
  NAND2_X1 U11325 ( .A1(n20533), .A2(n20564), .ZN(n20592) );
  AND2_X1 U11326 ( .A1(n10356), .A2(n14761), .ZN(n10133) );
  OAI211_X1 U11327 ( .C1(n16367), .C2(n16364), .A(n21529), .B(n21461), .ZN(
        n16389) );
  OAI21_X1 U11328 ( .B1(n12861), .B2(n10164), .A(n12872), .ZN(n10163) );
  AND2_X1 U11329 ( .A1(n14654), .A2(n10357), .ZN(n10356) );
  NAND2_X1 U11330 ( .A1(n9930), .A2(n10838), .ZN(n10840) );
  NAND2_X1 U11331 ( .A1(n9881), .A2(n12800), .ZN(n14535) );
  NOR2_X2 U11332 ( .A1(n20629), .A2(n20628), .ZN(n20684) );
  NOR2_X2 U11333 ( .A1(n20562), .A2(n20500), .ZN(n20383) );
  OR2_X1 U11334 ( .A1(n12860), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12861) );
  NAND2_X1 U11335 ( .A1(n19280), .A2(n10157), .ZN(n19230) );
  OR2_X1 U11336 ( .A1(n16533), .A2(n11482), .ZN(n11021) );
  OAI21_X1 U11337 ( .B1(n10193), .B2(n10167), .A(n12805), .ZN(n14599) );
  NAND2_X1 U11338 ( .A1(n21743), .A2(n10031), .ZN(n21293) );
  NAND2_X1 U11339 ( .A1(n12772), .A2(n12771), .ZN(n14601) );
  NOR2_X1 U11340 ( .A1(n21743), .A2(n14659), .ZN(n21494) );
  AOI21_X1 U11341 ( .B1(n14751), .B2(n15043), .A(n14750), .ZN(n14769) );
  OR2_X1 U11342 ( .A1(n9688), .A2(n16279), .ZN(n16055) );
  AND2_X1 U11343 ( .A1(n12824), .A2(n12846), .ZN(n10511) );
  AND2_X1 U11344 ( .A1(n18919), .A2(n11854), .ZN(n18915) );
  XNOR2_X1 U11345 ( .A(n12799), .B(n12995), .ZN(n13795) );
  NOR2_X1 U11346 ( .A1(n16201), .A2(n10255), .ZN(n16192) );
  OR2_X1 U11347 ( .A1(n16194), .A2(n16182), .ZN(n16174) );
  NOR2_X1 U11348 ( .A1(n15570), .A2(n15571), .ZN(n13088) );
  AND2_X1 U11349 ( .A1(n17406), .A2(n11405), .ZN(n17383) );
  XNOR2_X1 U11350 ( .A(n12867), .B(n12853), .ZN(n14752) );
  NAND2_X1 U11351 ( .A1(n12798), .A2(n12797), .ZN(n12799) );
  AND2_X1 U11352 ( .A1(n13895), .A2(n13774), .ZN(n12244) );
  NOR2_X1 U11353 ( .A1(n18124), .A2(n18339), .ZN(n18113) );
  AND2_X1 U11354 ( .A1(n10256), .A2(n17892), .ZN(n16201) );
  INV_X1 U11356 ( .A(n15650), .ZN(n13073) );
  OR2_X1 U11357 ( .A1(n16234), .A2(n10257), .ZN(n10256) );
  AND2_X1 U11358 ( .A1(n10784), .A2(n10056), .ZN(n20291) );
  NOR2_X1 U11359 ( .A1(n16223), .A2(n16224), .ZN(n16210) );
  NAND2_X1 U11360 ( .A1(n17440), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17433) );
  NAND2_X1 U11361 ( .A1(n13066), .A2(n13065), .ZN(n15650) );
  OR2_X1 U11362 ( .A1(n13155), .A2(n16240), .ZN(n16234) );
  AND2_X1 U11363 ( .A1(n10775), .A2(n14582), .ZN(n20622) );
  AND2_X2 U11364 ( .A1(n10773), .A2(n14582), .ZN(n10910) );
  AND2_X1 U11365 ( .A1(n10775), .A2(n17183), .ZN(n10820) );
  AND2_X1 U11366 ( .A1(n10773), .A2(n17183), .ZN(n20689) );
  INV_X1 U11367 ( .A(n19116), .ZN(n19096) );
  AND2_X1 U11368 ( .A1(n10181), .A2(n10180), .ZN(n17440) );
  AND2_X1 U11369 ( .A1(n10788), .A2(n17183), .ZN(n10789) );
  CLKBUF_X1 U11370 ( .A(n15825), .Z(n15875) );
  OR2_X1 U11371 ( .A1(n11009), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11013) );
  AND2_X1 U11372 ( .A1(n12214), .A2(n9719), .ZN(n10775) );
  OR2_X1 U11373 ( .A1(n12214), .A2(n10771), .ZN(n10770) );
  XNOR2_X1 U11374 ( .A(n12680), .B(n12679), .ZN(n12775) );
  AND2_X1 U11375 ( .A1(n13151), .A2(n13150), .ZN(n16296) );
  AND2_X1 U11376 ( .A1(n12214), .A2(n10772), .ZN(n10773) );
  NAND2_X1 U11377 ( .A1(n17886), .A2(n16297), .ZN(n16259) );
  AND2_X1 U11378 ( .A1(n13166), .A2(n13165), .ZN(n16219) );
  AND2_X1 U11379 ( .A1(n14582), .A2(n16635), .ZN(n10783) );
  AOI21_X1 U11380 ( .B1(n10198), .B2(n21638), .A(n9767), .ZN(n13680) );
  INV_X1 U11381 ( .A(n12214), .ZN(n9691) );
  NOR2_X1 U11382 ( .A1(n21189), .A2(n14468), .ZN(n21603) );
  NOR2_X1 U11383 ( .A1(n21189), .A2(n14459), .ZN(n21597) );
  NAND2_X1 U11384 ( .A1(n11099), .A2(n9987), .ZN(n9986) );
  NOR2_X1 U11385 ( .A1(n21189), .A2(n14473), .ZN(n21591) );
  NOR2_X1 U11386 ( .A1(n21189), .A2(n14445), .ZN(n21577) );
  NAND2_X1 U11387 ( .A1(n13146), .A2(n13754), .ZN(n16297) );
  AND2_X1 U11388 ( .A1(n13146), .A2(n13140), .ZN(n13164) );
  AND2_X1 U11389 ( .A1(n13146), .A2(n13751), .ZN(n21180) );
  NOR2_X1 U11390 ( .A1(n21189), .A2(n14561), .ZN(n21609) );
  CLKBUF_X1 U11391 ( .A(n14505), .Z(n21453) );
  NAND2_X1 U11392 ( .A1(n15088), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15226) );
  NOR2_X2 U11393 ( .A1(n20226), .A2(n13780), .ZN(n12194) );
  OR2_X1 U11394 ( .A1(n12733), .A2(n12735), .ZN(n12736) );
  NOR2_X1 U11395 ( .A1(n21189), .A2(n14657), .ZN(n21615) );
  NOR2_X1 U11396 ( .A1(n21189), .A2(n14770), .ZN(n21621) );
  NOR2_X1 U11397 ( .A1(n21189), .A2(n14771), .ZN(n21627) );
  XNOR2_X1 U11398 ( .A(n12103), .B(n10106), .ZN(n19056) );
  AND2_X1 U11399 ( .A1(n12976), .A2(n13618), .ZN(n13146) );
  XNOR2_X1 U11400 ( .A(n10782), .B(n10767), .ZN(n16635) );
  NOR2_X2 U11401 ( .A1(n21169), .A2(n12924), .ZN(n21161) );
  NAND2_X1 U11402 ( .A1(n19062), .A2(n12101), .ZN(n12103) );
  NAND2_X1 U11403 ( .A1(n15390), .A2(n15389), .ZN(n21757) );
  AOI21_X1 U11404 ( .B1(n14346), .B2(n12193), .A(n14802), .ZN(n16897) );
  INV_X1 U11405 ( .A(n11837), .ZN(n10155) );
  OR2_X1 U11406 ( .A1(n10763), .A2(n10762), .ZN(n10768) );
  NAND2_X1 U11407 ( .A1(n11242), .A2(n11241), .ZN(n14777) );
  OR2_X1 U11408 ( .A1(n12659), .A2(n12660), .ZN(n12658) );
  OR3_X1 U11409 ( .A1(n13753), .A2(n13297), .A3(n20982), .ZN(n15390) );
  OR3_X2 U11410 ( .A1(n13753), .A2(n17840), .A3(n13521), .ZN(n20989) );
  NAND2_X1 U11411 ( .A1(n10042), .A2(n9961), .ZN(n10746) );
  NAND2_X1 U11412 ( .A1(n10319), .A2(n10318), .ZN(n14410) );
  AND2_X1 U11413 ( .A1(n9944), .A2(n12681), .ZN(n12729) );
  INV_X2 U11414 ( .A(n18590), .ZN(n18586) );
  AND2_X1 U11415 ( .A1(n9943), .A2(n9821), .ZN(n9944) );
  INV_X1 U11416 ( .A(n19049), .ZN(n10156) );
  AND2_X1 U11417 ( .A1(n10262), .A2(n10260), .ZN(n10258) );
  NAND2_X2 U11418 ( .A1(n11842), .A2(n17632), .ZN(n18950) );
  NAND2_X1 U11419 ( .A1(n10003), .A2(n12654), .ZN(n12662) );
  AND2_X1 U11420 ( .A1(n13431), .A2(n13327), .ZN(n18587) );
  NAND2_X1 U11421 ( .A1(n10634), .A2(n10644), .ZN(n10882) );
  AND2_X1 U11422 ( .A1(n13017), .A2(n13016), .ZN(n14773) );
  AND4_X1 U11423 ( .A1(n10743), .A2(n10742), .A3(n10741), .A4(n10740), .ZN(
        n10745) );
  AND2_X1 U11424 ( .A1(n12927), .A2(n12926), .ZN(n12936) );
  AND2_X1 U11425 ( .A1(n13136), .A2(n13142), .ZN(n9876) );
  NAND2_X1 U11426 ( .A1(n10132), .A2(n10131), .ZN(n10634) );
  CLKBUF_X1 U11427 ( .A(n12991), .Z(n12992) );
  XNOR2_X1 U11428 ( .A(n11820), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19107) );
  NAND2_X1 U11429 ( .A1(n12639), .A2(n15772), .ZN(n13136) );
  NAND2_X1 U11430 ( .A1(n10086), .A2(n10088), .ZN(n13121) );
  AND2_X1 U11431 ( .A1(n13619), .A2(n9700), .ZN(n15443) );
  NAND2_X1 U11432 ( .A1(n12994), .A2(n9700), .ZN(n13490) );
  NAND2_X1 U11433 ( .A1(n11823), .A2(n13511), .ZN(n11828) );
  NAND2_X1 U11434 ( .A1(n13610), .A2(n9700), .ZN(n13104) );
  NAND2_X1 U11435 ( .A1(n11819), .A2(n10016), .ZN(n11820) );
  AND2_X1 U11436 ( .A1(n10733), .A2(n11396), .ZN(n11092) );
  AND2_X1 U11437 ( .A1(n10691), .A2(n13389), .ZN(n10692) );
  NAND2_X1 U11438 ( .A1(n12745), .A2(n12744), .ZN(n12959) );
  AND2_X1 U11439 ( .A1(n11186), .A2(n13780), .ZN(n10677) );
  INV_X1 U11440 ( .A(n13035), .ZN(n13060) );
  AND2_X1 U11441 ( .A1(n12743), .A2(n12694), .ZN(n12712) );
  AND2_X1 U11443 ( .A1(n12587), .A2(n10510), .ZN(n10091) );
  NAND2_X1 U11444 ( .A1(n13458), .A2(n12089), .ZN(n10016) );
  OR2_X1 U11445 ( .A1(n12588), .A2(n13035), .ZN(n13736) );
  INV_X1 U11446 ( .A(n13496), .ZN(n13744) );
  AND3_X1 U11447 ( .A1(n11747), .A2(n11746), .A3(n11745), .ZN(n13608) );
  NAND4_X1 U11448 ( .A1(n11943), .A2(n11942), .A3(n11941), .A4(n11940), .ZN(
        n18681) );
  AND3_X1 U11449 ( .A1(n11960), .A2(n11959), .A3(n11958), .ZN(n19426) );
  NAND2_X1 U11450 ( .A1(n10158), .A2(n9766), .ZN(n12089) );
  OR2_X1 U11451 ( .A1(n11731), .A2(n11730), .ZN(n13511) );
  CLKBUF_X3 U11452 ( .A(n9989), .Z(n13223) );
  NAND2_X1 U11453 ( .A1(n9891), .A2(n9888), .ZN(n10837) );
  NAND2_X1 U11454 ( .A1(n9990), .A2(n20298), .ZN(n9988) );
  NOR2_X1 U11455 ( .A1(n13912), .A2(n11219), .ZN(n10721) );
  NAND2_X1 U11456 ( .A1(n9956), .A2(n11220), .ZN(n10876) );
  NAND2_X1 U11457 ( .A1(n15394), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12744) );
  NAND2_X2 U11458 ( .A1(n10107), .A2(n11713), .ZN(n13458) );
  NAND4_X1 U11459 ( .A1(n11923), .A2(n11922), .A3(n11921), .A4(n11920), .ZN(
        n19440) );
  NAND3_X1 U11461 ( .A1(n9717), .A2(n11878), .A3(n9768), .ZN(n19443) );
  OR2_X1 U11462 ( .A1(n10631), .A2(n10630), .ZN(n11062) );
  INV_X1 U11463 ( .A(n11219), .ZN(n11207) );
  CLKBUF_X2 U11464 ( .A(n10712), .Z(n11389) );
  BUF_X2 U11465 ( .A(n11208), .Z(n13780) );
  OR2_X1 U11466 ( .A1(n17495), .A2(n11220), .ZN(n20964) );
  OR2_X1 U11468 ( .A1(n12706), .A2(n12705), .ZN(n12769) );
  NAND4_X1 U11469 ( .A1(n11816), .A2(n11815), .A3(n11814), .A4(n11813), .ZN(
        n13441) );
  INV_X2 U11470 ( .A(U212), .ZN(n17979) );
  OR2_X1 U11471 ( .A1(n12693), .A2(n12692), .ZN(n12862) );
  NAND2_X2 U11472 ( .A1(n10597), .A2(n10596), .ZN(n17495) );
  AND2_X2 U11473 ( .A1(n10708), .A2(n9923), .ZN(n20298) );
  NAND2_X1 U11474 ( .A1(n12545), .A2(n9751), .ZN(n14469) );
  OR2_X2 U11475 ( .A1(n12600), .A2(n12599), .ZN(n14449) );
  NOR2_X2 U11476 ( .A1(n15837), .A2(n16117), .ZN(n14437) );
  NOR2_X1 U11477 ( .A1(n10551), .A2(n12616), .ZN(n12623) );
  AND4_X1 U11478 ( .A1(n12609), .A2(n12608), .A3(n12607), .A4(n12606), .ZN(
        n12624) );
  NAND3_X1 U11479 ( .A1(n10590), .A2(n10549), .A3(n10589), .ZN(n10597) );
  AND4_X1 U11480 ( .A1(n12540), .A2(n12539), .A3(n12538), .A4(n12537), .ZN(
        n12545) );
  AND4_X1 U11481 ( .A1(n12580), .A2(n12579), .A3(n12578), .A4(n12577), .ZN(
        n12586) );
  AND4_X1 U11482 ( .A1(n12553), .A2(n12552), .A3(n12551), .A4(n12550), .ZN(
        n12565) );
  NAND2_X2 U11483 ( .A1(n19996), .A2(n19943), .ZN(n19999) );
  AND2_X1 U11484 ( .A1(n10587), .A2(n10586), .ZN(n10590) );
  NAND4_X1 U11485 ( .A1(n10595), .A2(n10594), .A3(n10593), .A4(n10592), .ZN(
        n10596) );
  AND4_X1 U11486 ( .A1(n12530), .A2(n12529), .A3(n12528), .A4(n12527), .ZN(
        n10566) );
  AND4_X1 U11487 ( .A1(n12549), .A2(n12548), .A3(n12547), .A4(n12546), .ZN(
        n12566) );
  NOR2_X2 U11488 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19635), .ZN(
        n19656) );
  BUF_X2 U11489 ( .A(n15283), .Z(n15354) );
  INV_X2 U11490 ( .A(n19942), .ZN(n20002) );
  AND2_X1 U11491 ( .A1(n10683), .A2(n10682), .ZN(n10684) );
  BUF_X2 U11492 ( .A(n12612), .Z(n15362) );
  AND2_X2 U11493 ( .A1(n12316), .A2(n14353), .ZN(n10802) );
  NAND2_X2 U11495 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20979), .ZN(n20899) );
  NAND2_X2 U11496 ( .A1(n20979), .A2(n20846), .ZN(n20898) );
  BUF_X2 U11497 ( .A(n10606), .Z(n10697) );
  INV_X2 U11498 ( .A(n20026), .ZN(n19996) );
  NAND2_X2 U11499 ( .A1(n18409), .A2(n13539), .ZN(n18539) );
  AND2_X2 U11500 ( .A1(n12325), .A2(n14353), .ZN(n10804) );
  AND2_X1 U11501 ( .A1(n11682), .A2(n11673), .ZN(n13351) );
  AND2_X2 U11502 ( .A1(n12319), .A2(n14353), .ZN(n12355) );
  INV_X2 U11504 ( .A(n18027), .ZN(n18029) );
  BUF_X4 U11506 ( .A(n10606), .Z(n9696) );
  CLKBUF_X1 U11508 ( .A(n10575), .Z(n14354) );
  AND2_X1 U11509 ( .A1(n14012), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11684) );
  AND2_X1 U11510 ( .A1(n13539), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11673) );
  NOR2_X2 U11513 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11683) );
  NOR2_X2 U11514 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13393) );
  CLKBUF_X1 U11516 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n21737) );
  AND2_X2 U11517 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10275) );
  XNOR2_X1 U11518 ( .A(n11836), .B(n11834), .ZN(n19065) );
  NAND2_X1 U11519 ( .A1(n11836), .A2(n11835), .ZN(n11837) );
  NOR2_X2 U11520 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18334), .ZN(n18312) );
  NAND2_X2 U11521 ( .A1(n18830), .A2(n11857), .ZN(n18861) );
  AND2_X1 U11522 ( .A1(n12517), .A2(n12519), .ZN(n15302) );
  AND2_X2 U11523 ( .A1(n12048), .A2(n12047), .ZN(n19306) );
  INV_X4 U11524 ( .A(n21013), .ZN(n9697) );
  INV_X1 U11525 ( .A(n9697), .ZN(n9698) );
  INV_X1 U11526 ( .A(n21013), .ZN(n21094) );
  AOI211_X2 U11527 ( .C1(n16248), .C2(n21041), .A(n15637), .B(n15636), .ZN(
        n15638) );
  NOR2_X2 U11528 ( .A1(n12636), .A2(n15823), .ZN(n13495) );
  NAND3_X1 U11529 ( .A1(n12636), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n14449), 
        .ZN(n12940) );
  INV_X2 U11530 ( .A(n12632), .ZN(n13500) );
  NAND2_X4 U11531 ( .A1(n12526), .A2(n12525), .ZN(n12632) );
  NOR2_X2 U11533 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18118), .ZN(n18102) );
  NOR2_X2 U11534 ( .A1(n18922), .A2(n18926), .ZN(n18908) );
  NOR2_X4 U11535 ( .A1(n12775), .A2(n12774), .ZN(n10502) );
  AND2_X4 U11536 ( .A1(n12510), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14287) );
  NAND2_X1 U11537 ( .A1(n10502), .A2(n12757), .ZN(n12811) );
  INV_X1 U11538 ( .A(n10502), .ZN(n12801) );
  NAND2_X2 U11539 ( .A1(n10502), .A2(n9784), .ZN(n12867) );
  INV_X1 U11540 ( .A(n13060), .ZN(n9700) );
  INV_X2 U11541 ( .A(n13060), .ZN(n9701) );
  AND2_X1 U11542 ( .A1(n12520), .A2(n10275), .ZN(n9702) );
  AND2_X1 U11543 ( .A1(n14287), .A2(n12518), .ZN(n9703) );
  AND2_X2 U11544 ( .A1(n14290), .A2(n12520), .ZN(n9706) );
  AND2_X4 U11545 ( .A1(n14290), .A2(n12520), .ZN(n12617) );
  AND2_X1 U11546 ( .A1(n14287), .A2(n14304), .ZN(n9707) );
  AND2_X1 U11547 ( .A1(n14287), .A2(n14304), .ZN(n12665) );
  NAND2_X2 U11548 ( .A1(n9904), .A2(n9903), .ZN(n12243) );
  NAND2_X1 U11549 ( .A1(n10460), .A2(n14353), .ZN(n9904) );
  NAND2_X1 U11550 ( .A1(n10459), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9903) );
  INV_X1 U11551 ( .A(n17495), .ZN(n13389) );
  AOI21_X1 U11552 ( .B1(n21761), .B2(n12636), .A(n13131), .ZN(n12643) );
  AND2_X1 U11553 ( .A1(n21641), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15378) );
  NAND2_X1 U11554 ( .A1(n11221), .A2(n9989), .ZN(n13916) );
  AND2_X1 U11555 ( .A1(n11219), .A2(n17491), .ZN(n11221) );
  AND4_X1 U11556 ( .A1(n10867), .A2(n10866), .A3(n10865), .A4(n10864), .ZN(
        n10868) );
  AND4_X1 U11557 ( .A1(n10863), .A2(n10862), .A3(n10861), .A4(n10860), .ZN(
        n10869) );
  CLKBUF_X2 U11558 ( .A(n12630), .Z(n15772) );
  NOR2_X1 U11559 ( .A1(n12241), .A2(n12240), .ZN(n12242) );
  OR2_X1 U11560 ( .A1(n12244), .A2(n10559), .ZN(n10126) );
  INV_X1 U11561 ( .A(n13775), .ZN(n12240) );
  NAND2_X1 U11562 ( .A1(n10426), .A2(n10424), .ZN(n10423) );
  NOR2_X1 U11563 ( .A1(n16420), .A2(n12506), .ZN(n10424) );
  AND2_X1 U11564 ( .A1(n9743), .A2(n17202), .ZN(n10186) );
  NAND2_X1 U11565 ( .A1(n17032), .A2(n14875), .ZN(n10187) );
  XNOR2_X1 U11566 ( .A(n12229), .B(n12230), .ZN(n13905) );
  XNOR2_X1 U11567 ( .A(n13775), .B(n13773), .ZN(n13894) );
  INV_X1 U11568 ( .A(n13774), .ZN(n13773) );
  NAND2_X1 U11569 ( .A1(n20324), .A2(n20944), .ZN(n20500) );
  NAND2_X1 U11570 ( .A1(n10267), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10266) );
  NAND2_X1 U11571 ( .A1(n16259), .A2(n13160), .ZN(n10267) );
  NAND2_X1 U11572 ( .A1(n10234), .A2(n10232), .ZN(n10237) );
  NAND2_X1 U11573 ( .A1(n10500), .A2(n10233), .ZN(n10232) );
  INV_X1 U11574 ( .A(n12756), .ZN(n10233) );
  NAND2_X1 U11575 ( .A1(n10504), .A2(n10503), .ZN(n12733) );
  AOI21_X1 U11576 ( .B1(n10506), .B2(n12707), .A(n12865), .ZN(n10503) );
  AOI21_X1 U11577 ( .B1(n12708), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10507), 
        .ZN(n10506) );
  INV_X1 U11578 ( .A(n11382), .ZN(n9990) );
  NAND2_X1 U11579 ( .A1(n11371), .A2(n9779), .ZN(n10450) );
  NAND2_X1 U11580 ( .A1(n10719), .A2(n9777), .ZN(n10451) );
  OAI21_X1 U11581 ( .B1(n10713), .B2(n11207), .A(n11388), .ZN(n10714) );
  INV_X1 U11582 ( .A(n20298), .ZN(n11388) );
  NAND2_X1 U11583 ( .A1(n10659), .A2(n14353), .ZN(n10666) );
  NOR2_X1 U11584 ( .A1(n11828), .A2(n13608), .ZN(n11832) );
  AND2_X1 U11585 ( .A1(n11832), .A2(n12083), .ZN(n11838) );
  NOR2_X1 U11586 ( .A1(n14460), .A2(n14469), .ZN(n13496) );
  NOR2_X1 U11587 ( .A1(n15501), .A2(n15517), .ZN(n10360) );
  NOR2_X1 U11588 ( .A1(n15196), .A2(n10377), .ZN(n10376) );
  INV_X1 U11589 ( .A(n15086), .ZN(n10377) );
  NAND2_X1 U11590 ( .A1(n10358), .A2(n10133), .ZN(n14941) );
  INV_X1 U11591 ( .A(n13878), .ZN(n15565) );
  INV_X1 U11592 ( .A(n10263), .ZN(n10262) );
  OAI21_X1 U11593 ( .B1(n12955), .B2(n9759), .A(n12961), .ZN(n10263) );
  NAND2_X1 U11594 ( .A1(n12960), .A2(n12959), .ZN(n12961) );
  OR2_X1 U11595 ( .A1(n12957), .A2(n10259), .ZN(n10261) );
  OR2_X1 U11596 ( .A1(n9759), .A2(n12956), .ZN(n10259) );
  NAND2_X1 U11597 ( .A1(n10279), .A2(n10513), .ZN(n10140) );
  NAND2_X1 U11598 ( .A1(n10527), .A2(n15719), .ZN(n10526) );
  AND3_X2 U11599 ( .A1(n12643), .A2(n12637), .A3(n13736), .ZN(n13145) );
  AND2_X1 U11600 ( .A1(n10560), .A2(n20298), .ZN(n10717) );
  NAND2_X1 U11602 ( .A1(n10346), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10345) );
  INV_X1 U11603 ( .A(n10347), .ZN(n10346) );
  NOR2_X1 U11604 ( .A1(n10968), .A2(n10967), .ZN(n10975) );
  OR2_X1 U11605 ( .A1(n10932), .A2(n10931), .ZN(n10937) );
  NAND2_X1 U11606 ( .A1(n10880), .A2(n10879), .ZN(n10881) );
  NAND2_X1 U11607 ( .A1(n11473), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10879) );
  INV_X1 U11608 ( .A(n17495), .ZN(n9956) );
  INV_X1 U11610 ( .A(n11586), .ZN(n11153) );
  NAND2_X1 U11611 ( .A1(n10413), .A2(n10412), .ZN(n10411) );
  OR2_X1 U11612 ( .A1(n20080), .A2(n11482), .ZN(n11017) );
  NAND2_X1 U11613 ( .A1(n17080), .A2(n17081), .ZN(n17046) );
  NOR2_X1 U11614 ( .A1(n10899), .A2(n9931), .ZN(n9924) );
  NAND2_X1 U11615 ( .A1(n11075), .A2(n9711), .ZN(n10934) );
  INV_X1 U11616 ( .A(n9988), .ZN(n11386) );
  NAND2_X1 U11617 ( .A1(n10040), .A2(n10041), .ZN(n9957) );
  NAND2_X1 U11618 ( .A1(n12494), .A2(n11382), .ZN(n10040) );
  INV_X1 U11619 ( .A(n9948), .ZN(n9947) );
  OAI211_X1 U11620 ( .C1(n11102), .C2(n16619), .A(n10750), .B(n10749), .ZN(
        n9948) );
  NAND2_X1 U11621 ( .A1(n10188), .A2(n10200), .ZN(n11075) );
  AND2_X1 U11622 ( .A1(n10841), .A2(n11072), .ZN(n10188) );
  NAND2_X1 U11623 ( .A1(n9797), .A2(n10746), .ZN(n9960) );
  NAND2_X2 U11624 ( .A1(n10023), .A2(n10024), .ZN(n11208) );
  AND2_X1 U11625 ( .A1(n12220), .A2(n16694), .ZN(n14249) );
  AND2_X1 U11626 ( .A1(n14582), .A2(n14360), .ZN(n10784) );
  AND2_X1 U11627 ( .A1(n12214), .A2(n10780), .ZN(n10788) );
  NAND2_X1 U11628 ( .A1(n12039), .A2(n12040), .ZN(n12138) );
  NAND2_X1 U11629 ( .A1(n12062), .A2(n12068), .ZN(n12147) );
  NAND2_X1 U11630 ( .A1(n11684), .A2(n10249), .ZN(n17767) );
  NAND2_X1 U11631 ( .A1(n19043), .A2(n11846), .ZN(n12112) );
  AND2_X1 U11632 ( .A1(n11838), .A2(n12081), .ZN(n11842) );
  AND2_X1 U11633 ( .A1(n19431), .A2(n19448), .ZN(n12074) );
  XNOR2_X1 U11634 ( .A(n11838), .B(n12081), .ZN(n11839) );
  NAND3_X1 U11635 ( .A1(n12153), .A2(n9763), .A3(n12074), .ZN(n13367) );
  AND2_X1 U11636 ( .A1(n17854), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13618) );
  OAI211_X1 U11637 ( .C1(n14601), .C2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n14535), .B(n9995), .ZN(n12809) );
  NAND2_X1 U11638 ( .A1(n10030), .A2(n13882), .ZN(n13883) );
  INV_X1 U11639 ( .A(n13612), .ZN(n17840) );
  AOI21_X1 U11640 ( .B1(n16439), .B2(n10322), .A(n16942), .ZN(n16442) );
  NAND2_X1 U11641 ( .A1(n15422), .A2(n11573), .ZN(n11575) );
  NOR2_X1 U11642 ( .A1(n14388), .A2(n14802), .ZN(n11644) );
  AOI21_X1 U11643 ( .B1(n14778), .B2(n10387), .A(n10385), .ZN(n10384) );
  INV_X1 U11644 ( .A(n13980), .ZN(n10385) );
  AND2_X1 U11646 ( .A1(n11515), .A2(n9858), .ZN(n10405) );
  NAND2_X1 U11647 ( .A1(n10209), .A2(n10408), .ZN(n14901) );
  AOI21_X1 U11648 ( .B1(n10060), .B2(n10063), .A(n11438), .ZN(n10059) );
  NAND2_X1 U11649 ( .A1(n14852), .A2(n9755), .ZN(n10058) );
  NAND2_X1 U11650 ( .A1(n10062), .A2(n10065), .ZN(n14824) );
  NAND2_X1 U11651 ( .A1(n10203), .A2(n17104), .ZN(n10020) );
  INV_X1 U11652 ( .A(n16886), .ZN(n11241) );
  INV_X1 U11653 ( .A(n16597), .ZN(n11242) );
  AND2_X1 U11654 ( .A1(n11236), .A2(n11235), .ZN(n16598) );
  NAND2_X1 U11655 ( .A1(n9905), .A2(n12228), .ZN(n13904) );
  OAI21_X1 U11656 ( .B1(n14582), .B2(n12239), .A(n12238), .ZN(n13775) );
  NAND2_X1 U11657 ( .A1(n13894), .A2(n13895), .ZN(n13899) );
  NAND2_X1 U11658 ( .A1(n11181), .A2(n11573), .ZN(n10318) );
  NAND2_X1 U11659 ( .A1(n10171), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10319) );
  NAND2_X1 U11660 ( .A1(n10172), .A2(n10320), .ZN(n10171) );
  NAND2_X1 U11662 ( .A1(n18915), .A2(n9969), .ZN(n18914) );
  AOI21_X1 U11663 ( .B1(n11856), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9969) );
  NOR2_X1 U11664 ( .A1(n19879), .A2(n17632), .ZN(n19263) );
  AND2_X1 U11665 ( .A1(n12033), .A2(n19426), .ZN(n13372) );
  AND2_X1 U11666 ( .A1(n19426), .A2(n19440), .ZN(n12153) );
  NAND2_X1 U11667 ( .A1(n16159), .A2(n9775), .ZN(n16141) );
  NAND2_X1 U11668 ( .A1(n11059), .A2(n14498), .ZN(n13219) );
  NAND2_X1 U11669 ( .A1(n12190), .A2(n12189), .ZN(n14909) );
  OR2_X1 U11670 ( .A1(n12188), .A2(n12187), .ZN(n12190) );
  XNOR2_X1 U11671 ( .A(n11641), .B(n11559), .ZN(n15429) );
  XNOR2_X1 U11672 ( .A(n10190), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16908) );
  INV_X1 U11673 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20947) );
  NOR2_X1 U11674 ( .A1(n12229), .A2(n13915), .ZN(n20944) );
  INV_X1 U11675 ( .A(n19448), .ZN(n18576) );
  OR2_X1 U11676 ( .A1(n12675), .A2(n12674), .ZN(n12677) );
  NAND3_X1 U11677 ( .A1(n10578), .A2(n10577), .A3(n10579), .ZN(n9892) );
  INV_X1 U11678 ( .A(n10576), .ZN(n9893) );
  NAND2_X1 U11679 ( .A1(n10571), .A2(n10569), .ZN(n9890) );
  NAND2_X1 U11680 ( .A1(n10916), .A2(n10914), .ZN(n9926) );
  NAND2_X1 U11681 ( .A1(n20927), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10873) );
  OAI22_X1 U11682 ( .A1(n12052), .A2(n12056), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n14012), .ZN(n12053) );
  AOI21_X1 U11683 ( .B1(n21737), .B2(n12902), .A(n12904), .ZN(n12915) );
  NOR2_X1 U11684 ( .A1(n12903), .A2(n12905), .ZN(n12904) );
  INV_X1 U11685 ( .A(n12906), .ZN(n12903) );
  INV_X1 U11686 ( .A(n10515), .ZN(n10512) );
  OR2_X1 U11687 ( .A1(n12755), .A2(n12754), .ZN(n12804) );
  AND3_X1 U11688 ( .A1(n12728), .A2(n12727), .A3(n12726), .ZN(n12734) );
  INV_X1 U11689 ( .A(n12677), .ZN(n12778) );
  NAND2_X1 U11690 ( .A1(n10003), .A2(n12641), .ZN(n10002) );
  NAND2_X1 U11691 ( .A1(n12655), .A2(n9773), .ZN(n9998) );
  NAND2_X1 U11692 ( .A1(n10874), .A2(n10873), .ZN(n10895) );
  XNOR2_X1 U11693 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10894) );
  AND4_X1 U11695 ( .A1(n10779), .A2(n10778), .A3(n10777), .A4(n10776), .ZN(
        n10787) );
  OR2_X1 U11696 ( .A1(n10796), .A2(n10795), .ZN(n10117) );
  AND2_X1 U11697 ( .A1(n11382), .A2(n20298), .ZN(n9922) );
  INV_X1 U11698 ( .A(n15548), .ZN(n10375) );
  INV_X1 U11699 ( .A(n15375), .ZN(n15348) );
  NAND2_X1 U11700 ( .A1(n10193), .A2(n12805), .ZN(n10191) );
  NAND2_X1 U11701 ( .A1(n10502), .A2(n10237), .ZN(n12846) );
  INV_X1 U11702 ( .A(n15565), .ZN(n15562) );
  AND2_X1 U11703 ( .A1(n10088), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14325) );
  OAI21_X1 U11704 ( .B1(n12890), .B2(n12881), .A(n10545), .ZN(n10279) );
  INV_X1 U11705 ( .A(n15688), .ZN(n13053) );
  NOR2_X1 U11706 ( .A1(n13039), .A2(n16341), .ZN(n10527) );
  INV_X1 U11707 ( .A(n17872), .ZN(n10228) );
  NAND2_X1 U11708 ( .A1(n13011), .A2(n10523), .ZN(n10522) );
  INV_X1 U11709 ( .A(n14773), .ZN(n10523) );
  AND2_X1 U11710 ( .A1(n12630), .A2(n12929), .ZN(n10085) );
  OAI21_X1 U11711 ( .B1(n21765), .B2(n14314), .A(n14313), .ZN(n14448) );
  INV_X1 U11712 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21575) );
  INV_X1 U11713 ( .A(n10713), .ZN(n10710) );
  OR2_X1 U11714 ( .A1(n11041), .A2(n11042), .ZN(n11049) );
  NAND2_X1 U11715 ( .A1(n11013), .A2(n11456), .ZN(n11015) );
  NAND2_X1 U11716 ( .A1(n10979), .A2(n14568), .ZN(n10991) );
  NAND2_X1 U11717 ( .A1(n9886), .A2(n9885), .ZN(n11031) );
  NAND2_X1 U11718 ( .A1(n10876), .A2(n11166), .ZN(n9885) );
  NAND2_X1 U11719 ( .A1(n10725), .A2(n10724), .ZN(n10043) );
  AOI21_X1 U11720 ( .B1(n11412), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10723), 
        .ZN(n10724) );
  AND2_X1 U11721 ( .A1(n20959), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10723) );
  NAND2_X1 U11722 ( .A1(n9848), .A2(n10123), .ZN(n10122) );
  INV_X1 U11723 ( .A(n10125), .ZN(n10123) );
  INV_X1 U11724 ( .A(n16734), .ZN(n10468) );
  NOR2_X1 U11725 ( .A1(n13871), .A2(n10393), .ZN(n10392) );
  INV_X1 U11726 ( .A(n13876), .ZN(n10393) );
  NAND2_X1 U11727 ( .A1(n9956), .A2(n9780), .ZN(n10730) );
  NAND2_X1 U11728 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10344) );
  NOR2_X1 U11729 ( .A1(n17126), .A2(n10352), .ZN(n10351) );
  NOR2_X1 U11730 ( .A1(n14794), .A2(n10427), .ZN(n10426) );
  INV_X1 U11731 ( .A(n14893), .ZN(n10427) );
  INV_X1 U11732 ( .A(n14813), .ZN(n10406) );
  INV_X1 U11733 ( .A(n16424), .ZN(n10407) );
  INV_X1 U11734 ( .A(n9786), .ZN(n10213) );
  NOR2_X1 U11735 ( .A1(n16989), .A2(n9825), .ZN(n10130) );
  NOR2_X1 U11736 ( .A1(n11437), .A2(n11436), .ZN(n10129) );
  AND2_X1 U11737 ( .A1(n14858), .A2(n11432), .ZN(n9901) );
  AND2_X1 U11738 ( .A1(n10396), .A2(n14872), .ZN(n10395) );
  OR2_X1 U11739 ( .A1(n16493), .A2(n11482), .ZN(n11439) );
  NOR2_X1 U11740 ( .A1(n11523), .A2(n10420), .ZN(n10419) );
  INV_X1 U11741 ( .A(n10421), .ZN(n10420) );
  OR2_X1 U11742 ( .A1(n16499), .A2(n11522), .ZN(n11523) );
  AND2_X1 U11743 ( .A1(n11366), .A2(n10397), .ZN(n10396) );
  INV_X1 U11744 ( .A(n16502), .ZN(n10397) );
  INV_X1 U11745 ( .A(n11368), .ZN(n11366) );
  INV_X1 U11746 ( .A(n16534), .ZN(n11367) );
  NAND2_X1 U11747 ( .A1(n9765), .A2(n11477), .ZN(n11029) );
  NOR2_X1 U11748 ( .A1(n16989), .A2(n11437), .ZN(n10444) );
  NAND2_X1 U11749 ( .A1(n11012), .A2(n11435), .ZN(n10067) );
  AND2_X1 U11750 ( .A1(n10402), .A2(n10400), .ZN(n10399) );
  INV_X1 U11751 ( .A(n14846), .ZN(n10400) );
  OR2_X1 U11752 ( .A1(n20089), .A2(n11482), .ZN(n11011) );
  NOR2_X1 U11753 ( .A1(n14624), .A2(n10403), .ZN(n10402) );
  INV_X1 U11754 ( .A(n10561), .ZN(n10403) );
  INV_X1 U11755 ( .A(n11137), .ZN(n10416) );
  INV_X1 U11756 ( .A(n17378), .ZN(n17303) );
  INV_X1 U11757 ( .A(n13870), .ZN(n10391) );
  INV_X1 U11758 ( .A(n11555), .ZN(n11542) );
  AOI21_X1 U11759 ( .B1(n16592), .B2(n11477), .A(n17405), .ZN(n10214) );
  INV_X1 U11760 ( .A(n16592), .ZN(n10215) );
  AND2_X1 U11761 ( .A1(n10480), .A2(n17170), .ZN(n10479) );
  NAND2_X1 U11762 ( .A1(n10482), .A2(n10484), .ZN(n10480) );
  INV_X1 U11763 ( .A(n10482), .ZN(n10477) );
  NOR2_X1 U11764 ( .A1(n10481), .A2(n11482), .ZN(n10476) );
  OR2_X1 U11765 ( .A1(n10810), .A2(n10809), .ZN(n10877) );
  AND2_X1 U11766 ( .A1(n10746), .A2(n10760), .ZN(n10110) );
  AND2_X1 U11767 ( .A1(n9908), .A2(n11097), .ZN(n9987) );
  INV_X1 U11768 ( .A(n10760), .ZN(n9908) );
  CLKBUF_X1 U11769 ( .A(n11186), .Z(n11187) );
  NAND2_X1 U11770 ( .A1(n20951), .A2(n11182), .ZN(n10316) );
  NAND2_X1 U11771 ( .A1(n14410), .A2(n11183), .ZN(n10317) );
  NAND2_X1 U11772 ( .A1(n11415), .A2(n11397), .ZN(n11399) );
  AND2_X1 U11773 ( .A1(n14249), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12230) );
  AND3_X1 U11774 ( .A1(n10714), .A2(n10716), .A3(n10715), .ZN(n10068) );
  AND2_X1 U11775 ( .A1(n14337), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11054) );
  NAND2_X1 U11776 ( .A1(n12318), .A2(n14353), .ZN(n10554) );
  AND2_X1 U11777 ( .A1(n14249), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12221) );
  NAND2_X1 U11778 ( .A1(n9691), .A2(n9719), .ZN(n10774) );
  NAND2_X1 U11779 ( .A1(n10789), .A2(n16635), .ZN(n10947) );
  INV_X1 U11780 ( .A(n19436), .ZN(n13322) );
  AND2_X1 U11781 ( .A1(n11858), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10304) );
  OR2_X1 U11782 ( .A1(n11838), .A2(n11833), .ZN(n11834) );
  NAND3_X1 U11783 ( .A1(n9973), .A2(n11831), .A3(n9971), .ZN(n11836) );
  AND2_X1 U11784 ( .A1(n12031), .A2(n12030), .ZN(n12045) );
  NAND2_X1 U11785 ( .A1(n13362), .A2(n13373), .ZN(n13377) );
  AND2_X1 U11786 ( .A1(n12142), .A2(n12141), .ZN(n13366) );
  INV_X1 U11787 ( .A(n19883), .ZN(n18039) );
  NAND2_X1 U11788 ( .A1(n13617), .A2(n13616), .ZN(n13758) );
  OR2_X1 U11789 ( .A1(n13753), .A2(n13614), .ZN(n13617) );
  AND2_X1 U11790 ( .A1(n13613), .A2(n13742), .ZN(n13614) );
  NAND2_X1 U11791 ( .A1(n10370), .A2(n15380), .ZN(n10369) );
  INV_X1 U11792 ( .A(n15448), .ZN(n10370) );
  INV_X1 U11793 ( .A(n15480), .ZN(n10359) );
  NAND2_X1 U11794 ( .A1(n15273), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15313) );
  NAND2_X1 U11795 ( .A1(n15656), .A2(n10376), .ZN(n15568) );
  INV_X1 U11796 ( .A(n15079), .ZN(n14977) );
  INV_X1 U11797 ( .A(n14559), .ZN(n14557) );
  INV_X1 U11798 ( .A(n13885), .ZN(n13884) );
  NAND2_X1 U11799 ( .A1(n13689), .A2(n13688), .ZN(n13885) );
  INV_X1 U11800 ( .A(n15928), .ZN(n10100) );
  AND2_X1 U11801 ( .A1(n16103), .A2(n16158), .ZN(n10146) );
  AND3_X1 U11802 ( .A1(n15928), .A2(n15938), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10141) );
  NAND2_X1 U11803 ( .A1(n10148), .A2(n16103), .ZN(n10144) );
  NAND2_X1 U11804 ( .A1(n10166), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15977) );
  INV_X1 U11805 ( .A(n16012), .ZN(n10166) );
  NAND2_X1 U11806 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10257) );
  NAND2_X1 U11807 ( .A1(n10165), .A2(n12890), .ZN(n15997) );
  INV_X1 U11808 ( .A(n15977), .ZN(n10165) );
  AND2_X1 U11809 ( .A1(n13023), .A2(n13022), .ZN(n14764) );
  NAND3_X1 U11810 ( .A1(n9996), .A2(n12809), .A3(n12808), .ZN(n10197) );
  INV_X1 U11811 ( .A(n17878), .ZN(n10196) );
  AND2_X1 U11812 ( .A1(n13145), .A2(n13144), .ZN(n13754) );
  NAND2_X1 U11813 ( .A1(n14665), .A2(n13517), .ZN(n12788) );
  NAND2_X1 U11814 ( .A1(n9946), .A2(n12642), .ZN(n10274) );
  INV_X1 U11815 ( .A(n13751), .ZN(n14293) );
  OR2_X1 U11816 ( .A1(n14303), .A2(n14302), .ZN(n17843) );
  OR2_X1 U11817 ( .A1(n11027), .A2(n11026), .ZN(n11428) );
  NAND2_X1 U11818 ( .A1(n10340), .A2(n16513), .ZN(n16516) );
  NAND2_X1 U11819 ( .A1(n10322), .A2(n9781), .ZN(n10340) );
  INV_X1 U11820 ( .A(n16993), .ZN(n10339) );
  NAND2_X1 U11821 ( .A1(n9896), .A2(n11024), .ZN(n11023) );
  INV_X1 U11822 ( .A(n11027), .ZN(n9896) );
  OR2_X2 U11823 ( .A1(n10970), .A2(n11473), .ZN(n11456) );
  INV_X1 U11824 ( .A(n10881), .ZN(n9898) );
  INV_X1 U11825 ( .A(n10882), .ZN(n9897) );
  INV_X1 U11826 ( .A(n20180), .ZN(n20150) );
  NAND2_X1 U11827 ( .A1(n12454), .A2(n12455), .ZN(n12458) );
  NOR2_X1 U11828 ( .A1(n13870), .A2(n10389), .ZN(n14433) );
  NAND2_X1 U11829 ( .A1(n10390), .A2(n10550), .ZN(n10389) );
  AND3_X1 U11830 ( .A1(n11264), .A2(n11263), .A3(n11262), .ZN(n13981) );
  INV_X1 U11831 ( .A(n10382), .ZN(n10381) );
  OAI21_X1 U11832 ( .B1(n10384), .B2(n9709), .A(n13977), .ZN(n10382) );
  AOI22_X1 U11833 ( .A1(n14410), .A2(n12192), .B1(n12191), .B2(n14389), .ZN(
        n14346) );
  INV_X1 U11834 ( .A(n16875), .ZN(n16850) );
  AND2_X1 U11835 ( .A1(n11635), .A2(n11633), .ZN(n16415) );
  INV_X1 U11836 ( .A(n11600), .ZN(n11155) );
  INV_X1 U11837 ( .A(n11591), .ZN(n11154) );
  NAND2_X1 U11838 ( .A1(n11479), .A2(n9914), .ZN(n9913) );
  OR2_X1 U11839 ( .A1(n10409), .A2(n11485), .ZN(n9914) );
  NAND2_X1 U11840 ( .A1(n10127), .A2(n10562), .ZN(n16929) );
  NOR2_X1 U11841 ( .A1(n16973), .A2(n16976), .ZN(n14857) );
  NAND2_X1 U11842 ( .A1(n10066), .A2(n10444), .ZN(n10063) );
  AND2_X1 U11843 ( .A1(n17033), .A2(n10453), .ZN(n16991) );
  NOR2_X1 U11844 ( .A1(n10454), .A2(n17277), .ZN(n10453) );
  INV_X1 U11845 ( .A(n10455), .ZN(n10454) );
  NAND2_X1 U11846 ( .A1(n14836), .A2(n10421), .ZN(n16526) );
  AND2_X1 U11847 ( .A1(n14836), .A2(n14837), .ZN(n16528) );
  OR2_X1 U11848 ( .A1(n11011), .A2(n17007), .ZN(n11435) );
  NAND2_X1 U11849 ( .A1(n17033), .A2(n10457), .ZN(n14834) );
  AND2_X1 U11850 ( .A1(n10434), .A2(n17016), .ZN(n10433) );
  OR2_X1 U11851 ( .A1(n10437), .A2(n10435), .ZN(n10434) );
  NAND2_X1 U11852 ( .A1(n10401), .A2(n10402), .ZN(n14847) );
  NAND2_X1 U11853 ( .A1(n10415), .A2(n9713), .ZN(n16755) );
  AND2_X1 U11854 ( .A1(n17099), .A2(n9870), .ZN(n17056) );
  AND2_X1 U11855 ( .A1(n17099), .A2(n17301), .ZN(n17074) );
  BUF_X1 U11856 ( .A(n17032), .Z(n17099) );
  NAND2_X1 U11857 ( .A1(n9801), .A2(n9934), .ZN(n17105) );
  CLKBUF_X1 U11858 ( .A(n17104), .Z(n17107) );
  NAND2_X1 U11859 ( .A1(n10940), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10226) );
  NAND2_X1 U11860 ( .A1(n10224), .A2(n10050), .ZN(n17133) );
  AOI21_X1 U11861 ( .B1(n9687), .B2(n10022), .A(n9849), .ZN(n10050) );
  NAND2_X1 U11862 ( .A1(n10225), .A2(n9836), .ZN(n10224) );
  NOR2_X1 U11863 ( .A1(n11477), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10022) );
  AND3_X1 U11864 ( .A1(n11246), .A2(n11245), .A3(n11244), .ZN(n14778) );
  AND2_X1 U11865 ( .A1(n10053), .A2(n10052), .ZN(n11076) );
  OR2_X1 U11866 ( .A1(n11071), .A2(n17432), .ZN(n10052) );
  NAND2_X1 U11867 ( .A1(n17177), .A2(n9958), .ZN(n10445) );
  AND2_X1 U11868 ( .A1(n11071), .A2(n17432), .ZN(n9958) );
  NAND2_X1 U11869 ( .A1(n10443), .A2(n17423), .ZN(n17144) );
  NAND3_X1 U11870 ( .A1(n10934), .A2(n11084), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17146) );
  AOI22_X1 U11871 ( .A1(n17156), .A2(n17157), .B1(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n20188), .ZN(n17141) );
  OAI21_X1 U11872 ( .B1(n11099), .B2(n11098), .A(n11097), .ZN(n11101) );
  INV_X1 U11873 ( .A(n17439), .ZN(n10314) );
  AND2_X1 U11874 ( .A1(n11237), .A2(n11231), .ZN(n10404) );
  INV_X1 U11875 ( .A(n16598), .ZN(n11237) );
  INV_X1 U11876 ( .A(n17178), .ZN(n10449) );
  NAND2_X1 U11877 ( .A1(n10872), .A2(n11482), .ZN(n10474) );
  AND2_X1 U11878 ( .A1(n10483), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10482) );
  OR2_X1 U11879 ( .A1(n10484), .A2(n11482), .ZN(n10483) );
  NAND2_X1 U11880 ( .A1(n13900), .A2(n13901), .ZN(n13903) );
  NAND2_X1 U11881 ( .A1(n10792), .A2(n14360), .ZN(n10900) );
  BUF_X1 U11882 ( .A(n10911), .Z(n20456) );
  AND2_X1 U11883 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20504) );
  OR2_X1 U11884 ( .A1(n20921), .A2(n20912), .ZN(n20506) );
  NAND2_X1 U11885 ( .A1(n20584), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n9953) );
  NOR2_X1 U11886 ( .A1(n20536), .A2(n20563), .ZN(n9952) );
  AOI21_X1 U11887 ( .B1(n20534), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n9955) );
  NOR2_X1 U11888 ( .A1(n9951), .A2(n20563), .ZN(n9950) );
  INV_X1 U11889 ( .A(n9953), .ZN(n9951) );
  NAND2_X1 U11890 ( .A1(n20557), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n9954) );
  NAND2_X1 U11891 ( .A1(n20921), .A2(n20912), .ZN(n20562) );
  NAND2_X1 U11892 ( .A1(n10789), .A2(n14360), .ZN(n20655) );
  OR3_X1 U11893 ( .A1(n20689), .A2(n20720), .A3(n20939), .ZN(n20696) );
  OR2_X1 U11894 ( .A1(n20921), .A2(n20931), .ZN(n20695) );
  INV_X1 U11895 ( .A(n10947), .ZN(n17503) );
  OR2_X1 U11896 ( .A1(n20969), .A2(n17482), .ZN(n17483) );
  AOI21_X1 U11897 ( .B1(n12064), .B2(n12063), .A(n12147), .ZN(n19878) );
  AND2_X1 U11898 ( .A1(n14235), .A2(n14234), .ZN(n19884) );
  INV_X1 U11899 ( .A(n13429), .ZN(n14234) );
  XNOR2_X1 U11900 ( .A(n12127), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n18064) );
  NAND2_X1 U11901 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18569), .ZN(n18563) );
  OR2_X1 U11902 ( .A1(n11775), .A2(n11774), .ZN(n12081) );
  AND3_X1 U11903 ( .A1(n10159), .A2(n11680), .A3(n11679), .ZN(n10158) );
  NAND2_X1 U11904 ( .A1(n13363), .A2(n13377), .ZN(n13429) );
  NOR2_X1 U11905 ( .A1(n18039), .A2(n20032), .ZN(n10084) );
  AND4_X1 U11906 ( .A1(n11939), .A2(n11938), .A3(n11937), .A4(n11936), .ZN(
        n11940) );
  NAND2_X1 U11907 ( .A1(n17599), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17600) );
  NAND2_X1 U11908 ( .A1(n18908), .A2(n9757), .ZN(n18848) );
  NOR2_X1 U11909 ( .A1(n18892), .A2(n10295), .ZN(n10294) );
  AND2_X1 U11910 ( .A1(n19281), .A2(n10157), .ZN(n18813) );
  NAND2_X1 U11911 ( .A1(n18971), .A2(n10289), .ZN(n18922) );
  AND2_X1 U11912 ( .A1(n18968), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10289) );
  OR2_X1 U11913 ( .A1(n13458), .A2(n19379), .ZN(n11817) );
  NAND2_X1 U11915 ( .A1(n10152), .A2(n10302), .ZN(n11865) );
  NAND4_X2 U11916 ( .A1(n11982), .A2(n11981), .A3(n11980), .A4(n11979), .ZN(
        n20031) );
  AND3_X1 U11917 ( .A1(n11974), .A2(n11973), .A3(n11972), .ZN(n11980) );
  AOI22_X1 U11918 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11981) );
  NAND2_X1 U11919 ( .A1(n18830), .A2(n10025), .ZN(n18815) );
  AND2_X1 U11920 ( .A1(n11862), .A2(n10160), .ZN(n10025) );
  INV_X1 U11921 ( .A(n18951), .ZN(n10028) );
  INV_X1 U11922 ( .A(n19387), .ZN(n19875) );
  NAND4_X1 U11923 ( .A1(n11796), .A2(n11795), .A3(n11794), .A4(n11793), .ZN(
        n17632) );
  NOR2_X1 U11924 ( .A1(n19041), .A2(n19040), .ZN(n19039) );
  NAND2_X1 U11925 ( .A1(n9985), .A2(n9983), .ZN(n9981) );
  NAND2_X1 U11926 ( .A1(n19065), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n19067) );
  INV_X1 U11927 ( .A(n19093), .ZN(n9975) );
  NAND2_X1 U11928 ( .A1(n11827), .A2(n9976), .ZN(n9970) );
  INV_X1 U11929 ( .A(n19306), .ZN(n19283) );
  NOR2_X1 U11930 ( .A1(n18039), .A2(n19914), .ZN(n18742) );
  AND4_X1 U11931 ( .A1(n11948), .A2(n11947), .A3(n11946), .A4(n11945), .ZN(
        n11960) );
  NOR2_X1 U11932 ( .A1(n19920), .A2(n20047), .ZN(n20038) );
  OR2_X1 U11933 ( .A1(n11469), .A2(n11468), .ZN(n14789) );
  AND2_X1 U11934 ( .A1(n21116), .A2(n15824), .ZN(n21111) );
  INV_X1 U11935 ( .A(n21116), .ZN(n15818) );
  NOR2_X1 U11936 ( .A1(n9732), .A2(n15380), .ZN(n10364) );
  NOR2_X1 U11937 ( .A1(n10373), .A2(n10372), .ZN(n10371) );
  NOR2_X1 U11938 ( .A1(n15822), .A2(n17937), .ZN(n10373) );
  INV_X1 U11939 ( .A(n15420), .ZN(n10372) );
  NAND2_X1 U11940 ( .A1(n15448), .A2(n10364), .ZN(n10363) );
  OR2_X1 U11941 ( .A1(n10369), .A2(n9732), .ZN(n10366) );
  NAND2_X1 U11942 ( .A1(n10136), .A2(n15715), .ZN(n16085) );
  NAND2_X1 U11943 ( .A1(n10138), .A2(n10137), .ZN(n10136) );
  INV_X1 U11944 ( .A(n15716), .ZN(n10137) );
  INV_X1 U11945 ( .A(n15717), .ZN(n10138) );
  NAND2_X1 U11946 ( .A1(n20989), .A2(n13524), .ZN(n17885) );
  NOR2_X1 U11947 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n10265), .ZN(
        n10264) );
  INV_X1 U11948 ( .A(n16131), .ZN(n10265) );
  AND2_X1 U11949 ( .A1(n16259), .A2(n16165), .ZN(n10268) );
  INV_X1 U11950 ( .A(n17899), .ZN(n17906) );
  AND2_X1 U11951 ( .A1(n13146), .A2(n13122), .ZN(n17922) );
  INV_X1 U11952 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21422) );
  INV_X1 U11953 ( .A(n21586), .ZN(n21584) );
  NAND2_X1 U11954 ( .A1(n11645), .A2(n11644), .ZN(n13221) );
  NAND2_X1 U11955 ( .A1(n12499), .A2(n17819), .ZN(n12500) );
  AOI21_X1 U11956 ( .B1(n10322), .B2(n10330), .A(n10333), .ZN(n10329) );
  NAND2_X1 U11957 ( .A1(n10322), .A2(n10322), .ZN(n10331) );
  OAI21_X1 U11958 ( .B1(n10336), .B2(n20147), .A(n10334), .ZN(n10333) );
  NAND2_X1 U11959 ( .A1(n20180), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20145) );
  AND2_X1 U11960 ( .A1(n12251), .A2(n9847), .ZN(n10470) );
  AOI21_X1 U11961 ( .B1(n11650), .B2(n12189), .A(n11649), .ZN(n16773) );
  NOR2_X1 U11962 ( .A1(n20227), .A2(n12194), .ZN(n14700) );
  AOI21_X1 U11963 ( .B1(n14892), .B2(n9968), .A(n9964), .ZN(n9962) );
  NAND2_X1 U11964 ( .A1(n17196), .A2(n9965), .ZN(n9964) );
  NAND2_X1 U11965 ( .A1(n11549), .A2(n9968), .ZN(n9965) );
  OR2_X1 U11966 ( .A1(n14798), .A2(n17166), .ZN(n9992) );
  NAND2_X1 U11967 ( .A1(n9933), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10116) );
  AND2_X1 U11968 ( .A1(n11089), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10055) );
  AND2_X1 U11969 ( .A1(n17187), .A2(n13341), .ZN(n17190) );
  INV_X1 U11970 ( .A(n17187), .ZN(n17172) );
  AND2_X1 U11971 ( .A1(n11090), .A2(n13223), .ZN(n17196) );
  OR2_X1 U11972 ( .A1(n13219), .A2(n13223), .ZN(n17181) );
  NAND2_X1 U11973 ( .A1(n17187), .A2(n20929), .ZN(n17166) );
  XNOR2_X1 U11974 ( .A(n11648), .B(n11518), .ZN(n16764) );
  NAND2_X1 U11975 ( .A1(n10220), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10218) );
  AND2_X1 U11976 ( .A1(n10219), .A2(n11483), .ZN(n10217) );
  NOR3_X1 U11977 ( .A1(n17216), .A2(n11563), .A3(n10175), .ZN(n10179) );
  OAI211_X1 U11978 ( .C1(n14901), .C2(n9915), .A(n9912), .B(n9910), .ZN(n15428) );
  NAND2_X1 U11979 ( .A1(n11479), .A2(n9916), .ZN(n9915) );
  NAND2_X1 U11980 ( .A1(n14901), .A2(n9911), .ZN(n9910) );
  OAI21_X1 U11981 ( .B1(n11485), .B2(n11479), .A(n9913), .ZN(n9912) );
  XNOR2_X1 U11982 ( .A(n10019), .B(n12179), .ZN(n16910) );
  OAI21_X1 U11983 ( .B1(n10209), .B2(n10410), .A(n10017), .ZN(n10019) );
  INV_X1 U11984 ( .A(n10018), .ZN(n10017) );
  OAI21_X1 U11985 ( .B1(n14892), .B2(n11549), .A(n9968), .ZN(n9963) );
  NOR2_X1 U11986 ( .A1(n14902), .A2(n14887), .ZN(n10189) );
  OAI21_X1 U11987 ( .B1(n14909), .B2(n17444), .A(n14908), .ZN(n14910) );
  XNOR2_X1 U11988 ( .A(n14901), .B(n9764), .ZN(n16919) );
  NOR2_X1 U11989 ( .A1(n14798), .A2(n17429), .ZN(n10185) );
  NAND2_X1 U11990 ( .A1(n14892), .A2(n9993), .ZN(n14812) );
  NAND2_X1 U11991 ( .A1(n9994), .A2(n14887), .ZN(n9993) );
  INV_X1 U11992 ( .A(n16922), .ZN(n9994) );
  NAND2_X1 U11993 ( .A1(n10491), .A2(n10487), .ZN(n10486) );
  NAND2_X1 U11994 ( .A1(n10113), .A2(n9933), .ZN(n10114) );
  AND2_X1 U11995 ( .A1(n16966), .A2(n9737), .ZN(n10113) );
  OAI211_X1 U11996 ( .C1(n17032), .C2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n17021), .B(n10054), .ZN(n17295) );
  NAND2_X1 U11997 ( .A1(n14835), .A2(n10458), .ZN(n10054) );
  XNOR2_X1 U11998 ( .A(n10432), .B(n17018), .ZN(n17299) );
  AOI21_X1 U11999 ( .B1(n10431), .B2(n10437), .A(n10436), .ZN(n10432) );
  NAND2_X1 U12000 ( .A1(n11415), .A2(n11414), .ZN(n17429) );
  INV_X1 U12001 ( .A(n17461), .ZN(n17444) );
  NAND2_X1 U12002 ( .A1(n11415), .A2(n11204), .ZN(n17458) );
  NOR2_X2 U12003 ( .A1(n11402), .A2(n20953), .ZN(n17454) );
  INV_X1 U12004 ( .A(n17429), .ZN(n17456) );
  INV_X1 U12005 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20938) );
  INV_X1 U12006 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20927) );
  NAND2_X1 U12007 ( .A1(n17455), .A2(n12225), .ZN(n12227) );
  NAND2_X1 U12008 ( .A1(n13899), .A2(n13776), .ZN(n13777) );
  NAND2_X1 U12009 ( .A1(n14410), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17484) );
  INV_X1 U12010 ( .A(n20555), .ZN(n20557) );
  NOR2_X1 U12011 ( .A1(n19884), .A2(n18033), .ZN(n20051) );
  INV_X1 U12012 ( .A(n18742), .ZN(n18033) );
  XNOR2_X1 U12013 ( .A(n18083), .B(n10292), .ZN(n10291) );
  INV_X1 U12014 ( .A(n18084), .ZN(n10292) );
  OR2_X1 U12015 ( .A1(n18086), .A2(n18085), .ZN(n10290) );
  INV_X1 U12016 ( .A(n18416), .ZN(n18436) );
  NAND2_X1 U12017 ( .A1(n18505), .A2(n10245), .ZN(n18492) );
  AND2_X1 U12018 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n10246), .ZN(n10245) );
  NOR2_X1 U12019 ( .A1(n18448), .A2(n10247), .ZN(n10246) );
  NAND2_X1 U12020 ( .A1(n13359), .A2(n9742), .ZN(n13579) );
  INV_X1 U12021 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n18564) );
  NOR2_X1 U12022 ( .A1(n12001), .A2(n12000), .ZN(n12002) );
  OR2_X2 U12023 ( .A1(n13457), .A2(n18576), .ZN(n18662) );
  OR2_X1 U12024 ( .A1(n13457), .A2(n13433), .ZN(n18638) );
  OR2_X1 U12025 ( .A1(n13457), .A2(n19448), .ZN(n18636) );
  INV_X1 U12026 ( .A(n18813), .ZN(n19236) );
  AND2_X1 U12027 ( .A1(n19119), .A2(n17632), .ZN(n19015) );
  INV_X1 U12028 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18678) );
  NOR2_X1 U12029 ( .A1(n19174), .A2(n9841), .ZN(n19186) );
  NAND2_X1 U12030 ( .A1(n12912), .A2(n12901), .ZN(n12906) );
  NOR2_X1 U12031 ( .A1(n10236), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10235) );
  INV_X1 U12032 ( .A(n10500), .ZN(n10236) );
  NOR2_X1 U12033 ( .A1(n12810), .A2(n9843), .ZN(n10500) );
  NAND2_X1 U12034 ( .A1(n12948), .A2(n12921), .ZN(n12952) );
  INV_X1 U12035 ( .A(n12783), .ZN(n10507) );
  NOR2_X1 U12036 ( .A1(n12640), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10001) );
  AND4_X1 U12037 ( .A1(n10944), .A2(n10943), .A3(n10942), .A4(n10941), .ZN(
        n10954) );
  NAND2_X1 U12038 ( .A1(n20537), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10817) );
  INV_X1 U12039 ( .A(n11384), .ZN(n10694) );
  AND2_X2 U12040 ( .A1(n14370), .A2(n10575), .ZN(n10606) );
  NAND2_X1 U12041 ( .A1(n12319), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10682) );
  OR2_X1 U12042 ( .A1(n12907), .A2(n12919), .ZN(n12909) );
  AND2_X1 U12043 ( .A1(n12909), .A2(n12897), .ZN(n12911) );
  OR2_X1 U12044 ( .A1(n12821), .A2(n12820), .ZN(n12828) );
  INV_X1 U12045 ( .A(n12743), .ZN(n12745) );
  NOR2_X1 U12046 ( .A1(n12878), .A2(n13061), .ZN(n10007) );
  OR2_X1 U12047 ( .A1(n12724), .A2(n12723), .ZN(n12789) );
  NAND2_X1 U12048 ( .A1(n13145), .A2(n9876), .ZN(n9875) );
  INV_X1 U12049 ( .A(n15823), .ZN(n12929) );
  NAND2_X1 U12050 ( .A1(n12635), .A2(n14469), .ZN(n12648) );
  OAI21_X1 U12051 ( .B1(n12636), .B2(n12632), .A(n14464), .ZN(n10509) );
  NAND2_X1 U12052 ( .A1(n14460), .A2(n12588), .ZN(n12587) );
  AND2_X2 U12053 ( .A1(n13503), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12517) );
  AND2_X1 U12054 ( .A1(n12971), .A2(n12970), .ZN(n13134) );
  NAND2_X1 U12055 ( .A1(n9921), .A2(n11208), .ZN(n10713) );
  NAND2_X1 U12056 ( .A1(n10611), .A2(n14353), .ZN(n10495) );
  NAND2_X1 U12057 ( .A1(n10616), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10494) );
  NOR2_X1 U12058 ( .A1(n10730), .A2(n9988), .ZN(n10733) );
  NAND2_X1 U12059 ( .A1(n10570), .A2(n10572), .ZN(n9889) );
  NAND2_X1 U12060 ( .A1(n9932), .A2(n10920), .ZN(n9925) );
  NAND2_X1 U12061 ( .A1(n9691), .A2(n10780), .ZN(n10048) );
  NAND2_X1 U12062 ( .A1(n10792), .A2(n16635), .ZN(n10903) );
  NAND2_X1 U12063 ( .A1(n10582), .A2(n10581), .ZN(n10585) );
  OR2_X1 U12064 ( .A1(n11172), .A2(n11046), .ZN(n10582) );
  AND2_X1 U12065 ( .A1(n10873), .A2(n10583), .ZN(n10584) );
  NAND2_X1 U12066 ( .A1(n10585), .A2(n10584), .ZN(n10874) );
  NAND2_X1 U12067 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20947), .ZN(
        n11046) );
  AOI21_X1 U12068 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n19890), .A(
        n12061), .ZN(n12068) );
  AND2_X1 U12069 ( .A1(n11687), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11685) );
  INV_X1 U12070 ( .A(n11827), .ZN(n9972) );
  INV_X1 U12071 ( .A(n10016), .ZN(n11823) );
  AND2_X1 U12072 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11686) );
  AND4_X1 U12073 ( .A1(n10855), .A2(n10854), .A3(n10853), .A4(n10852), .ZN(
        n10870) );
  AOI221_X1 U12074 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12915), 
        .C1(n13764), .C2(n12915), .A(n12914), .ZN(n12960) );
  NOR2_X1 U12075 ( .A1(n14449), .A2(n15395), .ZN(n12630) );
  NOR2_X2 U12076 ( .A1(n15122), .A2(n15588), .ZN(n15088) );
  AND2_X1 U12077 ( .A1(n15085), .A2(n15657), .ZN(n15086) );
  AND2_X1 U12078 ( .A1(n14548), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14647) );
  INV_X1 U12079 ( .A(n15492), .ZN(n10534) );
  NOR2_X1 U12080 ( .A1(n10536), .A2(n15505), .ZN(n10535) );
  INV_X1 U12081 ( .A(n15519), .ZN(n10536) );
  NAND2_X1 U12082 ( .A1(n16103), .A2(n12882), .ZN(n10516) );
  INV_X1 U12083 ( .A(n12885), .ZN(n10514) );
  INV_X1 U12084 ( .A(n9861), .ZN(n10530) );
  AND2_X1 U12085 ( .A1(n10532), .A2(n13072), .ZN(n10531) );
  INV_X1 U12086 ( .A(n15610), .ZN(n10532) );
  NAND2_X1 U12087 ( .A1(n16103), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10092) );
  AND2_X1 U12088 ( .A1(n10519), .A2(n13053), .ZN(n10518) );
  INV_X1 U12089 ( .A(n15669), .ZN(n10519) );
  INV_X1 U12090 ( .A(n10163), .ZN(n10162) );
  NAND2_X1 U12091 ( .A1(n10277), .A2(n9712), .ZN(n10009) );
  NAND2_X1 U12092 ( .A1(n12832), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12833) );
  AND2_X1 U12093 ( .A1(n12638), .A2(n13126), .ZN(n12969) );
  INV_X1 U12094 ( .A(n12626), .ZN(n12966) );
  INV_X1 U12095 ( .A(n12965), .ZN(n10260) );
  NAND2_X1 U12096 ( .A1(n13680), .A2(n13679), .ZN(n12737) );
  INV_X1 U12097 ( .A(n21737), .ZN(n14299) );
  INV_X1 U12098 ( .A(n12588), .ZN(n13126) );
  NAND2_X1 U12099 ( .A1(n12731), .A2(n12730), .ZN(n14666) );
  AOI22_X1 U12100 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12589), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12591) );
  NAND2_X1 U12101 ( .A1(n12687), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12603) );
  AOI22_X1 U12102 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12605), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12513) );
  NAND2_X1 U12103 ( .A1(n11449), .A2(n9844), .ZN(n11461) );
  NAND2_X1 U12104 ( .A1(n11461), .A2(n11456), .ZN(n11464) );
  AOI21_X1 U12105 ( .B1(n10322), .B2(n10325), .A(n10324), .ZN(n10323) );
  INV_X1 U12106 ( .A(n17815), .ZN(n10324) );
  NOR2_X1 U12107 ( .A1(n10964), .A2(n10963), .ZN(n11247) );
  INV_X1 U12108 ( .A(n20964), .ZN(n11651) );
  NAND2_X1 U12109 ( .A1(n10748), .A2(n10747), .ZN(n10765) );
  CLKBUF_X1 U12110 ( .A(n12325), .Z(n16657) );
  CLKBUF_X1 U12111 ( .A(n12316), .Z(n16658) );
  CLKBUF_X1 U12112 ( .A(n12317), .Z(n16664) );
  CLKBUF_X1 U12113 ( .A(n12319), .Z(n16663) );
  CLKBUF_X1 U12114 ( .A(n9696), .Z(n16662) );
  CLKBUF_X1 U12115 ( .A(n12324), .Z(n16656) );
  CLKBUF_X1 U12116 ( .A(n12379), .Z(n12329) );
  AND2_X1 U12117 ( .A1(n12284), .A2(n16745), .ZN(n10469) );
  NAND2_X1 U12118 ( .A1(n16749), .A2(n16758), .ZN(n10125) );
  INV_X1 U12119 ( .A(n16759), .ZN(n10124) );
  NOR2_X1 U12120 ( .A1(n9709), .A2(n10388), .ZN(n10379) );
  AND2_X1 U12121 ( .A1(n11571), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11611) );
  NAND2_X1 U12122 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10349) );
  OR2_X1 U12123 ( .A1(n10349), .A2(n10348), .ZN(n10347) );
  NOR2_X1 U12124 ( .A1(n10410), .A2(n12178), .ZN(n10409) );
  AND2_X1 U12125 ( .A1(n11470), .A2(n14791), .ZN(n10408) );
  NOR2_X1 U12126 ( .A1(n17230), .A2(n11563), .ZN(n14815) );
  INV_X1 U12127 ( .A(n10063), .ZN(n10061) );
  INV_X1 U12128 ( .A(n9755), .ZN(n10060) );
  AND2_X1 U12129 ( .A1(n14837), .A2(n16527), .ZN(n10421) );
  NOR2_X1 U12130 ( .A1(n17007), .A2(n10458), .ZN(n10457) );
  OR2_X1 U12131 ( .A1(n11006), .A2(n10436), .ZN(n10435) );
  NOR2_X1 U12132 ( .A1(n10435), .A2(n17038), .ZN(n10430) );
  AND2_X1 U12133 ( .A1(n9815), .A2(n9934), .ZN(n10202) );
  INV_X1 U12134 ( .A(n14431), .ZN(n10401) );
  OR2_X1 U12135 ( .A1(n14701), .A2(n14589), .ZN(n11137) );
  AND2_X1 U12136 ( .A1(n10392), .A2(n9864), .ZN(n10390) );
  AND3_X1 U12137 ( .A1(n11279), .A2(n11278), .A3(n11277), .ZN(n13871) );
  NAND2_X1 U12138 ( .A1(n9942), .A2(n11085), .ZN(n11087) );
  NAND2_X1 U12139 ( .A1(n9941), .A2(n11482), .ZN(n9940) );
  NAND2_X1 U12140 ( .A1(n9942), .A2(n9939), .ZN(n9938) );
  AND2_X1 U12141 ( .A1(n11085), .A2(n11477), .ZN(n9939) );
  NAND2_X1 U12142 ( .A1(n9687), .A2(n11482), .ZN(n10225) );
  AND2_X1 U12143 ( .A1(n11389), .A2(n11208), .ZN(n11372) );
  NAND2_X1 U12144 ( .A1(n11096), .A2(n10765), .ZN(n11097) );
  NAND3_X2 U12145 ( .A1(n9928), .A2(n9929), .A3(n10811), .ZN(n10841) );
  INV_X1 U12146 ( .A(n10757), .ZN(n9909) );
  AOI21_X1 U12147 ( .B1(n10753), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10752), .ZN(n10757) );
  AND2_X1 U12148 ( .A1(n20959), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10752) );
  AND2_X1 U12149 ( .A1(n10711), .A2(n10722), .ZN(n11371) );
  NAND2_X1 U12150 ( .A1(n11045), .A2(n10709), .ZN(n10711) );
  NAND2_X1 U12151 ( .A1(n10739), .A2(n10738), .ZN(n10763) );
  AND2_X2 U12152 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14331) );
  AND2_X1 U12153 ( .A1(n10721), .A2(n13780), .ZN(n10051) );
  OAI21_X1 U12154 ( .B1(n11179), .B2(n11178), .A(n10173), .ZN(n10172) );
  AOI21_X1 U12155 ( .B1(n9887), .B2(n11178), .A(n10174), .ZN(n10173) );
  NAND2_X1 U12156 ( .A1(n10174), .A2(n13389), .ZN(n10320) );
  INV_X1 U12157 ( .A(n10048), .ZN(n10056) );
  NAND2_X1 U12158 ( .A1(n11673), .A2(n13393), .ZN(n17769) );
  AND2_X1 U12159 ( .A1(n11685), .A2(n11684), .ZN(n13345) );
  INV_X1 U12160 ( .A(n11703), .ZN(n12012) );
  NAND2_X1 U12161 ( .A1(n12113), .A2(n13191), .ZN(n10299) );
  NOR2_X1 U12162 ( .A1(n11971), .A2(n11970), .ZN(n11982) );
  NAND3_X1 U12163 ( .A1(n9758), .A2(n10538), .A3(n19043), .ZN(n18938) );
  NOR2_X1 U12164 ( .A1(n19039), .A2(n19317), .ZN(n12105) );
  INV_X1 U12165 ( .A(n9983), .ZN(n9980) );
  NAND2_X1 U12166 ( .A1(n19089), .A2(n12097), .ZN(n12098) );
  NAND2_X1 U12167 ( .A1(n19448), .A2(n10081), .ZN(n12034) );
  NOR2_X1 U12168 ( .A1(n12034), .A2(n12032), .ZN(n12040) );
  NOR2_X1 U12169 ( .A1(n13537), .A2(n13539), .ZN(n17797) );
  NAND2_X1 U12170 ( .A1(n11682), .A2(n11686), .ZN(n17799) );
  INV_X1 U12171 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n21017) );
  NAND2_X1 U12172 ( .A1(n21074), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15777) );
  INV_X1 U12173 ( .A(n14769), .ZN(n10357) );
  NAND2_X1 U12174 ( .A1(n14760), .A2(n14759), .ZN(n14761) );
  NAND2_X1 U12175 ( .A1(n15353), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15381) );
  INV_X1 U12176 ( .A(n15352), .ZN(n15353) );
  OAI21_X1 U12177 ( .B1(n15923), .B2(n15565), .A(n15333), .ZN(n15480) );
  AND2_X1 U12178 ( .A1(n15272), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15273) );
  NAND2_X1 U12179 ( .A1(n15295), .A2(n15294), .ZN(n15501) );
  OR2_X1 U12180 ( .A1(n15942), .A2(n15565), .ZN(n15295) );
  AND2_X1 U12181 ( .A1(n15227), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15228) );
  INV_X1 U12182 ( .A(n15226), .ZN(n15227) );
  NAND2_X1 U12183 ( .A1(n15228), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15271) );
  AND2_X1 U12184 ( .A1(n9771), .A2(n15534), .ZN(n10374) );
  AND2_X1 U12185 ( .A1(n15656), .A2(n9771), .ZN(n15547) );
  INV_X1 U12186 ( .A(n15568), .ZN(n10034) );
  AND2_X1 U12187 ( .A1(n15596), .A2(n15608), .ZN(n10039) );
  INV_X1 U12188 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15186) );
  AND2_X1 U12189 ( .A1(n15087), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15187) );
  AND3_X1 U12190 ( .A1(n15156), .A2(n15155), .A3(n15154), .ZN(n15639) );
  OR2_X1 U12191 ( .A1(n15658), .A2(n15639), .ZN(n15641) );
  NAND2_X1 U12192 ( .A1(n14980), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15153) );
  AND2_X1 U12193 ( .A1(n14979), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14980) );
  INV_X1 U12194 ( .A(n15031), .ZN(n14979) );
  NAND2_X1 U12195 ( .A1(n15656), .A2(n15086), .ZN(n15658) );
  NAND2_X1 U12196 ( .A1(n15656), .A2(n15657), .ZN(n15674) );
  NOR2_X1 U12197 ( .A1(n15063), .A2(n14978), .ZN(n15027) );
  NAND2_X1 U12198 ( .A1(n15027), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15031) );
  NAND2_X1 U12199 ( .A1(n14997), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15063) );
  INV_X1 U12200 ( .A(n14975), .ZN(n14976) );
  NOR2_X1 U12201 ( .A1(n14958), .A2(n14957), .ZN(n15893) );
  INV_X1 U12202 ( .A(n15656), .ZN(n15741) );
  NAND2_X1 U12203 ( .A1(n14952), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14975) );
  NOR2_X2 U12204 ( .A1(n14753), .A2(n21017), .ZN(n14952) );
  NAND2_X1 U12205 ( .A1(n12806), .A2(n14601), .ZN(n12808) );
  NAND2_X1 U12206 ( .A1(n10194), .A2(n12773), .ZN(n12806) );
  INV_X1 U12207 ( .A(n12805), .ZN(n10192) );
  NAND2_X1 U12208 ( .A1(n10358), .A2(n14654), .ZN(n14768) );
  NAND2_X1 U12209 ( .A1(n14321), .A2(n14320), .ZN(n14330) );
  AND2_X1 U12210 ( .A1(n14327), .A2(n14326), .ZN(n14328) );
  NOR2_X1 U12211 ( .A1(n10498), .A2(n10497), .ZN(n10496) );
  NAND2_X1 U12212 ( .A1(n15967), .A2(n10283), .ZN(n10282) );
  NAND2_X1 U12213 ( .A1(n12890), .A2(n15936), .ZN(n10283) );
  AND2_X1 U12214 ( .A1(n15518), .A2(n9838), .ZN(n15491) );
  NAND2_X1 U12215 ( .A1(n15518), .A2(n10535), .ZN(n15503) );
  NAND2_X1 U12216 ( .A1(n10094), .A2(n10093), .ZN(n15947) );
  NOR2_X1 U12217 ( .A1(n10515), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10093) );
  NAND2_X1 U12218 ( .A1(n15975), .A2(n10513), .ZN(n10094) );
  AND2_X1 U12219 ( .A1(n13073), .A2(n9839), .ZN(n15599) );
  NAND2_X1 U12220 ( .A1(n13073), .A2(n13072), .ZN(n15628) );
  NAND2_X1 U12221 ( .A1(n15975), .A2(n16013), .ZN(n16012) );
  INV_X1 U12222 ( .A(n15648), .ZN(n13065) );
  INV_X1 U12223 ( .A(n15647), .ZN(n13066) );
  INV_X1 U12224 ( .A(n12878), .ZN(n10005) );
  NOR2_X1 U12225 ( .A1(n16074), .A2(n16072), .ZN(n16054) );
  AND2_X1 U12226 ( .A1(n13052), .A2(n13051), .ZN(n15688) );
  INV_X1 U12227 ( .A(n10526), .ZN(n10524) );
  NOR2_X1 U12228 ( .A1(n15761), .A2(n10526), .ZN(n15721) );
  INV_X1 U12229 ( .A(n10527), .ZN(n10525) );
  NAND2_X1 U12230 ( .A1(n10528), .A2(n10529), .ZN(n16343) );
  NAND2_X1 U12231 ( .A1(n10521), .A2(n14764), .ZN(n10520) );
  INV_X1 U12232 ( .A(n10522), .ZN(n10521) );
  NAND2_X1 U12233 ( .A1(n13795), .A2(n13794), .ZN(n9881) );
  NAND2_X1 U12234 ( .A1(n13750), .A2(n13113), .ZN(n12981) );
  INV_X1 U12235 ( .A(n13737), .ZN(n10086) );
  XNOR2_X1 U12236 ( .A(n13679), .B(n13680), .ZN(n14438) );
  NAND2_X1 U12237 ( .A1(n12801), .A2(n10015), .ZN(n12802) );
  INV_X1 U12238 ( .A(n13766), .ZN(n16350) );
  NAND2_X1 U12239 ( .A1(n10014), .A2(n12658), .ZN(n10161) );
  AND2_X1 U12240 ( .A1(n21294), .A2(n21586), .ZN(n21298) );
  OAI21_X1 U12241 ( .B1(n21384), .B2(n14711), .A(n21742), .ZN(n14717) );
  OAI21_X1 U12242 ( .B1(n21452), .B2(n21518), .A(n21742), .ZN(n21460) );
  NOR2_X1 U12243 ( .A1(n21455), .A2(n21189), .ZN(n21529) );
  NAND2_X1 U12244 ( .A1(n21186), .A2(n21185), .ZN(n21492) );
  OR2_X1 U12245 ( .A1(n13753), .A2(n21530), .ZN(n14313) );
  NOR2_X1 U12246 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20959) );
  NAND3_X1 U12247 ( .A1(n10717), .A2(n10710), .A3(n11382), .ZN(n11045) );
  NAND2_X1 U12248 ( .A1(n10876), .A2(n11048), .ZN(n10875) );
  OR2_X1 U12249 ( .A1(n14343), .A2(n11379), .ZN(n14387) );
  INV_X1 U12250 ( .A(n16914), .ZN(n10334) );
  NAND2_X1 U12252 ( .A1(n11464), .A2(n11459), .ZN(n11463) );
  INV_X1 U12253 ( .A(n10337), .ZN(n10336) );
  OAI21_X1 U12254 ( .B1(n20147), .B2(n10338), .A(n16398), .ZN(n10337) );
  INV_X1 U12255 ( .A(n16415), .ZN(n10338) );
  NOR2_X1 U12256 ( .A1(n11450), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10269) );
  NAND2_X1 U12257 ( .A1(n11449), .A2(n11448), .ZN(n16461) );
  AND2_X1 U12258 ( .A1(n11507), .A2(n11506), .ZN(n16457) );
  NAND2_X1 U12259 ( .A1(n10326), .A2(n16489), .ZN(n17814) );
  NAND2_X1 U12260 ( .A1(n16488), .A2(n10322), .ZN(n10326) );
  NAND2_X1 U12261 ( .A1(n10988), .A2(n9787), .ZN(n11009) );
  NAND2_X1 U12262 ( .A1(n10988), .A2(n9714), .ZN(n11003) );
  NAND2_X1 U12263 ( .A1(n10988), .A2(n10989), .ZN(n11000) );
  OR2_X1 U12264 ( .A1(n10271), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10270) );
  OR2_X1 U12265 ( .A1(n10971), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10271) );
  OR2_X1 U12266 ( .A1(n10970), .A2(n10971), .ZN(n10978) );
  NAND2_X1 U12267 ( .A1(n11207), .A2(n16619), .ZN(n10131) );
  NAND2_X1 U12268 ( .A1(n11031), .A2(n10878), .ZN(n10132) );
  INV_X1 U12269 ( .A(n16649), .ZN(n16616) );
  NOR2_X1 U12270 ( .A1(n10466), .A2(n16681), .ZN(n10465) );
  AND4_X1 U12271 ( .A1(n14249), .A2(n14491), .A3(n12250), .A4(n12249), .ZN(
        n12251) );
  AND2_X1 U12272 ( .A1(n11514), .A2(n11513), .ZN(n14813) );
  NOR2_X1 U12273 ( .A1(n16707), .A2(n12431), .ZN(n16692) );
  NOR2_X1 U12274 ( .A1(n10122), .A2(n9863), .ZN(n10121) );
  AND2_X1 U12275 ( .A1(n11365), .A2(n11364), .ZN(n11368) );
  NAND2_X1 U12276 ( .A1(n16744), .A2(n10469), .ZN(n16739) );
  INV_X1 U12277 ( .A(n13981), .ZN(n11265) );
  INV_X1 U12278 ( .A(n10730), .ZN(n10729) );
  NAND2_X1 U12279 ( .A1(n11618), .A2(n9739), .ZN(n11632) );
  INV_X1 U12280 ( .A(n11618), .ZN(n11621) );
  NOR2_X1 U12281 ( .A1(n10456), .A2(n11376), .ZN(n10455) );
  INV_X1 U12282 ( .A(n10457), .ZN(n10456) );
  NOR2_X1 U12283 ( .A1(n10344), .A2(n10343), .ZN(n10342) );
  AND2_X1 U12284 ( .A1(n9727), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10350) );
  INV_X1 U12285 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17126) );
  INV_X1 U12286 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11579) );
  INV_X1 U12287 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13332) );
  NAND2_X1 U12288 ( .A1(n9760), .A2(n10178), .ZN(n10177) );
  INV_X1 U12289 ( .A(n15421), .ZN(n10178) );
  OR2_X1 U12290 ( .A1(n17362), .A2(n11483), .ZN(n10310) );
  AND2_X1 U12291 ( .A1(n10409), .A2(n11485), .ZN(n9911) );
  INV_X1 U12292 ( .A(n14900), .ZN(n11478) );
  INV_X1 U12293 ( .A(n11485), .ZN(n9916) );
  NOR2_X1 U12294 ( .A1(n14919), .A2(n10311), .ZN(n12181) );
  INV_X1 U12295 ( .A(n10312), .ZN(n10311) );
  AOI21_X1 U12296 ( .B1(n17220), .B2(n14902), .A(n11564), .ZN(n10312) );
  OAI21_X1 U12297 ( .B1(n10408), .B2(n10410), .A(n14900), .ZN(n10018) );
  AND2_X1 U12298 ( .A1(n9805), .A2(n10211), .ZN(n10210) );
  OR2_X1 U12299 ( .A1(n14889), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10211) );
  INV_X1 U12300 ( .A(n14794), .ZN(n10425) );
  INV_X1 U12301 ( .A(n10426), .ZN(n10422) );
  AOI21_X1 U12302 ( .B1(n14815), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17362), .ZN(n14919) );
  NOR2_X1 U12303 ( .A1(n16405), .A2(n11482), .ZN(n14889) );
  NAND2_X1 U12304 ( .A1(n10071), .A2(n10487), .ZN(n10069) );
  NAND2_X1 U12305 ( .A1(n10127), .A2(n10070), .ZN(n10485) );
  NOR2_X1 U12306 ( .A1(n10071), .A2(n14885), .ZN(n10070) );
  INV_X1 U12307 ( .A(n10428), .ZN(n10553) );
  NAND2_X1 U12308 ( .A1(n9804), .A2(n10412), .ZN(n10223) );
  NAND2_X1 U12309 ( .A1(n10411), .A2(n10213), .ZN(n10212) );
  INV_X1 U12310 ( .A(n16823), .ZN(n10394) );
  AOI21_X1 U12311 ( .B1(n10414), .B2(n9804), .A(n10413), .ZN(n10473) );
  INV_X1 U12312 ( .A(n11422), .ZN(n10414) );
  AND2_X1 U12313 ( .A1(n10419), .A2(n14865), .ZN(n10418) );
  AND2_X1 U12314 ( .A1(n11497), .A2(n11496), .ZN(n16502) );
  NAND2_X1 U12315 ( .A1(n10399), .A2(n14840), .ZN(n10398) );
  NAND2_X1 U12316 ( .A1(n14839), .A2(n16535), .ZN(n16534) );
  NOR2_X1 U12317 ( .A1(n11021), .A2(n17277), .ZN(n16989) );
  AND2_X1 U12318 ( .A1(n11358), .A2(n11357), .ZN(n14846) );
  INV_X1 U12319 ( .A(n16756), .ZN(n11143) );
  OR2_X1 U12320 ( .A1(n11005), .A2(n10458), .ZN(n17017) );
  INV_X1 U12321 ( .A(n17026), .ZN(n10436) );
  AND2_X1 U12322 ( .A1(n10438), .A2(n17027), .ZN(n10437) );
  AOI21_X1 U12323 ( .B1(n10441), .B2(n10440), .A(n10439), .ZN(n10438) );
  INV_X1 U12324 ( .A(n17039), .ZN(n10439) );
  AND2_X1 U12325 ( .A1(n10997), .A2(n10440), .ZN(n10049) );
  INV_X1 U12326 ( .A(n11426), .ZN(n10441) );
  NOR2_X1 U12327 ( .A1(n17046), .A2(n11433), .ZN(n10997) );
  CLKBUF_X1 U12328 ( .A(n14425), .Z(n14562) );
  AOI21_X1 U12329 ( .B1(n11422), .B2(n17049), .A(n17048), .ZN(n17064) );
  AND2_X1 U12330 ( .A1(n11119), .A2(n9762), .ZN(n10417) );
  NAND2_X1 U12331 ( .A1(n11422), .A2(n17080), .ZN(n17125) );
  NAND2_X1 U12332 ( .A1(n10313), .A2(n10315), .ZN(n17404) );
  AND2_X1 U12333 ( .A1(n11404), .A2(n10314), .ZN(n10313) );
  NAND2_X1 U12334 ( .A1(n17142), .A2(n17146), .ZN(n11078) );
  AND3_X1 U12335 ( .A1(n11240), .A2(n11239), .A3(n11238), .ZN(n16886) );
  INV_X1 U12336 ( .A(n17161), .ZN(n11107) );
  INV_X1 U12337 ( .A(n10475), .ZN(n9917) );
  AOI21_X1 U12338 ( .B1(n10479), .B2(n10477), .A(n10476), .ZN(n10475) );
  AOI21_X1 U12339 ( .B1(n14828), .B2(n14276), .A(n14281), .ZN(n10180) );
  OAI211_X1 U12340 ( .C1(n11361), .C2(n20071), .A(n11210), .B(n11209), .ZN(
        n13921) );
  NAND2_X1 U12341 ( .A1(n13909), .A2(n13908), .ZN(n13911) );
  NAND2_X1 U12342 ( .A1(n12215), .A2(n17491), .ZN(n12237) );
  INV_X1 U12343 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14358) );
  NAND2_X1 U12344 ( .A1(n10719), .A2(n17495), .ZN(n11393) );
  AND2_X1 U12345 ( .A1(n14249), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13774) );
  INV_X1 U12346 ( .A(n12222), .ZN(n13772) );
  CLKBUF_X1 U12347 ( .A(n11184), .Z(n11185) );
  CLKBUF_X1 U12348 ( .A(n10812), .Z(n10909) );
  INV_X1 U12349 ( .A(n20629), .ZN(n20913) );
  NAND2_X1 U12350 ( .A1(n20324), .A2(n17499), .ZN(n20424) );
  OR2_X1 U12351 ( .A1(n20324), .A2(n20944), .ZN(n20650) );
  NOR2_X1 U12352 ( .A1(n20650), .A2(n20695), .ZN(n20656) );
  OR2_X1 U12353 ( .A1(n20324), .A2(n17499), .ZN(n20628) );
  NOR2_X2 U12354 ( .A1(n17490), .A2(n17489), .ZN(n20314) );
  NOR2_X2 U12355 ( .A1(n17488), .A2(n17489), .ZN(n20315) );
  CLKBUF_X1 U12356 ( .A(n13912), .Z(n13913) );
  OR2_X1 U12357 ( .A1(n20650), .A2(n20506), .ZN(n17509) );
  NAND2_X1 U12358 ( .A1(n11180), .A2(n11051), .ZN(n14388) );
  NOR2_X1 U12359 ( .A1(n14351), .A2(n14350), .ZN(n14803) );
  NAND2_X1 U12360 ( .A1(n12147), .A2(n12146), .ZN(n19883) );
  NAND2_X1 U12361 ( .A1(n12078), .A2(n12077), .ZN(n19870) );
  OR2_X1 U12362 ( .A1(n19387), .A2(n13368), .ZN(n12078) );
  NOR2_X1 U12363 ( .A1(n18090), .A2(n18092), .ZN(n18091) );
  NOR2_X1 U12364 ( .A1(n18113), .A2(n18114), .ZN(n18112) );
  NAND2_X1 U12365 ( .A1(n18135), .A2(n18140), .ZN(n18123) );
  INV_X1 U12366 ( .A(n18796), .ZN(n10284) );
  NOR2_X1 U12367 ( .A1(n18161), .A2(P3_EBX_REG_24__SCAN_IN), .ZN(n18135) );
  NOR2_X1 U12368 ( .A1(n18150), .A2(n18339), .ZN(n18133) );
  NOR2_X1 U12369 ( .A1(n18133), .A2(n18134), .ZN(n18132) );
  NOR2_X1 U12370 ( .A1(n18167), .A2(n18339), .ZN(n18158) );
  NOR2_X1 U12371 ( .A1(n18158), .A2(n18833), .ZN(n18157) );
  INV_X1 U12372 ( .A(n10249), .ZN(n13394) );
  INV_X1 U12373 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n10247) );
  NOR2_X1 U12374 ( .A1(n18227), .A2(n10252), .ZN(n10251) );
  INV_X1 U12375 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n10252) );
  NOR2_X1 U12376 ( .A1(n18686), .A2(n18688), .ZN(n10078) );
  AND2_X1 U12377 ( .A1(n17797), .A2(n11687), .ZN(n9867) );
  OR2_X1 U12378 ( .A1(n11761), .A2(n11760), .ZN(n12083) );
  AOI22_X1 U12379 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11815) );
  NOR2_X1 U12380 ( .A1(n14235), .A2(n19934), .ZN(n18679) );
  NAND3_X1 U12381 ( .A1(n12074), .A2(n12038), .A3(n12037), .ZN(n18745) );
  NOR2_X1 U12382 ( .A1(n10081), .A2(n19443), .ZN(n12037) );
  INV_X1 U12383 ( .A(n18339), .ZN(n18406) );
  NAND2_X1 U12384 ( .A1(n12118), .A2(n9731), .ZN(n17572) );
  AND2_X1 U12385 ( .A1(n12118), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18058) );
  NAND2_X1 U12386 ( .A1(n18908), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18890) );
  INV_X1 U12387 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18987) );
  NAND2_X1 U12388 ( .A1(n10286), .A2(n10287), .ZN(n14574) );
  NOR2_X1 U12389 ( .A1(n19068), .A2(n10288), .ZN(n10287) );
  INV_X1 U12390 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10288) );
  AND2_X1 U12391 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n19080) );
  NAND2_X1 U12392 ( .A1(n12168), .A2(n10074), .ZN(n10073) );
  NAND2_X1 U12393 ( .A1(n18966), .A2(n13381), .ZN(n10298) );
  NAND2_X1 U12394 ( .A1(n10026), .A2(n9862), .ZN(n17565) );
  OAI21_X1 U12395 ( .B1(n17644), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11866), .ZN(n10026) );
  AND2_X1 U12396 ( .A1(n18807), .A2(n17566), .ZN(n17639) );
  NAND2_X1 U12397 ( .A1(n10302), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10300) );
  NAND2_X1 U12398 ( .A1(n18966), .A2(n19140), .ZN(n10076) );
  NAND2_X1 U12399 ( .A1(n18816), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10077) );
  INV_X1 U12400 ( .A(n10152), .ZN(n10301) );
  INV_X1 U12401 ( .A(n19230), .ZN(n18807) );
  OR2_X1 U12403 ( .A1(n11856), .A2(n19157), .ZN(n11857) );
  CLKBUF_X1 U12404 ( .A(n18951), .Z(n18963) );
  INV_X1 U12405 ( .A(n19382), .ZN(n19876) );
  AND2_X1 U12406 ( .A1(n18994), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n19281) );
  INV_X1 U12407 ( .A(n18950), .ZN(n18966) );
  NAND2_X1 U12408 ( .A1(n19055), .A2(n12104), .ZN(n19040) );
  INV_X1 U12409 ( .A(n12102), .ZN(n10106) );
  NAND2_X1 U12410 ( .A1(n19056), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19055) );
  XNOR2_X1 U12411 ( .A(n12098), .B(n10102), .ZN(n19082) );
  INV_X1 U12412 ( .A(n12099), .ZN(n10102) );
  NAND2_X1 U12413 ( .A1(n19105), .A2(n12096), .ZN(n19090) );
  NAND2_X1 U12414 ( .A1(n19090), .A2(n19091), .ZN(n19089) );
  AND2_X1 U12415 ( .A1(n12045), .A2(n12040), .ZN(n13362) );
  INV_X1 U12416 ( .A(n19879), .ZN(n19391) );
  INV_X1 U12417 ( .A(n13537), .ZN(n13529) );
  OR2_X1 U12418 ( .A1(n20046), .A2(n13367), .ZN(n19382) );
  NOR2_X1 U12419 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19414), .ZN(n19765) );
  OR2_X1 U12420 ( .A1(n12019), .A2(n12018), .ZN(n19431) );
  INV_X1 U12421 ( .A(n19765), .ZN(n19455) );
  AOI21_X1 U12422 ( .B1(n15468), .B2(n9700), .A(n13115), .ZN(n13118) );
  NAND2_X1 U12423 ( .A1(n15595), .A2(n10038), .ZN(n10032) );
  NAND2_X1 U12424 ( .A1(n13584), .A2(n12992), .ZN(n13802) );
  INV_X1 U12425 ( .A(n21111), .ZN(n15821) );
  NAND2_X1 U12426 ( .A1(n13499), .A2(n13498), .ZN(n21116) );
  OR2_X1 U12427 ( .A1(n13620), .A2(n13497), .ZN(n13498) );
  INV_X1 U12429 ( .A(n15822), .ZN(n15872) );
  NOR2_X1 U12430 ( .A1(n15889), .A2(n13623), .ZN(n15890) );
  OR2_X1 U12431 ( .A1(n13620), .A2(n13619), .ZN(n13621) );
  NAND2_X1 U12432 ( .A1(n13758), .A2(n13618), .ZN(n13622) );
  INV_X1 U12433 ( .A(n15890), .ZN(n15901) );
  AND2_X1 U12434 ( .A1(n13414), .A2(n17847), .ZN(n21132) );
  NAND2_X1 U12435 ( .A1(n10032), .A2(n10033), .ZN(n15985) );
  NAND2_X1 U12436 ( .A1(n13883), .A2(n14320), .ZN(n13886) );
  INV_X1 U12437 ( .A(n17877), .ZN(n17880) );
  XNOR2_X1 U12438 ( .A(n9936), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16145) );
  OAI21_X1 U12439 ( .B1(n15927), .B2(n12891), .A(n9883), .ZN(n9936) );
  NAND2_X1 U12440 ( .A1(n15927), .A2(n10199), .ZN(n9883) );
  NOR2_X1 U12441 ( .A1(n16103), .A2(n10497), .ZN(n10199) );
  NAND2_X1 U12442 ( .A1(n10150), .A2(n10141), .ZN(n10149) );
  NAND2_X1 U12443 ( .A1(n15927), .A2(n10146), .ZN(n10145) );
  AND2_X1 U12444 ( .A1(n16259), .A2(n13171), .ZN(n10255) );
  OAI21_X1 U12445 ( .B1(n15975), .B2(n12882), .A(n16103), .ZN(n15978) );
  NAND2_X1 U12446 ( .A1(n10239), .A2(n10238), .ZN(n15990) );
  NAND2_X1 U12447 ( .A1(n15996), .A2(n16224), .ZN(n10238) );
  NAND2_X1 U12448 ( .A1(n15997), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10239) );
  INV_X1 U12449 ( .A(n10256), .ZN(n16221) );
  OR2_X1 U12450 ( .A1(n17886), .A2(n13799), .ZN(n16301) );
  OR2_X1 U12451 ( .A1(n13523), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17899) );
  NAND2_X1 U12452 ( .A1(n10277), .A2(n17872), .ZN(n17864) );
  INV_X1 U12453 ( .A(n21175), .ZN(n17907) );
  NAND2_X1 U12454 ( .A1(n10505), .A2(n12708), .ZN(n10276) );
  NAND2_X1 U12455 ( .A1(n10012), .A2(n14441), .ZN(n10011) );
  OAI21_X1 U12456 ( .B1(n14315), .B2(n17932), .A(n21189), .ZN(n21747) );
  NOR2_X1 U12457 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21733) );
  OAI221_X1 U12458 ( .B1(n21586), .B2(n21501), .C1(n21584), .C2(n21500), .A(
        n21582), .ZN(n21519) );
  INV_X1 U12459 ( .A(n21291), .ZN(n21578) );
  INV_X1 U12460 ( .A(n21304), .ZN(n21592) );
  INV_X1 U12461 ( .A(n21308), .ZN(n21598) );
  INV_X1 U12462 ( .A(n21312), .ZN(n21604) );
  INV_X1 U12463 ( .A(n21316), .ZN(n21610) );
  INV_X1 U12464 ( .A(n21320), .ZN(n21616) );
  INV_X1 U12465 ( .A(n21324), .ZN(n21622) );
  INV_X1 U12466 ( .A(n21328), .ZN(n21630) );
  AOI221_X1 U12467 ( .B1(n21638), .B2(n13237), .C1(n17853), .C2(n13237), .A(
        n17930), .ZN(n17855) );
  AND2_X1 U12468 ( .A1(n13237), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17854) );
  INV_X1 U12469 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21530) );
  INV_X1 U12470 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21657) );
  INV_X1 U12471 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n21666) );
  INV_X1 U12472 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n21672) );
  OR2_X1 U12474 ( .A1(n11458), .A2(n11472), .ZN(n16405) );
  AND2_X1 U12475 ( .A1(n11463), .A2(n11457), .ZN(n11458) );
  NAND2_X1 U12476 ( .A1(n10332), .A2(n10336), .ZN(n16400) );
  NAND2_X1 U12477 ( .A1(n16414), .A2(n10322), .ZN(n10332) );
  AOI21_X1 U12478 ( .B1(n16414), .B2(n10322), .A(n16415), .ZN(n16397) );
  NAND2_X1 U12479 ( .A1(n11023), .A2(n9895), .ZN(n9894) );
  AND2_X1 U12480 ( .A1(n11473), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n9895) );
  NAND2_X1 U12481 ( .A1(n16529), .A2(n16993), .ZN(n16515) );
  NAND2_X1 U12482 ( .A1(n10322), .A2(n11607), .ZN(n16529) );
  AND2_X1 U12483 ( .A1(n10988), .A2(n9725), .ZN(n11008) );
  OR2_X1 U12484 ( .A1(n20053), .A2(n11656), .ZN(n20180) );
  INV_X1 U12485 ( .A(n20182), .ZN(n20169) );
  NOR2_X1 U12486 ( .A1(n9900), .A2(n9899), .ZN(n10939) );
  INV_X1 U12487 ( .A(n10935), .ZN(n9900) );
  AND2_X1 U12488 ( .A1(n20053), .A2(n14403), .ZN(n20185) );
  INV_X1 U12489 ( .A(n20185), .ZN(n20171) );
  AND2_X1 U12490 ( .A1(n13213), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20197) );
  INV_X1 U12491 ( .A(n20189), .ZN(n20129) );
  INV_X1 U12492 ( .A(n20145), .ZN(n20186) );
  NAND2_X1 U12493 ( .A1(n10322), .A2(n20197), .ZN(n16649) );
  CLKBUF_X1 U12494 ( .A(n15429), .Z(n15430) );
  OR2_X1 U12495 ( .A1(n11315), .A2(n11314), .ZN(n14595) );
  OR2_X1 U12496 ( .A1(n11289), .A2(n11288), .ZN(n14422) );
  CLKBUF_X1 U12497 ( .A(n20207), .Z(n16760) );
  INV_X1 U12498 ( .A(n20944), .ZN(n17499) );
  NAND2_X1 U12499 ( .A1(n10464), .A2(n10467), .ZN(n10461) );
  NOR2_X2 U12500 ( .A1(n20226), .A2(n12207), .ZN(n16875) );
  NAND2_X1 U12501 ( .A1(n12206), .A2(n17488), .ZN(n16878) );
  INV_X1 U12502 ( .A(n10380), .ZN(n13978) );
  AOI21_X1 U12503 ( .B1(n10386), .B2(n10384), .A(n9709), .ZN(n10380) );
  NAND2_X1 U12504 ( .A1(n14777), .A2(n10387), .ZN(n10386) );
  INV_X2 U12505 ( .A(n16897), .ZN(n20226) );
  INV_X1 U12506 ( .A(n20271), .ZN(n20240) );
  OAI21_X1 U12507 ( .B1(n14349), .B2(n13388), .A(n13387), .ZN(n20260) );
  INV_X1 U12508 ( .A(n20260), .ZN(n20276) );
  AOI21_X1 U12509 ( .B1(n16733), .B2(n17182), .A(n11161), .ZN(n11162) );
  NAND2_X1 U12510 ( .A1(n17033), .A2(n10455), .ZN(n17002) );
  INV_X1 U12511 ( .A(n14834), .ZN(n17003) );
  INV_X1 U12512 ( .A(n17166), .ZN(n17182) );
  INV_X1 U12513 ( .A(n17181), .ZN(n17193) );
  NAND2_X1 U12514 ( .A1(n14916), .A2(n14915), .ZN(n16402) );
  NAND2_X1 U12515 ( .A1(n16929), .A2(n16937), .ZN(n16920) );
  NAND2_X1 U12516 ( .A1(n16965), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16956) );
  NOR2_X1 U12517 ( .A1(n16966), .A2(n9783), .ZN(n14881) );
  AOI21_X1 U12518 ( .B1(n16975), .B2(n14857), .A(n9825), .ZN(n14861) );
  INV_X1 U12519 ( .A(n10187), .ZN(n16979) );
  AND2_X1 U12520 ( .A1(n16975), .A2(n16974), .ZN(n16978) );
  XNOR2_X1 U12521 ( .A(n11030), .B(n10537), .ZN(n11421) );
  NOR2_X1 U12522 ( .A1(n11022), .A2(n16988), .ZN(n11030) );
  NAND2_X1 U12523 ( .A1(n10058), .A2(n10063), .ZN(n11022) );
  AOI21_X1 U12524 ( .B1(n17033), .B2(n9832), .A(n9716), .ZN(n14849) );
  INV_X1 U12525 ( .A(n14843), .ZN(n10207) );
  NAND2_X1 U12526 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n11376), .ZN(
        n10208) );
  NAND2_X1 U12527 ( .A1(n10064), .A2(n11435), .ZN(n14825) );
  OR2_X1 U12528 ( .A1(n14852), .A2(n11012), .ZN(n10064) );
  AOI21_X1 U12529 ( .B1(n14834), .B2(n14833), .A(n14832), .ZN(n14856) );
  NAND2_X1 U12530 ( .A1(n9716), .A2(n17007), .ZN(n10169) );
  AND2_X1 U12531 ( .A1(n9832), .A2(n17007), .ZN(n10170) );
  NOR2_X1 U12532 ( .A1(n17074), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10021) );
  NAND4_X1 U12533 ( .A1(n10314), .A2(n11404), .A3(n9792), .A4(n10315), .ZN(
        n17378) );
  INV_X1 U12534 ( .A(n17105), .ZN(n17106) );
  INV_X1 U12535 ( .A(n17458), .ZN(n17412) );
  OR2_X1 U12536 ( .A1(n14777), .A2(n14778), .ZN(n10383) );
  AND2_X1 U12537 ( .A1(n10446), .A2(n10445), .ZN(n17143) );
  AND2_X1 U12538 ( .A1(n10315), .A2(n10314), .ZN(n17431) );
  NAND2_X1 U12539 ( .A1(n17177), .A2(n11071), .ZN(n17160) );
  NAND2_X1 U12540 ( .A1(n13903), .A2(n11231), .ZN(n16599) );
  OAI21_X1 U12541 ( .B1(n10872), .B2(n10484), .A(n10482), .ZN(n17169) );
  INV_X1 U12542 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20920) );
  NAND2_X1 U12543 ( .A1(n13904), .A2(n13907), .ZN(n20931) );
  NAND2_X1 U12544 ( .A1(n13899), .A2(n13898), .ZN(n20921) );
  NAND2_X1 U12545 ( .A1(n13897), .A2(n13896), .ZN(n13898) );
  NOR2_X1 U12546 ( .A1(n20562), .A2(n20424), .ZN(n20346) );
  INV_X1 U12547 ( .A(n20339), .ZN(n20352) );
  OAI21_X1 U12548 ( .B1(n20396), .B2(n20395), .A(n20394), .ZN(n20413) );
  INV_X1 U12549 ( .A(n20443), .ZN(n20446) );
  OAI21_X1 U12550 ( .B1(n20563), .B2(n20423), .A(n20422), .ZN(n20445) );
  OAI21_X1 U12551 ( .B1(n20459), .B2(n20458), .A(n20457), .ZN(n20477) );
  AOI21_X1 U12552 ( .B1(n20939), .B2(n17494), .A(n17493), .ZN(n20496) );
  OR2_X1 U12553 ( .A1(n20500), .A2(n20695), .ZN(n17480) );
  OAI21_X1 U12554 ( .B1(n20916), .B2(n20513), .A(n20512), .ZN(n20530) );
  NAND2_X1 U12555 ( .A1(n20502), .A2(n20501), .ZN(n20555) );
  AOI21_X1 U12556 ( .B1(n9798), .B2(n9954), .A(n9949), .ZN(n20535) );
  INV_X1 U12557 ( .A(n9955), .ZN(n9949) );
  NAND2_X1 U12558 ( .A1(n9954), .A2(n9950), .ZN(n20540) );
  OAI21_X1 U12559 ( .B1(n20571), .B2(n20570), .A(n20569), .ZN(n20588) );
  OAI21_X1 U12560 ( .B1(n20654), .B2(n20658), .A(n20653), .ZN(n20683) );
  AND2_X1 U12561 ( .A1(n20696), .A2(n20690), .ZN(n20721) );
  OR2_X1 U12562 ( .A1(n20628), .A2(n20695), .ZN(n17507) );
  INV_X1 U12563 ( .A(n20666), .ZN(n20728) );
  OAI21_X1 U12564 ( .B1(n17502), .B2(n17505), .A(n17501), .ZN(n20748) );
  INV_X1 U12565 ( .A(n20701), .ZN(n20757) );
  INV_X1 U12566 ( .A(n20669), .ZN(n20766) );
  INV_X1 U12567 ( .A(n20707), .ZN(n20767) );
  INV_X1 U12568 ( .A(n20672), .ZN(n20777) );
  INV_X1 U12569 ( .A(n20713), .ZN(n20787) );
  OR2_X1 U12570 ( .A1(n17521), .A2(n17520), .ZN(n20816) );
  INV_X1 U12571 ( .A(n20678), .ZN(n20797) );
  INV_X1 U12572 ( .A(n20681), .ZN(n20807) );
  INV_X1 U12573 ( .A(n20285), .ZN(n20819) );
  NOR2_X1 U12574 ( .A1(n14407), .A2(n14413), .ZN(n14504) );
  NAND2_X1 U12575 ( .A1(n20051), .A2(n18681), .ZN(n20049) );
  XNOR2_X1 U12576 ( .A(n19420), .B(n18681), .ZN(n20046) );
  INV_X1 U12577 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n20035) );
  NOR2_X1 U12578 ( .A1(n18123), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n18122) );
  NAND2_X1 U12579 ( .A1(n18122), .A2(n18447), .ZN(n18118) );
  NOR2_X1 U12580 ( .A1(n18204), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n18191) );
  NAND2_X1 U12581 ( .A1(n18191), .A2(n18537), .ZN(n18185) );
  NOR2_X1 U12582 ( .A1(n18189), .A2(n18339), .ZN(n18180) );
  NOR2_X1 U12583 ( .A1(n18180), .A2(n18181), .ZN(n18179) );
  NOR2_X1 U12584 ( .A1(n18339), .A2(n18061), .ZN(n18190) );
  NOR2_X1 U12585 ( .A1(n18190), .A2(n18873), .ZN(n18189) );
  NAND2_X1 U12586 ( .A1(n18210), .A2(n18205), .ZN(n18204) );
  NOR2_X1 U12587 ( .A1(n18226), .A2(P3_EBX_REG_18__SCAN_IN), .ZN(n18210) );
  NOR2_X1 U12588 ( .A1(n18282), .A2(P3_EBX_REG_14__SCAN_IN), .ZN(n18259) );
  NAND2_X1 U12589 ( .A1(n18259), .A2(n18258), .ZN(n18255) );
  NAND2_X1 U12590 ( .A1(n18287), .A2(n18285), .ZN(n18282) );
  NOR2_X1 U12591 ( .A1(n18306), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n18287) );
  NOR2_X1 U12592 ( .A1(n18381), .A2(P3_EBX_REG_6__SCAN_IN), .ZN(n18366) );
  NAND2_X1 U12593 ( .A1(n18366), .A2(n18564), .ZN(n18359) );
  INV_X1 U12594 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n18382) );
  NAND2_X1 U12595 ( .A1(n18387), .A2(n18382), .ZN(n18381) );
  NOR2_X1 U12596 ( .A1(n18415), .A2(P3_EBX_REG_4__SCAN_IN), .ZN(n18387) );
  INV_X1 U12597 ( .A(n18435), .ZN(n18402) );
  AND3_X1 U12598 ( .A1(n9879), .A2(n9878), .A3(n9877), .ZN(n18419) );
  INV_X1 U12599 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n9879) );
  NOR2_X2 U12600 ( .A1(n20049), .A2(n19903), .ZN(n18432) );
  NOR2_X1 U12601 ( .A1(n14236), .A2(n20051), .ZN(n18385) );
  NOR2_X1 U12602 ( .A1(n18447), .A2(n10247), .ZN(n10244) );
  NOR2_X1 U12603 ( .A1(n18172), .A2(n17679), .ZN(n18511) );
  NAND2_X1 U12604 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17549), .ZN(n18533) );
  AND2_X1 U12605 ( .A1(n13890), .A2(n10250), .ZN(n17549) );
  AND2_X1 U12606 ( .A1(n9744), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U12607 ( .A1(n13890), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n14485) );
  NAND4_X1 U12608 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .A4(n13720), .ZN(n13721) );
  AND2_X1 U12609 ( .A1(n13359), .A2(n10240), .ZN(n13720) );
  NOR2_X1 U12610 ( .A1(n18307), .A2(n10242), .ZN(n10240) );
  NOR2_X1 U12611 ( .A1(n18573), .A2(n18382), .ZN(n18569) );
  AND2_X1 U12612 ( .A1(n18587), .A2(n10254), .ZN(n18574) );
  INV_X1 U12613 ( .A(n18578), .ZN(n10254) );
  NAND2_X1 U12614 ( .A1(n18574), .A2(P3_EBX_REG_4__SCAN_IN), .ZN(n18573) );
  INV_X1 U12615 ( .A(n18602), .ZN(n18598) );
  NAND2_X1 U12616 ( .A1(n18614), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n18610) );
  NOR2_X1 U12617 ( .A1(n18690), .A2(n18619), .ZN(n18614) );
  INV_X1 U12618 ( .A(n18624), .ZN(n18620) );
  NOR2_X1 U12619 ( .A1(n18594), .A2(n10079), .ZN(n18630) );
  NAND2_X1 U12620 ( .A1(n10080), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n10079) );
  INV_X1 U12621 ( .A(n18634), .ZN(n10080) );
  NAND2_X1 U12622 ( .A1(n18630), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n18629) );
  NOR2_X1 U12623 ( .A1(n18661), .A2(n18794), .ZN(n13545) );
  NAND2_X1 U12624 ( .A1(n13545), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n18594) );
  NOR2_X1 U12625 ( .A1(n18662), .A2(n13434), .ZN(n18674) );
  INV_X1 U12626 ( .A(n18662), .ZN(n18677) );
  AND4_X1 U12627 ( .A1(n11735), .A2(n11734), .A3(n11733), .A4(n11732), .ZN(
        n11747) );
  AND4_X1 U12628 ( .A1(n11707), .A2(n11706), .A3(n11705), .A4(n11704), .ZN(
        n11713) );
  INV_X1 U12629 ( .A(n18636), .ZN(n13488) );
  NAND2_X1 U12630 ( .A1(n10082), .A2(n20038), .ZN(n13457) );
  NAND2_X1 U12631 ( .A1(n10083), .A2(n9845), .ZN(n10082) );
  NAND2_X1 U12632 ( .A1(n13429), .A2(n10084), .ZN(n10083) );
  INV_X1 U12633 ( .A(n18638), .ZN(n18673) );
  INV_X1 U12634 ( .A(n18674), .ZN(n13793) );
  NAND2_X1 U12635 ( .A1(n18742), .A2(n18679), .ZN(n18736) );
  INV_X1 U12636 ( .A(n18736), .ZN(n18738) );
  NOR2_X1 U12637 ( .A1(n18790), .A2(n19420), .ZN(n18791) );
  INV_X1 U12638 ( .A(n18924), .ZN(n18891) );
  INV_X1 U12639 ( .A(n18849), .ZN(n10293) );
  AND2_X1 U12640 ( .A1(n18908), .A2(n10294), .ZN(n18869) );
  NAND2_X1 U12641 ( .A1(n19043), .A2(n9758), .ZN(n14569) );
  INV_X1 U12642 ( .A(n19636), .ZN(n19801) );
  NOR2_X1 U12643 ( .A1(n19069), .A2(n19068), .ZN(n19054) );
  INV_X1 U12644 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n19095) );
  NAND2_X1 U12645 ( .A1(n19765), .A2(n19408), .ZN(n19636) );
  NAND2_X1 U12646 ( .A1(n18985), .A2(n18868), .ZN(n19122) );
  INV_X1 U12647 ( .A(n19121), .ZN(n19112) );
  INV_X1 U12648 ( .A(n11866), .ZN(n17633) );
  NAND2_X1 U12649 ( .A1(n18830), .A2(n11862), .ZN(n17597) );
  AOI21_X1 U12650 ( .B1(n19186), .B2(n9840), .A(n19302), .ZN(n19193) );
  AOI21_X1 U12651 ( .B1(n19230), .B2(n19875), .A(n9778), .ZN(n19223) );
  NOR2_X1 U12652 ( .A1(n19234), .A2(n19197), .ZN(n19273) );
  AND2_X1 U12653 ( .A1(n19370), .A2(n17632), .ZN(n19297) );
  INV_X1 U12654 ( .A(n13371), .ZN(n12047) );
  NAND2_X1 U12655 ( .A1(n19067), .A2(n11837), .ZN(n19050) );
  NAND2_X1 U12656 ( .A1(n9857), .A2(n9974), .ZN(n19075) );
  OR2_X1 U12657 ( .A1(n12155), .A2(n12154), .ZN(n19341) );
  AND2_X1 U12658 ( .A1(n19341), .A2(n19391), .ZN(n19370) );
  INV_X1 U12659 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19409) );
  INV_X1 U12660 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19890) );
  OR2_X1 U12661 ( .A1(n19902), .A2(n19901), .ZN(n19904) );
  INV_X1 U12662 ( .A(n20038), .ZN(n19914) );
  NOR2_X1 U12663 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20016), .ZN(
        n19909) );
  INV_X1 U12664 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n20016) );
  AND2_X2 U12665 ( .A1(n13186), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n15837)
         );
  CLKBUF_X1 U12666 ( .A(n18016), .Z(n18025) );
  NOR2_X1 U12667 ( .A1(n17987), .A2(n17936), .ZN(n17992) );
  AND2_X1 U12668 ( .A1(n14789), .A2(n16937), .ZN(n14791) );
  NAND2_X1 U12669 ( .A1(n10127), .A2(n10492), .ZN(n10491) );
  NAND2_X1 U12670 ( .A1(n10037), .A2(n10035), .ZN(P1_U2850) );
  INV_X1 U12671 ( .A(n10036), .ZN(n10035) );
  NAND2_X1 U12672 ( .A1(n10032), .A2(n9774), .ZN(n10037) );
  OAI22_X1 U12673 ( .A1(n16208), .A2(n15821), .B1(n15805), .B2(n21116), .ZN(
        n10036) );
  AOI21_X1 U12674 ( .B1(n15447), .B2(n10364), .A(n10362), .ZN(n10361) );
  NAND2_X1 U12675 ( .A1(n10371), .A2(n10363), .ZN(n10362) );
  OAI21_X1 U12676 ( .B1(n16085), .B2(n16117), .A(n9796), .ZN(P1_U2987) );
  NOR2_X1 U12677 ( .A1(n16089), .A2(n16088), .ZN(n10134) );
  OR2_X1 U12678 ( .A1(n16311), .A2(n20989), .ZN(n10135) );
  NOR2_X1 U12679 ( .A1(n16130), .A2(n10264), .ZN(n16132) );
  OR2_X1 U12680 ( .A1(n16916), .A2(n20189), .ZN(n12507) );
  AOI211_X1 U12681 ( .C1(n20187), .C2(n12504), .A(n12503), .B(n12502), .ZN(
        n12508) );
  OAI21_X1 U12682 ( .B1(n15428), .B2(n17181), .A(n15427), .ZN(P2_U2983) );
  AOI21_X1 U12683 ( .B1(n16908), .B2(n17196), .A(n16907), .ZN(n16909) );
  AND2_X1 U12684 ( .A1(n9967), .A2(n9966), .ZN(n16918) );
  INV_X1 U12685 ( .A(n9991), .ZN(n14799) );
  OAI211_X1 U12686 ( .C1(n14812), .C2(n17139), .A(n14797), .B(n9992), .ZN(
        n9991) );
  AOI21_X1 U12687 ( .B1(n10027), .B2(n17196), .A(n16954), .ZN(n16955) );
  OAI21_X1 U12688 ( .B1(n10112), .B2(n9723), .A(n10116), .ZN(n10027) );
  AND3_X1 U12689 ( .A1(n11569), .A2(n11568), .A3(n11567), .ZN(n11570) );
  NAND2_X1 U12690 ( .A1(n16908), .A2(n17454), .ZN(n12185) );
  INV_X1 U12691 ( .A(n12184), .ZN(n12186) );
  INV_X1 U12692 ( .A(n14910), .ZN(n14912) );
  NOR2_X1 U12693 ( .A1(n10185), .A2(n14821), .ZN(n10184) );
  AND3_X1 U12694 ( .A1(n10115), .A2(n10114), .A3(n9806), .ZN(n17238) );
  NAND2_X1 U12695 ( .A1(n9933), .A2(n9734), .ZN(n10115) );
  OAI211_X1 U12696 ( .C1(n17006), .C2(n17458), .A(n10205), .B(n10204), .ZN(
        P2_U3029) );
  INV_X1 U12697 ( .A(n10206), .ZN(n10205) );
  NAND2_X1 U12698 ( .A1(n14844), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10204) );
  OAI21_X1 U12699 ( .B1(n14849), .B2(n10208), .A(n10207), .ZN(n10206) );
  NOR2_X1 U12700 ( .A1(n17295), .A2(n17415), .ZN(n17296) );
  OAI211_X1 U12701 ( .C1(n17379), .C2(n17458), .A(n10046), .B(n10045), .ZN(
        P2_U3037) );
  NOR2_X1 U12702 ( .A1(n17377), .A2(n10047), .ZN(n10046) );
  NAND2_X1 U12703 ( .A1(n17376), .A2(n17454), .ZN(n10045) );
  AND2_X1 U12704 ( .A1(n17378), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10047) );
  OR2_X1 U12705 ( .A1(n18096), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9882) );
  AOI21_X1 U12706 ( .B1(n10291), .B2(n18414), .A(n10290), .ZN(n18089) );
  NAND2_X1 U12707 ( .A1(n18492), .A2(n10248), .ZN(n18491) );
  NOR2_X1 U12708 ( .A1(n18590), .A2(n18098), .ZN(n10248) );
  AND2_X1 U12709 ( .A1(n13359), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n13360) );
  INV_X1 U12710 ( .A(n18587), .ZN(n18589) );
  OAI21_X1 U12711 ( .B1(n17622), .B2(n19034), .A(n17564), .ZN(P3_U2800) );
  NAND2_X1 U12712 ( .A1(n10105), .A2(n10103), .ZN(P3_U2843) );
  NAND2_X1 U12713 ( .A1(n19193), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10105) );
  AOI21_X1 U12714 ( .B1(n19192), .B2(n19191), .A(n10104), .ZN(n10103) );
  OAI21_X1 U12715 ( .B1(n19195), .B2(n19311), .A(n19194), .ZN(n10104) );
  BUF_X1 U12716 ( .A(n13351), .Z(n17783) );
  AND3_X1 U12717 ( .A1(n10090), .A2(n9718), .A3(n14449), .ZN(n13119) );
  INV_X1 U12718 ( .A(n9933), .ZN(n16948) );
  NAND2_X1 U12719 ( .A1(n17032), .A2(n9743), .ZN(n9933) );
  NAND2_X1 U12720 ( .A1(n15270), .A2(n9754), .ZN(n15478) );
  NAND2_X1 U12721 ( .A1(n15270), .A2(n15269), .ZN(n15500) );
  NAND2_X2 U12722 ( .A1(n10306), .A2(n10307), .ZN(n11220) );
  AND2_X1 U12723 ( .A1(n9731), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9708) );
  AND2_X2 U12724 ( .A1(n11054), .A2(n14354), .ZN(n10624) );
  INV_X1 U12725 ( .A(n11225), .ZN(n11232) );
  NAND2_X1 U12726 ( .A1(n11682), .A2(n11683), .ZN(n11693) );
  NAND2_X1 U12727 ( .A1(n14250), .A2(n12251), .ZN(n14419) );
  NOR2_X1 U12728 ( .A1(n13916), .A2(n11482), .ZN(n9709) );
  NAND2_X1 U12729 ( .A1(n10391), .A2(n10390), .ZN(n9710) );
  NOR2_X1 U12730 ( .A1(n10124), .A2(n10125), .ZN(n16744) );
  NAND2_X1 U12731 ( .A1(n10391), .A2(n10392), .ZN(n13875) );
  NAND2_X1 U12732 ( .A1(n11367), .A2(n10395), .ZN(n14870) );
  INV_X2 U12733 ( .A(n12762), .ZN(n12718) );
  NAND2_X1 U12734 ( .A1(n9925), .A2(n10933), .ZN(n9711) );
  AND2_X1 U12735 ( .A1(n10227), .A2(n12869), .ZN(n9712) );
  AND2_X1 U12736 ( .A1(n10416), .A2(n14642), .ZN(n9713) );
  AND2_X1 U12737 ( .A1(n10552), .A2(n10989), .ZN(n9714) );
  AND2_X1 U12738 ( .A1(n10745), .A2(n10744), .ZN(n9715) );
  AND2_X1 U12739 ( .A1(n17291), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9716) );
  AND2_X1 U12740 ( .A1(n11367), .A2(n10396), .ZN(n14871) );
  AND4_X1 U12741 ( .A1(n11882), .A2(n11881), .A3(n11880), .A4(n11879), .ZN(
        n9717) );
  AND2_X1 U12742 ( .A1(n14464), .A2(n13500), .ZN(n9718) );
  INV_X1 U12743 ( .A(n10876), .ZN(n9887) );
  NOR2_X1 U12744 ( .A1(n16921), .A2(n10493), .ZN(n10492) );
  INV_X1 U12745 ( .A(n10492), .ZN(n10071) );
  INV_X1 U12746 ( .A(n9809), .ZN(n10878) );
  AND2_X1 U12747 ( .A1(n10764), .A2(n10768), .ZN(n9719) );
  AND2_X1 U12748 ( .A1(n12658), .A2(n10013), .ZN(n9720) );
  AND2_X1 U12749 ( .A1(n12461), .A2(n9850), .ZN(n9721) );
  AND2_X1 U12750 ( .A1(n9713), .A2(n11143), .ZN(n9722) );
  NAND2_X1 U12751 ( .A1(n13054), .A2(n13053), .ZN(n15668) );
  INV_X1 U12752 ( .A(n10481), .ZN(n10478) );
  OR2_X1 U12753 ( .A1(n10484), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10481) );
  NAND2_X1 U12754 ( .A1(n9933), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9723) );
  AND2_X1 U12755 ( .A1(n10489), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9724) );
  AND2_X1 U12756 ( .A1(n9714), .A2(n9846), .ZN(n9725) );
  AND2_X1 U12757 ( .A1(n17495), .A2(n20298), .ZN(n9726) );
  INV_X1 U12758 ( .A(n12243), .ZN(n13912) );
  AND2_X1 U12759 ( .A1(n10351), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9727) );
  OR2_X1 U12760 ( .A1(n11029), .A2(n11028), .ZN(n10128) );
  AND2_X1 U12761 ( .A1(n10518), .A2(n15654), .ZN(n9728) );
  AND2_X1 U12762 ( .A1(n10524), .A2(n13047), .ZN(n9729) );
  AND2_X1 U12763 ( .A1(n9724), .A2(n10069), .ZN(n9730) );
  NAND2_X1 U12764 ( .A1(n14611), .A2(n9762), .ZN(n14253) );
  AND2_X1 U12765 ( .A1(n12119), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9731) );
  NAND2_X1 U12766 ( .A1(n15899), .A2(n15824), .ZN(n9732) );
  OR2_X1 U12767 ( .A1(n11026), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n9733) );
  AND2_X1 U12768 ( .A1(n17454), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9734) );
  AND2_X1 U12769 ( .A1(n13054), .A2(n10518), .ZN(n15653) );
  AND2_X1 U12770 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9735) );
  AND2_X1 U12771 ( .A1(n9735), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9736) );
  AND2_X1 U12772 ( .A1(n17454), .A2(n9871), .ZN(n9737) );
  OR2_X1 U12773 ( .A1(n9733), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n9738) );
  AND2_X1 U12774 ( .A1(n9736), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9739) );
  AND2_X1 U12775 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9740) );
  INV_X1 U12776 ( .A(n9899), .ZN(n10936) );
  AND2_X1 U12777 ( .A1(n18966), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9741) );
  INV_X1 U12778 ( .A(n12493), .ZN(n10466) );
  AND2_X1 U12779 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .ZN(n9742) );
  AND2_X1 U12780 ( .A1(n14875), .A2(n9868), .ZN(n9743) );
  AND2_X1 U12781 ( .A1(n10251), .A2(P3_EBX_REG_18__SCAN_IN), .ZN(n9744) );
  INV_X1 U12782 ( .A(n14902), .ZN(n10176) );
  INV_X1 U12783 ( .A(n10181), .ZN(n17452) );
  AND2_X2 U12784 ( .A1(n12379), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10617) );
  AND2_X2 U12785 ( .A1(n12325), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10618) );
  NAND2_X1 U12786 ( .A1(n11449), .A2(n10269), .ZN(n9745) );
  BUF_X1 U12787 ( .A(n12558), .Z(n15278) );
  NAND2_X1 U12788 ( .A1(n13393), .A2(n11683), .ZN(n9746) );
  NOR2_X1 U12789 ( .A1(n10122), .A2(n10124), .ZN(n16723) );
  INV_X1 U12790 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11687) );
  AND2_X1 U12791 ( .A1(n15656), .A2(n15740), .ZN(n9747) );
  INV_X1 U12792 ( .A(n16967), .ZN(n10412) );
  NAND2_X1 U12793 ( .A1(n16744), .A2(n16745), .ZN(n16738) );
  AND2_X1 U12794 ( .A1(n10428), .A2(n10425), .ZN(n14793) );
  NAND2_X1 U12795 ( .A1(n15518), .A2(n15519), .ZN(n15502) );
  INV_X1 U12796 ( .A(n14899), .ZN(n10410) );
  AND2_X1 U12797 ( .A1(n18505), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n9748) );
  NAND2_X1 U12798 ( .A1(n11153), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11585) );
  NAND2_X1 U12799 ( .A1(n10181), .A2(n11398), .ZN(n10315) );
  INV_X1 U12800 ( .A(n12089), .ZN(n12079) );
  NAND2_X1 U12801 ( .A1(n13393), .A2(n11686), .ZN(n9749) );
  AND2_X1 U12802 ( .A1(n14469), .A2(n15395), .ZN(n9750) );
  AND4_X1 U12803 ( .A1(n12544), .A2(n12543), .A3(n12542), .A4(n12541), .ZN(
        n9751) );
  NAND2_X1 U12804 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n9752) );
  INV_X1 U12805 ( .A(n10328), .ZN(n15437) );
  OAI21_X1 U12806 ( .B1(n16442), .B2(n10331), .A(n10329), .ZN(n10328) );
  AND2_X1 U12807 ( .A1(n18614), .A2(n10078), .ZN(n9753) );
  AND2_X1 U12808 ( .A1(n10360), .A2(n15490), .ZN(n9754) );
  NAND2_X1 U12809 ( .A1(n16922), .A2(n10189), .ZN(n10190) );
  AND2_X1 U12810 ( .A1(n10444), .A2(n11435), .ZN(n9755) );
  INV_X1 U12811 ( .A(n12869), .ZN(n10164) );
  AND2_X1 U12812 ( .A1(n10294), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9757) );
  AND2_X1 U12813 ( .A1(n11846), .A2(n10305), .ZN(n9758) );
  AND2_X1 U12814 ( .A1(n12960), .A2(n12958), .ZN(n9759) );
  NAND2_X1 U12815 ( .A1(n14558), .A2(n14557), .ZN(n14646) );
  AND2_X1 U12816 ( .A1(n15537), .A2(n15536), .ZN(n15518) );
  AND2_X1 U12817 ( .A1(n14836), .A2(n10419), .ZN(n14863) );
  OR2_X1 U12818 ( .A1(n12181), .A2(n10310), .ZN(n9760) );
  AND3_X1 U12819 ( .A1(n9689), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9761) );
  NAND2_X1 U12820 ( .A1(n10009), .A2(n10162), .ZN(n16020) );
  NAND2_X1 U12821 ( .A1(n11153), .A2(n10351), .ZN(n10353) );
  AND2_X1 U12822 ( .A1(n14254), .A2(n14260), .ZN(n9762) );
  AOI21_X1 U12823 ( .B1(n11422), .B2(n10997), .A(n10441), .ZN(n17037) );
  NOR2_X1 U12824 ( .A1(n19443), .A2(n13322), .ZN(n9763) );
  NAND2_X1 U12825 ( .A1(n10431), .A2(n10438), .ZN(n17025) );
  AND2_X1 U12826 ( .A1(n10197), .A2(n10195), .ZN(n17871) );
  AND2_X1 U12827 ( .A1(n14900), .A2(n14899), .ZN(n9764) );
  AND2_X1 U12828 ( .A1(n11428), .A2(n9894), .ZN(n9765) );
  INV_X1 U12829 ( .A(n11844), .ZN(n9985) );
  NAND2_X1 U12830 ( .A1(n17866), .A2(n12861), .ZN(n16090) );
  AND4_X1 U12831 ( .A1(n11692), .A2(n11691), .A3(n11690), .A4(n11689), .ZN(
        n9766) );
  AND2_X1 U12832 ( .A1(n12743), .A2(n12789), .ZN(n9767) );
  AND3_X1 U12834 ( .A1(n11875), .A2(n11876), .A3(n11877), .ZN(n9768) );
  AND2_X1 U12835 ( .A1(n10090), .A2(n9718), .ZN(n13750) );
  NOR3_X1 U12836 ( .A1(n11664), .A2(n11482), .A3(n11564), .ZN(n9769) );
  OR3_X1 U12837 ( .A1(n17216), .A2(n11563), .A3(n14887), .ZN(n9770) );
  AND2_X1 U12838 ( .A1(n10376), .A2(n10375), .ZN(n9771) );
  NAND2_X1 U12839 ( .A1(n12737), .A2(n12736), .ZN(n12774) );
  XNOR2_X1 U12840 ( .A(n12733), .B(n12734), .ZN(n13679) );
  INV_X1 U12841 ( .A(n12652), .ZN(n10003) );
  INV_X1 U12842 ( .A(n16341), .ZN(n10529) );
  OR2_X1 U12843 ( .A1(n16425), .A2(n16424), .ZN(n9772) );
  AND2_X1 U12844 ( .A1(n12652), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9773) );
  NOR2_X1 U12845 ( .A1(n11463), .A2(n11457), .ZN(n11472) );
  AND2_X1 U12846 ( .A1(n10033), .A2(n21112), .ZN(n9774) );
  OR2_X1 U12847 ( .A1(n13159), .A2(n16137), .ZN(n9775) );
  AND4_X1 U12848 ( .A1(n10951), .A2(n10950), .A3(n10949), .A4(n10948), .ZN(
        n9776) );
  INV_X1 U12849 ( .A(n10112), .ZN(n16965) );
  AND2_X1 U12850 ( .A1(n17495), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9777) );
  AND2_X1 U12851 ( .A1(n19236), .A2(n19263), .ZN(n9778) );
  AND2_X1 U12852 ( .A1(n13389), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9779) );
  INV_X1 U12853 ( .A(n12631), .ZN(n10088) );
  AND2_X1 U12854 ( .A1(n11220), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9780) );
  OR2_X1 U12856 ( .A1(n11607), .A2(n10339), .ZN(n9781) );
  NOR2_X1 U12857 ( .A1(n11017), .A2(n11376), .ZN(n11437) );
  OR2_X1 U12858 ( .A1(n10479), .A2(n10478), .ZN(n9782) );
  AND2_X1 U12859 ( .A1(n10187), .A2(n14862), .ZN(n9783) );
  AND2_X1 U12860 ( .A1(n10237), .A2(n12844), .ZN(n9784) );
  AND2_X1 U12861 ( .A1(n9940), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9785) );
  AND3_X1 U12862 ( .A1(n17822), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n11477), .ZN(n9786) );
  AND2_X1 U12863 ( .A1(n9725), .A2(n11007), .ZN(n9787) );
  OR3_X1 U12864 ( .A1(n16131), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12892), .ZN(n9788) );
  OR2_X1 U12865 ( .A1(n16967), .A2(n9786), .ZN(n9789) );
  INV_X1 U12866 ( .A(n10513), .ZN(n10278) );
  NAND2_X1 U12867 ( .A1(n12890), .A2(n10514), .ZN(n10513) );
  NAND2_X1 U12868 ( .A1(n10008), .A2(n10005), .ZN(n9791) );
  OR2_X1 U12869 ( .A1(n17452), .A2(n11406), .ZN(n9792) );
  OR2_X1 U12870 ( .A1(n10882), .A2(n10881), .ZN(n9899) );
  INV_X1 U12871 ( .A(n15517), .ZN(n15269) );
  OR2_X1 U12872 ( .A1(n15447), .A2(n10366), .ZN(n9793) );
  AND3_X1 U12873 ( .A1(n9898), .A2(n9897), .A3(n10938), .ZN(n9794) );
  NAND2_X1 U12874 ( .A1(n11043), .A2(n11042), .ZN(n11180) );
  INV_X1 U12875 ( .A(n11180), .ZN(n10174) );
  NAND2_X1 U12876 ( .A1(n10231), .A2(n12756), .ZN(n12757) );
  AND2_X1 U12877 ( .A1(n11386), .A2(n11372), .ZN(n9795) );
  NAND2_X1 U12878 ( .A1(n10767), .A2(n10782), .ZN(n10761) );
  AND2_X1 U12879 ( .A1(n10135), .A2(n10134), .ZN(n9796) );
  AND2_X1 U12880 ( .A1(n10966), .A2(n10965), .ZN(n11085) );
  INV_X1 U12881 ( .A(n11085), .ZN(n9941) );
  NOR2_X1 U12882 ( .A1(n16436), .A2(n10423), .ZN(n11640) );
  AND2_X1 U12883 ( .A1(n10043), .A2(n10044), .ZN(n9797) );
  NAND2_X1 U12884 ( .A1(n10666), .A2(n10665), .ZN(n10712) );
  AND2_X1 U12885 ( .A1(n9953), .A2(n9952), .ZN(n9798) );
  NAND2_X1 U12886 ( .A1(n10474), .A2(n10478), .ZN(n9799) );
  NAND2_X1 U12887 ( .A1(n11530), .A2(n11529), .ZN(n16451) );
  INV_X1 U12888 ( .A(n12891), .ZN(n10243) );
  OR2_X1 U12889 ( .A1(n9688), .A2(n16146), .ZN(n12891) );
  NAND2_X1 U12890 ( .A1(n15894), .A2(n15893), .ZN(n9800) );
  AND2_X1 U12891 ( .A1(n15270), .A2(n10360), .ZN(n15489) );
  AND2_X1 U12892 ( .A1(n9938), .A2(n9940), .ZN(n9801) );
  INV_X1 U12893 ( .A(n10128), .ZN(n11438) );
  AND2_X1 U12894 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9802) );
  INV_X1 U12895 ( .A(n10066), .ZN(n10065) );
  NAND2_X1 U12896 ( .A1(n10540), .A2(n10067), .ZN(n10066) );
  NOR3_X1 U12897 ( .A1(n11087), .A2(n11482), .A3(n17384), .ZN(n9803) );
  AND2_X1 U12898 ( .A1(n14857), .A2(n9901), .ZN(n9804) );
  AND2_X1 U12899 ( .A1(n11467), .A2(n10562), .ZN(n9805) );
  NOR2_X1 U12900 ( .A1(n17236), .A2(n17237), .ZN(n9806) );
  NOR2_X1 U12901 ( .A1(n10970), .A2(n10271), .ZN(n9807) );
  AND2_X1 U12902 ( .A1(n12042), .A2(n13363), .ZN(n9808) );
  AND2_X1 U12903 ( .A1(n10494), .A2(n10495), .ZN(n9809) );
  AND2_X1 U12904 ( .A1(n10129), .A2(n10128), .ZN(n9810) );
  AND2_X1 U12905 ( .A1(n10190), .A2(n9963), .ZN(n9811) );
  AND2_X1 U12906 ( .A1(n10358), .A2(n10356), .ZN(n9812) );
  AND2_X1 U12907 ( .A1(n18861), .A2(n11858), .ZN(n9813) );
  AND2_X1 U12908 ( .A1(n9757), .A2(n10293), .ZN(n9814) );
  AND2_X1 U12909 ( .A1(n9938), .A2(n9785), .ZN(n9815) );
  INV_X1 U12910 ( .A(n12642), .ZN(n9945) );
  AND2_X1 U12911 ( .A1(n10461), .A2(n10466), .ZN(n9816) );
  AND2_X1 U12912 ( .A1(n10359), .A2(n9754), .ZN(n9817) );
  AND2_X1 U12913 ( .A1(n10243), .A2(n13160), .ZN(n9818) );
  OR2_X1 U12914 ( .A1(n16259), .A2(n13797), .ZN(n17892) );
  AND2_X1 U12915 ( .A1(n10449), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9819) );
  NAND2_X1 U12916 ( .A1(n10462), .A2(n9816), .ZN(n9820) );
  OR2_X1 U12917 ( .A1(n9945), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9821) );
  NAND2_X1 U12918 ( .A1(n18815), .A2(n18950), .ZN(n9822) );
  INV_X1 U12919 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14012) );
  NOR2_X1 U12920 ( .A1(n13375), .A2(n10249), .ZN(n9823) );
  INV_X1 U12921 ( .A(n10488), .ZN(n10487) );
  NAND2_X1 U12922 ( .A1(n14791), .A2(n14885), .ZN(n10488) );
  AND2_X2 U12923 ( .A1(n12379), .A2(n14353), .ZN(n10803) );
  AND2_X1 U12924 ( .A1(n13890), .A2(n10251), .ZN(n9824) );
  AND2_X1 U12925 ( .A1(n11442), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9825) );
  NAND2_X1 U12926 ( .A1(n9794), .A2(n10935), .ZN(n10968) );
  NOR2_X1 U12927 ( .A1(n15549), .A2(n15550), .ZN(n15537) );
  NOR2_X1 U12928 ( .A1(n13870), .A2(n13871), .ZN(n13869) );
  AND2_X1 U12929 ( .A1(n18908), .A2(n9814), .ZN(n17599) );
  NOR2_X1 U12930 ( .A1(n15761), .A2(n10525), .ZN(n9826) );
  OR2_X1 U12931 ( .A1(n11602), .A2(n10347), .ZN(n9827) );
  NOR2_X1 U12932 ( .A1(n14431), .A2(n14624), .ZN(n9828) );
  AND2_X1 U12933 ( .A1(n16759), .A2(n16758), .ZN(n9829) );
  OR2_X1 U12934 ( .A1(n11594), .A2(n10344), .ZN(n9830) );
  OR2_X1 U12935 ( .A1(n11602), .A2(n10349), .ZN(n9831) );
  AND2_X1 U12936 ( .A1(n17454), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9832) );
  INV_X1 U12937 ( .A(n12810), .ZN(n10501) );
  AND2_X1 U12938 ( .A1(n10401), .A2(n10399), .ZN(n9833) );
  NOR2_X1 U12939 ( .A1(n14431), .A2(n10398), .ZN(n14839) );
  AND2_X1 U12940 ( .A1(n14611), .A2(n14260), .ZN(n14252) );
  NOR2_X1 U12941 ( .A1(n14590), .A2(n11137), .ZN(n14641) );
  NAND2_X1 U12942 ( .A1(n11155), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11602) );
  NAND2_X1 U12943 ( .A1(n11266), .A2(n11265), .ZN(n13870) );
  NAND2_X1 U12944 ( .A1(n10341), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11596) );
  OR2_X1 U12945 ( .A1(n11602), .A2(n17020), .ZN(n9834) );
  OR2_X1 U12946 ( .A1(n10353), .A2(n11589), .ZN(n9835) );
  NOR2_X1 U12947 ( .A1(n12632), .A2(n21641), .ZN(n15043) );
  AOI21_X1 U12948 ( .B1(n9918), .B2(n9782), .A(n9917), .ZN(n17156) );
  AND2_X1 U12949 ( .A1(n16592), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9836) );
  INV_X1 U12950 ( .A(n14441), .ZN(n10013) );
  AND2_X1 U12952 ( .A1(n18795), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12118) );
  OR2_X1 U12953 ( .A1(n10893), .A2(n10892), .ZN(n11072) );
  NOR2_X1 U12954 ( .A1(n14584), .A2(n10520), .ZN(n14762) );
  NAND2_X1 U12955 ( .A1(n10383), .A2(n10387), .ZN(n13979) );
  AND2_X1 U12956 ( .A1(n10535), .A2(n10534), .ZN(n9838) );
  AND2_X1 U12957 ( .A1(n10531), .A2(n10530), .ZN(n9839) );
  OR2_X1 U12958 ( .A1(n14584), .A2(n17913), .ZN(n14772) );
  INV_X1 U12959 ( .A(n15761), .ZN(n10528) );
  OR2_X1 U12960 ( .A1(n19286), .A2(n19185), .ZN(n9840) );
  OR2_X1 U12961 ( .A1(n19175), .A2(n19399), .ZN(n9841) );
  NAND2_X1 U12962 ( .A1(n11367), .A2(n11366), .ZN(n11498) );
  OAI22_X1 U12963 ( .A1(n10126), .A2(n12242), .B1(n13772), .B2(n10559), .ZN(
        n16889) );
  AND2_X1 U12965 ( .A1(n13890), .A2(n9744), .ZN(n9842) );
  AND2_X1 U12966 ( .A1(n12823), .A2(n12822), .ZN(n9843) );
  OR2_X1 U12967 ( .A1(n19222), .A2(n19245), .ZN(n12163) );
  INV_X1 U12968 ( .A(n12163), .ZN(n10157) );
  AND2_X1 U12969 ( .A1(n10269), .A2(n10547), .ZN(n9844) );
  INV_X1 U12970 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10352) );
  NAND2_X1 U12971 ( .A1(n13073), .A2(n10531), .ZN(n10533) );
  NAND2_X1 U12972 ( .A1(n13431), .A2(n13430), .ZN(n9845) );
  INV_X1 U12973 ( .A(n17038), .ZN(n10440) );
  NAND2_X1 U12974 ( .A1(n11473), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n9846) );
  AND4_X1 U12975 ( .A1(n14706), .A2(n14595), .A3(n14564), .A4(n14422), .ZN(
        n9847) );
  INV_X1 U12976 ( .A(n10322), .ZN(n20147) );
  INV_X1 U12977 ( .A(n10388), .ZN(n10387) );
  NOR2_X1 U12978 ( .A1(n11247), .A2(n13916), .ZN(n10388) );
  INV_X1 U12979 ( .A(n15569), .ZN(n10038) );
  AND2_X1 U12980 ( .A1(n15104), .A2(n15103), .ZN(n15569) );
  AND2_X1 U12981 ( .A1(n11367), .A2(n9851), .ZN(n16470) );
  INV_X1 U12982 ( .A(n9918), .ZN(n10872) );
  NAND2_X1 U12983 ( .A1(n10842), .A2(n11073), .ZN(n9918) );
  NAND2_X1 U12984 ( .A1(n11154), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11594) );
  AND2_X1 U12985 ( .A1(n10469), .A2(n10468), .ZN(n9848) );
  NOR2_X1 U12986 ( .A1(n16592), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9849) );
  AND2_X1 U12987 ( .A1(n10465), .A2(n16686), .ZN(n9850) );
  AND2_X1 U12988 ( .A1(n15823), .A2(n15395), .ZN(n12921) );
  OR2_X1 U12989 ( .A1(n16103), .A2(n16158), .ZN(n10148) );
  NOR2_X1 U12990 ( .A1(n14584), .A2(n10522), .ZN(n14763) );
  INV_X1 U12991 ( .A(n10933), .ZN(n9931) );
  AND2_X1 U12992 ( .A1(n10395), .A2(n10394), .ZN(n9851) );
  AND2_X1 U12993 ( .A1(n9838), .A2(n15477), .ZN(n9852) );
  AND2_X1 U12994 ( .A1(n9708), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9853) );
  AND2_X1 U12995 ( .A1(n9839), .A2(n13083), .ZN(n9854) );
  INV_X1 U12996 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10343) );
  AND2_X1 U12997 ( .A1(n14449), .A2(n15395), .ZN(n13113) );
  AND2_X1 U12998 ( .A1(n12118), .A2(n9708), .ZN(n9855) );
  NAND2_X1 U12999 ( .A1(n11631), .A2(n9740), .ZN(n11637) );
  NAND2_X1 U13001 ( .A1(n14537), .A2(n14585), .ZN(n14584) );
  NAND2_X1 U13002 ( .A1(n11631), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9856) );
  NAND2_X1 U13003 ( .A1(n11618), .A2(n9736), .ZN(n11627) );
  AND2_X1 U13004 ( .A1(n9970), .A2(n19076), .ZN(n9857) );
  NOR2_X1 U13005 ( .A1(n13800), .A2(n14536), .ZN(n14537) );
  AND2_X1 U13006 ( .A1(n18587), .A2(n19448), .ZN(n18590) );
  INV_X1 U13007 ( .A(n16489), .ZN(n10325) );
  INV_X1 U13008 ( .A(n16924), .ZN(n10330) );
  AND3_X1 U13009 ( .A1(n10407), .A2(n16448), .A3(n10406), .ZN(n9858) );
  INV_X1 U13010 ( .A(n15380), .ZN(n10368) );
  NAND2_X1 U13011 ( .A1(n11618), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11620) );
  NAND2_X1 U13012 ( .A1(n11618), .A2(n9735), .ZN(n9859) );
  AND2_X1 U13013 ( .A1(n13359), .A2(n10241), .ZN(n9860) );
  AND2_X1 U13014 ( .A1(n13080), .A2(n13079), .ZN(n9861) );
  OR2_X1 U13015 ( .A1(n18950), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9862) );
  INV_X1 U13016 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10348) );
  NAND2_X1 U13017 ( .A1(n10528), .A2(n9729), .ZN(n15708) );
  INV_X1 U13018 ( .A(n15708), .ZN(n13054) );
  INV_X1 U13019 ( .A(n16681), .ZN(n10467) );
  NAND2_X1 U13020 ( .A1(n16724), .A2(n16728), .ZN(n9863) );
  NAND3_X1 U13021 ( .A1(n11305), .A2(n11304), .A3(n11303), .ZN(n9864) );
  INV_X1 U13022 ( .A(n10242), .ZN(n10241) );
  NAND2_X1 U13023 ( .A1(n9742), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n10242) );
  AND2_X1 U13024 ( .A1(n16686), .A2(n10467), .ZN(n9865) );
  AND2_X1 U13025 ( .A1(n9740), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9866) );
  INV_X1 U13026 ( .A(n17785), .ZN(n13314) );
  INV_X1 U13027 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n9877) );
  INV_X1 U13028 ( .A(n16117), .ZN(n17882) );
  AND4_X1 U13029 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n9868) );
  INV_X1 U13030 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19858) );
  AND2_X1 U13031 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n9869) );
  INV_X1 U13032 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n9878) );
  INV_X1 U13033 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n9968) );
  INV_X1 U13034 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18405) );
  INV_X1 U13035 ( .A(n16137), .ZN(n10497) );
  AND2_X1 U13036 ( .A1(n17301), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9870) );
  INV_X1 U13037 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10160) );
  INV_X1 U13038 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10458) );
  AND2_X1 U13039 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n9871) );
  INV_X1 U13040 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n10253) );
  INV_X1 U13041 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10295) );
  INV_X1 U13042 ( .A(n10220), .ZN(n10219) );
  NAND2_X1 U13043 ( .A1(n11488), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10220) );
  AND2_X1 U13044 ( .A1(n10078), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U13045 ( .A1(n13516), .A2(n21586), .ZN(n16117) );
  AND3_X1 U13046 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21638), .A3(n14448), 
        .ZN(n14479) );
  NAND2_X1 U13047 ( .A1(n21638), .A2(n14448), .ZN(n21189) );
  NAND2_X1 U13048 ( .A1(n21739), .A2(n21638), .ZN(n10231) );
  NOR2_X1 U13049 ( .A1(n12709), .A2(n21638), .ZN(n12865) );
  NOR2_X1 U13050 ( .A1(n12636), .A2(n21638), .ZN(n12743) );
  CLKBUF_X1 U13051 ( .A(n21356), .Z(n9873) );
  NOR2_X2 U13052 ( .A1(n20317), .A2(n9990), .ZN(n20772) );
  NAND2_X1 U13053 ( .A1(n20697), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20317) );
  NAND2_X2 U13054 ( .A1(n10029), .A2(n12652), .ZN(n12655) );
  NAND2_X2 U13055 ( .A1(n9874), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12652) );
  NAND4_X1 U13056 ( .A1(n12977), .A2(n13121), .A3(n10089), .A4(n12981), .ZN(
        n9874) );
  NAND2_X1 U13057 ( .A1(n10087), .A2(n12638), .ZN(n12977) );
  NAND2_X2 U13058 ( .A1(n9875), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10029) );
  NAND2_X2 U13059 ( .A1(n10230), .A2(n10095), .ZN(n15975) );
  NAND2_X2 U13060 ( .A1(n9880), .A2(n10009), .ZN(n10230) );
  NAND3_X1 U13061 ( .A1(n18088), .A2(n18089), .A3(n9882), .ZN(P3_U2641) );
  NAND2_X2 U13062 ( .A1(n15928), .A2(n15938), .ZN(n15927) );
  NAND2_X2 U13063 ( .A1(n9884), .A2(n15946), .ZN(n15928) );
  AND2_X4 U13064 ( .A1(n14331), .A2(n10573), .ZN(n12319) );
  NAND2_X2 U13065 ( .A1(n16930), .A2(n11454), .ZN(n10127) );
  NAND2_X1 U13066 ( .A1(n10837), .A2(n9887), .ZN(n9886) );
  NOR2_X1 U13067 ( .A1(n9890), .A2(n9889), .ZN(n9888) );
  NOR2_X1 U13068 ( .A1(n9893), .A2(n9892), .ZN(n9891) );
  NAND2_X2 U13069 ( .A1(n10991), .A2(n11456), .ZN(n10988) );
  NOR2_X4 U13070 ( .A1(n14705), .A2(n14643), .ZN(n16759) );
  NAND2_X2 U13071 ( .A1(n14250), .A2(n10470), .ZN(n14705) );
  NAND2_X2 U13072 ( .A1(n16889), .A2(n12246), .ZN(n14250) );
  AND2_X1 U13073 ( .A1(n12458), .A2(n12461), .ZN(n16687) );
  NAND2_X1 U13074 ( .A1(n9721), .A2(n12458), .ZN(n9902) );
  AND2_X2 U13075 ( .A1(n13904), .A2(n12233), .ZN(n13895) );
  INV_X1 U13076 ( .A(n13906), .ZN(n9905) );
  NAND2_X2 U13077 ( .A1(n13912), .A2(n11219), .ZN(n10726) );
  NAND2_X2 U13079 ( .A1(n9906), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10756) );
  NAND3_X1 U13080 ( .A1(n10728), .A2(n10727), .A3(n14333), .ZN(n9906) );
  NAND3_X2 U13081 ( .A1(n9957), .A2(n9795), .A3(n9692), .ZN(n14333) );
  NOR2_X2 U13082 ( .A1(n9907), .A2(n11184), .ZN(n10728) );
  AND2_X1 U13084 ( .A1(n11390), .A2(n10051), .ZN(n9907) );
  OAI21_X2 U13085 ( .B1(n11091), .B2(n10751), .A(n9947), .ZN(n11096) );
  XNOR2_X2 U13086 ( .A(n9909), .B(n11100), .ZN(n10760) );
  NAND2_X1 U13087 ( .A1(n10689), .A2(n14353), .ZN(n9919) );
  NAND2_X1 U13088 ( .A1(n10688), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9920) );
  NAND3_X1 U13089 ( .A1(n9685), .A2(n10710), .A3(n9922), .ZN(n10722) );
  NAND2_X1 U13090 ( .A1(n10707), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9923) );
  INV_X2 U13091 ( .A(n10840), .ZN(n10200) );
  NOR2_X1 U13092 ( .A1(n9927), .A2(n9926), .ZN(n9932) );
  NAND4_X1 U13093 ( .A1(n10919), .A2(n10915), .A3(n10913), .A4(n10918), .ZN(
        n9927) );
  NAND2_X1 U13094 ( .A1(n10118), .A2(n16694), .ZN(n9928) );
  NAND2_X1 U13095 ( .A1(n10117), .A2(n16694), .ZN(n9929) );
  NAND3_X1 U13096 ( .A1(n10836), .A2(n10835), .A3(n10834), .ZN(n9930) );
  INV_X1 U13097 ( .A(n9942), .ZN(n9935) );
  NAND2_X1 U13098 ( .A1(n9935), .A2(n11482), .ZN(n9934) );
  INV_X1 U13099 ( .A(n9937), .ZN(n11396) );
  NAND2_X1 U13100 ( .A1(n10690), .A2(n10721), .ZN(n9937) );
  NAND2_X1 U13101 ( .A1(n9937), .A2(n9990), .ZN(n10691) );
  NAND3_X1 U13102 ( .A1(n10029), .A2(n12642), .A3(n12652), .ZN(n9943) );
  NAND2_X1 U13103 ( .A1(n12655), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9946) );
  AND2_X2 U13104 ( .A1(n17032), .A2(n11089), .ZN(n17033) );
  INV_X1 U13105 ( .A(n16635), .ZN(n14360) );
  NAND3_X2 U13106 ( .A1(n9986), .A2(n10108), .A3(n10109), .ZN(n12214) );
  XNOR2_X2 U13107 ( .A(n13772), .B(n13777), .ZN(n20324) );
  NAND2_X1 U13108 ( .A1(n11374), .A2(n9957), .ZN(n14356) );
  INV_X1 U13109 ( .A(n10043), .ZN(n9961) );
  OAI21_X2 U13110 ( .B1(n11091), .B2(n11060), .A(n9715), .ZN(n10762) );
  AND2_X2 U13111 ( .A1(n9960), .A2(n9959), .ZN(n11099) );
  NAND3_X1 U13112 ( .A1(n10746), .A2(n10763), .A3(n10762), .ZN(n9959) );
  NAND2_X1 U13113 ( .A1(n10190), .A2(n9962), .ZN(n9967) );
  INV_X1 U13114 ( .A(n16917), .ZN(n9966) );
  NAND2_X1 U13115 ( .A1(n9972), .A2(n19076), .ZN(n9971) );
  NAND3_X1 U13116 ( .A1(n19093), .A2(n19076), .A3(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n9973) );
  NAND2_X1 U13117 ( .A1(n9975), .A2(n11827), .ZN(n9974) );
  INV_X1 U13118 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n9976) );
  NAND2_X1 U13119 ( .A1(n19092), .A2(n11827), .ZN(n19077) );
  NAND2_X1 U13120 ( .A1(n19093), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n19092) );
  OAI211_X1 U13121 ( .C1(n19052), .C2(n9985), .A(n9977), .B(n9983), .ZN(n19044) );
  NAND2_X1 U13122 ( .A1(n19052), .A2(n9982), .ZN(n9977) );
  NAND2_X1 U13123 ( .A1(n19052), .A2(n9979), .ZN(n9978) );
  NOR2_X1 U13124 ( .A1(n9982), .A2(n9980), .ZN(n9979) );
  NAND2_X1 U13125 ( .A1(n19052), .A2(n11841), .ZN(n11845) );
  NOR2_X1 U13126 ( .A1(n11844), .A2(n9984), .ZN(n9982) );
  NAND2_X1 U13127 ( .A1(n11844), .A2(n9984), .ZN(n9983) );
  INV_X1 U13128 ( .A(n11841), .ZN(n9984) );
  NAND3_X1 U13129 ( .A1(n10302), .A2(n10152), .A3(n9741), .ZN(n11866) );
  NOR2_X2 U13130 ( .A1(n11863), .A2(n11864), .ZN(n10302) );
  NOR2_X2 U13131 ( .A1(n10774), .A2(n17183), .ZN(n20393) );
  INV_X2 U13132 ( .A(n11220), .ZN(n9989) );
  OAI211_X2 U13133 ( .C1(n10756), .C2(n11398), .A(n10755), .B(n10754), .ZN(
        n11100) );
  OR2_X1 U13134 ( .A1(n14599), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9995) );
  AND2_X1 U13135 ( .A1(n12807), .A2(n12833), .ZN(n9996) );
  NAND2_X1 U13136 ( .A1(n14599), .A2(n9869), .ZN(n12807) );
  OAI21_X1 U13137 ( .B1(n16145), .B2(n21175), .A(n9997), .ZN(P1_U3002) );
  OAI211_X2 U13138 ( .C1(n12655), .C2(n10002), .A(n9999), .B(n9998), .ZN(
        n14442) );
  OAI21_X1 U13139 ( .B1(n12652), .B2(n10001), .A(n10000), .ZN(n9999) );
  NAND2_X1 U13140 ( .A1(n12652), .A2(n12641), .ZN(n10000) );
  NAND2_X1 U13141 ( .A1(n10004), .A2(n9688), .ZN(n10006) );
  NAND2_X1 U13142 ( .A1(n10008), .A2(n10007), .ZN(n10004) );
  NAND2_X1 U13143 ( .A1(n16022), .A2(n16033), .ZN(n10008) );
  NAND2_X1 U13144 ( .A1(n10277), .A2(n10227), .ZN(n17866) );
  OAI211_X2 U13145 ( .C1(n10014), .C2(n10013), .A(n10011), .B(n10010), .ZN(
        n21739) );
  NAND2_X1 U13146 ( .A1(n10014), .A2(n9720), .ZN(n10010) );
  INV_X1 U13147 ( .A(n12658), .ZN(n10012) );
  NAND2_X2 U13148 ( .A1(n12732), .A2(n12662), .ZN(n10014) );
  INV_X1 U13149 ( .A(n12757), .ZN(n10015) );
  AOI21_X2 U13150 ( .B1(n11837), .B2(n19356), .A(n10156), .ZN(n10154) );
  NOR2_X1 U13151 ( .A1(n17056), .A2(n10021), .ZN(n17340) );
  NAND2_X1 U13152 ( .A1(n10676), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10024) );
  NAND2_X1 U13153 ( .A1(n10671), .A2(n14353), .ZN(n10023) );
  NAND2_X2 U13154 ( .A1(n10028), .A2(n10157), .ZN(n11856) );
  AND2_X2 U13155 ( .A1(n12801), .A2(n12776), .ZN(n14659) );
  NAND3_X1 U13156 ( .A1(n12801), .A2(n12776), .A3(n15043), .ZN(n10030) );
  NAND2_X1 U13157 ( .A1(n14659), .A2(n12921), .ZN(n12782) );
  NAND2_X1 U13158 ( .A1(n14659), .A2(n12757), .ZN(n21581) );
  NAND2_X1 U13159 ( .A1(n14659), .A2(n10015), .ZN(n21365) );
  INV_X1 U13160 ( .A(n14659), .ZN(n10031) );
  XNOR2_X1 U13161 ( .A(n14659), .B(n21580), .ZN(n14512) );
  AND2_X2 U13162 ( .A1(n15758), .A2(n14959), .ZN(n15656) );
  NOR2_X2 U13163 ( .A1(n14941), .A2(n15760), .ZN(n15758) );
  NAND2_X1 U13164 ( .A1(n17495), .A2(n11220), .ZN(n20968) );
  NAND3_X1 U13165 ( .A1(n9685), .A2(n9990), .A3(n17495), .ZN(n10041) );
  XNOR2_X2 U13166 ( .A(n10042), .B(n10043), .ZN(n10767) );
  OAI211_X2 U13167 ( .C1(n10756), .C2(n13332), .A(n10731), .B(n10732), .ZN(
        n10044) );
  XNOR2_X1 U13168 ( .A(n17099), .B(n17348), .ZN(n17376) );
  NAND2_X1 U13169 ( .A1(n11422), .A2(n10049), .ZN(n10431) );
  NAND2_X2 U13170 ( .A1(n17132), .A2(n17133), .ZN(n11422) );
  NAND3_X1 U13171 ( .A1(n10842), .A2(n11073), .A3(n9819), .ZN(n10053) );
  NAND2_X1 U13172 ( .A1(n17032), .A2(n10055), .ZN(n17021) );
  NAND3_X1 U13173 ( .A1(n10784), .A2(n10056), .A3(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10822) );
  OR2_X1 U13174 ( .A1(n14852), .A2(n10061), .ZN(n10057) );
  NAND2_X1 U13175 ( .A1(n10057), .A2(n10059), .ZN(n16975) );
  NAND2_X1 U13176 ( .A1(n14852), .A2(n11435), .ZN(n10062) );
  NAND2_X1 U13177 ( .A1(n10068), .A2(n10718), .ZN(n10719) );
  OAI211_X1 U13178 ( .C1(n10127), .C2(n10488), .A(n10485), .B(n9730), .ZN(
        n10221) );
  OAI22_X1 U13179 ( .A1(n10072), .A2(n17565), .B1(n10297), .B2(n10298), .ZN(
        n10075) );
  INV_X1 U13180 ( .A(n10299), .ZN(n10074) );
  AOI21_X2 U13181 ( .B1(n11871), .B2(n11870), .A(n10075), .ZN(n12156) );
  AND3_X2 U13182 ( .A1(n9822), .A2(n10077), .A3(n10076), .ZN(n18798) );
  NAND2_X1 U13183 ( .A1(n18614), .A2(n9872), .ZN(n18602) );
  NAND2_X1 U13185 ( .A1(n13496), .A2(n10085), .ZN(n13737) );
  AND3_X2 U13186 ( .A1(n10091), .A2(n12648), .A3(n10508), .ZN(n12638) );
  NAND4_X1 U13187 ( .A1(n14449), .A2(n10090), .A3(n9718), .A4(n12917), .ZN(
        n10089) );
  INV_X1 U13188 ( .A(n13750), .ZN(n12962) );
  AND2_X2 U13189 ( .A1(n13495), .A2(n13130), .ZN(n10090) );
  NOR2_X2 U13190 ( .A1(n12880), .A2(n16034), .ZN(n16022) );
  NOR2_X1 U13191 ( .A1(n12890), .A2(n16260), .ZN(n16034) );
  NAND2_X1 U13192 ( .A1(n16055), .A2(n10092), .ZN(n12880) );
  NAND2_X1 U13193 ( .A1(n12893), .A2(n10096), .ZN(n12895) );
  NAND2_X1 U13194 ( .A1(n10098), .A2(n10097), .ZN(n10096) );
  INV_X1 U13195 ( .A(n10099), .ZN(n10097) );
  NAND2_X1 U13196 ( .A1(n10100), .A2(n10496), .ZN(n10098) );
  OAI21_X1 U13197 ( .B1(n15938), .B2(n10101), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10099) );
  NAND2_X1 U13198 ( .A1(n15927), .A2(n10496), .ZN(n15903) );
  INV_X1 U13199 ( .A(n10496), .ZN(n10101) );
  NAND2_X1 U13200 ( .A1(n16957), .A2(n16958), .ZN(n16930) );
  AOI22_X1 U13201 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10912), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10776) );
  NAND3_X2 U13202 ( .A1(n10452), .A2(n10451), .A3(n10450), .ZN(n10753) );
  AND2_X4 U13203 ( .A1(n12511), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14290) );
  NAND2_X1 U13204 ( .A1(n13441), .A2(n13458), .ZN(n12090) );
  NAND2_X2 U13205 ( .A1(n14571), .A2(n12110), .ZN(n19280) );
  OAI21_X1 U13206 ( .B1(n10760), .B2(n10759), .A(n10111), .ZN(n10108) );
  NAND3_X1 U13207 ( .A1(n10758), .A2(n10761), .A3(n10110), .ZN(n10109) );
  NAND2_X1 U13208 ( .A1(n11097), .A2(n10760), .ZN(n10111) );
  NAND2_X1 U13209 ( .A1(n16966), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10112) );
  NAND3_X1 U13210 ( .A1(n10787), .A2(n10786), .A3(n10785), .ZN(n10118) );
  XNOR2_X2 U13211 ( .A(n10119), .B(n17384), .ZN(n17109) );
  NOR2_X2 U13212 ( .A1(n11087), .A2(n11482), .ZN(n10119) );
  NAND2_X1 U13213 ( .A1(n9820), .A2(n10120), .ZN(n12495) );
  NOR2_X1 U13214 ( .A1(n16675), .A2(n16883), .ZN(n10120) );
  NAND3_X1 U13215 ( .A1(n14859), .A2(n10130), .A3(n9810), .ZN(n10413) );
  NAND2_X2 U13216 ( .A1(n11015), .A2(n11014), .ZN(n11027) );
  NAND2_X1 U13217 ( .A1(n13883), .A2(n10139), .ZN(n14321) );
  AND2_X1 U13218 ( .A1(n13884), .A2(n14320), .ZN(n10139) );
  NAND2_X1 U13219 ( .A1(n15928), .A2(n9689), .ZN(n10150) );
  OAI211_X1 U13220 ( .C1(n15928), .C2(n10143), .A(n10144), .B(n10142), .ZN(
        n10147) );
  NAND2_X1 U13221 ( .A1(n15928), .A2(n10143), .ZN(n10142) );
  NOR2_X1 U13222 ( .A1(n16103), .A2(n16158), .ZN(n10143) );
  NAND3_X1 U13223 ( .A1(n10149), .A2(n10147), .A3(n10145), .ZN(n16163) );
  OAI21_X2 U13224 ( .B1(n15947), .B2(n12887), .A(n16103), .ZN(n15938) );
  OR2_X1 U13225 ( .A1(n10301), .A2(n10153), .ZN(n19129) );
  NOR2_X1 U13226 ( .A1(n18798), .A2(n18799), .ZN(n10153) );
  OAI21_X2 U13227 ( .B1(n19065), .B2(n10155), .A(n10154), .ZN(n19052) );
  AND2_X1 U13228 ( .A1(n11678), .A2(n11681), .ZN(n10159) );
  NAND2_X1 U13229 ( .A1(n11818), .A2(n12079), .ZN(n11819) );
  NAND2_X2 U13230 ( .A1(n9802), .A2(n10249), .ZN(n18541) );
  NAND3_X1 U13231 ( .A1(n10161), .A2(n12664), .A3(n21638), .ZN(n10355) );
  NAND2_X1 U13232 ( .A1(n10161), .A2(n12664), .ZN(n21391) );
  OR2_X1 U13233 ( .A1(n10161), .A2(n10013), .ZN(n13762) );
  INV_X1 U13234 ( .A(n12802), .ZN(n10167) );
  NAND2_X1 U13235 ( .A1(n12811), .A2(n12921), .ZN(n10193) );
  NAND2_X1 U13236 ( .A1(n17033), .A2(n10170), .ZN(n10168) );
  NAND2_X1 U13237 ( .A1(n10168), .A2(n10169), .ZN(n14850) );
  NOR2_X2 U13238 ( .A1(n17253), .A2(n17242), .ZN(n17231) );
  NOR2_X1 U13239 ( .A1(n17216), .A2(n11563), .ZN(n14818) );
  NAND4_X1 U13240 ( .A1(n10176), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n11483), .ZN(n10175) );
  NOR2_X1 U13241 ( .A1(n10179), .A2(n10177), .ZN(n11565) );
  NAND2_X1 U13242 ( .A1(n10934), .A2(n11084), .ZN(n10443) );
  INV_X1 U13243 ( .A(n17146), .ZN(n11081) );
  OAI21_X1 U13244 ( .B1(n14822), .B2(n17458), .A(n10182), .ZN(P2_U3019) );
  INV_X1 U13245 ( .A(n10183), .ZN(n10182) );
  OAI21_X1 U13246 ( .B1(n14812), .B2(n17415), .A(n10184), .ZN(n10183) );
  AND2_X2 U13247 ( .A1(n17032), .A2(n10186), .ZN(n16922) );
  NAND2_X1 U13248 ( .A1(n16922), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14892) );
  OAI211_X1 U13249 ( .C1(n12802), .C2(n10192), .A(n10191), .B(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10194) );
  NAND3_X1 U13250 ( .A1(n10197), .A2(n10195), .A3(n17873), .ZN(n10277) );
  NAND3_X1 U13251 ( .A1(n12808), .A2(n12809), .A3(n12807), .ZN(n17879) );
  NAND2_X1 U13252 ( .A1(n10196), .A2(n12833), .ZN(n10195) );
  INV_X1 U13253 ( .A(n14505), .ZN(n10198) );
  NAND2_X1 U13254 ( .A1(n10447), .A2(n11083), .ZN(n17104) );
  AOI21_X1 U13255 ( .B1(n10202), .B2(n17109), .A(n9803), .ZN(n10201) );
  AOI21_X2 U13256 ( .B1(n10544), .B2(n10412), .A(n10212), .ZN(n10222) );
  NAND2_X1 U13257 ( .A1(n16922), .A2(n10217), .ZN(n10216) );
  OAI211_X1 U13258 ( .C1(n16922), .C2(n11483), .A(n10218), .B(n10216), .ZN(
        n15426) );
  NAND2_X1 U13259 ( .A1(n14886), .A2(n10221), .ZN(n14891) );
  NAND2_X1 U13260 ( .A1(n10442), .A2(n14784), .ZN(n10940) );
  OAI21_X2 U13261 ( .B1(n10230), .B2(n10278), .A(n10229), .ZN(n15918) );
  NAND2_X1 U13262 ( .A1(n21739), .A2(n10235), .ZN(n10234) );
  NAND2_X1 U13263 ( .A1(n15904), .A2(n12892), .ZN(n12893) );
  NAND3_X1 U13264 ( .A1(n15938), .A2(n15928), .A3(n9818), .ZN(n15904) );
  AND2_X1 U13265 ( .A1(n18505), .A2(n10244), .ZN(n18496) );
  NAND2_X1 U13266 ( .A1(n10261), .A2(n10258), .ZN(n12967) );
  NAND2_X1 U13267 ( .A1(n10261), .A2(n10262), .ZN(n13753) );
  NOR2_X2 U13268 ( .A1(n16178), .A2(n10268), .ZN(n16159) );
  NOR2_X1 U13269 ( .A1(n11027), .A2(n9733), .ZN(n11430) );
  OR2_X2 U13270 ( .A1(n11027), .A2(n9738), .ZN(n11445) );
  NAND2_X1 U13271 ( .A1(n11445), .A2(n11456), .ZN(n11444) );
  NOR2_X2 U13272 ( .A1(n10970), .A2(n10270), .ZN(n10979) );
  NAND2_X1 U13273 ( .A1(n10273), .A2(n10272), .ZN(n15434) );
  NAND2_X1 U13274 ( .A1(n11481), .A2(n10878), .ZN(n10272) );
  OAI21_X1 U13275 ( .B1(n11480), .B2(P2_EBX_REG_30__SCAN_IN), .A(n11473), .ZN(
        n10273) );
  NAND2_X1 U13276 ( .A1(n11472), .A2(n11471), .ZN(n11480) );
  XNOR2_X2 U13277 ( .A(n10274), .B(n12682), .ZN(n13502) );
  AND2_X2 U13278 ( .A1(n12520), .A2(n10275), .ZN(n12717) );
  AND2_X2 U13279 ( .A1(n12517), .A2(n10275), .ZN(n15283) );
  XNOR2_X2 U13280 ( .A(n10276), .B(n12783), .ZN(n14665) );
  INV_X1 U13281 ( .A(n10285), .ZN(n18125) );
  OR2_X1 U13282 ( .A1(n18132), .A2(n18339), .ZN(n10285) );
  INV_X1 U13283 ( .A(n19069), .ZN(n10286) );
  NOR2_X1 U13284 ( .A1(n18091), .A2(n18339), .ZN(n18083) );
  NAND2_X1 U13285 ( .A1(n12118), .A2(n9853), .ZN(n12127) );
  INV_X1 U13286 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10296) );
  NAND2_X2 U13287 ( .A1(n18815), .A2(n10303), .ZN(n18816) );
  AND2_X2 U13288 ( .A1(n18861), .A2(n10304), .ZN(n10303) );
  INV_X1 U13289 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10305) );
  NAND2_X1 U13290 ( .A1(n10308), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10306) );
  NAND2_X1 U13291 ( .A1(n10309), .A2(n14353), .ZN(n10307) );
  NAND4_X1 U13292 ( .A1(n10599), .A2(n10598), .A3(n10600), .A4(n10601), .ZN(
        n10308) );
  NAND4_X1 U13293 ( .A1(n10605), .A2(n10604), .A3(n10602), .A4(n10603), .ZN(
        n10309) );
  AOI21_X1 U13294 ( .B1(n10317), .B2(n10316), .A(n13223), .ZN(n11201) );
  NAND2_X1 U13295 ( .A1(n16488), .A2(n10322), .ZN(n10321) );
  NAND2_X1 U13296 ( .A1(n10321), .A2(n10323), .ZN(n16476) );
  NAND2_X1 U13297 ( .A1(n11631), .A2(n9866), .ZN(n11572) );
  INV_X1 U13298 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10327) );
  NAND3_X1 U13299 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11580) );
  INV_X1 U13300 ( .A(n11594), .ZN(n10341) );
  NAND2_X1 U13301 ( .A1(n10341), .A2(n10342), .ZN(n11600) );
  NAND2_X1 U13302 ( .A1(n11153), .A2(n10350), .ZN(n11591) );
  INV_X1 U13303 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10354) );
  NAND2_X2 U13304 ( .A1(n13500), .A2(n15823), .ZN(n12635) );
  NAND3_X1 U13305 ( .A1(n13495), .A2(n13130), .A3(n13500), .ZN(n13302) );
  NAND2_X1 U13306 ( .A1(n10355), .A2(n12676), .ZN(n12680) );
  OAI21_X1 U13307 ( .B1(n15447), .B2(n15448), .A(n10368), .ZN(n10367) );
  NAND2_X1 U13308 ( .A1(n9793), .A2(n10361), .ZN(P1_U2873) );
  NOR2_X1 U13309 ( .A1(n15447), .A2(n15448), .ZN(n15446) );
  NAND2_X1 U13310 ( .A1(n15656), .A2(n10374), .ZN(n15515) );
  NAND2_X1 U13311 ( .A1(n14777), .A2(n10379), .ZN(n10378) );
  NAND2_X1 U13312 ( .A1(n10378), .A2(n10381), .ZN(n13976) );
  NAND2_X1 U13313 ( .A1(n13903), .A2(n10404), .ZN(n16597) );
  AND2_X1 U13314 ( .A1(n16447), .A2(n9858), .ZN(n14914) );
  NAND2_X1 U13315 ( .A1(n16447), .A2(n10405), .ZN(n11648) );
  NAND2_X1 U13316 ( .A1(n16447), .A2(n16448), .ZN(n16425) );
  INV_X2 U13317 ( .A(n14590), .ZN(n10415) );
  NAND2_X1 U13318 ( .A1(n14611), .A2(n10417), .ZN(n14492) );
  NAND2_X1 U13319 ( .A1(n14836), .A2(n10418), .ZN(n14864) );
  NOR2_X1 U13320 ( .A1(n16436), .A2(n16420), .ZN(n10428) );
  OR3_X1 U13321 ( .A1(n16436), .A2(n10422), .A3(n16420), .ZN(n12505) );
  INV_X2 U13322 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10575) );
  NAND2_X1 U13323 ( .A1(n10429), .A2(n10433), .ZN(n14852) );
  NAND3_X1 U13324 ( .A1(n11422), .A2(n10430), .A3(n10997), .ZN(n10429) );
  NAND3_X1 U13325 ( .A1(n10934), .A2(n11084), .A3(n11482), .ZN(n10442) );
  NAND2_X1 U13326 ( .A1(n14824), .A2(n11018), .ZN(n14823) );
  AND2_X2 U13327 ( .A1(n10056), .A2(n10783), .ZN(n20361) );
  NAND2_X1 U13328 ( .A1(n11076), .A2(n17158), .ZN(n10446) );
  NAND3_X1 U13329 ( .A1(n10446), .A2(n10445), .A3(n17144), .ZN(n17142) );
  OAI21_X1 U13330 ( .B1(n11080), .B2(n9790), .A(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10447) );
  NAND2_X1 U13331 ( .A1(n10448), .A2(n11082), .ZN(n17131) );
  NAND2_X1 U13332 ( .A1(n11083), .A2(n11080), .ZN(n10448) );
  INV_X1 U13333 ( .A(n11082), .ZN(n9790) );
  NAND3_X1 U13334 ( .A1(n10696), .A2(n10695), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10452) );
  NAND4_X1 U13335 ( .A1(n10654), .A2(n10653), .A3(n10651), .A4(n10652), .ZN(
        n10459) );
  NAND4_X1 U13336 ( .A1(n10650), .A2(n10647), .A3(n10648), .A4(n10649), .ZN(
        n10460) );
  NAND2_X1 U13337 ( .A1(n16687), .A2(n9865), .ZN(n10462) );
  NAND2_X1 U13338 ( .A1(n16687), .A2(n16686), .ZN(n16685) );
  INV_X1 U13339 ( .A(n12461), .ZN(n10464) );
  INV_X1 U13340 ( .A(n10544), .ZN(n10472) );
  NAND2_X1 U13341 ( .A1(n10473), .A2(n10472), .ZN(n10471) );
  XNOR2_X1 U13342 ( .A(n10471), .B(n9789), .ZN(n17261) );
  INV_X1 U13343 ( .A(n16601), .ZN(n10484) );
  NAND3_X1 U13344 ( .A1(n10486), .A2(n10489), .A3(n10485), .ZN(n14888) );
  NAND2_X1 U13345 ( .A1(n10491), .A2(n14791), .ZN(n14884) );
  NAND2_X1 U13346 ( .A1(n10490), .A2(n14792), .ZN(n10489) );
  INV_X1 U13347 ( .A(n14791), .ZN(n10490) );
  INV_X1 U13348 ( .A(n10562), .ZN(n10493) );
  NAND2_X1 U13349 ( .A1(n12890), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10498) );
  NAND3_X1 U13350 ( .A1(n10502), .A2(n12757), .A3(n10501), .ZN(n10499) );
  NAND2_X1 U13351 ( .A1(n13502), .A2(n10506), .ZN(n10504) );
  NAND2_X1 U13352 ( .A1(n13502), .A2(n21638), .ZN(n10505) );
  INV_X1 U13353 ( .A(n10509), .ZN(n10508) );
  NAND2_X1 U13354 ( .A1(n14464), .A2(n12632), .ZN(n12631) );
  NAND2_X1 U13355 ( .A1(n12636), .A2(n14464), .ZN(n12634) );
  NAND3_X1 U13356 ( .A1(n12966), .A2(n15823), .A3(n12632), .ZN(n10510) );
  NAND3_X1 U13357 ( .A1(n13584), .A2(n13000), .A3(n12992), .ZN(n13800) );
  NAND3_X1 U13358 ( .A1(n12824), .A2(n12846), .A3(n12921), .ZN(n12831) );
  AOI21_X1 U13359 ( .B1(n10511), .B2(n15043), .A(n14653), .ZN(n14655) );
  INV_X1 U13360 ( .A(n12884), .ZN(n10517) );
  NAND2_X1 U13361 ( .A1(n13054), .A2(n9728), .ZN(n15647) );
  NAND2_X1 U13362 ( .A1(n13073), .A2(n9854), .ZN(n15570) );
  INV_X1 U13363 ( .A(n10533), .ZN(n15609) );
  NAND2_X1 U13364 ( .A1(n15518), .A2(n9852), .ZN(n15459) );
  NAND2_X1 U13365 ( .A1(n11130), .A2(n11129), .ZN(n14590) );
  INV_X1 U13366 ( .A(n14425), .ZN(n11130) );
  AOI21_X1 U13367 ( .B1(n14907), .B2(n17456), .A(n14906), .ZN(n14908) );
  XNOR2_X1 U13368 ( .A(n16978), .B(n16977), .ZN(n17275) );
  INV_X1 U13369 ( .A(n15515), .ZN(n15270) );
  AND3_X1 U13370 ( .A1(n13134), .A2(n13130), .A3(n12972), .ZN(n13612) );
  INV_X1 U13371 ( .A(n13976), .ZN(n11266) );
  NOR2_X2 U13372 ( .A1(n14492), .A2(n14493), .ZN(n14424) );
  INV_X1 U13373 ( .A(n14655), .ZN(n14654) );
  INV_X1 U13374 ( .A(n14864), .ZN(n11530) );
  NAND2_X1 U13375 ( .A1(n10726), .A2(n11389), .ZN(n11186) );
  CLKBUF_X1 U13376 ( .A(n14941), .Z(n15759) );
  NOR2_X1 U13377 ( .A1(n11389), .A2(n11208), .ZN(n10690) );
  NOR2_X2 U13378 ( .A1(n16753), .A2(n14845), .ZN(n14836) );
  AND2_X1 U13379 ( .A1(n20298), .A2(n11220), .ZN(n10709) );
  OAI21_X1 U13381 ( .B1(n15429), .B2(n17429), .A(n11565), .ZN(n11566) );
  CLKBUF_X1 U13382 ( .A(n16957), .Z(n16959) );
  INV_X1 U13383 ( .A(n14665), .ZN(n21185) );
  NAND2_X1 U13384 ( .A1(n21186), .A2(n14665), .ZN(n21451) );
  NAND2_X1 U13385 ( .A1(n14914), .A2(n11647), .ZN(n12189) );
  NAND2_X1 U13386 ( .A1(n16705), .A2(n16706), .ZN(n16707) );
  NOR2_X1 U13387 ( .A1(n11419), .A2(n11418), .ZN(n11420) );
  AOI22_X1 U13388 ( .A1(n12319), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12317), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U13389 ( .A1(n12319), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12317), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10662) );
  AOI22_X1 U13390 ( .A1(n12319), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12317), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10655) );
  AOI22_X1 U13391 ( .A1(n12319), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12317), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U13392 ( .A1(n12317), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10588) );
  NAND2_X4 U13393 ( .A1(n10566), .A2(n12535), .ZN(n15823) );
  NAND2_X2 U13394 ( .A1(n12984), .A2(n14449), .ZN(n12994) );
  NAND2_X1 U13395 ( .A1(n14666), .A2(n12732), .ZN(n14505) );
  AND2_X1 U13396 ( .A1(n10128), .A2(n11423), .ZN(n10537) );
  INV_X1 U13397 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n11573) );
  AND3_X1 U13398 ( .A1(n11849), .A2(n11848), .A3(n11847), .ZN(n10538) );
  NAND2_X1 U13399 ( .A1(n16470), .A2(n11505), .ZN(n16456) );
  AND4_X1 U13400 ( .A1(n19245), .A2(n11852), .A3(n11851), .A4(n11850), .ZN(
        n10539) );
  AND2_X1 U13401 ( .A1(n11018), .A2(n14826), .ZN(n10540) );
  AND3_X1 U13402 ( .A1(n12007), .A2(n12006), .A3(n12005), .ZN(n10541) );
  AND4_X1 U13403 ( .A1(n13174), .A2(n10546), .A3(n13173), .A4(n9788), .ZN(
        n10542) );
  AND2_X1 U13404 ( .A1(n13033), .A2(n13032), .ZN(n10543) );
  AND2_X1 U13405 ( .A1(n16032), .A2(n16044), .ZN(n10545) );
  OR3_X1 U13406 ( .A1(n16130), .A2(n13161), .A3(n12894), .ZN(n10546) );
  AND2_X1 U13407 ( .A1(n16437), .A2(n16699), .ZN(n10547) );
  INV_X1 U13408 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17090) );
  AND2_X2 U13409 ( .A1(n14287), .A2(n12517), .ZN(n12610) );
  AND4_X1 U13410 ( .A1(n10642), .A2(n10641), .A3(n10640), .A4(n10639), .ZN(
        n10548) );
  AND2_X1 U13411 ( .A1(n10588), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10549) );
  NAND3_X1 U13412 ( .A1(n11318), .A2(n11317), .A3(n11316), .ZN(n10550) );
  AND2_X1 U13413 ( .A1(n12589), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10551) );
  AND2_X2 U13414 ( .A1(n10782), .A2(n10768), .ZN(n17455) );
  NAND2_X1 U13415 ( .A1(n11444), .A2(n11443), .ZN(n11447) );
  INV_X1 U13416 ( .A(n15758), .ZN(n15894) );
  INV_X1 U13417 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n13237) );
  INV_X1 U13418 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17029) );
  INV_X1 U13419 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11483) );
  INV_X1 U13420 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17071) );
  INV_X1 U13421 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13764) );
  INV_X1 U13422 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11849) );
  NAND2_X1 U13423 ( .A1(n11473), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10552) );
  NOR2_X2 U13424 ( .A1(n10322), .A2(n20177), .ZN(n20107) );
  NOR2_X1 U13425 ( .A1(n20628), .A2(n20562), .ZN(n10555) );
  NOR2_X1 U13426 ( .A1(n21522), .A2(n21574), .ZN(n10556) );
  NOR2_X1 U13427 ( .A1(n21522), .A2(n21361), .ZN(n10557) );
  INV_X1 U13428 ( .A(n11156), .ZN(n11571) );
  NAND2_X1 U13429 ( .A1(n11157), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11156) );
  INV_X1 U13430 ( .A(n10900), .ZN(n10945) );
  AND4_X1 U13431 ( .A1(n10638), .A2(n10637), .A3(n10636), .A4(n10635), .ZN(
        n10558) );
  NAND2_X1 U13432 ( .A1(n19116), .A2(n17601), .ZN(n18868) );
  AND2_X1 U13433 ( .A1(n12243), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10559) );
  AND2_X1 U13434 ( .A1(n11219), .A2(n12243), .ZN(n10560) );
  INV_X1 U13435 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n11055) );
  NAND2_X1 U13436 ( .A1(n12457), .A2(n12456), .ZN(n12461) );
  NAND3_X1 U13437 ( .A1(n11356), .A2(n11355), .A3(n11354), .ZN(n10561) );
  INV_X1 U13438 ( .A(n14885), .ZN(n14792) );
  NAND2_X1 U13439 ( .A1(n16945), .A2(n11455), .ZN(n10562) );
  NAND2_X1 U13440 ( .A1(n13918), .A2(n13919), .ZN(n10563) );
  NOR2_X1 U13441 ( .A1(n20650), .A2(n20629), .ZN(n10564) );
  INV_X1 U13442 ( .A(n17480), .ZN(n20476) );
  INV_X1 U13443 ( .A(n14464), .ZN(n15824) );
  AND2_X2 U13444 ( .A1(n14304), .A2(n12519), .ZN(n12696) );
  AND4_X1 U13445 ( .A1(n12585), .A2(n12584), .A3(n12583), .A4(n12582), .ZN(
        n10565) );
  NAND2_X1 U13446 ( .A1(n20361), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10816) );
  NAND2_X1 U13447 ( .A1(n10817), .A2(n10816), .ZN(n10818) );
  INV_X1 U13448 ( .A(n12911), .ZN(n12900) );
  NAND2_X1 U13449 ( .A1(n21392), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12901) );
  INV_X1 U13450 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12902) );
  INV_X1 U13451 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12510) );
  NAND2_X1 U13452 ( .A1(n12900), .A2(n12899), .ZN(n12912) );
  INV_X1 U13453 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12511) );
  AOI22_X1 U13454 ( .A1(n12959), .A2(n12825), .B1(n12948), .B2(
        P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12810) );
  OR2_X1 U13455 ( .A1(n12768), .A2(n12767), .ZN(n12825) );
  INV_X1 U13456 ( .A(n12769), .ZN(n12790) );
  NAND2_X1 U13457 ( .A1(n11036), .A2(n10878), .ZN(n10880) );
  INV_X1 U13458 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11847) );
  INV_X1 U13459 ( .A(n15153), .ZN(n15087) );
  OR2_X1 U13460 ( .A1(n12843), .A2(n12842), .ZN(n12855) );
  NOR2_X1 U13461 ( .A1(n12890), .A2(n16202), .ZN(n12884) );
  INV_X1 U13462 ( .A(n9750), .ZN(n13035) );
  INV_X1 U13463 ( .A(n13801), .ZN(n13000) );
  AND2_X1 U13464 ( .A1(n13744), .A2(n15776), .ZN(n13142) );
  INV_X1 U13465 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13740) );
  NAND2_X1 U13466 ( .A1(n12657), .A2(n12656), .ZN(n12659) );
  AOI22_X1 U13467 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n12319), .B1(
        n12317), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10674) );
  INV_X1 U13468 ( .A(n10717), .ZN(n10718) );
  INV_X1 U13469 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n12049) );
  NOR2_X1 U13470 ( .A1(n18950), .A2(n17652), .ZN(n11864) );
  OR2_X1 U13471 ( .A1(n11842), .A2(n17632), .ZN(n11843) );
  AND2_X1 U13472 ( .A1(n12950), .A2(n12951), .ZN(n12949) );
  INV_X1 U13473 ( .A(n15461), .ZN(n13114) );
  INV_X1 U13474 ( .A(n15271), .ZN(n15272) );
  INV_X1 U13475 ( .A(n15893), .ZN(n14959) );
  AND2_X2 U13476 ( .A1(n14977), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14997) );
  INV_X1 U13477 ( .A(n11450), .ZN(n11448) );
  INV_X1 U13478 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11598) );
  AND2_X1 U13479 ( .A1(n11473), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10971) );
  OR2_X1 U13480 ( .A1(n11041), .A2(n11040), .ZN(n11043) );
  XNOR2_X1 U13481 ( .A(n16707), .B(n12431), .ZN(n16691) );
  AND4_X1 U13482 ( .A1(n10846), .A2(n10845), .A3(n10844), .A4(n10843), .ZN(
        n10871) );
  INV_X1 U13483 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15588) );
  NAND2_X1 U13484 ( .A1(n13917), .A2(n11234), .ZN(n13920) );
  AND2_X1 U13485 ( .A1(n10591), .A2(n14353), .ZN(n10595) );
  AND2_X1 U13486 ( .A1(n12049), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12065) );
  INV_X1 U13487 ( .A(n17572), .ZN(n12122) );
  OR2_X1 U13488 ( .A1(n18545), .A2(n12013), .ZN(n12014) );
  AND2_X1 U13489 ( .A1(n21074), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21082) );
  OR3_X1 U13490 ( .A1(n13753), .A2(n20982), .A3(n14293), .ZN(n13413) );
  NAND2_X1 U13491 ( .A1(n12696), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12601) );
  NAND2_X1 U13492 ( .A1(n16350), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n15375) );
  NAND2_X1 U13493 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n14976), .ZN(
        n15079) );
  INV_X1 U13494 ( .A(n15630), .ZN(n13072) );
  OR3_X1 U13495 ( .A1(n13759), .A2(n13758), .A3(n13757), .ZN(n17825) );
  NAND2_X1 U13496 ( .A1(n12742), .A2(n12741), .ZN(n14441) );
  INV_X1 U13497 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21392) );
  INV_X1 U13498 ( .A(n11157), .ZN(n11610) );
  INV_X1 U13499 ( .A(n16720), .ZN(n11529) );
  INV_X1 U13500 ( .A(n14563), .ZN(n11129) );
  OR2_X1 U13501 ( .A1(n11261), .A2(n11260), .ZN(n12249) );
  OAI21_X1 U13502 ( .B1(n14360), .B2(n12239), .A(n12224), .ZN(n13906) );
  XNOR2_X1 U13503 ( .A(n11096), .B(n10765), .ZN(n10766) );
  AND2_X1 U13504 ( .A1(n10998), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17038) );
  NAND2_X1 U13505 ( .A1(n14424), .A2(n14426), .ZN(n14425) );
  NAND2_X1 U13506 ( .A1(n17142), .A2(n11079), .ZN(n11080) );
  INV_X1 U13507 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11181) );
  OR2_X1 U13508 ( .A1(n18868), .A2(n19125), .ZN(n12124) );
  OR2_X1 U13509 ( .A1(n12112), .A2(n18966), .ZN(n18994) );
  AND4_X1 U13510 ( .A1(n11978), .A2(n11977), .A3(n11976), .A4(n11975), .ZN(
        n11979) );
  OR2_X1 U13511 ( .A1(n12139), .A2(n12076), .ZN(n19879) );
  AND4_X1 U13512 ( .A1(n11895), .A2(n11894), .A3(n11893), .A4(n11892), .ZN(
        n11901) );
  AND4_X1 U13513 ( .A1(n11919), .A2(n11918), .A3(n11917), .A4(n11916), .ZN(
        n11920) );
  OR3_X1 U13514 ( .A1(n21087), .A2(n21674), .A3(n15766), .ZN(n15747) );
  NAND2_X1 U13515 ( .A1(n14752), .A2(n15043), .ZN(n14760) );
  AND2_X1 U13516 ( .A1(n15121), .A2(n15120), .ZN(n15584) );
  INV_X1 U13517 ( .A(n15043), .ZN(n15082) );
  AND2_X1 U13518 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n14322), .ZN(
        n14548) );
  NOR2_X1 U13519 ( .A1(n16174), .A2(n16165), .ZN(n16156) );
  INV_X1 U13520 ( .A(n16034), .ZN(n16044) );
  OR2_X1 U13521 ( .A1(n16301), .A2(n14539), .ZN(n17891) );
  INV_X1 U13522 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13745) );
  OR2_X1 U13523 ( .A1(n21365), .A2(n21492), .ZN(n21397) );
  NOR2_X1 U13524 ( .A1(n21190), .A2(n21189), .ZN(n21463) );
  INV_X1 U13525 ( .A(n21494), .ZN(n21499) );
  INV_X1 U13526 ( .A(n14670), .ZN(n14695) );
  AOI21_X1 U13527 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21422), .A(n21189), 
        .ZN(n21582) );
  NAND2_X1 U13528 ( .A1(n11195), .A2(n13389), .ZN(n11643) );
  INV_X1 U13529 ( .A(n20126), .ZN(n20182) );
  OR2_X1 U13530 ( .A1(n16453), .A2(n16485), .ZN(n11537) );
  NOR2_X1 U13531 ( .A1(n12491), .A2(n12492), .ZN(n16650) );
  INV_X1 U13532 ( .A(n14387), .ZN(n12192) );
  INV_X1 U13533 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17020) );
  INV_X1 U13534 ( .A(n17190), .ZN(n17175) );
  NAND2_X1 U13535 ( .A1(n13219), .A2(n11152), .ZN(n17187) );
  NAND2_X1 U13536 ( .A1(n16991), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16981) );
  AND3_X1 U13537 ( .A1(n11343), .A2(n11342), .A3(n11341), .ZN(n14624) );
  NAND2_X1 U13538 ( .A1(n10558), .A2(n10548), .ZN(n13917) );
  AND4_X1 U13539 ( .A1(n13913), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13914), 
        .A4(n17491), .ZN(n13915) );
  OR3_X1 U13540 ( .A1(n20622), .A2(n20644), .A3(n20939), .ZN(n20626) );
  NAND3_X1 U13541 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20958), .A3(n20697), 
        .ZN(n17489) );
  OR2_X1 U13542 ( .A1(n20628), .A2(n20506), .ZN(n20285) );
  INV_X1 U13543 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20939) );
  NOR2_X1 U13544 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18255), .ZN(n18233) );
  INV_X1 U13545 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19025) );
  INV_X1 U13546 ( .A(n13836), .ZN(n18635) );
  NAND2_X1 U13547 ( .A1(n14569), .A2(n18951), .ZN(n14570) );
  INV_X1 U13548 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19068) );
  AOI21_X1 U13549 ( .B1(n20034), .B2(n19400), .A(n19909), .ZN(n19414) );
  INV_X1 U13550 ( .A(n19688), .ZN(n19689) );
  OR2_X1 U13551 ( .A1(n13298), .A2(n20982), .ZN(n15389) );
  INV_X1 U13552 ( .A(n13618), .ZN(n20982) );
  AND2_X1 U13553 ( .A1(n15724), .A2(n15618), .ZN(n15682) );
  NOR2_X1 U13554 ( .A1(n15747), .A2(n15600), .ZN(n15724) );
  AND2_X2 U13555 ( .A1(n15453), .A2(n15452), .ZN(n21013) );
  AND2_X1 U13556 ( .A1(n21116), .A2(n14464), .ZN(n21112) );
  INV_X1 U13557 ( .A(n13933), .ZN(n21170) );
  INV_X1 U13558 ( .A(n15837), .ZN(n14436) );
  INV_X1 U13559 ( .A(n17885), .ZN(n17870) );
  NAND2_X1 U13560 ( .A1(n14747), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14753) );
  AND2_X1 U13561 ( .A1(n14321), .A2(n13887), .ZN(n21097) );
  INV_X1 U13562 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12894) );
  NAND2_X1 U13563 ( .A1(n16219), .A2(n13168), .ZN(n16292) );
  NOR2_X1 U13564 ( .A1(n17925), .A2(n16304), .ZN(n17910) );
  OAI22_X1 U13565 ( .A1(n21199), .A2(n21198), .B1(n21395), .B2(n21197), .ZN(
        n21222) );
  OAI211_X1 U13566 ( .C1(n21195), .C2(n21530), .A(n21463), .B(n21194), .ZN(
        n21223) );
  OR2_X1 U13567 ( .A1(n21186), .A2(n14665), .ZN(n21429) );
  OAI22_X1 U13568 ( .A1(n21261), .A2(n21260), .B1(n21259), .B2(n21395), .ZN(
        n21285) );
  OAI22_X1 U13569 ( .A1(n21301), .A2(n21300), .B1(n21641), .B2(n21299), .ZN(
        n21331) );
  INV_X1 U13570 ( .A(n21349), .ZN(n21357) );
  OR2_X1 U13571 ( .A1(n21186), .A2(n21185), .ZN(n21389) );
  NOR2_X2 U13572 ( .A1(n21365), .A2(n21429), .ZN(n21384) );
  OAI211_X1 U13573 ( .C1(n21586), .C2(n14714), .A(n14444), .B(n21582), .ZN(
        n14477) );
  INV_X1 U13574 ( .A(n21397), .ZN(n21418) );
  OAI221_X1 U13575 ( .B1(n21586), .B2(n21428), .C1(n21584), .C2(n21427), .A(
        n21582), .ZN(n21446) );
  NOR2_X2 U13576 ( .A1(n21499), .A2(n21429), .ZN(n21486) );
  NOR2_X2 U13577 ( .A1(n21499), .A2(n21451), .ZN(n21518) );
  INV_X1 U13578 ( .A(n21524), .ZN(n21564) );
  OAI21_X1 U13579 ( .B1(n14664), .B2(n14667), .A(n21582), .ZN(n14693) );
  NOR2_X2 U13580 ( .A1(n21581), .A2(n21429), .ZN(n16393) );
  NOR2_X2 U13581 ( .A1(n16117), .A2(n14436), .ZN(n14478) );
  AND2_X1 U13582 ( .A1(n21645), .A2(n12629), .ZN(n12917) );
  INV_X1 U13583 ( .A(n11643), .ZN(n11645) );
  INV_X1 U13584 ( .A(n20181), .ZN(n20167) );
  INV_X1 U13585 ( .A(n20165), .ZN(n20187) );
  OR2_X1 U13586 ( .A1(n11301), .A2(n11300), .ZN(n14564) );
  INV_X1 U13587 ( .A(n16752), .ZN(n16757) );
  NOR2_X1 U13588 ( .A1(n14344), .A2(n14335), .ZN(n13779) );
  INV_X1 U13589 ( .A(n16883), .ZN(n20227) );
  NOR2_X2 U13590 ( .A1(n20260), .A2(n20273), .ZN(n20272) );
  INV_X1 U13591 ( .A(n13270), .ZN(n20277) );
  INV_X2 U13592 ( .A(n13296), .ZN(n20281) );
  INV_X1 U13593 ( .A(n11162), .ZN(n11163) );
  NAND2_X1 U13594 ( .A1(n11417), .A2(n11416), .ZN(n11418) );
  INV_X1 U13595 ( .A(n14831), .ZN(n14832) );
  OAI21_X2 U13596 ( .B1(n17484), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n17483), 
        .ZN(n20697) );
  NAND2_X1 U13597 ( .A1(n20293), .A2(n20292), .ZN(n20320) );
  INV_X1 U13598 ( .A(n20417), .ZN(n20405) );
  NAND2_X1 U13599 ( .A1(n20921), .A2(n20931), .ZN(n20629) );
  INV_X1 U13600 ( .A(n20481), .ZN(n20470) );
  INV_X1 U13601 ( .A(n20482), .ZN(n20497) );
  NOR2_X2 U13602 ( .A1(n20506), .A2(n20424), .ZN(n20529) );
  INV_X1 U13603 ( .A(n20506), .ZN(n20501) );
  OAI21_X1 U13604 ( .B1(n20601), .B2(n20600), .A(n20599), .ZN(n20617) );
  AND2_X1 U13605 ( .A1(n20626), .A2(n20623), .ZN(n20645) );
  INV_X1 U13606 ( .A(n20697), .ZN(n20510) );
  INV_X1 U13607 ( .A(n20710), .ZN(n20776) );
  INV_X1 U13608 ( .A(n20688), .ZN(n20818) );
  NOR2_X1 U13609 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n18185), .ZN(n18171) );
  NOR2_X1 U13610 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18359), .ZN(n18338) );
  INV_X1 U13611 ( .A(n18437), .ZN(n18392) );
  INV_X1 U13612 ( .A(n18385), .ZN(n18441) );
  NAND2_X1 U13613 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n18620), .ZN(n18619) );
  NOR2_X1 U13614 ( .A1(n18635), .A2(n18749), .ZN(n18655) );
  AND2_X1 U13615 ( .A1(n18576), .A2(n13642), .ZN(n13836) );
  NOR2_X1 U13616 ( .A1(n13457), .A2(n13435), .ZN(n13544) );
  INV_X1 U13617 ( .A(n18793), .ZN(n18785) );
  OR2_X1 U13618 ( .A1(n19008), .A2(n18678), .ZN(n18985) );
  INV_X1 U13619 ( .A(n18985), .ZN(n18977) );
  NAND2_X1 U13620 ( .A1(n13194), .A2(n13193), .ZN(n19031) );
  AND2_X1 U13621 ( .A1(n19167), .A2(n19341), .ZN(n19192) );
  NOR2_X1 U13622 ( .A1(n19399), .A2(n19273), .ZN(n19301) );
  OR2_X1 U13623 ( .A1(n19318), .A2(n20031), .ZN(n19387) );
  INV_X1 U13624 ( .A(n19360), .ZN(n19396) );
  CLKBUF_X1 U13625 ( .A(n19517), .Z(n19505) );
  INV_X1 U13626 ( .A(n19556), .ZN(n19560) );
  INV_X1 U13627 ( .A(n19752), .ZN(n19756) );
  AND2_X1 U13628 ( .A1(n19801), .A2(BUF2_REG_21__SCAN_IN), .ZN(n19835) );
  INV_X1 U13629 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n20047) );
  INV_X1 U13630 ( .A(n20040), .ZN(n20032) );
  INV_X1 U13631 ( .A(n17490), .ZN(n17488) );
  INV_X1 U13632 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21426) );
  NAND2_X1 U13633 ( .A1(n15408), .A2(n15396), .ZN(n21086) );
  INV_X1 U13634 ( .A(n15994), .ZN(n15856) );
  INV_X1 U13635 ( .A(n16010), .ZN(n15864) );
  NAND2_X1 U13636 ( .A1(n13622), .A2(n13621), .ZN(n15899) );
  INV_X1 U13637 ( .A(n13826), .ZN(n21139) );
  INV_X1 U13638 ( .A(n21132), .ZN(n21151) );
  INV_X1 U13639 ( .A(n21169), .ZN(n13853) );
  NAND2_X1 U13640 ( .A1(n17885), .A2(n13714), .ZN(n17877) );
  INV_X1 U13641 ( .A(n17922), .ZN(n21174) );
  OR2_X2 U13642 ( .A1(n13149), .A2(n12982), .ZN(n21175) );
  OR2_X1 U13643 ( .A1(n21293), .A2(n21389), .ZN(n21251) );
  OR2_X1 U13644 ( .A1(n21293), .A2(n21429), .ZN(n21283) );
  OR2_X1 U13645 ( .A1(n21293), .A2(n21451), .ZN(n21335) );
  OR2_X1 U13646 ( .A1(n21293), .A2(n21492), .ZN(n21349) );
  OR2_X1 U13647 ( .A1(n21365), .A2(n21389), .ZN(n21388) );
  AOI22_X1 U13648 ( .A1(n14717), .A2(n14713), .B1(n21190), .B2(n21258), .ZN(
        n14746) );
  OR2_X1 U13649 ( .A1(n21365), .A2(n21451), .ZN(n14742) );
  NAND2_X1 U13650 ( .A1(n21494), .A2(n21390), .ZN(n21449) );
  AOI22_X1 U13651 ( .A1(n21460), .A2(n21457), .B1(n21456), .B2(n21455), .ZN(
        n21491) );
  NAND2_X1 U13652 ( .A1(n21494), .A2(n21493), .ZN(n21569) );
  NAND2_X1 U13653 ( .A1(n14660), .A2(n14665), .ZN(n21524) );
  INV_X1 U13654 ( .A(n21632), .ZN(n16396) );
  OR2_X1 U13655 ( .A1(n21581), .A2(n21492), .ZN(n21636) );
  INV_X1 U13656 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21638) );
  INV_X1 U13657 ( .A(n21730), .ZN(n21726) );
  INV_X1 U13658 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n21661) );
  INV_X1 U13659 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n21694) );
  INV_X1 U13660 ( .A(n21755), .ZN(n21716) );
  NAND2_X1 U13661 ( .A1(n21657), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21755) );
  NAND2_X1 U13662 ( .A1(n20190), .A2(n13221), .ZN(n20053) );
  INV_X1 U13663 ( .A(n11667), .ZN(n11668) );
  INV_X1 U13664 ( .A(n20107), .ZN(n17819) );
  NAND2_X1 U13665 ( .A1(n20053), .A2(n11646), .ZN(n20189) );
  NOR2_X1 U13666 ( .A1(n13779), .A2(n14802), .ZN(n20207) );
  INV_X1 U13667 ( .A(n20931), .ZN(n20912) );
  OR2_X1 U13668 ( .A1(n16730), .A2(n16729), .ZN(n16846) );
  AND2_X1 U13669 ( .A1(n16850), .A2(n13873), .ZN(n20232) );
  INV_X1 U13670 ( .A(n20272), .ZN(n20271) );
  OR2_X1 U13671 ( .A1(n13221), .A2(n16694), .ZN(n13296) );
  NOR2_X1 U13672 ( .A1(n11164), .A2(n11163), .ZN(n11165) );
  INV_X1 U13673 ( .A(n17196), .ZN(n17139) );
  AOI211_X1 U13674 ( .C1(n14923), .C2(n17454), .A(n14922), .B(n14921), .ZN(
        n14924) );
  INV_X1 U13675 ( .A(n17454), .ZN(n17415) );
  AND2_X1 U13676 ( .A1(n20328), .A2(n20327), .ZN(n20339) );
  NAND2_X1 U13677 ( .A1(n20356), .A2(n20913), .ZN(n20417) );
  OR2_X1 U13678 ( .A1(n20500), .A2(n20629), .ZN(n20443) );
  OR2_X1 U13679 ( .A1(n20424), .A2(n20695), .ZN(n20481) );
  INV_X1 U13680 ( .A(n10555), .ZN(n20621) );
  INV_X1 U13681 ( .A(n10564), .ZN(n20649) );
  INV_X1 U13682 ( .A(n20656), .ZN(n20725) );
  AOI211_X2 U13683 ( .C1(n17506), .C2(n17505), .A(n20510), .B(n17504), .ZN(
        n20752) );
  AOI211_X2 U13684 ( .C1(n17517), .C2(n17518), .A(n17521), .B(n17516), .ZN(
        n20825) );
  INV_X1 U13685 ( .A(n20909), .ZN(n20828) );
  OR2_X1 U13686 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20839), .ZN(n20976) );
  INV_X1 U13687 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18037) );
  OR2_X1 U13688 ( .A1(n20049), .A2(n14239), .ZN(n18437) );
  NAND2_X1 U13689 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18441), .ZN(n18435) );
  AND2_X1 U13690 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n13627), .ZN(n13711) );
  NOR2_X1 U13691 ( .A1(n18636), .A2(n13435), .ZN(n18659) );
  INV_X1 U13692 ( .A(n18703), .ZN(n18708) );
  OR2_X1 U13693 ( .A1(n20041), .A2(n18738), .ZN(n18733) );
  INV_X1 U13694 ( .A(n18791), .ZN(n18787) );
  INV_X1 U13695 ( .A(n18847), .ZN(n18933) );
  INV_X1 U13696 ( .A(n19015), .ZN(n19034) );
  INV_X1 U13697 ( .A(n19122), .ZN(n19084) );
  NAND2_X1 U13698 ( .A1(n18041), .A2(n12117), .ZN(n19116) );
  INV_X1 U13699 ( .A(n19297), .ZN(n19311) );
  INV_X1 U13700 ( .A(n19341), .ZN(n19399) );
  INV_X1 U13701 ( .A(n19583), .ZN(n19579) );
  INV_X1 U13702 ( .A(n19657), .ZN(n19844) );
  INV_X1 U13703 ( .A(n18414), .ZN(n19923) );
  INV_X1 U13704 ( .A(n20014), .ZN(n20011) );
  INV_X1 U13705 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19947) );
  NOR2_X1 U13706 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13189), .ZN(n18016)
         );
  INV_X1 U13707 ( .A(n17992), .ZN(n17989) );
  OAI211_X1 U13708 ( .C1(n14909), .C2(n12497), .A(n12496), .B(n12495), .ZN(
        P2_U2890) );
  INV_X1 U13709 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10567) );
  AND2_X2 U13710 ( .A1(n10567), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10568) );
  AND2_X4 U13711 ( .A1(n10568), .A2(n10575), .ZN(n12379) );
  AOI22_X1 U13712 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10572) );
  AND2_X4 U13713 ( .A1(n10568), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12316) );
  AOI22_X1 U13715 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10571) );
  INV_X2 U13716 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14811) );
  AND3_X4 U13717 ( .A1(n10575), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        n14811), .ZN(n12325) );
  AOI22_X1 U13718 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10570) );
  NOR2_X4 U13719 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14370) );
  AND2_X4 U13720 ( .A1(n14370), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12324) );
  AOI22_X1 U13721 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10569) );
  AND2_X2 U13722 ( .A1(n12324), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10921) );
  AND2_X2 U13723 ( .A1(n10697), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10926) );
  AOI22_X1 U13724 ( .A1(n10921), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10579) );
  AND2_X4 U13725 ( .A1(n14331), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12318) );
  INV_X2 U13726 ( .A(n10554), .ZN(n12309) );
  AND2_X2 U13727 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10574) );
  AND2_X4 U13728 ( .A1(n10574), .A2(n10575), .ZN(n12317) );
  AOI22_X1 U13730 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10578) );
  INV_X1 U13731 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10573) );
  AOI22_X1 U13733 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10577) );
  AND2_X2 U13734 ( .A1(n11054), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12356) );
  AND2_X2 U13735 ( .A1(n12319), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10797) );
  AOI22_X1 U13736 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10576) );
  NAND2_X1 U13737 ( .A1(n20938), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10581) );
  NAND2_X1 U13738 ( .A1(n14358), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10580) );
  NAND2_X1 U13739 ( .A1(n10581), .A2(n10580), .ZN(n11172) );
  NAND2_X1 U13740 ( .A1(n14811), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10583) );
  OAI21_X1 U13741 ( .B1(n10585), .B2(n10584), .A(n10874), .ZN(n11170) );
  INV_X1 U13742 ( .A(n11170), .ZN(n11166) );
  AOI22_X1 U13743 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12324), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10587) );
  AOI22_X1 U13744 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12325), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10586) );
  AOI22_X1 U13745 ( .A1(n9696), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12318), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U13746 ( .A1(n12319), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12317), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10591) );
  AOI22_X1 U13747 ( .A1(n9696), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12318), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10594) );
  AOI22_X1 U13748 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12325), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U13749 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12324), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10592) );
  AOI22_X1 U13750 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12324), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10601) );
  AOI22_X1 U13751 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12325), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10600) );
  AOI22_X1 U13752 ( .A1(n10697), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12317), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10599) );
  AOI22_X1 U13753 ( .A1(n12318), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12319), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10598) );
  AOI22_X1 U13754 ( .A1(n10697), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12318), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10605) );
  AOI22_X1 U13755 ( .A1(n12319), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12317), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10604) );
  AOI22_X1 U13756 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12324), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U13757 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12325), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10602) );
  INV_X1 U13758 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n16619) );
  AOI22_X1 U13759 ( .A1(n9696), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12318), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U13760 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12325), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10609) );
  AOI22_X1 U13761 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12324), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10608) );
  AOI22_X1 U13762 ( .A1(n12319), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12317), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10607) );
  NAND4_X1 U13763 ( .A1(n10610), .A2(n10609), .A3(n10608), .A4(n10607), .ZN(
        n10611) );
  AOI22_X1 U13764 ( .A1(n9696), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12318), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U13765 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12325), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10614) );
  AOI22_X1 U13766 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12324), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10613) );
  AOI22_X1 U13767 ( .A1(n12319), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12317), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10612) );
  NAND4_X1 U13768 ( .A1(n10615), .A2(n10614), .A3(n10613), .A4(n10612), .ZN(
        n10616) );
  AOI22_X1 U13769 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10802), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10623) );
  AOI22_X1 U13770 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10622) );
  AOI22_X1 U13771 ( .A1(n10803), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10621) );
  AOI22_X1 U13772 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10804), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10620) );
  NAND4_X1 U13773 ( .A1(n10623), .A2(n10622), .A3(n10621), .A4(n10620), .ZN(
        n10631) );
  AOI22_X1 U13774 ( .A1(n10921), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10629) );
  AOI22_X1 U13775 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10628) );
  AOI22_X1 U13776 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10627) );
  AOI22_X1 U13777 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10626) );
  NAND4_X1 U13778 ( .A1(n10629), .A2(n10628), .A3(n10627), .A4(n10626), .ZN(
        n10630) );
  NAND2_X1 U13779 ( .A1(n10878), .A2(n11062), .ZN(n11213) );
  NOR2_X1 U13780 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10632) );
  NAND2_X1 U13781 ( .A1(n11207), .A2(n10632), .ZN(n10633) );
  NAND2_X1 U13782 ( .A1(n11213), .A2(n10633), .ZN(n10644) );
  OAI21_X1 U13783 ( .B1(n10634), .B2(n10644), .A(n10882), .ZN(n16623) );
  INV_X1 U13784 ( .A(n16623), .ZN(n10646) );
  XNOR2_X1 U13785 ( .A(n16623), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14265) );
  AOI22_X1 U13786 ( .A1(n10921), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10638) );
  AOI22_X1 U13787 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10637) );
  AOI22_X1 U13788 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12309), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10636) );
  AOI22_X1 U13789 ( .A1(n10624), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10635) );
  AOI22_X1 U13790 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10642) );
  AOI22_X1 U13791 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10641) );
  AOI22_X1 U13792 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10640) );
  AOI22_X1 U13793 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10639) );
  OAI21_X1 U13794 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20947), .A(
        n11046), .ZN(n11173) );
  INV_X1 U13795 ( .A(n11173), .ZN(n11168) );
  MUX2_X1 U13796 ( .A(n13917), .B(n11168), .S(n10876), .Z(n11033) );
  MUX2_X1 U13797 ( .A(n11033), .B(P2_EBX_REG_0__SCAN_IN), .S(n11473), .Z(
        n16641) );
  NAND2_X1 U13798 ( .A1(n16641), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13340) );
  AND2_X1 U13799 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13990) );
  NAND2_X1 U13800 ( .A1(n16641), .A2(n13990), .ZN(n10645) );
  INV_X1 U13801 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14247) );
  AND3_X1 U13802 ( .A1(n11473), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n10643) );
  OR2_X1 U13803 ( .A1(n10644), .A2(n10643), .ZN(n16628) );
  AOI22_X1 U13804 ( .A1(n13332), .A2(n13340), .B1(n10645), .B2(n16628), .ZN(
        n14264) );
  NAND2_X1 U13805 ( .A1(n14265), .A2(n14264), .ZN(n17192) );
  INV_X1 U13806 ( .A(n17192), .ZN(n14266) );
  AOI21_X1 U13807 ( .B1(n10646), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n14266), .ZN(n17170) );
  AOI22_X1 U13808 ( .A1(n9696), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12318), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10650) );
  AOI22_X1 U13809 ( .A1(n12319), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12317), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10649) );
  AOI22_X1 U13810 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12324), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U13811 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12325), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10647) );
  AOI22_X1 U13812 ( .A1(n9696), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12318), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10654) );
  AOI22_X1 U13813 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12324), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13814 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12325), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10651) );
  AOI22_X1 U13815 ( .A1(n9696), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12318), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U13816 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12325), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U13817 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12324), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10656) );
  NAND4_X1 U13818 ( .A1(n10658), .A2(n10657), .A3(n10656), .A4(n10655), .ZN(
        n10659) );
  AOI22_X1 U13819 ( .A1(n9696), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12318), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10663) );
  AOI22_X1 U13820 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12325), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10661) );
  AOI22_X1 U13821 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12324), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10660) );
  NAND4_X1 U13822 ( .A1(n10663), .A2(n10662), .A3(n10661), .A4(n10660), .ZN(
        n10664) );
  NAND2_X1 U13823 ( .A1(n10664), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10665) );
  AOI22_X1 U13824 ( .A1(n9696), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12318), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10670) );
  AOI22_X1 U13825 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12325), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10669) );
  AOI22_X1 U13826 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12324), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U13827 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12319), .B1(
        n12317), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10667) );
  NAND4_X1 U13828 ( .A1(n10670), .A2(n10669), .A3(n10668), .A4(n10667), .ZN(
        n10671) );
  AOI22_X1 U13829 ( .A1(n9696), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12318), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10675) );
  AOI22_X1 U13830 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12325), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U13831 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12324), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10672) );
  NAND4_X1 U13832 ( .A1(n10675), .A2(n10674), .A3(n10673), .A4(n10672), .ZN(
        n10676) );
  XNOR2_X1 U13833 ( .A(n9809), .B(n12243), .ZN(n11188) );
  NAND2_X1 U13834 ( .A1(n11188), .A2(n9921), .ZN(n11191) );
  NAND2_X1 U13835 ( .A1(n10677), .A2(n11191), .ZN(n11380) );
  AOI22_X1 U13836 ( .A1(n10697), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12318), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U13837 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12325), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U13838 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12324), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U13839 ( .A1(n12319), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12317), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10678) );
  NAND4_X1 U13840 ( .A1(n10681), .A2(n10680), .A3(n10679), .A4(n10678), .ZN(
        n10689) );
  AOI22_X1 U13841 ( .A1(n10697), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12318), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U13842 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12325), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U13843 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12324), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10685) );
  NAND2_X1 U13844 ( .A1(n12317), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10683) );
  NAND4_X1 U13845 ( .A1(n10687), .A2(n10686), .A3(n10685), .A4(n10684), .ZN(
        n10688) );
  NAND2_X1 U13846 ( .A1(n11380), .A2(n11382), .ZN(n10693) );
  NAND2_X1 U13847 ( .A1(n10693), .A2(n10692), .ZN(n10696) );
  NAND2_X1 U13848 ( .A1(n10726), .A2(n9989), .ZN(n11384) );
  NAND2_X1 U13849 ( .A1(n9937), .A2(n10694), .ZN(n10695) );
  AOI22_X1 U13850 ( .A1(n10697), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12318), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U13851 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12325), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10700) );
  AOI22_X1 U13852 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12324), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U13853 ( .A1(n12319), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12317), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10698) );
  NAND4_X1 U13854 ( .A1(n10701), .A2(n10700), .A3(n10699), .A4(n10698), .ZN(
        n10702) );
  NAND2_X1 U13855 ( .A1(n10702), .A2(n14353), .ZN(n10708) );
  AOI22_X1 U13856 ( .A1(n9696), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12318), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10706) );
  AOI22_X1 U13857 ( .A1(n12316), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12325), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10705) );
  AOI22_X1 U13858 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12324), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10704) );
  NAND4_X1 U13859 ( .A1(n10706), .A2(n10705), .A3(n10704), .A4(n10703), .ZN(
        n10707) );
  NAND2_X1 U13860 ( .A1(n10726), .A2(n11382), .ZN(n10716) );
  MUX2_X1 U13861 ( .A(n12243), .B(n11208), .S(n10712), .Z(n10715) );
  NAND2_X1 U13862 ( .A1(n10753), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10725) );
  AND2_X1 U13863 ( .A1(n17495), .A2(n11388), .ZN(n10720) );
  INV_X2 U13864 ( .A(n10722), .ZN(n11195) );
  NAND2_X1 U13865 ( .A1(n10728), .A2(n11643), .ZN(n11412) );
  NAND2_X1 U13866 ( .A1(n11195), .A2(n11651), .ZN(n10727) );
  AND2_X4 U13867 ( .A1(n11195), .A2(n10729), .ZN(n11555) );
  AOI22_X1 U13868 ( .A1(n11555), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10732) );
  NAND2_X1 U13869 ( .A1(n11092), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10731) );
  INV_X1 U13870 ( .A(n10753), .ZN(n10744) );
  INV_X1 U13871 ( .A(n10733), .ZN(n10734) );
  NAND2_X1 U13872 ( .A1(n10744), .A2(n10734), .ZN(n10736) );
  INV_X1 U13873 ( .A(n11092), .ZN(n11102) );
  NAND2_X1 U13874 ( .A1(n11102), .A2(n14354), .ZN(n10735) );
  NAND2_X1 U13875 ( .A1(n10736), .A2(n10735), .ZN(n10739) );
  INV_X1 U13876 ( .A(n20959), .ZN(n10741) );
  OAI22_X1 U13877 ( .A1(n14333), .A2(n11573), .B1(n20947), .B2(n10741), .ZN(
        n10737) );
  INV_X1 U13878 ( .A(n10737), .ZN(n10738) );
  BUF_X4 U13879 ( .A(n10756), .Z(n11091) );
  INV_X1 U13880 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n11060) );
  NAND2_X1 U13881 ( .A1(n11092), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10743) );
  NAND2_X1 U13882 ( .A1(n11555), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10742) );
  NAND2_X1 U13883 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10740) );
  NAND2_X1 U13884 ( .A1(n10753), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10748) );
  AOI21_X1 U13885 ( .B1(n11573), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10747) );
  INV_X1 U13886 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10751) );
  NAND2_X1 U13887 ( .A1(n11555), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10750) );
  NAND2_X1 U13888 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10749) );
  NOR2_X1 U13889 ( .A1(n10765), .A2(n11096), .ZN(n10759) );
  INV_X1 U13890 ( .A(n10759), .ZN(n10758) );
  INV_X1 U13891 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U13892 ( .A1(n11555), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10755) );
  NAND2_X1 U13893 ( .A1(n11092), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10754) );
  INV_X1 U13894 ( .A(n10761), .ZN(n10764) );
  XNOR2_X2 U13895 ( .A(n11099), .B(n10766), .ZN(n10781) );
  BUF_X4 U13896 ( .A(n10781), .Z(n14582) );
  AOI22_X1 U13897 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20393), .B1(
        n20622), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10779) );
  INV_X1 U13898 ( .A(n10767), .ZN(n10769) );
  NAND2_X1 U13899 ( .A1(n10769), .A2(n17455), .ZN(n10771) );
  NOR2_X1 U13900 ( .A1(n10770), .A2(n14582), .ZN(n10911) );
  AOI22_X1 U13901 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10911), .B1(
        n10812), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10778) );
  INV_X1 U13902 ( .A(n10771), .ZN(n10772) );
  AOI22_X1 U13903 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20689), .B1(
        n10910), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10777) );
  NOR2_X2 U13904 ( .A1(n10774), .A2(n14582), .ZN(n10912) );
  AND2_X2 U13905 ( .A1(n10788), .A2(n10783), .ZN(n10917) );
  AOI22_X1 U13906 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20291), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10786) );
  AND2_X2 U13907 ( .A1(n10788), .A2(n10784), .ZN(n20537) );
  AOI22_X1 U13908 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20361), .B1(
        n20537), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10785) );
  INV_X1 U13909 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10791) );
  INV_X1 U13910 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10790) );
  OAI22_X1 U13911 ( .A1(n10900), .A2(n10791), .B1(n10947), .B2(n10790), .ZN(
        n10796) );
  INV_X1 U13912 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10794) );
  INV_X1 U13913 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10793) );
  OAI22_X1 U13914 ( .A1(n20655), .A2(n10794), .B1(n10903), .B2(n10793), .ZN(
        n10795) );
  AOI22_X1 U13915 ( .A1(n10849), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10801) );
  AOI22_X1 U13916 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10800) );
  AOI22_X1 U13917 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10799) );
  AOI22_X1 U13918 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10798) );
  NAND4_X1 U13919 ( .A1(n10801), .A2(n10800), .A3(n10799), .A4(n10798), .ZN(
        n10810) );
  AOI22_X1 U13920 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U13921 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U13922 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U13923 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10921), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10805) );
  NAND4_X1 U13924 ( .A1(n10808), .A2(n10807), .A3(n10806), .A4(n10805), .ZN(
        n10809) );
  NAND2_X1 U13925 ( .A1(n9989), .A2(n10877), .ZN(n10811) );
  INV_X1 U13926 ( .A(n10841), .ZN(n10839) );
  INV_X1 U13927 ( .A(n10812), .ZN(n10815) );
  INV_X1 U13928 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10814) );
  NAND2_X1 U13929 ( .A1(n10917), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10813) );
  OAI211_X1 U13930 ( .C1(n10815), .C2(n10814), .A(n10813), .B(n16694), .ZN(
        n10819) );
  NOR2_X1 U13931 ( .A1(n10819), .A2(n10818), .ZN(n10836) );
  INV_X1 U13932 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10823) );
  NAND2_X1 U13933 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10821) );
  OAI211_X1 U13934 ( .C1(n10947), .C2(n10823), .A(n10822), .B(n10821), .ZN(
        n10827) );
  INV_X1 U13935 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10825) );
  INV_X1 U13936 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10824) );
  OAI22_X1 U13937 ( .A1(n10903), .A2(n10825), .B1(n20655), .B2(n10824), .ZN(
        n10826) );
  NOR2_X1 U13938 ( .A1(n10827), .A2(n10826), .ZN(n10835) );
  AOI22_X1 U13939 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10912), .B1(
        n10910), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10830) );
  AOI22_X1 U13940 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20689), .B1(
        n20622), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10829) );
  AOI22_X1 U13941 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10911), .B1(
        n20393), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10828) );
  NAND3_X1 U13942 ( .A1(n10830), .A2(n10829), .A3(n10828), .ZN(n10833) );
  INV_X1 U13943 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10831) );
  NOR2_X1 U13944 ( .A1(n10900), .A2(n10831), .ZN(n10832) );
  NOR2_X1 U13945 ( .A1(n10833), .A2(n10832), .ZN(n10834) );
  NAND3_X1 U13946 ( .A1(n13223), .A2(n13917), .A3(n11062), .ZN(n11066) );
  INV_X1 U13947 ( .A(n10837), .ZN(n11222) );
  NAND2_X1 U13948 ( .A1(n11066), .A2(n11222), .ZN(n10838) );
  NAND2_X1 U13949 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10846) );
  NAND2_X1 U13950 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10845) );
  NAND2_X1 U13951 ( .A1(n10803), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10844) );
  NAND2_X1 U13952 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10843) );
  NAND2_X1 U13953 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10855) );
  NAND2_X1 U13954 ( .A1(n10618), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10854) );
  INV_X1 U13955 ( .A(n12340), .ZN(n10848) );
  INV_X1 U13956 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10847) );
  OR2_X1 U13957 ( .A1(n10848), .A2(n10847), .ZN(n10853) );
  INV_X1 U13958 ( .A(n10849), .ZN(n10851) );
  INV_X1 U13959 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10850) );
  OR2_X1 U13960 ( .A1(n10851), .A2(n10850), .ZN(n10852) );
  INV_X1 U13961 ( .A(n10921), .ZN(n10857) );
  INV_X1 U13962 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10856) );
  OR2_X1 U13963 ( .A1(n10857), .A2(n10856), .ZN(n10863) );
  INV_X1 U13964 ( .A(n10926), .ZN(n10859) );
  INV_X1 U13965 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10858) );
  OR2_X1 U13966 ( .A1(n10859), .A2(n10858), .ZN(n10862) );
  NAND2_X1 U13967 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10861) );
  NAND2_X1 U13968 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10860) );
  NAND2_X1 U13969 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10867) );
  NAND2_X1 U13970 ( .A1(n10624), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10866) );
  NAND2_X1 U13971 ( .A1(n10625), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10865) );
  NAND2_X1 U13972 ( .A1(n10797), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10864) );
  XNOR2_X1 U13973 ( .A(n10895), .B(n10894), .ZN(n11048) );
  OAI21_X1 U13974 ( .B1(n10877), .B2(n10876), .A(n10875), .ZN(n11036) );
  NAND2_X1 U13975 ( .A1(n10882), .A2(n10881), .ZN(n10883) );
  NAND2_X1 U13976 ( .A1(n9899), .A2(n10883), .ZN(n16601) );
  AOI22_X1 U13977 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10887) );
  AOI22_X1 U13978 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10886) );
  AOI22_X1 U13979 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10885) );
  AOI22_X1 U13980 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10921), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10884) );
  NAND4_X1 U13981 ( .A1(n10887), .A2(n10886), .A3(n10885), .A4(n10884), .ZN(
        n10893) );
  AOI22_X1 U13982 ( .A1(n10849), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U13983 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10890) );
  AOI22_X1 U13984 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10889) );
  AOI22_X1 U13985 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10888) );
  NAND4_X1 U13986 ( .A1(n10891), .A2(n10890), .A3(n10889), .A4(n10888), .ZN(
        n10892) );
  NAND2_X1 U13987 ( .A1(n10895), .A2(n10894), .ZN(n10897) );
  NAND2_X1 U13988 ( .A1(n20920), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10896) );
  NAND2_X1 U13989 ( .A1(n10897), .A2(n10896), .ZN(n11041) );
  NAND2_X1 U13990 ( .A1(n11181), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11042) );
  MUX2_X1 U13991 ( .A(n11072), .B(n11049), .S(n10876), .Z(n11038) );
  INV_X1 U13992 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n11105) );
  MUX2_X1 U13993 ( .A(n11038), .B(n11105), .S(n11473), .Z(n10935) );
  XNOR2_X1 U13994 ( .A(n10936), .B(n10935), .ZN(n10898) );
  XNOR2_X1 U13995 ( .A(n10898), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17157) );
  INV_X1 U13996 ( .A(n10898), .ZN(n20188) );
  INV_X1 U13997 ( .A(n11072), .ZN(n10899) );
  INV_X1 U13998 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10902) );
  INV_X1 U13999 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10901) );
  OAI22_X1 U14000 ( .A1(n10900), .A2(n10902), .B1(n10947), .B2(n10901), .ZN(
        n10908) );
  INV_X1 U14001 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10906) );
  INV_X1 U14002 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10905) );
  OAI22_X1 U14003 ( .A1(n10903), .A2(n10906), .B1(n20655), .B2(n10905), .ZN(
        n10907) );
  NOR2_X1 U14004 ( .A1(n10908), .A2(n10907), .ZN(n10920) );
  AOI22_X1 U14005 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n10909), .B1(
        n20393), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U14006 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n10910), .B1(
        n20622), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U14007 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20456), .B1(
        n20689), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10914) );
  AOI22_X1 U14008 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n10912), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10913) );
  AOI22_X1 U14009 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n10917), .B1(
        n20537), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10919) );
  AOI22_X1 U14010 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20361), .B1(
        n20291), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10918) );
  AOI22_X1 U14011 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10925) );
  AOI22_X1 U14012 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U14013 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U14014 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10921), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10922) );
  NAND4_X1 U14015 ( .A1(n10925), .A2(n10924), .A3(n10923), .A4(n10922), .ZN(
        n10932) );
  AOI22_X1 U14016 ( .A1(n10849), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10930) );
  AOI22_X1 U14017 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U14018 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U14019 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10927) );
  NAND4_X1 U14020 ( .A1(n10930), .A2(n10929), .A3(n10928), .A4(n10927), .ZN(
        n10931) );
  INV_X1 U14021 ( .A(n10937), .ZN(n11243) );
  NAND2_X1 U14022 ( .A1(n11243), .A2(n13223), .ZN(n10933) );
  INV_X1 U14023 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n14613) );
  MUX2_X1 U14024 ( .A(n10937), .B(n14613), .S(n11473), .Z(n10938) );
  OAI21_X1 U14025 ( .B1(n10939), .B2(n10938), .A(n10968), .ZN(n14784) );
  INV_X1 U14026 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17423) );
  AOI22_X1 U14027 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20393), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U14028 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20456), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U14029 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20622), .B1(
        n10910), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U14030 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20689), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10941) );
  NAND2_X1 U14031 ( .A1(n10945), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10951) );
  INV_X1 U14032 ( .A(n10903), .ZN(n10946) );
  NAND2_X1 U14033 ( .A1(n10946), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10950) );
  INV_X1 U14034 ( .A(n20655), .ZN(n20652) );
  NAND2_X1 U14035 ( .A1(n20652), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10949) );
  NAND2_X1 U14036 ( .A1(n17503), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10948) );
  AOI22_X1 U14037 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20361), .B1(
        n20291), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10953) );
  AOI22_X1 U14038 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n10917), .B1(
        n20537), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10952) );
  NAND4_X1 U14039 ( .A1(n10954), .A2(n9776), .A3(n10953), .A4(n10952), .ZN(
        n10966) );
  AOI22_X1 U14040 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10958) );
  AOI22_X1 U14041 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U14042 ( .A1(n10803), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10804), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10956) );
  AOI22_X1 U14043 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10955) );
  NAND4_X1 U14044 ( .A1(n10958), .A2(n10957), .A3(n10956), .A4(n10955), .ZN(
        n10964) );
  AOI22_X1 U14045 ( .A1(n10921), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10962) );
  AOI22_X1 U14046 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12356), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U14047 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U14048 ( .A1(n10625), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10959) );
  NAND4_X1 U14049 ( .A1(n10962), .A2(n10961), .A3(n10960), .A4(n10959), .ZN(
        n10963) );
  NAND2_X1 U14050 ( .A1(n11247), .A2(n13223), .ZN(n10965) );
  MUX2_X1 U14051 ( .A(n11247), .B(P2_EBX_REG_6__SCAN_IN), .S(n11473), .Z(
        n10967) );
  XNOR2_X1 U14052 ( .A(n10968), .B(n10967), .ZN(n16592) );
  INV_X1 U14053 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17405) );
  INV_X1 U14054 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10969) );
  MUX2_X1 U14055 ( .A(n11477), .B(n10969), .S(n11473), .Z(n10974) );
  NAND2_X1 U14056 ( .A1(n10975), .A2(n10974), .ZN(n10970) );
  NAND2_X1 U14057 ( .A1(n10970), .A2(n10971), .ZN(n10972) );
  NAND2_X1 U14058 ( .A1(n10978), .A2(n10972), .ZN(n16578) );
  OR2_X1 U14059 ( .A1(n16578), .A2(n11482), .ZN(n10994) );
  INV_X1 U14060 ( .A(n10994), .ZN(n10973) );
  NAND2_X1 U14061 ( .A1(n10973), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17111) );
  OR2_X1 U14062 ( .A1(n10975), .A2(n10974), .ZN(n10976) );
  NAND2_X1 U14063 ( .A1(n10970), .A2(n10976), .ZN(n20166) );
  INV_X1 U14064 ( .A(n20166), .ZN(n10977) );
  NAND2_X1 U14065 ( .A1(n10977), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17123) );
  AND2_X1 U14066 ( .A1(n17111), .A2(n17123), .ZN(n17081) );
  INV_X1 U14067 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n14429) );
  INV_X1 U14068 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n14568) );
  NAND2_X1 U14069 ( .A1(n11473), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10980) );
  NOR2_X1 U14070 ( .A1(n10979), .A2(n10980), .ZN(n10981) );
  OR2_X1 U14071 ( .A1(n10988), .A2(n10981), .ZN(n16566) );
  OR2_X1 U14072 ( .A1(n16566), .A2(n11482), .ZN(n10996) );
  INV_X1 U14073 ( .A(n10996), .ZN(n10982) );
  NAND2_X1 U14074 ( .A1(n10982), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17066) );
  NAND2_X1 U14075 ( .A1(n11473), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10983) );
  OAI21_X1 U14076 ( .B1(n9807), .B2(n10983), .A(n11456), .ZN(n10984) );
  OR2_X1 U14077 ( .A1(n10984), .A2(n10979), .ZN(n20134) );
  INV_X1 U14078 ( .A(n20134), .ZN(n10986) );
  AND2_X1 U14079 ( .A1(n11477), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10985) );
  NAND2_X1 U14080 ( .A1(n10986), .A2(n10985), .ZN(n17085) );
  NAND2_X1 U14081 ( .A1(n11473), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10987) );
  XNOR2_X1 U14082 ( .A(n10978), .B(n10987), .ZN(n20151) );
  NAND2_X1 U14083 ( .A1(n20151), .A2(n11477), .ZN(n10995) );
  INV_X1 U14084 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17348) );
  OR2_X1 U14085 ( .A1(n10995), .A2(n17348), .ZN(n17096) );
  AND2_X1 U14086 ( .A1(n17085), .A2(n17096), .ZN(n17062) );
  NAND2_X1 U14087 ( .A1(n17066), .A2(n17062), .ZN(n17050) );
  NAND2_X1 U14088 ( .A1(n11473), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10989) );
  INV_X1 U14089 ( .A(n10989), .ZN(n10990) );
  NAND2_X1 U14090 ( .A1(n10991), .A2(n10990), .ZN(n10992) );
  NAND2_X1 U14091 ( .A1(n11000), .A2(n10992), .ZN(n16550) );
  OR2_X1 U14092 ( .A1(n16550), .A2(n11482), .ZN(n10993) );
  INV_X1 U14093 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17329) );
  NOR2_X1 U14094 ( .A1(n10993), .A2(n17329), .ZN(n17051) );
  OR2_X1 U14095 ( .A1(n17050), .A2(n17051), .ZN(n11433) );
  NAND2_X1 U14096 ( .A1(n10993), .A2(n17329), .ZN(n17052) );
  INV_X1 U14097 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17361) );
  OAI21_X1 U14098 ( .B1(n20134), .B2(n11482), .A(n17361), .ZN(n17086) );
  INV_X1 U14099 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17384) );
  NAND2_X1 U14100 ( .A1(n10994), .A2(n17384), .ZN(n17110) );
  INV_X1 U14101 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17397) );
  NAND2_X1 U14102 ( .A1(n20166), .A2(n17397), .ZN(n17122) );
  AND2_X1 U14103 ( .A1(n17110), .A2(n17122), .ZN(n17082) );
  NAND2_X1 U14104 ( .A1(n10995), .A2(n17348), .ZN(n17095) );
  AND3_X1 U14105 ( .A1(n17086), .A2(n17082), .A3(n17095), .ZN(n17047) );
  INV_X1 U14106 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17349) );
  NAND2_X1 U14107 ( .A1(n10996), .A2(n17349), .ZN(n17065) );
  AND3_X1 U14108 ( .A1(n17052), .A2(n17047), .A3(n17065), .ZN(n11426) );
  XNOR2_X1 U14109 ( .A(n11000), .B(n10552), .ZN(n16543) );
  NAND2_X1 U14110 ( .A1(n16543), .A2(n11477), .ZN(n10999) );
  INV_X1 U14111 ( .A(n10999), .ZN(n10998) );
  INV_X1 U14112 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17318) );
  NAND2_X1 U14113 ( .A1(n10999), .A2(n17318), .ZN(n17039) );
  XNOR2_X1 U14114 ( .A(n11003), .B(n9846), .ZN(n20123) );
  NAND2_X1 U14115 ( .A1(n20123), .A2(n11477), .ZN(n11001) );
  INV_X1 U14116 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17308) );
  NAND2_X1 U14117 ( .A1(n11001), .A2(n17308), .ZN(n17027) );
  AND2_X1 U14118 ( .A1(n11477), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11002) );
  NAND2_X1 U14119 ( .A1(n20123), .A2(n11002), .ZN(n17026) );
  NAND2_X1 U14120 ( .A1(n11473), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11007) );
  INV_X1 U14121 ( .A(n11007), .ZN(n11004) );
  XNOR2_X1 U14122 ( .A(n11008), .B(n11004), .ZN(n20106) );
  NAND2_X1 U14123 ( .A1(n20106), .A2(n11477), .ZN(n11005) );
  INV_X1 U14124 ( .A(n17017), .ZN(n11006) );
  NAND2_X1 U14125 ( .A1(n11005), .A2(n10458), .ZN(n17016) );
  NAND3_X1 U14126 ( .A1(n11009), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n11473), 
        .ZN(n11010) );
  NAND3_X1 U14127 ( .A1(n11013), .A2(n11456), .A3(n11010), .ZN(n20089) );
  XNOR2_X1 U14128 ( .A(n11011), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14853) );
  INV_X1 U14129 ( .A(n14853), .ZN(n11012) );
  INV_X1 U14130 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17007) );
  NAND2_X1 U14131 ( .A1(n11473), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11014) );
  OR2_X1 U14132 ( .A1(n11015), .A2(n11014), .ZN(n11016) );
  NAND2_X1 U14133 ( .A1(n11027), .A2(n11016), .ZN(n20080) );
  INV_X1 U14134 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11376) );
  INV_X1 U14135 ( .A(n11437), .ZN(n11018) );
  NAND2_X1 U14136 ( .A1(n11017), .A2(n11376), .ZN(n14826) );
  NAND2_X1 U14137 ( .A1(n11473), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11019) );
  MUX2_X1 U14138 ( .A(n11473), .B(n11019), .S(n11027), .Z(n11020) );
  NAND2_X1 U14139 ( .A1(n11020), .A2(n11023), .ZN(n16533) );
  INV_X1 U14140 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17277) );
  NAND2_X1 U14141 ( .A1(n11021), .A2(n17277), .ZN(n11424) );
  INV_X1 U14142 ( .A(n11424), .ZN(n16988) );
  INV_X1 U14143 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11024) );
  INV_X1 U14144 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n16737) );
  NAND2_X1 U14145 ( .A1(n11024), .A2(n16737), .ZN(n11025) );
  AND2_X1 U14146 ( .A1(n11473), .A2(n11025), .ZN(n11026) );
  INV_X1 U14147 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U14148 ( .A1(n11029), .A2(n11028), .ZN(n11423) );
  INV_X1 U14149 ( .A(n11031), .ZN(n11035) );
  INV_X1 U14150 ( .A(n11172), .ZN(n11032) );
  NAND2_X1 U14151 ( .A1(n11033), .A2(n11032), .ZN(n11034) );
  NAND2_X1 U14152 ( .A1(n11035), .A2(n11034), .ZN(n11039) );
  INV_X1 U14153 ( .A(n11036), .ZN(n11037) );
  NAND3_X1 U14154 ( .A1(n11039), .A2(n11038), .A3(n11037), .ZN(n11044) );
  NOR2_X1 U14155 ( .A1(n11181), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11040) );
  AND2_X1 U14156 ( .A1(n11044), .A2(n11180), .ZN(n20952) );
  OR2_X1 U14157 ( .A1(n11045), .A2(n17495), .ZN(n20950) );
  NOR2_X1 U14158 ( .A1(n20950), .A2(n16694), .ZN(n11205) );
  NAND2_X1 U14159 ( .A1(n20952), .A2(n11205), .ZN(n11199) );
  INV_X1 U14160 ( .A(n11045), .ZN(n11182) );
  INV_X1 U14161 ( .A(n11046), .ZN(n11047) );
  XNOR2_X1 U14162 ( .A(n11172), .B(n11047), .ZN(n11167) );
  INV_X1 U14163 ( .A(n11048), .ZN(n11050) );
  NAND2_X1 U14164 ( .A1(n11050), .A2(n11049), .ZN(n11178) );
  NOR2_X1 U14165 ( .A1(n11170), .A2(n11178), .ZN(n11052) );
  NAND2_X1 U14166 ( .A1(n11167), .A2(n11052), .ZN(n11051) );
  AOI21_X1 U14167 ( .B1(n11168), .B2(n11052), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n11053) );
  INV_X1 U14168 ( .A(n11053), .ZN(n11057) );
  INV_X1 U14169 ( .A(n11054), .ZN(n14338) );
  NAND2_X1 U14170 ( .A1(n14338), .A2(n11181), .ZN(n14392) );
  INV_X1 U14171 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n14104) );
  OAI21_X1 U14172 ( .B1(n10619), .B2(n14392), .A(n14104), .ZN(n11056) );
  NAND2_X1 U14173 ( .A1(n11056), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20940) );
  OAI21_X1 U14174 ( .B1(n14388), .B2(n11057), .A(n20940), .ZN(n20951) );
  NAND3_X1 U14175 ( .A1(n11182), .A2(n9887), .A3(n20951), .ZN(n11058) );
  NAND2_X1 U14176 ( .A1(n11199), .A2(n11058), .ZN(n11059) );
  NAND3_X1 U14177 ( .A1(n11055), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n14802) );
  INV_X1 U14178 ( .A(n14802), .ZN(n14498) );
  INV_X1 U14179 ( .A(n11062), .ZN(n11061) );
  NOR3_X1 U14180 ( .A1(n11061), .A2(n13917), .A3(n11060), .ZN(n11065) );
  NOR2_X1 U14181 ( .A1(n13917), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11063) );
  XNOR2_X1 U14182 ( .A(n11063), .B(n11062), .ZN(n13333) );
  AND2_X1 U14183 ( .A1(n13333), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11064) );
  NOR2_X1 U14184 ( .A1(n11065), .A2(n11064), .ZN(n11068) );
  XNOR2_X1 U14185 ( .A(n10751), .B(n11068), .ZN(n14274) );
  INV_X1 U14186 ( .A(n14274), .ZN(n11067) );
  XNOR2_X1 U14187 ( .A(n11066), .B(n11222), .ZN(n14272) );
  NAND2_X1 U14188 ( .A1(n11067), .A2(n14272), .ZN(n17197) );
  OR2_X1 U14189 ( .A1(n11068), .A2(n10751), .ZN(n11069) );
  NAND2_X1 U14190 ( .A1(n17197), .A2(n11069), .ZN(n11070) );
  XNOR2_X1 U14191 ( .A(n11070), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17178) );
  NAND2_X1 U14192 ( .A1(n11070), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11071) );
  NAND2_X1 U14193 ( .A1(n11073), .A2(n10899), .ZN(n11074) );
  NAND2_X1 U14194 ( .A1(n11075), .A2(n11074), .ZN(n17158) );
  INV_X1 U14195 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17432) );
  INV_X1 U14196 ( .A(n9687), .ZN(n11079) );
  NAND2_X1 U14197 ( .A1(n11078), .A2(n9687), .ZN(n11083) );
  NAND2_X1 U14198 ( .A1(n11081), .A2(n9941), .ZN(n11082) );
  NAND2_X1 U14199 ( .A1(n17105), .A2(n17397), .ZN(n11086) );
  AND2_X1 U14200 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17073) );
  AND2_X1 U14201 ( .A1(n17073), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17301) );
  NAND2_X1 U14202 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17304) );
  NOR2_X1 U14203 ( .A1(n17304), .A2(n17308), .ZN(n11088) );
  NAND2_X1 U14204 ( .A1(n17301), .A2(n11088), .ZN(n14835) );
  INV_X1 U14205 ( .A(n14835), .ZN(n11089) );
  OAI21_X1 U14206 ( .B1(n16991), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n16981), .ZN(n11206) );
  INV_X1 U14207 ( .A(n13219), .ZN(n11090) );
  NOR2_X1 U14208 ( .A1(n11206), .A2(n17139), .ZN(n11164) );
  INV_X1 U14209 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20880) );
  NAND2_X1 U14210 ( .A1(n11120), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11094) );
  NAND2_X1 U14211 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11093) );
  OAI211_X1 U14212 ( .C1(n11542), .C2(n20880), .A(n11094), .B(n11093), .ZN(
        n11095) );
  AOI21_X1 U14213 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11095), .ZN(n11522) );
  INV_X1 U14214 ( .A(n11096), .ZN(n11098) );
  NAND2_X1 U14215 ( .A1(n11101), .A2(n11100), .ZN(n17162) );
  INV_X1 U14216 ( .A(n17162), .ZN(n11108) );
  NAND2_X1 U14217 ( .A1(n11555), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11104) );
  NAND2_X1 U14218 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11103) );
  OAI211_X1 U14219 ( .C1(n11102), .C2(n11105), .A(n11104), .B(n11103), .ZN(
        n11106) );
  AOI21_X1 U14220 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n11106), .ZN(n17161) );
  NAND2_X1 U14221 ( .A1(n11108), .A2(n11107), .ZN(n14609) );
  INV_X1 U14222 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n17148) );
  NAND2_X1 U14223 ( .A1(n11120), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11110) );
  NAND2_X1 U14224 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11109) );
  OAI211_X1 U14225 ( .C1(n11542), .C2(n17148), .A(n11110), .B(n11109), .ZN(
        n11111) );
  AOI21_X1 U14226 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11111), .ZN(n14610) );
  NOR2_X2 U14227 ( .A1(n14609), .A2(n14610), .ZN(n14611) );
  AOI22_X1 U14228 ( .A1(n11555), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11113) );
  NAND2_X1 U14229 ( .A1(n11120), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11112) );
  OAI211_X1 U14230 ( .C1(n11091), .C2(n17405), .A(n11113), .B(n11112), .ZN(
        n14260) );
  AOI22_X1 U14231 ( .A1(n11555), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11115) );
  NAND2_X1 U14232 ( .A1(n11120), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11114) );
  OAI211_X1 U14233 ( .C1(n11091), .C2(n17397), .A(n11115), .B(n11114), .ZN(
        n14254) );
  INV_X1 U14234 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n17115) );
  NAND2_X1 U14235 ( .A1(n11120), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11117) );
  NAND2_X1 U14236 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11116) );
  OAI211_X1 U14237 ( .C1(n11542), .C2(n17115), .A(n11117), .B(n11116), .ZN(
        n11118) );
  AOI21_X1 U14238 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n11118), .ZN(n14628) );
  INV_X1 U14239 ( .A(n14628), .ZN(n11119) );
  INV_X1 U14240 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20861) );
  NAND2_X1 U14241 ( .A1(n11120), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11122) );
  NAND2_X1 U14242 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11121) );
  OAI211_X1 U14243 ( .C1(n11542), .C2(n20861), .A(n11122), .B(n11121), .ZN(
        n11123) );
  AOI21_X1 U14244 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11123), .ZN(n14493) );
  AOI22_X1 U14245 ( .A1(n11555), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11125) );
  NAND2_X1 U14246 ( .A1(n11120), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11124) );
  OAI211_X1 U14247 ( .C1(n11091), .C2(n17361), .A(n11125), .B(n11124), .ZN(
        n14426) );
  INV_X1 U14248 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n20865) );
  NAND2_X1 U14249 ( .A1(n11120), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11127) );
  NAND2_X1 U14250 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11126) );
  OAI211_X1 U14251 ( .C1(n11542), .C2(n20865), .A(n11127), .B(n11126), .ZN(
        n11128) );
  AOI21_X1 U14252 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11128), .ZN(n14563) );
  INV_X1 U14253 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n20869) );
  NAND2_X1 U14254 ( .A1(n11120), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11132) );
  NAND2_X1 U14255 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11131) );
  OAI211_X1 U14256 ( .C1(n11542), .C2(n20869), .A(n11132), .B(n11131), .ZN(
        n11133) );
  AOI21_X1 U14257 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11133), .ZN(n14701) );
  INV_X1 U14258 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20867) );
  NAND2_X1 U14259 ( .A1(n11120), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11135) );
  NAND2_X1 U14260 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11134) );
  OAI211_X1 U14261 ( .C1(n11542), .C2(n20867), .A(n11135), .B(n11134), .ZN(
        n11136) );
  AOI21_X1 U14262 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11136), .ZN(n14589) );
  AOI22_X1 U14263 ( .A1(n11555), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11139) );
  NAND2_X1 U14264 ( .A1(n11120), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11138) );
  OAI211_X1 U14265 ( .C1(n11091), .C2(n17308), .A(n11139), .B(n11138), .ZN(
        n14642) );
  INV_X1 U14266 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20873) );
  NAND2_X1 U14267 ( .A1(n11120), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11141) );
  NAND2_X1 U14268 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11140) );
  OAI211_X1 U14269 ( .C1(n11542), .C2(n20873), .A(n11141), .B(n11140), .ZN(
        n11142) );
  AOI21_X1 U14270 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n11142), .ZN(n16756) );
  INV_X1 U14271 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20875) );
  NAND2_X1 U14272 ( .A1(n11120), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11145) );
  NAND2_X1 U14273 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11144) );
  OAI211_X1 U14274 ( .C1(n11542), .C2(n20875), .A(n11145), .B(n11144), .ZN(
        n11146) );
  AOI21_X1 U14275 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11146), .ZN(n14845) );
  AOI22_X1 U14276 ( .A1(n11555), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11148) );
  NAND2_X1 U14277 ( .A1(n11120), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11147) );
  OAI211_X1 U14278 ( .C1(n11091), .C2(n11376), .A(n11148), .B(n11147), .ZN(
        n14837) );
  AOI22_X1 U14279 ( .A1(n11555), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11150) );
  NAND2_X1 U14280 ( .A1(n11120), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11149) );
  OAI211_X1 U14281 ( .C1(n11091), .C2(n17277), .A(n11150), .B(n11149), .ZN(
        n16527) );
  OR2_X1 U14282 ( .A1(n16526), .A2(n11522), .ZN(n16500) );
  INV_X1 U14283 ( .A(n16500), .ZN(n11151) );
  AOI21_X1 U14284 ( .B1(n11522), .B2(n16526), .A(n11151), .ZN(n16733) );
  NOR2_X2 U14285 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20958) );
  NOR2_X1 U14286 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20911) );
  OR2_X1 U14287 ( .A1(n20958), .A2(n20911), .ZN(n20943) );
  NAND2_X1 U14288 ( .A1(n20943), .A2(n11573), .ZN(n11152) );
  AND2_X1 U14289 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20929) );
  NAND2_X1 U14290 ( .A1(n11578), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11586) );
  INV_X1 U14291 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11608) );
  INV_X1 U14292 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16520) );
  NAND2_X1 U14293 ( .A1(n11610), .A2(n16520), .ZN(n11158) );
  NAND2_X1 U14294 ( .A1(n11156), .A2(n11158), .ZN(n16513) );
  NAND2_X1 U14295 ( .A1(n11573), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12239) );
  INV_X1 U14296 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20910) );
  NAND2_X1 U14297 ( .A1(n20910), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11159) );
  NAND2_X1 U14298 ( .A1(n12239), .A2(n11159), .ZN(n13341) );
  NOR2_X1 U14299 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n11639) );
  NAND2_X1 U14300 ( .A1(n20911), .A2(n11639), .ZN(n20181) );
  INV_X1 U14301 ( .A(n20167), .ZN(n17149) );
  NOR2_X1 U14302 ( .A1(n17149), .A2(n20880), .ZN(n11409) );
  AOI21_X1 U14303 ( .B1(n17172), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n11409), .ZN(n11160) );
  OAI21_X1 U14304 ( .B1(n16513), .B2(n17175), .A(n11160), .ZN(n11161) );
  OAI21_X1 U14305 ( .B1(n11421), .B2(n17181), .A(n11165), .ZN(P2_U2995) );
  MUX2_X1 U14306 ( .A(n20968), .B(n10876), .S(n11166), .Z(n11177) );
  OAI21_X1 U14307 ( .B1(n16694), .B2(n11168), .A(n11167), .ZN(n11169) );
  OAI21_X1 U14308 ( .B1(n11170), .B2(n16694), .A(n11169), .ZN(n11171) );
  NAND2_X1 U14309 ( .A1(n11171), .A2(n17495), .ZN(n11175) );
  OAI21_X1 U14310 ( .B1(n11173), .B2(n11172), .A(n9887), .ZN(n11174) );
  NAND2_X1 U14311 ( .A1(n11175), .A2(n11174), .ZN(n11176) );
  NAND2_X1 U14312 ( .A1(n11177), .A2(n11176), .ZN(n11179) );
  MUX2_X1 U14313 ( .A(n13389), .B(n13223), .S(n14410), .Z(n11202) );
  NAND2_X1 U14314 ( .A1(READY12_REG_SCAN_IN), .A2(READY21_REG_SCAN_IN), .ZN(
        n20966) );
  NOR2_X1 U14315 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n20838) );
  AOI211_X1 U14316 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n20838), .ZN(n20965) );
  INV_X1 U14317 ( .A(n20965), .ZN(n20834) );
  INV_X1 U14318 ( .A(n20834), .ZN(n20967) );
  AND2_X1 U14319 ( .A1(n20966), .A2(n20967), .ZN(n13215) );
  AND2_X1 U14320 ( .A1(n11388), .A2(n13215), .ZN(n11183) );
  INV_X1 U14321 ( .A(n11185), .ZN(n11370) );
  NAND2_X1 U14322 ( .A1(n11187), .A2(n20298), .ZN(n11194) );
  INV_X2 U14323 ( .A(n13780), .ZN(n20316) );
  OAI21_X1 U14324 ( .B1(n11188), .B2(n20316), .A(n11651), .ZN(n11381) );
  NAND2_X1 U14325 ( .A1(n9921), .A2(n17495), .ZN(n11189) );
  NAND3_X1 U14326 ( .A1(n20968), .A2(n11189), .A3(n13780), .ZN(n11190) );
  AOI21_X1 U14327 ( .B1(n20298), .B2(n11190), .A(n11386), .ZN(n11192) );
  NAND3_X1 U14328 ( .A1(n11381), .A2(n11192), .A3(n11191), .ZN(n11193) );
  AOI21_X1 U14329 ( .B1(n11370), .B2(n11194), .A(n11193), .ZN(n11378) );
  OAI21_X1 U14330 ( .B1(n20965), .B2(n16694), .A(n14404), .ZN(n11196) );
  OAI21_X1 U14331 ( .B1(n20298), .B2(n16694), .A(n11196), .ZN(n11197) );
  INV_X1 U14332 ( .A(n14388), .ZN(n14347) );
  NAND3_X1 U14333 ( .A1(n11197), .A2(n14347), .A3(n20966), .ZN(n11198) );
  NAND3_X1 U14334 ( .A1(n11378), .A2(n11199), .A3(n11198), .ZN(n11200) );
  NOR2_X2 U14335 ( .A1(n11203), .A2(n14802), .ZN(n11415) );
  NOR2_X1 U14336 ( .A1(n20950), .A2(n13223), .ZN(n11204) );
  INV_X1 U14337 ( .A(n11415), .ZN(n11402) );
  INV_X1 U14338 ( .A(n11205), .ZN(n20953) );
  NOR2_X1 U14339 ( .A1(n11206), .A2(n17415), .ZN(n11419) );
  AND2_X2 U14340 ( .A1(n11220), .A2(n17491), .ZN(n11225) );
  NAND2_X1 U14341 ( .A1(n12494), .A2(n11225), .ZN(n13918) );
  MUX2_X1 U14342 ( .A(n11208), .B(n20947), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n13919) );
  NAND4_X2 U14343 ( .A1(n11208), .A2(n11207), .A3(n9989), .A4(n17491), .ZN(
        n11361) );
  INV_X1 U14344 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n20071) );
  AOI21_X1 U14345 ( .B1(n11220), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11210) );
  NAND2_X1 U14346 ( .A1(n20316), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11209) );
  NAND2_X1 U14347 ( .A1(n10563), .A2(n13921), .ZN(n13924) );
  INV_X1 U14348 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20847) );
  NAND2_X1 U14349 ( .A1(n11225), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11212) );
  AND2_X2 U14350 ( .A1(n20316), .A2(n17491), .ZN(n11224) );
  NAND2_X1 U14351 ( .A1(n11224), .A2(P2_EAX_REG_1__SCAN_IN), .ZN(n11211) );
  OAI211_X1 U14352 ( .C1(n11361), .C2(n20847), .A(n11212), .B(n11211), .ZN(
        n11216) );
  XNOR2_X1 U14353 ( .A(n13924), .B(n11216), .ZN(n13909) );
  INV_X1 U14354 ( .A(n11213), .ZN(n11214) );
  AOI22_X1 U14355 ( .A1(n11214), .A2(n9989), .B1(n13780), .B2(n10726), .ZN(
        n11215) );
  MUX2_X1 U14356 ( .A(n20938), .B(n11215), .S(n17491), .Z(n13908) );
  INV_X1 U14357 ( .A(n11216), .ZN(n11217) );
  NAND2_X1 U14358 ( .A1(n13924), .A2(n11217), .ZN(n11218) );
  NAND2_X1 U14359 ( .A1(n13911), .A2(n11218), .ZN(n11230) );
  OR2_X1 U14360 ( .A1(n13916), .A2(n11222), .ZN(n11223) );
  OAI211_X1 U14361 ( .C1(n17491), .C2(n20927), .A(n11223), .B(n13918), .ZN(
        n11228) );
  XNOR2_X1 U14362 ( .A(n11230), .B(n11228), .ZN(n13900) );
  NAND2_X1 U14363 ( .A1(n11512), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11227) );
  AOI22_X1 U14364 ( .A1(n11224), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11225), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11226) );
  AND2_X1 U14365 ( .A1(n11227), .A2(n11226), .ZN(n13901) );
  INV_X1 U14366 ( .A(n11228), .ZN(n11229) );
  NAND2_X1 U14367 ( .A1(n11230), .A2(n11229), .ZN(n11231) );
  AOI22_X1 U14368 ( .A1(n11512), .A2(P2_REIP_REG_3__SCAN_IN), .B1(n11224), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n11236) );
  INV_X1 U14369 ( .A(n13916), .ZN(n11234) );
  OAI22_X1 U14370 ( .A1(n11232), .A2(n11398), .B1(n20920), .B2(n17491), .ZN(
        n11233) );
  AOI21_X1 U14371 ( .B1(n11234), .B2(n10877), .A(n11233), .ZN(n11235) );
  NAND2_X1 U14372 ( .A1(n11512), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11240) );
  OR2_X1 U14373 ( .A1(n13916), .A2(n10899), .ZN(n11239) );
  AOI22_X1 U14374 ( .A1(n11224), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11225), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11238) );
  NAND2_X1 U14375 ( .A1(n11512), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11246) );
  OR2_X1 U14376 ( .A1(n13916), .A2(n11243), .ZN(n11245) );
  AOI22_X1 U14377 ( .A1(n11224), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11225), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11244) );
  INV_X1 U14378 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20856) );
  NAND2_X1 U14379 ( .A1(n11225), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11249) );
  NAND2_X1 U14380 ( .A1(n11224), .A2(P2_EAX_REG_6__SCAN_IN), .ZN(n11248) );
  OAI211_X1 U14381 ( .C1(n11361), .C2(n20856), .A(n11249), .B(n11248), .ZN(
        n13980) );
  INV_X1 U14382 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20858) );
  NAND2_X1 U14383 ( .A1(n11225), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11251) );
  NAND2_X1 U14384 ( .A1(n11224), .A2(P2_EAX_REG_7__SCAN_IN), .ZN(n11250) );
  OAI211_X1 U14385 ( .C1(n11361), .C2(n20858), .A(n11251), .B(n11250), .ZN(
        n13977) );
  NAND2_X1 U14386 ( .A1(n11512), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11264) );
  AOI22_X1 U14387 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11255) );
  AOI22_X1 U14388 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14389 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11253) );
  AOI22_X1 U14390 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11252) );
  NAND4_X1 U14391 ( .A1(n11255), .A2(n11254), .A3(n11253), .A4(n11252), .ZN(
        n11261) );
  AOI22_X1 U14392 ( .A1(n10921), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11259) );
  AOI22_X1 U14393 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11258) );
  AOI22_X1 U14394 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11257) );
  AOI22_X1 U14395 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11256) );
  NAND4_X1 U14396 ( .A1(n11259), .A2(n11258), .A3(n11257), .A4(n11256), .ZN(
        n11260) );
  INV_X1 U14397 ( .A(n12249), .ZN(n14632) );
  OR2_X1 U14398 ( .A1(n13916), .A2(n14632), .ZN(n11263) );
  AOI22_X1 U14399 ( .A1(n11224), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11225), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11262) );
  NAND2_X1 U14400 ( .A1(n11512), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11279) );
  AOI22_X1 U14401 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11270) );
  AOI22_X1 U14402 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U14403 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11268) );
  AOI22_X1 U14404 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10921), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11267) );
  NAND4_X1 U14405 ( .A1(n11270), .A2(n11269), .A3(n11268), .A4(n11267), .ZN(
        n11276) );
  AOI22_X1 U14406 ( .A1(n10849), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11274) );
  AOI22_X1 U14407 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11273) );
  AOI22_X1 U14408 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11272) );
  AOI22_X1 U14409 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11271) );
  NAND4_X1 U14410 ( .A1(n11274), .A2(n11273), .A3(n11272), .A4(n11271), .ZN(
        n11275) );
  NOR2_X1 U14411 ( .A1(n11276), .A2(n11275), .ZN(n12247) );
  OR2_X1 U14412 ( .A1(n13916), .A2(n12247), .ZN(n11278) );
  AOI22_X1 U14413 ( .A1(n11224), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11225), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11277) );
  INV_X1 U14414 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20863) );
  AOI22_X1 U14415 ( .A1(n11224), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11291) );
  AOI22_X1 U14416 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11283) );
  AOI22_X1 U14417 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11282) );
  AOI22_X1 U14418 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11281) );
  AOI22_X1 U14419 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11280) );
  NAND4_X1 U14420 ( .A1(n11283), .A2(n11282), .A3(n11281), .A4(n11280), .ZN(
        n11289) );
  AOI22_X1 U14421 ( .A1(n10921), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11287) );
  AOI22_X1 U14422 ( .A1(n10624), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14423 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12309), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11285) );
  AOI22_X1 U14424 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11284) );
  NAND4_X1 U14425 ( .A1(n11287), .A2(n11286), .A3(n11285), .A4(n11284), .ZN(
        n11288) );
  INV_X1 U14426 ( .A(n14422), .ZN(n14420) );
  OR2_X1 U14427 ( .A1(n13916), .A2(n14420), .ZN(n11290) );
  OAI211_X1 U14428 ( .C1(n11361), .C2(n20863), .A(n11291), .B(n11290), .ZN(
        n13876) );
  NAND2_X1 U14429 ( .A1(n11512), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11305) );
  AOI22_X1 U14430 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11295) );
  AOI22_X1 U14431 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11294) );
  AOI22_X1 U14432 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11293) );
  AOI22_X1 U14433 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10921), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11292) );
  NAND4_X1 U14434 ( .A1(n11295), .A2(n11294), .A3(n11293), .A4(n11292), .ZN(
        n11301) );
  AOI22_X1 U14435 ( .A1(n10849), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11299) );
  AOI22_X1 U14436 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11298) );
  AOI22_X1 U14437 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11297) );
  AOI22_X1 U14438 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11296) );
  NAND4_X1 U14439 ( .A1(n11299), .A2(n11298), .A3(n11297), .A4(n11296), .ZN(
        n11300) );
  INV_X1 U14440 ( .A(n14564), .ZN(n11302) );
  OR2_X1 U14441 ( .A1(n13916), .A2(n11302), .ZN(n11304) );
  AOI22_X1 U14442 ( .A1(n11224), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11303) );
  NAND2_X1 U14443 ( .A1(n11512), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11318) );
  AOI22_X1 U14444 ( .A1(n10803), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11309) );
  AOI22_X1 U14445 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11308) );
  AOI22_X1 U14446 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11307) );
  AOI22_X1 U14447 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10804), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11306) );
  NAND4_X1 U14448 ( .A1(n11309), .A2(n11308), .A3(n11307), .A4(n11306), .ZN(
        n11315) );
  AOI22_X1 U14449 ( .A1(n10921), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11313) );
  AOI22_X1 U14450 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11312) );
  AOI22_X1 U14451 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12356), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11311) );
  AOI22_X1 U14452 ( .A1(n10625), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11310) );
  NAND4_X1 U14453 ( .A1(n11313), .A2(n11312), .A3(n11311), .A4(n11310), .ZN(
        n11314) );
  INV_X1 U14454 ( .A(n14595), .ZN(n14592) );
  OR2_X1 U14455 ( .A1(n13916), .A2(n14592), .ZN(n11317) );
  AOI22_X1 U14456 ( .A1(n11224), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11316) );
  AOI22_X1 U14457 ( .A1(n11224), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11330) );
  AOI22_X1 U14458 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11322) );
  AOI22_X1 U14459 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U14460 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11320) );
  AOI22_X1 U14461 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10921), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11319) );
  NAND4_X1 U14462 ( .A1(n11322), .A2(n11321), .A3(n11320), .A4(n11319), .ZN(
        n11328) );
  AOI22_X1 U14463 ( .A1(n10849), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14464 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14465 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U14466 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11323) );
  NAND4_X1 U14467 ( .A1(n11326), .A2(n11325), .A3(n11324), .A4(n11323), .ZN(
        n11327) );
  NOR2_X1 U14468 ( .A1(n11328), .A2(n11327), .ZN(n12252) );
  OR2_X1 U14469 ( .A1(n13916), .A2(n12252), .ZN(n11329) );
  OAI211_X1 U14470 ( .C1(n11361), .C2(n20869), .A(n11330), .B(n11329), .ZN(
        n14432) );
  NAND2_X1 U14471 ( .A1(n14433), .A2(n14432), .ZN(n14431) );
  NAND2_X1 U14472 ( .A1(n11512), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14473 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11334) );
  AOI22_X1 U14474 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14475 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14476 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11331) );
  NAND4_X1 U14477 ( .A1(n11334), .A2(n11333), .A3(n11332), .A4(n11331), .ZN(
        n11340) );
  AOI22_X1 U14478 ( .A1(n10921), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11338) );
  AOI22_X1 U14479 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U14480 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U14481 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11335) );
  NAND4_X1 U14482 ( .A1(n11338), .A2(n11337), .A3(n11336), .A4(n11335), .ZN(
        n11339) );
  NOR2_X1 U14483 ( .A1(n11340), .A2(n11339), .ZN(n14643) );
  OR2_X1 U14484 ( .A1(n13916), .A2(n14643), .ZN(n11342) );
  AOI22_X1 U14485 ( .A1(n11224), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11341) );
  NAND2_X1 U14486 ( .A1(n11512), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U14487 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U14488 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10803), .B1(
        n10802), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U14489 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11345) );
  AOI22_X1 U14490 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n10921), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11344) );
  NAND4_X1 U14491 ( .A1(n11347), .A2(n11346), .A3(n11345), .A4(n11344), .ZN(
        n11353) );
  AOI22_X1 U14492 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10849), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11351) );
  AOI22_X1 U14493 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n12309), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U14494 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12355), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11349) );
  AOI22_X1 U14495 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10797), .B1(
        n12356), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11348) );
  NAND4_X1 U14496 ( .A1(n11351), .A2(n11350), .A3(n11349), .A4(n11348), .ZN(
        n11352) );
  NOR2_X1 U14497 ( .A1(n11353), .A2(n11352), .ZN(n12253) );
  OR2_X1 U14498 ( .A1(n13916), .A2(n12253), .ZN(n11355) );
  AOI22_X1 U14499 ( .A1(n11224), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11354) );
  NAND2_X1 U14500 ( .A1(n11512), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14501 ( .A1(n11224), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11357) );
  INV_X1 U14502 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20877) );
  NAND2_X1 U14503 ( .A1(n11225), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11360) );
  NAND2_X1 U14504 ( .A1(n11224), .A2(P2_EAX_REG_17__SCAN_IN), .ZN(n11359) );
  OAI211_X1 U14505 ( .C1(n11361), .C2(n20877), .A(n11360), .B(n11359), .ZN(
        n14840) );
  INV_X1 U14506 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n16992) );
  NAND2_X1 U14507 ( .A1(n11225), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11363) );
  NAND2_X1 U14508 ( .A1(n11224), .A2(P2_EAX_REG_18__SCAN_IN), .ZN(n11362) );
  OAI211_X1 U14509 ( .C1(n11361), .C2(n16992), .A(n11363), .B(n11362), .ZN(
        n16535) );
  NAND2_X1 U14510 ( .A1(n11512), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11365) );
  AOI22_X1 U14511 ( .A1(n11224), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11364) );
  NAND2_X1 U14512 ( .A1(n16534), .A2(n11368), .ZN(n11369) );
  NAND2_X1 U14513 ( .A1(n11498), .A2(n11369), .ZN(n16855) );
  NAND2_X1 U14514 ( .A1(n11370), .A2(n11643), .ZN(n14389) );
  INV_X1 U14515 ( .A(n11372), .ZN(n11373) );
  NOR2_X1 U14516 ( .A1(n15442), .A2(n11373), .ZN(n11374) );
  NOR2_X1 U14517 ( .A1(n11371), .A2(n14356), .ZN(n13778) );
  AOI21_X1 U14518 ( .B1(n16694), .B2(n14389), .A(n13778), .ZN(n11375) );
  NOR2_X2 U14519 ( .A1(n11402), .A2(n11375), .ZN(n17461) );
  NOR3_X1 U14520 ( .A1(n17007), .A2(n10458), .A3(n11376), .ZN(n17278) );
  NAND2_X1 U14521 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17278), .ZN(
        n11377) );
  NOR2_X1 U14522 ( .A1(n14835), .A2(n11377), .ZN(n11487) );
  INV_X1 U14523 ( .A(n11378), .ZN(n14343) );
  NAND2_X1 U14524 ( .A1(n13223), .A2(n11389), .ZN(n11379) );
  NAND2_X1 U14525 ( .A1(n11380), .A2(n16694), .ZN(n14355) );
  NAND2_X1 U14526 ( .A1(n14355), .A2(n11381), .ZN(n11383) );
  NAND2_X1 U14527 ( .A1(n11383), .A2(n11382), .ZN(n11395) );
  NAND2_X1 U14528 ( .A1(n9937), .A2(n11384), .ZN(n11385) );
  NAND2_X1 U14529 ( .A1(n9692), .A2(n11385), .ZN(n11387) );
  NAND2_X1 U14530 ( .A1(n11387), .A2(n11386), .ZN(n11392) );
  AOI22_X1 U14531 ( .A1(n15442), .A2(n11389), .B1(n13389), .B2(n11388), .ZN(
        n11391) );
  NAND2_X1 U14532 ( .A1(n11396), .A2(n11390), .ZN(n12193) );
  AND3_X1 U14533 ( .A1(n11392), .A2(n11391), .A3(n12193), .ZN(n11394) );
  NAND3_X1 U14534 ( .A1(n11395), .A2(n11394), .A3(n11393), .ZN(n14363) );
  OR2_X1 U14535 ( .A1(n14363), .A2(n11396), .ZN(n11397) );
  INV_X1 U14536 ( .A(n11399), .ZN(n14830) );
  NAND2_X1 U14537 ( .A1(n13990), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14276) );
  NAND2_X1 U14538 ( .A1(n14830), .A2(n14276), .ZN(n14280) );
  INV_X1 U14539 ( .A(n14280), .ZN(n11401) );
  NOR2_X1 U14540 ( .A1(n13990), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14281) );
  INV_X1 U14541 ( .A(n14281), .ZN(n11400) );
  NOR2_X1 U14542 ( .A1(n14828), .A2(n11400), .ZN(n14270) );
  NOR2_X1 U14543 ( .A1(n11401), .A2(n14270), .ZN(n11403) );
  NAND2_X1 U14544 ( .A1(n11402), .A2(n20181), .ZN(n17451) );
  NAND2_X1 U14545 ( .A1(n11403), .A2(n17451), .ZN(n17439) );
  NOR2_X1 U14546 ( .A1(n17423), .A2(n17432), .ZN(n17417) );
  INV_X1 U14547 ( .A(n17417), .ZN(n11407) );
  NAND2_X1 U14548 ( .A1(n10181), .A2(n11407), .ZN(n11404) );
  AND2_X1 U14549 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11405) );
  AND2_X1 U14550 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n11405), .ZN(
        n11406) );
  OAI21_X1 U14551 ( .B1(n11487), .B2(n17452), .A(n17303), .ZN(n17281) );
  INV_X1 U14552 ( .A(n17370), .ZN(n17300) );
  NAND2_X1 U14553 ( .A1(n11487), .A2(n17300), .ZN(n17265) );
  NOR2_X1 U14554 ( .A1(n17265), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11408) );
  AOI211_X1 U14555 ( .C1(n17281), .C2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11409), .B(n11408), .ZN(n11410) );
  OAI21_X1 U14556 ( .B1(n16855), .B2(n17444), .A(n11410), .ZN(n11411) );
  INV_X1 U14557 ( .A(n11411), .ZN(n11417) );
  NAND2_X1 U14558 ( .A1(n11412), .A2(n13223), .ZN(n11413) );
  NAND2_X1 U14559 ( .A1(n11413), .A2(n14333), .ZN(n11414) );
  NAND2_X1 U14560 ( .A1(n16733), .A2(n17456), .ZN(n11416) );
  OAI21_X1 U14561 ( .B1(n11421), .B2(n17458), .A(n11420), .ZN(P2_U3027) );
  NAND2_X1 U14562 ( .A1(n11424), .A2(n11423), .ZN(n16973) );
  NAND2_X1 U14563 ( .A1(n11473), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11425) );
  XNOR2_X1 U14564 ( .A(n11428), .B(n11425), .ZN(n16503) );
  NAND2_X1 U14565 ( .A1(n16503), .A2(n11477), .ZN(n11441) );
  INV_X1 U14566 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16980) );
  AND2_X1 U14567 ( .A1(n11441), .A2(n16980), .ZN(n16976) );
  AND4_X1 U14568 ( .A1(n17016), .A2(n11426), .A3(n17027), .A4(n17039), .ZN(
        n11427) );
  AND3_X1 U14569 ( .A1(n14826), .A2(n14853), .A3(n11427), .ZN(n11432) );
  INV_X1 U14570 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n16726) );
  NAND2_X1 U14571 ( .A1(n11473), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11429) );
  NOR2_X1 U14572 ( .A1(n11430), .A2(n11429), .ZN(n11431) );
  OR2_X1 U14573 ( .A1(n11444), .A2(n11431), .ZN(n16493) );
  INV_X1 U14574 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14862) );
  NAND2_X1 U14575 ( .A1(n11439), .A2(n14862), .ZN(n14858) );
  NOR2_X1 U14576 ( .A1(n17038), .A2(n11433), .ZN(n11434) );
  NAND4_X1 U14577 ( .A1(n11435), .A2(n11434), .A3(n17017), .A4(n17026), .ZN(
        n11436) );
  INV_X1 U14578 ( .A(n11439), .ZN(n11440) );
  NAND2_X1 U14579 ( .A1(n11440), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14859) );
  INV_X1 U14580 ( .A(n11441), .ZN(n11442) );
  NAND2_X1 U14581 ( .A1(n11473), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11443) );
  INV_X1 U14582 ( .A(n11443), .ZN(n11446) );
  AOI21_X1 U14583 ( .B1(n11446), .B2(n11445), .A(n11449), .ZN(n17822) );
  AOI21_X1 U14584 ( .B1(n17822), .B2(n11477), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16967) );
  INV_X2 U14585 ( .A(n11447), .ZN(n11449) );
  AND2_X1 U14586 ( .A1(n11473), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11450) );
  NAND2_X1 U14587 ( .A1(n11447), .A2(n11450), .ZN(n11451) );
  NAND2_X1 U14588 ( .A1(n16461), .A2(n11451), .ZN(n16473) );
  OR2_X1 U14589 ( .A1(n16473), .A2(n11482), .ZN(n11452) );
  XNOR2_X1 U14590 ( .A(n11452), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16958) );
  INV_X1 U14591 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11453) );
  NOR3_X1 U14592 ( .A1(n16473), .A2(n11482), .A3(n11453), .ZN(n16931) );
  NAND2_X1 U14593 ( .A1(n11456), .A2(n11477), .ZN(n16945) );
  INV_X1 U14594 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16949) );
  NOR2_X1 U14595 ( .A1(n16945), .A2(n16949), .ZN(n16933) );
  NOR2_X1 U14596 ( .A1(n16931), .A2(n16933), .ZN(n11454) );
  NAND2_X1 U14597 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11455) );
  INV_X1 U14598 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n16437) );
  INV_X1 U14599 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n16699) );
  NAND2_X1 U14600 ( .A1(n11473), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11459) );
  AND2_X1 U14601 ( .A1(n11473), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11457) );
  INV_X1 U14602 ( .A(n11459), .ZN(n11460) );
  NAND2_X1 U14603 ( .A1(n11461), .A2(n11460), .ZN(n11462) );
  AND2_X1 U14604 ( .A1(n11463), .A2(n11462), .ZN(n16409) );
  NAND2_X1 U14605 ( .A1(n16409), .A2(n11477), .ZN(n14885) );
  INV_X1 U14606 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14887) );
  INV_X1 U14607 ( .A(n11481), .ZN(n11466) );
  OAI211_X1 U14608 ( .C1(n9745), .C2(P2_EBX_REG_25__SCAN_IN), .A(n11473), .B(
        P2_EBX_REG_26__SCAN_IN), .ZN(n11465) );
  AOI21_X1 U14609 ( .B1(n16429), .B2(n11477), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14788) );
  AOI21_X1 U14610 ( .B1(n14885), .B2(n14887), .A(n14788), .ZN(n11467) );
  OAI21_X1 U14611 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n14889), .ZN(n11470) );
  INV_X1 U14612 ( .A(n16429), .ZN(n11469) );
  NAND2_X1 U14613 ( .A1(n11477), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11468) );
  INV_X1 U14614 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17218) );
  OR2_X1 U14615 ( .A1(n16945), .A2(n17218), .ZN(n16937) );
  NAND2_X1 U14616 ( .A1(n11473), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11471) );
  XNOR2_X1 U14617 ( .A(n11472), .B(n11471), .ZN(n11476) );
  OAI21_X1 U14618 ( .B1(n11476), .B2(n11482), .A(n9968), .ZN(n14899) );
  NAND2_X1 U14619 ( .A1(n11473), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11474) );
  XNOR2_X1 U14620 ( .A(n11480), .B(n11474), .ZN(n11475) );
  AOI21_X1 U14621 ( .B1(n11475), .B2(n11477), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12178) );
  INV_X1 U14622 ( .A(n11475), .ZN(n11664) );
  INV_X1 U14623 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11564) );
  INV_X1 U14624 ( .A(n11476), .ZN(n12504) );
  NAND3_X1 U14625 ( .A1(n12504), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11477), .ZN(n14900) );
  AND2_X1 U14626 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11486) );
  AND2_X1 U14627 ( .A1(n11487), .A2(n11486), .ZN(n14875) );
  AND2_X1 U14628 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17202) );
  NAND2_X1 U14629 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14902) );
  NOR2_X1 U14630 ( .A1(n14902), .A2(n11564), .ZN(n11488) );
  NAND2_X1 U14631 ( .A1(n15426), .A2(n17454), .ZN(n11569) );
  NAND2_X1 U14632 ( .A1(n11512), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11490) );
  AOI22_X1 U14633 ( .A1(n11224), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11489) );
  AND2_X1 U14634 ( .A1(n11490), .A2(n11489), .ZN(n11650) );
  INV_X1 U14635 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20896) );
  NAND2_X1 U14636 ( .A1(n11225), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11492) );
  NAND2_X1 U14637 ( .A1(n11224), .A2(P2_EAX_REG_29__SCAN_IN), .ZN(n11491) );
  OAI211_X1 U14638 ( .C1(n11361), .C2(n20896), .A(n11492), .B(n11491), .ZN(
        n12187) );
  INV_X1 U14639 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n14894) );
  NAND2_X1 U14640 ( .A1(n11225), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11494) );
  NAND2_X1 U14641 ( .A1(n11224), .A2(P2_EAX_REG_28__SCAN_IN), .ZN(n11493) );
  OAI211_X1 U14642 ( .C1(n11361), .C2(n14894), .A(n11494), .B(n11493), .ZN(
        n14913) );
  AND2_X1 U14643 ( .A1(n12187), .A2(n14913), .ZN(n11647) );
  INV_X1 U14644 ( .A(n11647), .ZN(n11495) );
  NOR2_X1 U14645 ( .A1(n11650), .A2(n11495), .ZN(n11515) );
  NAND2_X1 U14646 ( .A1(n11512), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11497) );
  AOI22_X1 U14647 ( .A1(n11224), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11496) );
  INV_X1 U14648 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20883) );
  NAND2_X1 U14649 ( .A1(n11225), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11500) );
  NAND2_X1 U14650 ( .A1(n11224), .A2(P2_EAX_REG_21__SCAN_IN), .ZN(n11499) );
  OAI211_X1 U14651 ( .C1(n11361), .C2(n20883), .A(n11500), .B(n11499), .ZN(
        n14872) );
  NAND2_X1 U14652 ( .A1(n11512), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11502) );
  AOI22_X1 U14653 ( .A1(n11224), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11501) );
  AND2_X1 U14654 ( .A1(n11502), .A2(n11501), .ZN(n16823) );
  NAND2_X1 U14655 ( .A1(n11512), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14656 ( .A1(n11224), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11503) );
  AND2_X1 U14657 ( .A1(n11504), .A2(n11503), .ZN(n16471) );
  INV_X1 U14658 ( .A(n16471), .ZN(n11505) );
  NAND2_X1 U14659 ( .A1(n11512), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14660 ( .A1(n11224), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11506) );
  NOR2_X2 U14661 ( .A1(n16456), .A2(n16457), .ZN(n16447) );
  INV_X1 U14662 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20889) );
  NAND2_X1 U14663 ( .A1(n11225), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11509) );
  NAND2_X1 U14664 ( .A1(n11224), .A2(P2_EAX_REG_25__SCAN_IN), .ZN(n11508) );
  OAI211_X1 U14665 ( .C1(n11361), .C2(n20889), .A(n11509), .B(n11508), .ZN(
        n16448) );
  NAND2_X1 U14666 ( .A1(n11512), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14667 ( .A1(n11224), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11510) );
  AND2_X1 U14668 ( .A1(n11511), .A2(n11510), .ZN(n16424) );
  NAND2_X1 U14669 ( .A1(n11512), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U14670 ( .A1(n11224), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11225), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11513) );
  INV_X1 U14671 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n11561) );
  NAND2_X1 U14672 ( .A1(n11225), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11517) );
  NAND2_X1 U14673 ( .A1(n11224), .A2(P2_EAX_REG_31__SCAN_IN), .ZN(n11516) );
  OAI211_X1 U14674 ( .C1(n11361), .C2(n11561), .A(n11517), .B(n11516), .ZN(
        n11518) );
  NAND2_X1 U14675 ( .A1(n16764), .A2(n17461), .ZN(n11568) );
  INV_X1 U14676 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n16982) );
  NAND2_X1 U14677 ( .A1(n11120), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11520) );
  NAND2_X1 U14678 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11519) );
  OAI211_X1 U14679 ( .C1(n11542), .C2(n16982), .A(n11520), .B(n11519), .ZN(
        n11521) );
  AOI21_X1 U14680 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11521), .ZN(n16499) );
  AOI22_X1 U14681 ( .A1(n11555), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11525) );
  NAND2_X1 U14682 ( .A1(n11120), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11524) );
  OAI211_X1 U14683 ( .C1(n11091), .C2(n14862), .A(n11525), .B(n11524), .ZN(
        n14865) );
  INV_X1 U14684 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n16968) );
  NAND2_X1 U14685 ( .A1(n11120), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11527) );
  NAND2_X1 U14686 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11526) );
  OAI211_X1 U14687 ( .C1(n11542), .C2(n16968), .A(n11527), .B(n11526), .ZN(
        n11528) );
  AOI21_X1 U14688 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n11528), .ZN(n16720) );
  INV_X1 U14689 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n16950) );
  NAND2_X1 U14690 ( .A1(n11120), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11532) );
  NAND2_X1 U14691 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11531) );
  OAI211_X1 U14692 ( .C1(n11542), .C2(n16950), .A(n11532), .B(n11531), .ZN(
        n11533) );
  AOI21_X1 U14693 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11533), .ZN(n16453) );
  INV_X1 U14694 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20886) );
  NAND2_X1 U14695 ( .A1(n11120), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11535) );
  NAND2_X1 U14696 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11534) );
  OAI211_X1 U14697 ( .C1(n11542), .C2(n20886), .A(n11535), .B(n11534), .ZN(
        n11536) );
  AOI21_X1 U14698 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11536), .ZN(n16485) );
  NOR2_X2 U14699 ( .A1(n16451), .A2(n11537), .ZN(n16454) );
  AOI22_X1 U14700 ( .A1(n11555), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11539) );
  NAND2_X1 U14701 ( .A1(n11120), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11538) );
  OAI211_X1 U14702 ( .C1(n11091), .C2(n17218), .A(n11539), .B(n11538), .ZN(
        n16434) );
  NAND2_X1 U14703 ( .A1(n16454), .A2(n16434), .ZN(n16436) );
  INV_X1 U14704 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20891) );
  NAND2_X1 U14705 ( .A1(n11120), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11541) );
  NAND2_X1 U14706 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11540) );
  OAI211_X1 U14707 ( .C1(n11542), .C2(n20891), .A(n11541), .B(n11540), .ZN(
        n11543) );
  AOI21_X1 U14708 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11543), .ZN(n16420) );
  INV_X1 U14709 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U14710 ( .A1(n11555), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11544) );
  OAI21_X1 U14711 ( .B1(n11102), .B2(n11545), .A(n11544), .ZN(n11546) );
  AOI21_X1 U14712 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11546), .ZN(n14794) );
  INV_X1 U14713 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U14714 ( .A1(n11555), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11548) );
  NAND2_X1 U14715 ( .A1(n11120), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11547) );
  OAI211_X1 U14716 ( .C1(n11091), .C2(n11549), .A(n11548), .B(n11547), .ZN(
        n14893) );
  INV_X1 U14717 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U14718 ( .A1(n11555), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11550) );
  OAI21_X1 U14719 ( .B1(n11102), .B2(n11551), .A(n11550), .ZN(n11552) );
  AOI21_X1 U14720 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11552), .ZN(n12506) );
  AOI22_X1 U14721 ( .A1(n11555), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11554) );
  NAND2_X1 U14722 ( .A1(n11120), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11553) );
  OAI211_X1 U14723 ( .C1(n11091), .C2(n11564), .A(n11554), .B(n11553), .ZN(
        n11642) );
  NAND2_X1 U14724 ( .A1(n11640), .A2(n11642), .ZN(n11641) );
  INV_X1 U14725 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14726 ( .A1(n11555), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11556) );
  OAI21_X1 U14727 ( .B1(n11102), .B2(n11657), .A(n11556), .ZN(n11557) );
  AOI21_X1 U14728 ( .B1(n11558), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n11557), .ZN(n11559) );
  NAND2_X1 U14729 ( .A1(n17431), .A2(n17452), .ZN(n17220) );
  NAND2_X1 U14730 ( .A1(n14875), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11562) );
  OAI21_X1 U14731 ( .B1(n17378), .B2(n11562), .A(n17220), .ZN(n17241) );
  NAND2_X1 U14732 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17242) );
  AOI21_X1 U14733 ( .B1(n17220), .B2(n17242), .A(n16949), .ZN(n11560) );
  NAND2_X1 U14734 ( .A1(n17241), .A2(n11560), .ZN(n17230) );
  INV_X1 U14735 ( .A(n17202), .ZN(n11563) );
  INV_X1 U14736 ( .A(n17220), .ZN(n17362) );
  NOR2_X1 U14737 ( .A1(n17149), .A2(n11561), .ZN(n15421) );
  NAND2_X1 U14738 ( .A1(n17231), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17216) );
  INV_X1 U14739 ( .A(n11566), .ZN(n11567) );
  OAI21_X1 U14740 ( .B1(n15428), .B2(n17458), .A(n11570), .ZN(P2_U3015) );
  NAND2_X1 U14741 ( .A1(n11611), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11614) );
  INV_X1 U14742 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17813) );
  INV_X1 U14743 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16475) );
  INV_X1 U14744 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11624) );
  INV_X1 U14745 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16423) );
  INV_X1 U14746 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16412) );
  NAND2_X1 U14747 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11574) );
  MUX2_X1 U14748 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n16640) );
  INV_X1 U14749 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13336) );
  MUX2_X1 U14750 ( .A(n13336), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n14804) );
  NOR2_X1 U14751 ( .A1(n16640), .A2(n14804), .ZN(n16614) );
  OAI21_X1 U14752 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n9752), .ZN(n17184) );
  AND2_X1 U14753 ( .A1(n16614), .A2(n17184), .ZN(n16607) );
  INV_X1 U14754 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11576) );
  NAND2_X1 U14755 ( .A1(n9752), .A2(n11576), .ZN(n11577) );
  NAND2_X1 U14756 ( .A1(n11580), .A2(n11577), .ZN(n17174) );
  NAND2_X1 U14757 ( .A1(n16607), .A2(n17174), .ZN(n20192) );
  INV_X1 U14758 ( .A(n11578), .ZN(n11583) );
  NAND2_X1 U14759 ( .A1(n11580), .A2(n11579), .ZN(n11581) );
  AND2_X1 U14760 ( .A1(n11583), .A2(n11581), .ZN(n20195) );
  OR2_X1 U14761 ( .A1(n20192), .A2(n20195), .ZN(n20196) );
  INV_X1 U14762 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11582) );
  NAND2_X1 U14763 ( .A1(n11583), .A2(n11582), .ZN(n11584) );
  AND2_X1 U14764 ( .A1(n11586), .A2(n11584), .ZN(n17150) );
  NOR2_X1 U14765 ( .A1(n20196), .A2(n17150), .ZN(n16584) );
  NAND2_X1 U14766 ( .A1(n11586), .A2(n10352), .ZN(n11587) );
  NAND2_X1 U14767 ( .A1(n11585), .A2(n11587), .ZN(n17135) );
  NAND2_X1 U14768 ( .A1(n16584), .A2(n17135), .ZN(n20160) );
  NAND2_X1 U14769 ( .A1(n11585), .A2(n17126), .ZN(n11588) );
  AND2_X1 U14770 ( .A1(n10353), .A2(n11588), .ZN(n20161) );
  OR2_X1 U14771 ( .A1(n20160), .A2(n20161), .ZN(n20163) );
  INV_X1 U14772 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11589) );
  NAND2_X1 U14773 ( .A1(n10353), .A2(n11589), .ZN(n11590) );
  AND2_X1 U14774 ( .A1(n9835), .A2(n11590), .ZN(n17116) );
  NOR2_X1 U14775 ( .A1(n20163), .A2(n17116), .ZN(n20146) );
  INV_X1 U14776 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11592) );
  NAND2_X1 U14777 ( .A1(n9835), .A2(n11592), .ZN(n11593) );
  NAND2_X1 U14778 ( .A1(n11591), .A2(n11593), .ZN(n20149) );
  NAND2_X1 U14779 ( .A1(n20146), .A2(n20149), .ZN(n20136) );
  NAND2_X1 U14780 ( .A1(n11591), .A2(n17090), .ZN(n11595) );
  AND2_X1 U14781 ( .A1(n11594), .A2(n11595), .ZN(n20137) );
  OR2_X1 U14782 ( .A1(n20136), .A2(n20137), .ZN(n16560) );
  NAND2_X1 U14783 ( .A1(n11594), .A2(n17071), .ZN(n11597) );
  AND2_X1 U14784 ( .A1(n11596), .A2(n11597), .ZN(n17069) );
  NOR2_X1 U14785 ( .A1(n16560), .A2(n17069), .ZN(n16555) );
  NAND2_X1 U14786 ( .A1(n11596), .A2(n11598), .ZN(n11599) );
  NAND2_X1 U14787 ( .A1(n9830), .A2(n11599), .ZN(n17057) );
  AND2_X1 U14788 ( .A1(n16555), .A2(n17057), .ZN(n16544) );
  NAND2_X1 U14789 ( .A1(n9830), .A2(n10343), .ZN(n11601) );
  NAND2_X1 U14790 ( .A1(n11600), .A2(n11601), .ZN(n17041) );
  NAND2_X1 U14791 ( .A1(n16544), .A2(n17041), .ZN(n20118) );
  NAND2_X1 U14792 ( .A1(n11600), .A2(n17029), .ZN(n11603) );
  AND2_X1 U14793 ( .A1(n11602), .A2(n11603), .ZN(n20120) );
  OR2_X1 U14794 ( .A1(n20118), .A2(n20120), .ZN(n20121) );
  NAND2_X1 U14795 ( .A1(n11602), .A2(n17020), .ZN(n11604) );
  AND2_X1 U14796 ( .A1(n9834), .A2(n11604), .ZN(n20112) );
  NOR2_X1 U14797 ( .A1(n20121), .A2(n20112), .ZN(n20093) );
  NAND2_X1 U14798 ( .A1(n9831), .A2(n10348), .ZN(n11605) );
  NAND2_X1 U14799 ( .A1(n9827), .A2(n11605), .ZN(n20078) );
  INV_X1 U14800 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20102) );
  NAND2_X1 U14801 ( .A1(n9834), .A2(n20102), .ZN(n11606) );
  NAND2_X1 U14802 ( .A1(n9831), .A2(n11606), .ZN(n20095) );
  NAND3_X1 U14803 ( .A1(n20093), .A2(n20078), .A3(n20095), .ZN(n11607) );
  NAND2_X1 U14804 ( .A1(n9827), .A2(n11608), .ZN(n11609) );
  NAND2_X1 U14805 ( .A1(n11610), .A2(n11609), .ZN(n16993) );
  NAND2_X1 U14806 ( .A1(n16516), .A2(n10322), .ZN(n11613) );
  INV_X1 U14807 ( .A(n11611), .ZN(n11616) );
  INV_X1 U14808 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16506) );
  NAND2_X1 U14809 ( .A1(n11156), .A2(n16506), .ZN(n11612) );
  NAND2_X1 U14810 ( .A1(n11616), .A2(n11612), .ZN(n16983) );
  NAND2_X1 U14811 ( .A1(n11613), .A2(n16983), .ZN(n16488) );
  INV_X1 U14812 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11615) );
  NAND2_X1 U14813 ( .A1(n11616), .A2(n11615), .ZN(n11617) );
  NAND2_X1 U14814 ( .A1(n11614), .A2(n11617), .ZN(n16489) );
  NAND2_X1 U14815 ( .A1(n11614), .A2(n17813), .ZN(n11619) );
  NAND2_X1 U14816 ( .A1(n11621), .A2(n11619), .ZN(n17815) );
  NAND2_X1 U14817 ( .A1(n16476), .A2(n10322), .ZN(n11623) );
  NAND2_X1 U14818 ( .A1(n11621), .A2(n16475), .ZN(n11622) );
  NAND2_X1 U14819 ( .A1(n11620), .A2(n11622), .ZN(n16962) );
  NAND2_X1 U14820 ( .A1(n11623), .A2(n16962), .ZN(n16477) );
  NAND2_X1 U14821 ( .A1(n16477), .A2(n10322), .ZN(n11626) );
  NAND2_X1 U14822 ( .A1(n11620), .A2(n11624), .ZN(n11625) );
  NAND2_X1 U14823 ( .A1(n9859), .A2(n11625), .ZN(n16951) );
  NAND2_X1 U14824 ( .A1(n11626), .A2(n16951), .ZN(n16439) );
  NAND2_X1 U14825 ( .A1(n9859), .A2(n10354), .ZN(n11628) );
  AND2_X1 U14826 ( .A1(n11627), .A2(n11628), .ZN(n16942) );
  NAND2_X1 U14827 ( .A1(n11627), .A2(n16423), .ZN(n11630) );
  NAND2_X1 U14828 ( .A1(n11632), .A2(n11630), .ZN(n16924) );
  INV_X1 U14829 ( .A(n11631), .ZN(n11635) );
  NAND2_X1 U14830 ( .A1(n11632), .A2(n16412), .ZN(n11633) );
  INV_X1 U14831 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11634) );
  NAND2_X1 U14832 ( .A1(n11635), .A2(n11634), .ZN(n11636) );
  NAND2_X1 U14833 ( .A1(n9856), .A2(n11636), .ZN(n16398) );
  INV_X1 U14834 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16912) );
  NAND2_X1 U14835 ( .A1(n9856), .A2(n16912), .ZN(n11638) );
  AND2_X1 U14836 ( .A1(n11637), .A2(n11638), .ZN(n16914) );
  AND2_X1 U14837 ( .A1(n11639), .A2(n20910), .ZN(n13213) );
  INV_X1 U14838 ( .A(n20197), .ZN(n20177) );
  AOI21_X1 U14839 ( .B1(n15437), .B2(n20197), .A(n20107), .ZN(n11671) );
  XNOR2_X1 U14840 ( .A(n11637), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16904) );
  INV_X1 U14841 ( .A(n16904), .ZN(n11670) );
  NOR2_X1 U14842 ( .A1(n16649), .A2(n16904), .ZN(n15436) );
  NAND2_X1 U14843 ( .A1(n10328), .A2(n15436), .ZN(n11669) );
  OAI21_X1 U14844 ( .B1(n11640), .B2(n11642), .A(n11641), .ZN(n16906) );
  NAND2_X1 U14845 ( .A1(n11185), .A2(n11644), .ZN(n20190) );
  NAND2_X1 U14846 ( .A1(n20966), .A2(n20910), .ZN(n11658) );
  NOR2_X1 U14847 ( .A1(n10876), .A2(n11658), .ZN(n11646) );
  INV_X1 U14848 ( .A(n11648), .ZN(n11649) );
  AND2_X1 U14849 ( .A1(n20910), .A2(n13215), .ZN(n11660) );
  AND2_X1 U14850 ( .A1(n11651), .A2(n11660), .ZN(n14403) );
  NAND2_X1 U14851 ( .A1(n11658), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n11652) );
  NOR2_X1 U14852 ( .A1(n10876), .A2(n11652), .ZN(n11653) );
  NAND2_X1 U14853 ( .A1(n20053), .A2(n11653), .ZN(n20165) );
  NAND2_X1 U14854 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20939), .ZN(n14500) );
  NOR3_X1 U14855 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n17491), .A3(n14500), 
        .ZN(n14408) );
  INV_X1 U14856 ( .A(n14408), .ZN(n11654) );
  NAND2_X1 U14857 ( .A1(n20181), .A2(n11654), .ZN(n11655) );
  OR2_X1 U14858 ( .A1(n20197), .A2(n11655), .ZN(n11656) );
  NAND2_X1 U14859 ( .A1(n11658), .A2(n11657), .ZN(n11659) );
  OR2_X1 U14860 ( .A1(n13221), .A2(n11659), .ZN(n11661) );
  AOI21_X1 U14861 ( .B1(n13296), .B2(n11661), .A(n11660), .ZN(n20126) );
  AOI22_X1 U14862 ( .A1(n20150), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n20169), 
        .B2(P2_EBX_REG_30__SCAN_IN), .ZN(n11663) );
  NAND2_X1 U14863 ( .A1(n20186), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11662) );
  OAI211_X1 U14864 ( .C1(n11664), .C2(n20165), .A(n11663), .B(n11662), .ZN(
        n11665) );
  AOI21_X1 U14865 ( .B1(n16773), .B2(n20185), .A(n11665), .ZN(n11666) );
  OAI21_X1 U14866 ( .B1(n16906), .B2(n20189), .A(n11666), .ZN(n11667) );
  OAI211_X1 U14867 ( .C1(n11671), .C2(n11670), .A(n11669), .B(n11668), .ZN(
        P2_U2825) );
  AOI22_X1 U14868 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U14869 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11716), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11680) );
  NOR2_X1 U14870 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11672) );
  INV_X1 U14871 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11676) );
  AND2_X2 U14872 ( .A1(n11682), .A2(n11684), .ZN(n17785) );
  NAND2_X1 U14873 ( .A1(n17785), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11675) );
  NAND2_X1 U14874 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11674) );
  OAI211_X1 U14875 ( .C1(n9756), .C2(n11676), .A(n11675), .B(n11674), .ZN(
        n11677) );
  INV_X1 U14876 ( .A(n11677), .ZN(n11679) );
  INV_X2 U14877 ( .A(n11693), .ZN(n17782) );
  AOI22_X1 U14878 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11678) );
  AND2_X1 U14879 ( .A1(n11684), .A2(n13393), .ZN(n11703) );
  AOI22_X1 U14880 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11703), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11692) );
  AND2_X2 U14881 ( .A1(n11685), .A2(n11683), .ZN(n11725) );
  AOI22_X1 U14882 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11691) );
  INV_X2 U14883 ( .A(n9749), .ZN(n18543) );
  AOI22_X1 U14884 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11690) );
  INV_X1 U14885 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11688) );
  OR2_X1 U14886 ( .A1(n17765), .A2(n11688), .ZN(n11689) );
  NAND2_X1 U14887 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11697) );
  INV_X2 U14888 ( .A(n11693), .ZN(n12008) );
  NAND2_X1 U14889 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11696) );
  NAND2_X1 U14890 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11695) );
  NAND2_X1 U14891 ( .A1(n13472), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11694) );
  NAND4_X1 U14892 ( .A1(n11697), .A2(n11696), .A3(n11695), .A4(n11694), .ZN(
        n11702) );
  NAND2_X1 U14893 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11700) );
  INV_X2 U14894 ( .A(n9749), .ZN(n17699) );
  NAND2_X1 U14895 ( .A1(n17699), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11699) );
  NAND2_X1 U14896 ( .A1(n17784), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11698) );
  NAND3_X1 U14897 ( .A1(n11700), .A2(n11699), .A3(n11698), .ZN(n11701) );
  NOR2_X1 U14898 ( .A1(n11702), .A2(n11701), .ZN(n11715) );
  AOI22_X1 U14899 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11716), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11714) );
  NAND2_X1 U14900 ( .A1(n17682), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11707) );
  NAND2_X1 U14901 ( .A1(n17755), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11706) );
  NAND2_X1 U14902 ( .A1(n9690), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11705) );
  INV_X2 U14903 ( .A(n9746), .ZN(n17700) );
  NAND2_X1 U14904 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11704) );
  INV_X2 U14905 ( .A(n9867), .ZN(n17765) );
  INV_X1 U14906 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11710) );
  NAND2_X1 U14907 ( .A1(n17785), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11709) );
  NAND2_X1 U14908 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11708) );
  OAI211_X1 U14909 ( .C1(n17765), .C2(n11710), .A(n11709), .B(n11708), .ZN(
        n11711) );
  INV_X1 U14910 ( .A(n11711), .ZN(n11712) );
  AOI22_X1 U14911 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11716), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11724) );
  INV_X1 U14912 ( .A(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11719) );
  NAND2_X1 U14913 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11718) );
  NAND2_X1 U14914 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11717) );
  OAI211_X1 U14915 ( .C1(n9756), .C2(n11719), .A(n11718), .B(n11717), .ZN(
        n11720) );
  INV_X1 U14916 ( .A(n11720), .ZN(n11723) );
  AOI22_X1 U14917 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11722) );
  AOI22_X1 U14918 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17774), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11721) );
  NAND4_X1 U14919 ( .A1(n11724), .A2(n11723), .A3(n11722), .A4(n11721), .ZN(
        n11731) );
  INV_X2 U14920 ( .A(n13314), .ZN(n17762) );
  AOI22_X1 U14921 ( .A1(n17762), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11725), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11729) );
  AOI22_X1 U14922 ( .A1(n17682), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11728) );
  AOI22_X1 U14923 ( .A1(n9690), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11727) );
  INV_X1 U14924 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17766) );
  OR2_X1 U14925 ( .A1(n18545), .A2(n17766), .ZN(n11726) );
  NAND4_X1 U14926 ( .A1(n11729), .A2(n11728), .A3(n11727), .A4(n11726), .ZN(
        n11730) );
  AOI22_X1 U14927 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U14928 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11734) );
  AOI22_X1 U14929 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11733) );
  NAND2_X1 U14930 ( .A1(n17785), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11732) );
  INV_X1 U14931 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11738) );
  NAND2_X1 U14932 ( .A1(n9690), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11737) );
  NAND2_X1 U14933 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11736) );
  OAI211_X1 U14934 ( .C1(n17765), .C2(n11738), .A(n11737), .B(n11736), .ZN(
        n11744) );
  NAND2_X1 U14935 ( .A1(n17755), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11742) );
  NAND2_X1 U14936 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11741) );
  NAND2_X1 U14937 ( .A1(n17682), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11740) );
  NAND2_X1 U14938 ( .A1(n17699), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11739) );
  NAND4_X1 U14939 ( .A1(n11742), .A2(n11741), .A3(n11740), .A4(n11739), .ZN(
        n11743) );
  NOR2_X1 U14940 ( .A1(n11744), .A2(n11743), .ZN(n11746) );
  AOI22_X1 U14941 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11745) );
  INV_X2 U14942 ( .A(n18539), .ZN(n18523) );
  AOI22_X1 U14943 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11754) );
  NAND2_X1 U14944 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11750) );
  NAND2_X1 U14945 ( .A1(n17699), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11749) );
  NAND2_X1 U14946 ( .A1(n17784), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11748) );
  AND3_X1 U14947 ( .A1(n11750), .A2(n11749), .A3(n11748), .ZN(n11753) );
  BUF_X2 U14948 ( .A(n13351), .Z(n18550) );
  AOI22_X1 U14949 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U14950 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17774), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11751) );
  NAND4_X1 U14951 ( .A1(n11754), .A2(n11753), .A3(n11752), .A4(n11751), .ZN(
        n11761) );
  AOI22_X1 U14952 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11725), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11759) );
  AOI22_X1 U14953 ( .A1(n17762), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U14954 ( .A1(n17682), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11757) );
  INV_X1 U14955 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11755) );
  OR2_X1 U14956 ( .A1(n18545), .A2(n11755), .ZN(n11756) );
  NAND4_X1 U14957 ( .A1(n11759), .A2(n11758), .A3(n11757), .A4(n11756), .ZN(
        n11760) );
  AOI22_X1 U14958 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11769) );
  INV_X1 U14959 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11764) );
  NAND2_X1 U14960 ( .A1(n17785), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11763) );
  NAND2_X1 U14961 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11762) );
  OAI211_X1 U14962 ( .C1(n9756), .C2(n11764), .A(n11763), .B(n11762), .ZN(
        n11765) );
  INV_X1 U14963 ( .A(n11765), .ZN(n11768) );
  AOI22_X1 U14964 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11767) );
  AOI22_X1 U14965 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11766) );
  NAND4_X1 U14966 ( .A1(n11769), .A2(n11768), .A3(n11767), .A4(n11766), .ZN(
        n11775) );
  INV_X2 U14967 ( .A(n12012), .ZN(n18542) );
  AOI22_X1 U14968 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U14969 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11772) );
  AOI22_X1 U14970 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11771) );
  INV_X1 U14971 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18462) );
  OR2_X1 U14972 ( .A1(n18545), .A2(n18462), .ZN(n11770) );
  NAND4_X1 U14973 ( .A1(n11773), .A2(n11772), .A3(n11771), .A4(n11770), .ZN(
        n11774) );
  NAND2_X1 U14974 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11779) );
  NAND2_X1 U14975 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11778) );
  NAND2_X1 U14976 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11777) );
  NAND2_X1 U14977 ( .A1(n17755), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11776) );
  NAND4_X1 U14978 ( .A1(n11779), .A2(n11778), .A3(n11777), .A4(n11776), .ZN(
        n11784) );
  INV_X1 U14979 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11782) );
  NAND2_X1 U14980 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11781) );
  NAND2_X1 U14981 ( .A1(n13472), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11780) );
  OAI211_X1 U14982 ( .C1(n11782), .C2(n17769), .A(n11781), .B(n11780), .ZN(
        n11783) );
  NOR2_X1 U14983 ( .A1(n11784), .A2(n11783), .ZN(n11796) );
  INV_X1 U14984 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18471) );
  INV_X1 U14985 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11785) );
  OAI22_X1 U14986 ( .A1(n18464), .A2(n18471), .B1(n17767), .B2(n11785), .ZN(
        n11787) );
  INV_X1 U14987 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17727) );
  INV_X1 U14988 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14067) );
  OAI22_X1 U14989 ( .A1(n12012), .A2(n17727), .B1(n9749), .B2(n14067), .ZN(
        n11786) );
  NOR2_X1 U14990 ( .A1(n11787), .A2(n11786), .ZN(n11795) );
  INV_X1 U14991 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19453) );
  AOI22_X1 U14992 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18523), .B1(
        n18524), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11794) );
  INV_X1 U14993 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11788) );
  NOR2_X1 U14994 ( .A1(n17765), .A2(n11788), .ZN(n11792) );
  INV_X1 U14995 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11790) );
  INV_X1 U14996 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11789) );
  OAI22_X1 U14997 ( .A1(n13314), .A2(n11790), .B1(n9756), .B2(n11789), .ZN(
        n11791) );
  NOR2_X1 U14998 ( .A1(n11792), .A2(n11791), .ZN(n11793) );
  NAND2_X1 U14999 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11800) );
  NAND2_X1 U15000 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11799) );
  NAND2_X1 U15001 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11798) );
  NAND2_X1 U15002 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11797) );
  NAND4_X1 U15003 ( .A1(n11800), .A2(n11799), .A3(n11798), .A4(n11797), .ZN(
        n11805) );
  NAND2_X1 U15004 ( .A1(n17699), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11803) );
  NAND2_X1 U15005 ( .A1(n13472), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11802) );
  NAND2_X1 U15006 ( .A1(n17784), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11801) );
  NAND3_X1 U15007 ( .A1(n11803), .A2(n11802), .A3(n11801), .ZN(n11804) );
  NOR2_X1 U15008 ( .A1(n11805), .A2(n11804), .ZN(n11816) );
  NAND2_X1 U15009 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11809) );
  NAND2_X1 U15010 ( .A1(n17682), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11808) );
  NAND2_X1 U15011 ( .A1(n9690), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11807) );
  NAND2_X1 U15012 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11806) );
  AND4_X1 U15013 ( .A1(n11809), .A2(n11808), .A3(n11807), .A4(n11806), .ZN(
        n11814) );
  INV_X1 U15014 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14136) );
  NAND2_X1 U15015 ( .A1(n17785), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11811) );
  NAND2_X1 U15016 ( .A1(n17755), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11810) );
  OAI211_X1 U15017 ( .C1(n17765), .C2(n14136), .A(n11811), .B(n11810), .ZN(
        n11812) );
  INV_X1 U15018 ( .A(n11812), .ZN(n11813) );
  AND2_X1 U15019 ( .A1(n13441), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13447) );
  NAND2_X1 U15020 ( .A1(n13448), .A2(n13447), .ZN(n13446) );
  INV_X1 U15021 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19379) );
  NAND2_X1 U15022 ( .A1(n13446), .A2(n11817), .ZN(n19106) );
  INV_X1 U15023 ( .A(n13458), .ZN(n11818) );
  NAND2_X1 U15024 ( .A1(n19106), .A2(n19107), .ZN(n19109) );
  INV_X1 U15025 ( .A(n11820), .ZN(n11821) );
  NAND2_X1 U15026 ( .A1(n11821), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11822) );
  NAND2_X2 U15027 ( .A1(n19109), .A2(n11822), .ZN(n11826) );
  OAI21_X1 U15028 ( .B1(n11823), .B2(n13511), .A(n11828), .ZN(n11824) );
  XNOR2_X2 U15029 ( .A(n11826), .B(n11824), .ZN(n19093) );
  INV_X1 U15030 ( .A(n11824), .ZN(n11825) );
  NAND2_X1 U15031 ( .A1(n11826), .A2(n11825), .ZN(n11827) );
  XNOR2_X1 U15032 ( .A(n11828), .B(n13608), .ZN(n11829) );
  XNOR2_X1 U15033 ( .A(n11829), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19076) );
  INV_X1 U15034 ( .A(n11829), .ZN(n11830) );
  NAND2_X1 U15035 ( .A1(n11830), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11831) );
  NOR2_X1 U15036 ( .A1(n11832), .A2(n12083), .ZN(n11833) );
  INV_X1 U15037 ( .A(n11834), .ZN(n11835) );
  XNOR2_X1 U15038 ( .A(n11839), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19049) );
  INV_X1 U15039 ( .A(n11839), .ZN(n11840) );
  NAND2_X1 U15040 ( .A1(n11840), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11841) );
  NAND2_X1 U15041 ( .A1(n18950), .A2(n11843), .ZN(n11844) );
  NAND2_X1 U15042 ( .A1(n11845), .A2(n9985), .ZN(n11846) );
  INV_X1 U15043 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11848) );
  INV_X1 U15044 ( .A(n18938), .ZN(n18965) );
  INV_X1 U15045 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n19245) );
  INV_X1 U15046 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11852) );
  INV_X1 U15047 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11851) );
  INV_X1 U15048 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11850) );
  NAND2_X1 U15049 ( .A1(n18965), .A2(n10539), .ZN(n11853) );
  NAND2_X1 U15050 ( .A1(n11853), .A2(n18950), .ZN(n18919) );
  OR2_X1 U15051 ( .A1(n18950), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11854) );
  NOR2_X1 U15052 ( .A1(n11849), .A2(n11847), .ZN(n19287) );
  NAND2_X1 U15053 ( .A1(n19287), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n19272) );
  NOR2_X1 U15054 ( .A1(n19272), .A2(n11850), .ZN(n19247) );
  AND2_X1 U15055 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11855) );
  NAND2_X1 U15056 ( .A1(n19247), .A2(n11855), .ZN(n19222) );
  INV_X1 U15057 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n19210) );
  AND2_X1 U15058 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n19199) );
  INV_X1 U15059 ( .A(n19199), .ZN(n19157) );
  AND2_X1 U15060 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11859) );
  AND2_X1 U15061 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n19176) );
  AND3_X1 U15062 ( .A1(n11859), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n19176), .ZN(n11858) );
  AND3_X1 U15063 ( .A1(n19199), .A2(n19176), .A3(n11859), .ZN(n19168) );
  NAND2_X1 U15064 ( .A1(n19168), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18797) );
  INV_X1 U15065 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17672) );
  NOR2_X1 U15066 ( .A1(n18797), .A2(n17672), .ZN(n17671) );
  INV_X1 U15067 ( .A(n17671), .ZN(n17598) );
  INV_X1 U15068 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n19203) );
  AND2_X1 U15069 ( .A1(n18950), .A2(n19203), .ZN(n18901) );
  INV_X1 U15070 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18885) );
  NAND2_X1 U15071 ( .A1(n18901), .A2(n18885), .ZN(n11860) );
  NOR2_X1 U15072 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11860), .ZN(
        n18862) );
  INV_X1 U15073 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n19164) );
  INV_X1 U15074 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18855) );
  NAND4_X1 U15075 ( .A1(n18862), .A2(n17672), .A3(n19164), .A4(n18855), .ZN(
        n11861) );
  OAI21_X1 U15076 ( .B1(n11856), .B2(n17598), .A(n11861), .ZN(n11862) );
  INV_X1 U15077 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18799) );
  AND2_X1 U15078 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17652) );
  INV_X1 U15079 ( .A(n18821), .ZN(n11863) );
  INV_X1 U15080 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17662) );
  INV_X1 U15081 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13381) );
  NAND2_X1 U15082 ( .A1(n13381), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12157) );
  NAND3_X1 U15083 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17554) );
  NOR2_X2 U15084 ( .A1(n11866), .A2(n17554), .ZN(n17550) );
  INV_X1 U15085 ( .A(n17550), .ZN(n11867) );
  OAI211_X1 U15086 ( .C1(n17551), .C2(n18966), .A(n12157), .B(n11867), .ZN(
        n11871) );
  INV_X1 U15087 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11868) );
  NOR2_X1 U15088 ( .A1(n18950), .A2(n11868), .ZN(n11869) );
  MUX2_X1 U15089 ( .A(n18950), .B(n11869), .S(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .Z(n11870) );
  NOR2_X1 U15090 ( .A1(n13381), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12168) );
  AOI22_X1 U15091 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11878) );
  INV_X1 U15092 ( .A(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18463) );
  NAND2_X1 U15093 ( .A1(n17785), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11873) );
  NAND2_X1 U15094 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11872) );
  OAI211_X1 U15095 ( .C1(n9756), .C2(n18463), .A(n11873), .B(n11872), .ZN(
        n11874) );
  INV_X1 U15096 ( .A(n11874), .ZN(n11877) );
  AOI22_X1 U15097 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U15098 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U15099 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U15100 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U15101 ( .A1(n17755), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11880) );
  INV_X1 U15102 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17536) );
  OR2_X1 U15103 ( .A1(n18545), .A2(n17536), .ZN(n11879) );
  NAND2_X1 U15104 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11886) );
  NAND2_X1 U15105 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11885) );
  NAND2_X1 U15106 ( .A1(n17682), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11884) );
  NAND2_X1 U15107 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11883) );
  NAND4_X1 U15108 ( .A1(n11886), .A2(n11885), .A3(n11884), .A4(n11883), .ZN(
        n11891) );
  NAND2_X1 U15109 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11889) );
  NAND2_X1 U15110 ( .A1(n13472), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11888) );
  NAND2_X1 U15111 ( .A1(n17784), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11887) );
  NAND3_X1 U15112 ( .A1(n11889), .A2(n11888), .A3(n11887), .ZN(n11890) );
  NOR2_X1 U15113 ( .A1(n11891), .A2(n11890), .ZN(n11903) );
  AOI22_X1 U15114 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11716), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11902) );
  NAND2_X1 U15115 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11895) );
  NAND2_X1 U15116 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11894) );
  NAND2_X1 U15117 ( .A1(n9690), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11893) );
  NAND2_X1 U15118 ( .A1(n17699), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11892) );
  INV_X1 U15119 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11898) );
  INV_X1 U15120 ( .A(n13314), .ZN(n11944) );
  INV_X1 U15121 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n19652) );
  NAND2_X1 U15122 ( .A1(n11944), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11897) );
  NAND2_X1 U15123 ( .A1(n17755), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11896) );
  OAI211_X1 U15124 ( .C1(n17765), .C2(n11898), .A(n11897), .B(n11896), .ZN(
        n11899) );
  INV_X1 U15125 ( .A(n11899), .ZN(n11900) );
  NAND4_X1 U15126 ( .A1(n11903), .A2(n11902), .A3(n11901), .A4(n11900), .ZN(
        n19436) );
  NAND2_X1 U15127 ( .A1(n13546), .A2(n13322), .ZN(n12025) );
  INV_X1 U15128 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11906) );
  NAND2_X1 U15129 ( .A1(n11944), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11905) );
  NAND2_X1 U15130 ( .A1(n9690), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11904) );
  OAI211_X1 U15131 ( .C1(n18545), .C2(n11906), .A(n11905), .B(n11904), .ZN(
        n11912) );
  NAND2_X1 U15132 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11910) );
  NAND2_X1 U15133 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11909) );
  NAND2_X1 U15134 ( .A1(n17682), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11908) );
  NAND2_X1 U15135 ( .A1(n13472), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11907) );
  NAND4_X1 U15136 ( .A1(n11910), .A2(n11909), .A3(n11908), .A4(n11907), .ZN(
        n11911) );
  NOR2_X1 U15137 ( .A1(n11912), .A2(n11911), .ZN(n11923) );
  AOI22_X1 U15138 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11922) );
  INV_X1 U15139 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18518) );
  NAND2_X1 U15140 ( .A1(n17755), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11914) );
  NAND2_X1 U15141 ( .A1(n17784), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11913) );
  OAI211_X1 U15142 ( .C1(n11693), .C2(n18518), .A(n11914), .B(n11913), .ZN(
        n11915) );
  INV_X1 U15143 ( .A(n11915), .ZN(n11921) );
  NAND2_X1 U15144 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11919) );
  NAND2_X1 U15145 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11918) );
  NAND2_X1 U15146 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11917) );
  NAND2_X1 U15147 ( .A1(n17699), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11916) );
  NAND2_X1 U15148 ( .A1(n19443), .A2(n19440), .ZN(n12032) );
  NAND2_X1 U15149 ( .A1(n12025), .A2(n12032), .ZN(n11963) );
  INV_X1 U15150 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13547) );
  NAND2_X1 U15151 ( .A1(n9690), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11925) );
  NAND2_X1 U15152 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11924) );
  OAI211_X1 U15153 ( .C1(n17765), .C2(n13547), .A(n11925), .B(n11924), .ZN(
        n11931) );
  NAND2_X1 U15154 ( .A1(n17755), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11929) );
  NAND2_X1 U15155 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11928) );
  NAND2_X1 U15156 ( .A1(n17682), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11927) );
  NAND2_X1 U15157 ( .A1(n17699), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11926) );
  NAND4_X1 U15158 ( .A1(n11929), .A2(n11928), .A3(n11927), .A4(n11926), .ZN(
        n11930) );
  NOR2_X1 U15159 ( .A1(n11931), .A2(n11930), .ZN(n11943) );
  AOI22_X1 U15160 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11942) );
  INV_X1 U15161 ( .A(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11934) );
  INV_X1 U15162 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n19640) );
  NAND2_X1 U15163 ( .A1(n17785), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11933) );
  NAND2_X1 U15164 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11932) );
  OAI211_X1 U15165 ( .C1(n9756), .C2(n11934), .A(n11933), .B(n11932), .ZN(
        n11935) );
  INV_X1 U15166 ( .A(n11935), .ZN(n11941) );
  NAND2_X1 U15167 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11939) );
  NAND2_X1 U15168 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11938) );
  NAND2_X1 U15169 ( .A1(n13472), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11937) );
  NAND2_X1 U15170 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11936) );
  AOI22_X1 U15171 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U15172 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U15173 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11946) );
  INV_X1 U15174 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n19646) );
  NAND2_X1 U15175 ( .A1(n11944), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11945) );
  INV_X1 U15176 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11951) );
  NAND2_X1 U15177 ( .A1(n9690), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11950) );
  NAND2_X1 U15178 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11949) );
  OAI211_X1 U15179 ( .C1(n18545), .C2(n11951), .A(n11950), .B(n11949), .ZN(
        n11957) );
  NAND2_X1 U15180 ( .A1(n17755), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11955) );
  NAND2_X1 U15181 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11954) );
  NAND2_X1 U15182 ( .A1(n17682), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11953) );
  NAND2_X1 U15183 ( .A1(n17699), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11952) );
  NAND4_X1 U15184 ( .A1(n11955), .A2(n11954), .A3(n11953), .A4(n11952), .ZN(
        n11956) );
  NOR2_X1 U15185 ( .A1(n11957), .A2(n11956), .ZN(n11959) );
  AOI22_X1 U15186 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11958) );
  NAND2_X1 U15187 ( .A1(n10081), .A2(n19426), .ZN(n11961) );
  NAND2_X1 U15188 ( .A1(n13433), .A2(n11961), .ZN(n11962) );
  NAND2_X1 U15189 ( .A1(n11963), .A2(n11962), .ZN(n12024) );
  INV_X1 U15190 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13346) );
  NAND2_X1 U15191 ( .A1(n17785), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11965) );
  NAND2_X1 U15192 ( .A1(n9690), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11964) );
  OAI211_X1 U15193 ( .C1(n17765), .C2(n13346), .A(n11965), .B(n11964), .ZN(
        n11971) );
  NAND2_X1 U15194 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11969) );
  NAND2_X1 U15195 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11968) );
  NAND2_X1 U15196 ( .A1(n17682), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11967) );
  NAND2_X1 U15197 ( .A1(n17784), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11966) );
  NAND4_X1 U15198 ( .A1(n11969), .A2(n11968), .A3(n11967), .A4(n11966), .ZN(
        n11970) );
  NAND2_X1 U15199 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11974) );
  NAND2_X1 U15200 ( .A1(n17755), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11973) );
  NAND2_X1 U15201 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11972) );
  NAND2_X1 U15202 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11978) );
  NAND2_X1 U15203 ( .A1(n13472), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11977) );
  NAND2_X1 U15204 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11976) );
  NAND2_X1 U15205 ( .A1(n17699), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11975) );
  NAND2_X1 U15206 ( .A1(n10081), .A2(n20031), .ZN(n11983) );
  NAND2_X1 U15207 ( .A1(n11983), .A2(n19426), .ZN(n12071) );
  NAND2_X1 U15208 ( .A1(n12071), .A2(n12032), .ZN(n12023) );
  INV_X1 U15209 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11986) );
  NAND2_X1 U15210 ( .A1(n17762), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11985) );
  NAND2_X1 U15211 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11984) );
  OAI211_X1 U15212 ( .C1(n17765), .C2(n11986), .A(n11985), .B(n11984), .ZN(
        n11992) );
  NAND2_X1 U15213 ( .A1(n17682), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11990) );
  NAND2_X1 U15214 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11989) );
  NAND2_X1 U15215 ( .A1(n9690), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11988) );
  NAND2_X1 U15216 ( .A1(n17699), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11987) );
  NAND4_X1 U15217 ( .A1(n11990), .A2(n11989), .A3(n11988), .A4(n11987), .ZN(
        n11991) );
  NOR2_X1 U15218 ( .A1(n11992), .A2(n11991), .ZN(n12004) );
  AOI22_X1 U15219 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18524), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12003) );
  NAND2_X1 U15220 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11996) );
  NAND2_X1 U15221 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11995) );
  NAND2_X1 U15222 ( .A1(n17755), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11994) );
  NAND2_X1 U15223 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11993) );
  NAND4_X1 U15224 ( .A1(n11996), .A2(n11995), .A3(n11994), .A4(n11993), .ZN(
        n12001) );
  NAND2_X1 U15225 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11999) );
  NAND2_X1 U15226 ( .A1(n13472), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11998) );
  NAND2_X1 U15227 ( .A1(n17784), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11997) );
  NAND3_X1 U15228 ( .A1(n11999), .A2(n11998), .A3(n11997), .ZN(n12000) );
  AOI22_X1 U15229 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12011) );
  NAND2_X1 U15230 ( .A1(n9690), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12007) );
  NAND2_X1 U15231 ( .A1(n13472), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12006) );
  NAND2_X1 U15232 ( .A1(n17784), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12005) );
  AOI22_X1 U15233 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18552), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U15234 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17699), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12009) );
  NAND4_X1 U15235 ( .A1(n12011), .A2(n10541), .A3(n12010), .A4(n12009), .ZN(
        n12019) );
  INV_X1 U15236 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n19649) );
  BUF_X1 U15237 ( .A(n13345), .Z(n17705) );
  AOI22_X1 U15238 ( .A1(n17762), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17705), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U15239 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U15240 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12015) );
  INV_X1 U15241 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12013) );
  NAND4_X1 U15242 ( .A1(n12017), .A2(n12016), .A3(n12015), .A4(n12014), .ZN(
        n12018) );
  INV_X1 U15243 ( .A(n19431), .ZN(n12033) );
  NAND2_X1 U15244 ( .A1(n12034), .A2(n12033), .ZN(n12022) );
  NAND2_X1 U15245 ( .A1(n19448), .A2(n12032), .ZN(n12020) );
  NAND2_X1 U15246 ( .A1(n12020), .A2(n19436), .ZN(n12021) );
  NAND4_X1 U15247 ( .A1(n12024), .A2(n12023), .A3(n12022), .A4(n12021), .ZN(
        n12140) );
  INV_X1 U15248 ( .A(n12140), .ZN(n12031) );
  INV_X1 U15249 ( .A(n12025), .ZN(n12028) );
  NAND2_X1 U15250 ( .A1(n13433), .A2(n19448), .ZN(n12027) );
  AND2_X1 U15251 ( .A1(n19420), .A2(n18681), .ZN(n12026) );
  NAND2_X1 U15252 ( .A1(n12027), .A2(n12026), .ZN(n12141) );
  OAI21_X1 U15253 ( .B1(n12028), .B2(n12153), .A(n12141), .ZN(n12029) );
  NAND2_X1 U15254 ( .A1(n12029), .A2(n19431), .ZN(n12030) );
  INV_X1 U15255 ( .A(n19440), .ZN(n12036) );
  NAND2_X1 U15256 ( .A1(n12036), .A2(n19443), .ZN(n12073) );
  INV_X1 U15257 ( .A(n12073), .ZN(n13323) );
  INV_X1 U15258 ( .A(n12034), .ZN(n12035) );
  NAND4_X1 U15259 ( .A1(n13323), .A2(n13372), .A3(n19420), .A4(n12035), .ZN(
        n12042) );
  AND3_X1 U15260 ( .A1(n12036), .A2(n19426), .A3(n13322), .ZN(n12038) );
  NOR3_X1 U15261 ( .A1(n19426), .A2(n19431), .A3(n19436), .ZN(n12039) );
  NAND2_X1 U15262 ( .A1(n18745), .A2(n12138), .ZN(n18032) );
  INV_X1 U15263 ( .A(n18745), .ZN(n12041) );
  NAND2_X1 U15264 ( .A1(n12041), .A2(n20031), .ZN(n13363) );
  INV_X1 U15265 ( .A(n13373), .ZN(n12043) );
  OR2_X2 U15266 ( .A1(n13362), .A2(n12043), .ZN(n19160) );
  NOR2_X4 U15267 ( .A1(n19160), .A2(n19876), .ZN(n19289) );
  NAND2_X1 U15268 ( .A1(n13373), .A2(n13372), .ZN(n12048) );
  INV_X1 U15269 ( .A(n12074), .ZN(n12044) );
  NAND3_X1 U15270 ( .A1(n20031), .A2(n12044), .A3(n14235), .ZN(n12046) );
  NAND2_X1 U15271 ( .A1(n12046), .A2(n12045), .ZN(n13371) );
  MUX2_X1 U15272 ( .A(n19858), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12066) );
  NAND2_X1 U15273 ( .A1(n12066), .A2(n12065), .ZN(n12051) );
  NAND2_X1 U15274 ( .A1(n19858), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12050) );
  NAND2_X1 U15275 ( .A1(n12051), .A2(n12050), .ZN(n12057) );
  INV_X1 U15276 ( .A(n12057), .ZN(n12052) );
  MUX2_X1 U15277 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n19409), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12056) );
  OAI22_X1 U15278 ( .A1(n12053), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19890), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12059) );
  NOR2_X1 U15279 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19890), .ZN(
        n12054) );
  NAND2_X1 U15280 ( .A1(n12053), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12060) );
  AOI22_X1 U15281 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12059), .B1(
        n12054), .B2(n12060), .ZN(n12064) );
  AND2_X1 U15282 ( .A1(n11687), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12055) );
  NOR2_X1 U15283 ( .A1(n12065), .A2(n12055), .ZN(n12069) );
  AND2_X1 U15284 ( .A1(n12066), .A2(n12069), .ZN(n12063) );
  XNOR2_X1 U15285 ( .A(n12057), .B(n12056), .ZN(n12058) );
  NAND2_X1 U15286 ( .A1(n12064), .A2(n12058), .ZN(n12062) );
  AOI21_X1 U15287 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12060), .A(
        n12059), .ZN(n12061) );
  INV_X1 U15288 ( .A(n19878), .ZN(n13368) );
  XNOR2_X1 U15289 ( .A(n12066), .B(n12065), .ZN(n12067) );
  NAND2_X1 U15290 ( .A1(n12068), .A2(n12067), .ZN(n12146) );
  OR2_X1 U15291 ( .A1(n12146), .A2(n12069), .ZN(n12070) );
  NAND2_X1 U15292 ( .A1(n12070), .A2(n12147), .ZN(n19880) );
  INV_X1 U15293 ( .A(n12071), .ZN(n12075) );
  NAND2_X1 U15294 ( .A1(n13433), .A2(n19436), .ZN(n12072) );
  NAND4_X1 U15295 ( .A1(n12075), .A2(n12074), .A3(n12073), .A4(n12072), .ZN(
        n12139) );
  NAND2_X1 U15296 ( .A1(n19426), .A2(n20031), .ZN(n12148) );
  NOR2_X1 U15297 ( .A1(n12148), .A2(n13546), .ZN(n12137) );
  INV_X1 U15298 ( .A(n12137), .ZN(n12076) );
  NAND2_X1 U15299 ( .A1(n19880), .A2(n19391), .ZN(n12077) );
  NAND2_X1 U15300 ( .A1(n18678), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n19920) );
  NOR2_X4 U15301 ( .A1(n18041), .A2(n19420), .ZN(n19119) );
  NAND2_X1 U15302 ( .A1(n12156), .A2(n19015), .ZN(n12136) );
  NAND2_X1 U15303 ( .A1(n12079), .A2(n12090), .ZN(n12087) );
  NAND2_X1 U15304 ( .A1(n12087), .A2(n13511), .ZN(n12086) );
  NOR2_X1 U15305 ( .A1(n12086), .A2(n13608), .ZN(n12084) );
  NAND2_X1 U15306 ( .A1(n12084), .A2(n12083), .ZN(n12082) );
  INV_X1 U15307 ( .A(n12081), .ZN(n13698) );
  NOR2_X1 U15308 ( .A1(n12082), .A2(n13698), .ZN(n12080) );
  AND2_X1 U15309 ( .A1(n12080), .A2(n17632), .ZN(n12109) );
  INV_X1 U15310 ( .A(n17632), .ZN(n17608) );
  XNOR2_X1 U15311 ( .A(n12080), .B(n17608), .ZN(n19041) );
  XNOR2_X1 U15312 ( .A(n12082), .B(n12081), .ZN(n12102) );
  INV_X1 U15313 ( .A(n12083), .ZN(n13693) );
  XNOR2_X1 U15314 ( .A(n12084), .B(n13693), .ZN(n12085) );
  NAND2_X1 U15315 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12085), .ZN(
        n12101) );
  INV_X1 U15316 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n19356) );
  XNOR2_X1 U15317 ( .A(n19356), .B(n12085), .ZN(n19064) );
  XOR2_X1 U15318 ( .A(n13608), .B(n12086), .Z(n12099) );
  XNOR2_X1 U15319 ( .A(n12087), .B(n13511), .ZN(n12088) );
  OR2_X1 U15320 ( .A1(n12088), .A2(n9976), .ZN(n12097) );
  XNOR2_X1 U15321 ( .A(n12088), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n19091) );
  INV_X1 U15322 ( .A(n12092), .ZN(n12091) );
  NAND2_X1 U15323 ( .A1(n12091), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12096) );
  XNOR2_X1 U15324 ( .A(n12092), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19103) );
  INV_X1 U15325 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13464) );
  AOI21_X1 U15326 ( .B1(n13458), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12093) );
  MUX2_X1 U15327 ( .A(n12093), .B(n13458), .S(n13441), .Z(n12095) );
  NOR2_X1 U15328 ( .A1(n13458), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12094) );
  NOR2_X1 U15329 ( .A1(n12095), .A2(n12094), .ZN(n19102) );
  NAND2_X1 U15330 ( .A1(n19103), .A2(n19102), .ZN(n19105) );
  NAND2_X1 U15331 ( .A1(n12099), .A2(n12098), .ZN(n12100) );
  NAND2_X1 U15332 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n19082), .ZN(
        n19081) );
  NAND2_X1 U15333 ( .A1(n12100), .A2(n19081), .ZN(n19063) );
  NAND2_X1 U15334 ( .A1(n19064), .A2(n19063), .ZN(n19062) );
  NAND2_X1 U15335 ( .A1(n12102), .A2(n12103), .ZN(n12104) );
  INV_X1 U15336 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19317) );
  NAND2_X1 U15337 ( .A1(n12109), .A2(n12105), .ZN(n12110) );
  INV_X1 U15338 ( .A(n12105), .ZN(n12108) );
  NAND2_X1 U15339 ( .A1(n19041), .A2(n19040), .ZN(n12107) );
  NAND2_X1 U15340 ( .A1(n12109), .A2(n12108), .ZN(n12106) );
  OAI211_X1 U15341 ( .C1(n12109), .C2(n12108), .A(n12107), .B(n12106), .ZN(
        n14572) );
  NAND2_X1 U15342 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n14572), .ZN(
        n14571) );
  NAND2_X1 U15343 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n19133) );
  NOR2_X1 U15344 ( .A1(n18797), .A2(n19133), .ZN(n19141) );
  AND2_X1 U15345 ( .A1(n19141), .A2(n17652), .ZN(n17651) );
  AND2_X1 U15346 ( .A1(n17651), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17631) );
  AND2_X1 U15347 ( .A1(n17631), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17566) );
  NAND3_X1 U15348 ( .A1(n17639), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12111) );
  XOR2_X1 U15349 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12111), .Z(
        n12174) );
  NOR2_X2 U15350 ( .A1(n18041), .A2(n20031), .ZN(n19121) );
  INV_X1 U15351 ( .A(n17566), .ZN(n17636) );
  INV_X1 U15352 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12113) );
  NOR2_X1 U15353 ( .A1(n17636), .A2(n12113), .ZN(n12114) );
  NAND2_X1 U15354 ( .A1(n18813), .A2(n12114), .ZN(n17609) );
  NOR2_X1 U15355 ( .A1(n17609), .A2(n12157), .ZN(n12115) );
  AOI211_X1 U15356 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n17609), .A(
        n12168), .B(n12115), .ZN(n12160) );
  INV_X1 U15357 ( .A(n12160), .ZN(n12132) );
  AND2_X2 U15358 ( .A1(n19119), .A2(n17608), .ZN(n18978) );
  NAND2_X1 U15359 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n19400) );
  NAND2_X1 U15360 ( .A1(n20016), .A2(n19400), .ZN(n20037) );
  INV_X1 U15361 ( .A(n20037), .ZN(n12116) );
  NAND2_X1 U15362 ( .A1(n12116), .A2(n20035), .ZN(n12117) );
  AND2_X1 U15363 ( .A1(n20035), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17601) );
  INV_X1 U15364 ( .A(n18868), .ZN(n13199) );
  INV_X1 U15365 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12123) );
  NAND2_X1 U15366 ( .A1(n19080), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19069) );
  NAND2_X1 U15367 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n19024) );
  NOR2_X1 U15368 ( .A1(n19024), .A2(n19025), .ZN(n18997) );
  NAND3_X1 U15369 ( .A1(n18997), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18954) );
  INV_X1 U15370 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18973) );
  NAND2_X1 U15371 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18926) );
  NAND2_X1 U15372 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18892) );
  NAND2_X1 U15373 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18849) );
  NAND2_X1 U15374 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18809) );
  NOR2_X2 U15375 ( .A1(n17600), .A2(n18809), .ZN(n18795) );
  NAND2_X1 U15376 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17568) );
  INV_X1 U15377 ( .A(n17568), .ZN(n12119) );
  INV_X1 U15378 ( .A(n17601), .ZN(n18969) );
  AND2_X1 U15379 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n12119), .ZN(
        n12120) );
  AND2_X1 U15380 ( .A1(n12118), .A2(n12120), .ZN(n12125) );
  INV_X1 U15381 ( .A(n12125), .ZN(n12121) );
  NAND2_X1 U15382 ( .A1(n18678), .A2(n20047), .ZN(n20034) );
  NOR3_X1 U15383 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n18037), .ZN(n19408) );
  NAND2_X1 U15384 ( .A1(n12121), .A2(n19801), .ZN(n17569) );
  OAI211_X1 U15385 ( .C1(n12122), .C2(n18969), .A(n19116), .B(n17569), .ZN(
        n17571) );
  AOI21_X1 U15386 ( .B1(n13199), .B2(n12123), .A(n17571), .ZN(n17556) );
  INV_X1 U15387 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n18081) );
  INV_X1 U15388 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19125) );
  NAND2_X1 U15389 ( .A1(n12124), .A2(n19636), .ZN(n18924) );
  NAND2_X1 U15390 ( .A1(n18924), .A2(n12125), .ZN(n17560) );
  XOR2_X1 U15391 ( .A(n18081), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n12126) );
  OR2_X1 U15392 ( .A1(n17560), .A2(n12126), .ZN(n12130) );
  NAND2_X1 U15393 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n19079) );
  NAND2_X1 U15394 ( .A1(n19116), .A2(n19079), .ZN(n19008) );
  NOR2_X1 U15395 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n20048) );
  NOR2_X1 U15396 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n12128) );
  NAND2_X1 U15397 ( .A1(n20048), .A2(n12128), .ZN(n19110) );
  INV_X1 U15398 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n20000) );
  NOR2_X1 U15399 ( .A1(n19349), .A2(n20000), .ZN(n12167) );
  AOI21_X1 U15400 ( .B1(n18977), .B2(n18406), .A(n12167), .ZN(n12129) );
  OAI211_X1 U15401 ( .C1(n17556), .C2(n18081), .A(n12130), .B(n12129), .ZN(
        n12131) );
  AOI21_X1 U15402 ( .B1(n12132), .B2(n18978), .A(n12131), .ZN(n12133) );
  OAI21_X1 U15403 ( .B1(n12174), .B2(n19112), .A(n12133), .ZN(n12134) );
  INV_X1 U15404 ( .A(n12134), .ZN(n12135) );
  NAND2_X1 U15405 ( .A1(n12136), .A2(n12135), .ZN(P3_U2799) );
  NAND2_X1 U15406 ( .A1(n19880), .A2(n12137), .ZN(n12145) );
  OAI21_X1 U15407 ( .B1(n12140), .B2(n12139), .A(n12138), .ZN(n12142) );
  NAND2_X1 U15408 ( .A1(n12153), .A2(n19878), .ZN(n12143) );
  AND2_X1 U15409 ( .A1(n13366), .A2(n12143), .ZN(n12144) );
  AOI21_X1 U15410 ( .B1(n12145), .B2(n12144), .A(n19914), .ZN(n12155) );
  NAND2_X1 U15411 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n20040) );
  INV_X1 U15412 ( .A(n19426), .ZN(n12150) );
  INV_X1 U15413 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19930) );
  NAND2_X1 U15414 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19930), .ZN(n20026) );
  INV_X1 U15415 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19943) );
  NOR2_X1 U15416 ( .A1(n20026), .A2(n19943), .ZN(n19942) );
  NOR2_X1 U15417 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n19928) );
  NOR3_X1 U15418 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19942), .A3(n19928), 
        .ZN(n20030) );
  INV_X1 U15419 ( .A(n12148), .ZN(n12149) );
  AOI211_X1 U15420 ( .C1(n19420), .C2(n12150), .A(n20030), .B(n12149), .ZN(
        n12151) );
  NOR2_X1 U15421 ( .A1(n20032), .A2(n12151), .ZN(n18038) );
  NAND2_X1 U15422 ( .A1(n18742), .A2(n18038), .ZN(n12152) );
  NOR2_X1 U15423 ( .A1(n12153), .A2(n12152), .ZN(n12154) );
  NAND2_X1 U15424 ( .A1(n12156), .A2(n19297), .ZN(n12177) );
  OR2_X1 U15425 ( .A1(n19387), .A2(n19399), .ZN(n19377) );
  INV_X1 U15426 ( .A(n19263), .ZN(n19322) );
  AOI21_X1 U15427 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19313) );
  INV_X1 U15428 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19362) );
  NOR3_X1 U15429 ( .A1(n19362), .A2(n9976), .A3(n19356), .ZN(n19315) );
  NAND2_X1 U15430 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n19315), .ZN(
        n19331) );
  NOR2_X1 U15431 ( .A1(n19317), .A2(n19331), .ZN(n19320) );
  NAND2_X1 U15432 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n19320), .ZN(
        n19196) );
  NOR2_X1 U15433 ( .A1(n19313), .A2(n19196), .ZN(n19218) );
  NAND2_X1 U15434 ( .A1(n10157), .A2(n19218), .ZN(n19156) );
  AOI21_X1 U15435 ( .B1(n19283), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n19160), .ZN(n19378) );
  NAND2_X1 U15436 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19314) );
  NOR2_X1 U15437 ( .A1(n19196), .A2(n19314), .ZN(n19219) );
  NAND2_X1 U15438 ( .A1(n10157), .A2(n19219), .ZN(n19198) );
  OAI22_X1 U15439 ( .A1(n19382), .A2(n19156), .B1(n19378), .B2(n19198), .ZN(
        n19139) );
  INV_X1 U15440 ( .A(n12157), .ZN(n12158) );
  NAND4_X1 U15441 ( .A1(n19139), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n17566), .A4(n12158), .ZN(n12159) );
  OAI21_X1 U15442 ( .B1(n12160), .B2(n19322), .A(n12159), .ZN(n12172) );
  NAND2_X1 U15443 ( .A1(n19318), .A2(n19341), .ZN(n19361) );
  INV_X1 U15444 ( .A(n19361), .ZN(n12169) );
  INV_X1 U15445 ( .A(n19198), .ZN(n12161) );
  INV_X1 U15446 ( .A(n19160), .ZN(n19220) );
  AOI21_X1 U15447 ( .B1(n17651), .B2(n12161), .A(n19220), .ZN(n12165) );
  INV_X1 U15448 ( .A(n17651), .ZN(n17584) );
  NOR2_X1 U15449 ( .A1(n19156), .A2(n17584), .ZN(n12162) );
  NOR2_X1 U15450 ( .A1(n19382), .A2(n12162), .ZN(n17655) );
  NAND2_X1 U15451 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n19219), .ZN(
        n19282) );
  NOR2_X1 U15452 ( .A1(n12163), .A2(n19282), .ZN(n19217) );
  AOI21_X1 U15453 ( .B1(n17631), .B2(n19217), .A(n19306), .ZN(n12164) );
  NOR3_X1 U15454 ( .A1(n12165), .A2(n17655), .A3(n12164), .ZN(n17623) );
  NAND2_X1 U15455 ( .A1(n19399), .A2(n19110), .ZN(n19360) );
  OAI21_X1 U15456 ( .B1(n17623), .B2(n19399), .A(n19360), .ZN(n12166) );
  AOI21_X1 U15457 ( .B1(n12169), .B2(n17554), .A(n12166), .ZN(n17612) );
  AOI21_X1 U15458 ( .B1(n12169), .B2(n12168), .A(n12167), .ZN(n12170) );
  OAI21_X1 U15459 ( .B1(n17612), .B2(n13381), .A(n12170), .ZN(n12171) );
  AOI21_X1 U15460 ( .B1(n12172), .B2(n19341), .A(n12171), .ZN(n12173) );
  OAI21_X1 U15461 ( .B1(n12174), .B2(n19377), .A(n12173), .ZN(n12175) );
  INV_X1 U15462 ( .A(n12175), .ZN(n12176) );
  NAND2_X1 U15463 ( .A1(n12177), .A2(n12176), .ZN(P3_U2831) );
  NOR2_X1 U15464 ( .A1(n12178), .A2(n9769), .ZN(n12179) );
  INV_X1 U15465 ( .A(n9770), .ZN(n14903) );
  AOI21_X1 U15466 ( .B1(n14903), .B2(n10176), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12180) );
  NAND2_X1 U15467 ( .A1(n20167), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n16902) );
  OAI21_X1 U15468 ( .B1(n12181), .B2(n12180), .A(n16902), .ZN(n12182) );
  AOI21_X1 U15469 ( .B1(n16773), .B2(n17461), .A(n12182), .ZN(n12183) );
  OAI21_X1 U15470 ( .B1(n16906), .B2(n17429), .A(n12183), .ZN(n12184) );
  OAI211_X1 U15471 ( .C1(n16910), .C2(n17458), .A(n12186), .B(n12185), .ZN(
        P2_U3016) );
  AND2_X1 U15472 ( .A1(n14914), .A2(n14913), .ZN(n12188) );
  INV_X1 U15473 ( .A(n20966), .ZN(n20963) );
  OR2_X1 U15474 ( .A1(n15442), .A2(n20963), .ZN(n13217) );
  NOR2_X1 U15475 ( .A1(n13217), .A2(n14388), .ZN(n12191) );
  INV_X1 U15476 ( .A(n12194), .ZN(n12497) );
  AND2_X1 U15477 ( .A1(n12243), .A2(n13780), .ZN(n12195) );
  NAND2_X1 U15478 ( .A1(n16897), .A2(n12195), .ZN(n13873) );
  INV_X1 U15479 ( .A(n13873), .ZN(n12206) );
  NOR4_X1 U15480 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12199) );
  NOR4_X1 U15481 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12198) );
  NOR4_X1 U15482 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12197) );
  NOR4_X1 U15483 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12196) );
  AND4_X1 U15484 ( .A1(n12199), .A2(n12198), .A3(n12197), .A4(n12196), .ZN(
        n12204) );
  NOR4_X1 U15485 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12202) );
  NOR4_X1 U15486 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12201) );
  NOR4_X1 U15487 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12200) );
  INV_X1 U15488 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20852) );
  AND4_X1 U15489 ( .A1(n12202), .A2(n12201), .A3(n12200), .A4(n20852), .ZN(
        n12203) );
  NAND2_X1 U15490 ( .A1(n12204), .A2(n12203), .ZN(n12205) );
  AND2_X2 U15491 ( .A1(n12205), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n17490)
         );
  INV_X1 U15492 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n12212) );
  NOR2_X2 U15493 ( .A1(n13873), .A2(n17488), .ZN(n16873) );
  NAND2_X1 U15494 ( .A1(n16873), .A2(BUF1_REG_29__SCAN_IN), .ZN(n12211) );
  NAND2_X1 U15495 ( .A1(n11473), .A2(n13780), .ZN(n12207) );
  INV_X1 U15496 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n12209) );
  NAND2_X1 U15497 ( .A1(n17490), .A2(BUF1_REG_13__SCAN_IN), .ZN(n12208) );
  OAI21_X1 U15498 ( .B1(n17490), .B2(n12209), .A(n12208), .ZN(n14434) );
  AOI22_X1 U15499 ( .A1(n16875), .A2(n14434), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n20226), .ZN(n12210) );
  OAI211_X1 U15500 ( .C1(n16878), .C2(n12212), .A(n12211), .B(n12210), .ZN(
        n12213) );
  INV_X1 U15501 ( .A(n12213), .ZN(n12496) );
  INV_X1 U15502 ( .A(n12239), .ZN(n12225) );
  NAND2_X1 U15503 ( .A1(n17446), .A2(n12225), .ZN(n12219) );
  NAND2_X1 U15504 ( .A1(n12243), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12215) );
  AND2_X1 U15505 ( .A1(n20504), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12216) );
  NAND2_X1 U15506 ( .A1(n12216), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20814) );
  INV_X1 U15507 ( .A(n12216), .ZN(n12235) );
  NAND2_X1 U15508 ( .A1(n12235), .A2(n20920), .ZN(n12217) );
  AND3_X1 U15509 ( .A1(n20814), .A2(n20958), .A3(n12217), .ZN(n20651) );
  AOI21_X1 U15510 ( .B1(n12237), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n20651), .ZN(n12218) );
  NAND2_X1 U15511 ( .A1(n12219), .A2(n12218), .ZN(n12245) );
  NOR2_X1 U15512 ( .A1(n12243), .A2(n11573), .ZN(n12220) );
  NAND2_X1 U15513 ( .A1(n12245), .A2(n12221), .ZN(n16892) );
  OAI21_X1 U15514 ( .B1(n12245), .B2(n12221), .A(n16892), .ZN(n12222) );
  NAND2_X1 U15515 ( .A1(n20938), .A2(n20947), .ZN(n12223) );
  INV_X1 U15516 ( .A(n20504), .ZN(n20387) );
  AND2_X1 U15517 ( .A1(n12223), .A2(n20387), .ZN(n20419) );
  AND2_X1 U15518 ( .A1(n20419), .A2(n20958), .ZN(n20359) );
  AOI21_X1 U15519 ( .B1(n12237), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n20359), .ZN(n12224) );
  AOI22_X1 U15520 ( .A1(n12237), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20958), .B2(n20947), .ZN(n12226) );
  INV_X1 U15521 ( .A(n13905), .ZN(n12228) );
  INV_X1 U15522 ( .A(n12229), .ZN(n12232) );
  INV_X1 U15523 ( .A(n12230), .ZN(n12231) );
  NAND2_X1 U15524 ( .A1(n12232), .A2(n12231), .ZN(n12233) );
  NOR2_X1 U15525 ( .A1(n13895), .A2(n13774), .ZN(n12241) );
  INV_X1 U15526 ( .A(n20958), .ZN(n20563) );
  NAND2_X1 U15527 ( .A1(n20387), .A2(n20927), .ZN(n12234) );
  NAND2_X1 U15528 ( .A1(n12235), .A2(n12234), .ZN(n20418) );
  NOR2_X1 U15529 ( .A1(n20563), .A2(n20418), .ZN(n12236) );
  AOI21_X1 U15530 ( .B1(n12237), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12236), .ZN(n12238) );
  NAND2_X1 U15531 ( .A1(n12245), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12246) );
  INV_X1 U15532 ( .A(n12247), .ZN(n14491) );
  NAND2_X1 U15533 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14251) );
  NAND2_X1 U15534 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12248) );
  NOR2_X1 U15535 ( .A1(n14251), .A2(n12248), .ZN(n12250) );
  INV_X1 U15536 ( .A(n12252), .ZN(n14706) );
  INV_X1 U15537 ( .A(n12253), .ZN(n16758) );
  AOI22_X1 U15538 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12257) );
  AOI22_X1 U15539 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12256) );
  AOI22_X1 U15540 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U15541 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10921), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12254) );
  NAND4_X1 U15542 ( .A1(n12257), .A2(n12256), .A3(n12255), .A4(n12254), .ZN(
        n12263) );
  AOI22_X1 U15543 ( .A1(n10849), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U15544 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12260) );
  AOI22_X1 U15545 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12259) );
  AOI22_X1 U15546 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12258) );
  NAND4_X1 U15547 ( .A1(n12261), .A2(n12260), .A3(n12259), .A4(n12258), .ZN(
        n12262) );
  OR2_X1 U15548 ( .A1(n12263), .A2(n12262), .ZN(n16749) );
  AOI22_X1 U15549 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U15550 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U15551 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15552 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10921), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12264) );
  NAND4_X1 U15553 ( .A1(n12267), .A2(n12266), .A3(n12265), .A4(n12264), .ZN(
        n12273) );
  AOI22_X1 U15554 ( .A1(n10849), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12271) );
  AOI22_X1 U15555 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U15556 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15557 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12268) );
  NAND4_X1 U15558 ( .A1(n12271), .A2(n12270), .A3(n12269), .A4(n12268), .ZN(
        n12272) );
  OR2_X1 U15559 ( .A1(n12273), .A2(n12272), .ZN(n16745) );
  AOI22_X1 U15560 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U15561 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U15562 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U15563 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10921), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12274) );
  NAND4_X1 U15564 ( .A1(n12277), .A2(n12276), .A3(n12275), .A4(n12274), .ZN(
        n12283) );
  AOI22_X1 U15565 ( .A1(n10849), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12281) );
  AOI22_X1 U15566 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12280) );
  AOI22_X1 U15567 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12279) );
  AOI22_X1 U15568 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12278) );
  NAND4_X1 U15569 ( .A1(n12281), .A2(n12280), .A3(n12279), .A4(n12278), .ZN(
        n12282) );
  NOR2_X1 U15570 ( .A1(n12283), .A2(n12282), .ZN(n16741) );
  INV_X1 U15571 ( .A(n16741), .ZN(n12284) );
  AOI22_X1 U15572 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U15573 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U15574 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U15575 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10921), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12285) );
  NAND4_X1 U15576 ( .A1(n12288), .A2(n12287), .A3(n12286), .A4(n12285), .ZN(
        n12294) );
  AOI22_X1 U15577 ( .A1(n10849), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U15578 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U15579 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12290) );
  AOI22_X1 U15580 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12289) );
  NAND4_X1 U15581 ( .A1(n12292), .A2(n12291), .A3(n12290), .A4(n12289), .ZN(
        n12293) );
  NOR2_X1 U15582 ( .A1(n12294), .A2(n12293), .ZN(n16734) );
  AOI22_X1 U15583 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15584 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15585 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12296) );
  AOI22_X1 U15586 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10921), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12295) );
  NAND4_X1 U15587 ( .A1(n12298), .A2(n12297), .A3(n12296), .A4(n12295), .ZN(
        n12304) );
  AOI22_X1 U15588 ( .A1(n10849), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12302) );
  AOI22_X1 U15589 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12301) );
  AOI22_X1 U15590 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12300) );
  AOI22_X1 U15591 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12299) );
  NAND4_X1 U15592 ( .A1(n12302), .A2(n12301), .A3(n12300), .A4(n12299), .ZN(
        n12303) );
  OR2_X1 U15593 ( .A1(n12304), .A2(n12303), .ZN(n16724) );
  AOI22_X1 U15594 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U15595 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12307) );
  AOI22_X1 U15596 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15597 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10921), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12305) );
  NAND4_X1 U15598 ( .A1(n12308), .A2(n12307), .A3(n12306), .A4(n12305), .ZN(
        n12315) );
  AOI22_X1 U15599 ( .A1(n10849), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U15600 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15601 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U15602 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12310) );
  NAND4_X1 U15603 ( .A1(n12313), .A2(n12312), .A3(n12311), .A4(n12310), .ZN(
        n12314) );
  OR2_X1 U15604 ( .A1(n12315), .A2(n12314), .ZN(n16728) );
  INV_X1 U15605 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n20333) );
  AOI22_X1 U15606 ( .A1(n12329), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16658), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12328) );
  NAND2_X1 U15607 ( .A1(n16662), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12323) );
  NAND2_X1 U15608 ( .A1(n16664), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12322) );
  INV_X1 U15609 ( .A(n12318), .ZN(n14369) );
  INV_X1 U15610 ( .A(n14369), .ZN(n12330) );
  NAND2_X1 U15611 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12321) );
  NAND2_X1 U15612 ( .A1(n16663), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12320) );
  AND4_X1 U15613 ( .A1(n12323), .A2(n12322), .A3(n12321), .A4(n12320), .ZN(
        n12327) );
  AOI22_X1 U15614 ( .A1(n16656), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16657), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12326) );
  XNOR2_X1 U15615 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16653) );
  NAND4_X1 U15616 ( .A1(n12328), .A2(n12327), .A3(n12326), .A4(n16653), .ZN(
        n12339) );
  AOI22_X1 U15617 ( .A1(n12329), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16656), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12337) );
  NAND2_X1 U15618 ( .A1(n16662), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12334) );
  NAND2_X1 U15619 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12333) );
  NAND2_X1 U15620 ( .A1(n16664), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12332) );
  INV_X1 U15621 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n20760) );
  NAND2_X1 U15622 ( .A1(n16663), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12331) );
  AND4_X1 U15623 ( .A1(n12334), .A2(n12333), .A3(n12332), .A4(n12331), .ZN(
        n12336) );
  INV_X1 U15624 ( .A(n16653), .ZN(n16660) );
  AOI22_X1 U15625 ( .A1(n16658), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16657), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12335) );
  NAND4_X1 U15626 ( .A1(n12337), .A2(n12336), .A3(n16660), .A4(n12335), .ZN(
        n12338) );
  AND2_X1 U15627 ( .A1(n12339), .A2(n12338), .ZN(n12363) );
  NAND2_X1 U15628 ( .A1(n16694), .A2(n12363), .ZN(n12366) );
  AOI22_X1 U15629 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10802), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12344) );
  AOI22_X1 U15630 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12340), .B1(
        n10921), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12343) );
  AOI22_X1 U15631 ( .A1(n10619), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12342) );
  AOI22_X1 U15632 ( .A1(n10803), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10804), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12341) );
  NAND4_X1 U15633 ( .A1(n12344), .A2(n12343), .A3(n12342), .A4(n12341), .ZN(
        n12350) );
  AOI22_X1 U15634 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n10926), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12348) );
  AOI22_X1 U15635 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12355), .B1(
        n12309), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U15636 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10624), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U15637 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n10797), .B1(
        n12356), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12345) );
  NAND4_X1 U15638 ( .A1(n12348), .A2(n12347), .A3(n12346), .A4(n12345), .ZN(
        n12349) );
  OR2_X1 U15639 ( .A1(n12350), .A2(n12349), .ZN(n12387) );
  XNOR2_X1 U15640 ( .A(n12366), .B(n12387), .ZN(n16712) );
  AOI22_X1 U15641 ( .A1(n10617), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10619), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12354) );
  AOI22_X1 U15642 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12353) );
  AOI22_X1 U15643 ( .A1(n10804), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10618), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12352) );
  AOI22_X1 U15644 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10921), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12351) );
  NAND4_X1 U15645 ( .A1(n12354), .A2(n12353), .A3(n12352), .A4(n12351), .ZN(
        n12362) );
  AOI22_X1 U15646 ( .A1(n10849), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10926), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15647 ( .A1(n12309), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10625), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15648 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10624), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U15649 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10797), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12357) );
  NAND4_X1 U15650 ( .A1(n12360), .A2(n12359), .A3(n12358), .A4(n12357), .ZN(
        n12361) );
  OR2_X1 U15651 ( .A1(n12362), .A2(n12361), .ZN(n16717) );
  NAND2_X1 U15652 ( .A1(n16712), .A2(n16717), .ZN(n12365) );
  INV_X1 U15653 ( .A(n12363), .ZN(n12386) );
  NOR2_X1 U15654 ( .A1(n16694), .A2(n12386), .ZN(n16711) );
  NAND2_X1 U15655 ( .A1(n16712), .A2(n16711), .ZN(n12364) );
  INV_X1 U15656 ( .A(n12366), .ZN(n12367) );
  NAND2_X1 U15657 ( .A1(n12367), .A2(n12387), .ZN(n12385) );
  AOI22_X1 U15658 ( .A1(n12329), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n16656), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12374) );
  NAND2_X1 U15659 ( .A1(n16662), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12371) );
  NAND2_X1 U15660 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12370) );
  NAND2_X1 U15661 ( .A1(n16663), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12369) );
  NAND2_X1 U15662 ( .A1(n16664), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12368) );
  AND4_X1 U15663 ( .A1(n12371), .A2(n12370), .A3(n12369), .A4(n12368), .ZN(
        n12373) );
  AOI22_X1 U15664 ( .A1(n16658), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n16657), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12372) );
  NAND4_X1 U15665 ( .A1(n12374), .A2(n12373), .A3(n12372), .A4(n16653), .ZN(
        n12384) );
  AOI22_X1 U15666 ( .A1(n16658), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16656), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12382) );
  NAND2_X1 U15667 ( .A1(n16662), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12378) );
  NAND2_X1 U15668 ( .A1(n16664), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12377) );
  NAND2_X1 U15669 ( .A1(n16663), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12376) );
  NAND2_X1 U15670 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12375) );
  AND4_X1 U15671 ( .A1(n12378), .A2(n12377), .A3(n12376), .A4(n12375), .ZN(
        n12381) );
  AOI22_X1 U15672 ( .A1(n12329), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n16657), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12380) );
  NAND4_X1 U15673 ( .A1(n12382), .A2(n12381), .A3(n16660), .A4(n12380), .ZN(
        n12383) );
  NAND2_X1 U15674 ( .A1(n12384), .A2(n12383), .ZN(n12390) );
  NAND2_X1 U15675 ( .A1(n12385), .A2(n12390), .ZN(n12389) );
  NOR2_X1 U15676 ( .A1(n12390), .A2(n12386), .ZN(n12388) );
  NAND2_X1 U15677 ( .A1(n12388), .A2(n12387), .ZN(n12394) );
  NAND2_X1 U15678 ( .A1(n12389), .A2(n12394), .ZN(n12393) );
  INV_X1 U15679 ( .A(n12390), .ZN(n12391) );
  NAND2_X1 U15680 ( .A1(n13223), .A2(n12391), .ZN(n12392) );
  NAND2_X1 U15681 ( .A1(n12393), .A2(n12392), .ZN(n16706) );
  INV_X1 U15682 ( .A(n12394), .ZN(n12411) );
  INV_X1 U15683 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n20338) );
  AOI22_X1 U15684 ( .A1(n16658), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16656), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12401) );
  NAND2_X1 U15685 ( .A1(n16662), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n12398) );
  NAND2_X1 U15686 ( .A1(n16664), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12397) );
  NAND2_X1 U15687 ( .A1(n16663), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12396) );
  INV_X1 U15688 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14212) );
  NAND2_X1 U15689 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n12395) );
  AND4_X1 U15690 ( .A1(n12398), .A2(n12397), .A3(n12396), .A4(n12395), .ZN(
        n12400) );
  AOI22_X1 U15691 ( .A1(n12329), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16657), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12399) );
  NAND4_X1 U15692 ( .A1(n12401), .A2(n12400), .A3(n12399), .A4(n16653), .ZN(
        n12410) );
  AOI22_X1 U15693 ( .A1(n16658), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16656), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12408) );
  NAND2_X1 U15694 ( .A1(n16662), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n12405) );
  NAND2_X1 U15695 ( .A1(n16664), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12404) );
  NAND2_X1 U15696 ( .A1(n16663), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12403) );
  NAND2_X1 U15697 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12402) );
  AND4_X1 U15698 ( .A1(n12405), .A2(n12404), .A3(n12403), .A4(n12402), .ZN(
        n12407) );
  AOI22_X1 U15699 ( .A1(n12329), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16657), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12406) );
  NAND4_X1 U15700 ( .A1(n12408), .A2(n12407), .A3(n16660), .A4(n12406), .ZN(
        n12409) );
  AND2_X1 U15701 ( .A1(n12410), .A2(n12409), .ZN(n12412) );
  NAND2_X1 U15702 ( .A1(n12411), .A2(n12412), .ZN(n12436) );
  OAI211_X1 U15703 ( .C1(n12411), .C2(n12412), .A(n14249), .B(n12436), .ZN(
        n12431) );
  NAND2_X1 U15704 ( .A1(n13223), .A2(n12412), .ZN(n16702) );
  INV_X1 U15705 ( .A(n16702), .ZN(n12430) );
  AOI22_X1 U15706 ( .A1(n12329), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16656), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12419) );
  NAND2_X1 U15707 ( .A1(n16662), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12416) );
  NAND2_X1 U15708 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12415) );
  NAND2_X1 U15709 ( .A1(n16664), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12414) );
  NAND2_X1 U15710 ( .A1(n16663), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12413) );
  AND4_X1 U15711 ( .A1(n12416), .A2(n12415), .A3(n12414), .A4(n12413), .ZN(
        n12418) );
  AOI22_X1 U15712 ( .A1(n16658), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16657), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12417) );
  NAND4_X1 U15713 ( .A1(n12419), .A2(n12418), .A3(n12417), .A4(n16653), .ZN(
        n12428) );
  AOI22_X1 U15714 ( .A1(n12329), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16656), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12426) );
  NAND2_X1 U15715 ( .A1(n16662), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12423) );
  NAND2_X1 U15716 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12422) );
  NAND2_X1 U15717 ( .A1(n16664), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12421) );
  NAND2_X1 U15718 ( .A1(n16663), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12420) );
  AND4_X1 U15719 ( .A1(n12423), .A2(n12422), .A3(n12421), .A4(n12420), .ZN(
        n12425) );
  AOI22_X1 U15720 ( .A1(n16658), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16657), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12424) );
  NAND4_X1 U15721 ( .A1(n12426), .A2(n12425), .A3(n16660), .A4(n12424), .ZN(
        n12427) );
  NAND2_X1 U15722 ( .A1(n12428), .A2(n12427), .ZN(n16693) );
  INV_X1 U15723 ( .A(n16693), .ZN(n12429) );
  NAND2_X1 U15724 ( .A1(n12430), .A2(n12429), .ZN(n12435) );
  XNOR2_X1 U15725 ( .A(n12436), .B(n16693), .ZN(n12433) );
  INV_X1 U15726 ( .A(n14249), .ZN(n12432) );
  NOR2_X1 U15727 ( .A1(n12433), .A2(n12432), .ZN(n16696) );
  NAND2_X1 U15728 ( .A1(n16692), .A2(n16696), .ZN(n12434) );
  INV_X1 U15729 ( .A(n12457), .ZN(n12454) );
  NOR2_X1 U15730 ( .A1(n12436), .A2(n16693), .ZN(n12453) );
  AOI22_X1 U15731 ( .A1(n12329), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16656), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12443) );
  NAND2_X1 U15732 ( .A1(n16662), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12440) );
  NAND2_X1 U15733 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12439) );
  NAND2_X1 U15734 ( .A1(n16664), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12438) );
  NAND2_X1 U15735 ( .A1(n16663), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12437) );
  AND4_X1 U15736 ( .A1(n12440), .A2(n12439), .A3(n12438), .A4(n12437), .ZN(
        n12442) );
  AOI22_X1 U15737 ( .A1(n16658), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16657), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12441) );
  NAND4_X1 U15738 ( .A1(n12443), .A2(n12442), .A3(n12441), .A4(n16653), .ZN(
        n12452) );
  AOI22_X1 U15739 ( .A1(n12329), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16656), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12450) );
  NAND2_X1 U15740 ( .A1(n16662), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12447) );
  NAND2_X1 U15741 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12446) );
  NAND2_X1 U15742 ( .A1(n16664), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12445) );
  NAND2_X1 U15743 ( .A1(n16663), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12444) );
  AND4_X1 U15744 ( .A1(n12447), .A2(n12446), .A3(n12445), .A4(n12444), .ZN(
        n12449) );
  AOI22_X1 U15745 ( .A1(n16658), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16657), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12448) );
  NAND4_X1 U15746 ( .A1(n12450), .A2(n12449), .A3(n16660), .A4(n12448), .ZN(
        n12451) );
  AND2_X1 U15747 ( .A1(n12452), .A2(n12451), .ZN(n12459) );
  NAND2_X1 U15748 ( .A1(n12453), .A2(n12459), .ZN(n16679) );
  OAI211_X1 U15749 ( .C1(n12453), .C2(n12459), .A(n16679), .B(n14249), .ZN(
        n12455) );
  INV_X1 U15750 ( .A(n12455), .ZN(n12456) );
  INV_X1 U15751 ( .A(n12459), .ZN(n12460) );
  NOR2_X1 U15752 ( .A1(n16694), .A2(n12460), .ZN(n16686) );
  AOI22_X1 U15753 ( .A1(n12329), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16656), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12468) );
  NAND2_X1 U15754 ( .A1(n16662), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12465) );
  NAND2_X1 U15755 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12464) );
  NAND2_X1 U15756 ( .A1(n16664), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12463) );
  NAND2_X1 U15757 ( .A1(n16663), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12462) );
  AND4_X1 U15758 ( .A1(n12465), .A2(n12464), .A3(n12463), .A4(n12462), .ZN(
        n12467) );
  AOI22_X1 U15759 ( .A1(n16658), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n16657), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12466) );
  NAND4_X1 U15760 ( .A1(n12468), .A2(n12467), .A3(n12466), .A4(n16653), .ZN(
        n12478) );
  AOI22_X1 U15761 ( .A1(n12329), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16656), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12476) );
  NAND2_X1 U15762 ( .A1(n16662), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12473) );
  NAND2_X1 U15763 ( .A1(n12330), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12472) );
  NAND2_X1 U15764 ( .A1(n16664), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12471) );
  NAND2_X1 U15765 ( .A1(n16663), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12470) );
  AND4_X1 U15766 ( .A1(n12473), .A2(n12472), .A3(n12471), .A4(n12470), .ZN(
        n12475) );
  AOI22_X1 U15767 ( .A1(n16658), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16657), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12474) );
  NAND4_X1 U15768 ( .A1(n12476), .A2(n12475), .A3(n16660), .A4(n12474), .ZN(
        n12477) );
  NAND2_X1 U15769 ( .A1(n12478), .A2(n12477), .ZN(n16681) );
  AOI22_X1 U15770 ( .A1(n16662), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16664), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12480) );
  INV_X1 U15771 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14056) );
  AOI22_X1 U15772 ( .A1(n16663), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12330), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12479) );
  AND2_X1 U15773 ( .A1(n12480), .A2(n12479), .ZN(n12483) );
  AOI22_X1 U15774 ( .A1(n12329), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16657), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U15775 ( .A1(n16658), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16656), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12481) );
  NAND4_X1 U15776 ( .A1(n12483), .A2(n12482), .A3(n12481), .A4(n16653), .ZN(
        n12490) );
  AOI22_X1 U15777 ( .A1(n16662), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12330), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12485) );
  INV_X1 U15778 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14213) );
  AOI22_X1 U15779 ( .A1(n16663), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16664), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12484) );
  AND2_X1 U15780 ( .A1(n12485), .A2(n12484), .ZN(n12488) );
  AOI22_X1 U15781 ( .A1(n12329), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16658), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12487) );
  INV_X1 U15782 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n20745) );
  AOI22_X1 U15783 ( .A1(n16656), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16657), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12486) );
  NAND4_X1 U15784 ( .A1(n12488), .A2(n16660), .A3(n12487), .A4(n12486), .ZN(
        n12489) );
  NAND2_X1 U15785 ( .A1(n12490), .A2(n12489), .ZN(n12492) );
  OR3_X1 U15786 ( .A1(n16679), .A2(n13223), .A3(n16681), .ZN(n12491) );
  AOI21_X1 U15787 ( .B1(n12492), .B2(n12491), .A(n16650), .ZN(n12493) );
  NAND2_X1 U15788 ( .A1(n16897), .A2(n12494), .ZN(n16883) );
  AOI21_X1 U15789 ( .B1(n16400), .B2(n16914), .A(n20177), .ZN(n12498) );
  INV_X1 U15790 ( .A(n12498), .ZN(n12499) );
  NAND2_X1 U15791 ( .A1(n12500), .A2(n10328), .ZN(n12509) );
  AOI22_X1 U15792 ( .A1(n20150), .A2(P2_REIP_REG_29__SCAN_IN), .B1(n20169), 
        .B2(P2_EBX_REG_29__SCAN_IN), .ZN(n12501) );
  OAI21_X1 U15793 ( .B1(n16912), .B2(n20145), .A(n12501), .ZN(n12503) );
  NOR2_X1 U15794 ( .A1(n14909), .A2(n20171), .ZN(n12502) );
  AOI21_X1 U15795 ( .B1(n12506), .B2(n12505), .A(n11640), .ZN(n14907) );
  INV_X1 U15796 ( .A(n14907), .ZN(n16916) );
  NAND3_X1 U15797 ( .A1(n12509), .A2(n12508), .A3(n12507), .ZN(P2_U2826) );
  NOR2_X4 U15798 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12519) );
  AND2_X4 U15799 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12518) );
  AOI22_X1 U15800 ( .A1(n15302), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12515) );
  AOI22_X1 U15801 ( .A1(n12687), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15283), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12514) );
  NOR2_X4 U15802 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14304) );
  AOI22_X1 U15803 ( .A1(n12696), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12512) );
  INV_X1 U15804 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12516) );
  AND2_X2 U15805 ( .A1(n12516), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12520) );
  AOI22_X1 U15806 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12589), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12524) );
  AOI22_X1 U15807 ( .A1(n12536), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12523) );
  AND2_X2 U15808 ( .A1(n12519), .A2(n12518), .ZN(n12558) );
  AOI22_X1 U15809 ( .A1(n12717), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12558), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12522) );
  AND2_X2 U15810 ( .A1(n14290), .A2(n14304), .ZN(n12612) );
  AOI22_X1 U15811 ( .A1(n12611), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12521) );
  AOI22_X1 U15813 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12536), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12530) );
  AOI22_X1 U15814 ( .A1(n12687), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15283), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12529) );
  AOI22_X1 U15815 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12605), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12528) );
  AOI22_X1 U15816 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12527) );
  AOI22_X1 U15817 ( .A1(n12611), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12534) );
  AOI22_X1 U15818 ( .A1(n12617), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12589), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12533) );
  AOI22_X1 U15819 ( .A1(n9699), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12532) );
  AOI22_X1 U15820 ( .A1(n12717), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12558), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12531) );
  AND4_X2 U15821 ( .A1(n12534), .A2(n12533), .A3(n12532), .A4(n12531), .ZN(
        n12535) );
  AOI22_X1 U15822 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12589), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12540) );
  AOI22_X1 U15823 ( .A1(n12717), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12558), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12539) );
  AOI22_X1 U15824 ( .A1(n12611), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12538) );
  AOI22_X1 U15825 ( .A1(n12536), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12537) );
  AOI22_X1 U15826 ( .A1(n9699), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n9704), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12544) );
  AOI22_X1 U15827 ( .A1(n12687), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15283), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12543) );
  AOI22_X1 U15828 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12605), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12542) );
  AOI22_X1 U15829 ( .A1(n12696), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12541) );
  NAND2_X1 U15830 ( .A1(n12611), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12549) );
  NAND2_X1 U15831 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12548) );
  NAND2_X1 U15832 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12547) );
  NAND2_X1 U15833 ( .A1(n12589), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12546) );
  NAND2_X1 U15834 ( .A1(n9699), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12553) );
  NAND2_X1 U15835 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12552) );
  NAND2_X1 U15836 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12551) );
  NAND2_X1 U15837 ( .A1(n12696), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12550) );
  NAND2_X1 U15838 ( .A1(n12687), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12557) );
  NAND2_X1 U15839 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12556) );
  NAND2_X1 U15840 ( .A1(n15283), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12555) );
  NAND2_X1 U15841 ( .A1(n12594), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12554) );
  NAND2_X1 U15842 ( .A1(n12536), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12562) );
  NAND2_X1 U15843 ( .A1(n12617), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12561) );
  NAND2_X1 U15844 ( .A1(n12717), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12560) );
  NAND2_X1 U15845 ( .A1(n12558), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12559) );
  AND4_X2 U15846 ( .A1(n12562), .A2(n12561), .A3(n12560), .A4(n12559), .ZN(
        n12563) );
  AND4_X4 U15847 ( .A1(n12566), .A2(n12565), .A3(n12564), .A4(n12563), .ZN(
        n12695) );
  INV_X2 U15848 ( .A(n12695), .ZN(n12636) );
  AOI22_X1 U15849 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15283), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12570) );
  AOI22_X1 U15850 ( .A1(n9707), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12569) );
  AOI22_X1 U15851 ( .A1(n12589), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12717), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12568) );
  AOI22_X1 U15852 ( .A1(n12687), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12567) );
  NAND4_X1 U15853 ( .A1(n12570), .A2(n12569), .A3(n12568), .A4(n12567), .ZN(
        n12576) );
  AOI22_X1 U15854 ( .A1(n12536), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12611), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12574) );
  AOI22_X1 U15855 ( .A1(n9699), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12605), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12573) );
  AOI22_X1 U15856 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12572) );
  AOI22_X1 U15857 ( .A1(n12617), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12558), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12571) );
  NAND4_X1 U15858 ( .A1(n12574), .A2(n12573), .A3(n12572), .A4(n12571), .ZN(
        n12575) );
  AOI22_X1 U15859 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12589), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12580) );
  AOI22_X1 U15860 ( .A1(n12611), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12579) );
  AOI22_X1 U15861 ( .A1(n12717), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12558), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12578) );
  AOI22_X1 U15862 ( .A1(n12536), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12577) );
  AOI22_X1 U15863 ( .A1(n9699), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U15864 ( .A1(n12687), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15283), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12584) );
  AOI22_X1 U15865 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12605), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12583) );
  AOI22_X1 U15866 ( .A1(n12696), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12582) );
  NAND2_X1 U15867 ( .A1(n12586), .A2(n10565), .ZN(n12626) );
  AOI22_X1 U15868 ( .A1(n12611), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12593) );
  AOI22_X1 U15869 ( .A1(n12536), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12592) );
  AOI22_X1 U15870 ( .A1(n12717), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12558), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12590) );
  NAND4_X1 U15871 ( .A1(n12593), .A2(n12592), .A3(n12591), .A4(n12590), .ZN(
        n12600) );
  AOI22_X1 U15872 ( .A1(n15302), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12598) );
  AOI22_X1 U15873 ( .A1(n12687), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15283), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12597) );
  AOI22_X1 U15874 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12605), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U15875 ( .A1(n12696), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12595) );
  NAND4_X1 U15876 ( .A1(n12598), .A2(n12597), .A3(n12596), .A4(n12595), .ZN(
        n12599) );
  NAND2_X1 U15877 ( .A1(n15283), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12604) );
  NAND2_X1 U15878 ( .A1(n9707), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12609) );
  NAND2_X1 U15879 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12608) );
  NAND2_X1 U15880 ( .A1(n9699), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12607) );
  NAND2_X1 U15881 ( .A1(n12605), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12606) );
  NAND2_X1 U15882 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12615) );
  NAND2_X1 U15883 ( .A1(n12611), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12614) );
  NAND2_X1 U15884 ( .A1(n12612), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12613) );
  NAND3_X1 U15885 ( .A1(n12615), .A2(n12614), .A3(n12613), .ZN(n12616) );
  NAND2_X1 U15886 ( .A1(n12536), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12621) );
  NAND2_X1 U15887 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12620) );
  NAND2_X1 U15888 ( .A1(n9702), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12619) );
  NAND2_X1 U15889 ( .A1(n12558), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12618) );
  NAND4_X4 U15890 ( .A1(n12625), .A2(n12624), .A3(n12623), .A4(n12622), .ZN(
        n15395) );
  AND2_X2 U15891 ( .A1(n12966), .A2(n14469), .ZN(n13130) );
  INV_X1 U15892 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n12628) );
  INV_X1 U15893 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n12627) );
  NAND2_X1 U15894 ( .A1(n12628), .A2(n12627), .ZN(n21645) );
  NAND2_X1 U15895 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12629) );
  NAND2_X1 U15896 ( .A1(n12929), .A2(n12632), .ZN(n12633) );
  NAND2_X1 U15897 ( .A1(n12633), .A2(n14464), .ZN(n12647) );
  INV_X1 U15898 ( .A(n12647), .ZN(n12971) );
  NAND3_X1 U15899 ( .A1(n12971), .A2(n12695), .A3(n12635), .ZN(n12973) );
  NAND2_X1 U15900 ( .A1(n12973), .A2(n13766), .ZN(n12637) );
  INV_X2 U15901 ( .A(n15395), .ZN(n12924) );
  AND2_X4 U15902 ( .A1(n12924), .A2(n14449), .ZN(n21761) );
  AND2_X1 U15903 ( .A1(n14449), .A2(n14460), .ZN(n13131) );
  INV_X1 U15904 ( .A(n12638), .ZN(n12639) );
  NAND2_X1 U15905 ( .A1(n15394), .A2(n15395), .ZN(n15776) );
  NAND2_X1 U15906 ( .A1(n21733), .A2(n21638), .ZN(n13523) );
  NAND2_X1 U15907 ( .A1(n21575), .A2(n21422), .ZN(n21522) );
  NAND2_X1 U15908 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21571) );
  NAND2_X1 U15909 ( .A1(n21522), .A2(n21571), .ZN(n21393) );
  OR2_X1 U15910 ( .A1(n17854), .A2(n21575), .ZN(n12653) );
  OAI21_X1 U15911 ( .B1(n13523), .B2(n21393), .A(n12653), .ZN(n12640) );
  INV_X1 U15912 ( .A(n12640), .ZN(n12641) );
  MUX2_X1 U15913 ( .A(n17854), .B(n13523), .S(n21422), .Z(n12642) );
  INV_X1 U15914 ( .A(n12643), .ZN(n12645) );
  INV_X1 U15915 ( .A(n13145), .ZN(n12644) );
  OAI21_X1 U15916 ( .B1(n12645), .B2(n15395), .A(n12644), .ZN(n12651) );
  OR2_X1 U15917 ( .A1(n13744), .A2(n12632), .ZN(n13139) );
  NAND2_X1 U15918 ( .A1(n21733), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20985) );
  INV_X1 U15919 ( .A(n20985), .ZN(n12646) );
  AND3_X1 U15920 ( .A1(n13139), .A2(n12646), .A3(n15776), .ZN(n12650) );
  INV_X1 U15921 ( .A(n15772), .ZN(n13619) );
  AOI22_X1 U15922 ( .A1(n15443), .A2(n12648), .B1(n12647), .B2(n21761), .ZN(
        n12649) );
  NAND4_X1 U15923 ( .A1(n12651), .A2(n13136), .A3(n12650), .A4(n12649), .ZN(
        n12681) );
  NAND2_X1 U15924 ( .A1(n12653), .A2(n13740), .ZN(n12654) );
  NAND2_X1 U15925 ( .A1(n12655), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12657) );
  INV_X1 U15926 ( .A(n13523), .ZN(n12740) );
  XNOR2_X1 U15927 ( .A(n21571), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14712) );
  NAND2_X1 U15928 ( .A1(n12740), .A2(n14712), .ZN(n12656) );
  NOR2_X1 U15929 ( .A1(n17854), .A2(n21392), .ZN(n12660) );
  INV_X1 U15930 ( .A(n12659), .ZN(n12663) );
  INV_X1 U15931 ( .A(n12660), .ZN(n12661) );
  NAND4_X1 U15932 ( .A1(n12732), .A2(n12663), .A3(n12662), .A4(n12661), .ZN(
        n12664) );
  AOI22_X1 U15933 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(n9704), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12669) );
  INV_X1 U15934 ( .A(n12687), .ZN(n12762) );
  AOI22_X1 U15935 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12668) );
  INV_X1 U15936 ( .A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14102) );
  AOI22_X1 U15937 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12667) );
  AOI22_X1 U15938 ( .A1(n15341), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12666) );
  NAND4_X1 U15939 ( .A1(n12669), .A2(n12668), .A3(n12667), .A4(n12666), .ZN(
        n12675) );
  AOI22_X1 U15940 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12673) );
  AOI22_X1 U15941 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12672) );
  AOI22_X1 U15942 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12671) );
  AOI22_X1 U15943 ( .A1(n12717), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12670) );
  NAND4_X1 U15944 ( .A1(n12673), .A2(n12672), .A3(n12671), .A4(n12670), .ZN(
        n12674) );
  NAND2_X1 U15945 ( .A1(n12743), .A2(n12677), .ZN(n12676) );
  INV_X1 U15946 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12678) );
  OAI22_X1 U15947 ( .A1(n12778), .A2(n12744), .B1(n12940), .B2(n12678), .ZN(
        n12679) );
  INV_X1 U15948 ( .A(n12681), .ZN(n12682) );
  AOI22_X1 U15949 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12612), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12686) );
  AOI22_X1 U15950 ( .A1(n12536), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12685) );
  AOI22_X1 U15951 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U15952 ( .A1(n12717), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12683) );
  NAND4_X1 U15953 ( .A1(n12686), .A2(n12685), .A3(n12684), .A4(n12683), .ZN(
        n12693) );
  AOI22_X1 U15954 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12691) );
  AOI22_X1 U15955 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12690) );
  AOI22_X1 U15956 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12689) );
  AOI22_X1 U15957 ( .A1(n12696), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12688) );
  NAND4_X1 U15958 ( .A1(n12691), .A2(n12690), .A3(n12689), .A4(n12688), .ZN(
        n12692) );
  INV_X1 U15959 ( .A(n12862), .ZN(n12694) );
  NAND2_X1 U15960 ( .A1(n12695), .A2(n12862), .ZN(n12709) );
  AOI22_X1 U15961 ( .A1(n9699), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12700) );
  AOI22_X1 U15962 ( .A1(n12536), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12699) );
  AOI22_X1 U15963 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12698) );
  AOI22_X1 U15964 ( .A1(n15362), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12697) );
  NAND4_X1 U15965 ( .A1(n12700), .A2(n12699), .A3(n12698), .A4(n12697), .ZN(
        n12706) );
  AOI22_X1 U15966 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12704) );
  AOI22_X1 U15967 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12703) );
  AOI22_X1 U15968 ( .A1(n12717), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12702) );
  AOI22_X1 U15969 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12701) );
  NAND4_X1 U15970 ( .A1(n12704), .A2(n12703), .A3(n12702), .A4(n12701), .ZN(
        n12705) );
  MUX2_X1 U15971 ( .A(n12712), .B(n12865), .S(n12790), .Z(n12707) );
  INV_X1 U15972 ( .A(n12707), .ZN(n12708) );
  INV_X1 U15973 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12711) );
  AOI21_X1 U15974 ( .B1(n15394), .B2(n12769), .A(n21638), .ZN(n12710) );
  OAI211_X1 U15975 ( .C1(n12940), .C2(n12711), .A(n12710), .B(n12709), .ZN(
        n12783) );
  INV_X1 U15976 ( .A(n12712), .ZN(n12728) );
  NAND2_X1 U15977 ( .A1(n12948), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12727) );
  INV_X1 U15978 ( .A(n12744), .ZN(n12725) );
  AOI22_X1 U15979 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9694), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12716) );
  AOI22_X1 U15980 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12715) );
  AOI22_X1 U15981 ( .A1(n15362), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15341), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12714) );
  AOI22_X1 U15982 ( .A1(n12617), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12713) );
  NAND4_X1 U15983 ( .A1(n12716), .A2(n12715), .A3(n12714), .A4(n12713), .ZN(
        n12724) );
  AOI22_X1 U15984 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U15985 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12717), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U15986 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12720) );
  AOI22_X1 U15987 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12719) );
  NAND4_X1 U15988 ( .A1(n12722), .A2(n12721), .A3(n12720), .A4(n12719), .ZN(
        n12723) );
  NAND2_X1 U15989 ( .A1(n12725), .A2(n12789), .ZN(n12726) );
  INV_X1 U15990 ( .A(n14442), .ZN(n12731) );
  INV_X1 U15991 ( .A(n12729), .ZN(n12730) );
  INV_X1 U15992 ( .A(n12734), .ZN(n12735) );
  NAND2_X1 U15993 ( .A1(n12655), .A2(n21737), .ZN(n12742) );
  OAI21_X1 U15994 ( .B1(n21571), .B2(n21392), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12739) );
  INV_X1 U15995 ( .A(n21571), .ZN(n21289) );
  NAND2_X1 U15996 ( .A1(n12902), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n21361) );
  INV_X1 U15997 ( .A(n21361), .ZN(n12738) );
  NAND2_X1 U15998 ( .A1(n21289), .A2(n12738), .ZN(n14480) );
  NAND2_X1 U15999 ( .A1(n12739), .A2(n14480), .ZN(n21394) );
  INV_X1 U16000 ( .A(n17854), .ZN(n17848) );
  AOI22_X1 U16001 ( .A1(n12740), .A2(n21394), .B1(n17848), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U16002 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U16003 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12748) );
  AOI22_X1 U16004 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12747) );
  AOI22_X1 U16005 ( .A1(n12717), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12746) );
  NAND4_X1 U16006 ( .A1(n12749), .A2(n12748), .A3(n12747), .A4(n12746), .ZN(
        n12755) );
  AOI22_X1 U16007 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12753) );
  AOI22_X1 U16008 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12752) );
  AOI22_X1 U16009 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U16010 ( .A1(n15341), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12750) );
  NAND4_X1 U16011 ( .A1(n12753), .A2(n12752), .A3(n12751), .A4(n12750), .ZN(
        n12754) );
  AOI22_X1 U16012 ( .A1(n12959), .A2(n12804), .B1(n12948), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U16013 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12761) );
  AOI22_X1 U16014 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U16015 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U16016 ( .A1(n12717), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12758) );
  NAND4_X1 U16017 ( .A1(n12761), .A2(n12760), .A3(n12759), .A4(n12758), .ZN(
        n12768) );
  AOI22_X1 U16018 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n9694), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12766) );
  AOI22_X1 U16019 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12718), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12765) );
  INV_X1 U16020 ( .A(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14182) );
  AOI22_X1 U16021 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12764) );
  AOI22_X1 U16022 ( .A1(n15341), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12763) );
  NAND4_X1 U16023 ( .A1(n12766), .A2(n12765), .A3(n12764), .A4(n12763), .ZN(
        n12767) );
  XNOR2_X1 U16024 ( .A(n12811), .B(n10501), .ZN(n14547) );
  NAND2_X1 U16025 ( .A1(n14547), .A2(n12921), .ZN(n12772) );
  NAND2_X1 U16026 ( .A1(n12769), .A2(n12789), .ZN(n12777) );
  NAND2_X1 U16027 ( .A1(n12777), .A2(n12778), .ZN(n12803) );
  NAND2_X1 U16028 ( .A1(n12803), .A2(n12804), .ZN(n12827) );
  XNOR2_X1 U16029 ( .A(n12827), .B(n12825), .ZN(n12770) );
  NAND2_X1 U16030 ( .A1(n12770), .A2(n21761), .ZN(n12771) );
  INV_X1 U16031 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12773) );
  NAND2_X1 U16032 ( .A1(n12775), .A2(n12774), .ZN(n12776) );
  INV_X1 U16033 ( .A(n12921), .ZN(n13518) );
  OAI21_X1 U16034 ( .B1(n12778), .B2(n12777), .A(n12803), .ZN(n12780) );
  NAND2_X1 U16035 ( .A1(n15394), .A2(n14469), .ZN(n12784) );
  INV_X1 U16036 ( .A(n12784), .ZN(n12779) );
  AOI21_X1 U16037 ( .B1(n12780), .B2(n21761), .A(n12779), .ZN(n12781) );
  NAND2_X1 U16038 ( .A1(n12782), .A2(n12781), .ZN(n13794) );
  NAND2_X1 U16039 ( .A1(n21761), .A2(n12790), .ZN(n12785) );
  AND2_X1 U16040 ( .A1(n12785), .A2(n12784), .ZN(n13517) );
  AND2_X1 U16041 ( .A1(n13518), .A2(n12784), .ZN(n12786) );
  INV_X1 U16042 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13765) );
  AOI21_X1 U16043 ( .B1(n12786), .B2(n12785), .A(n13765), .ZN(n12787) );
  NAND2_X1 U16044 ( .A1(n13680), .A2(n15395), .ZN(n12794) );
  XNOR2_X1 U16045 ( .A(n12790), .B(n12789), .ZN(n12791) );
  NAND2_X1 U16046 ( .A1(n12791), .A2(n21761), .ZN(n12792) );
  AND3_X1 U16047 ( .A1(n13130), .A2(n12792), .A3(n15823), .ZN(n12793) );
  NAND2_X1 U16048 ( .A1(n12794), .A2(n12793), .ZN(n12795) );
  NAND2_X1 U16049 ( .A1(n13583), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12798) );
  INV_X1 U16050 ( .A(n12795), .ZN(n12796) );
  OR2_X1 U16051 ( .A1(n12796), .A2(n13519), .ZN(n12797) );
  INV_X1 U16052 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12995) );
  NAND2_X1 U16053 ( .A1(n12799), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12800) );
  OAI211_X1 U16054 ( .C1(n12804), .C2(n12803), .A(n12827), .B(n21761), .ZN(
        n12805) );
  AOI22_X1 U16055 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12815) );
  AOI22_X1 U16056 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12814) );
  AOI22_X1 U16057 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12813) );
  AOI22_X1 U16058 ( .A1(n12717), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12812) );
  NAND4_X1 U16059 ( .A1(n12815), .A2(n12814), .A3(n12813), .A4(n12812), .ZN(
        n12821) );
  AOI22_X1 U16060 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12819) );
  AOI22_X1 U16061 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U16062 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12817) );
  AOI22_X1 U16063 ( .A1(n15341), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12816) );
  NAND4_X1 U16064 ( .A1(n12819), .A2(n12818), .A3(n12817), .A4(n12816), .ZN(
        n12820) );
  NAND2_X1 U16065 ( .A1(n12959), .A2(n12828), .ZN(n12823) );
  NAND2_X1 U16066 ( .A1(n12948), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12822) );
  NAND2_X1 U16067 ( .A1(n10499), .A2(n9843), .ZN(n12824) );
  INV_X1 U16068 ( .A(n12825), .ZN(n12826) );
  NOR2_X1 U16069 ( .A1(n12827), .A2(n12826), .ZN(n12829) );
  NAND2_X1 U16070 ( .A1(n12829), .A2(n12828), .ZN(n12854) );
  OAI211_X1 U16071 ( .C1(n12829), .C2(n12828), .A(n12854), .B(n21761), .ZN(
        n12830) );
  NAND2_X1 U16072 ( .A1(n12831), .A2(n12830), .ZN(n12832) );
  INV_X1 U16073 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17917) );
  XNOR2_X1 U16074 ( .A(n12832), .B(n17917), .ZN(n17878) );
  AOI22_X1 U16075 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12837) );
  AOI22_X1 U16076 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12836) );
  AOI22_X1 U16077 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U16078 ( .A1(n15361), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12834) );
  NAND4_X1 U16079 ( .A1(n12837), .A2(n12836), .A3(n12835), .A4(n12834), .ZN(
        n12843) );
  AOI22_X1 U16080 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(n9704), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12841) );
  AOI22_X1 U16081 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12840) );
  INV_X1 U16082 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14076) );
  AOI22_X1 U16083 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12839) );
  AOI22_X1 U16084 ( .A1(n15341), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12838) );
  NAND4_X1 U16085 ( .A1(n12841), .A2(n12840), .A3(n12839), .A4(n12838), .ZN(
        n12842) );
  AOI22_X1 U16086 ( .A1(n12959), .A2(n12855), .B1(n12948), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12845) );
  INV_X1 U16087 ( .A(n12845), .ZN(n12844) );
  NAND2_X1 U16088 ( .A1(n12846), .A2(n12845), .ZN(n14751) );
  NAND3_X1 U16089 ( .A1(n12867), .A2(n14751), .A3(n12921), .ZN(n12849) );
  XNOR2_X1 U16090 ( .A(n12854), .B(n12855), .ZN(n12847) );
  NAND2_X1 U16091 ( .A1(n12847), .A2(n21761), .ZN(n12848) );
  NAND2_X1 U16092 ( .A1(n12849), .A2(n12848), .ZN(n12850) );
  OR2_X1 U16093 ( .A1(n12850), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17873) );
  NAND2_X1 U16094 ( .A1(n12850), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17872) );
  NAND2_X1 U16095 ( .A1(n12959), .A2(n12862), .ZN(n12852) );
  NAND2_X1 U16096 ( .A1(n12948), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12851) );
  NAND2_X1 U16097 ( .A1(n12852), .A2(n12851), .ZN(n12853) );
  NAND2_X1 U16098 ( .A1(n14752), .A2(n12921), .ZN(n12859) );
  INV_X1 U16099 ( .A(n12854), .ZN(n12856) );
  NAND2_X1 U16100 ( .A1(n12856), .A2(n12855), .ZN(n12864) );
  XNOR2_X1 U16101 ( .A(n12864), .B(n12862), .ZN(n12857) );
  NAND2_X1 U16102 ( .A1(n12857), .A2(n21761), .ZN(n12858) );
  NAND2_X1 U16103 ( .A1(n12859), .A2(n12858), .ZN(n12860) );
  XNOR2_X1 U16104 ( .A(n12860), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17863) );
  NAND2_X1 U16105 ( .A1(n21761), .A2(n12862), .ZN(n12863) );
  OR2_X1 U16106 ( .A1(n12864), .A2(n12863), .ZN(n16091) );
  AND2_X1 U16107 ( .A1(n12865), .A2(n12921), .ZN(n12866) );
  OAI21_X1 U16108 ( .B1(n16091), .B2(n17898), .A(n12890), .ZN(n12868) );
  OAI21_X1 U16109 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n12868), .ZN(n12869) );
  NAND2_X1 U16110 ( .A1(n16091), .A2(n17898), .ZN(n12870) );
  NAND2_X1 U16111 ( .A1(n12870), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12871) );
  NAND2_X1 U16112 ( .A1(n12890), .A2(n12871), .ZN(n12872) );
  INV_X1 U16113 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16279) );
  NAND2_X1 U16114 ( .A1(n9689), .A2(n16279), .ZN(n12873) );
  NAND2_X1 U16115 ( .A1(n16055), .A2(n12873), .ZN(n16074) );
  INV_X1 U16116 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16070) );
  AND2_X1 U16117 ( .A1(n9689), .A2(n16070), .ZN(n16072) );
  NAND2_X1 U16118 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12874) );
  NAND2_X1 U16119 ( .A1(n12890), .A2(n12874), .ZN(n16065) );
  INV_X1 U16120 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16287) );
  NAND2_X1 U16121 ( .A1(n9689), .A2(n16287), .ZN(n12875) );
  AND2_X1 U16122 ( .A1(n16065), .A2(n12875), .ZN(n12876) );
  NAND2_X1 U16123 ( .A1(n16054), .A2(n12876), .ZN(n16033) );
  OR2_X1 U16124 ( .A1(n12890), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16024) );
  NAND2_X1 U16125 ( .A1(n12890), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12877) );
  NAND2_X1 U16126 ( .A1(n16024), .A2(n12877), .ZN(n16037) );
  INV_X1 U16127 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16260) );
  NAND2_X1 U16128 ( .A1(n9689), .A2(n16260), .ZN(n16047) );
  NAND2_X1 U16129 ( .A1(n16037), .A2(n16047), .ZN(n12878) );
  INV_X1 U16130 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16331) );
  INV_X1 U16131 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16316) );
  AND3_X1 U16132 ( .A1(n16070), .A2(n16331), .A3(n16316), .ZN(n12879) );
  NOR2_X1 U16133 ( .A1(n9689), .A2(n12879), .ZN(n16021) );
  NOR2_X1 U16134 ( .A1(n12880), .A2(n16021), .ZN(n16032) );
  NOR2_X1 U16135 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12881) );
  INV_X1 U16136 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16224) );
  INV_X1 U16137 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16212) );
  INV_X1 U16138 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15986) );
  INV_X1 U16139 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16246) );
  NAND4_X1 U16140 ( .A1(n16224), .A2(n16212), .A3(n15986), .A4(n16246), .ZN(
        n12882) );
  NAND3_X1 U16141 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12883) );
  NAND2_X1 U16142 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15976) );
  NOR2_X1 U16143 ( .A1(n12883), .A2(n15976), .ZN(n12885) );
  INV_X1 U16144 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16202) );
  INV_X1 U16145 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12886) );
  INV_X1 U16146 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15916) );
  INV_X1 U16147 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15959) );
  NAND2_X1 U16148 ( .A1(n15916), .A2(n15959), .ZN(n12887) );
  AND2_X1 U16149 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13157) );
  NAND2_X1 U16150 ( .A1(n13157), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15936) );
  NAND2_X1 U16151 ( .A1(n15918), .A2(n15936), .ZN(n12889) );
  NAND2_X1 U16152 ( .A1(n12888), .A2(n12890), .ZN(n15946) );
  AND2_X1 U16153 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16137) );
  INV_X1 U16154 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16158) );
  INV_X1 U16155 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15920) );
  NAND2_X1 U16156 ( .A1(n16158), .A2(n15920), .ZN(n16146) );
  INV_X1 U16157 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13160) );
  INV_X1 U16158 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12892) );
  XNOR2_X1 U16159 ( .A(n12895), .B(n12894), .ZN(n15387) );
  NAND2_X1 U16160 ( .A1(n21575), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12897) );
  NAND2_X1 U16161 ( .A1(n13740), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12896) );
  NAND2_X1 U16162 ( .A1(n12897), .A2(n12896), .ZN(n12907) );
  NAND2_X1 U16163 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21422), .ZN(
        n12919) );
  NAND2_X1 U16164 ( .A1(n13745), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12898) );
  NAND2_X1 U16165 ( .A1(n12901), .A2(n12898), .ZN(n12910) );
  INV_X1 U16166 ( .A(n12910), .ZN(n12899) );
  MUX2_X1 U16167 ( .A(n12902), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        n14299), .Z(n12905) );
  NAND3_X1 U16168 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12915), .A3(
        n13764), .ZN(n12950) );
  XNOR2_X1 U16169 ( .A(n12906), .B(n12905), .ZN(n12951) );
  NAND2_X1 U16170 ( .A1(n12907), .A2(n12919), .ZN(n12908) );
  NAND2_X1 U16171 ( .A1(n12909), .A2(n12908), .ZN(n12928) );
  NAND2_X1 U16172 ( .A1(n12911), .A2(n12910), .ZN(n12913) );
  NAND2_X1 U16173 ( .A1(n12913), .A2(n12912), .ZN(n12939) );
  NOR2_X1 U16174 ( .A1(n12928), .A2(n12939), .ZN(n12916) );
  INV_X1 U16175 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21184) );
  NOR2_X1 U16176 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21184), .ZN(
        n12914) );
  AOI21_X1 U16177 ( .B1(n12949), .B2(n12916), .A(n12960), .ZN(n13615) );
  NAND2_X1 U16178 ( .A1(n12917), .A2(n21657), .ZN(n15398) );
  NAND2_X1 U16179 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21759) );
  INV_X1 U16180 ( .A(n21759), .ZN(n13209) );
  AOI21_X1 U16181 ( .B1(n15395), .B2(n15398), .A(n13209), .ZN(n12918) );
  NAND2_X1 U16182 ( .A1(n13615), .A2(n12918), .ZN(n12968) );
  OAI21_X1 U16183 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21422), .A(
        n12919), .ZN(n12923) );
  INV_X1 U16184 ( .A(n12923), .ZN(n12920) );
  NAND2_X1 U16185 ( .A1(n12959), .A2(n12920), .ZN(n12922) );
  NAND2_X1 U16186 ( .A1(n12922), .A2(n12952), .ZN(n12927) );
  NAND2_X1 U16187 ( .A1(n12929), .A2(n14449), .ZN(n12925) );
  NAND2_X1 U16188 ( .A1(n12925), .A2(n12924), .ZN(n12943) );
  OAI211_X1 U16189 ( .C1(n12588), .C2(n15394), .A(n12920), .B(n12943), .ZN(
        n12926) );
  INV_X1 U16190 ( .A(n12928), .ZN(n12933) );
  NAND2_X1 U16191 ( .A1(n12959), .A2(n15395), .ZN(n12930) );
  NAND2_X1 U16192 ( .A1(n12929), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12931) );
  OAI211_X1 U16193 ( .C1(n12933), .C2(n12940), .A(n12930), .B(n12931), .ZN(
        n12935) );
  NAND2_X1 U16194 ( .A1(n12931), .A2(n15395), .ZN(n12932) );
  NOR2_X1 U16195 ( .A1(n12959), .A2(n12932), .ZN(n12934) );
  OAI22_X1 U16196 ( .A1(n12936), .A2(n12935), .B1(n12934), .B2(n12933), .ZN(
        n12938) );
  NAND2_X1 U16197 ( .A1(n12936), .A2(n12935), .ZN(n12937) );
  NAND2_X1 U16198 ( .A1(n12938), .A2(n12937), .ZN(n12947) );
  INV_X1 U16199 ( .A(n12939), .ZN(n12941) );
  NAND2_X1 U16200 ( .A1(n12959), .A2(n12941), .ZN(n12942) );
  OAI211_X1 U16201 ( .C1(n12941), .C2(n12940), .A(n12942), .B(n12943), .ZN(
        n12946) );
  INV_X1 U16202 ( .A(n12942), .ZN(n12945) );
  INV_X1 U16203 ( .A(n12943), .ZN(n12944) );
  AOI22_X1 U16204 ( .A1(n12947), .A2(n12946), .B1(n12945), .B2(n12944), .ZN(
        n12957) );
  NOR2_X1 U16205 ( .A1(n12949), .A2(n12948), .ZN(n12956) );
  INV_X1 U16206 ( .A(n12952), .ZN(n12958) );
  INV_X1 U16207 ( .A(n12950), .ZN(n12954) );
  OAI22_X1 U16208 ( .A1(n12952), .A2(n12951), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n13764), .ZN(n12953) );
  AOI21_X1 U16209 ( .B1(n12958), .B2(n12954), .A(n12953), .ZN(n12955) );
  NOR2_X1 U16210 ( .A1(n12962), .A2(n13209), .ZN(n13611) );
  OR2_X1 U16211 ( .A1(n13611), .A2(n15394), .ZN(n12964) );
  NAND2_X1 U16212 ( .A1(n21761), .A2(n15398), .ZN(n12963) );
  AOI21_X1 U16213 ( .B1(n12964), .B2(n12963), .A(n10088), .ZN(n12965) );
  MUX2_X1 U16214 ( .A(n12968), .B(n12967), .S(n12966), .Z(n12975) );
  AND2_X1 U16215 ( .A1(n12969), .A2(n15394), .ZN(n13236) );
  INV_X1 U16216 ( .A(n13236), .ZN(n13304) );
  OR2_X1 U16217 ( .A1(n12635), .A2(n12636), .ZN(n12970) );
  NAND2_X1 U16218 ( .A1(n13766), .A2(n15394), .ZN(n12972) );
  OR2_X1 U16219 ( .A1(n12635), .A2(n12924), .ZN(n13141) );
  AND3_X1 U16220 ( .A1(n12973), .A2(n14449), .A3(n13141), .ZN(n13129) );
  AOI21_X1 U16221 ( .B1(n13304), .B2(n17840), .A(n13129), .ZN(n13756) );
  NAND3_X1 U16222 ( .A1(n13753), .A2(n16350), .A3(n15395), .ZN(n12974) );
  NAND3_X1 U16223 ( .A1(n12975), .A2(n13756), .A3(n12974), .ZN(n12976) );
  INV_X1 U16224 ( .A(n13146), .ZN(n13149) );
  OR2_X1 U16225 ( .A1(n13126), .A2(n15772), .ZN(n12978) );
  NAND2_X1 U16226 ( .A1(n13612), .A2(n12978), .ZN(n13301) );
  INV_X1 U16227 ( .A(n13121), .ZN(n12979) );
  NAND2_X1 U16228 ( .A1(n12979), .A2(n12636), .ZN(n12980) );
  AND4_X1 U16229 ( .A1(n12981), .A2(n12977), .A3(n13301), .A4(n12980), .ZN(
        n12982) );
  NAND2_X1 U16230 ( .A1(n9750), .A2(n13113), .ZN(n12993) );
  OR2_X1 U16231 ( .A1(n12993), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n12988) );
  INV_X1 U16232 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12983) );
  NAND2_X1 U16233 ( .A1(n13113), .A2(n12983), .ZN(n12986) );
  INV_X1 U16234 ( .A(n14469), .ZN(n12984) );
  INV_X1 U16235 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13582) );
  NAND2_X1 U16236 ( .A1(n12994), .A2(n13582), .ZN(n12985) );
  NAND3_X1 U16237 ( .A1(n12986), .A2(n12985), .A3(n9701), .ZN(n12987) );
  NAND2_X1 U16238 ( .A1(n12988), .A2(n12987), .ZN(n12991) );
  NAND2_X1 U16239 ( .A1(n12994), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12990) );
  INV_X1 U16240 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13510) );
  NAND2_X1 U16241 ( .A1(n9700), .A2(n13510), .ZN(n12989) );
  NAND2_X1 U16242 ( .A1(n12990), .A2(n12989), .ZN(n13491) );
  XNOR2_X1 U16243 ( .A(n12991), .B(n13491), .ZN(n13585) );
  NAND2_X1 U16244 ( .A1(n13585), .A2(n13610), .ZN(n13584) );
  OR2_X1 U16245 ( .A1(n12993), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n12999) );
  NAND2_X1 U16246 ( .A1(n12994), .A2(n12995), .ZN(n12997) );
  INV_X1 U16247 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n21090) );
  NAND2_X1 U16248 ( .A1(n13610), .A2(n21090), .ZN(n12996) );
  NAND3_X1 U16249 ( .A1(n12997), .A2(n9701), .A3(n12996), .ZN(n12998) );
  AND2_X1 U16250 ( .A1(n12999), .A2(n12998), .ZN(n13801) );
  MUX2_X1 U16251 ( .A(n13104), .B(n9701), .S(P1_EBX_REG_3__SCAN_IN), .Z(n13001) );
  OAI21_X1 U16252 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13490), .A(
        n13001), .ZN(n14536) );
  OR2_X1 U16253 ( .A1(n12993), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n13007) );
  NAND2_X1 U16254 ( .A1(n9700), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13002) );
  NAND2_X1 U16255 ( .A1(n12994), .A2(n13002), .ZN(n13005) );
  INV_X1 U16256 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13003) );
  NAND2_X1 U16257 ( .A1(n13610), .A2(n13003), .ZN(n13004) );
  NAND2_X1 U16258 ( .A1(n13005), .A2(n13004), .ZN(n13006) );
  NAND2_X1 U16259 ( .A1(n13007), .A2(n13006), .ZN(n14585) );
  INV_X1 U16260 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n21108) );
  NAND2_X1 U16261 ( .A1(n13610), .A2(n21108), .ZN(n13009) );
  NAND2_X1 U16262 ( .A1(n9701), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13008) );
  NAND3_X1 U16263 ( .A1(n13009), .A2(n12994), .A3(n13008), .ZN(n13010) );
  OAI21_X1 U16264 ( .B1(n13104), .B2(P1_EBX_REG_5__SCAN_IN), .A(n13010), .ZN(
        n17913) );
  INV_X1 U16265 ( .A(n17913), .ZN(n13011) );
  OR2_X1 U16266 ( .A1(n12993), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n13017) );
  NAND2_X1 U16267 ( .A1(n9700), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13012) );
  NAND2_X1 U16268 ( .A1(n12994), .A2(n13012), .ZN(n13015) );
  INV_X1 U16269 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n13013) );
  NAND2_X1 U16270 ( .A1(n13610), .A2(n13013), .ZN(n13014) );
  NAND2_X1 U16271 ( .A1(n13015), .A2(n13014), .ZN(n13016) );
  INV_X1 U16272 ( .A(n13104), .ZN(n13018) );
  INV_X1 U16273 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13019) );
  NAND2_X1 U16274 ( .A1(n13018), .A2(n13019), .ZN(n13023) );
  NAND2_X1 U16275 ( .A1(n13610), .A2(n13019), .ZN(n13021) );
  NAND2_X1 U16276 ( .A1(n9701), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13020) );
  NAND3_X1 U16277 ( .A1(n13021), .A2(n12994), .A3(n13020), .ZN(n13022) );
  OR2_X1 U16278 ( .A1(n12993), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n13028) );
  NAND2_X1 U16279 ( .A1(n9700), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13024) );
  NAND2_X1 U16280 ( .A1(n12994), .A2(n13024), .ZN(n13026) );
  INV_X1 U16281 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n15767) );
  NAND2_X1 U16282 ( .A1(n13610), .A2(n15767), .ZN(n13025) );
  NAND2_X1 U16283 ( .A1(n13026), .A2(n13025), .ZN(n13027) );
  NAND2_X1 U16284 ( .A1(n13028), .A2(n13027), .ZN(n15762) );
  NAND2_X1 U16285 ( .A1(n14762), .A2(n15762), .ZN(n15761) );
  INV_X1 U16286 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n21104) );
  NAND2_X1 U16287 ( .A1(n13610), .A2(n21104), .ZN(n13030) );
  NAND2_X1 U16288 ( .A1(n9701), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13029) );
  NAND3_X1 U16289 ( .A1(n13030), .A2(n12994), .A3(n13029), .ZN(n13031) );
  OAI21_X1 U16290 ( .B1(n13104), .B2(P1_EBX_REG_9__SCAN_IN), .A(n13031), .ZN(
        n16341) );
  MUX2_X1 U16291 ( .A(n13104), .B(n9700), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13033) );
  OR2_X1 U16292 ( .A1(n13490), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13032) );
  OR2_X1 U16293 ( .A1(n12993), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n13038) );
  NAND2_X1 U16294 ( .A1(n12994), .A2(n16331), .ZN(n13036) );
  INV_X1 U16295 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15751) );
  NAND2_X1 U16296 ( .A1(n13610), .A2(n15751), .ZN(n13034) );
  NAND3_X1 U16297 ( .A1(n13036), .A2(n9700), .A3(n13034), .ZN(n13037) );
  NAND2_X1 U16298 ( .A1(n13038), .A2(n13037), .ZN(n15743) );
  NAND2_X1 U16299 ( .A1(n10543), .A2(n15743), .ZN(n13039) );
  OR2_X1 U16300 ( .A1(n12993), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n13044) );
  NAND2_X1 U16301 ( .A1(n9701), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13040) );
  NAND2_X1 U16302 ( .A1(n12994), .A2(n13040), .ZN(n13042) );
  INV_X1 U16303 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15815) );
  NAND2_X1 U16304 ( .A1(n13610), .A2(n15815), .ZN(n13041) );
  NAND2_X1 U16305 ( .A1(n13042), .A2(n13041), .ZN(n13043) );
  NAND2_X1 U16306 ( .A1(n13044), .A2(n13043), .ZN(n15719) );
  MUX2_X1 U16307 ( .A(n13104), .B(n9700), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n13046) );
  OR2_X1 U16308 ( .A1(n13490), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13045) );
  NAND2_X1 U16309 ( .A1(n13046), .A2(n13045), .ZN(n15710) );
  INV_X1 U16310 ( .A(n15710), .ZN(n13047) );
  OR2_X1 U16311 ( .A1(n12993), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n13052) );
  NAND2_X1 U16312 ( .A1(n12994), .A2(n16287), .ZN(n13050) );
  INV_X1 U16313 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n13048) );
  NAND2_X1 U16314 ( .A1(n13610), .A2(n13048), .ZN(n13049) );
  NAND3_X1 U16315 ( .A1(n13050), .A2(n9701), .A3(n13049), .ZN(n13051) );
  MUX2_X1 U16316 ( .A(n13104), .B(n9701), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n13055) );
  OAI21_X1 U16317 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n13490), .A(
        n13055), .ZN(n15669) );
  OR2_X1 U16318 ( .A1(n12993), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n13059) );
  INV_X1 U16319 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16261) );
  NAND2_X1 U16320 ( .A1(n12994), .A2(n16261), .ZN(n13057) );
  INV_X1 U16321 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15811) );
  NAND2_X1 U16322 ( .A1(n13610), .A2(n15811), .ZN(n13056) );
  NAND3_X1 U16323 ( .A1(n13057), .A2(n9701), .A3(n13056), .ZN(n13058) );
  NAND2_X1 U16324 ( .A1(n13059), .A2(n13058), .ZN(n15654) );
  MUX2_X1 U16325 ( .A(n13104), .B(n9700), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n13064) );
  INV_X1 U16326 ( .A(n13490), .ZN(n13062) );
  INV_X1 U16327 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13061) );
  NAND2_X1 U16328 ( .A1(n13062), .A2(n13061), .ZN(n13063) );
  NAND2_X1 U16329 ( .A1(n13064), .A2(n13063), .ZN(n15648) );
  OR2_X1 U16330 ( .A1(n12993), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n13071) );
  NAND2_X1 U16331 ( .A1(n12994), .A2(n16246), .ZN(n13069) );
  INV_X1 U16332 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n13067) );
  NAND2_X1 U16333 ( .A1(n13610), .A2(n13067), .ZN(n13068) );
  NAND3_X1 U16334 ( .A1(n13069), .A2(n9701), .A3(n13068), .ZN(n13070) );
  AND2_X1 U16335 ( .A1(n13071), .A2(n13070), .ZN(n15630) );
  MUX2_X1 U16336 ( .A(n13104), .B(n9701), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n13074) );
  OAI21_X1 U16337 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n13490), .A(
        n13074), .ZN(n15610) );
  OR2_X1 U16338 ( .A1(n12993), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n13080) );
  NAND2_X1 U16339 ( .A1(n9701), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13075) );
  NAND2_X1 U16340 ( .A1(n12994), .A2(n13075), .ZN(n13078) );
  INV_X1 U16341 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n13076) );
  NAND2_X1 U16342 ( .A1(n13610), .A2(n13076), .ZN(n13077) );
  NAND2_X1 U16343 ( .A1(n13078), .A2(n13077), .ZN(n13079) );
  MUX2_X1 U16344 ( .A(n13104), .B(n9701), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n13082) );
  OR2_X1 U16345 ( .A1(n13490), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13081) );
  NAND2_X1 U16346 ( .A1(n13082), .A2(n13081), .ZN(n15587) );
  INV_X1 U16347 ( .A(n15587), .ZN(n13083) );
  OR2_X1 U16348 ( .A1(n12993), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n13087) );
  NAND2_X1 U16349 ( .A1(n12994), .A2(n16202), .ZN(n13085) );
  INV_X1 U16350 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15805) );
  NAND2_X1 U16351 ( .A1(n13610), .A2(n15805), .ZN(n13084) );
  NAND3_X1 U16352 ( .A1(n13085), .A2(n9701), .A3(n13084), .ZN(n13086) );
  AND2_X1 U16353 ( .A1(n13087), .A2(n13086), .ZN(n15571) );
  INV_X1 U16354 ( .A(n13088), .ZN(n15549) );
  INV_X1 U16355 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15803) );
  NAND2_X1 U16356 ( .A1(n13610), .A2(n15803), .ZN(n13090) );
  NAND2_X1 U16357 ( .A1(n9700), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13089) );
  NAND3_X1 U16358 ( .A1(n13090), .A2(n12994), .A3(n13089), .ZN(n13091) );
  OAI21_X1 U16359 ( .B1(n13104), .B2(P1_EBX_REG_23__SCAN_IN), .A(n13091), .ZN(
        n15550) );
  OR2_X1 U16360 ( .A1(n12993), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n13096) );
  NAND2_X1 U16361 ( .A1(n12994), .A2(n15959), .ZN(n13094) );
  INV_X1 U16362 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n13092) );
  NAND2_X1 U16363 ( .A1(n13610), .A2(n13092), .ZN(n13093) );
  NAND3_X1 U16364 ( .A1(n13094), .A2(n9701), .A3(n13093), .ZN(n13095) );
  NAND2_X1 U16365 ( .A1(n13096), .A2(n13095), .ZN(n15536) );
  MUX2_X1 U16366 ( .A(n13104), .B(n9701), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n13098) );
  OR2_X1 U16367 ( .A1(n13490), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13097) );
  AND2_X1 U16368 ( .A1(n13098), .A2(n13097), .ZN(n15519) );
  OR2_X1 U16369 ( .A1(n12993), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n13103) );
  INV_X1 U16370 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15939) );
  NAND2_X1 U16371 ( .A1(n12994), .A2(n15939), .ZN(n13101) );
  INV_X1 U16372 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n13099) );
  NAND2_X1 U16373 ( .A1(n13610), .A2(n13099), .ZN(n13100) );
  NAND3_X1 U16374 ( .A1(n13101), .A2(n9701), .A3(n13100), .ZN(n13102) );
  AND2_X1 U16375 ( .A1(n13103), .A2(n13102), .ZN(n15505) );
  MUX2_X1 U16376 ( .A(n13104), .B(n9701), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n13105) );
  OAI21_X1 U16377 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13490), .A(
        n13105), .ZN(n15492) );
  OR2_X1 U16378 ( .A1(n12993), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n13109) );
  NAND2_X1 U16379 ( .A1(n12994), .A2(n15920), .ZN(n13107) );
  INV_X1 U16380 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n15798) );
  NAND2_X1 U16381 ( .A1(n13610), .A2(n15798), .ZN(n13106) );
  NAND3_X1 U16382 ( .A1(n13107), .A2(n9701), .A3(n13106), .ZN(n13108) );
  NAND2_X1 U16383 ( .A1(n13109), .A2(n13108), .ZN(n15477) );
  INV_X1 U16384 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15797) );
  NAND2_X1 U16385 ( .A1(n13610), .A2(n15797), .ZN(n13111) );
  OR2_X1 U16386 ( .A1(n13490), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13110) );
  NAND2_X1 U16387 ( .A1(n13110), .A2(n13111), .ZN(n15460) );
  MUX2_X1 U16388 ( .A(n13111), .B(n15460), .S(n9701), .Z(n15466) );
  NOR2_X2 U16389 ( .A1(n15459), .A2(n15466), .ZN(n13112) );
  INV_X1 U16390 ( .A(n13112), .ZN(n15468) );
  INV_X1 U16391 ( .A(n13113), .ZN(n13497) );
  AOI22_X1 U16392 ( .A1(n13490), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n13497), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15461) );
  AOI22_X1 U16393 ( .A1(n13490), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n13497), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13116) );
  INV_X1 U16394 ( .A(n13116), .ZN(n13117) );
  INV_X1 U16395 ( .A(n15388), .ZN(n13123) );
  NAND2_X1 U16396 ( .A1(n13119), .A2(n12924), .ZN(n13120) );
  OAI21_X1 U16397 ( .B1(n13121), .B2(n12636), .A(n13120), .ZN(n13122) );
  NAND2_X1 U16398 ( .A1(n13123), .A2(n17922), .ZN(n13174) );
  INV_X1 U16399 ( .A(n15776), .ZN(n13124) );
  AND2_X1 U16400 ( .A1(n12969), .A2(n13124), .ZN(n13751) );
  AOI21_X1 U16401 ( .B1(n13500), .B2(n14460), .A(n15824), .ZN(n13125) );
  OAI211_X1 U16402 ( .C1(n13126), .C2(n14449), .A(n13744), .B(n13125), .ZN(
        n13127) );
  AND2_X1 U16403 ( .A1(n13127), .A2(n15395), .ZN(n13128) );
  NOR2_X1 U16404 ( .A1(n13129), .A2(n13128), .ZN(n13138) );
  INV_X1 U16405 ( .A(n13130), .ZN(n13132) );
  AOI21_X1 U16406 ( .B1(n13132), .B2(n13490), .A(n13131), .ZN(n13133) );
  OAI21_X1 U16407 ( .B1(n13134), .B2(n9700), .A(n13133), .ZN(n13135) );
  INV_X1 U16408 ( .A(n13135), .ZN(n13137) );
  AND3_X1 U16409 ( .A1(n13138), .A2(n13137), .A3(n13136), .ZN(n13739) );
  OAI211_X1 U16410 ( .C1(n13736), .C2(n14449), .A(n13739), .B(n13139), .ZN(
        n13140) );
  NOR2_X2 U16411 ( .A1(n21180), .A2(n13164), .ZN(n17886) );
  INV_X1 U16412 ( .A(n13141), .ZN(n13143) );
  AND2_X1 U16413 ( .A1(n13143), .A2(n13142), .ZN(n13144) );
  INV_X1 U16414 ( .A(n16259), .ZN(n13159) );
  NAND2_X1 U16415 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16165) );
  NAND2_X1 U16416 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13171) );
  NAND3_X1 U16417 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16327) );
  INV_X1 U16418 ( .A(n16327), .ZN(n16324) );
  AND3_X1 U16419 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16324), .ZN(n16317) );
  NAND2_X1 U16420 ( .A1(n16317), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16305) );
  NOR2_X1 U16421 ( .A1(n16070), .A2(n16305), .ZN(n13148) );
  INV_X1 U16422 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14544) );
  NOR2_X1 U16423 ( .A1(n12773), .A2(n14544), .ZN(n17887) );
  NAND2_X1 U16424 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17887), .ZN(
        n16304) );
  OAI21_X1 U16425 ( .B1(n13765), .B2(n13582), .A(n12995), .ZN(n14541) );
  INV_X1 U16426 ( .A(n14541), .ZN(n13147) );
  NOR2_X1 U16427 ( .A1(n16304), .A2(n13147), .ZN(n16329) );
  NAND2_X1 U16428 ( .A1(n13148), .A2(n16329), .ZN(n16280) );
  INV_X1 U16429 ( .A(n16280), .ZN(n13153) );
  NAND2_X1 U16430 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14539) );
  NOR2_X1 U16431 ( .A1(n16304), .A2(n14539), .ZN(n16298) );
  NAND2_X1 U16432 ( .A1(n16298), .A2(n13148), .ZN(n13162) );
  INV_X1 U16433 ( .A(n13162), .ZN(n13167) );
  OR2_X1 U16434 ( .A1(n17886), .A2(n13167), .ZN(n13152) );
  NAND2_X1 U16435 ( .A1(n13164), .A2(n13765), .ZN(n13151) );
  NAND2_X1 U16436 ( .A1(n13149), .A2(n17899), .ZN(n13150) );
  OAI211_X1 U16437 ( .C1(n16297), .C2(n13153), .A(n13152), .B(n16296), .ZN(
        n16240) );
  NAND4_X1 U16438 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16241) );
  INV_X1 U16439 ( .A(n16241), .ZN(n16243) );
  AND2_X1 U16440 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13154) );
  NAND2_X1 U16441 ( .A1(n16243), .A2(n13154), .ZN(n16230) );
  AND2_X1 U16442 ( .A1(n16259), .A2(n16230), .ZN(n13155) );
  INV_X1 U16443 ( .A(n16296), .ZN(n13797) );
  INV_X1 U16444 ( .A(n17892), .ZN(n13161) );
  INV_X1 U16445 ( .A(n13164), .ZN(n13156) );
  NAND2_X1 U16446 ( .A1(n13156), .A2(n16297), .ZN(n21178) );
  INV_X1 U16447 ( .A(n13157), .ZN(n16182) );
  AOI22_X1 U16448 ( .A1(n21178), .A2(n16182), .B1(n21180), .B2(n15936), .ZN(
        n13158) );
  NAND2_X1 U16449 ( .A1(n16192), .A2(n13158), .ZN(n16178) );
  INV_X1 U16450 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21715) );
  NOR2_X1 U16451 ( .A1(n17899), .A2(n21715), .ZN(n15383) );
  INV_X1 U16452 ( .A(n15383), .ZN(n13173) );
  OR2_X1 U16453 ( .A1(n16297), .A2(n16280), .ZN(n13166) );
  NOR2_X1 U16454 ( .A1(n13765), .A2(n13162), .ZN(n13163) );
  NAND2_X1 U16455 ( .A1(n13164), .A2(n13163), .ZN(n13165) );
  NAND2_X1 U16456 ( .A1(n21180), .A2(n13167), .ZN(n13168) );
  INV_X1 U16457 ( .A(n16230), .ZN(n13169) );
  AND2_X1 U16458 ( .A1(n13169), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13170) );
  NAND2_X1 U16459 ( .A1(n16292), .A2(n13170), .ZN(n16223) );
  INV_X1 U16460 ( .A(n13171), .ZN(n13172) );
  NAND2_X1 U16461 ( .A1(n16210), .A2(n13172), .ZN(n16194) );
  NAND3_X1 U16462 ( .A1(n16156), .A2(n16137), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16131) );
  OAI21_X1 U16463 ( .B1(n15387), .B2(n21175), .A(n10542), .ZN(P1_U3000) );
  NOR2_X1 U16464 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13176) );
  NOR4_X1 U16465 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13175) );
  NAND4_X1 U16466 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13176), .A4(n13175), .ZN(n13189) );
  NOR4_X1 U16467 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13177) );
  NAND3_X1 U16468 ( .A1(n13177), .A2(n21666), .A3(n21694), .ZN(n13183) );
  NOR4_X1 U16469 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(
        P1_ADDRESS_REG_16__SCAN_IN), .A3(P1_ADDRESS_REG_15__SCAN_IN), .A4(
        P1_ADDRESS_REG_14__SCAN_IN), .ZN(n13181) );
  NOR4_X1 U16470 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_18__SCAN_IN), .ZN(n13180) );
  NOR4_X1 U16471 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(
        P1_ADDRESS_REG_8__SCAN_IN), .A3(P1_ADDRESS_REG_7__SCAN_IN), .A4(
        P1_ADDRESS_REG_5__SCAN_IN), .ZN(n13179) );
  NOR4_X1 U16472 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(
        P1_ADDRESS_REG_12__SCAN_IN), .A3(P1_ADDRESS_REG_11__SCAN_IN), .A4(
        P1_ADDRESS_REG_10__SCAN_IN), .ZN(n13178) );
  NAND4_X1 U16473 ( .A1(n13181), .A2(n13180), .A3(n13179), .A4(n13178), .ZN(
        n13182) );
  NOR4_X1 U16474 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(n13183), .A4(n13182), .ZN(n13185) );
  NAND2_X1 U16475 ( .A1(n21661), .A2(n21672), .ZN(n14021) );
  NOR4_X1 U16476 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_4__SCAN_IN), .A3(P1_ADDRESS_REG_1__SCAN_IN), .A4(n14021), .ZN(n13184) );
  NAND2_X1 U16477 ( .A1(n13185), .A2(n13184), .ZN(n13186) );
  INV_X1 U16478 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21756) );
  NOR3_X1 U16479 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n21756), .ZN(n13188) );
  NOR4_X1 U16480 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13187) );
  NAND4_X1 U16481 ( .A1(n15837), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13188), .A4(
        n13187), .ZN(U214) );
  NOR2_X1 U16482 ( .A1(n17488), .A2(n13189), .ZN(n17936) );
  NAND2_X1 U16483 ( .A1(n17936), .A2(U214), .ZN(U212) );
  INV_X1 U16484 ( .A(n17582), .ZN(n13190) );
  INV_X1 U16485 ( .A(n17644), .ZN(n17581) );
  AOI21_X1 U16486 ( .B1(n13190), .B2(n18966), .A(n17581), .ZN(n13192) );
  INV_X1 U16487 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13191) );
  XNOR2_X1 U16488 ( .A(n18950), .B(n13191), .ZN(n17642) );
  NOR2_X1 U16489 ( .A1(n13192), .A2(n17642), .ZN(n17634) );
  AOI211_X1 U16490 ( .C1(n13192), .C2(n17642), .A(n19034), .B(n17634), .ZN(
        n13208) );
  NAND2_X1 U16491 ( .A1(n19280), .A2(n19121), .ZN(n13194) );
  NAND2_X1 U16492 ( .A1(n19281), .A2(n18978), .ZN(n13193) );
  INV_X1 U16493 ( .A(n17631), .ZN(n13195) );
  NOR3_X1 U16494 ( .A1(n18933), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n13195), .ZN(n13207) );
  INV_X1 U16495 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13198) );
  INV_X1 U16496 ( .A(n19079), .ZN(n19404) );
  INV_X1 U16497 ( .A(n12118), .ZN(n17588) );
  OR2_X1 U16498 ( .A1(n19125), .A2(n17600), .ZN(n18066) );
  NOR2_X1 U16499 ( .A1(n18809), .A2(n18066), .ZN(n18057) );
  NOR2_X1 U16500 ( .A1(n18057), .A2(n18969), .ZN(n13196) );
  AOI211_X1 U16501 ( .C1(n19404), .C2(n17588), .A(n13196), .B(n19096), .ZN(
        n18806) );
  INV_X1 U16502 ( .A(n18806), .ZN(n13197) );
  AOI21_X1 U16503 ( .B1(n13199), .B2(n13198), .A(n13197), .ZN(n17591) );
  INV_X1 U16504 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13201) );
  OAI211_X1 U16505 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n12118), .B(n17568), .ZN(n13200) );
  OAI22_X1 U16506 ( .A1(n17591), .A2(n13201), .B1(n18891), .B2(n13200), .ZN(
        n13206) );
  INV_X1 U16507 ( .A(n18058), .ZN(n17586) );
  INV_X1 U16508 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18115) );
  NOR2_X1 U16509 ( .A1(n17586), .A2(n18115), .ZN(n17585) );
  OAI21_X1 U16510 ( .B1(n17585), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n17572), .ZN(n18056) );
  NAND2_X1 U16511 ( .A1(n18813), .A2(n17651), .ZN(n17653) );
  NAND2_X1 U16512 ( .A1(n17651), .A2(n18807), .ZN(n17660) );
  AOI22_X1 U16513 ( .A1(n18978), .A2(n17653), .B1(n19121), .B2(n17660), .ZN(
        n18800) );
  NAND2_X1 U16514 ( .A1(n18800), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17593) );
  INV_X1 U16515 ( .A(n18978), .ZN(n19004) );
  NAND2_X1 U16516 ( .A1(n19004), .A2(n19112), .ZN(n18843) );
  NAND3_X1 U16517 ( .A1(n17593), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n18843), .ZN(n13204) );
  INV_X1 U16518 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n13202) );
  NOR2_X1 U16519 ( .A1(n19110), .A2(n13202), .ZN(n17645) );
  INV_X1 U16520 ( .A(n17645), .ZN(n13203) );
  OAI211_X1 U16521 ( .C1(n18985), .C2(n18056), .A(n13204), .B(n13203), .ZN(
        n13205) );
  OR4_X1 U16522 ( .A1(n13208), .A2(n13207), .A3(n13206), .A4(n13205), .ZN(
        P3_U2802) );
  INV_X1 U16523 ( .A(HOLD), .ZN(n21647) );
  NOR2_X1 U16524 ( .A1(n12627), .A2(n21647), .ZN(n13211) );
  AOI22_X1 U16525 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n13210) );
  NAND2_X1 U16526 ( .A1(n13209), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21644) );
  OAI211_X1 U16527 ( .C1(n13211), .C2(n13210), .A(n15398), .B(n21644), .ZN(
        P1_U3195) );
  NOR2_X1 U16528 ( .A1(n20966), .A2(n14500), .ZN(n14409) );
  NAND2_X1 U16529 ( .A1(n11055), .A2(n20939), .ZN(n14411) );
  INV_X1 U16530 ( .A(n14411), .ZN(n13212) );
  NAND2_X1 U16531 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n13390) );
  INV_X1 U16532 ( .A(n13390), .ZN(n17482) );
  NAND2_X1 U16533 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17482), .ZN(n17860) );
  INV_X1 U16534 ( .A(n17860), .ZN(n14800) );
  NOR4_X1 U16535 ( .A1(n13213), .A2(n14409), .A3(n13212), .A4(n14800), .ZN(
        P2_U3178) );
  INV_X1 U16536 ( .A(n20190), .ZN(n16645) );
  INV_X1 U16537 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n20978) );
  NOR2_X1 U16538 ( .A1(n14411), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15440) );
  INV_X1 U16539 ( .A(n15440), .ZN(n13214) );
  OAI211_X1 U16540 ( .C1(n16645), .C2(n20978), .A(n13221), .B(n13214), .ZN(
        P2_U2814) );
  NOR2_X1 U16541 ( .A1(n14388), .A2(n13215), .ZN(n13216) );
  AND2_X1 U16542 ( .A1(n13217), .A2(n13216), .ZN(n13218) );
  NAND2_X1 U16543 ( .A1(n14389), .A2(n13218), .ZN(n14396) );
  AND2_X1 U16544 ( .A1(n14396), .A2(n14498), .ZN(n20956) );
  OAI21_X1 U16545 ( .B1(n20956), .B2(n14104), .A(n13219), .ZN(P2_U2819) );
  INV_X1 U16546 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13673) );
  NOR3_X4 U16547 ( .A1(n13221), .A2(n13223), .A3(n20963), .ZN(n20279) );
  INV_X1 U16548 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n18780) );
  NAND2_X1 U16549 ( .A1(n17490), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13220) );
  OAI21_X1 U16550 ( .B1(n17490), .B2(n18780), .A(n13220), .ZN(n16791) );
  NAND2_X1 U16551 ( .A1(n20279), .A2(n16791), .ZN(n13231) );
  INV_X1 U16552 ( .A(n13221), .ZN(n13222) );
  OAI21_X1 U16553 ( .B1(n13223), .B2(n20966), .A(n13222), .ZN(n20282) );
  NAND2_X1 U16554 ( .A1(n20282), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13224) );
  OAI211_X1 U16555 ( .C1(n13673), .C2(n13296), .A(n13231), .B(n13224), .ZN(
        P2_U2962) );
  INV_X1 U16556 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13456) );
  INV_X1 U16557 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n13226) );
  NAND2_X1 U16558 ( .A1(n17490), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13225) );
  OAI21_X1 U16559 ( .B1(n17490), .B2(n13226), .A(n13225), .ZN(n16768) );
  NAND2_X1 U16560 ( .A1(n20279), .A2(n16768), .ZN(n13229) );
  NAND2_X1 U16561 ( .A1(n20282), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13227) );
  OAI211_X1 U16562 ( .C1(n13456), .C2(n13296), .A(n13229), .B(n13227), .ZN(
        P2_U2966) );
  INV_X1 U16563 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n20242) );
  NAND2_X1 U16564 ( .A1(n20282), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13228) );
  OAI211_X1 U16565 ( .C1(n20242), .C2(n13296), .A(n13229), .B(n13228), .ZN(
        P2_U2981) );
  INV_X1 U16566 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n20251) );
  NAND2_X1 U16567 ( .A1(n20282), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13230) );
  OAI211_X1 U16568 ( .C1(n20251), .C2(n13296), .A(n13231), .B(n13230), .ZN(
        P2_U2977) );
  INV_X1 U16569 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13235) );
  INV_X1 U16570 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13234) );
  INV_X1 U16571 ( .A(n20282), .ZN(n13270) );
  INV_X1 U16572 ( .A(n20279), .ZN(n13233) );
  INV_X1 U16573 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n13232) );
  INV_X1 U16574 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13675) );
  MUX2_X1 U16575 ( .A(n13232), .B(n13675), .S(n17490), .Z(n14699) );
  OAI222_X1 U16576 ( .A1(n13296), .A2(n13235), .B1(n13234), .B2(n13270), .C1(
        n13233), .C2(n14699), .ZN(P2_U2982) );
  INV_X1 U16577 ( .A(n13119), .ZN(n13297) );
  NAND2_X1 U16578 ( .A1(n13615), .A2(n13236), .ZN(n13298) );
  NOR2_X2 U16579 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21586) );
  AND2_X1 U16580 ( .A1(n21586), .A2(n13237), .ZN(n15611) );
  AOI21_X1 U16581 ( .B1(n15389), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n15611), 
        .ZN(n13238) );
  NAND2_X1 U16582 ( .A1(n15390), .A2(n13238), .ZN(P1_U2801) );
  AOI22_X1 U16583 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n20282), .B1(n20281), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13241) );
  NAND2_X1 U16584 ( .A1(n17488), .A2(BUF2_REG_7__SCAN_IN), .ZN(n13240) );
  NAND2_X1 U16585 ( .A1(n17490), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13239) );
  AND2_X1 U16586 ( .A1(n13240), .A2(n13239), .ZN(n20319) );
  INV_X1 U16587 ( .A(n20319), .ZN(n16814) );
  NAND2_X1 U16588 ( .A1(n20279), .A2(n16814), .ZN(n13288) );
  NAND2_X1 U16589 ( .A1(n13241), .A2(n13288), .ZN(P2_U2959) );
  AOI22_X1 U16590 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n20282), .B1(n20281), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n13244) );
  INV_X1 U16591 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n13243) );
  NAND2_X1 U16592 ( .A1(n17490), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13242) );
  OAI21_X1 U16593 ( .B1(n17490), .B2(n13243), .A(n13242), .ZN(n16824) );
  NAND2_X1 U16594 ( .A1(n20279), .A2(n16824), .ZN(n13290) );
  NAND2_X1 U16595 ( .A1(n13244), .A2(n13290), .ZN(P2_U2958) );
  AOI22_X1 U16596 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13247) );
  NAND2_X1 U16597 ( .A1(n17488), .A2(BUF2_REG_1__SCAN_IN), .ZN(n13246) );
  NAND2_X1 U16598 ( .A1(n17490), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13245) );
  AND2_X1 U16599 ( .A1(n13246), .A2(n13245), .ZN(n20225) );
  INV_X1 U16600 ( .A(n20225), .ZN(n16865) );
  NAND2_X1 U16601 ( .A1(n20279), .A2(n16865), .ZN(n13265) );
  NAND2_X1 U16602 ( .A1(n13247), .A2(n13265), .ZN(P2_U2968) );
  AOI22_X1 U16603 ( .A1(P2_UWORD_REG_9__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n13249) );
  INV_X1 U16604 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n18778) );
  NAND2_X1 U16605 ( .A1(n17490), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13248) );
  OAI21_X1 U16606 ( .B1(n17490), .B2(n18778), .A(n13248), .ZN(n16799) );
  NAND2_X1 U16607 ( .A1(n20279), .A2(n16799), .ZN(n13295) );
  NAND2_X1 U16608 ( .A1(n13249), .A2(n13295), .ZN(P2_U2961) );
  AOI22_X1 U16609 ( .A1(P2_LWORD_REG_0__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n13252) );
  NAND2_X1 U16610 ( .A1(n17488), .A2(BUF2_REG_0__SCAN_IN), .ZN(n13251) );
  NAND2_X1 U16611 ( .A1(n17490), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13250) );
  AND2_X1 U16612 ( .A1(n13251), .A2(n13250), .ZN(n20233) );
  INV_X1 U16613 ( .A(n20233), .ZN(n16874) );
  NAND2_X1 U16614 ( .A1(n20279), .A2(n16874), .ZN(n13286) );
  NAND2_X1 U16615 ( .A1(n13252), .A2(n13286), .ZN(P2_U2967) );
  AOI22_X1 U16616 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13256) );
  NAND2_X1 U16617 ( .A1(n17488), .A2(BUF2_REG_3__SCAN_IN), .ZN(n13254) );
  NAND2_X1 U16618 ( .A1(n17490), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13253) );
  AND2_X1 U16619 ( .A1(n13254), .A2(n13253), .ZN(n20302) );
  INV_X1 U16620 ( .A(n20302), .ZN(n13255) );
  NAND2_X1 U16621 ( .A1(n20279), .A2(n13255), .ZN(n13278) );
  NAND2_X1 U16622 ( .A1(n13256), .A2(n13278), .ZN(P2_U2955) );
  AOI22_X1 U16623 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13259) );
  NAND2_X1 U16624 ( .A1(n17488), .A2(BUF2_REG_5__SCAN_IN), .ZN(n13258) );
  NAND2_X1 U16625 ( .A1(n17490), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13257) );
  AND2_X1 U16626 ( .A1(n13258), .A2(n13257), .ZN(n20308) );
  INV_X1 U16627 ( .A(n20308), .ZN(n16832) );
  NAND2_X1 U16628 ( .A1(n20279), .A2(n16832), .ZN(n13276) );
  NAND2_X1 U16629 ( .A1(n13259), .A2(n13276), .ZN(P2_U2957) );
  AOI22_X1 U16630 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n13261) );
  INV_X1 U16631 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n19424) );
  NAND2_X1 U16632 ( .A1(n17490), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13260) );
  OAI21_X1 U16633 ( .B1(n17490), .B2(n19424), .A(n13260), .ZN(n16857) );
  NAND2_X1 U16634 ( .A1(n20279), .A2(n16857), .ZN(n13271) );
  NAND2_X1 U16635 ( .A1(n13261), .A2(n13271), .ZN(P2_U2954) );
  AOI22_X1 U16636 ( .A1(P2_UWORD_REG_8__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n13264) );
  INV_X1 U16637 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n13263) );
  NAND2_X1 U16638 ( .A1(n17490), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13262) );
  OAI21_X1 U16639 ( .B1(n17490), .B2(n13263), .A(n13262), .ZN(n16805) );
  NAND2_X1 U16640 ( .A1(n20279), .A2(n16805), .ZN(n13284) );
  NAND2_X1 U16641 ( .A1(n13264), .A2(n13284), .ZN(P2_U2960) );
  AOI22_X1 U16642 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13266) );
  NAND2_X1 U16643 ( .A1(n13266), .A2(n13265), .ZN(P2_U2953) );
  AOI22_X1 U16644 ( .A1(P2_UWORD_REG_13__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n13267) );
  NAND2_X1 U16645 ( .A1(n20279), .A2(n14434), .ZN(n13282) );
  NAND2_X1 U16646 ( .A1(n13267), .A2(n13282), .ZN(P2_U2965) );
  AOI22_X1 U16647 ( .A1(P2_UWORD_REG_11__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n13269) );
  NAND2_X1 U16648 ( .A1(n17490), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13268) );
  OAI21_X1 U16649 ( .B1(n17490), .B2(n18782), .A(n13268), .ZN(n16783) );
  NAND2_X1 U16650 ( .A1(n20279), .A2(n16783), .ZN(n13280) );
  NAND2_X1 U16651 ( .A1(n13269), .A2(n13280), .ZN(P2_U2963) );
  AOI22_X1 U16652 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n20282), .B1(n20281), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13272) );
  NAND2_X1 U16653 ( .A1(n13272), .A2(n13271), .ZN(P2_U2969) );
  AOI22_X1 U16654 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n20282), .B1(n20281), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13275) );
  NAND2_X1 U16655 ( .A1(n17488), .A2(BUF2_REG_4__SCAN_IN), .ZN(n13274) );
  NAND2_X1 U16656 ( .A1(n17490), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13273) );
  AND2_X1 U16657 ( .A1(n13274), .A2(n13273), .ZN(n20305) );
  INV_X1 U16658 ( .A(n20305), .ZN(n16840) );
  NAND2_X1 U16659 ( .A1(n20279), .A2(n16840), .ZN(n13292) );
  NAND2_X1 U16660 ( .A1(n13275), .A2(n13292), .ZN(P2_U2971) );
  AOI22_X1 U16661 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n20282), .B1(n20281), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13277) );
  NAND2_X1 U16662 ( .A1(n13277), .A2(n13276), .ZN(P2_U2972) );
  AOI22_X1 U16663 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n13279) );
  NAND2_X1 U16664 ( .A1(n13279), .A2(n13278), .ZN(P2_U2970) );
  AOI22_X1 U16665 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13281) );
  NAND2_X1 U16666 ( .A1(n13281), .A2(n13280), .ZN(P2_U2978) );
  AOI22_X1 U16667 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13283) );
  NAND2_X1 U16668 ( .A1(n13283), .A2(n13282), .ZN(P2_U2980) );
  AOI22_X1 U16669 ( .A1(P2_LWORD_REG_8__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n13285) );
  NAND2_X1 U16670 ( .A1(n13285), .A2(n13284), .ZN(P2_U2975) );
  AOI22_X1 U16671 ( .A1(P2_UWORD_REG_0__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n13287) );
  NAND2_X1 U16672 ( .A1(n13287), .A2(n13286), .ZN(P2_U2952) );
  AOI22_X1 U16673 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13289) );
  NAND2_X1 U16674 ( .A1(n13289), .A2(n13288), .ZN(P2_U2974) );
  AOI22_X1 U16675 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13291) );
  NAND2_X1 U16676 ( .A1(n13291), .A2(n13290), .ZN(P2_U2973) );
  AOI22_X1 U16677 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n13293) );
  NAND2_X1 U16678 ( .A1(n13293), .A2(n13292), .ZN(P2_U2956) );
  INV_X1 U16679 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n20253) );
  NAND2_X1 U16680 ( .A1(n20277), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13294) );
  OAI211_X1 U16681 ( .C1(n20253), .C2(n13296), .A(n13295), .B(n13294), .ZN(
        P2_U2976) );
  AND2_X1 U16682 ( .A1(n13298), .A2(n13297), .ZN(n13299) );
  AOI21_X1 U16683 ( .B1(n13753), .B2(n13619), .A(n13299), .ZN(n20981) );
  NAND3_X1 U16684 ( .A1(n13619), .A2(n13497), .A3(n15398), .ZN(n13300) );
  NAND2_X1 U16685 ( .A1(n13300), .A2(n21759), .ZN(n21762) );
  AND2_X1 U16686 ( .A1(n20981), .A2(n21762), .ZN(n17837) );
  NOR2_X1 U16687 ( .A1(n17837), .A2(n20982), .ZN(n20991) );
  INV_X1 U16688 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13309) );
  OAI21_X1 U16689 ( .B1(n15394), .B2(n13302), .A(n13301), .ZN(n13303) );
  MUX2_X1 U16690 ( .A(n13754), .B(n13303), .S(n13753), .Z(n13306) );
  NOR2_X1 U16691 ( .A1(n13304), .A2(n13615), .ZN(n13305) );
  OAI21_X1 U16692 ( .B1(n13306), .B2(n13305), .A(n14464), .ZN(n17839) );
  INV_X1 U16693 ( .A(n17839), .ZN(n13307) );
  NAND2_X1 U16694 ( .A1(n20991), .A2(n13307), .ZN(n13308) );
  OAI21_X1 U16695 ( .B1(n20991), .B2(n13309), .A(n13308), .ZN(P1_U3484) );
  INV_X1 U16696 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13551) );
  AOI22_X1 U16697 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13313) );
  AOI22_X1 U16698 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13312) );
  AOI22_X1 U16699 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13311) );
  INV_X1 U16700 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19419) );
  OR2_X1 U16701 ( .A1(n18545), .A2(n19419), .ZN(n13310) );
  AND4_X1 U16702 ( .A1(n13313), .A2(n13312), .A3(n13311), .A4(n13310), .ZN(
        n13321) );
  AOI22_X1 U16703 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13320) );
  AOI22_X1 U16704 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13318) );
  AOI22_X1 U16705 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13317) );
  AOI22_X1 U16706 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13316) );
  NAND2_X1 U16707 ( .A1(n17762), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13315) );
  AND4_X1 U16708 ( .A1(n13318), .A2(n13317), .A3(n13316), .A4(n13315), .ZN(
        n13319) );
  AND3_X1 U16709 ( .A1(n13321), .A2(n13320), .A3(n13319), .ZN(n13438) );
  NAND4_X1 U16710 ( .A1(n13323), .A2(n13372), .A3(n18576), .A4(n13322), .ZN(
        n13326) );
  INV_X1 U16711 ( .A(n13367), .ZN(n13324) );
  NAND2_X1 U16712 ( .A1(n13324), .A2(n19878), .ZN(n13325) );
  NAND2_X1 U16713 ( .A1(n13326), .A2(n13325), .ZN(n13431) );
  AND3_X1 U16714 ( .A1(n20031), .A2(n18681), .A3(n20038), .ZN(n13327) );
  NAND4_X1 U16715 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_2__SCAN_IN), 
        .A3(P3_EBX_REG_0__SCAN_IN), .A4(P3_EBX_REG_1__SCAN_IN), .ZN(n18578) );
  NOR2_X2 U16716 ( .A1(n18564), .A2(n18563), .ZN(n13359) );
  INV_X1 U16717 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n13328) );
  NAND3_X1 U16718 ( .A1(n13359), .A2(n18576), .A3(n13328), .ZN(n13330) );
  NOR2_X1 U16719 ( .A1(n18590), .A2(n13359), .ZN(n18565) );
  NAND2_X1 U16720 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18565), .ZN(n13329) );
  OAI211_X1 U16721 ( .C1(n13438), .C2(n18586), .A(n13330), .B(n13329), .ZN(
        P3_U2695) );
  XNOR2_X1 U16722 ( .A(n16628), .B(n13332), .ZN(n13331) );
  XNOR2_X1 U16723 ( .A(n13340), .B(n13331), .ZN(n13986) );
  NOR2_X1 U16724 ( .A1(n17181), .A2(n13986), .ZN(n13338) );
  XNOR2_X1 U16725 ( .A(n13333), .B(n13332), .ZN(n13989) );
  NAND2_X1 U16726 ( .A1(n17196), .A2(n13989), .ZN(n13335) );
  NOR2_X1 U16727 ( .A1(n20181), .A2(n20847), .ZN(n13988) );
  INV_X1 U16728 ( .A(n13988), .ZN(n13334) );
  OAI211_X1 U16729 ( .C1(n17187), .C2(n13336), .A(n13335), .B(n13334), .ZN(
        n13337) );
  AOI211_X1 U16730 ( .C1(n13336), .C2(n17190), .A(n13338), .B(n13337), .ZN(
        n13339) );
  OAI21_X1 U16731 ( .B1(n14360), .B2(n17166), .A(n13339), .ZN(P2_U3013) );
  XNOR2_X1 U16732 ( .A(n13917), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17453) );
  NOR2_X1 U16733 ( .A1(n20181), .A2(n20071), .ZN(n17460) );
  OAI21_X1 U16734 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n16641), .A(
        n13340), .ZN(n17457) );
  OAI21_X1 U16735 ( .B1(n17172), .B2(n13341), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13342) );
  OAI21_X1 U16736 ( .B1(n17457), .B2(n17181), .A(n13342), .ZN(n13343) );
  AOI211_X1 U16737 ( .C1(n17453), .C2(n17196), .A(n17460), .B(n13343), .ZN(
        n13344) );
  OAI21_X1 U16738 ( .B1(n10780), .B2(n17166), .A(n13344), .ZN(P2_U3014) );
  AOI22_X1 U16739 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13350) );
  AOI22_X1 U16740 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13349) );
  AOI22_X1 U16741 ( .A1(n17705), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17699), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13348) );
  INV_X1 U16742 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19423) );
  OR2_X1 U16743 ( .A1(n18545), .A2(n19423), .ZN(n13347) );
  AND4_X1 U16744 ( .A1(n13350), .A2(n13349), .A3(n13348), .A4(n13347), .ZN(
        n13358) );
  INV_X1 U16745 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n19643) );
  AOI22_X1 U16746 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11716), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13357) );
  AOI22_X1 U16747 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13355) );
  AOI22_X1 U16748 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13354) );
  AOI22_X1 U16749 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13353) );
  NAND2_X1 U16750 ( .A1(n17762), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13352) );
  AND4_X1 U16751 ( .A1(n13355), .A2(n13354), .A3(n13353), .A4(n13352), .ZN(
        n13356) );
  AND3_X1 U16752 ( .A1(n13358), .A2(n13357), .A3(n13356), .ZN(n13566) );
  OAI211_X1 U16753 ( .C1(n13360), .C2(P3_EBX_REG_9__SCAN_IN), .A(n18586), .B(
        n13579), .ZN(n13361) );
  OAI21_X1 U16754 ( .B1(n13566), .B2(n18586), .A(n13361), .ZN(P3_U2694) );
  INV_X1 U16755 ( .A(n20030), .ZN(n19934) );
  NOR2_X1 U16756 ( .A1(n18039), .A2(n20032), .ZN(n13364) );
  OAI21_X1 U16757 ( .B1(n18679), .B2(n13429), .A(n13364), .ZN(n13365) );
  OAI211_X1 U16758 ( .C1(n13368), .C2(n13367), .A(n13366), .B(n13365), .ZN(
        n19897) );
  INV_X1 U16759 ( .A(n19897), .ZN(n13369) );
  INV_X1 U16760 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n19401) );
  NAND3_X1 U16761 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n20015)
         );
  OR2_X1 U16762 ( .A1(n19401), .A2(n20015), .ZN(n17800) );
  NAND2_X1 U16763 ( .A1(n20035), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19415) );
  OAI211_X1 U16764 ( .C1(n19914), .C2(n13369), .A(n17800), .B(n19415), .ZN(
        n17809) );
  INV_X1 U16765 ( .A(n17809), .ZN(n13541) );
  NAND2_X1 U16766 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19283), .ZN(
        n13370) );
  AOI21_X1 U16767 ( .B1(n13373), .B2(n13370), .A(n13404), .ZN(n13376) );
  AOI21_X1 U16768 ( .B1(n9763), .B2(n13372), .A(n13371), .ZN(n13535) );
  OAI21_X1 U16769 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n13373), .A(
        n13535), .ZN(n13374) );
  INV_X1 U16770 ( .A(n13374), .ZN(n13375) );
  MUX2_X1 U16771 ( .A(n13376), .B(n9823), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13380) );
  INV_X1 U16772 ( .A(n18409), .ZN(n13530) );
  NAND2_X1 U16773 ( .A1(n13394), .A2(n14012), .ZN(n13534) );
  NAND2_X1 U16774 ( .A1(n13530), .A2(n13534), .ZN(n18424) );
  INV_X1 U16775 ( .A(n18424), .ZN(n13382) );
  INV_X1 U16776 ( .A(n13377), .ZN(n17806) );
  OAI21_X1 U16777 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n17806), .ZN(n13378) );
  OAI22_X1 U16778 ( .A1(n19382), .A2(n13382), .B1(n13529), .B2(n13378), .ZN(
        n13379) );
  NOR2_X1 U16779 ( .A1(n13380), .A2(n13379), .ZN(n19856) );
  INV_X1 U16780 ( .A(n20048), .ZN(n18442) );
  NOR2_X1 U16781 ( .A1(n18678), .A2(n13464), .ZN(n13400) );
  AOI22_X1 U16782 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n19379), .B2(n13381), .ZN(
        n13398) );
  AOI22_X1 U16783 ( .A1(n19909), .A2(n13382), .B1(n13400), .B2(n13398), .ZN(
        n13383) );
  OAI211_X1 U16784 ( .C1(n19856), .C2(n18442), .A(n17809), .B(n13383), .ZN(
        n13384) );
  INV_X1 U16785 ( .A(n13384), .ZN(n13385) );
  AOI21_X1 U16786 ( .B1(n13541), .B2(n14012), .A(n13385), .ZN(P3_U3288) );
  INV_X1 U16787 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13392) );
  AND2_X1 U16788 ( .A1(n11185), .A2(n16694), .ZN(n13386) );
  NAND2_X1 U16789 ( .A1(n14410), .A2(n13386), .ZN(n14349) );
  NAND2_X1 U16790 ( .A1(n20965), .A2(n14498), .ZN(n13388) );
  NAND2_X1 U16791 ( .A1(n20281), .A2(n20967), .ZN(n13387) );
  NAND2_X1 U16792 ( .A1(n20260), .A2(n13389), .ZN(n20235) );
  OR2_X1 U16793 ( .A1(n13390), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20962) );
  INV_X2 U16794 ( .A(n20962), .ZN(n20273) );
  AOI22_X1 U16795 ( .A1(n20273), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n20272), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13391) );
  OAI21_X1 U16796 ( .B1(n13392), .B2(n20235), .A(n13391), .ZN(P2_U2924) );
  NAND2_X1 U16797 ( .A1(n19160), .A2(n13404), .ZN(n13397) );
  NAND2_X1 U16798 ( .A1(n19306), .A2(n13433), .ZN(n13463) );
  INV_X1 U16799 ( .A(n13393), .ZN(n13395) );
  NAND2_X1 U16800 ( .A1(n13395), .A2(n13394), .ZN(n14246) );
  INV_X1 U16801 ( .A(n14246), .ZN(n13401) );
  NAND2_X1 U16802 ( .A1(n13463), .A2(n13401), .ZN(n13396) );
  NAND2_X1 U16803 ( .A1(n13397), .A2(n13396), .ZN(n19859) );
  INV_X1 U16804 ( .A(n13398), .ZN(n13399) );
  AOI22_X1 U16805 ( .A1(n19909), .A2(n13401), .B1(n13400), .B2(n13399), .ZN(
        n13402) );
  INV_X1 U16806 ( .A(n13402), .ZN(n13403) );
  AOI21_X1 U16807 ( .B1(n19859), .B2(n20048), .A(n13403), .ZN(n13405) );
  AOI22_X1 U16808 ( .A1(n17809), .A2(n13405), .B1(n13541), .B2(n13404), .ZN(
        P3_U3289) );
  AOI21_X1 U16809 ( .B1(n19341), .B2(n19160), .A(n19396), .ZN(n13412) );
  NOR2_X1 U16810 ( .A1(n13441), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13445) );
  NOR2_X1 U16811 ( .A1(n13445), .A2(n13447), .ZN(n13653) );
  INV_X1 U16812 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n13406) );
  NOR2_X1 U16813 ( .A1(n19110), .A2(n13406), .ZN(n13649) );
  NOR2_X1 U16814 ( .A1(n19876), .A2(n19283), .ZN(n19187) );
  NOR2_X1 U16815 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n19187), .ZN(
        n13407) );
  NAND2_X1 U16816 ( .A1(n19341), .A2(n13407), .ZN(n13449) );
  INV_X1 U16817 ( .A(n13449), .ZN(n13408) );
  AOI211_X1 U16818 ( .C1(n19370), .C2(n13653), .A(n13649), .B(n13408), .ZN(
        n13411) );
  INV_X1 U16819 ( .A(n19377), .ZN(n19351) );
  INV_X1 U16820 ( .A(n13653), .ZN(n13409) );
  NAND2_X1 U16821 ( .A1(n19351), .A2(n13409), .ZN(n13410) );
  OAI211_X1 U16822 ( .C1(n13412), .C2(n13464), .A(n13411), .B(n13410), .ZN(
        P3_U2862) );
  INV_X1 U16823 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14079) );
  OAI21_X1 U16824 ( .B1(n15390), .B2(n15395), .A(n13413), .ZN(n13414) );
  INV_X1 U16825 ( .A(n15398), .ZN(n17847) );
  NAND2_X1 U16826 ( .A1(n21132), .A2(n14449), .ZN(n21117) );
  INV_X2 U16827 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21641) );
  NOR2_X1 U16828 ( .A1(n21641), .A2(n13237), .ZN(n14314) );
  INV_X1 U16829 ( .A(n14314), .ZN(n17928) );
  OR2_X1 U16830 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17928), .ZN(n21142) );
  INV_X2 U16831 ( .A(n21142), .ZN(n21760) );
  NOR2_X4 U16832 ( .A1(n21132), .A2(n21760), .ZN(n13826) );
  AOI22_X1 U16833 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13415) );
  OAI21_X1 U16834 ( .B1(n14079), .B2(n21117), .A(n13415), .ZN(P1_U2913) );
  INV_X1 U16835 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U16836 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13416) );
  OAI21_X1 U16837 ( .B1(n13417), .B2(n21117), .A(n13416), .ZN(P1_U2910) );
  INV_X1 U16838 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13419) );
  AOI22_X1 U16839 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13418) );
  OAI21_X1 U16840 ( .B1(n13419), .B2(n21117), .A(n13418), .ZN(P1_U2914) );
  INV_X1 U16841 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13421) );
  AOI22_X1 U16842 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13420) );
  OAI21_X1 U16843 ( .B1(n13421), .B2(n21117), .A(n13420), .ZN(P1_U2916) );
  INV_X1 U16844 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13423) );
  AOI22_X1 U16845 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13422) );
  OAI21_X1 U16846 ( .B1(n13423), .B2(n21117), .A(n13422), .ZN(P1_U2917) );
  INV_X1 U16847 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13425) );
  AOI22_X1 U16848 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13424) );
  OAI21_X1 U16849 ( .B1(n13425), .B2(n21117), .A(n13424), .ZN(P1_U2915) );
  INV_X1 U16850 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13427) );
  AOI22_X1 U16851 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13426) );
  OAI21_X1 U16852 ( .B1(n13427), .B2(n21117), .A(n13426), .ZN(P1_U2912) );
  AOI22_X1 U16853 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13428) );
  OAI21_X1 U16854 ( .B1(n15263), .B2(n21117), .A(n13428), .ZN(P1_U2911) );
  NOR2_X1 U16855 ( .A1(n20031), .A2(n18681), .ZN(n13430) );
  INV_X1 U16856 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18768) );
  INV_X1 U16857 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18766) );
  NOR2_X1 U16858 ( .A1(n18768), .A2(n18766), .ZN(n13487) );
  AND4_X1 U16859 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n13432) );
  NAND4_X1 U16860 ( .A1(n13487), .A2(P3_EAX_REG_5__SCAN_IN), .A3(
        P3_EAX_REG_6__SCAN_IN), .A4(n13432), .ZN(n13435) );
  INV_X1 U16861 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18776) );
  OR3_X1 U16862 ( .A1(n18677), .A2(n13544), .A3(n18776), .ZN(n13437) );
  INV_X1 U16863 ( .A(n13433), .ZN(n13434) );
  AOI22_X1 U16864 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18674), .B1(n18659), .B2(
        n18776), .ZN(n13436) );
  OAI211_X1 U16865 ( .C1(n13438), .C2(n18638), .A(n13437), .B(n13436), .ZN(
        P3_U2727) );
  INV_X1 U16866 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n13564) );
  INV_X1 U16867 ( .A(n13457), .ZN(n13439) );
  OAI22_X1 U16868 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18636), .B1(n13439), .B2(
        n18766), .ZN(n13440) );
  AOI21_X1 U16869 ( .B1(n18673), .B2(n13441), .A(n13440), .ZN(n13442) );
  OAI21_X1 U16870 ( .B1(n13793), .B2(n13564), .A(n13442), .ZN(P3_U2735) );
  INV_X1 U16871 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13444) );
  INV_X1 U16872 ( .A(P2_UWORD_REG_8__SCAN_IN), .ZN(n14193) );
  INV_X1 U16873 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n13443) );
  OAI222_X1 U16874 ( .A1(n20235), .A2(n13444), .B1(n20962), .B2(n14193), .C1(
        n20271), .C2(n13443), .ZN(P2_U2927) );
  XOR2_X1 U16875 ( .A(n13445), .B(n13448), .Z(n19120) );
  INV_X1 U16876 ( .A(n19370), .ZN(n19343) );
  OAI21_X1 U16877 ( .B1(n13448), .B2(n13447), .A(n13446), .ZN(n19117) );
  INV_X1 U16878 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n20018) );
  OAI22_X1 U16879 ( .A1(n19343), .A2(n19117), .B1(n20018), .B2(n19110), .ZN(
        n13454) );
  NAND2_X1 U16880 ( .A1(n19360), .A2(n13449), .ZN(n13452) );
  NOR2_X1 U16881 ( .A1(n19160), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13450) );
  NOR2_X1 U16882 ( .A1(n19361), .A2(n13450), .ZN(n13451) );
  MUX2_X1 U16883 ( .A(n13452), .B(n13451), .S(n19379), .Z(n13453) );
  AOI211_X1 U16884 ( .C1(n19120), .C2(n19351), .A(n13454), .B(n13453), .ZN(
        n13455) );
  INV_X1 U16885 ( .A(n13455), .ZN(P3_U2861) );
  INV_X1 U16886 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n18024) );
  INV_X1 U16887 ( .A(P2_UWORD_REG_14__SCAN_IN), .ZN(n14179) );
  OAI222_X1 U16888 ( .A1(n20271), .A2(n18024), .B1(n20235), .B2(n13456), .C1(
        n14179), .C2(n20962), .ZN(P2_U2921) );
  INV_X1 U16889 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n13462) );
  AOI22_X1 U16890 ( .A1(n18673), .A2(n13458), .B1(n13457), .B2(
        P3_EAX_REG_1__SCAN_IN), .ZN(n13461) );
  INV_X1 U16891 ( .A(n13487), .ZN(n13459) );
  OAI211_X1 U16892 ( .C1(P3_EAX_REG_0__SCAN_IN), .C2(P3_EAX_REG_1__SCAN_IN), 
        .A(n13488), .B(n13459), .ZN(n13460) );
  OAI211_X1 U16893 ( .C1(n13793), .C2(n13462), .A(n13461), .B(n13460), .ZN(
        P3_U2734) );
  MUX2_X1 U16894 ( .A(n19160), .B(n13463), .S(n11687), .Z(n19861) );
  AOI22_X1 U16895 ( .A1(n19861), .A2(n20048), .B1(P3_STATE2_REG_1__SCAN_IN), 
        .B2(n13464), .ZN(n13465) );
  AOI22_X1 U16896 ( .A1(n17809), .A2(n13465), .B1(n13541), .B2(n11687), .ZN(
        n13467) );
  INV_X1 U16897 ( .A(n19909), .ZN(n13531) );
  NOR3_X1 U16898 ( .A1(n13531), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        n13541), .ZN(n13466) );
  OR2_X1 U16899 ( .A1(n13467), .A2(n13466), .ZN(P3_U3290) );
  AOI22_X1 U16900 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11716), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13476) );
  INV_X1 U16901 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13470) );
  NAND2_X1 U16902 ( .A1(n17762), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13469) );
  NAND2_X1 U16903 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n13468) );
  OAI211_X1 U16904 ( .C1(n9756), .C2(n13470), .A(n13469), .B(n13468), .ZN(
        n13471) );
  INV_X1 U16905 ( .A(n13471), .ZN(n13475) );
  AOI22_X1 U16906 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13474) );
  AOI22_X1 U16907 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13473) );
  NAND4_X1 U16908 ( .A1(n13476), .A2(n13475), .A3(n13474), .A4(n13473), .ZN(
        n13482) );
  AOI22_X1 U16909 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13480) );
  AOI22_X1 U16910 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13479) );
  AOI22_X1 U16911 ( .A1(n17705), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13478) );
  INV_X1 U16912 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19429) );
  OR2_X1 U16913 ( .A1(n18545), .A2(n19429), .ZN(n13477) );
  NAND4_X1 U16914 ( .A1(n13480), .A2(n13479), .A3(n13478), .A4(n13477), .ZN(
        n13481) );
  OR2_X1 U16915 ( .A1(n13482), .A2(n13481), .ZN(n18672) );
  NOR3_X1 U16916 ( .A1(n19448), .A2(n13579), .A3(P3_EBX_REG_10__SCAN_IN), .ZN(
        n13485) );
  INV_X1 U16917 ( .A(n13579), .ZN(n13483) );
  INV_X1 U16918 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n18317) );
  NOR3_X1 U16919 ( .A1(n18590), .A2(n13483), .A3(n18317), .ZN(n13484) );
  AOI211_X1 U16920 ( .C1(n18590), .C2(n18672), .A(n13485), .B(n13484), .ZN(
        n13486) );
  INV_X1 U16921 ( .A(n13486), .ZN(P3_U2693) );
  NAND3_X1 U16922 ( .A1(n13488), .A2(P3_EAX_REG_2__SCAN_IN), .A3(n13487), .ZN(
        n13513) );
  INV_X1 U16923 ( .A(n13513), .ZN(n13512) );
  AOI22_X1 U16924 ( .A1(n13488), .A2(n13487), .B1(P3_EAX_REG_2__SCAN_IN), .B2(
        n18662), .ZN(n13489) );
  OAI222_X1 U16925 ( .A1(n13793), .A2(n19424), .B1(n13512), .B2(n13489), .C1(
        n18638), .C2(n12079), .ZN(P3_U2733) );
  OR2_X1 U16926 ( .A1(n13490), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13492) );
  AND2_X1 U16927 ( .A1(n13492), .A2(n13491), .ZN(n15786) );
  INV_X1 U16928 ( .A(n15786), .ZN(n21173) );
  AND2_X1 U16929 ( .A1(n13754), .A2(n13618), .ZN(n13493) );
  NAND2_X1 U16930 ( .A1(n13753), .A2(n13493), .ZN(n13499) );
  NOR2_X1 U16931 ( .A1(n14464), .A2(n20982), .ZN(n13494) );
  NAND4_X1 U16932 ( .A1(n13496), .A2(n13495), .A3(n13494), .A4(n12632), .ZN(
        n13620) );
  NAND2_X1 U16933 ( .A1(n14665), .A2(n13500), .ZN(n13501) );
  NAND2_X1 U16934 ( .A1(n13501), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13508) );
  INV_X1 U16935 ( .A(n13508), .ZN(n13509) );
  INV_X1 U16936 ( .A(n14325), .ZN(n14554) );
  INV_X1 U16937 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13503) );
  NAND2_X1 U16938 ( .A1(n21641), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13505) );
  NAND2_X1 U16939 ( .A1(n15379), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n13504) );
  OAI211_X1 U16940 ( .C1(n14554), .C2(n13503), .A(n13505), .B(n13504), .ZN(
        n13506) );
  AOI21_X1 U16941 ( .B1(n13502), .B2(n15043), .A(n13506), .ZN(n13507) );
  INV_X1 U16942 ( .A(n13507), .ZN(n13685) );
  OR2_X1 U16943 ( .A1(n13508), .A2(n13507), .ZN(n13687) );
  OAI21_X1 U16944 ( .B1(n13509), .B2(n13685), .A(n13687), .ZN(n15793) );
  INV_X2 U16945 ( .A(n21112), .ZN(n15817) );
  OAI222_X1 U16946 ( .A1(n21173), .A2(n15821), .B1(n21116), .B2(n13510), .C1(
        n15793), .C2(n15817), .ZN(P1_U2872) );
  INV_X1 U16947 ( .A(n13511), .ZN(n13515) );
  INV_X1 U16948 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n19430) );
  AOI21_X1 U16949 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n18662), .A(n13512), .ZN(
        n13514) );
  INV_X1 U16950 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18731) );
  NOR2_X1 U16951 ( .A1(n18731), .A2(n13513), .ZN(n13607) );
  OAI222_X1 U16952 ( .A1(n18638), .A2(n13515), .B1(n13793), .B2(n19430), .C1(
        n13514), .C2(n13607), .ZN(P3_U2732) );
  NAND3_X1 U16953 ( .A1(n21638), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17927) );
  INV_X1 U16954 ( .A(n17927), .ZN(n13516) );
  OAI211_X1 U16955 ( .C1(n14665), .C2(n13518), .A(n13517), .B(n13765), .ZN(
        n13520) );
  NAND2_X1 U16956 ( .A1(n13520), .A2(n13519), .ZN(n21176) );
  OR2_X1 U16957 ( .A1(n12588), .A2(n20982), .ZN(n13521) );
  INV_X1 U16958 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13522) );
  OR2_X1 U16959 ( .A1(n17899), .A2(n13522), .ZN(n21182) );
  NAND2_X1 U16960 ( .A1(n21584), .A2(n13523), .ZN(n21758) );
  NAND2_X1 U16961 ( .A1(n21758), .A2(n21638), .ZN(n13524) );
  NAND2_X1 U16962 ( .A1(n21638), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17849) );
  NAND2_X1 U16963 ( .A1(n21426), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13525) );
  NAND2_X1 U16964 ( .A1(n17849), .A2(n13525), .ZN(n13714) );
  OAI21_X1 U16965 ( .B1(n17870), .B2(n13714), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13526) );
  OAI211_X1 U16966 ( .C1(n21176), .C2(n20989), .A(n21182), .B(n13526), .ZN(
        n13527) );
  INV_X1 U16967 ( .A(n13527), .ZN(n13528) );
  OAI21_X1 U16968 ( .B1(n15793), .B2(n16117), .A(n13528), .ZN(P1_U2999) );
  AOI221_X1 U16969 ( .B1(n13534), .B2(n19876), .C1(n13529), .C2(n19160), .A(
        n18409), .ZN(n19893) );
  NOR3_X1 U16970 ( .A1(n19893), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n18442), .ZN(n13533) );
  NOR3_X1 U16971 ( .A1(n13531), .A2(n18524), .A3(n13530), .ZN(n13532) );
  NOR2_X1 U16972 ( .A1(n13533), .A2(n13532), .ZN(n13542) );
  OAI21_X1 U16973 ( .B1(n13535), .B2(n18409), .A(n13534), .ZN(n13536) );
  AOI21_X1 U16974 ( .B1(n19160), .B2(n13537), .A(n13536), .ZN(n19894) );
  NOR2_X1 U16975 ( .A1(n19894), .A2(n18442), .ZN(n13538) );
  AOI211_X1 U16976 ( .C1(n19909), .C2(n18541), .A(n13541), .B(n13538), .ZN(
        n13540) );
  OAI22_X1 U16977 ( .A1(n13542), .A2(n13541), .B1(n13540), .B2(n13539), .ZN(
        P3_U3285) );
  NOR2_X2 U16978 ( .A1(n18662), .A2(n19440), .ZN(n18648) );
  INV_X1 U16979 ( .A(n18648), .ZN(n18658) );
  INV_X1 U16980 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18794) );
  NAND3_X1 U16981 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .A3(P3_EAX_REG_9__SCAN_IN), .ZN(n13593) );
  NAND4_X1 U16982 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(P3_EAX_REG_14__SCAN_IN), .A4(P3_EAX_REG_13__SCAN_IN), .ZN(n13543)
         );
  NOR2_X1 U16983 ( .A1(n13593), .A2(n13543), .ZN(n18660) );
  NAND2_X1 U16984 ( .A1(n13544), .A2(n18660), .ZN(n18661) );
  OAI211_X1 U16985 ( .C1(n13545), .C2(P3_EAX_REG_16__SCAN_IN), .A(n18594), .B(
        n18662), .ZN(n13563) );
  NOR2_X2 U16986 ( .A1(n18662), .A2(n13546), .ZN(n18653) );
  INV_X1 U16987 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13548) );
  OAI22_X1 U16988 ( .A1(n18464), .A2(n13548), .B1(n17767), .B2(n13547), .ZN(
        n13549) );
  AOI21_X1 U16989 ( .B1(n9867), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(n13549), .ZN(n13561) );
  INV_X1 U16990 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13550) );
  OAI22_X1 U16991 ( .A1(n13551), .A2(n18539), .B1(n18541), .B2(n13550), .ZN(
        n13557) );
  AOI22_X1 U16992 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13555) );
  AOI22_X1 U16993 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13554) );
  AOI22_X1 U16994 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13553) );
  NAND2_X1 U16995 ( .A1(n11944), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n13552) );
  NAND4_X1 U16996 ( .A1(n13555), .A2(n13554), .A3(n13553), .A4(n13552), .ZN(
        n13556) );
  NOR2_X1 U16997 ( .A1(n13557), .A2(n13556), .ZN(n13560) );
  AOI22_X1 U16998 ( .A1(n17705), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13559) );
  AOI22_X1 U16999 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13558) );
  NAND4_X1 U17000 ( .A1(n13561), .A2(n13560), .A3(n13559), .A4(n13558), .ZN(
        n13891) );
  AOI22_X1 U17001 ( .A1(n18653), .A2(BUF2_REG_16__SCAN_IN), .B1(n18673), .B2(
        n13891), .ZN(n13562) );
  OAI211_X1 U17002 ( .C1(n18658), .C2(n13564), .A(n13563), .B(n13562), .ZN(
        P3_U2719) );
  INV_X1 U17003 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18720) );
  NAND2_X1 U17004 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18659), .ZN(n13592) );
  NOR2_X1 U17005 ( .A1(n18720), .A2(n13592), .ZN(n18671) );
  INV_X1 U17006 ( .A(n13592), .ZN(n13565) );
  AOI21_X1 U17007 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n18662), .A(n13565), .ZN(
        n13567) );
  OAI222_X1 U17008 ( .A1(n18778), .A2(n13793), .B1(n18671), .B2(n13567), .C1(
        n18638), .C2(n13566), .ZN(P3_U2726) );
  AOI22_X1 U17009 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13571) );
  AOI22_X1 U17010 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13570) );
  AOI22_X1 U17011 ( .A1(n17705), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17699), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13569) );
  INV_X1 U17012 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19434) );
  OR2_X1 U17013 ( .A1(n18545), .A2(n19434), .ZN(n13568) );
  AND4_X1 U17014 ( .A1(n13571), .A2(n13570), .A3(n13569), .A4(n13568), .ZN(
        n13578) );
  AOI22_X1 U17015 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13577) );
  AOI22_X1 U17016 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13575) );
  AOI22_X1 U17017 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13574) );
  AOI22_X1 U17018 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13573) );
  NAND2_X1 U17019 ( .A1(n17762), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13572) );
  AND4_X1 U17020 ( .A1(n13575), .A2(n13574), .A3(n13573), .A4(n13572), .ZN(
        n13576) );
  AND3_X1 U17021 ( .A1(n13578), .A2(n13577), .A3(n13576), .ZN(n13629) );
  INV_X1 U17022 ( .A(n13720), .ZN(n13580) );
  OAI211_X1 U17023 ( .C1(n9860), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18586), .B(
        n13580), .ZN(n13581) );
  OAI21_X1 U17024 ( .B1(n13629), .B2(n18586), .A(n13581), .ZN(P3_U2692) );
  XNOR2_X1 U17025 ( .A(n13583), .B(n13582), .ZN(n13717) );
  INV_X1 U17026 ( .A(n13717), .ZN(n13591) );
  OAI21_X1 U17027 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n16297), .A(
        n16296), .ZN(n21179) );
  INV_X1 U17028 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21660) );
  NOR2_X1 U17029 ( .A1(n17899), .A2(n21660), .ZN(n13716) );
  OAI21_X1 U17030 ( .B1(n13585), .B2(n13610), .A(n13584), .ZN(n15782) );
  INV_X1 U17031 ( .A(n15782), .ZN(n13586) );
  NOR2_X1 U17032 ( .A1(n21174), .A2(n13586), .ZN(n13587) );
  AOI211_X1 U17033 ( .C1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n21179), .A(
        n13716), .B(n13587), .ZN(n13590) );
  NOR2_X1 U17034 ( .A1(n21180), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13799) );
  INV_X1 U17035 ( .A(n13799), .ZN(n13588) );
  NAND3_X1 U17036 ( .A1(n16259), .A2(n13582), .A3(n13588), .ZN(n13589) );
  OAI211_X1 U17037 ( .C1(n13591), .C2(n21175), .A(n13590), .B(n13589), .ZN(
        P1_U3030) );
  INV_X1 U17038 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n18784) );
  NOR2_X1 U17039 ( .A1(n13593), .A2(n13592), .ZN(n13627) );
  AOI21_X1 U17040 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18662), .A(n13627), .ZN(
        n13606) );
  AOI22_X1 U17041 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13598) );
  AOI22_X1 U17042 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13597) );
  AOI22_X1 U17043 ( .A1(n17705), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13596) );
  INV_X1 U17044 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13594) );
  OR2_X1 U17045 ( .A1(n18545), .A2(n13594), .ZN(n13595) );
  AND4_X1 U17046 ( .A1(n13598), .A2(n13597), .A3(n13596), .A4(n13595), .ZN(
        n13605) );
  AOI22_X1 U17047 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13604) );
  AOI22_X1 U17048 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13602) );
  INV_X1 U17049 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14065) );
  AOI22_X1 U17050 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13601) );
  AOI22_X1 U17051 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13600) );
  NAND2_X1 U17052 ( .A1(n17762), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n13599) );
  AND4_X1 U17053 ( .A1(n13602), .A2(n13601), .A3(n13600), .A4(n13599), .ZN(
        n13603) );
  AND3_X1 U17054 ( .A1(n13605), .A2(n13604), .A3(n13603), .ZN(n13648) );
  OAI222_X1 U17055 ( .A1(n13793), .A2(n18784), .B1(n13711), .B2(n13606), .C1(
        n18638), .C2(n13648), .ZN(P3_U2723) );
  INV_X1 U17056 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n19435) );
  NAND2_X1 U17057 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n13607), .ZN(n13695) );
  INV_X1 U17058 ( .A(n13695), .ZN(n13694) );
  AOI21_X1 U17059 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n18662), .A(n13607), .ZN(
        n13609) );
  OAI222_X1 U17060 ( .A1(n13793), .A2(n19435), .B1(n13694), .B2(n13609), .C1(
        n18638), .C2(n13608), .ZN(P3_U2731) );
  NAND2_X1 U17061 ( .A1(n13611), .A2(n13610), .ZN(n13613) );
  NAND2_X1 U17062 ( .A1(n13612), .A2(n15772), .ZN(n13742) );
  INV_X1 U17063 ( .A(n12977), .ZN(n14306) );
  NAND3_X1 U17064 ( .A1(n13615), .A2(n14306), .A3(n21759), .ZN(n13616) );
  NAND2_X1 U17065 ( .A1(n12635), .A2(n14464), .ZN(n13623) );
  NAND2_X2 U17066 ( .A1(n15899), .A2(n13623), .ZN(n15897) );
  INV_X1 U17067 ( .A(DATAI_0_), .ZN(n13624) );
  OR2_X1 U17068 ( .A1(n15837), .A2(n13624), .ZN(n13626) );
  NAND2_X1 U17069 ( .A1(n15837), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13625) );
  NAND2_X1 U17070 ( .A1(n13626), .A2(n13625), .ZN(n15874) );
  INV_X1 U17071 ( .A(n15874), .ZN(n14445) );
  INV_X1 U17072 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n21152) );
  OAI222_X1 U17073 ( .A1(n15793), .A2(n15897), .B1(n15901), .B2(n14445), .C1(
        n15899), .C2(n21152), .ZN(P1_U2904) );
  INV_X1 U17074 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n18782) );
  AOI22_X1 U17075 ( .A1(n18671), .A2(P3_EAX_REG_10__SCAN_IN), .B1(
        P3_EAX_REG_11__SCAN_IN), .B2(n18662), .ZN(n13628) );
  OAI222_X1 U17076 ( .A1(n13793), .A2(n18782), .B1(n18638), .B2(n13629), .C1(
        n13628), .C2(n13627), .ZN(P3_U2724) );
  AOI22_X1 U17077 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13634) );
  AOI22_X1 U17078 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13633) );
  AOI22_X1 U17079 ( .A1(n17705), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17699), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13632) );
  INV_X1 U17080 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13630) );
  OR2_X1 U17081 ( .A1(n18545), .A2(n13630), .ZN(n13631) );
  AND4_X1 U17082 ( .A1(n13634), .A2(n13633), .A3(n13632), .A4(n13631), .ZN(
        n13641) );
  AOI22_X1 U17083 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13640) );
  AOI22_X1 U17084 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13638) );
  AOI22_X1 U17085 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13637) );
  AOI22_X1 U17086 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13636) );
  NAND2_X1 U17087 ( .A1(n11944), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n13635) );
  AND4_X1 U17088 ( .A1(n13638), .A2(n13637), .A3(n13636), .A4(n13635), .ZN(
        n13639) );
  AND3_X1 U17089 ( .A1(n13641), .A2(n13640), .A3(n13639), .ZN(n14489) );
  INV_X1 U17090 ( .A(n18594), .ZN(n13642) );
  INV_X1 U17091 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18749) );
  NOR3_X1 U17092 ( .A1(n18677), .A2(n13836), .A3(n18749), .ZN(n13643) );
  AOI21_X1 U17093 ( .B1(n13836), .B2(n18749), .A(n13643), .ZN(n13645) );
  AOI22_X1 U17094 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n18653), .B1(n18648), .B2(
        BUF2_REG_1__SCAN_IN), .ZN(n13644) );
  OAI211_X1 U17095 ( .C1(n14489), .C2(n18638), .A(n13645), .B(n13644), .ZN(
        P3_U2718) );
  NAND2_X1 U17096 ( .A1(n18576), .A2(n13720), .ZN(n13786) );
  NAND3_X1 U17097 ( .A1(n18586), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n13786), 
        .ZN(n13647) );
  OR2_X1 U17098 ( .A1(n13786), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n13646) );
  OAI211_X1 U17099 ( .C1(n18586), .C2(n13648), .A(n13647), .B(n13646), .ZN(
        P3_U2691) );
  NAND3_X1 U17100 ( .A1(n18678), .A2(n18969), .A3(n19116), .ZN(n13650) );
  AOI21_X1 U17101 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n13650), .A(
        n13649), .ZN(n13652) );
  NAND2_X1 U17102 ( .A1(n19119), .A2(n13653), .ZN(n13651) );
  OAI211_X1 U17103 ( .C1(n19112), .C2(n13653), .A(n13652), .B(n13651), .ZN(
        P3_U2830) );
  INV_X1 U17104 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n16849) );
  AOI22_X1 U17105 ( .A1(n20273), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n20240), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13654) );
  OAI21_X1 U17106 ( .B1(n16849), .B2(n20235), .A(n13654), .ZN(P2_U2932) );
  INV_X1 U17107 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n14057) );
  AOI22_X1 U17108 ( .A1(n20273), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n20240), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13655) );
  OAI21_X1 U17109 ( .B1(n14057), .B2(n20235), .A(n13655), .ZN(P2_U2928) );
  INV_X1 U17110 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13657) );
  AOI22_X1 U17111 ( .A1(n20273), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n20240), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13656) );
  OAI21_X1 U17112 ( .B1(n13657), .B2(n20235), .A(n13656), .ZN(P2_U2934) );
  INV_X1 U17113 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13659) );
  AOI22_X1 U17114 ( .A1(n20273), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n20240), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13658) );
  OAI21_X1 U17115 ( .B1(n13659), .B2(n20235), .A(n13658), .ZN(P2_U2931) );
  INV_X1 U17116 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13661) );
  AOI22_X1 U17117 ( .A1(n20273), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n20240), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13660) );
  OAI21_X1 U17118 ( .B1(n13661), .B2(n20235), .A(n13660), .ZN(P2_U2933) );
  INV_X1 U17119 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13663) );
  AOI22_X1 U17120 ( .A1(n20273), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n20240), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13662) );
  OAI21_X1 U17121 ( .B1(n13663), .B2(n20235), .A(n13662), .ZN(P2_U2929) );
  INV_X1 U17122 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13665) );
  AOI22_X1 U17123 ( .A1(n20273), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n20240), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13664) );
  OAI21_X1 U17124 ( .B1(n13665), .B2(n20235), .A(n13664), .ZN(P2_U2922) );
  INV_X1 U17125 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13667) );
  AOI22_X1 U17126 ( .A1(n20273), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n20240), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13666) );
  OAI21_X1 U17127 ( .B1(n13667), .B2(n20235), .A(n13666), .ZN(P2_U2935) );
  INV_X1 U17128 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13669) );
  AOI22_X1 U17129 ( .A1(n20273), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n20240), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13668) );
  OAI21_X1 U17130 ( .B1(n13669), .B2(n20235), .A(n13668), .ZN(P2_U2926) );
  INV_X1 U17131 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13671) );
  AOI22_X1 U17132 ( .A1(n20273), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n20240), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13670) );
  OAI21_X1 U17133 ( .B1(n13671), .B2(n20235), .A(n13670), .ZN(P2_U2930) );
  AOI22_X1 U17134 ( .A1(n20273), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n20240), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13672) );
  OAI21_X1 U17135 ( .B1(n13673), .B2(n20235), .A(n13672), .ZN(P2_U2925) );
  NOR2_X1 U17136 ( .A1(n21761), .A2(n21759), .ZN(n13674) );
  OR2_X2 U17137 ( .A1(n15390), .A2(n13674), .ZN(n21169) );
  OR2_X1 U17138 ( .A1(n21169), .A2(n15395), .ZN(n13933) );
  INV_X1 U17139 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n21124) );
  INV_X1 U17140 ( .A(n21161), .ZN(n13678) );
  NOR2_X1 U17141 ( .A1(n14436), .A2(n13675), .ZN(n13676) );
  AOI21_X1 U17142 ( .B1(DATAI_15_), .B2(n14436), .A(n13676), .ZN(n15879) );
  INV_X1 U17143 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13677) );
  OAI222_X1 U17144 ( .A1(n13933), .A2(n21124), .B1(n13678), .B2(n15879), .C1(
        n13677), .C2(n13853), .ZN(P1_U2967) );
  NAND2_X1 U17145 ( .A1(n14438), .A2(n15043), .ZN(n13684) );
  INV_X1 U17146 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n13681) );
  INV_X1 U17147 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15778) );
  OAI22_X1 U17148 ( .A1(n15329), .A2(n13681), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15778), .ZN(n13682) );
  AOI21_X1 U17149 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n14325), .A(
        n13682), .ZN(n13683) );
  NAND2_X1 U17150 ( .A1(n13684), .A2(n13683), .ZN(n13689) );
  NOR2_X1 U17151 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13878) );
  OR2_X1 U17152 ( .A1(n13685), .A2(n15565), .ZN(n13686) );
  OAI21_X1 U17153 ( .B1(n13689), .B2(n13688), .A(n13885), .ZN(n15785) );
  AOI22_X1 U17154 ( .A1(n21111), .A2(n15782), .B1(n15818), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13690) );
  OAI21_X1 U17155 ( .B1(n15785), .B2(n15817), .A(n13690), .ZN(P1_U2871) );
  INV_X1 U17156 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n19439) );
  AOI21_X1 U17157 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n18662), .A(n13694), .ZN(
        n13692) );
  INV_X1 U17158 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18727) );
  NOR2_X1 U17159 ( .A1(n18727), .A2(n13695), .ZN(n13691) );
  OAI222_X1 U17160 ( .A1(n18638), .A2(n13693), .B1(n13793), .B2(n19439), .C1(
        n13692), .C2(n13691), .ZN(P3_U2730) );
  AOI22_X1 U17161 ( .A1(n13694), .A2(P3_EAX_REG_5__SCAN_IN), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n18662), .ZN(n13697) );
  NAND2_X1 U17162 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .ZN(n13696) );
  NOR2_X1 U17163 ( .A1(n13696), .A2(n13695), .ZN(n13791) );
  OAI222_X1 U17164 ( .A1(n18638), .A2(n13698), .B1(n13793), .B2(n13243), .C1(
        n13697), .C2(n13791), .ZN(P3_U2729) );
  INV_X1 U17165 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n19655) );
  OAI22_X1 U17166 ( .A1(n19655), .A2(n18539), .B1(n18541), .B2(n18518), .ZN(
        n13710) );
  AOI22_X1 U17167 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13703) );
  AOI22_X1 U17168 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13702) );
  AOI22_X1 U17169 ( .A1(n17705), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17699), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13701) );
  INV_X1 U17170 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13699) );
  OR2_X1 U17171 ( .A1(n18545), .A2(n13699), .ZN(n13700) );
  NAND4_X1 U17172 ( .A1(n13703), .A2(n13702), .A3(n13701), .A4(n13700), .ZN(
        n13709) );
  AOI22_X1 U17173 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13707) );
  AOI22_X1 U17174 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13706) );
  AOI22_X1 U17175 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13705) );
  NAND2_X1 U17176 ( .A1(n11944), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n13704) );
  NAND4_X1 U17177 ( .A1(n13707), .A2(n13706), .A3(n13705), .A4(n13704), .ZN(
        n13708) );
  NOR3_X1 U17178 ( .A1(n13710), .A2(n13709), .A3(n13708), .ZN(n13788) );
  AOI21_X1 U17179 ( .B1(n18662), .B2(P3_EAX_REG_13__SCAN_IN), .A(n13711), .ZN(
        n13713) );
  NAND2_X1 U17180 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n13711), .ZN(n18670) );
  INV_X1 U17181 ( .A(n18670), .ZN(n13712) );
  OAI222_X1 U17182 ( .A1(n18638), .A2(n13788), .B1(n13793), .B2(n12209), .C1(
        n13713), .C2(n13712), .ZN(P3_U2722) );
  NOR2_X1 U17183 ( .A1(n17885), .A2(n15778), .ZN(n13715) );
  AOI211_X1 U17184 ( .C1(n17880), .C2(n15778), .A(n13716), .B(n13715), .ZN(
        n13719) );
  INV_X1 U17185 ( .A(n20989), .ZN(n17883) );
  NAND2_X1 U17186 ( .A1(n13717), .A2(n17883), .ZN(n13718) );
  OAI211_X1 U17187 ( .C1(n15785), .C2(n16117), .A(n13719), .B(n13718), .ZN(
        P1_U2998) );
  INV_X1 U17188 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n18258) );
  INV_X1 U17189 ( .A(n13721), .ZN(n13722) );
  OAI21_X1 U17190 ( .B1(n13722), .B2(P3_EBX_REG_15__SCAN_IN), .A(n18586), .ZN(
        n13735) );
  INV_X1 U17191 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13723) );
  OAI22_X1 U17192 ( .A1(n13723), .A2(n18541), .B1(n18539), .B2(n17727), .ZN(
        n13734) );
  AOI22_X1 U17193 ( .A1(n17762), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11725), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13727) );
  AOI22_X1 U17194 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n17774), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13726) );
  AOI22_X1 U17195 ( .A1(n9690), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13725) );
  OR2_X1 U17196 ( .A1(n18545), .A2(n19453), .ZN(n13724) );
  NAND4_X1 U17197 ( .A1(n13727), .A2(n13726), .A3(n13725), .A4(n13724), .ZN(
        n13733) );
  AOI22_X1 U17198 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17782), .B1(
        n17705), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13731) );
  AOI22_X1 U17199 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13730) );
  AOI22_X1 U17200 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13729) );
  NAND2_X1 U17201 ( .A1(n13472), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n13728) );
  NAND4_X1 U17202 ( .A1(n13731), .A2(n13730), .A3(n13729), .A4(n13728), .ZN(
        n13732) );
  NOR3_X1 U17203 ( .A1(n13734), .A2(n13733), .A3(n13732), .ZN(n18663) );
  OAI22_X1 U17204 ( .A1(n13890), .A2(n13735), .B1(n18663), .B2(n18586), .ZN(
        P3_U2688) );
  INV_X1 U17205 ( .A(n21391), .ZN(n21192) );
  AND3_X1 U17206 ( .A1(n12962), .A2(n13737), .A3(n13736), .ZN(n13738) );
  NAND3_X1 U17207 ( .A1(n13739), .A2(n13738), .A3(n12977), .ZN(n14283) );
  AND2_X1 U17208 ( .A1(n13751), .A2(n13740), .ZN(n16349) );
  NOR2_X1 U17209 ( .A1(n14293), .A2(n13740), .ZN(n13741) );
  MUX2_X1 U17210 ( .A(n16349), .B(n13741), .S(n13745), .Z(n13747) );
  INV_X1 U17211 ( .A(n13754), .ZN(n13743) );
  NAND2_X1 U17212 ( .A1(n13743), .A2(n13742), .ZN(n14288) );
  NOR2_X1 U17213 ( .A1(n14283), .A2(n13744), .ZN(n14296) );
  XNOR2_X1 U17214 ( .A(n12518), .B(n13745), .ZN(n13749) );
  MUX2_X1 U17215 ( .A(n14288), .B(n14296), .S(n13749), .Z(n13746) );
  AOI211_X1 U17216 ( .C1(n21192), .C2(n14283), .A(n13747), .B(n13746), .ZN(
        n13748) );
  INV_X1 U17217 ( .A(n13748), .ZN(n14282) );
  AOI22_X1 U17218 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13582), .B2(n12894), .ZN(
        n16353) );
  NOR2_X1 U17219 ( .A1(n13237), .A2(n13765), .ZN(n16355) );
  INV_X1 U17220 ( .A(n14313), .ZN(n21732) );
  AOI222_X1 U17221 ( .A1(n14282), .A2(n21733), .B1(n16353), .B2(n16355), .C1(
        n21732), .C2(n13749), .ZN(n13761) );
  OAI211_X1 U17222 ( .C1(n13751), .C2(n13750), .A(n17847), .B(n21759), .ZN(
        n13752) );
  INV_X1 U17223 ( .A(n13752), .ZN(n13755) );
  MUX2_X1 U17224 ( .A(n13755), .B(n13754), .S(n13753), .Z(n13759) );
  OAI21_X1 U17225 ( .B1(n14460), .B2(n15776), .A(n13756), .ZN(n13757) );
  INV_X1 U17226 ( .A(n17825), .ZN(n14305) );
  NAND2_X1 U17227 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14314), .ZN(n17932) );
  INV_X1 U17228 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20990) );
  OAI22_X1 U17229 ( .A1(n14305), .A2(n20982), .B1(n17932), .B2(n20990), .ZN(
        n13768) );
  AOI21_X1 U17230 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21638), .A(n13768), 
        .ZN(n21736) );
  NAND2_X1 U17231 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21736), .ZN(
        n13760) );
  OAI21_X1 U17232 ( .B1(n13761), .B2(n21736), .A(n13760), .ZN(P1_U3472) );
  INV_X1 U17233 ( .A(n21736), .ZN(n16360) );
  XNOR2_X1 U17234 ( .A(n13762), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n21053) );
  NAND4_X1 U17235 ( .A1(n21053), .A2(n13768), .A3(n21733), .A4(n14306), .ZN(
        n13763) );
  OAI21_X1 U17236 ( .B1(n13764), .B2(n16360), .A(n13763), .ZN(P1_U3468) );
  AOI22_X1 U17237 ( .A1(n21732), .A2(n13503), .B1(P1_STATE2_REG_1__SCAN_IN), 
        .B2(n13765), .ZN(n13771) );
  INV_X1 U17238 ( .A(n13502), .ZN(n15789) );
  INV_X1 U17239 ( .A(n14283), .ZN(n16352) );
  MUX2_X1 U17240 ( .A(n13766), .B(n14293), .S(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n13767) );
  OAI21_X1 U17241 ( .B1(n15789), .B2(n16352), .A(n13767), .ZN(n17827) );
  NAND3_X1 U17242 ( .A1(n13768), .A2(n21733), .A3(n17827), .ZN(n13770) );
  NAND2_X1 U17243 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21736), .ZN(
        n13769) );
  OAI211_X1 U17244 ( .C1(n21736), .C2(n13771), .A(n13770), .B(n13769), .ZN(
        P1_U3474) );
  NAND2_X1 U17245 ( .A1(n13775), .A2(n13774), .ZN(n13776) );
  INV_X1 U17246 ( .A(n13778), .ZN(n14386) );
  NOR2_X1 U17247 ( .A1(n14410), .A2(n14386), .ZN(n14344) );
  NOR2_X1 U17248 ( .A1(n14363), .A2(n9937), .ZN(n14335) );
  NAND2_X1 U17249 ( .A1(n20207), .A2(n13780), .ZN(n16752) );
  INV_X1 U17250 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n16602) );
  NOR2_X1 U17251 ( .A1(n20207), .A2(n16602), .ZN(n13781) );
  AOI21_X1 U17252 ( .B1(n17446), .B2(n20207), .A(n13781), .ZN(n13782) );
  OAI21_X1 U17253 ( .B1(n20324), .B2(n16752), .A(n13782), .ZN(P2_U2884) );
  INV_X1 U17254 ( .A(DATAI_1_), .ZN(n13783) );
  OR2_X1 U17255 ( .A1(n15837), .A2(n13783), .ZN(n13785) );
  NAND2_X1 U17256 ( .A1(n15837), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13784) );
  NAND2_X1 U17257 ( .A1(n13785), .A2(n13784), .ZN(n15869) );
  INV_X1 U17258 ( .A(n15869), .ZN(n14473) );
  OAI222_X1 U17259 ( .A1(n15785), .A2(n15897), .B1(n15901), .B2(n14473), .C1(
        n15899), .C2(n13681), .ZN(P1_U2903) );
  INV_X1 U17260 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n18294) );
  NOR2_X1 U17261 ( .A1(n18294), .A2(n13786), .ZN(n13787) );
  AOI21_X1 U17262 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n18586), .A(n13787), .ZN(
        n13790) );
  NAND2_X1 U17263 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n13787), .ZN(n13825) );
  INV_X1 U17264 ( .A(n13825), .ZN(n13789) );
  OAI22_X1 U17265 ( .A1(n13790), .A2(n13789), .B1(n13788), .B2(n18586), .ZN(
        P3_U2690) );
  INV_X1 U17266 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n19446) );
  AOI21_X1 U17267 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n18662), .A(n13791), .ZN(
        n13792) );
  OAI222_X1 U17268 ( .A1(n18638), .A2(n17608), .B1(n13793), .B2(n19446), .C1(
        n13792), .C2(n18659), .ZN(P3_U2728) );
  XNOR2_X1 U17269 ( .A(n13795), .B(n13794), .ZN(n13975) );
  NAND2_X1 U17270 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13796) );
  OAI22_X1 U17271 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17886), .B1(
        n13796), .B2(n16297), .ZN(n13798) );
  OAI21_X1 U17272 ( .B1(n13798), .B2(n13797), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13807) );
  AND2_X1 U17273 ( .A1(n17906), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n13971) );
  NOR3_X1 U17274 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13582), .A3(
        n16301), .ZN(n13805) );
  NAND2_X1 U17275 ( .A1(n13802), .A2(n13801), .ZN(n13803) );
  NAND2_X1 U17276 ( .A1(n13800), .A2(n13803), .ZN(n21085) );
  OAI22_X1 U17277 ( .A1(n16297), .A2(n14541), .B1(n21174), .B2(n21085), .ZN(
        n13804) );
  NOR3_X1 U17278 ( .A1(n13971), .A2(n13805), .A3(n13804), .ZN(n13806) );
  OAI211_X1 U17279 ( .C1(n13975), .C2(n21175), .A(n13807), .B(n13806), .ZN(
        P1_U3029) );
  NAND3_X1 U17280 ( .A1(n18586), .A2(n13825), .A3(P3_EBX_REG_14__SCAN_IN), 
        .ZN(n13824) );
  AOI22_X1 U17281 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13815) );
  INV_X1 U17282 ( .A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13810) );
  NAND2_X1 U17283 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n13809) );
  NAND2_X1 U17284 ( .A1(n9690), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13808) );
  OAI211_X1 U17285 ( .C1(n9756), .C2(n13810), .A(n13809), .B(n13808), .ZN(
        n13811) );
  INV_X1 U17286 ( .A(n13811), .ZN(n13814) );
  INV_X1 U17287 ( .A(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n19514) );
  AOI22_X1 U17288 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18552), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13813) );
  AOI22_X1 U17289 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13812) );
  NAND4_X1 U17290 ( .A1(n13815), .A2(n13814), .A3(n13813), .A4(n13812), .ZN(
        n13822) );
  AOI22_X1 U17291 ( .A1(n17705), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11725), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13820) );
  AOI22_X1 U17292 ( .A1(n17762), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13819) );
  AOI22_X1 U17293 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17699), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13818) );
  INV_X1 U17294 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13816) );
  OR2_X1 U17295 ( .A1(n18545), .A2(n13816), .ZN(n13817) );
  NAND4_X1 U17296 ( .A1(n13820), .A2(n13819), .A3(n13818), .A4(n13817), .ZN(
        n13821) );
  OR2_X1 U17297 ( .A1(n13822), .A2(n13821), .ZN(n18667) );
  NAND2_X1 U17298 ( .A1(n18590), .A2(n18667), .ZN(n13823) );
  OAI211_X1 U17299 ( .C1(n13825), .C2(P3_EBX_REG_14__SCAN_IN), .A(n13824), .B(
        n13823), .ZN(P3_U2689) );
  INV_X1 U17300 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14971) );
  AOI22_X1 U17301 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13827) );
  OAI21_X1 U17302 ( .B1(n14971), .B2(n21117), .A(n13827), .ZN(P1_U2920) );
  INV_X1 U17303 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13829) );
  AOI22_X1 U17304 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13828) );
  OAI21_X1 U17305 ( .B1(n13829), .B2(n21117), .A(n13828), .ZN(P1_U2908) );
  INV_X1 U17306 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13831) );
  AOI22_X1 U17307 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13830) );
  OAI21_X1 U17308 ( .B1(n13831), .B2(n21117), .A(n13830), .ZN(P1_U2907) );
  INV_X1 U17309 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13833) );
  AOI22_X1 U17310 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13832) );
  OAI21_X1 U17311 ( .B1(n13833), .B2(n21117), .A(n13832), .ZN(P1_U2906) );
  INV_X1 U17312 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13835) );
  AOI22_X1 U17313 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13834) );
  OAI21_X1 U17314 ( .B1(n13835), .B2(n21117), .A(n13834), .ZN(P1_U2909) );
  NAND2_X1 U17315 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18655), .ZN(n18654) );
  INV_X1 U17316 ( .A(n18654), .ZN(n13837) );
  AOI21_X1 U17317 ( .B1(P3_EAX_REG_19__SCAN_IN), .B2(n18662), .A(n13837), .ZN(
        n13852) );
  NAND2_X1 U17318 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n13837), .ZN(n14530) );
  INV_X1 U17319 ( .A(n14530), .ZN(n13851) );
  INV_X1 U17320 ( .A(n18653), .ZN(n18640) );
  INV_X1 U17321 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n16848) );
  INV_X1 U17322 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17764) );
  INV_X1 U17323 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17752) );
  OAI22_X1 U17324 ( .A1(n18541), .A2(n17764), .B1(n18539), .B2(n17752), .ZN(
        n13848) );
  AOI22_X1 U17325 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13841) );
  AOI22_X1 U17326 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13840) );
  AOI22_X1 U17327 ( .A1(n17705), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17699), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13839) );
  INV_X1 U17328 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17761) );
  OR2_X1 U17329 ( .A1(n18545), .A2(n17761), .ZN(n13838) );
  NAND4_X1 U17330 ( .A1(n13841), .A2(n13840), .A3(n13839), .A4(n13838), .ZN(
        n13847) );
  AOI22_X1 U17331 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13845) );
  AOI22_X1 U17332 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13844) );
  AOI22_X1 U17333 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13843) );
  NAND2_X1 U17334 ( .A1(n11944), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n13842) );
  NAND4_X1 U17335 ( .A1(n13845), .A2(n13844), .A3(n13843), .A4(n13842), .ZN(
        n13846) );
  NOR3_X1 U17336 ( .A1(n13848), .A2(n13847), .A3(n13846), .ZN(n17547) );
  OAI22_X1 U17337 ( .A1(n18640), .A2(n16848), .B1(n17547), .B2(n18638), .ZN(
        n13849) );
  AOI21_X1 U17338 ( .B1(BUF2_REG_3__SCAN_IN), .B2(n18648), .A(n13849), .ZN(
        n13850) );
  OAI21_X1 U17339 ( .B1(n13852), .B2(n13851), .A(n13850), .ZN(P3_U2716) );
  INV_X1 U17340 ( .A(n13933), .ZN(n21155) );
  AOI22_X1 U17341 ( .A1(n21155), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n21169), .ZN(n13854) );
  MUX2_X1 U17342 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n15837), .Z(
        n15881) );
  NAND2_X1 U17343 ( .A1(n21161), .A2(n15881), .ZN(n13938) );
  NAND2_X1 U17344 ( .A1(n13854), .A2(n13938), .ZN(P1_U2966) );
  AOI22_X1 U17345 ( .A1(n21155), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n21169), .ZN(n13855) );
  MUX2_X1 U17346 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n15837), .Z(
        n15895) );
  NAND2_X1 U17347 ( .A1(n21161), .A2(n15895), .ZN(n13954) );
  NAND2_X1 U17348 ( .A1(n13855), .A2(n13954), .ZN(P1_U2961) );
  AOI22_X1 U17349 ( .A1(n21155), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n21169), .ZN(n13856) );
  MUX2_X1 U17350 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n15837), .Z(
        n15898) );
  NAND2_X1 U17351 ( .A1(n21161), .A2(n15898), .ZN(n13944) );
  NAND2_X1 U17352 ( .A1(n13856), .A2(n13944), .ZN(P1_U2960) );
  AOI22_X1 U17353 ( .A1(n21155), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n21169), .ZN(n13860) );
  INV_X1 U17354 ( .A(DATAI_7_), .ZN(n13857) );
  OR2_X1 U17355 ( .A1(n15837), .A2(n13857), .ZN(n13859) );
  NAND2_X1 U17356 ( .A1(n15837), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13858) );
  NAND2_X1 U17357 ( .A1(n13859), .A2(n13858), .ZN(n15846) );
  NAND2_X1 U17358 ( .A1(n21161), .A2(n15846), .ZN(n13942) );
  NAND2_X1 U17359 ( .A1(n13860), .A2(n13942), .ZN(P1_U2959) );
  AOI22_X1 U17360 ( .A1(n21155), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n21169), .ZN(n13864) );
  INV_X1 U17361 ( .A(DATAI_6_), .ZN(n13861) );
  OR2_X1 U17362 ( .A1(n15837), .A2(n13861), .ZN(n13863) );
  NAND2_X1 U17363 ( .A1(n15837), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13862) );
  NAND2_X1 U17364 ( .A1(n13863), .A2(n13862), .ZN(n15850) );
  NAND2_X1 U17365 ( .A1(n21161), .A2(n15850), .ZN(n13940) );
  NAND2_X1 U17366 ( .A1(n13864), .A2(n13940), .ZN(P1_U2958) );
  AOI22_X1 U17367 ( .A1(n21155), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n21169), .ZN(n13868) );
  INV_X1 U17368 ( .A(DATAI_5_), .ZN(n13865) );
  OR2_X1 U17369 ( .A1(n15837), .A2(n13865), .ZN(n13867) );
  NAND2_X1 U17370 ( .A1(n15837), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13866) );
  NAND2_X1 U17371 ( .A1(n13867), .A2(n13866), .ZN(n15853) );
  NAND2_X1 U17372 ( .A1(n21161), .A2(n15853), .ZN(n13935) );
  NAND2_X1 U17373 ( .A1(n13868), .A2(n13935), .ZN(P1_U2957) );
  AND2_X1 U17374 ( .A1(n13870), .A2(n13871), .ZN(n13872) );
  NOR2_X1 U17375 ( .A1(n13869), .A2(n13872), .ZN(n17373) );
  INV_X1 U17376 ( .A(n17373), .ZN(n20154) );
  INV_X1 U17377 ( .A(n20232), .ZN(n14625) );
  AOI22_X1 U17378 ( .A1(n14625), .A2(n16799), .B1(P2_EAX_REG_9__SCAN_IN), .B2(
        n20226), .ZN(n13874) );
  OAI21_X1 U17379 ( .B1(n20154), .B2(n14700), .A(n13874), .ZN(P2_U2910) );
  OAI21_X1 U17380 ( .B1(n13869), .B2(n13876), .A(n13875), .ZN(n20139) );
  AOI22_X1 U17381 ( .A1(n14625), .A2(n16791), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n20226), .ZN(n13877) );
  OAI21_X1 U17382 ( .B1(n20139), .B2(n14700), .A(n13877), .ZN(P2_U2909) );
  INV_X1 U17383 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n13880) );
  XNOR2_X1 U17384 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21093) );
  AOI21_X1 U17385 ( .B1(n13878), .B2(n21093), .A(n15378), .ZN(n13879) );
  OAI21_X1 U17386 ( .B1(n15329), .B2(n13880), .A(n13879), .ZN(n13881) );
  AOI21_X1 U17387 ( .B1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n14325), .A(
        n13881), .ZN(n13882) );
  NAND2_X1 U17388 ( .A1(n15378), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14320) );
  NAND2_X1 U17389 ( .A1(n13886), .A2(n13885), .ZN(n13887) );
  INV_X1 U17390 ( .A(n21097), .ZN(n13970) );
  INV_X1 U17391 ( .A(n21085), .ZN(n13888) );
  AOI22_X1 U17392 ( .A1(n21111), .A2(n13888), .B1(n15818), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13889) );
  OAI21_X1 U17393 ( .B1(n13970), .B2(n15817), .A(n13889), .ZN(P1_U2870) );
  OAI21_X1 U17394 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n13890), .A(n14485), .ZN(
        n13893) );
  NAND2_X1 U17395 ( .A1(n18590), .A2(n13891), .ZN(n13892) );
  OAI21_X1 U17396 ( .B1(n13893), .B2(n18590), .A(n13892), .ZN(P3_U2687) );
  INV_X1 U17397 ( .A(n16857), .ZN(n20299) );
  INV_X1 U17398 ( .A(n13894), .ZN(n13897) );
  INV_X1 U17399 ( .A(n13895), .ZN(n13896) );
  OR2_X1 U17400 ( .A1(n13900), .A2(n13901), .ZN(n13902) );
  NAND2_X1 U17401 ( .A1(n13903), .A2(n13902), .ZN(n20923) );
  XNOR2_X1 U17402 ( .A(n20921), .B(n20923), .ZN(n13929) );
  NAND2_X1 U17403 ( .A1(n13906), .A2(n13905), .ZN(n13907) );
  OR2_X1 U17404 ( .A1(n13909), .A2(n13908), .ZN(n13910) );
  NAND2_X1 U17405 ( .A1(n13911), .A2(n13910), .ZN(n20934) );
  NOR2_X1 U17406 ( .A1(n20931), .A2(n20934), .ZN(n13926) );
  AOI21_X1 U17407 ( .B1(n20931), .B2(n20934), .A(n13926), .ZN(n20221) );
  NAND2_X1 U17408 ( .A1(n16694), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13914) );
  AND3_X1 U17409 ( .A1(n13920), .A2(n13919), .A3(n13918), .ZN(n13923) );
  INV_X1 U17410 ( .A(n13921), .ZN(n13922) );
  NAND2_X1 U17411 ( .A1(n13923), .A2(n13922), .ZN(n13925) );
  AND2_X1 U17412 ( .A1(n13925), .A2(n13924), .ZN(n20229) );
  NAND2_X1 U17413 ( .A1(n20944), .A2(n20229), .ZN(n20228) );
  NAND2_X1 U17414 ( .A1(n20221), .A2(n20228), .ZN(n20220) );
  INV_X1 U17415 ( .A(n13926), .ZN(n13927) );
  NAND2_X1 U17416 ( .A1(n20220), .A2(n13927), .ZN(n13928) );
  NAND2_X1 U17417 ( .A1(n13928), .A2(n13929), .ZN(n16884) );
  OAI21_X1 U17418 ( .B1(n13929), .B2(n13928), .A(n16884), .ZN(n13930) );
  NAND2_X1 U17419 ( .A1(n13930), .A2(n20227), .ZN(n13932) );
  AOI22_X1 U17420 ( .A1(n12194), .A2(n20923), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n20226), .ZN(n13931) );
  OAI211_X1 U17421 ( .C1(n20232), .C2(n20299), .A(n13932), .B(n13931), .ZN(
        P2_U2917) );
  AOI22_X1 U17422 ( .A1(n21170), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n21169), .ZN(n13934) );
  NAND2_X1 U17423 ( .A1(n21161), .A2(n15874), .ZN(n13958) );
  NAND2_X1 U17424 ( .A1(n13934), .A2(n13958), .ZN(P1_U2937) );
  AOI22_X1 U17425 ( .A1(n21170), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n21169), .ZN(n13936) );
  NAND2_X1 U17426 ( .A1(n13936), .A2(n13935), .ZN(P1_U2942) );
  AOI22_X1 U17427 ( .A1(n21170), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n21169), .ZN(n13937) );
  NAND2_X1 U17428 ( .A1(n21161), .A2(n15869), .ZN(n13960) );
  NAND2_X1 U17429 ( .A1(n13937), .A2(n13960), .ZN(P1_U2938) );
  AOI22_X1 U17430 ( .A1(n21170), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n21169), .ZN(n13939) );
  NAND2_X1 U17431 ( .A1(n13939), .A2(n13938), .ZN(P1_U2951) );
  AOI22_X1 U17432 ( .A1(n21170), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n21169), .ZN(n13941) );
  NAND2_X1 U17433 ( .A1(n13941), .A2(n13940), .ZN(P1_U2943) );
  AOI22_X1 U17434 ( .A1(n21170), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n21169), .ZN(n13943) );
  NAND2_X1 U17435 ( .A1(n13943), .A2(n13942), .ZN(P1_U2944) );
  AOI22_X1 U17436 ( .A1(n21170), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n21169), .ZN(n13945) );
  NAND2_X1 U17437 ( .A1(n13945), .A2(n13944), .ZN(P1_U2945) );
  AOI22_X1 U17438 ( .A1(n21170), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n21169), .ZN(n13949) );
  INV_X1 U17439 ( .A(DATAI_3_), .ZN(n13946) );
  OR2_X1 U17440 ( .A1(n15837), .A2(n13946), .ZN(n13948) );
  NAND2_X1 U17441 ( .A1(n15837), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13947) );
  NAND2_X1 U17442 ( .A1(n13948), .A2(n13947), .ZN(n15861) );
  NAND2_X1 U17443 ( .A1(n21161), .A2(n15861), .ZN(n13962) );
  NAND2_X1 U17444 ( .A1(n13949), .A2(n13962), .ZN(P1_U2940) );
  AOI22_X1 U17445 ( .A1(n21170), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n21169), .ZN(n13953) );
  INV_X1 U17446 ( .A(DATAI_4_), .ZN(n13950) );
  OR2_X1 U17447 ( .A1(n15837), .A2(n13950), .ZN(n13952) );
  NAND2_X1 U17448 ( .A1(n15837), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13951) );
  NAND2_X1 U17449 ( .A1(n13952), .A2(n13951), .ZN(n15857) );
  NAND2_X1 U17450 ( .A1(n21161), .A2(n15857), .ZN(n13956) );
  NAND2_X1 U17451 ( .A1(n13953), .A2(n13956), .ZN(P1_U2941) );
  AOI22_X1 U17452 ( .A1(n21170), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n21169), .ZN(n13955) );
  NAND2_X1 U17453 ( .A1(n13955), .A2(n13954), .ZN(P1_U2946) );
  AOI22_X1 U17454 ( .A1(n21170), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n21169), .ZN(n13957) );
  NAND2_X1 U17455 ( .A1(n13957), .A2(n13956), .ZN(P1_U2956) );
  AOI22_X1 U17456 ( .A1(n21170), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n21169), .ZN(n13959) );
  NAND2_X1 U17457 ( .A1(n13959), .A2(n13958), .ZN(P1_U2952) );
  AOI22_X1 U17458 ( .A1(n21170), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n21169), .ZN(n13961) );
  NAND2_X1 U17459 ( .A1(n13961), .A2(n13960), .ZN(P1_U2953) );
  AOI22_X1 U17460 ( .A1(n21170), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n21169), .ZN(n13963) );
  NAND2_X1 U17461 ( .A1(n13963), .A2(n13962), .ZN(P1_U2955) );
  AOI22_X1 U17462 ( .A1(n21170), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n21169), .ZN(n13967) );
  INV_X1 U17463 ( .A(DATAI_2_), .ZN(n13964) );
  OR2_X1 U17464 ( .A1(n15837), .A2(n13964), .ZN(n13966) );
  NAND2_X1 U17465 ( .A1(n15837), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13965) );
  NAND2_X1 U17466 ( .A1(n13966), .A2(n13965), .ZN(n15865) );
  NAND2_X1 U17467 ( .A1(n21161), .A2(n15865), .ZN(n13968) );
  NAND2_X1 U17468 ( .A1(n13967), .A2(n13968), .ZN(P1_U2954) );
  AOI22_X1 U17469 ( .A1(n21170), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n21169), .ZN(n13969) );
  NAND2_X1 U17470 ( .A1(n13969), .A2(n13968), .ZN(P1_U2939) );
  INV_X1 U17471 ( .A(n15865), .ZN(n14459) );
  OAI222_X1 U17472 ( .A1(n13970), .A2(n15897), .B1(n15901), .B2(n14459), .C1(
        n15899), .C2(n13880), .ZN(P1_U2902) );
  AOI21_X1 U17473 ( .B1(n17870), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13971), .ZN(n13972) );
  OAI21_X1 U17474 ( .B1(n21093), .B2(n17877), .A(n13972), .ZN(n13973) );
  AOI21_X1 U17475 ( .B1(n21097), .B2(n17882), .A(n13973), .ZN(n13974) );
  OAI21_X1 U17476 ( .B1(n20989), .B2(n13975), .A(n13974), .ZN(P1_U2997) );
  OAI21_X1 U17477 ( .B1(n13978), .B2(n13977), .A(n13976), .ZN(n20172) );
  INV_X1 U17478 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n20257) );
  OAI222_X1 U17479 ( .A1(n20172), .A2(n14700), .B1(n20257), .B2(n16897), .C1(
        n20232), .C2(n20319), .ZN(P2_U2912) );
  XNOR2_X1 U17480 ( .A(n13979), .B(n13980), .ZN(n17408) );
  INV_X1 U17481 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n20259) );
  INV_X1 U17482 ( .A(n16824), .ZN(n20311) );
  OAI222_X1 U17483 ( .A1(n17408), .A2(n14700), .B1(n20259), .B2(n16897), .C1(
        n20232), .C2(n20311), .ZN(P2_U2913) );
  NAND2_X1 U17484 ( .A1(n13976), .A2(n13981), .ZN(n13982) );
  NAND2_X1 U17485 ( .A1(n13870), .A2(n13982), .ZN(n17380) );
  INV_X1 U17486 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n20255) );
  INV_X1 U17487 ( .A(n16805), .ZN(n13983) );
  OAI222_X1 U17488 ( .A1(n17380), .A2(n14700), .B1(n16897), .B2(n20255), .C1(
        n20232), .C2(n13983), .ZN(P2_U2911) );
  INV_X1 U17489 ( .A(n13875), .ZN(n13984) );
  OAI21_X1 U17490 ( .B1(n13984), .B2(n9864), .A(n9710), .ZN(n17347) );
  INV_X1 U17491 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n20249) );
  INV_X1 U17492 ( .A(n16783), .ZN(n13985) );
  OAI222_X1 U17493 ( .A1(n17347), .A2(n14700), .B1(n16897), .B2(n20249), .C1(
        n20232), .C2(n13985), .ZN(P2_U2908) );
  OAI22_X1 U17494 ( .A1(n14360), .A2(n17429), .B1(n17458), .B2(n13986), .ZN(
        n13987) );
  AOI211_X1 U17495 ( .C1(n17461), .C2(n20934), .A(n13988), .B(n13987), .ZN(
        n13994) );
  INV_X1 U17496 ( .A(n17451), .ZN(n14271) );
  AOI22_X1 U17497 ( .A1(n14271), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n17454), .B2(n13989), .ZN(n13993) );
  INV_X1 U17498 ( .A(n13990), .ZN(n13991) );
  OAI211_X1 U17499 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n10181), .B(n13991), .ZN(n13992) );
  NAND3_X1 U17500 ( .A1(n13994), .A2(n13993), .A3(n13992), .ZN(n14233) );
  INV_X1 U17501 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n14231) );
  NOR4_X1 U17502 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(
        P3_BYTEENABLE_REG_3__SCAN_IN), .A3(n14182), .A4(n20869), .ZN(n13995)
         );
  NAND3_X1 U17503 ( .A1(P3_BYTEENABLE_REG_2__SCAN_IN), .A2(
        P1_DATAO_REG_6__SCAN_IN), .A3(n13995), .ZN(n14007) );
  INV_X1 U17504 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13996) );
  NAND4_X1 U17505 ( .A1(n13996), .A2(n20858), .A3(BUF1_REG_20__SCAN_IN), .A4(
        DATAI_17_), .ZN(n13998) );
  INV_X1 U17506 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n13997) );
  NOR3_X1 U17507 ( .A1(n13998), .A2(P3_LWORD_REG_0__SCAN_IN), .A3(n13997), 
        .ZN(n14005) );
  INV_X1 U17508 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n17959) );
  NAND2_X1 U17509 ( .A1(n19646), .A2(n17959), .ZN(n13999) );
  NOR4_X1 U17510 ( .A1(n17672), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A3(
        P1_INSTQUEUE_REG_3__2__SCAN_IN), .A4(n13999), .ZN(n14000) );
  INV_X1 U17511 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n20243) );
  NAND4_X1 U17512 ( .A1(n14000), .A2(n20243), .A3(P3_DATAO_REG_18__SCAN_IN), 
        .A4(P2_DATAO_REG_28__SCAN_IN), .ZN(n14003) );
  INV_X1 U17513 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19967) );
  NAND4_X1 U17514 ( .A1(DATAI_23_), .A2(DATAI_27_), .A3(n14136), .A4(n19967), 
        .ZN(n14002) );
  INV_X1 U17515 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14164) );
  NAND4_X1 U17516 ( .A1(DATAI_6_), .A2(P3_DATAO_REG_2__SCAN_IN), .A3(n16158), 
        .A4(n14164), .ZN(n14001) );
  NOR3_X1 U17517 ( .A1(n14003), .A2(n14002), .A3(n14001), .ZN(n14004) );
  INV_X1 U17518 ( .A(DATAI_25_), .ZN(n14201) );
  NAND4_X1 U17519 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n14005), .A3(
        n14004), .A4(n14201), .ZN(n14006) );
  NOR4_X1 U17520 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n21666), .A3(
        n14007), .A4(n14006), .ZN(n14041) );
  NAND4_X1 U17521 ( .A1(P1_EAX_REG_4__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .A3(P2_MEMORYFETCH_REG_SCAN_IN), 
        .A4(n11589), .ZN(n14011) );
  INV_X1 U17522 ( .A(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14053) );
  NAND4_X1 U17523 ( .A1(P2_EAX_REG_23__SCAN_IN), .A2(P1_EBX_REG_23__SCAN_IN), 
        .A3(P3_UWORD_REG_4__SCAN_IN), .A4(n14053), .ZN(n14010) );
  NAND4_X1 U17524 ( .A1(P2_EAX_REG_19__SCAN_IN), .A2(P3_UWORD_REG_3__SCAN_IN), 
        .A3(n17007), .A4(n14076), .ZN(n14009) );
  NAND4_X1 U17525 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_7__4__SCAN_IN), .A3(n16246), .A4(n14067), .ZN(n14008)
         );
  NOR4_X1 U17526 ( .A1(n14011), .A2(n14010), .A3(n14009), .A4(n14008), .ZN(
        n14040) );
  INV_X1 U17527 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14152) );
  INV_X1 U17528 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n17978) );
  NAND4_X1 U17529 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_14__SCAN_IN), .A3(n14152), .A4(n17978), .ZN(n14016)
         );
  NAND4_X1 U17530 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(
        P3_EBX_REG_6__SCAN_IN), .A3(P3_ADDRESS_REG_16__SCAN_IN), .A4(n15588), 
        .ZN(n14015) );
  NAND4_X1 U17531 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), 
        .A4(P3_BE_N_REG_1__SCAN_IN), .ZN(n14014) );
  NAND4_X1 U17532 ( .A1(n14012), .A2(n16331), .A3(
        P1_INSTQUEUE_REG_14__6__SCAN_IN), .A4(P3_REIP_REG_16__SCAN_IN), .ZN(
        n14013) );
  NOR4_X1 U17533 ( .A1(n14016), .A2(n14015), .A3(n14014), .A4(n14013), .ZN(
        n14039) );
  NOR4_X1 U17534 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_REIP_REG_0__SCAN_IN), .A3(DATAI_20_), .A4(n14104), .ZN(n14020) );
  NOR4_X1 U17535 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .A3(P2_INSTQUEUE_REG_8__3__SCAN_IN), 
        .A4(n14212), .ZN(n14019) );
  INV_X1 U17536 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14178) );
  NOR4_X1 U17537 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n14178), .A3(n20856), 
        .A4(n14179), .ZN(n14018) );
  INV_X1 U17538 ( .A(P1_LWORD_REG_7__SCAN_IN), .ZN(n21138) );
  NOR4_X1 U17539 ( .A1(BUF2_REG_16__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(n14193), .A4(n21138), .ZN(n14017) );
  NAND4_X1 U17540 ( .A1(n14020), .A2(n14019), .A3(n14018), .A4(n14017), .ZN(
        n14037) );
  INV_X1 U17541 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14167) );
  NOR4_X1 U17542 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n14167), .A3(
        n14213), .A4(n14056), .ZN(n14024) );
  INV_X1 U17543 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n20800) );
  INV_X1 U17544 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14091) );
  NOR4_X1 U17545 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_11__7__SCAN_IN), .A3(n20800), .A4(n14091), .ZN(n14023) );
  NOR2_X1 U17546 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20058) );
  INV_X1 U17547 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14166) );
  INV_X1 U17548 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15028) );
  NOR4_X1 U17549 ( .A1(n14021), .A2(n14166), .A3(n14354), .A4(n15028), .ZN(
        n14022) );
  NAND4_X1 U17550 ( .A1(n14024), .A2(n14023), .A3(n20058), .A4(n14022), .ZN(
        n14036) );
  INV_X1 U17551 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n17958) );
  NOR4_X1 U17552 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        BUF2_REG_25__SCAN_IN), .A3(n17958), .A4(n18727), .ZN(n14028) );
  INV_X1 U17553 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21665) );
  NOR4_X1 U17554 ( .A1(P1_ADDRESS_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_10__SCAN_IN), .A3(P3_DATAO_REG_23__SCAN_IN), .A4(
        n21665), .ZN(n14027) );
  INV_X1 U17555 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n21122) );
  NOR4_X1 U17556 ( .A1(BUF1_REG_13__SCAN_IN), .A2(P2_LWORD_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(n21122), .ZN(n14026) );
  INV_X1 U17557 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19960) );
  NOR4_X1 U17558 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_REIP_REG_22__SCAN_IN), .A3(P1_LWORD_REG_10__SCAN_IN), .A4(n19960), 
        .ZN(n14025) );
  NAND4_X1 U17559 ( .A1(n14028), .A2(n14027), .A3(n14026), .A4(n14025), .ZN(
        n14035) );
  NOR4_X1 U17560 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_EAX_REG_14__SCAN_IN), .A3(P1_EAX_REG_23__SCAN_IN), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n14033) );
  INV_X1 U17561 ( .A(DATAI_12_), .ZN(n14029) );
  NOR4_X1 U17562 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_11__4__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A4(n14029), .ZN(n14032) );
  NOR4_X1 U17563 ( .A1(P3_ADDRESS_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(n13675), .A4(n14102), .ZN(n14031)
         );
  INV_X1 U17564 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14095) );
  INV_X1 U17565 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n17986) );
  NOR4_X1 U17566 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(P2_REIP_REG_14__SCAN_IN), 
        .A3(n14095), .A4(n17986), .ZN(n14030) );
  NAND4_X1 U17567 ( .A1(n14033), .A2(n14032), .A3(n14031), .A4(n14030), .ZN(
        n14034) );
  NOR4_X1 U17568 ( .A1(n14037), .A2(n14036), .A3(n14035), .A4(n14034), .ZN(
        n14038) );
  NAND4_X1 U17569 ( .A1(n14041), .A2(n14040), .A3(n14039), .A4(n14038), .ZN(
        n14230) );
  INV_X1 U17570 ( .A(P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(n19926) );
  INV_X1 U17571 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n20006) );
  AOI22_X1 U17572 ( .A1(n19926), .A2(keyinput9), .B1(keyinput20), .B2(n20006), 
        .ZN(n14042) );
  OAI221_X1 U17573 ( .B1(n19926), .B2(keyinput9), .C1(n20006), .C2(keyinput20), 
        .A(n14042), .ZN(n14051) );
  INV_X1 U17574 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n14044) );
  AOI22_X1 U17575 ( .A1(n15588), .A2(keyinput6), .B1(keyinput105), .B2(n14044), 
        .ZN(n14043) );
  OAI221_X1 U17576 ( .B1(n15588), .B2(keyinput6), .C1(n14044), .C2(keyinput105), .A(n14043), .ZN(n14050) );
  XOR2_X1 U17577 ( .A(n12995), .B(keyinput79), .Z(n14047) );
  XNOR2_X1 U17578 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B(keyinput99), .ZN(
        n14046) );
  XNOR2_X1 U17579 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(keyinput63), 
        .ZN(n14045) );
  NAND3_X1 U17580 ( .A1(n14047), .A2(n14046), .A3(n14045), .ZN(n14049) );
  INV_X1 U17581 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19975) );
  XNOR2_X1 U17582 ( .A(n19975), .B(keyinput11), .ZN(n14048) );
  NOR4_X1 U17583 ( .A1(n14051), .A2(n14050), .A3(n14049), .A4(n14048), .ZN(
        n14089) );
  INV_X1 U17584 ( .A(P3_UWORD_REG_4__SCAN_IN), .ZN(n14054) );
  AOI22_X1 U17585 ( .A1(n14054), .A2(keyinput13), .B1(n14053), .B2(keyinput100), .ZN(n14052) );
  OAI221_X1 U17586 ( .B1(n14054), .B2(keyinput13), .C1(n14053), .C2(
        keyinput100), .A(n14052), .ZN(n14063) );
  AOI22_X1 U17587 ( .A1(n14057), .A2(keyinput47), .B1(n14056), .B2(keyinput49), 
        .ZN(n14055) );
  OAI221_X1 U17588 ( .B1(n14057), .B2(keyinput47), .C1(n14056), .C2(keyinput49), .A(n14055), .ZN(n14062) );
  INV_X1 U17589 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n21145) );
  AOI22_X1 U17590 ( .A1(n15803), .A2(keyinput26), .B1(n21145), .B2(keyinput122), .ZN(n14058) );
  OAI221_X1 U17591 ( .B1(n15803), .B2(keyinput26), .C1(n21145), .C2(
        keyinput122), .A(n14058), .ZN(n14061) );
  AOI22_X1 U17592 ( .A1(n11589), .A2(keyinput60), .B1(keyinput56), .B2(n11785), 
        .ZN(n14059) );
  OAI221_X1 U17593 ( .B1(n11589), .B2(keyinput60), .C1(n11785), .C2(keyinput56), .A(n14059), .ZN(n14060) );
  NOR4_X1 U17594 ( .A1(n14063), .A2(n14062), .A3(n14061), .A4(n14060), .ZN(
        n14088) );
  AOI22_X1 U17595 ( .A1(n20978), .A2(keyinput75), .B1(n14065), .B2(keyinput66), 
        .ZN(n14064) );
  OAI221_X1 U17596 ( .B1(n20978), .B2(keyinput75), .C1(n14065), .C2(keyinput66), .A(n14064), .ZN(n14073) );
  AOI22_X1 U17597 ( .A1(n14067), .A2(keyinput32), .B1(n21672), .B2(keyinput59), 
        .ZN(n14066) );
  OAI221_X1 U17598 ( .B1(n14067), .B2(keyinput32), .C1(n21672), .C2(keyinput59), .A(n14066), .ZN(n14072) );
  INV_X1 U17599 ( .A(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n19500) );
  AOI22_X1 U17600 ( .A1(n19500), .A2(keyinput44), .B1(n16246), .B2(keyinput111), .ZN(n14068) );
  OAI221_X1 U17601 ( .B1(n19500), .B2(keyinput44), .C1(n16246), .C2(
        keyinput111), .A(n14068), .ZN(n14071) );
  AOI22_X1 U17602 ( .A1(n17007), .A2(keyinput1), .B1(keyinput90), .B2(n16849), 
        .ZN(n14069) );
  OAI221_X1 U17603 ( .B1(n17007), .B2(keyinput1), .C1(n16849), .C2(keyinput90), 
        .A(n14069), .ZN(n14070) );
  NOR4_X1 U17604 ( .A1(n14073), .A2(n14072), .A3(n14071), .A4(n14070), .ZN(
        n14087) );
  INV_X1 U17605 ( .A(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17780) );
  AOI22_X1 U17606 ( .A1(n17780), .A2(keyinput38), .B1(n21694), .B2(keyinput113), .ZN(n14074) );
  OAI221_X1 U17607 ( .B1(n17780), .B2(keyinput38), .C1(n21694), .C2(
        keyinput113), .A(n14074), .ZN(n14085) );
  INV_X1 U17608 ( .A(P3_UWORD_REG_3__SCAN_IN), .ZN(n14077) );
  AOI22_X1 U17609 ( .A1(n14077), .A2(keyinput5), .B1(n14076), .B2(keyinput42), 
        .ZN(n14075) );
  OAI221_X1 U17610 ( .B1(n14077), .B2(keyinput5), .C1(n14076), .C2(keyinput42), 
        .A(n14075), .ZN(n14084) );
  INV_X1 U17611 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n19228) );
  AOI22_X1 U17612 ( .A1(n19228), .A2(keyinput35), .B1(n14079), .B2(keyinput101), .ZN(n14078) );
  OAI221_X1 U17613 ( .B1(n19228), .B2(keyinput35), .C1(n14079), .C2(
        keyinput101), .A(n14078), .ZN(n14083) );
  XNOR2_X1 U17614 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput88), 
        .ZN(n14081) );
  XNOR2_X1 U17615 ( .A(DATAI_12_), .B(keyinput68), .ZN(n14080) );
  NAND2_X1 U17616 ( .A1(n14081), .A2(n14080), .ZN(n14082) );
  NOR4_X1 U17617 ( .A1(n14085), .A2(n14084), .A3(n14083), .A4(n14082), .ZN(
        n14086) );
  NAND4_X1 U17618 ( .A1(n14089), .A2(n14088), .A3(n14087), .A4(n14086), .ZN(
        n14228) );
  AOI22_X1 U17619 ( .A1(n14091), .A2(keyinput53), .B1(keyinput72), .B2(n18678), 
        .ZN(n14090) );
  OAI221_X1 U17620 ( .B1(n14091), .B2(keyinput53), .C1(n18678), .C2(keyinput72), .A(n14090), .ZN(n14099) );
  INV_X1 U17621 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n21126) );
  AOI22_X1 U17622 ( .A1(n21126), .A2(keyinput50), .B1(n16212), .B2(keyinput52), 
        .ZN(n14092) );
  OAI221_X1 U17623 ( .B1(n21126), .B2(keyinput50), .C1(n16212), .C2(keyinput52), .A(n14092), .ZN(n14098) );
  INV_X1 U17624 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20871) );
  AOI22_X1 U17625 ( .A1(n17986), .A2(keyinput65), .B1(n20871), .B2(keyinput43), 
        .ZN(n14093) );
  OAI221_X1 U17626 ( .B1(n17986), .B2(keyinput65), .C1(n20871), .C2(keyinput43), .A(n14093), .ZN(n14097) );
  AOI22_X1 U17627 ( .A1(n14095), .A2(keyinput93), .B1(n20865), .B2(keyinput54), 
        .ZN(n14094) );
  OAI221_X1 U17628 ( .B1(n14095), .B2(keyinput93), .C1(n20865), .C2(keyinput54), .A(n14094), .ZN(n14096) );
  NOR4_X1 U17629 ( .A1(n14099), .A2(n14098), .A3(n14097), .A4(n14096), .ZN(
        n14129) );
  INV_X1 U17630 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19978) );
  AOI22_X1 U17631 ( .A1(n19978), .A2(keyinput78), .B1(n13675), .B2(keyinput39), 
        .ZN(n14100) );
  OAI221_X1 U17632 ( .B1(n19978), .B2(keyinput78), .C1(n13675), .C2(keyinput39), .A(n14100), .ZN(n14109) );
  INV_X1 U17633 ( .A(P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n21643) );
  AOI22_X1 U17634 ( .A1(n14102), .A2(keyinput81), .B1(keyinput51), .B2(n21643), 
        .ZN(n14101) );
  OAI221_X1 U17635 ( .B1(n14102), .B2(keyinput81), .C1(n21643), .C2(keyinput51), .A(n14101), .ZN(n14108) );
  AOI22_X1 U17636 ( .A1(n21665), .A2(keyinput112), .B1(n14104), .B2(keyinput86), .ZN(n14103) );
  OAI221_X1 U17637 ( .B1(n21665), .B2(keyinput112), .C1(n14104), .C2(
        keyinput86), .A(n14103), .ZN(n14107) );
  INV_X1 U17638 ( .A(P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19927) );
  INV_X1 U17639 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n21717) );
  AOI22_X1 U17640 ( .A1(n19927), .A2(keyinput69), .B1(n21717), .B2(keyinput21), 
        .ZN(n14105) );
  OAI221_X1 U17641 ( .B1(n19927), .B2(keyinput69), .C1(n21717), .C2(keyinput21), .A(n14105), .ZN(n14106) );
  NOR4_X1 U17642 ( .A1(n14109), .A2(n14108), .A3(n14107), .A4(n14106), .ZN(
        n14128) );
  INV_X1 U17643 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n18695) );
  AOI22_X1 U17644 ( .A1(n18695), .A2(keyinput104), .B1(n17958), .B2(keyinput77), .ZN(n14110) );
  OAI221_X1 U17645 ( .B1(n18695), .B2(keyinput104), .C1(n17958), .C2(
        keyinput77), .A(n14110), .ZN(n14117) );
  INV_X1 U17646 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18018) );
  AOI22_X1 U17647 ( .A1(n11624), .A2(keyinput19), .B1(keyinput48), .B2(n18018), 
        .ZN(n14111) );
  OAI221_X1 U17648 ( .B1(n11624), .B2(keyinput19), .C1(n18018), .C2(keyinput48), .A(n14111), .ZN(n14116) );
  AOI22_X1 U17649 ( .A1(n18727), .A2(keyinput74), .B1(keyinput127), .B2(n19960), .ZN(n14112) );
  OAI221_X1 U17650 ( .B1(n18727), .B2(keyinput74), .C1(n19960), .C2(
        keyinput127), .A(n14112), .ZN(n14115) );
  INV_X1 U17651 ( .A(P1_LWORD_REG_10__SCAN_IN), .ZN(n21134) );
  AOI22_X1 U17652 ( .A1(n21134), .A2(keyinput84), .B1(n18987), .B2(keyinput34), 
        .ZN(n14113) );
  OAI221_X1 U17653 ( .B1(n21134), .B2(keyinput84), .C1(n18987), .C2(keyinput34), .A(n14113), .ZN(n14114) );
  NOR4_X1 U17654 ( .A1(n14117), .A2(n14116), .A3(n14115), .A4(n14114), .ZN(
        n14127) );
  INV_X1 U17655 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19985) );
  INV_X1 U17656 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n17966) );
  AOI22_X1 U17657 ( .A1(n19985), .A2(keyinput119), .B1(n17966), .B2(keyinput92), .ZN(n14118) );
  OAI221_X1 U17658 ( .B1(n19985), .B2(keyinput119), .C1(n17966), .C2(
        keyinput92), .A(n14118), .ZN(n14125) );
  INV_X1 U17659 ( .A(P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20827) );
  AOI22_X1 U17660 ( .A1(n20800), .A2(keyinput28), .B1(keyinput94), .B2(n20827), 
        .ZN(n14119) );
  OAI221_X1 U17661 ( .B1(n20800), .B2(keyinput28), .C1(n20827), .C2(keyinput94), .A(n14119), .ZN(n14124) );
  INV_X1 U17662 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n20268) );
  INV_X1 U17663 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n21721) );
  AOI22_X1 U17664 ( .A1(n20268), .A2(keyinput3), .B1(keyinput106), .B2(n21721), 
        .ZN(n14120) );
  OAI221_X1 U17665 ( .B1(n20268), .B2(keyinput3), .C1(n21721), .C2(keyinput106), .A(n14120), .ZN(n14123) );
  AOI22_X1 U17666 ( .A1(n21122), .A2(keyinput82), .B1(n15028), .B2(keyinput125), .ZN(n14121) );
  OAI221_X1 U17667 ( .B1(n21122), .B2(keyinput82), .C1(n15028), .C2(
        keyinput125), .A(n14121), .ZN(n14122) );
  NOR4_X1 U17668 ( .A1(n14125), .A2(n14124), .A3(n14123), .A4(n14122), .ZN(
        n14126) );
  NAND4_X1 U17669 ( .A1(n14129), .A2(n14128), .A3(n14127), .A4(n14126), .ZN(
        n14227) );
  INV_X1 U17670 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n18705) );
  AOI22_X1 U17671 ( .A1(n18705), .A2(keyinput80), .B1(n17959), .B2(keyinput33), 
        .ZN(n14130) );
  OAI221_X1 U17672 ( .B1(n18705), .B2(keyinput80), .C1(n17959), .C2(keyinput33), .A(n14130), .ZN(n14140) );
  AOI22_X1 U17673 ( .A1(n20243), .A2(keyinput124), .B1(n20071), .B2(
        keyinput118), .ZN(n14131) );
  OAI221_X1 U17674 ( .B1(n20243), .B2(keyinput124), .C1(n20071), .C2(
        keyinput118), .A(n14131), .ZN(n14139) );
  INV_X1 U17675 ( .A(DATAI_23_), .ZN(n14133) );
  AOI22_X1 U17676 ( .A1(n14133), .A2(keyinput58), .B1(keyinput87), .B2(n19967), 
        .ZN(n14132) );
  OAI221_X1 U17677 ( .B1(n14133), .B2(keyinput58), .C1(n19967), .C2(keyinput87), .A(n14132), .ZN(n14138) );
  INV_X1 U17678 ( .A(DATAI_27_), .ZN(n14135) );
  AOI22_X1 U17679 ( .A1(n14136), .A2(keyinput91), .B1(n14135), .B2(keyinput121), .ZN(n14134) );
  OAI221_X1 U17680 ( .B1(n14136), .B2(keyinput91), .C1(n14135), .C2(
        keyinput121), .A(n14134), .ZN(n14137) );
  NOR4_X1 U17681 ( .A1(n14140), .A2(n14139), .A3(n14138), .A4(n14137), .ZN(
        n14176) );
  INV_X1 U17682 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n20238) );
  AOI22_X1 U17683 ( .A1(n20238), .A2(keyinput85), .B1(n19646), .B2(keyinput62), 
        .ZN(n14141) );
  OAI221_X1 U17684 ( .B1(n20238), .B2(keyinput85), .C1(n19646), .C2(keyinput62), .A(n14141), .ZN(n14150) );
  INV_X1 U17685 ( .A(DATAI_17_), .ZN(n14143) );
  AOI22_X1 U17686 ( .A1(n14143), .A2(keyinput15), .B1(keyinput22), .B2(n13997), 
        .ZN(n14142) );
  OAI221_X1 U17687 ( .B1(n14143), .B2(keyinput15), .C1(n13997), .C2(keyinput22), .A(n14142), .ZN(n14149) );
  XNOR2_X1 U17688 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B(keyinput114), .ZN(
        n14147) );
  XNOR2_X1 U17689 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(keyinput117), 
        .ZN(n14146) );
  XNOR2_X1 U17690 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(keyinput67), 
        .ZN(n14145) );
  XNOR2_X1 U17691 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B(keyinput110), .ZN(
        n14144) );
  NAND4_X1 U17692 ( .A1(n14147), .A2(n14146), .A3(n14145), .A4(n14144), .ZN(
        n14148) );
  NOR3_X1 U17693 ( .A1(n14150), .A2(n14149), .A3(n14148), .ZN(n14175) );
  AOI22_X1 U17694 ( .A1(n14152), .A2(keyinput0), .B1(keyinput116), .B2(n17978), 
        .ZN(n14151) );
  OAI221_X1 U17695 ( .B1(n14152), .B2(keyinput0), .C1(n17978), .C2(keyinput116), .A(n14151), .ZN(n14161) );
  INV_X1 U17696 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19973) );
  AOI22_X1 U17697 ( .A1(n19973), .A2(keyinput2), .B1(n16331), .B2(keyinput97), 
        .ZN(n14153) );
  OAI221_X1 U17698 ( .B1(n19973), .B2(keyinput2), .C1(n16331), .C2(keyinput97), 
        .A(n14153), .ZN(n14160) );
  INV_X1 U17699 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14154) );
  XOR2_X1 U17700 ( .A(n14154), .B(keyinput4), .Z(n14158) );
  XNOR2_X1 U17701 ( .A(keyinput57), .B(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14157) );
  XNOR2_X1 U17702 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B(keyinput17), .ZN(
        n14156) );
  XNOR2_X1 U17703 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(keyinput8), 
        .ZN(n14155) );
  NAND4_X1 U17704 ( .A1(n14158), .A2(n14157), .A3(n14156), .A4(n14155), .ZN(
        n14159) );
  NOR3_X1 U17705 ( .A1(n14161), .A2(n14160), .A3(n14159), .ZN(n14174) );
  AOI22_X1 U17706 ( .A1(n13861), .A2(keyinput109), .B1(n16158), .B2(
        keyinput108), .ZN(n14162) );
  OAI221_X1 U17707 ( .B1(n13861), .B2(keyinput109), .C1(n16158), .C2(
        keyinput108), .A(n14162), .ZN(n14172) );
  INV_X1 U17708 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n18734) );
  AOI22_X1 U17709 ( .A1(n14164), .A2(keyinput71), .B1(keyinput37), .B2(n18734), 
        .ZN(n14163) );
  OAI221_X1 U17710 ( .B1(n14164), .B2(keyinput71), .C1(n18734), .C2(keyinput37), .A(n14163), .ZN(n14171) );
  AOI22_X1 U17711 ( .A1(n14167), .A2(keyinput89), .B1(n14166), .B2(keyinput102), .ZN(n14165) );
  OAI221_X1 U17712 ( .B1(n14167), .B2(keyinput89), .C1(n14166), .C2(
        keyinput102), .A(n14165), .ZN(n14170) );
  INV_X1 U17713 ( .A(P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n21642) );
  AOI22_X1 U17714 ( .A1(n21642), .A2(keyinput95), .B1(n18768), .B2(keyinput27), 
        .ZN(n14168) );
  OAI221_X1 U17715 ( .B1(n21642), .B2(keyinput95), .C1(n18768), .C2(keyinput27), .A(n14168), .ZN(n14169) );
  NOR4_X1 U17716 ( .A1(n14172), .A2(n14171), .A3(n14170), .A4(n14169), .ZN(
        n14173) );
  NAND4_X1 U17717 ( .A1(n14176), .A2(n14175), .A3(n14174), .A4(n14173), .ZN(
        n14226) );
  AOI22_X1 U17718 ( .A1(n14179), .A2(keyinput30), .B1(n14178), .B2(keyinput61), 
        .ZN(n14177) );
  OAI221_X1 U17719 ( .B1(n14179), .B2(keyinput30), .C1(n14178), .C2(keyinput61), .A(n14177), .ZN(n14187) );
  INV_X1 U17720 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n20003) );
  AOI22_X1 U17721 ( .A1(n21661), .A2(keyinput29), .B1(keyinput25), .B2(n20003), 
        .ZN(n14180) );
  OAI221_X1 U17722 ( .B1(n21661), .B2(keyinput29), .C1(n20003), .C2(keyinput25), .A(n14180), .ZN(n14186) );
  INV_X1 U17723 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20004) );
  AOI22_X1 U17724 ( .A1(n20004), .A2(keyinput10), .B1(n14182), .B2(keyinput36), 
        .ZN(n14181) );
  OAI221_X1 U17725 ( .B1(n20004), .B2(keyinput10), .C1(n14182), .C2(keyinput36), .A(n14181), .ZN(n14185) );
  INV_X1 U17726 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n21119) );
  AOI22_X1 U17727 ( .A1(n20856), .A2(keyinput115), .B1(keyinput14), .B2(n21119), .ZN(n14183) );
  OAI221_X1 U17728 ( .B1(n20856), .B2(keyinput115), .C1(n21119), .C2(
        keyinput14), .A(n14183), .ZN(n14184) );
  NOR4_X1 U17729 ( .A1(n14187), .A2(n14186), .A3(n14185), .A4(n14184), .ZN(
        n14224) );
  INV_X1 U17730 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19416) );
  INV_X1 U17731 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14189) );
  AOI22_X1 U17732 ( .A1(n19416), .A2(keyinput98), .B1(n14189), .B2(keyinput55), 
        .ZN(n14188) );
  OAI221_X1 U17733 ( .B1(n19416), .B2(keyinput98), .C1(n14189), .C2(keyinput55), .A(n14188), .ZN(n14199) );
  INV_X1 U17734 ( .A(P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n20826) );
  INV_X1 U17735 ( .A(DATAI_20_), .ZN(n14191) );
  AOI22_X1 U17736 ( .A1(n20826), .A2(keyinput70), .B1(n14191), .B2(keyinput76), 
        .ZN(n14190) );
  OAI221_X1 U17737 ( .B1(n20826), .B2(keyinput70), .C1(n14191), .C2(keyinput76), .A(n14190), .ZN(n14198) );
  AOI22_X1 U17738 ( .A1(keyinput23), .A2(n14193), .B1(keyinput83), .B2(n14231), 
        .ZN(n14192) );
  OAI21_X1 U17739 ( .B1(n14193), .B2(keyinput23), .A(n14192), .ZN(n14197) );
  XOR2_X1 U17740 ( .A(n21138), .B(keyinput31), .Z(n14195) );
  XNOR2_X1 U17741 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B(keyinput64), .ZN(
        n14194) );
  NAND2_X1 U17742 ( .A1(n14195), .A2(n14194), .ZN(n14196) );
  NOR4_X1 U17743 ( .A1(n14199), .A2(n14198), .A3(n14197), .A4(n14196), .ZN(
        n14223) );
  AOI22_X1 U17744 ( .A1(n20858), .A2(keyinput96), .B1(keyinput41), .B2(n14201), 
        .ZN(n14200) );
  OAI221_X1 U17745 ( .B1(n20858), .B2(keyinput96), .C1(n14201), .C2(keyinput41), .A(n14200), .ZN(n14209) );
  INV_X1 U17746 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n17956) );
  AOI22_X1 U17747 ( .A1(n19095), .A2(keyinput73), .B1(keyinput126), .B2(n17956), .ZN(n14202) );
  OAI221_X1 U17748 ( .B1(n19095), .B2(keyinput73), .C1(n17956), .C2(
        keyinput126), .A(n14202), .ZN(n14208) );
  INV_X1 U17749 ( .A(P3_LWORD_REG_0__SCAN_IN), .ZN(n18740) );
  AOI22_X1 U17750 ( .A1(n10343), .A2(keyinput12), .B1(keyinput16), .B2(n18740), 
        .ZN(n14203) );
  OAI221_X1 U17751 ( .B1(n10343), .B2(keyinput12), .C1(n18740), .C2(keyinput16), .A(n14203), .ZN(n14207) );
  XNOR2_X1 U17752 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B(keyinput24), .ZN(
        n14205) );
  XNOR2_X1 U17753 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B(keyinput45), .ZN(
        n14204) );
  NAND2_X1 U17754 ( .A1(n14205), .A2(n14204), .ZN(n14206) );
  NOR4_X1 U17755 ( .A1(n14209), .A2(n14208), .A3(n14207), .A4(n14206), .ZN(
        n14222) );
  INV_X1 U17756 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20021) );
  INV_X1 U17757 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n21140) );
  AOI22_X1 U17758 ( .A1(n20021), .A2(keyinput40), .B1(keyinput107), .B2(n21140), .ZN(n14210) );
  OAI221_X1 U17759 ( .B1(n20021), .B2(keyinput40), .C1(n21140), .C2(
        keyinput107), .A(n14210), .ZN(n14220) );
  AOI22_X1 U17760 ( .A1(n14213), .A2(keyinput46), .B1(n14212), .B2(keyinput7), 
        .ZN(n14211) );
  OAI221_X1 U17761 ( .B1(n14213), .B2(keyinput46), .C1(n14212), .C2(keyinput7), 
        .A(n14211), .ZN(n14219) );
  AOI22_X1 U17762 ( .A1(n20869), .A2(keyinput123), .B1(keyinput18), .B2(n21666), .ZN(n14214) );
  OAI221_X1 U17763 ( .B1(n20869), .B2(keyinput123), .C1(n21666), .C2(
        keyinput18), .A(n14214), .ZN(n14218) );
  INV_X1 U17764 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14216) );
  AOI22_X1 U17765 ( .A1(n9877), .A2(keyinput120), .B1(n14216), .B2(keyinput103), .ZN(n14215) );
  OAI221_X1 U17766 ( .B1(n9877), .B2(keyinput120), .C1(n14216), .C2(
        keyinput103), .A(n14215), .ZN(n14217) );
  NOR4_X1 U17767 ( .A1(n14220), .A2(n14219), .A3(n14218), .A4(n14217), .ZN(
        n14221) );
  NAND4_X1 U17768 ( .A1(n14224), .A2(n14223), .A3(n14222), .A4(n14221), .ZN(
        n14225) );
  NOR4_X1 U17769 ( .A1(n14228), .A2(n14227), .A3(n14226), .A4(n14225), .ZN(
        n14229) );
  OAI221_X1 U17770 ( .B1(keyinput83), .B2(n14231), .C1(keyinput83), .C2(n14230), .A(n14229), .ZN(n14232) );
  XNOR2_X1 U17771 ( .A(n14233), .B(n14232), .ZN(P2_U3045) );
  NAND2_X1 U17772 ( .A1(n20051), .A2(n10081), .ZN(n18445) );
  INV_X1 U17773 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18324) );
  NAND3_X1 U17774 ( .A1(n20035), .A2(n20047), .A3(n18037), .ZN(n19925) );
  NOR2_X1 U17775 ( .A1(n18678), .A2(n19925), .ZN(n18414) );
  NAND2_X1 U17776 ( .A1(n18406), .A2(n18414), .ZN(n18247) );
  NOR2_X1 U17777 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n20016), .ZN(n19918) );
  INV_X1 U17778 ( .A(n19918), .ZN(n19907) );
  OAI211_X1 U17779 ( .C1(n19920), .C2(n19907), .A(n19923), .B(n19110), .ZN(
        n14236) );
  OAI21_X1 U17780 ( .B1(n18324), .B2(n18247), .A(n18435), .ZN(n14243) );
  AOI21_X1 U17781 ( .B1(n18406), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n19923), .ZN(n18276) );
  INV_X1 U17782 ( .A(n18276), .ZN(n18367) );
  OR2_X1 U17783 ( .A1(n20031), .A2(n20030), .ZN(n14238) );
  NOR2_X1 U17784 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(n20032), .ZN(n14237) );
  NAND2_X1 U17785 ( .A1(n14238), .A2(n14237), .ZN(n19903) );
  NAND2_X1 U17786 ( .A1(n20031), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n14240) );
  NAND2_X1 U17787 ( .A1(n19903), .A2(n14240), .ZN(n14239) );
  OAI22_X1 U17788 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18367), .B1(
        n9878), .B2(n18437), .ZN(n14242) );
  AOI211_X4 U17789 ( .C1(n18037), .C2(n20040), .A(n20049), .B(n14240), .ZN(
        n18416) );
  OR2_X1 U17790 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(
        n18420) );
  NAND2_X1 U17791 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n18581) );
  NAND2_X1 U17792 ( .A1(n18420), .A2(n18581), .ZN(n18588) );
  OAI22_X1 U17793 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18408), .B1(n18436), 
        .B2(n18588), .ZN(n14241) );
  AOI211_X1 U17794 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n14243), .A(
        n14242), .B(n14241), .ZN(n14245) );
  NAND2_X1 U17795 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18385), .ZN(n14244) );
  OAI211_X1 U17796 ( .C1(n18445), .C2(n14246), .A(n14245), .B(n14244), .ZN(
        P3_U2670) );
  MUX2_X1 U17797 ( .A(n14247), .B(n14360), .S(n16760), .Z(n14248) );
  OAI21_X1 U17798 ( .B1(n20912), .B2(n16752), .A(n14248), .ZN(P2_U2886) );
  AND2_X1 U17799 ( .A1(n14249), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n16890) );
  NAND2_X1 U17800 ( .A1(n14250), .A2(n16890), .ZN(n16894) );
  NOR2_X1 U17801 ( .A1(n16894), .A2(n14251), .ZN(n14490) );
  XNOR2_X1 U17802 ( .A(n14490), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14256) );
  OAI21_X1 U17803 ( .B1(n14252), .B2(n14254), .A(n14253), .ZN(n20173) );
  MUX2_X1 U17804 ( .A(n10969), .B(n20173), .S(n16760), .Z(n14255) );
  OAI21_X1 U17805 ( .B1(n14256), .B2(n16752), .A(n14255), .ZN(P2_U2880) );
  INV_X1 U17806 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n16588) );
  INV_X1 U17807 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14257) );
  NOR2_X1 U17808 ( .A1(n16894), .A2(n14257), .ZN(n14259) );
  INV_X1 U17809 ( .A(n14490), .ZN(n14258) );
  OAI211_X1 U17810 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n14259), .A(
        n14258), .B(n16757), .ZN(n14263) );
  NOR2_X1 U17811 ( .A1(n14611), .A2(n14260), .ZN(n14261) );
  OR2_X1 U17812 ( .A1(n14252), .A2(n14261), .ZN(n17409) );
  INV_X1 U17813 ( .A(n17409), .ZN(n16594) );
  NAND2_X1 U17814 ( .A1(n16594), .A2(n16760), .ZN(n14262) );
  OAI211_X1 U17815 ( .C1(n20207), .C2(n16588), .A(n14263), .B(n14262), .ZN(
        P2_U2881) );
  NOR2_X1 U17816 ( .A1(n14265), .A2(n14264), .ZN(n17191) );
  NOR3_X1 U17817 ( .A1(n17458), .A2(n14266), .A3(n17191), .ZN(n14267) );
  AOI21_X1 U17818 ( .B1(n17461), .B2(n20923), .A(n14267), .ZN(n14268) );
  INV_X1 U17819 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20849) );
  OR2_X1 U17820 ( .A1(n17149), .A2(n20849), .ZN(n17185) );
  OAI211_X1 U17821 ( .C1(n17429), .C2(n14582), .A(n14268), .B(n17185), .ZN(
        n14269) );
  AOI211_X1 U17822 ( .C1(n14271), .C2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n14270), .B(n14269), .ZN(n14279) );
  INV_X1 U17823 ( .A(n14272), .ZN(n14273) );
  NAND2_X1 U17824 ( .A1(n14274), .A2(n14273), .ZN(n17195) );
  NAND3_X1 U17825 ( .A1(n17454), .A2(n17197), .A3(n17195), .ZN(n14275) );
  OAI21_X1 U17826 ( .B1(n14828), .B2(n14276), .A(n14275), .ZN(n14277) );
  INV_X1 U17827 ( .A(n14277), .ZN(n14278) );
  OAI211_X1 U17828 ( .C1(n14281), .C2(n14280), .A(n14279), .B(n14278), .ZN(
        P2_U3044) );
  NOR2_X1 U17829 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13237), .ZN(n14309) );
  MUX2_X1 U17830 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14282), .S(
        n17825), .Z(n17832) );
  AOI22_X1 U17831 ( .A1(n14309), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n17832), .B2(n13237), .ZN(n14303) );
  NAND2_X1 U17832 ( .A1(n21739), .A2(n14283), .ZN(n14298) );
  NAND2_X1 U17833 ( .A1(n12518), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14285) );
  NAND2_X1 U17834 ( .A1(n14285), .A2(n21737), .ZN(n14286) );
  NAND2_X1 U17835 ( .A1(n12762), .A2(n14286), .ZN(n21731) );
  AOI21_X1 U17836 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n14290), .A(
        n14287), .ZN(n14294) );
  MUX2_X1 U17837 ( .A(n14287), .B(n14299), .S(n12518), .Z(n14289) );
  OAI21_X1 U17838 ( .B1(n14290), .B2(n14289), .A(n14288), .ZN(n14292) );
  NAND2_X1 U17839 ( .A1(n16349), .A2(n21737), .ZN(n14291) );
  OAI211_X1 U17840 ( .C1(n14294), .C2(n14293), .A(n14292), .B(n14291), .ZN(
        n14295) );
  AOI21_X1 U17841 ( .B1(n14296), .B2(n21731), .A(n14295), .ZN(n14297) );
  NAND2_X1 U17842 ( .A1(n14298), .A2(n14297), .ZN(n21734) );
  NOR2_X1 U17843 ( .A1(n17825), .A2(n14299), .ZN(n14300) );
  AOI21_X1 U17844 ( .B1(n21734), .B2(n17825), .A(n14300), .ZN(n17833) );
  INV_X1 U17845 ( .A(n17833), .ZN(n14301) );
  AOI22_X1 U17846 ( .A1(n14301), .A2(n13237), .B1(n21737), .B2(n14309), .ZN(
        n14302) );
  AOI21_X1 U17847 ( .B1(n21053), .B2(n14306), .A(n14305), .ZN(n14308) );
  OAI21_X1 U17848 ( .B1(n17825), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13237), .ZN(n14307) );
  OR2_X1 U17849 ( .A1(n14308), .A2(n14307), .ZN(n14311) );
  NAND2_X1 U17850 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n14309), .ZN(
        n14310) );
  NAND2_X1 U17851 ( .A1(n14311), .A2(n14310), .ZN(n17842) );
  INV_X1 U17852 ( .A(n17842), .ZN(n14312) );
  OAI21_X1 U17853 ( .B1(n17843), .B2(n14304), .A(n14312), .ZN(n14316) );
  NOR2_X1 U17854 ( .A1(n14316), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n14315) );
  NOR2_X1 U17855 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21765) );
  OR2_X1 U17856 ( .A1(n14316), .A2(n17928), .ZN(n17858) );
  INV_X1 U17857 ( .A(n17858), .ZN(n14318) );
  NOR2_X1 U17858 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n13237), .ZN(n21740) );
  OAI22_X1 U17859 ( .A1(n14665), .A2(n21584), .B1(n21740), .B2(n15789), .ZN(
        n14317) );
  OAI21_X1 U17860 ( .B1(n14318), .B2(n14317), .A(n21747), .ZN(n14319) );
  OAI21_X1 U17861 ( .B1(n21747), .B2(n21422), .A(n14319), .ZN(P1_U3478) );
  AND2_X2 U17862 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14322) );
  NOR2_X1 U17863 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n14322), .ZN(
        n14323) );
  NOR2_X1 U17864 ( .A1(n14548), .A2(n14323), .ZN(n21066) );
  INV_X1 U17865 ( .A(n15378), .ZN(n15149) );
  INV_X1 U17866 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n21069) );
  OAI22_X1 U17867 ( .A1(n21066), .A2(n15565), .B1(n15149), .B2(n21069), .ZN(
        n14324) );
  AOI21_X1 U17868 ( .B1(n15379), .B2(P1_EAX_REG_3__SCAN_IN), .A(n14324), .ZN(
        n14327) );
  NAND2_X1 U17869 ( .A1(n14325), .A2(n21737), .ZN(n14326) );
  OAI21_X2 U17870 ( .B1(n21743), .B2(n15082), .A(n14328), .ZN(n14329) );
  NAND2_X1 U17871 ( .A1(n14330), .A2(n14329), .ZN(n14546) );
  OAI21_X1 U17872 ( .B1(n14330), .B2(n14329), .A(n14546), .ZN(n21073) );
  INV_X1 U17873 ( .A(n15861), .ZN(n14468) );
  INV_X1 U17874 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n21147) );
  OAI222_X1 U17875 ( .A1(n21073), .A2(n15897), .B1(n15901), .B2(n14468), .C1(
        n15899), .C2(n21147), .ZN(P1_U2901) );
  AND2_X1 U17876 ( .A1(n14387), .A2(n14386), .ZN(n14367) );
  INV_X1 U17877 ( .A(n14331), .ZN(n14332) );
  NAND2_X1 U17878 ( .A1(n14332), .A2(n14811), .ZN(n14368) );
  XNOR2_X1 U17879 ( .A(n14368), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14341) );
  INV_X1 U17880 ( .A(n14333), .ZN(n14334) );
  OR2_X1 U17881 ( .A1(n14335), .A2(n14334), .ZN(n14375) );
  OAI21_X1 U17882 ( .B1(n12330), .B2(n14353), .A(n10554), .ZN(n14336) );
  NAND2_X1 U17883 ( .A1(n14375), .A2(n14336), .ZN(n14340) );
  OAI211_X1 U17884 ( .C1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n14337), .A(
        n11412), .B(n14338), .ZN(n14339) );
  OAI211_X1 U17885 ( .C1(n14367), .C2(n14341), .A(n14340), .B(n14339), .ZN(
        n14342) );
  AOI21_X1 U17886 ( .B1(n17446), .B2(n14363), .A(n14342), .ZN(n17474) );
  NOR2_X1 U17887 ( .A1(n14344), .A2(n14343), .ZN(n14345) );
  NAND2_X1 U17888 ( .A1(n14346), .A2(n14345), .ZN(n14351) );
  NAND2_X1 U17889 ( .A1(n14404), .A2(n14347), .ZN(n14348) );
  AOI211_X1 U17890 ( .C1(n14349), .C2(n14348), .A(n20963), .B(n20834), .ZN(
        n14350) );
  INV_X1 U17891 ( .A(n14803), .ZN(n14352) );
  MUX2_X1 U17892 ( .A(n14353), .B(n17474), .S(n14352), .Z(n14400) );
  INV_X1 U17893 ( .A(n14363), .ZN(n14378) );
  AOI21_X1 U17894 ( .B1(n14354), .B2(n14358), .A(n14331), .ZN(n14357) );
  NAND2_X1 U17895 ( .A1(n14356), .A2(n14355), .ZN(n14361) );
  AOI22_X1 U17896 ( .A1(n11412), .A2(n14358), .B1(n14357), .B2(n14361), .ZN(
        n14359) );
  OAI21_X1 U17897 ( .B1(n14360), .B2(n14378), .A(n14359), .ZN(n17469) );
  MUX2_X1 U17898 ( .A(n14361), .B(n11412), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n14362) );
  AOI21_X1 U17899 ( .B1(n17455), .B2(n14363), .A(n14362), .ZN(n17465) );
  NAND2_X1 U17900 ( .A1(n17465), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n14364) );
  OAI21_X1 U17901 ( .B1(n17469), .B2(n14364), .A(n20938), .ZN(n14366) );
  NAND2_X1 U17902 ( .A1(n17469), .A2(n14364), .ZN(n14365) );
  AOI21_X1 U17903 ( .B1(n14366), .B2(n14365), .A(n14803), .ZN(n14382) );
  INV_X1 U17904 ( .A(n14367), .ZN(n14372) );
  NAND2_X1 U17905 ( .A1(n14369), .A2(n14368), .ZN(n14373) );
  NOR2_X1 U17906 ( .A1(n14370), .A2(n14337), .ZN(n14371) );
  AOI22_X1 U17907 ( .A1(n14372), .A2(n14373), .B1(n14371), .B2(n11412), .ZN(
        n14377) );
  INV_X1 U17908 ( .A(n14373), .ZN(n14374) );
  NAND2_X1 U17909 ( .A1(n14375), .A2(n14374), .ZN(n14376) );
  OAI211_X1 U17910 ( .C1(n14582), .C2(n14378), .A(n14377), .B(n14376), .ZN(
        n14806) );
  OR2_X1 U17911 ( .A1(n14806), .A2(n14803), .ZN(n14380) );
  NAND2_X1 U17912 ( .A1(n14803), .A2(n14811), .ZN(n14379) );
  NAND2_X1 U17913 ( .A1(n14380), .A2(n14379), .ZN(n14399) );
  INV_X1 U17914 ( .A(n14399), .ZN(n14381) );
  OAI21_X1 U17915 ( .B1(n14382), .B2(n20927), .A(n14381), .ZN(n14383) );
  NAND2_X1 U17916 ( .A1(n14382), .A2(n20927), .ZN(n14384) );
  AND3_X1 U17917 ( .A1(n14400), .A2(n14383), .A3(n14384), .ZN(n14385) );
  OAI22_X1 U17918 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n14385), .B1(
        n14400), .B2(n14384), .ZN(n14402) );
  INV_X1 U17919 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17862) );
  MUX2_X1 U17920 ( .A(n14387), .B(n14386), .S(n14410), .Z(n14391) );
  NAND2_X1 U17921 ( .A1(n14389), .A2(n14388), .ZN(n14390) );
  NAND2_X1 U17922 ( .A1(n14391), .A2(n14390), .ZN(n20955) );
  NOR2_X1 U17923 ( .A1(P2_MORE_REG_SCAN_IN), .A2(P2_FLUSH_REG_SCAN_IN), .ZN(
        n14395) );
  INV_X1 U17924 ( .A(n14392), .ZN(n14393) );
  NOR2_X1 U17925 ( .A1(n16694), .A2(n14393), .ZN(n14394) );
  NAND2_X1 U17926 ( .A1(n11185), .A2(n14394), .ZN(n17477) );
  OAI211_X1 U17927 ( .C1(n14396), .C2(n14395), .A(n20950), .B(n17477), .ZN(
        n14397) );
  AOI211_X1 U17928 ( .C1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n14803), .A(
        n20955), .B(n14397), .ZN(n14398) );
  OAI21_X1 U17929 ( .B1(n14400), .B2(n14399), .A(n14398), .ZN(n14401) );
  AOI21_X1 U17930 ( .B1(n14402), .B2(n17862), .A(n14401), .ZN(n14416) );
  AOI21_X1 U17931 ( .B1(n14416), .B2(n11055), .A(n11573), .ZN(n14407) );
  NAND2_X1 U17932 ( .A1(n14404), .A2(n14403), .ZN(n14406) );
  NOR2_X1 U17933 ( .A1(n20959), .A2(n20939), .ZN(n14405) );
  NAND2_X1 U17934 ( .A1(n14406), .A2(n14405), .ZN(n14413) );
  AOI211_X1 U17935 ( .C1(n20951), .C2(n14800), .A(n14409), .B(n14408), .ZN(
        n14415) );
  INV_X1 U17936 ( .A(n17484), .ZN(n17470) );
  NAND2_X1 U17937 ( .A1(n14411), .A2(n11573), .ZN(n20969) );
  OAI21_X1 U17938 ( .B1(n17470), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n20969), 
        .ZN(n14412) );
  OAI21_X1 U17939 ( .B1(n14413), .B2(n20966), .A(n14412), .ZN(n14414) );
  OAI211_X1 U17940 ( .C1(n14416), .C2(n14802), .A(n14415), .B(n14414), .ZN(
        n14417) );
  AOI21_X1 U17941 ( .B1(n14504), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n14417), 
        .ZN(n14418) );
  INV_X1 U17942 ( .A(n14418), .ZN(P2_U3176) );
  INV_X1 U17943 ( .A(n14419), .ZN(n14423) );
  NOR2_X1 U17944 ( .A1(n14419), .A2(n14420), .ZN(n14565) );
  INV_X1 U17945 ( .A(n14565), .ZN(n14421) );
  OAI211_X1 U17946 ( .C1(n14423), .C2(n14422), .A(n14421), .B(n16757), .ZN(
        n14428) );
  OAI21_X1 U17947 ( .B1(n14424), .B2(n14426), .A(n14562), .ZN(n20140) );
  INV_X1 U17948 ( .A(n20140), .ZN(n17366) );
  NAND2_X1 U17949 ( .A1(n17366), .A2(n16760), .ZN(n14427) );
  OAI211_X1 U17950 ( .C1(n16760), .C2(n14429), .A(n14428), .B(n14427), .ZN(
        P2_U2877) );
  OAI21_X1 U17951 ( .B1(n14504), .B2(n11573), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n14430) );
  NAND2_X1 U17952 ( .A1(n14430), .A2(n17860), .ZN(P2_U3593) );
  OAI21_X1 U17953 ( .B1(n14433), .B2(n14432), .A(n14431), .ZN(n16540) );
  INV_X1 U17954 ( .A(n14434), .ZN(n14435) );
  INV_X1 U17955 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n20244) );
  OAI222_X1 U17956 ( .A1(n16540), .A2(n14700), .B1(n14435), .B2(n20232), .C1(
        n20244), .C2(n16897), .ZN(P2_U2906) );
  AOI22_X1 U17957 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n14478), .B1(DATAI_24_), 
        .B2(n14437), .ZN(n21538) );
  NOR2_X1 U17958 ( .A1(n21575), .A2(n21361), .ZN(n14714) );
  INV_X1 U17959 ( .A(n21365), .ZN(n14440) );
  NAND2_X1 U17960 ( .A1(n21186), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21580) );
  INV_X1 U17961 ( .A(n21580), .ZN(n14439) );
  NAND2_X1 U17962 ( .A1(n14440), .A2(n14439), .ZN(n14661) );
  OR2_X1 U17963 ( .A1(n21391), .A2(n14441), .ZN(n21338) );
  INV_X1 U17964 ( .A(n21338), .ZN(n21362) );
  AND2_X1 U17965 ( .A1(n14442), .A2(n13502), .ZN(n21572) );
  INV_X1 U17966 ( .A(n14480), .ZN(n14443) );
  AOI21_X1 U17967 ( .B1(n21362), .B2(n21572), .A(n14443), .ZN(n14446) );
  NAND3_X1 U17968 ( .A1(n14661), .A2(n21586), .A3(n14446), .ZN(n14444) );
  NAND2_X1 U17969 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n14452) );
  AOI22_X1 U17970 ( .A1(DATAI_16_), .A2(n14437), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n14478), .ZN(n21590) );
  INV_X1 U17971 ( .A(n21590), .ZN(n21523) );
  INV_X1 U17972 ( .A(n21577), .ZN(n21466) );
  INV_X1 U17973 ( .A(n14446), .ZN(n14447) );
  AOI22_X1 U17974 ( .A1(n14447), .A2(n21586), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14714), .ZN(n14481) );
  NAND2_X1 U17975 ( .A1(n14479), .A2(n14449), .ZN(n21291) );
  OAI22_X1 U17976 ( .A1(n21466), .A2(n14481), .B1(n14480), .B2(n21291), .ZN(
        n14450) );
  AOI21_X1 U17977 ( .B1(n21418), .B2(n21523), .A(n14450), .ZN(n14451) );
  OAI211_X1 U17978 ( .C1(n21538), .C2(n14742), .A(n14452), .B(n14451), .ZN(
        P1_U3089) );
  AOI22_X1 U17979 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n14478), .B1(DATAI_30_), 
        .B2(n14437), .ZN(n21562) );
  NAND2_X1 U17980 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n14455) );
  AOI22_X1 U17981 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n14478), .B1(DATAI_22_), 
        .B2(n14437), .ZN(n21626) );
  INV_X1 U17982 ( .A(n21626), .ZN(n21559) );
  INV_X1 U17983 ( .A(n15850), .ZN(n14770) );
  INV_X1 U17984 ( .A(n21621), .ZN(n21484) );
  NAND2_X1 U17985 ( .A1(n14479), .A2(n12632), .ZN(n21324) );
  OAI22_X1 U17986 ( .A1(n21484), .A2(n14481), .B1(n14480), .B2(n21324), .ZN(
        n14453) );
  AOI21_X1 U17987 ( .B1(n21418), .B2(n21559), .A(n14453), .ZN(n14454) );
  OAI211_X1 U17988 ( .C1(n21562), .C2(n14742), .A(n14455), .B(n14454), .ZN(
        P1_U3095) );
  AOI22_X1 U17989 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n14478), .B1(DATAI_29_), 
        .B2(n14437), .ZN(n21558) );
  NAND2_X1 U17990 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14458) );
  AOI22_X1 U17991 ( .A1(DATAI_21_), .A2(n14437), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n14478), .ZN(n21620) );
  INV_X1 U17992 ( .A(n21620), .ZN(n21555) );
  INV_X1 U17993 ( .A(n15853), .ZN(n14657) );
  INV_X1 U17994 ( .A(n21615), .ZN(n21481) );
  NAND2_X1 U17995 ( .A1(n14479), .A2(n15823), .ZN(n21320) );
  OAI22_X1 U17996 ( .A1(n21481), .A2(n14481), .B1(n14480), .B2(n21320), .ZN(
        n14456) );
  AOI21_X1 U17997 ( .B1(n21418), .B2(n21555), .A(n14456), .ZN(n14457) );
  OAI211_X1 U17998 ( .C1(n21558), .C2(n14742), .A(n14458), .B(n14457), .ZN(
        P1_U3094) );
  AOI22_X1 U17999 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n14478), .B1(DATAI_26_), 
        .B2(n14437), .ZN(n21546) );
  NAND2_X1 U18000 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14463) );
  AOI22_X1 U18001 ( .A1(DATAI_18_), .A2(n14437), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n14478), .ZN(n21602) );
  INV_X1 U18002 ( .A(n21602), .ZN(n21543) );
  INV_X1 U18003 ( .A(n21597), .ZN(n21472) );
  NAND2_X1 U18004 ( .A1(n14479), .A2(n14460), .ZN(n21308) );
  OAI22_X1 U18005 ( .A1(n21472), .A2(n14481), .B1(n14480), .B2(n21308), .ZN(
        n14461) );
  AOI21_X1 U18006 ( .B1(n21418), .B2(n21543), .A(n14461), .ZN(n14462) );
  OAI211_X1 U18007 ( .C1(n21546), .C2(n14742), .A(n14463), .B(n14462), .ZN(
        P1_U3091) );
  AOI22_X1 U18008 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n14478), .B1(DATAI_31_), 
        .B2(n14437), .ZN(n21570) );
  NAND2_X1 U18009 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14467) );
  AOI22_X1 U18010 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n14478), .B1(DATAI_23_), 
        .B2(n14437), .ZN(n21637) );
  INV_X1 U18011 ( .A(n21637), .ZN(n21563) );
  INV_X1 U18012 ( .A(n15846), .ZN(n14771) );
  INV_X1 U18013 ( .A(n21627), .ZN(n21490) );
  NAND2_X1 U18014 ( .A1(n14479), .A2(n14464), .ZN(n21328) );
  OAI22_X1 U18015 ( .A1(n21490), .A2(n14481), .B1(n14480), .B2(n21328), .ZN(
        n14465) );
  AOI21_X1 U18016 ( .B1(n21418), .B2(n21563), .A(n14465), .ZN(n14466) );
  OAI211_X1 U18017 ( .C1(n21570), .C2(n14742), .A(n14467), .B(n14466), .ZN(
        P1_U3096) );
  AOI22_X1 U18018 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n14478), .B1(DATAI_27_), 
        .B2(n14437), .ZN(n21550) );
  NAND2_X1 U18019 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14472) );
  AOI22_X1 U18020 ( .A1(DATAI_19_), .A2(n14437), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n14478), .ZN(n21608) );
  INV_X1 U18021 ( .A(n21608), .ZN(n21547) );
  INV_X1 U18022 ( .A(n21603), .ZN(n21475) );
  NAND2_X1 U18023 ( .A1(n14479), .A2(n14469), .ZN(n21312) );
  OAI22_X1 U18024 ( .A1(n21475), .A2(n14481), .B1(n14480), .B2(n21312), .ZN(
        n14470) );
  AOI21_X1 U18025 ( .B1(n21418), .B2(n21547), .A(n14470), .ZN(n14471) );
  OAI211_X1 U18026 ( .C1(n21550), .C2(n14742), .A(n14472), .B(n14471), .ZN(
        P1_U3092) );
  AOI22_X1 U18027 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n14478), .B1(DATAI_25_), 
        .B2(n14437), .ZN(n21542) );
  NAND2_X1 U18028 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n14476) );
  AOI22_X1 U18029 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n14478), .B1(DATAI_17_), 
        .B2(n14437), .ZN(n21596) );
  INV_X1 U18030 ( .A(n21596), .ZN(n21539) );
  INV_X1 U18031 ( .A(n21591), .ZN(n21469) );
  NAND2_X1 U18032 ( .A1(n14479), .A2(n15395), .ZN(n21304) );
  OAI22_X1 U18033 ( .A1(n21469), .A2(n14481), .B1(n14480), .B2(n21304), .ZN(
        n14474) );
  AOI21_X1 U18034 ( .B1(n21418), .B2(n21539), .A(n14474), .ZN(n14475) );
  OAI211_X1 U18035 ( .C1(n21542), .C2(n14742), .A(n14476), .B(n14475), .ZN(
        P1_U3090) );
  AOI22_X1 U18036 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n14478), .B1(DATAI_28_), 
        .B2(n14437), .ZN(n21554) );
  NAND2_X1 U18037 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14484) );
  AOI22_X1 U18038 ( .A1(DATAI_20_), .A2(n14437), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n14478), .ZN(n21614) );
  INV_X1 U18039 ( .A(n21614), .ZN(n21551) );
  INV_X1 U18040 ( .A(n15857), .ZN(n14561) );
  INV_X1 U18041 ( .A(n21609), .ZN(n21478) );
  NAND2_X1 U18042 ( .A1(n14479), .A2(n12636), .ZN(n21316) );
  OAI22_X1 U18043 ( .A1(n21478), .A2(n14481), .B1(n14480), .B2(n21316), .ZN(
        n14482) );
  AOI21_X1 U18044 ( .B1(n21418), .B2(n21551), .A(n14482), .ZN(n14483) );
  OAI211_X1 U18045 ( .C1(n21554), .C2(n14742), .A(n14484), .B(n14483), .ZN(
        P1_U3093) );
  INV_X1 U18046 ( .A(n14485), .ZN(n14487) );
  INV_X1 U18047 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n18227) );
  NOR2_X1 U18048 ( .A1(n9824), .A2(n18590), .ZN(n14486) );
  OAI21_X1 U18049 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n14487), .A(n14486), .ZN(
        n14488) );
  OAI21_X1 U18050 ( .B1(n14489), .B2(n18586), .A(n14488), .ZN(P3_U2686) );
  INV_X1 U18051 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n20153) );
  NAND2_X1 U18052 ( .A1(n14490), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14631) );
  NOR2_X1 U18053 ( .A1(n14631), .A2(n14632), .ZN(n14630) );
  OAI211_X1 U18054 ( .C1(n14630), .C2(n14491), .A(n16757), .B(n14419), .ZN(
        n14497) );
  AND2_X1 U18055 ( .A1(n14492), .A2(n14493), .ZN(n14494) );
  OR2_X1 U18056 ( .A1(n14494), .A2(n14424), .ZN(n20155) );
  INV_X1 U18057 ( .A(n20155), .ZN(n14495) );
  NAND2_X1 U18058 ( .A1(n14495), .A2(n16760), .ZN(n14496) );
  OAI211_X1 U18059 ( .C1(n16760), .C2(n20153), .A(n14497), .B(n14496), .ZN(
        P2_U2878) );
  NAND2_X1 U18060 ( .A1(n20911), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20055) );
  INV_X1 U18061 ( .A(n20055), .ZN(n14499) );
  AOI21_X1 U18062 ( .B1(n14499), .B2(n20966), .A(n14498), .ZN(n14503) );
  INV_X1 U18063 ( .A(n14500), .ZN(n14501) );
  OAI211_X1 U18064 ( .C1(n14504), .C2(n14501), .A(n20963), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n14502) );
  OAI211_X1 U18065 ( .C1(n14504), .C2(n14503), .A(n14502), .B(n20177), .ZN(
        P2_U3177) );
  INV_X1 U18066 ( .A(n21747), .ZN(n14515) );
  INV_X1 U18067 ( .A(n21740), .ZN(n14511) );
  INV_X1 U18068 ( .A(n21453), .ZN(n21526) );
  NOR2_X1 U18069 ( .A1(n21584), .A2(n21426), .ZN(n14507) );
  NAND2_X1 U18070 ( .A1(n21586), .A2(n21426), .ZN(n21742) );
  INV_X1 U18071 ( .A(n21742), .ZN(n14506) );
  MUX2_X1 U18072 ( .A(n14507), .B(n14506), .S(n21186), .Z(n14508) );
  AOI21_X1 U18073 ( .B1(n14511), .B2(n21526), .A(n14508), .ZN(n14510) );
  NAND2_X1 U18074 ( .A1(n14515), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n14509) );
  OAI21_X1 U18075 ( .B1(n14515), .B2(n14510), .A(n14509), .ZN(P1_U3477) );
  AOI22_X1 U18076 ( .A1(n14512), .A2(n21586), .B1(n21192), .B2(n14511), .ZN(
        n14514) );
  NAND2_X1 U18077 ( .A1(n14515), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14513) );
  OAI21_X1 U18078 ( .B1(n14515), .B2(n14514), .A(n14513), .ZN(P1_U3476) );
  XNOR2_X1 U18079 ( .A(n9710), .B(n10550), .ZN(n17335) );
  INV_X1 U18080 ( .A(n14700), .ZN(n16899) );
  NAND2_X1 U18081 ( .A1(n17490), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14516) );
  OAI21_X1 U18082 ( .B1(n17490), .B2(n18784), .A(n14516), .ZN(n20278) );
  AOI222_X1 U18083 ( .A1(n17335), .A2(n16899), .B1(n20226), .B2(
        P2_EAX_REG_12__SCAN_IN), .C1(n14625), .C2(n20278), .ZN(n14517) );
  INV_X1 U18084 ( .A(n14517), .ZN(P2_U2907) );
  AOI22_X1 U18085 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14522) );
  AOI22_X1 U18086 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14521) );
  AOI22_X1 U18087 ( .A1(n17705), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14520) );
  INV_X1 U18088 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14518) );
  OR2_X1 U18089 ( .A1(n18545), .A2(n14518), .ZN(n14519) );
  AND4_X1 U18090 ( .A1(n14522), .A2(n14521), .A3(n14520), .A4(n14519), .ZN(
        n14529) );
  AOI22_X1 U18091 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14528) );
  AOI22_X1 U18092 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14526) );
  AOI22_X1 U18093 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14525) );
  AOI22_X1 U18094 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14524) );
  NAND2_X1 U18095 ( .A1(n17762), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n14523) );
  AND4_X1 U18096 ( .A1(n14526), .A2(n14525), .A3(n14524), .A4(n14523), .ZN(
        n14527) );
  AND3_X1 U18097 ( .A1(n14529), .A2(n14528), .A3(n14527), .ZN(n17545) );
  INV_X1 U18098 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18701) );
  NOR2_X1 U18099 ( .A1(n18701), .A2(n14530), .ZN(n18647) );
  INV_X1 U18100 ( .A(n18647), .ZN(n14532) );
  OAI21_X1 U18101 ( .B1(n18677), .B2(n18701), .A(n14530), .ZN(n14531) );
  AOI22_X1 U18102 ( .A1(n14532), .A2(n14531), .B1(n18648), .B2(
        BUF2_REG_4__SCAN_IN), .ZN(n14534) );
  NAND2_X1 U18103 ( .A1(n18653), .A2(BUF2_REG_20__SCAN_IN), .ZN(n14533) );
  OAI211_X1 U18104 ( .C1(n17545), .C2(n18638), .A(n14534), .B(n14533), .ZN(
        P3_U2715) );
  XOR2_X1 U18105 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n14535), .Z(
        n14600) );
  XNOR2_X1 U18106 ( .A(n14600), .B(n14599), .ZN(n14640) );
  NAND2_X1 U18107 ( .A1(n17891), .A2(n16297), .ZN(n16334) );
  NAND2_X1 U18108 ( .A1(n16334), .A2(n14541), .ZN(n17925) );
  INV_X1 U18109 ( .A(n17925), .ZN(n14620) );
  AND2_X1 U18110 ( .A1(n13800), .A2(n14536), .ZN(n14538) );
  OR2_X1 U18111 ( .A1(n14538), .A2(n14537), .ZN(n21109) );
  NAND2_X1 U18112 ( .A1(n17906), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n14636) );
  INV_X1 U18113 ( .A(n14539), .ZN(n17888) );
  OR2_X1 U18114 ( .A1(n17886), .A2(n17888), .ZN(n14540) );
  AND2_X1 U18115 ( .A1(n14540), .A2(n16296), .ZN(n16325) );
  OAI21_X1 U18116 ( .B1(n16297), .B2(n14541), .A(n16325), .ZN(n14618) );
  NAND2_X1 U18117 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14618), .ZN(
        n14542) );
  OAI211_X1 U18118 ( .C1(n21174), .C2(n21109), .A(n14636), .B(n14542), .ZN(
        n14543) );
  AOI21_X1 U18119 ( .B1(n14620), .B2(n14544), .A(n14543), .ZN(n14545) );
  OAI21_X1 U18120 ( .B1(n14640), .B2(n21175), .A(n14545), .ZN(P1_U3028) );
  INV_X1 U18121 ( .A(n14546), .ZN(n14558) );
  INV_X1 U18122 ( .A(n14647), .ZN(n14648) );
  INV_X1 U18123 ( .A(n14548), .ZN(n14550) );
  INV_X1 U18124 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n14549) );
  NAND2_X1 U18125 ( .A1(n14550), .A2(n14549), .ZN(n14551) );
  NAND2_X1 U18126 ( .A1(n14648), .A2(n14551), .ZN(n21065) );
  NAND2_X1 U18127 ( .A1(n21641), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14553) );
  NAND2_X1 U18128 ( .A1(n15379), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n14552) );
  OAI211_X1 U18129 ( .C1(n14554), .C2(n13764), .A(n14553), .B(n14552), .ZN(
        n14555) );
  MUX2_X1 U18130 ( .A(n21065), .B(n14555), .S(n15565), .Z(n14556) );
  AOI21_X1 U18131 ( .B1(n14547), .B2(n15043), .A(n14556), .ZN(n14559) );
  NAND2_X1 U18132 ( .A1(n14546), .A2(n14559), .ZN(n14560) );
  AND2_X1 U18133 ( .A1(n14646), .A2(n14560), .ZN(n21062) );
  INV_X1 U18134 ( .A(n21062), .ZN(n14587) );
  OAI222_X1 U18135 ( .A1(n14587), .A2(n15897), .B1(n15901), .B2(n14561), .C1(
        n15899), .C2(n21145), .ZN(P1_U2900) );
  AOI21_X1 U18136 ( .B1(n14563), .B2(n14562), .A(n10415), .ZN(n17352) );
  NAND2_X1 U18137 ( .A1(n17352), .A2(n16760), .ZN(n14567) );
  NAND2_X1 U18138 ( .A1(n14565), .A2(n14564), .ZN(n14593) );
  OAI211_X1 U18139 ( .C1(n14565), .C2(n14564), .A(n14593), .B(n16757), .ZN(
        n14566) );
  OAI211_X1 U18140 ( .C1(n16760), .C2(n14568), .A(n14567), .B(n14566), .ZN(
        P2_U2876) );
  XNOR2_X1 U18141 ( .A(n14570), .B(n18966), .ZN(n19327) );
  OAI21_X1 U18142 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n14572), .A(
        n14571), .ZN(n14573) );
  INV_X1 U18143 ( .A(n14573), .ZN(n19324) );
  INV_X1 U18144 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14577) );
  OR2_X1 U18145 ( .A1(n19125), .A2(n19069), .ZN(n18388) );
  NOR2_X1 U18146 ( .A1(n19068), .A2(n18388), .ZN(n18373) );
  NAND2_X1 U18147 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18373), .ZN(
        n18363) );
  INV_X1 U18148 ( .A(n18363), .ZN(n18352) );
  NAND2_X1 U18149 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18352), .ZN(
        n18351) );
  NOR2_X1 U18150 ( .A1(n14577), .A2(n18351), .ZN(n18325) );
  AOI21_X1 U18151 ( .B1(n14577), .B2(n18351), .A(n18325), .ZN(n18344) );
  AOI21_X1 U18152 ( .B1(n19404), .B2(n14574), .A(n19096), .ZN(n19035) );
  INV_X1 U18153 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19036) );
  NOR2_X1 U18154 ( .A1(n14574), .A2(n19036), .ZN(n18341) );
  OAI211_X1 U18155 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18341), .A(
        n19801), .B(n19024), .ZN(n14576) );
  INV_X2 U18156 ( .A(n19110), .ZN(n19302) );
  NAND2_X1 U18157 ( .A1(n19302), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n14575) );
  OAI211_X1 U18158 ( .C1(n14577), .C2(n19035), .A(n14576), .B(n14575), .ZN(
        n14578) );
  AOI21_X1 U18159 ( .B1(n18344), .B2(n19122), .A(n14578), .ZN(n14579) );
  OAI21_X1 U18160 ( .B1(n14570), .B2(n19004), .A(n14579), .ZN(n14580) );
  AOI21_X1 U18161 ( .B1(n19324), .B2(n19121), .A(n14580), .ZN(n14581) );
  OAI21_X1 U18162 ( .B1(n19327), .B2(n19034), .A(n14581), .ZN(P3_U2822) );
  INV_X2 U18163 ( .A(n16760), .ZN(n20204) );
  MUX2_X1 U18164 ( .A(n14582), .B(n16619), .S(n20204), .Z(n14583) );
  OAI21_X1 U18165 ( .B1(n20921), .B2(n16752), .A(n14583), .ZN(P2_U2885) );
  OR2_X1 U18166 ( .A1(n14537), .A2(n14585), .ZN(n14586) );
  NAND2_X1 U18167 ( .A1(n14584), .A2(n14586), .ZN(n21056) );
  OAI222_X1 U18168 ( .A1(n21056), .A2(n15821), .B1(n21116), .B2(n13003), .C1(
        n15817), .C2(n14587), .ZN(P1_U2868) );
  INV_X1 U18169 ( .A(n14589), .ZN(n14588) );
  NAND2_X1 U18170 ( .A1(n10415), .A2(n14588), .ZN(n14702) );
  NAND2_X1 U18171 ( .A1(n14590), .A2(n14589), .ZN(n14591) );
  NAND2_X1 U18172 ( .A1(n14702), .A2(n14591), .ZN(n17338) );
  INV_X1 U18173 ( .A(n14593), .ZN(n14596) );
  NOR2_X1 U18174 ( .A1(n14593), .A2(n14592), .ZN(n14707) );
  INV_X1 U18175 ( .A(n14707), .ZN(n14594) );
  OAI211_X1 U18176 ( .C1(n14596), .C2(n14595), .A(n14594), .B(n16757), .ZN(
        n14598) );
  NAND2_X1 U18177 ( .A1(n20204), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14597) );
  OAI211_X1 U18178 ( .C1(n17338), .C2(n20204), .A(n14598), .B(n14597), .ZN(
        P2_U2875) );
  AOI22_X1 U18179 ( .A1(n14600), .A2(n14599), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14535), .ZN(n14603) );
  XNOR2_X1 U18180 ( .A(n14601), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14602) );
  XNOR2_X1 U18181 ( .A(n14603), .B(n14602), .ZN(n14623) );
  INV_X1 U18182 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21667) );
  NOR2_X1 U18183 ( .A1(n17899), .A2(n21667), .ZN(n14617) );
  AOI21_X1 U18184 ( .B1(n17870), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n14617), .ZN(n14604) );
  OAI21_X1 U18185 ( .B1(n21065), .B2(n17877), .A(n14604), .ZN(n14605) );
  AOI21_X1 U18186 ( .B1(n21062), .B2(n17882), .A(n14605), .ZN(n14606) );
  OAI21_X1 U18187 ( .B1(n14623), .B2(n20989), .A(n14606), .ZN(P1_U2995) );
  NOR2_X1 U18188 ( .A1(n20204), .A2(n10780), .ZN(n14607) );
  AOI21_X1 U18189 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n20204), .A(n14607), .ZN(
        n14608) );
  OAI21_X1 U18190 ( .B1(n17499), .B2(n16752), .A(n14608), .ZN(P2_U2887) );
  XOR2_X1 U18191 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n16894), .Z(n14615)
         );
  AND2_X1 U18192 ( .A1(n14609), .A2(n14610), .ZN(n14612) );
  OR2_X1 U18193 ( .A1(n14612), .A2(n14611), .ZN(n17153) );
  MUX2_X1 U18194 ( .A(n17153), .B(n14613), .S(n20204), .Z(n14614) );
  OAI21_X1 U18195 ( .B1(n14615), .B2(n16752), .A(n14614), .ZN(P2_U2882) );
  NOR2_X1 U18196 ( .A1(n21174), .A2(n21056), .ZN(n14616) );
  AOI211_X1 U18197 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n14618), .A(
        n14617), .B(n14616), .ZN(n14622) );
  INV_X1 U18198 ( .A(n17887), .ZN(n14619) );
  OAI211_X1 U18199 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n14620), .B(n14619), .ZN(n14621) );
  OAI211_X1 U18200 ( .C1(n14623), .C2(n21175), .A(n14622), .B(n14621), .ZN(
        P1_U3027) );
  AOI21_X1 U18201 ( .B1(n14624), .B2(n14431), .A(n9828), .ZN(n20128) );
  INV_X1 U18202 ( .A(n20128), .ZN(n14627) );
  AOI22_X1 U18203 ( .A1(n14625), .A2(n16768), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n20226), .ZN(n14626) );
  OAI21_X1 U18204 ( .B1(n14627), .B2(n14700), .A(n14626), .ZN(P2_U2905) );
  NAND2_X1 U18205 ( .A1(n14253), .A2(n14628), .ZN(n14629) );
  NAND2_X1 U18206 ( .A1(n14492), .A2(n14629), .ZN(n17386) );
  NOR2_X1 U18207 ( .A1(n17386), .A2(n20204), .ZN(n14634) );
  AOI211_X1 U18208 ( .C1(n14632), .C2(n14631), .A(n16752), .B(n14630), .ZN(
        n14633) );
  AOI211_X1 U18209 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n20204), .A(n14634), .B(
        n14633), .ZN(n14635) );
  INV_X1 U18210 ( .A(n14635), .ZN(P2_U2879) );
  OAI21_X1 U18211 ( .B1(n17885), .B2(n21069), .A(n14636), .ZN(n14638) );
  NOR2_X1 U18212 ( .A1(n21073), .A2(n16117), .ZN(n14637) );
  AOI211_X1 U18213 ( .C1(n17880), .C2(n21066), .A(n14638), .B(n14637), .ZN(
        n14639) );
  OAI21_X1 U18214 ( .B1(n20989), .B2(n14640), .A(n14639), .ZN(P1_U2996) );
  OAI21_X1 U18215 ( .B1(n14641), .B2(n14642), .A(n16755), .ZN(n20127) );
  AOI211_X1 U18216 ( .C1(n14643), .C2(n14705), .A(n16752), .B(n16759), .ZN(
        n14644) );
  AOI21_X1 U18217 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n20204), .A(n14644), .ZN(
        n14645) );
  OAI21_X1 U18218 ( .B1(n20204), .B2(n20127), .A(n14645), .ZN(P2_U2873) );
  INV_X1 U18219 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n14652) );
  AND2_X2 U18220 ( .A1(n14647), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14747) );
  INV_X1 U18221 ( .A(n14747), .ZN(n14650) );
  INV_X1 U18222 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n21044) );
  NAND2_X1 U18223 ( .A1(n14648), .A2(n21044), .ZN(n14649) );
  NAND2_X1 U18224 ( .A1(n14650), .A2(n14649), .ZN(n21051) );
  AOI22_X1 U18225 ( .A1(n21051), .A2(n15562), .B1(n15378), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n14651) );
  OAI21_X1 U18226 ( .B1(n15329), .B2(n14652), .A(n14651), .ZN(n14653) );
  NAND2_X1 U18227 ( .A1(n14655), .A2(n14646), .ZN(n14656) );
  AND2_X1 U18228 ( .A1(n14768), .A2(n14656), .ZN(n21106) );
  INV_X1 U18229 ( .A(n21106), .ZN(n14658) );
  OAI222_X1 U18230 ( .A1(n14658), .A2(n15897), .B1(n15901), .B2(n14657), .C1(
        n15899), .C2(n14652), .ZN(P1_U2899) );
  NOR2_X1 U18231 ( .A1(n21581), .A2(n21186), .ZN(n14660) );
  OAI21_X1 U18232 ( .B1(n21494), .B2(n14660), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14662) );
  AOI21_X1 U18233 ( .B1(n14662), .B2(n14661), .A(n21584), .ZN(n21745) );
  INV_X1 U18234 ( .A(n21745), .ZN(n14663) );
  NOR2_X1 U18235 ( .A1(n14663), .A2(n21581), .ZN(n14664) );
  NAND2_X1 U18236 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21574) );
  NOR2_X1 U18237 ( .A1(n21574), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n14667) );
  NAND2_X1 U18238 ( .A1(n14693), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n14674) );
  OR2_X1 U18239 ( .A1(n21391), .A2(n10013), .ZN(n21527) );
  INV_X1 U18240 ( .A(n21527), .ZN(n21573) );
  INV_X1 U18241 ( .A(n14666), .ZN(n21423) );
  NOR3_X1 U18242 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21422), .A3(
        n21574), .ZN(n14671) );
  AOI21_X1 U18243 ( .B1(n21573), .B2(n21423), .A(n14671), .ZN(n14669) );
  INV_X1 U18244 ( .A(n14667), .ZN(n14668) );
  OAI22_X1 U18245 ( .A1(n14669), .A2(n21584), .B1(n14668), .B2(n21641), .ZN(
        n14670) );
  INV_X1 U18246 ( .A(n14671), .ZN(n14694) );
  OAI22_X1 U18247 ( .A1(n21484), .A2(n14695), .B1(n21324), .B2(n14694), .ZN(
        n14672) );
  AOI21_X1 U18248 ( .B1(n16393), .B2(n21559), .A(n14672), .ZN(n14673) );
  OAI211_X1 U18249 ( .C1(n21562), .C2(n21524), .A(n14674), .B(n14673), .ZN(
        P1_U3143) );
  NAND2_X1 U18250 ( .A1(n14693), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n14677) );
  OAI22_X1 U18251 ( .A1(n21490), .A2(n14695), .B1(n21328), .B2(n14694), .ZN(
        n14675) );
  AOI21_X1 U18252 ( .B1(n16393), .B2(n21563), .A(n14675), .ZN(n14676) );
  OAI211_X1 U18253 ( .C1(n21570), .C2(n21524), .A(n14677), .B(n14676), .ZN(
        P1_U3144) );
  NAND2_X1 U18254 ( .A1(n14693), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n14680) );
  OAI22_X1 U18255 ( .A1(n21472), .A2(n14695), .B1(n21308), .B2(n14694), .ZN(
        n14678) );
  AOI21_X1 U18256 ( .B1(n16393), .B2(n21543), .A(n14678), .ZN(n14679) );
  OAI211_X1 U18257 ( .C1(n21546), .C2(n21524), .A(n14680), .B(n14679), .ZN(
        P1_U3139) );
  NAND2_X1 U18258 ( .A1(n14693), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n14683) );
  OAI22_X1 U18259 ( .A1(n21478), .A2(n14695), .B1(n21316), .B2(n14694), .ZN(
        n14681) );
  AOI21_X1 U18260 ( .B1(n16393), .B2(n21551), .A(n14681), .ZN(n14682) );
  OAI211_X1 U18261 ( .C1(n21554), .C2(n21524), .A(n14683), .B(n14682), .ZN(
        P1_U3141) );
  NAND2_X1 U18262 ( .A1(n14693), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n14686) );
  OAI22_X1 U18263 ( .A1(n21466), .A2(n14695), .B1(n21291), .B2(n14694), .ZN(
        n14684) );
  AOI21_X1 U18264 ( .B1(n16393), .B2(n21523), .A(n14684), .ZN(n14685) );
  OAI211_X1 U18265 ( .C1(n21538), .C2(n21524), .A(n14686), .B(n14685), .ZN(
        P1_U3137) );
  NAND2_X1 U18266 ( .A1(n14693), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n14689) );
  OAI22_X1 U18267 ( .A1(n21469), .A2(n14695), .B1(n21304), .B2(n14694), .ZN(
        n14687) );
  AOI21_X1 U18268 ( .B1(n16393), .B2(n21539), .A(n14687), .ZN(n14688) );
  OAI211_X1 U18269 ( .C1(n21542), .C2(n21524), .A(n14689), .B(n14688), .ZN(
        P1_U3138) );
  NAND2_X1 U18270 ( .A1(n14693), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n14692) );
  OAI22_X1 U18271 ( .A1(n21481), .A2(n14695), .B1(n21320), .B2(n14694), .ZN(
        n14690) );
  AOI21_X1 U18272 ( .B1(n16393), .B2(n21555), .A(n14690), .ZN(n14691) );
  OAI211_X1 U18273 ( .C1(n21558), .C2(n21524), .A(n14692), .B(n14691), .ZN(
        P1_U3142) );
  NAND2_X1 U18274 ( .A1(n14693), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n14698) );
  OAI22_X1 U18275 ( .A1(n21475), .A2(n14695), .B1(n21312), .B2(n14694), .ZN(
        n14696) );
  AOI21_X1 U18276 ( .B1(n16393), .B2(n21547), .A(n14696), .ZN(n14697) );
  OAI211_X1 U18277 ( .C1(n21550), .C2(n21524), .A(n14698), .B(n14697), .ZN(
        P1_U3140) );
  OAI21_X1 U18278 ( .B1(n9828), .B2(n10561), .A(n14847), .ZN(n20108) );
  OAI222_X1 U18279 ( .A1(n20108), .A2(n14700), .B1(n16897), .B2(n13235), .C1(
        n14699), .C2(n20232), .ZN(P2_U2904) );
  INV_X1 U18280 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n14710) );
  AND2_X1 U18281 ( .A1(n14702), .A2(n14701), .ZN(n14703) );
  OR2_X1 U18282 ( .A1(n14703), .A2(n14641), .ZN(n17323) );
  INV_X1 U18283 ( .A(n17323), .ZN(n14704) );
  NAND2_X1 U18284 ( .A1(n14704), .A2(n16760), .ZN(n14709) );
  OAI211_X1 U18285 ( .C1(n14707), .C2(n14706), .A(n16757), .B(n14705), .ZN(
        n14708) );
  OAI211_X1 U18286 ( .C1(n16760), .C2(n14710), .A(n14709), .B(n14708), .ZN(
        P2_U2874) );
  NAND2_X1 U18287 ( .A1(n14742), .A2(n21586), .ZN(n14711) );
  NOR2_X1 U18288 ( .A1(n21338), .A2(n21453), .ZN(n14713) );
  NAND2_X1 U18289 ( .A1(n14712), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21533) );
  INV_X1 U18290 ( .A(n21533), .ZN(n21190) );
  NOR2_X1 U18291 ( .A1(n21393), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21258) );
  OR2_X1 U18292 ( .A1(n14712), .A2(n21641), .ZN(n21395) );
  INV_X1 U18293 ( .A(n21395), .ZN(n21455) );
  INV_X1 U18294 ( .A(n14713), .ZN(n14716) );
  INV_X1 U18295 ( .A(n14714), .ZN(n14715) );
  OR2_X1 U18296 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14715), .ZN(
        n14741) );
  AOI22_X1 U18297 ( .A1(n14717), .A2(n14716), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n14741), .ZN(n14718) );
  OAI21_X1 U18298 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n21393), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n21255) );
  NAND3_X1 U18299 ( .A1(n21529), .A2(n14718), .A3(n21255), .ZN(n14740) );
  NAND2_X1 U18300 ( .A1(n14740), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n14721) );
  INV_X1 U18301 ( .A(n21538), .ZN(n21587) );
  OAI22_X1 U18302 ( .A1(n14742), .A2(n21590), .B1(n14741), .B2(n21291), .ZN(
        n14719) );
  AOI21_X1 U18303 ( .B1(n21384), .B2(n21587), .A(n14719), .ZN(n14720) );
  OAI211_X1 U18304 ( .C1(n14746), .C2(n21466), .A(n14721), .B(n14720), .ZN(
        P1_U3081) );
  NAND2_X1 U18305 ( .A1(n14740), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n14724) );
  INV_X1 U18306 ( .A(n21558), .ZN(n21617) );
  OAI22_X1 U18307 ( .A1(n14742), .A2(n21620), .B1(n14741), .B2(n21320), .ZN(
        n14722) );
  AOI21_X1 U18308 ( .B1(n21384), .B2(n21617), .A(n14722), .ZN(n14723) );
  OAI211_X1 U18309 ( .C1(n14746), .C2(n21481), .A(n14724), .B(n14723), .ZN(
        P1_U3086) );
  NAND2_X1 U18310 ( .A1(n14740), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n14727) );
  INV_X1 U18311 ( .A(n21542), .ZN(n21593) );
  OAI22_X1 U18312 ( .A1(n14742), .A2(n21596), .B1(n14741), .B2(n21304), .ZN(
        n14725) );
  AOI21_X1 U18313 ( .B1(n21384), .B2(n21593), .A(n14725), .ZN(n14726) );
  OAI211_X1 U18314 ( .C1(n14746), .C2(n21469), .A(n14727), .B(n14726), .ZN(
        P1_U3082) );
  NAND2_X1 U18315 ( .A1(n14740), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n14730) );
  INV_X1 U18316 ( .A(n21562), .ZN(n21623) );
  OAI22_X1 U18317 ( .A1(n14742), .A2(n21626), .B1(n14741), .B2(n21324), .ZN(
        n14728) );
  AOI21_X1 U18318 ( .B1(n21384), .B2(n21623), .A(n14728), .ZN(n14729) );
  OAI211_X1 U18319 ( .C1(n14746), .C2(n21484), .A(n14730), .B(n14729), .ZN(
        P1_U3087) );
  NAND2_X1 U18320 ( .A1(n14740), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n14733) );
  INV_X1 U18321 ( .A(n21546), .ZN(n21599) );
  OAI22_X1 U18322 ( .A1(n14742), .A2(n21602), .B1(n14741), .B2(n21308), .ZN(
        n14731) );
  AOI21_X1 U18323 ( .B1(n21384), .B2(n21599), .A(n14731), .ZN(n14732) );
  OAI211_X1 U18324 ( .C1(n14746), .C2(n21472), .A(n14733), .B(n14732), .ZN(
        P1_U3083) );
  NAND2_X1 U18325 ( .A1(n14740), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n14736) );
  INV_X1 U18326 ( .A(n21570), .ZN(n21631) );
  OAI22_X1 U18327 ( .A1(n14742), .A2(n21637), .B1(n14741), .B2(n21328), .ZN(
        n14734) );
  AOI21_X1 U18328 ( .B1(n21384), .B2(n21631), .A(n14734), .ZN(n14735) );
  OAI211_X1 U18329 ( .C1(n14746), .C2(n21490), .A(n14736), .B(n14735), .ZN(
        P1_U3088) );
  NAND2_X1 U18330 ( .A1(n14740), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n14739) );
  INV_X1 U18331 ( .A(n21550), .ZN(n21605) );
  OAI22_X1 U18332 ( .A1(n14742), .A2(n21608), .B1(n14741), .B2(n21312), .ZN(
        n14737) );
  AOI21_X1 U18333 ( .B1(n21384), .B2(n21605), .A(n14737), .ZN(n14738) );
  OAI211_X1 U18334 ( .C1(n14746), .C2(n21475), .A(n14739), .B(n14738), .ZN(
        P1_U3084) );
  NAND2_X1 U18335 ( .A1(n14740), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n14745) );
  INV_X1 U18336 ( .A(n21554), .ZN(n21611) );
  OAI22_X1 U18337 ( .A1(n14742), .A2(n21614), .B1(n14741), .B2(n21316), .ZN(
        n14743) );
  AOI21_X1 U18338 ( .B1(n21384), .B2(n21611), .A(n14743), .ZN(n14744) );
  OAI211_X1 U18339 ( .C1(n14746), .C2(n21478), .A(n14745), .B(n14744), .ZN(
        P1_U3085) );
  INV_X1 U18340 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n14749) );
  OAI21_X1 U18341 ( .B1(n14747), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n14753), .ZN(n21039) );
  AOI22_X1 U18342 ( .A1(n21039), .A2(n15562), .B1(n15378), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n14748) );
  OAI21_X1 U18343 ( .B1(n15329), .B2(n14749), .A(n14748), .ZN(n14750) );
  INV_X1 U18344 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n14757) );
  INV_X1 U18345 ( .A(n14753), .ZN(n14755) );
  INV_X1 U18346 ( .A(n14952), .ZN(n14754) );
  OAI21_X1 U18347 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n14755), .A(
        n14754), .ZN(n21025) );
  AOI22_X1 U18348 ( .A1(n15562), .A2(n21025), .B1(n15378), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14756) );
  OAI21_X1 U18349 ( .B1(n15329), .B2(n14757), .A(n14756), .ZN(n14758) );
  INV_X1 U18350 ( .A(n14758), .ZN(n14759) );
  OAI21_X1 U18351 ( .B1(n9812), .B2(n14761), .A(n15759), .ZN(n17867) );
  NOR2_X1 U18352 ( .A1(n14763), .A2(n14764), .ZN(n14765) );
  OR2_X1 U18353 ( .A1(n14762), .A2(n14765), .ZN(n21020) );
  INV_X1 U18354 ( .A(n21020), .ZN(n14766) );
  AOI22_X1 U18355 ( .A1(n14766), .A2(n21111), .B1(n15818), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n14767) );
  OAI21_X1 U18356 ( .B1(n17867), .B2(n15817), .A(n14767), .ZN(P1_U2865) );
  XOR2_X1 U18357 ( .A(n14769), .B(n14768), .Z(n21037) );
  INV_X1 U18358 ( .A(n21037), .ZN(n14775) );
  OAI222_X1 U18359 ( .A1(n15897), .A2(n14775), .B1(n15901), .B2(n14770), .C1(
        n15899), .C2(n14749), .ZN(P1_U2898) );
  OAI222_X1 U18360 ( .A1(n17867), .A2(n15897), .B1(n15901), .B2(n14771), .C1(
        n15899), .C2(n14757), .ZN(P1_U2897) );
  AND2_X1 U18361 ( .A1(n14772), .A2(n14773), .ZN(n14774) );
  OR2_X1 U18362 ( .A1(n14774), .A2(n14763), .ZN(n21027) );
  OAI222_X1 U18363 ( .A1(n21027), .A2(n15821), .B1(n21116), .B2(n13013), .C1(
        n15817), .C2(n14775), .ZN(P1_U2866) );
  NAND2_X1 U18364 ( .A1(n10322), .A2(n20196), .ZN(n14776) );
  XOR2_X1 U18365 ( .A(n14776), .B(n17150), .Z(n14787) );
  INV_X1 U18366 ( .A(n17153), .ZN(n17420) );
  INV_X1 U18367 ( .A(n14778), .ZN(n14779) );
  XNOR2_X1 U18368 ( .A(n14777), .B(n14779), .ZN(n17419) );
  NAND2_X1 U18369 ( .A1(n17419), .A2(n20185), .ZN(n14783) );
  AOI21_X1 U18370 ( .B1(n20169), .B2(P2_EBX_REG_5__SCAN_IN), .A(n20167), .ZN(
        n14780) );
  OAI21_X1 U18371 ( .B1(n17148), .B2(n20180), .A(n14780), .ZN(n14781) );
  AOI21_X1 U18372 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n20186), .A(
        n14781), .ZN(n14782) );
  OAI211_X1 U18373 ( .C1(n20165), .C2(n14784), .A(n14783), .B(n14782), .ZN(
        n14785) );
  AOI21_X1 U18374 ( .B1(n17420), .B2(n20129), .A(n14785), .ZN(n14786) );
  OAI21_X1 U18375 ( .B1(n14787), .B2(n20177), .A(n14786), .ZN(P2_U2850) );
  INV_X1 U18376 ( .A(n14788), .ZN(n14790) );
  NAND2_X1 U18377 ( .A1(n14790), .A2(n14789), .ZN(n16921) );
  XNOR2_X1 U18378 ( .A(n14888), .B(n14887), .ZN(n14822) );
  AOI21_X1 U18379 ( .B1(n14794), .B2(n10553), .A(n14793), .ZN(n16688) );
  INV_X1 U18380 ( .A(n16688), .ZN(n14798) );
  NAND2_X1 U18381 ( .A1(n16415), .A2(n17190), .ZN(n14795) );
  NAND2_X1 U18382 ( .A1(n20167), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n14814) );
  OAI211_X1 U18383 ( .C1(n16412), .C2(n17187), .A(n14795), .B(n14814), .ZN(
        n14796) );
  INV_X1 U18384 ( .A(n14796), .ZN(n14797) );
  OAI21_X1 U18385 ( .B1(n14822), .B2(n17181), .A(n14799), .ZN(P2_U2987) );
  AOI22_X1 U18386 ( .A1(n14800), .A2(P2_FLUSH_REG_SCAN_IN), .B1(
        P2_STATE2_REG_3__SCAN_IN), .B2(n11573), .ZN(n14801) );
  OAI21_X1 U18387 ( .B1(n14803), .B2(n14802), .A(n14801), .ZN(n17478) );
  AOI211_X1 U18388 ( .C1(n16640), .C2(n14804), .A(n16614), .B(n20147), .ZN(
        n16627) );
  AOI21_X1 U18389 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20147), .A(
        n16627), .ZN(n17468) );
  MUX2_X1 U18390 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n16640), .S(
        n10322), .Z(n17467) );
  INV_X1 U18391 ( .A(n17467), .ZN(n14805) );
  NOR3_X1 U18392 ( .A1(n17468), .A2(n14805), .A3(n11055), .ZN(n14809) );
  INV_X1 U18393 ( .A(n14806), .ZN(n14807) );
  INV_X1 U18394 ( .A(n20911), .ZN(n17476) );
  OAI22_X1 U18395 ( .A1(n20921), .A2(n17484), .B1(n14807), .B2(n17476), .ZN(
        n14808) );
  OAI21_X1 U18396 ( .B1(n14809), .B2(n14808), .A(n17478), .ZN(n14810) );
  OAI21_X1 U18397 ( .B1(n17478), .B2(n14811), .A(n14810), .ZN(P2_U3599) );
  AOI21_X1 U18398 ( .B1(n14813), .B2(n9772), .A(n14914), .ZN(n16788) );
  INV_X1 U18399 ( .A(n16788), .ZN(n14820) );
  INV_X1 U18400 ( .A(n14814), .ZN(n14817) );
  NOR3_X1 U18401 ( .A1(n14815), .A2(n17362), .A3(n14887), .ZN(n14816) );
  AOI211_X1 U18402 ( .C1(n14818), .C2(n14887), .A(n14817), .B(n14816), .ZN(
        n14819) );
  OAI21_X1 U18403 ( .B1(n14820), .B2(n17444), .A(n14819), .ZN(n14821) );
  INV_X1 U18404 ( .A(n14823), .ZN(n14827) );
  AOI22_X1 U18405 ( .A1(n14827), .A2(n14826), .B1(n14825), .B2(n14824), .ZN(
        n17006) );
  NAND2_X1 U18406 ( .A1(n17415), .A2(n14828), .ZN(n14833) );
  NAND2_X1 U18407 ( .A1(n10181), .A2(n14835), .ZN(n14829) );
  NAND2_X1 U18408 ( .A1(n17303), .A2(n14829), .ZN(n17292) );
  AOI21_X1 U18409 ( .B1(n10458), .B2(n14830), .A(n17292), .ZN(n14831) );
  OAI21_X1 U18410 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17452), .A(
        n14856), .ZN(n14844) );
  NOR2_X1 U18411 ( .A1(n14835), .A2(n17370), .ZN(n17291) );
  NOR2_X1 U18412 ( .A1(n14836), .A2(n14837), .ZN(n14838) );
  OR2_X1 U18413 ( .A1(n16528), .A2(n14838), .ZN(n20084) );
  NOR2_X1 U18414 ( .A1(n9833), .A2(n14840), .ZN(n14841) );
  OR2_X1 U18415 ( .A1(n14839), .A2(n14841), .ZN(n20083) );
  INV_X1 U18416 ( .A(n20083), .ZN(n16870) );
  NOR2_X1 U18417 ( .A1(n17149), .A2(n20877), .ZN(n16998) );
  AOI21_X1 U18418 ( .B1(n16870), .B2(n17461), .A(n16998), .ZN(n14842) );
  OAI21_X1 U18419 ( .B1(n20084), .B2(n17429), .A(n14842), .ZN(n14843) );
  AOI21_X1 U18420 ( .B1(n14845), .B2(n16753), .A(n14836), .ZN(n17012) );
  AND2_X1 U18421 ( .A1(n14847), .A2(n14846), .ZN(n14848) );
  OR2_X1 U18422 ( .A1(n14848), .A2(n9833), .ZN(n20096) );
  NAND2_X1 U18423 ( .A1(n20167), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n17010) );
  OAI21_X1 U18424 ( .B1(n20096), .B2(n17444), .A(n17010), .ZN(n14851) );
  AOI211_X1 U18425 ( .C1(n17012), .C2(n17456), .A(n14851), .B(n14850), .ZN(
        n14855) );
  XNOR2_X1 U18426 ( .A(n14852), .B(n14853), .ZN(n17008) );
  NAND2_X1 U18427 ( .A1(n17008), .A2(n17412), .ZN(n14854) );
  OAI211_X1 U18428 ( .C1(n14856), .C2(n17007), .A(n14855), .B(n14854), .ZN(
        P2_U3030) );
  NAND2_X1 U18429 ( .A1(n14859), .A2(n14858), .ZN(n14860) );
  XNOR2_X1 U18430 ( .A(n14861), .B(n14860), .ZN(n14883) );
  OAI21_X1 U18431 ( .B1(n14863), .B2(n14865), .A(n14864), .ZN(n16725) );
  NOR2_X1 U18432 ( .A1(n17149), .A2(n20883), .ZN(n14874) );
  NOR2_X1 U18433 ( .A1(n16489), .A2(n17175), .ZN(n14866) );
  AOI211_X1 U18434 ( .C1(n17172), .C2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n14874), .B(n14866), .ZN(n14867) );
  OAI21_X1 U18435 ( .B1(n16725), .B2(n17166), .A(n14867), .ZN(n14868) );
  AOI21_X1 U18436 ( .B1(n14881), .B2(n17196), .A(n14868), .ZN(n14869) );
  OAI21_X1 U18437 ( .B1(n14883), .B2(n17181), .A(n14869), .ZN(P2_U2993) );
  NOR2_X1 U18438 ( .A1(n16725), .A2(n17429), .ZN(n14880) );
  OR2_X1 U18439 ( .A1(n14871), .A2(n14872), .ZN(n14873) );
  NAND2_X1 U18440 ( .A1(n14870), .A2(n14873), .ZN(n16831) );
  INV_X1 U18441 ( .A(n14874), .ZN(n14878) );
  NAND2_X1 U18442 ( .A1(n14875), .A2(n17300), .ZN(n14876) );
  MUX2_X1 U18443 ( .A(n14876), .B(n17241), .S(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .Z(n14877) );
  OAI211_X1 U18444 ( .C1(n16831), .C2(n17444), .A(n14878), .B(n14877), .ZN(
        n14879) );
  AOI211_X1 U18445 ( .C1(n14881), .C2(n17454), .A(n14880), .B(n14879), .ZN(
        n14882) );
  OAI21_X1 U18446 ( .B1(n14883), .B2(n17458), .A(n14882), .ZN(P2_U3025) );
  NAND2_X1 U18447 ( .A1(n14884), .A2(n14792), .ZN(n14886) );
  XOR2_X1 U18448 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14889), .Z(
        n14890) );
  XNOR2_X1 U18449 ( .A(n14891), .B(n14890), .ZN(n14925) );
  XNOR2_X1 U18450 ( .A(n14892), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14923) );
  OAI21_X1 U18451 ( .B1(n14793), .B2(n14893), .A(n12505), .ZN(n16682) );
  NOR2_X1 U18452 ( .A1(n17149), .A2(n14894), .ZN(n14918) );
  NOR2_X1 U18453 ( .A1(n16398), .A2(n17175), .ZN(n14895) );
  AOI211_X1 U18454 ( .C1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17172), .A(
        n14918), .B(n14895), .ZN(n14896) );
  OAI21_X1 U18455 ( .B1(n16682), .B2(n17166), .A(n14896), .ZN(n14897) );
  AOI21_X1 U18456 ( .B1(n17196), .B2(n14923), .A(n14897), .ZN(n14898) );
  OAI21_X1 U18457 ( .B1(n14925), .B2(n17181), .A(n14898), .ZN(P2_U2986) );
  INV_X1 U18458 ( .A(n14919), .ZN(n14905) );
  NAND2_X1 U18459 ( .A1(n20167), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n16911) );
  OAI211_X1 U18460 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(n14903), .B(n14902), .ZN(
        n14904) );
  OAI211_X1 U18461 ( .C1(n14905), .C2(n9968), .A(n16911), .B(n14904), .ZN(
        n14906) );
  NAND2_X1 U18462 ( .A1(n9811), .A2(n17454), .ZN(n14911) );
  OAI211_X1 U18463 ( .C1(n16919), .C2(n17458), .A(n14912), .B(n14911), .ZN(
        P2_U3017) );
  NOR2_X1 U18464 ( .A1(n16682), .A2(n17429), .ZN(n14922) );
  NAND2_X1 U18465 ( .A1(n14914), .A2(n14913), .ZN(n14916) );
  OR2_X1 U18466 ( .A1(n14914), .A2(n14913), .ZN(n14915) );
  NOR2_X1 U18467 ( .A1(n9770), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14917) );
  OAI21_X1 U18468 ( .B1(n16402), .B2(n17444), .A(n14920), .ZN(n14921) );
  OAI21_X1 U18469 ( .B1(n14925), .B2(n17458), .A(n14924), .ZN(P2_U3018) );
  INV_X1 U18470 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n14927) );
  XNOR2_X1 U18471 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n14952), .ZN(
        n16124) );
  AOI22_X1 U18472 ( .A1(n15562), .A2(n16124), .B1(n15378), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14926) );
  OAI21_X1 U18473 ( .B1(n15329), .B2(n14927), .A(n14926), .ZN(n14940) );
  AOI22_X1 U18474 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14931) );
  AOI22_X1 U18475 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9705), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14930) );
  AOI22_X1 U18476 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14929) );
  AOI22_X1 U18477 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14928) );
  NAND4_X1 U18478 ( .A1(n14931), .A2(n14930), .A3(n14929), .A4(n14928), .ZN(
        n14937) );
  AOI22_X1 U18479 ( .A1(n15354), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14935) );
  AOI22_X1 U18480 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15361), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14934) );
  AOI22_X1 U18481 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15341), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14933) );
  AOI22_X1 U18482 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14932) );
  NAND4_X1 U18483 ( .A1(n14935), .A2(n14934), .A3(n14933), .A4(n14932), .ZN(
        n14936) );
  NOR2_X1 U18484 ( .A1(n14937), .A2(n14936), .ZN(n14938) );
  NOR2_X1 U18485 ( .A1(n15082), .A2(n14938), .ZN(n14939) );
  NOR2_X1 U18486 ( .A1(n14940), .A2(n14939), .ZN(n15760) );
  AOI22_X1 U18487 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9694), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14945) );
  AOI22_X1 U18488 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14944) );
  AOI22_X1 U18489 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14943) );
  AOI22_X1 U18490 ( .A1(n15360), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14942) );
  NAND4_X1 U18491 ( .A1(n14945), .A2(n14944), .A3(n14943), .A4(n14942), .ZN(
        n14951) );
  AOI22_X1 U18492 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n15202), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14949) );
  AOI22_X1 U18493 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15361), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14948) );
  AOI22_X1 U18494 ( .A1(n15362), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15341), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14947) );
  AOI22_X1 U18495 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14946) );
  NAND4_X1 U18496 ( .A1(n14949), .A2(n14948), .A3(n14947), .A4(n14946), .ZN(
        n14950) );
  NOR2_X1 U18497 ( .A1(n14951), .A2(n14950), .ZN(n14955) );
  XNOR2_X1 U18498 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n14975), .ZN(
        n21012) );
  INV_X1 U18499 ( .A(n21012), .ZN(n14953) );
  AOI22_X1 U18500 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n15378), .B1(
        n15562), .B2(n14953), .ZN(n14954) );
  OAI21_X1 U18501 ( .B1(n15082), .B2(n14955), .A(n14954), .ZN(n14958) );
  INV_X1 U18502 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n14956) );
  NOR2_X1 U18503 ( .A1(n15329), .A2(n14956), .ZN(n14957) );
  AOI22_X1 U18504 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9704), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14963) );
  AOI22_X1 U18505 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9705), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14962) );
  AOI22_X1 U18506 ( .A1(n15360), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15361), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14961) );
  AOI22_X1 U18507 ( .A1(n15362), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15341), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14960) );
  NAND4_X1 U18508 ( .A1(n14963), .A2(n14962), .A3(n14961), .A4(n14960), .ZN(
        n14969) );
  AOI22_X1 U18509 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14967) );
  AOI22_X1 U18510 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14966) );
  AOI22_X1 U18511 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12558), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14965) );
  AOI22_X1 U18512 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14964) );
  NAND4_X1 U18513 ( .A1(n14967), .A2(n14966), .A3(n14965), .A4(n14964), .ZN(
        n14968) );
  NOR2_X1 U18514 ( .A1(n14969), .A2(n14968), .ZN(n14974) );
  OAI21_X1 U18515 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n21426), .A(
        n21641), .ZN(n14970) );
  OAI21_X1 U18516 ( .B1(n15329), .B2(n14971), .A(n14970), .ZN(n14972) );
  INV_X1 U18517 ( .A(n14972), .ZN(n14973) );
  OAI21_X1 U18518 ( .B1(n15375), .B2(n14974), .A(n14973), .ZN(n14985) );
  NAND2_X1 U18519 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14978) );
  INV_X1 U18520 ( .A(n14980), .ZN(n14982) );
  INV_X1 U18521 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14981) );
  NAND2_X1 U18522 ( .A1(n14982), .A2(n14981), .ZN(n14983) );
  NAND2_X1 U18523 ( .A1(n15153), .A2(n14983), .ZN(n16039) );
  OR2_X1 U18524 ( .A1(n16039), .A2(n15565), .ZN(n14984) );
  NAND2_X1 U18525 ( .A1(n14985), .A2(n14984), .ZN(n15660) );
  INV_X1 U18526 ( .A(n15660), .ZN(n15085) );
  AOI22_X1 U18527 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14989) );
  AOI22_X1 U18528 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9705), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14988) );
  AOI22_X1 U18529 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14987) );
  AOI22_X1 U18530 ( .A1(n15361), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14986) );
  NAND4_X1 U18531 ( .A1(n14989), .A2(n14988), .A3(n14987), .A4(n14986), .ZN(
        n14995) );
  AOI22_X1 U18532 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14993) );
  AOI22_X1 U18533 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14992) );
  AOI22_X1 U18534 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15341), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14991) );
  AOI22_X1 U18535 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14990) );
  NAND4_X1 U18536 ( .A1(n14993), .A2(n14992), .A3(n14991), .A4(n14990), .ZN(
        n14994) );
  NOR2_X1 U18537 ( .A1(n14995), .A2(n14994), .ZN(n14996) );
  NOR2_X1 U18538 ( .A1(n15082), .A2(n14996), .ZN(n15729) );
  INV_X1 U18539 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n15886) );
  INV_X1 U18540 ( .A(n14997), .ZN(n14999) );
  INV_X1 U18541 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n14998) );
  NAND2_X1 U18542 ( .A1(n14999), .A2(n14998), .ZN(n15000) );
  NAND2_X1 U18543 ( .A1(n15063), .A2(n15000), .ZN(n16098) );
  AOI22_X1 U18544 ( .A1(n16098), .A2(n15562), .B1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n15378), .ZN(n15001) );
  OAI21_X1 U18545 ( .B1(n15329), .B2(n15886), .A(n15001), .ZN(n15698) );
  AOI22_X1 U18546 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(n9704), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15005) );
  AOI22_X1 U18547 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9705), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15004) );
  AOI22_X1 U18548 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15003) );
  AOI22_X1 U18549 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12558), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15002) );
  NAND4_X1 U18550 ( .A1(n15005), .A2(n15004), .A3(n15003), .A4(n15002), .ZN(
        n15011) );
  AOI22_X1 U18551 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15009) );
  AOI22_X1 U18552 ( .A1(n15362), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15008) );
  AOI22_X1 U18553 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15361), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15007) );
  AOI22_X1 U18554 ( .A1(n15341), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15006) );
  NAND4_X1 U18555 ( .A1(n15009), .A2(n15008), .A3(n15007), .A4(n15006), .ZN(
        n15010) );
  OAI21_X1 U18556 ( .B1(n15011), .B2(n15010), .A(n15043), .ZN(n15016) );
  NAND2_X1 U18557 ( .A1(n15379), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n15015) );
  INV_X1 U18558 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15012) );
  XNOR2_X1 U18559 ( .A(n15031), .B(n15012), .ZN(n16050) );
  NAND2_X1 U18560 ( .A1(n16050), .A2(n15562), .ZN(n15014) );
  NAND2_X1 U18561 ( .A1(n15378), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15013) );
  NAND4_X1 U18562 ( .A1(n15016), .A2(n15015), .A3(n15014), .A4(n15013), .ZN(
        n15673) );
  AOI22_X1 U18563 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9694), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15020) );
  AOI22_X1 U18564 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15019) );
  AOI22_X1 U18565 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15341), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15018) );
  AOI22_X1 U18566 ( .A1(n15361), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12558), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15017) );
  NAND4_X1 U18567 ( .A1(n15020), .A2(n15019), .A3(n15018), .A4(n15017), .ZN(
        n15026) );
  AOI22_X1 U18568 ( .A1(n15362), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15024) );
  AOI22_X1 U18569 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15023) );
  AOI22_X1 U18570 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15022) );
  AOI22_X1 U18571 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15021) );
  NAND4_X1 U18572 ( .A1(n15024), .A2(n15023), .A3(n15022), .A4(n15021), .ZN(
        n15025) );
  NOR2_X1 U18573 ( .A1(n15026), .A2(n15025), .ZN(n15034) );
  NAND2_X1 U18574 ( .A1(n15379), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n15033) );
  INV_X1 U18575 ( .A(n15027), .ZN(n15029) );
  NAND2_X1 U18576 ( .A1(n15029), .A2(n15028), .ZN(n15030) );
  NAND2_X1 U18577 ( .A1(n15031), .A2(n15030), .ZN(n16060) );
  AOI22_X1 U18578 ( .A1(n16060), .A2(n15562), .B1(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n15378), .ZN(n15032) );
  OAI211_X1 U18579 ( .C1(n15034), .C2(n15082), .A(n15033), .B(n15032), .ZN(
        n15686) );
  OAI211_X1 U18580 ( .C1(n15729), .C2(n15698), .A(n15673), .B(n15686), .ZN(
        n15067) );
  AOI22_X1 U18581 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15202), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15038) );
  AOI22_X1 U18582 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15037) );
  AOI22_X1 U18583 ( .A1(n12617), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15361), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15036) );
  AOI22_X1 U18584 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15341), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15035) );
  NAND4_X1 U18585 ( .A1(n15038), .A2(n15037), .A3(n15036), .A4(n15035), .ZN(
        n15045) );
  AOI22_X1 U18586 ( .A1(n15362), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15042) );
  AOI22_X1 U18587 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15041) );
  AOI22_X1 U18588 ( .A1(n15360), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15040) );
  AOI22_X1 U18589 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15039) );
  NAND4_X1 U18590 ( .A1(n15042), .A2(n15041), .A3(n15040), .A4(n15039), .ZN(
        n15044) );
  OAI21_X1 U18591 ( .B1(n15045), .B2(n15044), .A(n15043), .ZN(n15052) );
  NAND2_X1 U18592 ( .A1(n15379), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n15051) );
  NAND2_X1 U18593 ( .A1(n15378), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15050) );
  INV_X1 U18594 ( .A(n15063), .ZN(n15046) );
  NAND2_X1 U18595 ( .A1(n15046), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15048) );
  INV_X1 U18596 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15047) );
  XNOR2_X1 U18597 ( .A(n15048), .B(n15047), .ZN(n16077) );
  NAND2_X1 U18598 ( .A1(n16077), .A2(n15562), .ZN(n15049) );
  NAND4_X1 U18599 ( .A1(n15052), .A2(n15051), .A3(n15050), .A4(n15049), .ZN(
        n15701) );
  AOI22_X1 U18600 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12718), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15056) );
  AOI22_X1 U18601 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15055) );
  AOI22_X1 U18602 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15361), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15054) );
  AOI22_X1 U18603 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15053) );
  NAND4_X1 U18604 ( .A1(n15056), .A2(n15055), .A3(n15054), .A4(n15053), .ZN(
        n15062) );
  AOI22_X1 U18605 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n15202), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15060) );
  AOI22_X1 U18606 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15059) );
  AOI22_X1 U18607 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12581), .B1(
        n15341), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15058) );
  AOI22_X1 U18608 ( .A1(n12617), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12558), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15057) );
  NAND4_X1 U18609 ( .A1(n15060), .A2(n15059), .A3(n15058), .A4(n15057), .ZN(
        n15061) );
  NOR2_X1 U18610 ( .A1(n15062), .A2(n15061), .ZN(n15066) );
  NAND2_X1 U18611 ( .A1(n15379), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n15065) );
  INV_X1 U18612 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16087) );
  XNOR2_X1 U18613 ( .A(n15063), .B(n16087), .ZN(n16086) );
  AOI22_X1 U18614 ( .A1(n16086), .A2(n15562), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n15378), .ZN(n15064) );
  OAI211_X1 U18615 ( .C1(n15066), .C2(n15082), .A(n15065), .B(n15064), .ZN(
        n15716) );
  NAND2_X1 U18616 ( .A1(n15701), .A2(n15716), .ZN(n15671) );
  NOR2_X1 U18617 ( .A1(n15067), .A2(n15671), .ZN(n15084) );
  AOI22_X1 U18618 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15071) );
  AOI22_X1 U18619 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15070) );
  AOI22_X1 U18620 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15069) );
  AOI22_X1 U18621 ( .A1(n15361), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15068) );
  NAND4_X1 U18622 ( .A1(n15071), .A2(n15070), .A3(n15069), .A4(n15068), .ZN(
        n15077) );
  AOI22_X1 U18623 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9705), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15075) );
  AOI22_X1 U18624 ( .A1(n12617), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15074) );
  AOI22_X1 U18625 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15341), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15073) );
  AOI22_X1 U18626 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15072) );
  NAND4_X1 U18627 ( .A1(n15075), .A2(n15074), .A3(n15073), .A4(n15072), .ZN(
        n15076) );
  NOR2_X1 U18628 ( .A1(n15077), .A2(n15076), .ZN(n15083) );
  NAND2_X1 U18629 ( .A1(n15379), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n15081) );
  INV_X1 U18630 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15078) );
  XNOR2_X1 U18631 ( .A(n15079), .B(n15078), .ZN(n16111) );
  AOI22_X1 U18632 ( .A1(n16111), .A2(n15562), .B1(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n15378), .ZN(n15080) );
  OAI211_X1 U18633 ( .C1(n15083), .C2(n15082), .A(n15081), .B(n15080), .ZN(
        n15740) );
  AND2_X1 U18634 ( .A1(n15084), .A2(n15740), .ZN(n15657) );
  INV_X1 U18635 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16001) );
  OR3_X4 U18636 ( .A1(n15191), .A2(n15186), .A3(n16001), .ZN(n15122) );
  INV_X1 U18637 ( .A(n15088), .ZN(n15106) );
  INV_X1 U18638 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15574) );
  NAND2_X1 U18639 ( .A1(n15106), .A2(n15574), .ZN(n15089) );
  NAND2_X1 U18640 ( .A1(n15226), .A2(n15089), .ZN(n15981) );
  OR2_X1 U18641 ( .A1(n15981), .A2(n15565), .ZN(n15104) );
  AOI22_X1 U18642 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9694), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15093) );
  AOI22_X1 U18643 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15092) );
  AOI22_X1 U18644 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15091) );
  AOI22_X1 U18645 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12558), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15090) );
  NAND4_X1 U18646 ( .A1(n15093), .A2(n15092), .A3(n15091), .A4(n15090), .ZN(
        n15099) );
  AOI22_X1 U18647 ( .A1(n15362), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15097) );
  AOI22_X1 U18648 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15361), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15096) );
  AOI22_X1 U18649 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15341), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15095) );
  AOI22_X1 U18650 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15094) );
  NAND4_X1 U18651 ( .A1(n15097), .A2(n15096), .A3(n15095), .A4(n15094), .ZN(
        n15098) );
  NOR2_X1 U18652 ( .A1(n15099), .A2(n15098), .ZN(n15102) );
  OAI21_X1 U18653 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21426), .A(
        n21641), .ZN(n15101) );
  NAND2_X1 U18654 ( .A1(n15379), .A2(P1_EAX_REG_22__SCAN_IN), .ZN(n15100) );
  OAI211_X1 U18655 ( .C1(n15375), .C2(n15102), .A(n15101), .B(n15100), .ZN(
        n15103) );
  NAND2_X1 U18656 ( .A1(n15122), .A2(n15588), .ZN(n15105) );
  NAND2_X1 U18657 ( .A1(n15106), .A2(n15105), .ZN(n15992) );
  OR2_X1 U18658 ( .A1(n15992), .A2(n15565), .ZN(n15121) );
  AOI22_X1 U18659 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15110) );
  AOI22_X1 U18660 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15109) );
  AOI22_X1 U18661 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15361), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15108) );
  AOI22_X1 U18662 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9686), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15107) );
  NAND4_X1 U18663 ( .A1(n15110), .A2(n15109), .A3(n15108), .A4(n15107), .ZN(
        n15116) );
  AOI22_X1 U18664 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15114) );
  AOI22_X1 U18665 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15113) );
  AOI22_X1 U18666 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15341), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15112) );
  AOI22_X1 U18667 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12558), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15111) );
  NAND4_X1 U18668 ( .A1(n15114), .A2(n15113), .A3(n15112), .A4(n15111), .ZN(
        n15115) );
  NOR2_X1 U18669 ( .A1(n15116), .A2(n15115), .ZN(n15119) );
  AOI21_X1 U18670 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15588), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n15117) );
  AOI21_X1 U18671 ( .B1(n15379), .B2(P1_EAX_REG_21__SCAN_IN), .A(n15117), .ZN(
        n15118) );
  OAI21_X1 U18672 ( .B1(n15375), .B2(n15119), .A(n15118), .ZN(n15120) );
  OAI21_X1 U18673 ( .B1(n15191), .B2(n15186), .A(n16001), .ZN(n15123) );
  AND2_X1 U18674 ( .A1(n15123), .A2(n15122), .ZN(n15999) );
  NAND2_X1 U18675 ( .A1(n15999), .A2(n15562), .ZN(n15138) );
  AOI22_X1 U18676 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n9694), .B1(
        n12581), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15127) );
  AOI22_X1 U18677 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n15202), .B1(
        n9705), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15126) );
  AOI22_X1 U18678 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15125) );
  AOI22_X1 U18679 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n9706), .B1(
        n12558), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15124) );
  NAND4_X1 U18680 ( .A1(n15127), .A2(n15126), .A3(n15125), .A4(n15124), .ZN(
        n15133) );
  AOI22_X1 U18681 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n15354), .B1(
        n12718), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15131) );
  AOI22_X1 U18682 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15130) );
  AOI22_X1 U18683 ( .A1(n15360), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15361), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15129) );
  AOI22_X1 U18684 ( .A1(n15341), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15128) );
  NAND4_X1 U18685 ( .A1(n15131), .A2(n15130), .A3(n15129), .A4(n15128), .ZN(
        n15132) );
  NOR2_X1 U18686 ( .A1(n15133), .A2(n15132), .ZN(n15136) );
  OAI21_X1 U18687 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21426), .A(
        n21641), .ZN(n15135) );
  NAND2_X1 U18688 ( .A1(n15379), .A2(P1_EAX_REG_20__SCAN_IN), .ZN(n15134) );
  OAI211_X1 U18689 ( .C1(n15375), .C2(n15136), .A(n15135), .B(n15134), .ZN(
        n15137) );
  NAND2_X1 U18690 ( .A1(n15138), .A2(n15137), .ZN(n15564) );
  AOI22_X1 U18691 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15142) );
  AOI22_X1 U18692 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15141) );
  AOI22_X1 U18693 ( .A1(n15362), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15341), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15140) );
  AOI22_X1 U18694 ( .A1(n15361), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12558), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15139) );
  NAND4_X1 U18695 ( .A1(n15142), .A2(n15141), .A3(n15140), .A4(n15139), .ZN(
        n15148) );
  AOI22_X1 U18696 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n9704), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15146) );
  AOI22_X1 U18697 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15145) );
  AOI22_X1 U18698 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15144) );
  AOI22_X1 U18699 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15143) );
  NAND4_X1 U18700 ( .A1(n15146), .A2(n15145), .A3(n15144), .A4(n15143), .ZN(
        n15147) );
  OAI21_X1 U18701 ( .B1(n15148), .B2(n15147), .A(n15348), .ZN(n15156) );
  INV_X1 U18702 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n15150) );
  INV_X1 U18703 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15152) );
  OAI22_X1 U18704 ( .A1(n15329), .A2(n15150), .B1(n15152), .B2(n15149), .ZN(
        n15151) );
  INV_X1 U18705 ( .A(n15151), .ZN(n15155) );
  XNOR2_X1 U18706 ( .A(n15153), .B(n15152), .ZN(n16028) );
  NAND2_X1 U18707 ( .A1(n16028), .A2(n15562), .ZN(n15154) );
  NOR2_X1 U18708 ( .A1(n15564), .A2(n15639), .ZN(n15195) );
  AOI22_X1 U18709 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n9703), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15160) );
  AOI22_X1 U18710 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15159) );
  AOI22_X1 U18711 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15158) );
  AOI22_X1 U18712 ( .A1(n15341), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15157) );
  NAND4_X1 U18713 ( .A1(n15160), .A2(n15159), .A3(n15158), .A4(n15157), .ZN(
        n15166) );
  AOI22_X1 U18714 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15164) );
  AOI22_X1 U18715 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15163) );
  AOI22_X1 U18716 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15162) );
  AOI22_X1 U18717 ( .A1(n15361), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12558), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15161) );
  NAND4_X1 U18718 ( .A1(n15164), .A2(n15163), .A3(n15162), .A4(n15161), .ZN(
        n15165) );
  OR2_X1 U18719 ( .A1(n15166), .A2(n15165), .ZN(n15167) );
  NAND2_X1 U18720 ( .A1(n15348), .A2(n15167), .ZN(n15171) );
  INV_X1 U18721 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n15168) );
  INV_X1 U18722 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15188) );
  OAI22_X1 U18723 ( .A1(n15329), .A2(n15168), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15188), .ZN(n15169) );
  INV_X1 U18724 ( .A(n15169), .ZN(n15170) );
  NAND2_X1 U18725 ( .A1(n15171), .A2(n15170), .ZN(n15563) );
  AOI22_X1 U18726 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15175) );
  AOI22_X1 U18727 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9705), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15174) );
  AOI22_X1 U18728 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15173) );
  AOI22_X1 U18729 ( .A1(n12617), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15172) );
  NAND4_X1 U18730 ( .A1(n15175), .A2(n15174), .A3(n15173), .A4(n15172), .ZN(
        n15181) );
  AOI22_X1 U18731 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15179) );
  AOI22_X1 U18732 ( .A1(n15360), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15361), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15178) );
  AOI22_X1 U18733 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15341), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15177) );
  AOI22_X1 U18734 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15176) );
  NAND4_X1 U18735 ( .A1(n15179), .A2(n15178), .A3(n15177), .A4(n15176), .ZN(
        n15180) );
  OR2_X1 U18736 ( .A1(n15181), .A2(n15180), .ZN(n15182) );
  NAND2_X1 U18737 ( .A1(n15348), .A2(n15182), .ZN(n15185) );
  OAI22_X1 U18738 ( .A1(n15329), .A2(n13423), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15186), .ZN(n15183) );
  INV_X1 U18739 ( .A(n15183), .ZN(n15184) );
  NAND2_X1 U18740 ( .A1(n15185), .A2(n15184), .ZN(n15566) );
  NAND3_X1 U18741 ( .A1(n15563), .A2(n15566), .A3(n15565), .ZN(n15193) );
  XNOR2_X1 U18742 ( .A(n15191), .B(n15186), .ZN(n16008) );
  INV_X1 U18743 ( .A(n15187), .ZN(n15189) );
  NAND2_X1 U18744 ( .A1(n15189), .A2(n15188), .ZN(n15190) );
  NAND2_X1 U18745 ( .A1(n15191), .A2(n15190), .ZN(n16016) );
  NAND3_X1 U18746 ( .A1(n16008), .A2(n15562), .A3(n16016), .ZN(n15192) );
  NAND2_X1 U18747 ( .A1(n15193), .A2(n15192), .ZN(n15194) );
  NAND4_X1 U18748 ( .A1(n15569), .A2(n15584), .A3(n15195), .A4(n15194), .ZN(
        n15196) );
  XNOR2_X1 U18749 ( .A(n15226), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15969) );
  NAND2_X1 U18750 ( .A1(n15969), .A2(n15562), .ZN(n15225) );
  AOI22_X1 U18751 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n9704), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15201) );
  AOI22_X1 U18752 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15200) );
  AOI22_X1 U18753 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15199) );
  AOI22_X1 U18754 ( .A1(n15341), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15198) );
  NAND4_X1 U18755 ( .A1(n15201), .A2(n15200), .A3(n15199), .A4(n15198), .ZN(
        n15208) );
  AOI22_X1 U18756 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15206) );
  AOI22_X1 U18757 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15205) );
  AOI22_X1 U18758 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15204) );
  AOI22_X1 U18759 ( .A1(n15361), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12558), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15203) );
  NAND4_X1 U18760 ( .A1(n15206), .A2(n15205), .A3(n15204), .A4(n15203), .ZN(
        n15207) );
  NOR2_X1 U18761 ( .A1(n15208), .A2(n15207), .ZN(n15231) );
  AOI22_X1 U18762 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15283), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15212) );
  AOI22_X1 U18763 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15341), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15211) );
  AOI22_X1 U18764 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15210) );
  AOI22_X1 U18765 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15209) );
  NAND4_X1 U18766 ( .A1(n15212), .A2(n15211), .A3(n15210), .A4(n15209), .ZN(
        n15218) );
  AOI22_X1 U18767 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15216) );
  AOI22_X1 U18768 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15215) );
  AOI22_X1 U18769 ( .A1(n12536), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15361), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15214) );
  AOI22_X1 U18770 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15213) );
  NAND4_X1 U18771 ( .A1(n15216), .A2(n15215), .A3(n15214), .A4(n15213), .ZN(
        n15217) );
  NOR2_X1 U18772 ( .A1(n15218), .A2(n15217), .ZN(n15232) );
  XOR2_X1 U18773 ( .A(n15231), .B(n15232), .Z(n15219) );
  NAND2_X1 U18774 ( .A1(n15219), .A2(n15348), .ZN(n15223) );
  NAND2_X1 U18775 ( .A1(n21641), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15220) );
  OAI211_X1 U18776 ( .C1(n15329), .C2(n14079), .A(n15565), .B(n15220), .ZN(
        n15221) );
  INV_X1 U18777 ( .A(n15221), .ZN(n15222) );
  NAND2_X1 U18778 ( .A1(n15223), .A2(n15222), .ZN(n15224) );
  NAND2_X1 U18779 ( .A1(n15225), .A2(n15224), .ZN(n15548) );
  INV_X1 U18780 ( .A(n15228), .ZN(n15229) );
  INV_X1 U18781 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15961) );
  NAND2_X1 U18782 ( .A1(n15229), .A2(n15961), .ZN(n15230) );
  AND2_X1 U18783 ( .A1(n15271), .A2(n15230), .ZN(n15965) );
  NOR2_X1 U18784 ( .A1(n15232), .A2(n15231), .ZN(n15249) );
  AOI22_X1 U18785 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15236) );
  AOI22_X1 U18786 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15235) );
  AOI22_X1 U18787 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15234) );
  AOI22_X1 U18788 ( .A1(n15361), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15233) );
  NAND4_X1 U18789 ( .A1(n15236), .A2(n15235), .A3(n15234), .A4(n15233), .ZN(
        n15242) );
  AOI22_X1 U18790 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n9704), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15240) );
  AOI22_X1 U18791 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15283), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15239) );
  AOI22_X1 U18792 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15238) );
  AOI22_X1 U18793 ( .A1(n15341), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15237) );
  NAND4_X1 U18794 ( .A1(n15240), .A2(n15239), .A3(n15238), .A4(n15237), .ZN(
        n15241) );
  OR2_X1 U18795 ( .A1(n15242), .A2(n15241), .ZN(n15248) );
  INV_X1 U18796 ( .A(n15248), .ZN(n15243) );
  XNOR2_X1 U18797 ( .A(n15249), .B(n15243), .ZN(n15246) );
  NAND2_X1 U18798 ( .A1(n21641), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15244) );
  OAI211_X1 U18799 ( .C1(n15329), .C2(n13427), .A(n15565), .B(n15244), .ZN(
        n15245) );
  AOI21_X1 U18800 ( .B1(n15246), .B2(n15348), .A(n15245), .ZN(n15247) );
  AOI21_X1 U18801 ( .B1(n15965), .B2(n15562), .A(n15247), .ZN(n15534) );
  XNOR2_X1 U18802 ( .A(n15271), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15950) );
  NAND2_X1 U18803 ( .A1(n15950), .A2(n15562), .ZN(n15268) );
  NAND2_X1 U18804 ( .A1(n15249), .A2(n15248), .ZN(n15276) );
  AOI22_X1 U18805 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15283), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15253) );
  AOI22_X1 U18806 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15252) );
  AOI22_X1 U18807 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15251) );
  AOI22_X1 U18808 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15250) );
  NAND4_X1 U18809 ( .A1(n15253), .A2(n15252), .A3(n15251), .A4(n15250), .ZN(
        n15260) );
  AOI22_X1 U18810 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15258) );
  AOI22_X1 U18811 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15361), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15257) );
  AOI22_X1 U18812 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15256) );
  AOI22_X1 U18813 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15255) );
  NAND4_X1 U18814 ( .A1(n15258), .A2(n15257), .A3(n15256), .A4(n15255), .ZN(
        n15259) );
  NOR2_X1 U18815 ( .A1(n15260), .A2(n15259), .ZN(n15277) );
  XOR2_X1 U18816 ( .A(n15276), .B(n15277), .Z(n15261) );
  NAND2_X1 U18817 ( .A1(n15261), .A2(n15348), .ZN(n15266) );
  INV_X1 U18818 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n15263) );
  NAND2_X1 U18819 ( .A1(n21641), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15262) );
  OAI211_X1 U18820 ( .C1(n15329), .C2(n15263), .A(n15565), .B(n15262), .ZN(
        n15264) );
  INV_X1 U18821 ( .A(n15264), .ZN(n15265) );
  NAND2_X1 U18822 ( .A1(n15266), .A2(n15265), .ZN(n15267) );
  NAND2_X1 U18823 ( .A1(n15268), .A2(n15267), .ZN(n15517) );
  INV_X1 U18824 ( .A(n15273), .ZN(n15274) );
  INV_X1 U18825 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15508) );
  NAND2_X1 U18826 ( .A1(n15274), .A2(n15508), .ZN(n15275) );
  NAND2_X1 U18827 ( .A1(n15313), .A2(n15275), .ZN(n15942) );
  NOR2_X1 U18828 ( .A1(n15277), .A2(n15276), .ZN(n15297) );
  AOI22_X1 U18829 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15282) );
  AOI22_X1 U18830 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15281) );
  AOI22_X1 U18831 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15280) );
  AOI22_X1 U18832 ( .A1(n15361), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15279) );
  NAND4_X1 U18833 ( .A1(n15282), .A2(n15281), .A3(n15280), .A4(n15279), .ZN(
        n15289) );
  AOI22_X1 U18834 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n9703), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15287) );
  AOI22_X1 U18835 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15283), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15286) );
  AOI22_X1 U18836 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15285) );
  AOI22_X1 U18837 ( .A1(n15341), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15284) );
  NAND4_X1 U18838 ( .A1(n15287), .A2(n15286), .A3(n15285), .A4(n15284), .ZN(
        n15288) );
  OR2_X1 U18839 ( .A1(n15289), .A2(n15288), .ZN(n15296) );
  XNOR2_X1 U18840 ( .A(n15297), .B(n15296), .ZN(n15293) );
  NAND2_X1 U18841 ( .A1(n21641), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15290) );
  OAI211_X1 U18842 ( .C1(n15329), .C2(n13417), .A(n15565), .B(n15290), .ZN(
        n15291) );
  INV_X1 U18843 ( .A(n15291), .ZN(n15292) );
  OAI21_X1 U18844 ( .B1(n15293), .B2(n15375), .A(n15292), .ZN(n15294) );
  XNOR2_X1 U18845 ( .A(n15313), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15931) );
  NAND2_X1 U18846 ( .A1(n15297), .A2(n15296), .ZN(n15316) );
  AOI22_X1 U18847 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n15354), .B1(
        n12718), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15301) );
  AOI22_X1 U18848 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15300) );
  AOI22_X1 U18849 ( .A1(n15360), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15361), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15299) );
  AOI22_X1 U18850 ( .A1(n15341), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15298) );
  NAND4_X1 U18851 ( .A1(n15301), .A2(n15300), .A3(n15299), .A4(n15298), .ZN(
        n15308) );
  AOI22_X1 U18852 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15202), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15306) );
  AOI22_X1 U18853 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n9694), .B1(n9704), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15305) );
  AOI22_X1 U18854 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15304) );
  AOI22_X1 U18855 ( .A1(n12617), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15303) );
  NAND4_X1 U18856 ( .A1(n15306), .A2(n15305), .A3(n15304), .A4(n15303), .ZN(
        n15307) );
  NOR2_X1 U18857 ( .A1(n15308), .A2(n15307), .ZN(n15317) );
  XOR2_X1 U18858 ( .A(n15316), .B(n15317), .Z(n15311) );
  OAI21_X1 U18859 ( .B1(n21426), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n21641), .ZN(n15309) );
  OAI21_X1 U18860 ( .B1(n15329), .B2(n13835), .A(n15309), .ZN(n15310) );
  AOI21_X1 U18861 ( .B1(n15311), .B2(n15348), .A(n15310), .ZN(n15312) );
  AOI21_X1 U18862 ( .B1(n15931), .B2(n15562), .A(n15312), .ZN(n15490) );
  INV_X1 U18863 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15929) );
  OR2_X2 U18864 ( .A1(n15313), .A2(n15929), .ZN(n15314) );
  INV_X1 U18865 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15481) );
  OR2_X2 U18866 ( .A1(n15314), .A2(n15481), .ZN(n15352) );
  NAND2_X1 U18867 ( .A1(n15314), .A2(n15481), .ZN(n15315) );
  NAND2_X1 U18868 ( .A1(n15352), .A2(n15315), .ZN(n15923) );
  NOR2_X1 U18869 ( .A1(n15317), .A2(n15316), .ZN(n15336) );
  AOI22_X1 U18870 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15321) );
  AOI22_X1 U18871 ( .A1(n15202), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12617), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15320) );
  AOI22_X1 U18872 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15319) );
  AOI22_X1 U18873 ( .A1(n15361), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15318) );
  NAND4_X1 U18874 ( .A1(n15321), .A2(n15320), .A3(n15319), .A4(n15318), .ZN(
        n15327) );
  AOI22_X1 U18875 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n9704), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15325) );
  AOI22_X1 U18876 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15324) );
  AOI22_X1 U18877 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15323) );
  AOI22_X1 U18878 ( .A1(n15341), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15322) );
  NAND4_X1 U18879 ( .A1(n15325), .A2(n15324), .A3(n15323), .A4(n15322), .ZN(
        n15326) );
  OR2_X1 U18880 ( .A1(n15327), .A2(n15326), .ZN(n15335) );
  XNOR2_X1 U18881 ( .A(n15336), .B(n15335), .ZN(n15332) );
  NAND2_X1 U18882 ( .A1(n21641), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15328) );
  OAI211_X1 U18883 ( .C1(n15329), .C2(n13829), .A(n15565), .B(n15328), .ZN(
        n15330) );
  INV_X1 U18884 ( .A(n15330), .ZN(n15331) );
  OAI21_X1 U18885 ( .B1(n15332), .B2(n15375), .A(n15331), .ZN(n15333) );
  XNOR2_X1 U18886 ( .A(n15352), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15469) );
  INV_X1 U18887 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15470) );
  AOI21_X1 U18888 ( .B1(n15470), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n15334) );
  AOI21_X1 U18889 ( .B1(n15379), .B2(P1_EAX_REG_29__SCAN_IN), .A(n15334), .ZN(
        n15351) );
  NAND2_X1 U18890 ( .A1(n15336), .A2(n15335), .ZN(n15369) );
  AOI22_X1 U18891 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9694), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15340) );
  AOI22_X1 U18892 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15339) );
  AOI22_X1 U18893 ( .A1(n12536), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15338) );
  AOI22_X1 U18894 ( .A1(n12581), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15337) );
  NAND4_X1 U18895 ( .A1(n15340), .A2(n15339), .A3(n15338), .A4(n15337), .ZN(
        n15347) );
  AOI22_X1 U18896 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15362), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15345) );
  AOI22_X1 U18897 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15344) );
  AOI22_X1 U18898 ( .A1(n15341), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15343) );
  AOI22_X1 U18899 ( .A1(n15361), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15342) );
  NAND4_X1 U18900 ( .A1(n15345), .A2(n15344), .A3(n15343), .A4(n15342), .ZN(
        n15346) );
  NOR2_X1 U18901 ( .A1(n15347), .A2(n15346), .ZN(n15370) );
  XOR2_X1 U18902 ( .A(n15369), .B(n15370), .Z(n15349) );
  NAND2_X1 U18903 ( .A1(n15349), .A2(n15348), .ZN(n15350) );
  AOI22_X1 U18904 ( .A1(n15469), .A2(n15562), .B1(n15351), .B2(n15350), .ZN(
        n15465) );
  INV_X1 U18905 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15454) );
  XNOR2_X1 U18906 ( .A(n15381), .B(n15454), .ZN(n15907) );
  AOI22_X1 U18907 ( .A1(n15254), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9704), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15359) );
  AOI22_X1 U18908 ( .A1(n9705), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15354), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15358) );
  AOI22_X1 U18909 ( .A1(n12718), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12594), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15357) );
  AOI22_X1 U18910 ( .A1(n15355), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15278), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15356) );
  NAND4_X1 U18911 ( .A1(n15359), .A2(n15358), .A3(n15357), .A4(n15356), .ZN(
        n15368) );
  AOI22_X1 U18912 ( .A1(n12536), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15360), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15366) );
  AOI22_X1 U18913 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15361), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15365) );
  AOI22_X1 U18914 ( .A1(n15362), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15364) );
  AOI22_X1 U18915 ( .A1(n9694), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15197), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15363) );
  NAND4_X1 U18916 ( .A1(n15366), .A2(n15365), .A3(n15364), .A4(n15363), .ZN(
        n15367) );
  NOR2_X1 U18917 ( .A1(n15368), .A2(n15367), .ZN(n15372) );
  NOR2_X1 U18918 ( .A1(n15370), .A2(n15369), .ZN(n15371) );
  XOR2_X1 U18919 ( .A(n15372), .B(n15371), .Z(n15376) );
  AOI21_X1 U18920 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n21641), .A(
        n15562), .ZN(n15374) );
  NAND2_X1 U18921 ( .A1(n15379), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n15373) );
  OAI211_X1 U18922 ( .C1(n15376), .C2(n15375), .A(n15374), .B(n15373), .ZN(
        n15377) );
  OAI21_X1 U18923 ( .B1(n15907), .B2(n15565), .A(n15377), .ZN(n15448) );
  AOI22_X1 U18924 ( .A1(n15379), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n15378), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15380) );
  OR2_X2 U18925 ( .A1(n15381), .A2(n15454), .ZN(n15382) );
  INV_X1 U18926 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15409) );
  XNOR2_X2 U18927 ( .A(n15382), .B(n15409), .ZN(n15453) );
  AOI21_X1 U18928 ( .B1(n17870), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15383), .ZN(n15384) );
  OAI21_X1 U18929 ( .B1(n15453), .B2(n17877), .A(n15384), .ZN(n15385) );
  AOI21_X1 U18930 ( .B1(n15418), .B2(n17882), .A(n15385), .ZN(n15386) );
  OAI21_X1 U18931 ( .B1(n15387), .B2(n20989), .A(n15386), .ZN(P1_U2968) );
  INV_X1 U18932 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15410) );
  OAI22_X1 U18933 ( .A1(n15388), .A2(n15821), .B1(n15410), .B2(n21116), .ZN(
        P1_U2841) );
  NAND2_X1 U18934 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21765), .ZN(n17852) );
  AND2_X1 U18935 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21638), .ZN(n15391) );
  NAND2_X1 U18936 ( .A1(n15562), .A2(n15391), .ZN(n15392) );
  OAI21_X1 U18937 ( .B1(n17852), .B2(n21638), .A(n15392), .ZN(n15393) );
  OR3_X4 U18938 ( .A1(n21757), .A2(n17906), .A3(n15393), .ZN(n21074) );
  NOR2_X1 U18939 ( .A1(n15777), .A2(n15394), .ZN(n15408) );
  NAND2_X1 U18940 ( .A1(n15395), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n15404) );
  AND2_X1 U18941 ( .A1(n21759), .A2(n21426), .ZN(n17846) );
  NOR2_X1 U18942 ( .A1(n15404), .A2(n17846), .ZN(n15396) );
  NAND2_X1 U18943 ( .A1(n21074), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15451) );
  NAND2_X1 U18944 ( .A1(n15418), .A2(n21036), .ZN(n15416) );
  INV_X1 U18945 ( .A(n17846), .ZN(n15397) );
  AOI21_X1 U18946 ( .B1(n12924), .B2(n15398), .A(n15397), .ZN(n15406) );
  NAND2_X2 U18947 ( .A1(n15408), .A2(n15406), .ZN(n21087) );
  NAND2_X1 U18948 ( .A1(n21087), .A2(n21074), .ZN(n15791) );
  INV_X1 U18949 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21706) );
  INV_X1 U18950 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21702) );
  INV_X1 U18951 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21699) );
  INV_X1 U18952 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21674) );
  INV_X1 U18953 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21668) );
  NAND3_X1 U18954 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n21052) );
  NOR2_X1 U18955 ( .A1(n21667), .A2(n21052), .ZN(n21047) );
  NAND2_X1 U18956 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n21047), .ZN(n21028) );
  NOR2_X1 U18957 ( .A1(n21668), .A2(n21028), .ZN(n21029) );
  NAND2_X1 U18958 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n21029), .ZN(n15766) );
  NOR2_X1 U18959 ( .A1(n21674), .A2(n15766), .ZN(n15764) );
  NAND3_X1 U18960 ( .A1(n15764), .A2(P1_REIP_REG_10__SCAN_IN), .A3(
        P1_REIP_REG_9__SCAN_IN), .ZN(n15616) );
  NAND3_X1 U18961 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n15620) );
  NAND2_X1 U18962 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n15399) );
  NOR2_X1 U18963 ( .A1(n15620), .A2(n15399), .ZN(n15601) );
  INV_X1 U18964 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21682) );
  NAND3_X1 U18965 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .ZN(n15689) );
  NOR2_X1 U18966 ( .A1(n21682), .A2(n15689), .ZN(n15618) );
  NAND3_X1 U18967 ( .A1(n15601), .A2(P1_REIP_REG_20__SCAN_IN), .A3(n15618), 
        .ZN(n15400) );
  NOR2_X1 U18968 ( .A1(n15616), .A2(n15400), .ZN(n15590) );
  NAND2_X1 U18969 ( .A1(n15590), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15575) );
  NOR2_X1 U18970 ( .A1(n21699), .A2(n15575), .ZN(n15552) );
  NAND2_X1 U18971 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n15552), .ZN(n15540) );
  NOR2_X1 U18972 ( .A1(n21702), .A2(n15540), .ZN(n15525) );
  NAND2_X1 U18973 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n15525), .ZN(n15506) );
  NOR2_X1 U18974 ( .A1(n21706), .A2(n15506), .ZN(n15507) );
  NAND2_X1 U18975 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n15507), .ZN(n15411) );
  INV_X1 U18976 ( .A(n15411), .ZN(n15401) );
  NAND3_X1 U18977 ( .A1(n21074), .A2(P1_REIP_REG_28__SCAN_IN), .A3(n15401), 
        .ZN(n15402) );
  NAND2_X1 U18978 ( .A1(n15791), .A2(n15402), .ZN(n15483) );
  NAND2_X1 U18979 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n15412) );
  NAND2_X1 U18980 ( .A1(n15791), .A2(n15412), .ZN(n15403) );
  NAND2_X1 U18981 ( .A1(n15483), .A2(n15403), .ZN(n15457) );
  INV_X1 U18982 ( .A(n15404), .ZN(n15405) );
  NOR2_X1 U18983 ( .A1(n15406), .A2(n15405), .ZN(n15407) );
  NAND2_X1 U18984 ( .A1(n15408), .A2(n15407), .ZN(n21089) );
  OAI22_X1 U18985 ( .A1(n21089), .A2(n15410), .B1(n15409), .B2(n21068), .ZN(
        n15414) );
  NOR2_X1 U18986 ( .A1(n21087), .A2(n15411), .ZN(n15482) );
  NAND2_X1 U18987 ( .A1(n15482), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15471) );
  NOR3_X1 U18988 ( .A1(n15471), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n15412), 
        .ZN(n15413) );
  AOI211_X1 U18989 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n15457), .A(n15414), 
        .B(n15413), .ZN(n15415) );
  OAI211_X1 U18990 ( .C1(n15388), .C2(n21086), .A(n15416), .B(n15415), .ZN(
        P1_U2809) );
  AND2_X1 U18991 ( .A1(n15837), .A2(n10088), .ZN(n15417) );
  NAND2_X1 U18992 ( .A1(n15899), .A2(n15417), .ZN(n15822) );
  INV_X1 U18993 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n17937) );
  NOR3_X1 U18994 ( .A1(n15889), .A2(n15837), .A3(n12631), .ZN(n15419) );
  AOI22_X1 U18995 ( .A1(n15873), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15889), .ZN(n15420) );
  AOI21_X1 U18996 ( .B1(n17172), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15421), .ZN(n15424) );
  NAND2_X1 U18997 ( .A1(n15422), .A2(n17190), .ZN(n15423) );
  OAI211_X1 U18998 ( .C1(n15429), .C2(n17166), .A(n15424), .B(n15423), .ZN(
        n15425) );
  AOI21_X1 U18999 ( .B1(n17196), .B2(n15426), .A(n15425), .ZN(n15427) );
  NAND2_X1 U19000 ( .A1(n20204), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n15431) );
  OAI21_X1 U19001 ( .B1(n15430), .B2(n20204), .A(n15431), .ZN(P2_U2856) );
  AOI22_X1 U19002 ( .A1(n20150), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n20169), 
        .B2(P2_EBX_REG_31__SCAN_IN), .ZN(n15433) );
  NAND2_X1 U19003 ( .A1(n20186), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15432) );
  OAI211_X1 U19004 ( .C1(n15434), .C2(n20165), .A(n15433), .B(n15432), .ZN(
        n15435) );
  AOI21_X1 U19005 ( .B1(n15437), .B2(n15436), .A(n15435), .ZN(n15439) );
  NAND2_X1 U19006 ( .A1(n16764), .A2(n20185), .ZN(n15438) );
  OAI211_X1 U19007 ( .C1(n15430), .C2(n20189), .A(n15439), .B(n15438), .ZN(
        P2_U2824) );
  INV_X1 U19008 ( .A(n20053), .ZN(n20961) );
  OAI21_X1 U19009 ( .B1(P2_READREQUEST_REG_SCAN_IN), .B2(n15440), .A(n20961), 
        .ZN(n15441) );
  OAI21_X1 U19010 ( .B1(n20961), .B2(n15442), .A(n15441), .ZN(P2_U3612) );
  OR2_X1 U19011 ( .A1(n15611), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n15445) );
  INV_X1 U19012 ( .A(n15443), .ZN(n15444) );
  MUX2_X1 U19013 ( .A(n15445), .B(n15444), .S(n21757), .Z(P1_U3487) );
  AOI21_X1 U19014 ( .B1(n15448), .B2(n15447), .A(n15446), .ZN(n15909) );
  INV_X1 U19015 ( .A(n15909), .ZN(n15828) );
  INV_X1 U19016 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21713) );
  INV_X1 U19017 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n15449) );
  OAI21_X1 U19018 ( .B1(n15471), .B2(n21713), .A(n15449), .ZN(n15458) );
  INV_X1 U19019 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n15450) );
  NOR2_X1 U19020 ( .A1(n21089), .A2(n15450), .ZN(n15456) );
  INV_X1 U19021 ( .A(n15451), .ZN(n15452) );
  OAI22_X1 U19022 ( .A1(n9697), .A2(n15907), .B1(n15454), .B2(n21068), .ZN(
        n15455) );
  AOI211_X1 U19023 ( .C1(n15458), .C2(n15457), .A(n15456), .B(n15455), .ZN(
        n15464) );
  OAI22_X1 U19024 ( .A1(n13112), .A2(n9701), .B1(n15459), .B2(n15460), .ZN(
        n15462) );
  XNOR2_X1 U19025 ( .A(n15462), .B(n15461), .ZN(n16134) );
  NAND2_X1 U19026 ( .A1(n16134), .A2(n21041), .ZN(n15463) );
  OAI211_X1 U19027 ( .C1(n15828), .C2(n15775), .A(n15464), .B(n15463), .ZN(
        P1_U2810) );
  XOR2_X1 U19028 ( .A(n15465), .B(n15479), .Z(n15914) );
  INV_X1 U19029 ( .A(n15914), .ZN(n15831) );
  NAND2_X1 U19030 ( .A1(n15459), .A2(n15466), .ZN(n15467) );
  NAND2_X1 U19031 ( .A1(n15468), .A2(n15467), .ZN(n15796) );
  INV_X1 U19032 ( .A(n15796), .ZN(n16142) );
  INV_X1 U19033 ( .A(n15469), .ZN(n15912) );
  OAI22_X1 U19034 ( .A1(n9697), .A2(n15912), .B1(n15470), .B2(n21068), .ZN(
        n15473) );
  NOR2_X1 U19035 ( .A1(n15471), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15472) );
  AOI211_X1 U19036 ( .C1(P1_EBX_REG_29__SCAN_IN), .C2(n21040), .A(n15473), .B(
        n15472), .ZN(n15474) );
  OAI21_X1 U19037 ( .B1(n21713), .B2(n15483), .A(n15474), .ZN(n15475) );
  AOI21_X1 U19038 ( .B1(n16142), .B2(n21041), .A(n15475), .ZN(n15476) );
  OAI21_X1 U19039 ( .B1(n15831), .B2(n15775), .A(n15476), .ZN(P1_U2811) );
  OAI21_X1 U19040 ( .B1(n15491), .B2(n15477), .A(n15459), .ZN(n16150) );
  AOI21_X1 U19041 ( .B1(n15480), .B2(n15478), .A(n15479), .ZN(n15925) );
  NAND2_X1 U19042 ( .A1(n15925), .A2(n21036), .ZN(n15488) );
  OAI22_X1 U19043 ( .A1(n9697), .A2(n15923), .B1(n15481), .B2(n21068), .ZN(
        n15486) );
  INV_X1 U19044 ( .A(n15482), .ZN(n15484) );
  INV_X1 U19045 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n15921) );
  AOI21_X1 U19046 ( .B1(n15484), .B2(n15921), .A(n15483), .ZN(n15485) );
  AOI211_X1 U19047 ( .C1(n21040), .C2(P1_EBX_REG_28__SCAN_IN), .A(n15486), .B(
        n15485), .ZN(n15487) );
  OAI211_X1 U19048 ( .C1(n21086), .C2(n16150), .A(n15488), .B(n15487), .ZN(
        P1_U2812) );
  OAI21_X1 U19049 ( .B1(n15489), .B2(n15490), .A(n15478), .ZN(n15932) );
  AOI21_X1 U19050 ( .B1(n15492), .B2(n15503), .A(n15491), .ZN(n16161) );
  INV_X1 U19051 ( .A(n21087), .ZN(n21081) );
  INV_X1 U19052 ( .A(n15507), .ZN(n15493) );
  INV_X1 U19053 ( .A(n21074), .ZN(n21080) );
  AOI21_X1 U19054 ( .B1(n21081), .B2(n15493), .A(n21080), .ZN(n15512) );
  INV_X1 U19055 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21708) );
  INV_X1 U19056 ( .A(n15931), .ZN(n15494) );
  OAI22_X1 U19057 ( .A1(n9697), .A2(n15494), .B1(n15929), .B2(n21068), .ZN(
        n15495) );
  AOI21_X1 U19058 ( .B1(n21040), .B2(P1_EBX_REG_27__SCAN_IN), .A(n15495), .ZN(
        n15497) );
  NAND3_X1 U19059 ( .A1(n21081), .A2(n15507), .A3(n21708), .ZN(n15496) );
  OAI211_X1 U19060 ( .C1(n15512), .C2(n21708), .A(n15497), .B(n15496), .ZN(
        n15498) );
  AOI21_X1 U19061 ( .B1(n16161), .B2(n21041), .A(n15498), .ZN(n15499) );
  OAI21_X1 U19062 ( .B1(n15932), .B2(n15775), .A(n15499), .ZN(P1_U2813) );
  AOI21_X1 U19063 ( .B1(n15501), .B2(n15500), .A(n15489), .ZN(n15944) );
  INV_X1 U19064 ( .A(n15944), .ZN(n15840) );
  INV_X1 U19065 ( .A(n15503), .ZN(n15504) );
  AOI21_X1 U19066 ( .B1(n15505), .B2(n15502), .A(n15504), .ZN(n16169) );
  NOR3_X1 U19067 ( .A1(n21087), .A2(n15507), .A3(n15506), .ZN(n15510) );
  OAI22_X1 U19068 ( .A1(n9697), .A2(n15942), .B1(n15508), .B2(n21068), .ZN(
        n15509) );
  AOI211_X1 U19069 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n21040), .A(n15510), .B(
        n15509), .ZN(n15511) );
  OAI21_X1 U19070 ( .B1(n15512), .B2(n21706), .A(n15511), .ZN(n15513) );
  AOI21_X1 U19071 ( .B1(n16169), .B2(n21041), .A(n15513), .ZN(n15514) );
  OAI21_X1 U19072 ( .B1(n15840), .B2(n15775), .A(n15514), .ZN(P1_U2814) );
  INV_X1 U19073 ( .A(n15500), .ZN(n15516) );
  AOI21_X1 U19074 ( .B1(n15517), .B2(n15515), .A(n15516), .ZN(n15954) );
  INV_X1 U19075 ( .A(n15954), .ZN(n15843) );
  OR2_X1 U19076 ( .A1(n15518), .A2(n15519), .ZN(n15520) );
  NAND2_X1 U19077 ( .A1(n15502), .A2(n15520), .ZN(n16175) );
  INV_X1 U19078 ( .A(n16175), .ZN(n15532) );
  INV_X1 U19079 ( .A(n15950), .ZN(n15521) );
  INV_X1 U19080 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15952) );
  OAI22_X1 U19081 ( .A1(n9697), .A2(n15521), .B1(n15952), .B2(n21068), .ZN(
        n15530) );
  INV_X1 U19082 ( .A(n15540), .ZN(n15522) );
  NAND2_X1 U19083 ( .A1(n21074), .A2(n15522), .ZN(n15523) );
  NAND2_X1 U19084 ( .A1(n15791), .A2(n15523), .ZN(n15556) );
  INV_X1 U19085 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21704) );
  NOR2_X1 U19086 ( .A1(n15556), .A2(n21704), .ZN(n15529) );
  NAND2_X1 U19087 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n15524) );
  OAI21_X1 U19088 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n15525), .A(n15524), 
        .ZN(n15526) );
  NOR2_X1 U19089 ( .A1(n21087), .A2(n15526), .ZN(n15528) );
  INV_X1 U19090 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15801) );
  NOR2_X1 U19091 ( .A1(n21089), .A2(n15801), .ZN(n15527) );
  OR4_X1 U19092 ( .A1(n15530), .A2(n15529), .A3(n15528), .A4(n15527), .ZN(
        n15531) );
  AOI21_X1 U19093 ( .B1(n15532), .B2(n21041), .A(n15531), .ZN(n15533) );
  OAI21_X1 U19094 ( .B1(n15843), .B2(n15775), .A(n15533), .ZN(P1_U2815) );
  OR2_X1 U19095 ( .A1(n15547), .A2(n15534), .ZN(n15535) );
  NAND2_X1 U19096 ( .A1(n15515), .A2(n15535), .ZN(n15962) );
  INV_X1 U19097 ( .A(n15536), .ZN(n15539) );
  INV_X1 U19098 ( .A(n15537), .ZN(n15538) );
  AOI21_X1 U19099 ( .B1(n15539), .B2(n15538), .A(n15518), .ZN(n16189) );
  NOR3_X1 U19100 ( .A1(n21087), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n15540), 
        .ZN(n15543) );
  INV_X1 U19101 ( .A(n15965), .ZN(n15541) );
  OAI22_X1 U19102 ( .A1(n21094), .A2(n15541), .B1(n15961), .B2(n21068), .ZN(
        n15542) );
  AOI211_X1 U19103 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n21040), .A(n15543), .B(
        n15542), .ZN(n15544) );
  OAI21_X1 U19104 ( .B1(n21702), .B2(n15556), .A(n15544), .ZN(n15545) );
  AOI21_X1 U19105 ( .B1(n16189), .B2(n21041), .A(n15545), .ZN(n15546) );
  OAI21_X1 U19106 ( .B1(n15962), .B2(n15775), .A(n15546), .ZN(P1_U2816) );
  AOI21_X1 U19107 ( .B1(n15548), .B2(n15568), .A(n15547), .ZN(n15973) );
  INV_X1 U19108 ( .A(n15973), .ZN(n15849) );
  AND2_X1 U19109 ( .A1(n15549), .A2(n15550), .ZN(n15551) );
  NOR2_X1 U19110 ( .A1(n15537), .A2(n15551), .ZN(n16197) );
  AOI21_X1 U19111 ( .B1(n21081), .B2(n15552), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n15557) );
  INV_X1 U19112 ( .A(n15969), .ZN(n15553) );
  INV_X1 U19113 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15971) );
  OAI22_X1 U19114 ( .A1(n21094), .A2(n15553), .B1(n15971), .B2(n21068), .ZN(
        n15554) );
  AOI21_X1 U19115 ( .B1(n21040), .B2(P1_EBX_REG_23__SCAN_IN), .A(n15554), .ZN(
        n15555) );
  OAI21_X1 U19116 ( .B1(n15557), .B2(n15556), .A(n15555), .ZN(n15558) );
  AOI21_X1 U19117 ( .B1(n16197), .B2(n21041), .A(n15558), .ZN(n15559) );
  OAI21_X1 U19118 ( .B1(n15849), .B2(n15775), .A(n15559), .ZN(P1_U2817) );
  INV_X1 U19119 ( .A(n16016), .ZN(n15560) );
  NAND2_X1 U19120 ( .A1(n15560), .A2(n15562), .ZN(n15561) );
  OAI21_X1 U19121 ( .B1(n15563), .B2(n15562), .A(n15561), .ZN(n15627) );
  NOR2_X4 U19122 ( .A1(n15641), .A2(n15627), .ZN(n15626) );
  INV_X1 U19123 ( .A(n15564), .ZN(n15596) );
  MUX2_X1 U19124 ( .A(n16008), .B(n15566), .S(n15565), .Z(n15608) );
  INV_X1 U19125 ( .A(n15584), .ZN(n15567) );
  INV_X1 U19126 ( .A(n15570), .ZN(n15585) );
  INV_X1 U19127 ( .A(n15571), .ZN(n15572) );
  OAI21_X1 U19128 ( .B1(n15585), .B2(n15572), .A(n15549), .ZN(n16208) );
  INV_X1 U19129 ( .A(n16208), .ZN(n15582) );
  NAND2_X1 U19130 ( .A1(n21074), .A2(n15590), .ZN(n15573) );
  NAND2_X1 U19131 ( .A1(n15791), .A2(n15573), .ZN(n15604) );
  OAI22_X1 U19132 ( .A1(n21094), .A2(n15981), .B1(n15574), .B2(n21068), .ZN(
        n15579) );
  INV_X1 U19133 ( .A(n15575), .ZN(n15576) );
  NOR2_X1 U19134 ( .A1(n15576), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15577) );
  AOI211_X1 U19135 ( .C1(P1_REIP_REG_21__SCAN_IN), .C2(P1_REIP_REG_22__SCAN_IN), .A(n15577), .B(n21087), .ZN(n15578) );
  AOI211_X1 U19136 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n21040), .A(n15579), .B(
        n15578), .ZN(n15580) );
  OAI21_X1 U19137 ( .B1(n21699), .B2(n15604), .A(n15580), .ZN(n15581) );
  AOI21_X1 U19138 ( .B1(n15582), .B2(n21041), .A(n15581), .ZN(n15583) );
  OAI21_X1 U19139 ( .B1(n15985), .B2(n15775), .A(n15583), .ZN(P1_U2818) );
  XNOR2_X1 U19140 ( .A(n15595), .B(n15584), .ZN(n15994) );
  INV_X1 U19141 ( .A(n15599), .ZN(n15586) );
  AOI21_X1 U19142 ( .B1(n15587), .B2(n15586), .A(n15585), .ZN(n16215) );
  INV_X1 U19143 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21697) );
  OAI22_X1 U19144 ( .A1(n9697), .A2(n15992), .B1(n15588), .B2(n21068), .ZN(
        n15589) );
  AOI21_X1 U19145 ( .B1(n21040), .B2(P1_EBX_REG_21__SCAN_IN), .A(n15589), .ZN(
        n15592) );
  NAND3_X1 U19146 ( .A1(n21081), .A2(n15590), .A3(n21697), .ZN(n15591) );
  OAI211_X1 U19147 ( .C1(n15604), .C2(n21697), .A(n15592), .B(n15591), .ZN(
        n15593) );
  AOI21_X1 U19148 ( .B1(n16215), .B2(n21041), .A(n15593), .ZN(n15594) );
  OAI21_X1 U19149 ( .B1(n15856), .B2(n15775), .A(n15594), .ZN(P1_U2819) );
  INV_X1 U19150 ( .A(n15595), .ZN(n15598) );
  AOI21_X1 U19151 ( .B1(n15626), .B2(n15608), .A(n15596), .ZN(n15597) );
  NOR2_X1 U19152 ( .A1(n15598), .A2(n15597), .ZN(n16003) );
  INV_X1 U19153 ( .A(n16003), .ZN(n15860) );
  AOI21_X1 U19154 ( .B1(n9861), .B2(n10533), .A(n15599), .ZN(n16227) );
  NAND2_X1 U19155 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n15600) );
  AOI21_X1 U19156 ( .B1(n15682), .B2(n15601), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15605) );
  AOI22_X1 U19157 ( .A1(n9698), .A2(n15999), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21082), .ZN(n15603) );
  NAND2_X1 U19158 ( .A1(n21040), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n15602) );
  OAI211_X1 U19159 ( .C1(n15605), .C2(n15604), .A(n15603), .B(n15602), .ZN(
        n15606) );
  AOI21_X1 U19160 ( .B1(n16227), .B2(n21041), .A(n15606), .ZN(n15607) );
  OAI21_X1 U19161 ( .B1(n15860), .B2(n15775), .A(n15607), .ZN(P1_U2820) );
  XOR2_X1 U19162 ( .A(n15608), .B(n15626), .Z(n16010) );
  AOI21_X1 U19163 ( .B1(n15610), .B2(n15628), .A(n15609), .ZN(n16235) );
  NAND2_X1 U19164 ( .A1(n21074), .A2(n15611), .ZN(n21042) );
  NAND2_X1 U19165 ( .A1(n21082), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15612) );
  OAI211_X1 U19166 ( .C1(n9697), .C2(n16008), .A(n21042), .B(n15612), .ZN(
        n15614) );
  INV_X1 U19167 ( .A(n15682), .ZN(n15615) );
  INV_X1 U19168 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n16014) );
  NOR4_X1 U19169 ( .A1(n15615), .A2(P1_REIP_REG_19__SCAN_IN), .A3(n15620), 
        .A4(n16014), .ZN(n15613) );
  AOI211_X1 U19170 ( .C1(P1_EBX_REG_19__SCAN_IN), .C2(n21040), .A(n15614), .B(
        n15613), .ZN(n15623) );
  NOR3_X1 U19171 ( .A1(n15615), .A2(P1_REIP_REG_18__SCAN_IN), .A3(n15620), 
        .ZN(n15637) );
  INV_X1 U19172 ( .A(n15616), .ZN(n15617) );
  AND2_X1 U19173 ( .A1(n21074), .A2(n15617), .ZN(n15749) );
  NAND2_X1 U19174 ( .A1(n15749), .A2(n15618), .ZN(n15619) );
  NAND2_X1 U19175 ( .A1(n15791), .A2(n15619), .ZN(n15691) );
  NAND2_X1 U19176 ( .A1(n15791), .A2(n15620), .ZN(n15621) );
  NAND2_X1 U19177 ( .A1(n15691), .A2(n15621), .ZN(n15632) );
  OAI21_X1 U19178 ( .B1(n15637), .B2(n15632), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15622) );
  NAND2_X1 U19179 ( .A1(n15623), .A2(n15622), .ZN(n15624) );
  AOI21_X1 U19180 ( .B1(n16235), .B2(n21041), .A(n15624), .ZN(n15625) );
  OAI21_X1 U19181 ( .B1(n15864), .B2(n15775), .A(n15625), .ZN(P1_U2821) );
  AOI21_X1 U19182 ( .B1(n15627), .B2(n15641), .A(n15626), .ZN(n16018) );
  INV_X1 U19183 ( .A(n16018), .ZN(n15868) );
  INV_X1 U19184 ( .A(n15628), .ZN(n15629) );
  AOI21_X1 U19185 ( .B1(n15630), .B2(n15650), .A(n15629), .ZN(n16248) );
  NAND2_X1 U19186 ( .A1(n21082), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15631) );
  OAI211_X1 U19187 ( .C1(n21094), .C2(n16016), .A(n21042), .B(n15631), .ZN(
        n15634) );
  INV_X1 U19188 ( .A(n15632), .ZN(n15643) );
  NOR2_X1 U19189 ( .A1(n15643), .A2(n16014), .ZN(n15633) );
  INV_X1 U19190 ( .A(n15635), .ZN(n15636) );
  OAI21_X1 U19191 ( .B1(n15868), .B2(n15775), .A(n15638), .ZN(P1_U2822) );
  NAND2_X1 U19192 ( .A1(n15658), .A2(n15639), .ZN(n15640) );
  NAND2_X1 U19193 ( .A1(n15641), .A2(n15640), .ZN(n16026) );
  NAND2_X1 U19194 ( .A1(n21082), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15642) );
  OAI211_X1 U19195 ( .C1(n9697), .C2(n16028), .A(n21042), .B(n15642), .ZN(
        n15646) );
  NAND3_X1 U19196 ( .A1(n15682), .A2(P1_REIP_REG_16__SCAN_IN), .A3(
        P1_REIP_REG_15__SCAN_IN), .ZN(n15644) );
  INV_X1 U19197 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21690) );
  AOI21_X1 U19198 ( .B1(n15644), .B2(n21690), .A(n15643), .ZN(n15645) );
  AOI211_X1 U19199 ( .C1(P1_EBX_REG_17__SCAN_IN), .C2(n21040), .A(n15646), .B(
        n15645), .ZN(n15652) );
  NAND2_X1 U19200 ( .A1(n15647), .A2(n15648), .ZN(n15649) );
  AND2_X1 U19201 ( .A1(n15650), .A2(n15649), .ZN(n16256) );
  NAND2_X1 U19202 ( .A1(n16256), .A2(n21041), .ZN(n15651) );
  OAI211_X1 U19203 ( .C1(n16026), .C2(n15775), .A(n15652), .B(n15651), .ZN(
        P1_U2823) );
  OR2_X1 U19204 ( .A1(n15653), .A2(n15654), .ZN(n15655) );
  NAND2_X1 U19205 ( .A1(n15647), .A2(n15655), .ZN(n16265) );
  INV_X1 U19206 ( .A(n15658), .ZN(n15659) );
  AOI21_X1 U19207 ( .B1(n15660), .B2(n15674), .A(n15659), .ZN(n16041) );
  NAND2_X1 U19208 ( .A1(n16041), .A2(n21036), .ZN(n15667) );
  INV_X1 U19209 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n15681) );
  XNOR2_X1 U19210 ( .A(n15681), .B(P1_REIP_REG_16__SCAN_IN), .ZN(n15665) );
  INV_X1 U19211 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21688) );
  NAND2_X1 U19212 ( .A1(n21082), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15661) );
  OAI211_X1 U19213 ( .C1(n9697), .C2(n16039), .A(n21042), .B(n15661), .ZN(
        n15662) );
  AOI21_X1 U19214 ( .B1(n21040), .B2(P1_EBX_REG_16__SCAN_IN), .A(n15662), .ZN(
        n15663) );
  OAI21_X1 U19215 ( .B1(n21688), .B2(n15691), .A(n15663), .ZN(n15664) );
  AOI21_X1 U19216 ( .B1(n15682), .B2(n15665), .A(n15664), .ZN(n15666) );
  OAI211_X1 U19217 ( .C1(n16265), .C2(n21086), .A(n15667), .B(n15666), .ZN(
        P1_U2824) );
  AND2_X1 U19218 ( .A1(n15668), .A2(n15669), .ZN(n15670) );
  OR2_X1 U19219 ( .A1(n15653), .A2(n15670), .ZN(n16273) );
  NAND2_X1 U19220 ( .A1(n9747), .A2(n15729), .ZN(n15672) );
  AOI21_X2 U19221 ( .B1(n15699), .B2(n15672), .A(n15671), .ZN(n15702) );
  NAND2_X1 U19222 ( .A1(n15702), .A2(n15686), .ZN(n15685) );
  INV_X1 U19223 ( .A(n15673), .ZN(n15676) );
  INV_X1 U19224 ( .A(n15674), .ZN(n15675) );
  AOI21_X2 U19225 ( .B1(n15685), .B2(n15676), .A(n15675), .ZN(n16052) );
  NAND2_X1 U19226 ( .A1(n16052), .A2(n21036), .ZN(n15684) );
  NAND2_X1 U19227 ( .A1(n21082), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15677) );
  OAI211_X1 U19228 ( .C1(n9697), .C2(n16050), .A(n21042), .B(n15677), .ZN(
        n15678) );
  AOI21_X1 U19229 ( .B1(n21040), .B2(P1_EBX_REG_15__SCAN_IN), .A(n15678), .ZN(
        n15679) );
  OAI21_X1 U19230 ( .B1(n15681), .B2(n15691), .A(n15679), .ZN(n15680) );
  AOI21_X1 U19231 ( .B1(n15682), .B2(n15681), .A(n15680), .ZN(n15683) );
  OAI211_X1 U19232 ( .C1(n16273), .C2(n21086), .A(n15684), .B(n15683), .ZN(
        P1_U2825) );
  OAI21_X1 U19233 ( .B1(n15702), .B2(n15686), .A(n15685), .ZN(n16064) );
  INV_X1 U19234 ( .A(n15668), .ZN(n15687) );
  AOI21_X1 U19235 ( .B1(n15688), .B2(n15708), .A(n15687), .ZN(n16284) );
  INV_X1 U19236 ( .A(n15689), .ZN(n15690) );
  AOI21_X1 U19237 ( .B1(n15724), .B2(n15690), .A(P1_REIP_REG_14__SCAN_IN), 
        .ZN(n15692) );
  NOR2_X1 U19238 ( .A1(n15692), .A2(n15691), .ZN(n15696) );
  INV_X1 U19239 ( .A(n21042), .ZN(n21060) );
  AOI21_X1 U19240 ( .B1(n21082), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n21060), .ZN(n15694) );
  NAND2_X1 U19241 ( .A1(n21040), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n15693) );
  OAI211_X1 U19242 ( .C1(n9697), .C2(n16060), .A(n15694), .B(n15693), .ZN(
        n15695) );
  AOI211_X1 U19243 ( .C1(n16284), .C2(n21041), .A(n15696), .B(n15695), .ZN(
        n15697) );
  OAI21_X1 U19244 ( .B1(n16064), .B2(n15775), .A(n15697), .ZN(P1_U2826) );
  OAI21_X1 U19245 ( .B1(n9747), .B2(n15698), .A(n15699), .ZN(n15730) );
  INV_X1 U19246 ( .A(n15729), .ZN(n15700) );
  OAI21_X1 U19247 ( .B1(n15730), .B2(n15700), .A(n15699), .ZN(n15717) );
  NAND2_X1 U19248 ( .A1(n15717), .A2(n15716), .ZN(n15715) );
  INV_X1 U19249 ( .A(n15701), .ZN(n15703) );
  AOI21_X1 U19250 ( .B1(n15715), .B2(n15703), .A(n15702), .ZN(n16079) );
  INV_X1 U19251 ( .A(n16079), .ZN(n15884) );
  NAND2_X1 U19252 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n15711) );
  INV_X1 U19253 ( .A(n15711), .ZN(n15704) );
  INV_X1 U19254 ( .A(n15791), .ZN(n15734) );
  AOI21_X1 U19255 ( .B1(n15749), .B2(n15704), .A(n15734), .ZN(n15725) );
  AOI21_X1 U19256 ( .B1(n21082), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n21060), .ZN(n15706) );
  NAND2_X1 U19257 ( .A1(n21040), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n15705) );
  OAI211_X1 U19258 ( .C1(n9697), .C2(n16077), .A(n15706), .B(n15705), .ZN(
        n15707) );
  AOI21_X1 U19259 ( .B1(n15725), .B2(P1_REIP_REG_13__SCAN_IN), .A(n15707), 
        .ZN(n15714) );
  INV_X1 U19260 ( .A(n15721), .ZN(n15709) );
  AOI21_X1 U19261 ( .B1(n15710), .B2(n15709), .A(n13054), .ZN(n16290) );
  NOR2_X1 U19262 ( .A1(n15711), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15712) );
  AOI22_X1 U19263 ( .A1(n16290), .A2(n21041), .B1(n15724), .B2(n15712), .ZN(
        n15713) );
  OAI211_X1 U19264 ( .C1(n15884), .C2(n15775), .A(n15714), .B(n15713), .ZN(
        P1_U2827) );
  NAND2_X1 U19265 ( .A1(n21082), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15718) );
  OAI211_X1 U19266 ( .C1(n9697), .C2(n16086), .A(n21042), .B(n15718), .ZN(
        n15723) );
  NOR2_X1 U19267 ( .A1(n9826), .A2(n15719), .ZN(n15720) );
  OR2_X1 U19268 ( .A1(n15721), .A2(n15720), .ZN(n16303) );
  NOR2_X1 U19269 ( .A1(n16303), .A2(n21086), .ZN(n15722) );
  AOI211_X1 U19270 ( .C1(P1_EBX_REG_12__SCAN_IN), .C2(n21040), .A(n15723), .B(
        n15722), .ZN(n15728) );
  INV_X1 U19271 ( .A(n15724), .ZN(n15739) );
  INV_X1 U19272 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21680) );
  NOR2_X1 U19273 ( .A1(n15739), .A2(n21680), .ZN(n15726) );
  OAI21_X1 U19274 ( .B1(n15726), .B2(P1_REIP_REG_12__SCAN_IN), .A(n15725), 
        .ZN(n15727) );
  OAI211_X1 U19275 ( .C1(n16085), .C2(n15775), .A(n15728), .B(n15727), .ZN(
        P1_U2828) );
  XNOR2_X1 U19276 ( .A(n15730), .B(n15729), .ZN(n16100) );
  NAND2_X1 U19277 ( .A1(n16100), .A2(n21036), .ZN(n15738) );
  INV_X1 U19278 ( .A(n16343), .ZN(n15744) );
  AOI21_X1 U19279 ( .B1(n15744), .B2(n15743), .A(n10543), .ZN(n15731) );
  NOR2_X1 U19280 ( .A1(n15731), .A2(n9826), .ZN(n16315) );
  AOI21_X1 U19281 ( .B1(n21082), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n21060), .ZN(n15733) );
  NAND2_X1 U19282 ( .A1(n21040), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n15732) );
  OAI211_X1 U19283 ( .C1(n9697), .C2(n16098), .A(n15733), .B(n15732), .ZN(
        n15736) );
  NOR3_X1 U19284 ( .A1(n15734), .A2(n15749), .A3(n21680), .ZN(n15735) );
  AOI211_X1 U19285 ( .C1(n16315), .C2(n21041), .A(n15736), .B(n15735), .ZN(
        n15737) );
  OAI211_X1 U19286 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n15739), .A(n15738), 
        .B(n15737), .ZN(P1_U2829) );
  INV_X1 U19287 ( .A(n15740), .ZN(n15742) );
  AOI21_X1 U19288 ( .B1(n15742), .B2(n15741), .A(n9747), .ZN(n16113) );
  INV_X1 U19289 ( .A(n16113), .ZN(n15892) );
  XNOR2_X1 U19290 ( .A(n15744), .B(n15743), .ZN(n16323) );
  INV_X1 U19291 ( .A(n16323), .ZN(n15819) );
  NAND2_X1 U19292 ( .A1(n21082), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15745) );
  OAI211_X1 U19293 ( .C1(n9697), .C2(n16111), .A(n21042), .B(n15745), .ZN(
        n15746) );
  INV_X1 U19294 ( .A(n15746), .ZN(n15755) );
  INV_X1 U19295 ( .A(n15747), .ZN(n21010) );
  INV_X1 U19296 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21677) );
  NOR2_X1 U19297 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n21677), .ZN(n15748) );
  NAND2_X1 U19298 ( .A1(n21010), .A2(n15748), .ZN(n15754) );
  INV_X1 U19299 ( .A(n15749), .ZN(n15750) );
  NAND3_X1 U19300 ( .A1(n15791), .A2(P1_REIP_REG_10__SCAN_IN), .A3(n15750), 
        .ZN(n15753) );
  OR2_X1 U19301 ( .A1(n21089), .A2(n15751), .ZN(n15752) );
  NAND4_X1 U19302 ( .A1(n15755), .A2(n15754), .A3(n15753), .A4(n15752), .ZN(
        n15756) );
  AOI21_X1 U19303 ( .B1(n21041), .B2(n15819), .A(n15756), .ZN(n15757) );
  OAI21_X1 U19304 ( .B1(n15892), .B2(n15775), .A(n15757), .ZN(P1_U2830) );
  AOI21_X1 U19305 ( .B1(n15760), .B2(n15759), .A(n15758), .ZN(n16126) );
  INV_X1 U19306 ( .A(n16126), .ZN(n15902) );
  OR2_X1 U19307 ( .A1(n14762), .A2(n15762), .ZN(n15763) );
  NAND2_X1 U19308 ( .A1(n15761), .A2(n15763), .ZN(n17893) );
  OAI21_X1 U19309 ( .B1(n15764), .B2(n21087), .A(n21074), .ZN(n21009) );
  AOI22_X1 U19310 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n21082), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n21009), .ZN(n15765) );
  OAI211_X1 U19311 ( .C1(n21086), .C2(n17893), .A(n15765), .B(n21042), .ZN(
        n15770) );
  NOR3_X1 U19312 ( .A1(n21087), .A2(n15766), .A3(P1_REIP_REG_8__SCAN_IN), .ZN(
        n15769) );
  OAI22_X1 U19313 ( .A1(n9697), .A2(n16124), .B1(n15767), .B2(n21089), .ZN(
        n15768) );
  NOR3_X1 U19314 ( .A1(n15770), .A2(n15769), .A3(n15768), .ZN(n15771) );
  OAI21_X1 U19315 ( .B1(n15902), .B2(n15775), .A(n15771), .ZN(P1_U2832) );
  INV_X1 U19316 ( .A(n15777), .ZN(n15773) );
  NAND2_X1 U19317 ( .A1(n15773), .A2(n15772), .ZN(n15774) );
  NAND2_X1 U19318 ( .A1(n15775), .A2(n15774), .ZN(n21096) );
  INV_X1 U19319 ( .A(n21096), .ZN(n15794) );
  AOI22_X1 U19320 ( .A1(n21081), .A2(n21660), .B1(n21040), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n15784) );
  NOR2_X1 U19321 ( .A1(n15777), .A2(n15776), .ZN(n21083) );
  OAI22_X1 U19322 ( .A1(n21068), .A2(n15778), .B1(n21660), .B2(n21074), .ZN(
        n15779) );
  AOI21_X1 U19323 ( .B1(n21526), .B2(n21083), .A(n15779), .ZN(n15780) );
  OAI21_X1 U19324 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n9697), .A(
        n15780), .ZN(n15781) );
  AOI21_X1 U19325 ( .B1(n21041), .B2(n15782), .A(n15781), .ZN(n15783) );
  OAI211_X1 U19326 ( .C1(n15785), .C2(n15794), .A(n15784), .B(n15783), .ZN(
        P1_U2839) );
  INV_X1 U19327 ( .A(n21083), .ZN(n21054) );
  OAI21_X1 U19328 ( .B1(n9698), .B2(n21082), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15788) );
  AOI22_X1 U19329 ( .A1(n21041), .A2(n15786), .B1(n21040), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n15787) );
  OAI211_X1 U19330 ( .C1(n21054), .C2(n15789), .A(n15788), .B(n15787), .ZN(
        n15790) );
  AOI21_X1 U19331 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(n15791), .A(n15790), .ZN(
        n15792) );
  OAI21_X1 U19332 ( .B1(n15794), .B2(n15793), .A(n15792), .ZN(P1_U2840) );
  AOI22_X1 U19333 ( .A1(n16134), .A2(n21111), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n15818), .ZN(n15795) );
  OAI21_X1 U19334 ( .B1(n15828), .B2(n15817), .A(n15795), .ZN(P1_U2842) );
  OAI222_X1 U19335 ( .A1(n15797), .A2(n21116), .B1(n15821), .B2(n15796), .C1(
        n15817), .C2(n15831), .ZN(P1_U2843) );
  INV_X1 U19336 ( .A(n15925), .ZN(n15834) );
  OAI222_X1 U19337 ( .A1(n15798), .A2(n21116), .B1(n15821), .B2(n16150), .C1(
        n15834), .C2(n15817), .ZN(P1_U2844) );
  AOI22_X1 U19338 ( .A1(n16161), .A2(n21111), .B1(n15818), .B2(
        P1_EBX_REG_27__SCAN_IN), .ZN(n15799) );
  OAI21_X1 U19339 ( .B1(n15932), .B2(n15817), .A(n15799), .ZN(P1_U2845) );
  AOI22_X1 U19340 ( .A1(n16169), .A2(n21111), .B1(n15818), .B2(
        P1_EBX_REG_26__SCAN_IN), .ZN(n15800) );
  OAI21_X1 U19341 ( .B1(n15840), .B2(n15817), .A(n15800), .ZN(P1_U2846) );
  OAI222_X1 U19342 ( .A1(n15801), .A2(n21116), .B1(n15821), .B2(n16175), .C1(
        n15843), .C2(n15817), .ZN(P1_U2847) );
  AOI22_X1 U19343 ( .A1(n16189), .A2(n21111), .B1(n15818), .B2(
        P1_EBX_REG_24__SCAN_IN), .ZN(n15802) );
  OAI21_X1 U19344 ( .B1(n15962), .B2(n15817), .A(n15802), .ZN(P1_U2848) );
  INV_X1 U19345 ( .A(n16197), .ZN(n15804) );
  OAI222_X1 U19346 ( .A1(n15804), .A2(n15821), .B1(n15803), .B2(n21116), .C1(
        n15849), .C2(n15817), .ZN(P1_U2849) );
  AOI22_X1 U19347 ( .A1(n16215), .A2(n21111), .B1(n15818), .B2(
        P1_EBX_REG_21__SCAN_IN), .ZN(n15806) );
  OAI21_X1 U19348 ( .B1(n15856), .B2(n15817), .A(n15806), .ZN(P1_U2851) );
  AOI22_X1 U19349 ( .A1(n16227), .A2(n21111), .B1(n15818), .B2(
        P1_EBX_REG_20__SCAN_IN), .ZN(n15807) );
  OAI21_X1 U19350 ( .B1(n15860), .B2(n15817), .A(n15807), .ZN(P1_U2852) );
  AOI22_X1 U19351 ( .A1(n16235), .A2(n21111), .B1(n15818), .B2(
        P1_EBX_REG_19__SCAN_IN), .ZN(n15808) );
  OAI21_X1 U19352 ( .B1(n15864), .B2(n15817), .A(n15808), .ZN(P1_U2853) );
  AOI22_X1 U19353 ( .A1(n16248), .A2(n21111), .B1(n15818), .B2(
        P1_EBX_REG_18__SCAN_IN), .ZN(n15809) );
  OAI21_X1 U19354 ( .B1(n15868), .B2(n15817), .A(n15809), .ZN(P1_U2854) );
  AOI22_X1 U19355 ( .A1(n16256), .A2(n21111), .B1(n15818), .B2(
        P1_EBX_REG_17__SCAN_IN), .ZN(n15810) );
  OAI21_X1 U19356 ( .B1(n16026), .B2(n15817), .A(n15810), .ZN(P1_U2855) );
  INV_X1 U19357 ( .A(n16041), .ZN(n15878) );
  OAI222_X1 U19358 ( .A1(n16265), .A2(n15821), .B1(n15811), .B2(n21116), .C1(
        n15878), .C2(n15817), .ZN(P1_U2856) );
  INV_X1 U19359 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15812) );
  INV_X1 U19360 ( .A(n16052), .ZN(n15880) );
  OAI222_X1 U19361 ( .A1(n16273), .A2(n15821), .B1(n15812), .B2(n21116), .C1(
        n15880), .C2(n15817), .ZN(P1_U2857) );
  AOI22_X1 U19362 ( .A1(n16284), .A2(n21111), .B1(n15818), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n15813) );
  OAI21_X1 U19363 ( .B1(n16064), .B2(n15817), .A(n15813), .ZN(P1_U2858) );
  AOI22_X1 U19364 ( .A1(n16290), .A2(n21111), .B1(n15818), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n15814) );
  OAI21_X1 U19365 ( .B1(n15884), .B2(n15817), .A(n15814), .ZN(P1_U2859) );
  OAI222_X1 U19366 ( .A1(n16303), .A2(n15821), .B1(n15815), .B2(n21116), .C1(
        n16085), .C2(n15817), .ZN(P1_U2860) );
  INV_X1 U19367 ( .A(n16100), .ZN(n15888) );
  AOI22_X1 U19368 ( .A1(n16315), .A2(n21111), .B1(n15818), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15816) );
  OAI21_X1 U19369 ( .B1(n15888), .B2(n15817), .A(n15816), .ZN(P1_U2861) );
  AOI22_X1 U19370 ( .A1(n15819), .A2(n21111), .B1(n15818), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n15820) );
  OAI21_X1 U19371 ( .B1(n15892), .B2(n15817), .A(n15820), .ZN(P1_U2862) );
  OAI222_X1 U19372 ( .A1(n17893), .A2(n15821), .B1(n21116), .B2(n15767), .C1(
        n15817), .C2(n15902), .ZN(P1_U2864) );
  AOI22_X1 U19373 ( .A1(n15872), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n15889), .ZN(n15827) );
  NOR3_X1 U19374 ( .A1(n15889), .A2(n15824), .A3(n15823), .ZN(n15825) );
  AOI22_X1 U19375 ( .A1(n15875), .A2(n15881), .B1(n15873), .B2(DATAI_30_), 
        .ZN(n15826) );
  OAI211_X1 U19376 ( .C1(n15828), .C2(n15897), .A(n15827), .B(n15826), .ZN(
        P1_U2874) );
  AOI22_X1 U19377 ( .A1(n15872), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n15889), .ZN(n15830) );
  MUX2_X1 U19378 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n15837), .Z(
        n21160) );
  AOI22_X1 U19379 ( .A1(n15875), .A2(n21160), .B1(n15873), .B2(DATAI_29_), 
        .ZN(n15829) );
  OAI211_X1 U19380 ( .C1(n15831), .C2(n15897), .A(n15830), .B(n15829), .ZN(
        P1_U2875) );
  AOI22_X1 U19381 ( .A1(n15872), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n15889), .ZN(n15833) );
  MUX2_X1 U19382 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n15837), .Z(
        n21158) );
  AOI22_X1 U19383 ( .A1(n15875), .A2(n21158), .B1(n15873), .B2(DATAI_28_), 
        .ZN(n15832) );
  OAI211_X1 U19384 ( .C1(n15834), .C2(n15897), .A(n15833), .B(n15832), .ZN(
        P1_U2876) );
  AOI22_X1 U19385 ( .A1(n15872), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n15889), .ZN(n15836) );
  MUX2_X1 U19386 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n15837), .Z(
        n21156) );
  AOI22_X1 U19387 ( .A1(n15875), .A2(n21156), .B1(n15873), .B2(DATAI_27_), 
        .ZN(n15835) );
  OAI211_X1 U19388 ( .C1(n15932), .C2(n15897), .A(n15836), .B(n15835), .ZN(
        P1_U2877) );
  AOI22_X1 U19389 ( .A1(n15872), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n15889), .ZN(n15839) );
  MUX2_X1 U19390 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n15837), .Z(
        n21153) );
  AOI22_X1 U19391 ( .A1(n15875), .A2(n21153), .B1(n15873), .B2(DATAI_26_), 
        .ZN(n15838) );
  OAI211_X1 U19392 ( .C1(n15840), .C2(n15897), .A(n15839), .B(n15838), .ZN(
        P1_U2878) );
  AOI22_X1 U19393 ( .A1(n15872), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n15889), .ZN(n15842) );
  AOI22_X1 U19394 ( .A1(n15875), .A2(n15895), .B1(n15873), .B2(DATAI_25_), 
        .ZN(n15841) );
  OAI211_X1 U19395 ( .C1(n15843), .C2(n15897), .A(n15842), .B(n15841), .ZN(
        P1_U2879) );
  AOI22_X1 U19396 ( .A1(n15872), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n15889), .ZN(n15845) );
  AOI22_X1 U19397 ( .A1(n15875), .A2(n15898), .B1(n15873), .B2(DATAI_24_), 
        .ZN(n15844) );
  OAI211_X1 U19398 ( .C1(n15962), .C2(n15897), .A(n15845), .B(n15844), .ZN(
        P1_U2880) );
  AOI22_X1 U19399 ( .A1(n15872), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n15889), .ZN(n15848) );
  AOI22_X1 U19400 ( .A1(n15875), .A2(n15846), .B1(n15873), .B2(DATAI_23_), 
        .ZN(n15847) );
  OAI211_X1 U19401 ( .C1(n15849), .C2(n15897), .A(n15848), .B(n15847), .ZN(
        P1_U2881) );
  AOI22_X1 U19402 ( .A1(n15872), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n15889), .ZN(n15852) );
  AOI22_X1 U19403 ( .A1(n15875), .A2(n15850), .B1(n15873), .B2(DATAI_22_), 
        .ZN(n15851) );
  OAI211_X1 U19404 ( .C1(n15985), .C2(n15897), .A(n15852), .B(n15851), .ZN(
        P1_U2882) );
  AOI22_X1 U19405 ( .A1(n15872), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n15889), .ZN(n15855) );
  AOI22_X1 U19406 ( .A1(n15875), .A2(n15853), .B1(n15873), .B2(DATAI_21_), 
        .ZN(n15854) );
  OAI211_X1 U19407 ( .C1(n15856), .C2(n15897), .A(n15855), .B(n15854), .ZN(
        P1_U2883) );
  AOI22_X1 U19408 ( .A1(n15872), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n15889), .ZN(n15859) );
  AOI22_X1 U19409 ( .A1(n15875), .A2(n15857), .B1(n15873), .B2(DATAI_20_), 
        .ZN(n15858) );
  OAI211_X1 U19410 ( .C1(n15860), .C2(n15897), .A(n15859), .B(n15858), .ZN(
        P1_U2884) );
  AOI22_X1 U19411 ( .A1(n15872), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n15889), .ZN(n15863) );
  AOI22_X1 U19412 ( .A1(n15875), .A2(n15861), .B1(n15873), .B2(DATAI_19_), 
        .ZN(n15862) );
  OAI211_X1 U19413 ( .C1(n15864), .C2(n15897), .A(n15863), .B(n15862), .ZN(
        P1_U2885) );
  AOI22_X1 U19414 ( .A1(n15872), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n15889), .ZN(n15867) );
  AOI22_X1 U19415 ( .A1(n15875), .A2(n15865), .B1(n15873), .B2(DATAI_18_), 
        .ZN(n15866) );
  OAI211_X1 U19416 ( .C1(n15868), .C2(n15897), .A(n15867), .B(n15866), .ZN(
        P1_U2886) );
  AOI22_X1 U19417 ( .A1(n15872), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n15889), .ZN(n15871) );
  AOI22_X1 U19418 ( .A1(n15875), .A2(n15869), .B1(n15873), .B2(DATAI_17_), 
        .ZN(n15870) );
  OAI211_X1 U19419 ( .C1(n16026), .C2(n15897), .A(n15871), .B(n15870), .ZN(
        P1_U2887) );
  AOI22_X1 U19420 ( .A1(n15872), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n15889), .ZN(n15877) );
  AOI22_X1 U19421 ( .A1(n15875), .A2(n15874), .B1(n15873), .B2(DATAI_16_), 
        .ZN(n15876) );
  OAI211_X1 U19422 ( .C1(n15878), .C2(n15897), .A(n15877), .B(n15876), .ZN(
        P1_U2888) );
  OAI222_X1 U19423 ( .A1(n15880), .A2(n15897), .B1(n15901), .B2(n15879), .C1(
        n21124), .C2(n15899), .ZN(P1_U2889) );
  INV_X1 U19424 ( .A(n15881), .ZN(n15882) );
  OAI222_X1 U19425 ( .A1(n16064), .A2(n15897), .B1(n15901), .B2(n15882), .C1(
        n21126), .C2(n15899), .ZN(P1_U2890) );
  AOI22_X1 U19426 ( .A1(n15890), .A2(n21160), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15889), .ZN(n15883) );
  OAI21_X1 U19427 ( .B1(n15884), .B2(n15897), .A(n15883), .ZN(P1_U2891) );
  AOI22_X1 U19428 ( .A1(n15890), .A2(n21158), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n15889), .ZN(n15885) );
  OAI21_X1 U19429 ( .B1(n16085), .B2(n15897), .A(n15885), .ZN(P1_U2892) );
  INV_X1 U19430 ( .A(n21156), .ZN(n15887) );
  OAI222_X1 U19431 ( .A1(n15888), .A2(n15897), .B1(n15901), .B2(n15887), .C1(
        n15886), .C2(n15899), .ZN(P1_U2893) );
  AOI22_X1 U19432 ( .A1(n15890), .A2(n21153), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15889), .ZN(n15891) );
  OAI21_X1 U19433 ( .B1(n15892), .B2(n15897), .A(n15891), .ZN(P1_U2894) );
  INV_X1 U19434 ( .A(n15895), .ZN(n15896) );
  OAI222_X1 U19435 ( .A1(n21011), .A2(n15897), .B1(n15901), .B2(n15896), .C1(
        n15899), .C2(n14956), .ZN(P1_U2895) );
  INV_X1 U19436 ( .A(n15898), .ZN(n15900) );
  OAI222_X1 U19437 ( .A1(n15902), .A2(n15897), .B1(n15901), .B2(n15900), .C1(
        n15899), .C2(n14927), .ZN(P1_U2896) );
  NAND2_X1 U19438 ( .A1(n15904), .A2(n15903), .ZN(n15905) );
  XNOR2_X1 U19439 ( .A(n15905), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16136) );
  NAND2_X1 U19440 ( .A1(n17906), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n16129) );
  NAND2_X1 U19441 ( .A1(n17870), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15906) );
  OAI211_X1 U19442 ( .C1(n15907), .C2(n17877), .A(n16129), .B(n15906), .ZN(
        n15908) );
  AOI21_X1 U19443 ( .B1(n15909), .B2(n17882), .A(n15908), .ZN(n15910) );
  OAI21_X1 U19444 ( .B1(n16136), .B2(n20989), .A(n15910), .ZN(P1_U2969) );
  NOR2_X1 U19445 ( .A1(n17899), .A2(n21713), .ZN(n16140) );
  AOI21_X1 U19446 ( .B1(n17870), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16140), .ZN(n15911) );
  OAI21_X1 U19447 ( .B1(n15912), .B2(n17877), .A(n15911), .ZN(n15913) );
  AOI21_X1 U19448 ( .B1(n15914), .B2(n17882), .A(n15913), .ZN(n15915) );
  OAI21_X1 U19449 ( .B1(n16145), .B2(n20989), .A(n15915), .ZN(P1_U2970) );
  NAND2_X1 U19450 ( .A1(n15916), .A2(n15939), .ZN(n16164) );
  NOR4_X1 U19451 ( .A1(n16164), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15917) );
  NAND2_X1 U19452 ( .A1(n16103), .A2(n15917), .ZN(n15919) );
  NOR2_X1 U19453 ( .A1(n17899), .A2(n15921), .ZN(n16148) );
  AOI21_X1 U19454 ( .B1(n17870), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16148), .ZN(n15922) );
  OAI21_X1 U19455 ( .B1(n15923), .B2(n17877), .A(n15922), .ZN(n15924) );
  AOI21_X1 U19456 ( .B1(n15925), .B2(n17882), .A(n15924), .ZN(n15926) );
  OAI21_X1 U19457 ( .B1(n16154), .B2(n20989), .A(n15926), .ZN(P1_U2971) );
  NOR2_X1 U19458 ( .A1(n17899), .A2(n21708), .ZN(n16155) );
  NOR2_X1 U19459 ( .A1(n17885), .A2(n15929), .ZN(n15930) );
  AOI211_X1 U19460 ( .C1(n17880), .C2(n15931), .A(n16155), .B(n15930), .ZN(
        n15935) );
  INV_X1 U19461 ( .A(n15932), .ZN(n15933) );
  NAND2_X1 U19462 ( .A1(n15933), .A2(n17882), .ZN(n15934) );
  OAI211_X1 U19463 ( .C1(n16163), .C2(n20989), .A(n15935), .B(n15934), .ZN(
        P1_U2972) );
  OAI21_X1 U19464 ( .B1(n15956), .B2(n15936), .A(n9689), .ZN(n15937) );
  NAND2_X1 U19465 ( .A1(n15938), .A2(n15937), .ZN(n15940) );
  XNOR2_X1 U19466 ( .A(n15940), .B(n15939), .ZN(n16172) );
  NOR2_X1 U19467 ( .A1(n17899), .A2(n21706), .ZN(n16168) );
  AOI21_X1 U19468 ( .B1(n17870), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16168), .ZN(n15941) );
  OAI21_X1 U19469 ( .B1(n15942), .B2(n17877), .A(n15941), .ZN(n15943) );
  AOI21_X1 U19470 ( .B1(n15944), .B2(n17882), .A(n15943), .ZN(n15945) );
  OAI21_X1 U19471 ( .B1(n20989), .B2(n16172), .A(n15945), .ZN(P1_U2973) );
  NAND2_X1 U19472 ( .A1(n15946), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15958) );
  MUX2_X1 U19473 ( .A(n15947), .B(n15959), .S(n9688), .Z(n15948) );
  AOI21_X1 U19474 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15958), .A(
        n15948), .ZN(n15949) );
  XNOR2_X1 U19475 ( .A(n15949), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16180) );
  NAND2_X1 U19476 ( .A1(n17880), .A2(n15950), .ZN(n15951) );
  NAND2_X1 U19477 ( .A1(n17906), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n16173) );
  OAI211_X1 U19478 ( .C1(n17885), .C2(n15952), .A(n15951), .B(n16173), .ZN(
        n15953) );
  AOI21_X1 U19479 ( .B1(n15954), .B2(n17882), .A(n15953), .ZN(n15955) );
  OAI21_X1 U19480 ( .B1(n16180), .B2(n20989), .A(n15955), .ZN(P1_U2974) );
  NAND2_X1 U19481 ( .A1(n15956), .A2(n15958), .ZN(n15957) );
  MUX2_X1 U19482 ( .A(n15958), .B(n15957), .S(n16103), .Z(n15960) );
  XNOR2_X1 U19483 ( .A(n15960), .B(n15959), .ZN(n16191) );
  NAND2_X1 U19484 ( .A1(n17906), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n16181) );
  OAI21_X1 U19485 ( .B1(n17885), .B2(n15961), .A(n16181), .ZN(n15964) );
  NOR2_X1 U19486 ( .A1(n15962), .A2(n16117), .ZN(n15963) );
  AOI211_X1 U19487 ( .C1(n17880), .C2(n15965), .A(n15964), .B(n15963), .ZN(
        n15966) );
  OAI21_X1 U19488 ( .B1(n20989), .B2(n16191), .A(n15966), .ZN(P1_U2975) );
  XNOR2_X1 U19489 ( .A(n12890), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15968) );
  XNOR2_X1 U19490 ( .A(n15967), .B(n15968), .ZN(n16199) );
  NAND2_X1 U19491 ( .A1(n17880), .A2(n15969), .ZN(n15970) );
  NAND2_X1 U19492 ( .A1(n17906), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n16193) );
  OAI211_X1 U19493 ( .C1(n17885), .C2(n15971), .A(n15970), .B(n16193), .ZN(
        n15972) );
  AOI21_X1 U19494 ( .B1(n15973), .B2(n17882), .A(n15972), .ZN(n15974) );
  OAI21_X1 U19495 ( .B1(n16199), .B2(n20989), .A(n15974), .ZN(P1_U2976) );
  XNOR2_X1 U19496 ( .A(n12890), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16013) );
  OAI21_X1 U19497 ( .B1(n15977), .B2(n15976), .A(n12890), .ZN(n15979) );
  NAND2_X1 U19498 ( .A1(n15979), .A2(n15978), .ZN(n15980) );
  XNOR2_X1 U19499 ( .A(n15980), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16200) );
  NAND2_X1 U19500 ( .A1(n16200), .A2(n17883), .ZN(n15984) );
  NOR2_X1 U19501 ( .A1(n17899), .A2(n21699), .ZN(n16204) );
  NOR2_X1 U19502 ( .A1(n17877), .A2(n15981), .ZN(n15982) );
  AOI211_X1 U19503 ( .C1(n17870), .C2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16204), .B(n15982), .ZN(n15983) );
  OAI211_X1 U19504 ( .C1(n16117), .C2(n15985), .A(n15984), .B(n15983), .ZN(
        P1_U2977) );
  INV_X1 U19505 ( .A(n15975), .ZN(n15989) );
  NAND2_X1 U19506 ( .A1(n15986), .A2(n16246), .ZN(n15987) );
  NOR2_X1 U19507 ( .A1(n12890), .A2(n15987), .ZN(n15988) );
  NAND2_X1 U19508 ( .A1(n15989), .A2(n15988), .ZN(n15996) );
  XNOR2_X1 U19509 ( .A(n15990), .B(n16212), .ZN(n16217) );
  NOR2_X1 U19510 ( .A1(n17899), .A2(n21697), .ZN(n16209) );
  AOI21_X1 U19511 ( .B1(n17870), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16209), .ZN(n15991) );
  OAI21_X1 U19512 ( .B1(n15992), .B2(n17877), .A(n15991), .ZN(n15993) );
  AOI21_X1 U19513 ( .B1(n15994), .B2(n17882), .A(n15993), .ZN(n15995) );
  OAI21_X1 U19514 ( .B1(n16217), .B2(n20989), .A(n15995), .ZN(P1_U2978) );
  NAND2_X1 U19515 ( .A1(n15997), .A2(n15996), .ZN(n15998) );
  XNOR2_X1 U19516 ( .A(n15998), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16229) );
  NAND2_X1 U19517 ( .A1(n17880), .A2(n15999), .ZN(n16000) );
  NAND2_X1 U19518 ( .A1(n17906), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n16218) );
  OAI211_X1 U19519 ( .C1(n17885), .C2(n16001), .A(n16000), .B(n16218), .ZN(
        n16002) );
  AOI21_X1 U19520 ( .B1(n16003), .B2(n17882), .A(n16002), .ZN(n16004) );
  OAI21_X1 U19521 ( .B1(n16229), .B2(n20989), .A(n16004), .ZN(P1_U2979) );
  OAI21_X1 U19522 ( .B1(n16246), .B2(n9689), .A(n16012), .ZN(n16006) );
  XNOR2_X1 U19523 ( .A(n12890), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16005) );
  XNOR2_X1 U19524 ( .A(n16006), .B(n16005), .ZN(n16238) );
  INV_X1 U19525 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21693) );
  NOR2_X1 U19526 ( .A1(n17899), .A2(n21693), .ZN(n16233) );
  AOI21_X1 U19527 ( .B1(n17870), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16233), .ZN(n16007) );
  OAI21_X1 U19528 ( .B1(n16008), .B2(n17877), .A(n16007), .ZN(n16009) );
  AOI21_X1 U19529 ( .B1(n16010), .B2(n17882), .A(n16009), .ZN(n16011) );
  OAI21_X1 U19530 ( .B1(n16238), .B2(n20989), .A(n16011), .ZN(P1_U2980) );
  OAI21_X1 U19531 ( .B1(n15975), .B2(n16013), .A(n16012), .ZN(n16250) );
  NOR2_X1 U19532 ( .A1(n17899), .A2(n16014), .ZN(n16242) );
  AOI21_X1 U19533 ( .B1(n17870), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16242), .ZN(n16015) );
  OAI21_X1 U19534 ( .B1(n16016), .B2(n17877), .A(n16015), .ZN(n16017) );
  AOI21_X1 U19535 ( .B1(n16018), .B2(n17882), .A(n16017), .ZN(n16019) );
  OAI21_X1 U19536 ( .B1(n20989), .B2(n16250), .A(n16019), .ZN(P1_U2981) );
  INV_X1 U19537 ( .A(n16020), .ZN(n16094) );
  NOR2_X1 U19538 ( .A1(n16094), .A2(n16021), .ZN(n16057) );
  AOI21_X1 U19539 ( .B1(n16057), .B2(n16022), .A(n9791), .ZN(n16023) );
  MUX2_X1 U19540 ( .A(n16024), .B(n16103), .S(n16023), .Z(n16025) );
  XOR2_X1 U19541 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n16025), .Z(
        n16258) );
  INV_X1 U19542 ( .A(n16026), .ZN(n16030) );
  NOR2_X1 U19543 ( .A1(n17899), .A2(n21690), .ZN(n16255) );
  AOI21_X1 U19544 ( .B1(n17870), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16255), .ZN(n16027) );
  OAI21_X1 U19545 ( .B1(n16028), .B2(n17877), .A(n16027), .ZN(n16029) );
  AOI21_X1 U19546 ( .B1(n16030), .B2(n17882), .A(n16029), .ZN(n16031) );
  OAI21_X1 U19547 ( .B1(n16258), .B2(n20989), .A(n16031), .ZN(P1_U2982) );
  OAI21_X1 U19548 ( .B1(n16020), .B2(n16033), .A(n16032), .ZN(n16046) );
  NOR2_X1 U19549 ( .A1(n16046), .A2(n16034), .ZN(n16048) );
  INV_X1 U19550 ( .A(n16047), .ZN(n16035) );
  NOR2_X1 U19551 ( .A1(n16048), .A2(n16035), .ZN(n16036) );
  XOR2_X1 U19552 ( .A(n16037), .B(n16036), .Z(n16268) );
  INV_X1 U19553 ( .A(n16268), .ZN(n16043) );
  NAND2_X1 U19554 ( .A1(n17906), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n16264) );
  NAND2_X1 U19555 ( .A1(n17870), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16038) );
  OAI211_X1 U19556 ( .C1(n17877), .C2(n16039), .A(n16264), .B(n16038), .ZN(
        n16040) );
  AOI21_X1 U19557 ( .B1(n16041), .B2(n17882), .A(n16040), .ZN(n16042) );
  OAI21_X1 U19558 ( .B1(n16043), .B2(n20989), .A(n16042), .ZN(P1_U2983) );
  NAND2_X1 U19559 ( .A1(n16044), .A2(n16047), .ZN(n16045) );
  AOI22_X1 U19560 ( .A1(n16048), .A2(n16047), .B1(n16046), .B2(n16045), .ZN(
        n16277) );
  NAND2_X1 U19561 ( .A1(n17906), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n16272) );
  NAND2_X1 U19562 ( .A1(n17870), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16049) );
  OAI211_X1 U19563 ( .C1(n17877), .C2(n16050), .A(n16272), .B(n16049), .ZN(
        n16051) );
  AOI21_X1 U19564 ( .B1(n16052), .B2(n17882), .A(n16051), .ZN(n16053) );
  OAI21_X1 U19565 ( .B1(n16277), .B2(n20989), .A(n16053), .ZN(P1_U2984) );
  NAND2_X1 U19566 ( .A1(n16054), .A2(n16065), .ZN(n16056) );
  OAI21_X1 U19567 ( .B1(n16057), .B2(n16056), .A(n16055), .ZN(n16059) );
  XNOR2_X1 U19568 ( .A(n9689), .B(n16287), .ZN(n16058) );
  XNOR2_X1 U19569 ( .A(n16059), .B(n16058), .ZN(n16278) );
  NAND2_X1 U19570 ( .A1(n16278), .A2(n17883), .ZN(n16063) );
  NOR2_X1 U19571 ( .A1(n17899), .A2(n21682), .ZN(n16283) );
  NOR2_X1 U19572 ( .A1(n17877), .A2(n16060), .ZN(n16061) );
  AOI211_X1 U19573 ( .C1(n17870), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16283), .B(n16061), .ZN(n16062) );
  OAI211_X1 U19574 ( .C1(n16117), .C2(n16064), .A(n16063), .B(n16062), .ZN(
        P1_U2985) );
  INV_X1 U19575 ( .A(n16065), .ZN(n16066) );
  OR2_X1 U19576 ( .A1(n16020), .A2(n16066), .ZN(n16069) );
  NOR2_X1 U19577 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16067) );
  OR2_X1 U19578 ( .A1(n9688), .A2(n16067), .ZN(n16068) );
  NAND2_X1 U19579 ( .A1(n16069), .A2(n16068), .ZN(n16084) );
  NOR2_X1 U19580 ( .A1(n12890), .A2(n16070), .ZN(n16071) );
  OR2_X1 U19581 ( .A1(n16072), .A2(n16071), .ZN(n16083) );
  INV_X1 U19582 ( .A(n16072), .ZN(n16073) );
  NAND2_X1 U19583 ( .A1(n16081), .A2(n16073), .ZN(n16075) );
  XNOR2_X1 U19584 ( .A(n16075), .B(n16074), .ZN(n16295) );
  INV_X1 U19585 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21684) );
  NOR2_X1 U19586 ( .A1(n17899), .A2(n21684), .ZN(n16289) );
  AOI21_X1 U19587 ( .B1(n17870), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16289), .ZN(n16076) );
  OAI21_X1 U19588 ( .B1(n16077), .B2(n17877), .A(n16076), .ZN(n16078) );
  AOI21_X1 U19589 ( .B1(n16079), .B2(n17882), .A(n16078), .ZN(n16080) );
  OAI21_X1 U19590 ( .B1(n20989), .B2(n16295), .A(n16080), .ZN(P1_U2986) );
  INV_X1 U19591 ( .A(n16081), .ZN(n16082) );
  AOI21_X1 U19592 ( .B1(n16084), .B2(n16083), .A(n16082), .ZN(n16311) );
  NOR2_X1 U19593 ( .A1(n17877), .A2(n16086), .ZN(n16089) );
  NAND2_X1 U19594 ( .A1(n17906), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n16302) );
  OAI21_X1 U19595 ( .B1(n17885), .B2(n16087), .A(n16302), .ZN(n16088) );
  INV_X1 U19596 ( .A(n16090), .ZN(n16092) );
  NAND2_X1 U19597 ( .A1(n9688), .A2(n16091), .ZN(n16121) );
  OAI21_X1 U19598 ( .B1(n16092), .B2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n16121), .ZN(n16093) );
  OAI21_X1 U19599 ( .B1(n17898), .B2(n16090), .A(n16093), .ZN(n16116) );
  NOR2_X1 U19600 ( .A1(n16116), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16102) );
  NAND3_X1 U19601 ( .A1(n16102), .A2(n16103), .A3(n16331), .ZN(n16106) );
  NAND3_X1 U19602 ( .A1(n16094), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n9689), .ZN(n16095) );
  NAND2_X1 U19603 ( .A1(n16106), .A2(n16095), .ZN(n16096) );
  XNOR2_X1 U19604 ( .A(n16096), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16320) );
  NOR2_X1 U19605 ( .A1(n17899), .A2(n21680), .ZN(n16314) );
  AOI21_X1 U19606 ( .B1(n17870), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16314), .ZN(n16097) );
  OAI21_X1 U19607 ( .B1(n16098), .B2(n17877), .A(n16097), .ZN(n16099) );
  AOI21_X1 U19608 ( .B1(n16100), .B2(n17882), .A(n16099), .ZN(n16101) );
  OAI21_X1 U19609 ( .B1(n16320), .B2(n20989), .A(n16101), .ZN(P1_U2988) );
  XNOR2_X1 U19610 ( .A(n16020), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16105) );
  NOR2_X1 U19611 ( .A1(n16102), .A2(n16331), .ZN(n16104) );
  MUX2_X1 U19612 ( .A(n16105), .B(n16104), .S(n16103), .Z(n16108) );
  INV_X1 U19613 ( .A(n16106), .ZN(n16107) );
  NOR2_X1 U19614 ( .A1(n16108), .A2(n16107), .ZN(n16337) );
  INV_X1 U19615 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n16109) );
  OR2_X1 U19616 ( .A1(n17899), .A2(n16109), .ZN(n16322) );
  NAND2_X1 U19617 ( .A1(n17870), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16110) );
  OAI211_X1 U19618 ( .C1(n17877), .C2(n16111), .A(n16322), .B(n16110), .ZN(
        n16112) );
  AOI21_X1 U19619 ( .B1(n16113), .B2(n17882), .A(n16112), .ZN(n16114) );
  OAI21_X1 U19620 ( .B1(n16337), .B2(n20989), .A(n16114), .ZN(P1_U2989) );
  XNOR2_X1 U19621 ( .A(n9689), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16115) );
  XNOR2_X1 U19622 ( .A(n16116), .B(n16115), .ZN(n16338) );
  INV_X1 U19623 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n21007) );
  NAND2_X1 U19624 ( .A1(n17906), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n16344) );
  OAI21_X1 U19625 ( .B1(n17885), .B2(n21007), .A(n16344), .ZN(n16119) );
  NOR2_X1 U19626 ( .A1(n21011), .A2(n16117), .ZN(n16118) );
  AOI211_X1 U19627 ( .C1(n17880), .C2(n21012), .A(n16119), .B(n16118), .ZN(
        n16120) );
  OAI21_X1 U19628 ( .B1(n16338), .B2(n20989), .A(n16120), .ZN(P1_U2990) );
  XNOR2_X1 U19629 ( .A(n16121), .B(n17898), .ZN(n16122) );
  XNOR2_X1 U19630 ( .A(n16090), .B(n16122), .ZN(n17896) );
  INV_X1 U19631 ( .A(n17896), .ZN(n16128) );
  AOI22_X1 U19632 ( .A1(n17870), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n17906), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n16123) );
  OAI21_X1 U19633 ( .B1(n16124), .B2(n17877), .A(n16123), .ZN(n16125) );
  AOI21_X1 U19634 ( .B1(n16126), .B2(n17882), .A(n16125), .ZN(n16127) );
  OAI21_X1 U19635 ( .B1(n16128), .B2(n20989), .A(n16127), .ZN(P1_U2991) );
  INV_X1 U19636 ( .A(n16129), .ZN(n16133) );
  AOI211_X1 U19637 ( .C1(n16134), .C2(n17922), .A(n16133), .B(n16132), .ZN(
        n16135) );
  OAI21_X1 U19638 ( .B1(n16136), .B2(n21175), .A(n16135), .ZN(P1_U3001) );
  INV_X1 U19639 ( .A(n16156), .ZN(n16138) );
  NOR3_X1 U19640 ( .A1(n16138), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n10497), .ZN(n16139) );
  AOI211_X1 U19641 ( .C1(n16141), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16140), .B(n16139), .ZN(n16144) );
  NAND2_X1 U19642 ( .A1(n16142), .A2(n17922), .ZN(n16143) );
  INV_X1 U19643 ( .A(n16159), .ZN(n16149) );
  AND3_X1 U19644 ( .A1(n16156), .A2(n10497), .A3(n16146), .ZN(n16147) );
  AOI211_X1 U19645 ( .C1(n16149), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16148), .B(n16147), .ZN(n16153) );
  INV_X1 U19646 ( .A(n16150), .ZN(n16151) );
  NAND2_X1 U19647 ( .A1(n16151), .A2(n17922), .ZN(n16152) );
  OAI211_X1 U19648 ( .C1(n16154), .C2(n21175), .A(n16153), .B(n16152), .ZN(
        P1_U3003) );
  AOI21_X1 U19649 ( .B1(n16156), .B2(n16158), .A(n16155), .ZN(n16157) );
  OAI21_X1 U19650 ( .B1(n16159), .B2(n16158), .A(n16157), .ZN(n16160) );
  AOI21_X1 U19651 ( .B1(n16161), .B2(n17922), .A(n16160), .ZN(n16162) );
  OAI21_X1 U19652 ( .B1(n16163), .B2(n21175), .A(n16162), .ZN(P1_U3004) );
  INV_X1 U19653 ( .A(n16174), .ZN(n16166) );
  AND3_X1 U19654 ( .A1(n16166), .A2(n16165), .A3(n16164), .ZN(n16167) );
  AOI211_X1 U19655 ( .C1(n16178), .C2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16168), .B(n16167), .ZN(n16171) );
  NAND2_X1 U19656 ( .A1(n16169), .A2(n17922), .ZN(n16170) );
  OAI211_X1 U19657 ( .C1(n16172), .C2(n21175), .A(n16171), .B(n16170), .ZN(
        P1_U3005) );
  OAI21_X1 U19658 ( .B1(n16174), .B2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n16173), .ZN(n16177) );
  NOR2_X1 U19659 ( .A1(n16175), .A2(n21174), .ZN(n16176) );
  AOI211_X1 U19660 ( .C1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n16178), .A(
        n16177), .B(n16176), .ZN(n16179) );
  OAI21_X1 U19661 ( .B1(n16180), .B2(n21175), .A(n16179), .ZN(P1_U3006) );
  INV_X1 U19662 ( .A(n16181), .ZN(n16188) );
  INV_X1 U19663 ( .A(n16301), .ZN(n16183) );
  INV_X1 U19664 ( .A(n16297), .ZN(n16300) );
  OAI21_X1 U19665 ( .B1(n16183), .B2(n16300), .A(n16182), .ZN(n16186) );
  INV_X1 U19666 ( .A(n16194), .ZN(n16184) );
  AOI21_X1 U19667 ( .B1(n16184), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16185) );
  AOI21_X1 U19668 ( .B1(n16192), .B2(n16186), .A(n16185), .ZN(n16187) );
  AOI211_X1 U19669 ( .C1(n16189), .C2(n17922), .A(n16188), .B(n16187), .ZN(
        n16190) );
  OAI21_X1 U19670 ( .B1(n16191), .B2(n21175), .A(n16190), .ZN(P1_U3007) );
  NOR2_X1 U19671 ( .A1(n16192), .A2(n12886), .ZN(n16196) );
  OAI21_X1 U19672 ( .B1(n16194), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16193), .ZN(n16195) );
  AOI211_X1 U19673 ( .C1(n16197), .C2(n17922), .A(n16196), .B(n16195), .ZN(
        n16198) );
  OAI21_X1 U19674 ( .B1(n16199), .B2(n21175), .A(n16198), .ZN(P1_U3008) );
  NAND2_X1 U19675 ( .A1(n16200), .A2(n17907), .ZN(n16207) );
  XNOR2_X1 U19676 ( .A(n16202), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16205) );
  INV_X1 U19677 ( .A(n16201), .ZN(n16213) );
  NOR2_X1 U19678 ( .A1(n16213), .A2(n16202), .ZN(n16203) );
  AOI211_X1 U19679 ( .C1(n16210), .C2(n16205), .A(n16204), .B(n16203), .ZN(
        n16206) );
  OAI211_X1 U19680 ( .C1(n21174), .C2(n16208), .A(n16207), .B(n16206), .ZN(
        P1_U3009) );
  AOI21_X1 U19681 ( .B1(n16210), .B2(n16212), .A(n16209), .ZN(n16211) );
  OAI21_X1 U19682 ( .B1(n16213), .B2(n16212), .A(n16211), .ZN(n16214) );
  AOI21_X1 U19683 ( .B1(n16215), .B2(n17922), .A(n16214), .ZN(n16216) );
  OAI21_X1 U19684 ( .B1(n16217), .B2(n21175), .A(n16216), .ZN(P1_U3010) );
  INV_X1 U19685 ( .A(n16218), .ZN(n16226) );
  INV_X1 U19686 ( .A(n16219), .ZN(n16220) );
  NOR3_X1 U19687 ( .A1(n16234), .A2(n21180), .A3(n16220), .ZN(n16222) );
  AOI211_X1 U19688 ( .C1(n16224), .C2(n16223), .A(n16222), .B(n16221), .ZN(
        n16225) );
  AOI211_X1 U19689 ( .C1(n16227), .C2(n17922), .A(n16226), .B(n16225), .ZN(
        n16228) );
  OAI21_X1 U19690 ( .B1(n16229), .B2(n21175), .A(n16228), .ZN(P1_U3011) );
  INV_X1 U19691 ( .A(n16292), .ZN(n16231) );
  NOR3_X1 U19692 ( .A1(n16231), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n16230), .ZN(n16232) );
  AOI211_X1 U19693 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16234), .A(
        n16233), .B(n16232), .ZN(n16237) );
  NAND2_X1 U19694 ( .A1(n16235), .A2(n17922), .ZN(n16236) );
  OAI211_X1 U19695 ( .C1(n16238), .C2(n21175), .A(n16237), .B(n16236), .ZN(
        P1_U3012) );
  AND2_X1 U19696 ( .A1(n16259), .A2(n16279), .ZN(n16239) );
  OR2_X1 U19697 ( .A1(n16240), .A2(n16239), .ZN(n16291) );
  AOI21_X1 U19698 ( .B1(n16259), .B2(n16241), .A(n16291), .ZN(n16252) );
  INV_X1 U19699 ( .A(n16242), .ZN(n16245) );
  NAND4_X1 U19700 ( .A1(n16292), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n16243), .A4(n16246), .ZN(n16244) );
  OAI211_X1 U19701 ( .C1(n16252), .C2(n16246), .A(n16245), .B(n16244), .ZN(
        n16247) );
  AOI21_X1 U19702 ( .B1(n16248), .B2(n17922), .A(n16247), .ZN(n16249) );
  OAI21_X1 U19703 ( .B1(n16250), .B2(n21175), .A(n16249), .ZN(P1_U3013) );
  AND2_X1 U19704 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16251) );
  AND2_X1 U19705 ( .A1(n16292), .A2(n16251), .ZN(n16262) );
  NAND3_X1 U19706 ( .A1(n16262), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16253) );
  AOI21_X1 U19707 ( .B1(n13061), .B2(n16253), .A(n16252), .ZN(n16254) );
  AOI211_X1 U19708 ( .C1(n16256), .C2(n17922), .A(n16255), .B(n16254), .ZN(
        n16257) );
  OAI21_X1 U19709 ( .B1(n16258), .B2(n21175), .A(n16257), .ZN(P1_U3014) );
  AOI21_X1 U19710 ( .B1(n16287), .B2(n16259), .A(n16291), .ZN(n16270) );
  NAND2_X1 U19711 ( .A1(n16262), .A2(n16260), .ZN(n16271) );
  AOI21_X1 U19712 ( .B1(n16270), .B2(n16271), .A(n16261), .ZN(n16267) );
  NAND3_X1 U19713 ( .A1(n16262), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n16261), .ZN(n16263) );
  OAI211_X1 U19714 ( .C1(n16265), .C2(n21174), .A(n16264), .B(n16263), .ZN(
        n16266) );
  AOI211_X1 U19715 ( .C1(n16268), .C2(n17907), .A(n16267), .B(n16266), .ZN(
        n16269) );
  INV_X1 U19716 ( .A(n16269), .ZN(P1_U3015) );
  INV_X1 U19717 ( .A(n16270), .ZN(n16275) );
  OAI211_X1 U19718 ( .C1(n16273), .C2(n21174), .A(n16272), .B(n16271), .ZN(
        n16274) );
  AOI21_X1 U19719 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16275), .A(
        n16274), .ZN(n16276) );
  OAI21_X1 U19720 ( .B1(n16277), .B2(n21175), .A(n16276), .ZN(P1_U3016) );
  INV_X1 U19721 ( .A(n16291), .ZN(n16288) );
  NAND2_X1 U19722 ( .A1(n16278), .A2(n17907), .ZN(n16286) );
  INV_X1 U19723 ( .A(n16334), .ZN(n16281) );
  NOR4_X1 U19724 ( .A1(n16281), .A2(n16280), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(n16279), .ZN(n16282) );
  AOI211_X1 U19725 ( .C1(n17922), .C2(n16284), .A(n16283), .B(n16282), .ZN(
        n16285) );
  OAI211_X1 U19726 ( .C1(n16288), .C2(n16287), .A(n16286), .B(n16285), .ZN(
        P1_U3017) );
  AOI21_X1 U19727 ( .B1(n16290), .B2(n17922), .A(n16289), .ZN(n16294) );
  OAI21_X1 U19728 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16292), .A(
        n16291), .ZN(n16293) );
  OAI211_X1 U19729 ( .C1(n16295), .C2(n21175), .A(n16294), .B(n16293), .ZN(
        P1_U3018) );
  OAI21_X1 U19730 ( .B1(n16329), .B2(n16297), .A(n16296), .ZN(n17889) );
  AOI21_X1 U19731 ( .B1(n16317), .B2(n16298), .A(n17886), .ZN(n16299) );
  AOI211_X1 U19732 ( .C1(n16300), .C2(n16305), .A(n17889), .B(n16299), .ZN(
        n16312) );
  OAI21_X1 U19733 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16301), .A(
        n16312), .ZN(n16309) );
  OAI21_X1 U19734 ( .B1(n16303), .B2(n21174), .A(n16302), .ZN(n16308) );
  INV_X1 U19735 ( .A(n17910), .ZN(n16306) );
  NOR3_X1 U19736 ( .A1(n16306), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n16305), .ZN(n16307) );
  AOI211_X1 U19737 ( .C1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n16309), .A(
        n16308), .B(n16307), .ZN(n16310) );
  OAI21_X1 U19738 ( .B1(n16311), .B2(n21175), .A(n16310), .ZN(P1_U3019) );
  NOR2_X1 U19739 ( .A1(n16312), .A2(n16316), .ZN(n16313) );
  AOI211_X1 U19740 ( .C1(n17922), .C2(n16315), .A(n16314), .B(n16313), .ZN(
        n16319) );
  NAND3_X1 U19741 ( .A1(n17910), .A2(n16317), .A3(n16316), .ZN(n16318) );
  OAI211_X1 U19742 ( .C1(n16320), .C2(n21175), .A(n16319), .B(n16318), .ZN(
        P1_U3020) );
  INV_X1 U19743 ( .A(n16329), .ZN(n16321) );
  INV_X1 U19744 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16339) );
  NOR4_X1 U19745 ( .A1(n16321), .A2(n16327), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A4(n16339), .ZN(n16335) );
  OAI21_X1 U19746 ( .B1(n16323), .B2(n21174), .A(n16322), .ZN(n16333) );
  NAND3_X1 U19747 ( .A1(n16325), .A2(n16329), .A3(n16324), .ZN(n16326) );
  NAND2_X1 U19748 ( .A1(n16326), .A2(n17892), .ZN(n16340) );
  NOR2_X1 U19749 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16327), .ZN(
        n16328) );
  AND2_X1 U19750 ( .A1(n16329), .A2(n16328), .ZN(n16330) );
  NAND2_X1 U19751 ( .A1(n16334), .A2(n16330), .ZN(n16345) );
  AOI21_X1 U19752 ( .B1(n16340), .B2(n16345), .A(n16331), .ZN(n16332) );
  AOI211_X1 U19753 ( .C1(n16335), .C2(n16334), .A(n16333), .B(n16332), .ZN(
        n16336) );
  OAI21_X1 U19754 ( .B1(n16337), .B2(n21175), .A(n16336), .ZN(P1_U3021) );
  NOR2_X1 U19755 ( .A1(n16338), .A2(n21175), .ZN(n16348) );
  NOR2_X1 U19756 ( .A1(n16340), .A2(n16339), .ZN(n16347) );
  NAND2_X1 U19757 ( .A1(n15761), .A2(n16341), .ZN(n16342) );
  NAND2_X1 U19758 ( .A1(n16343), .A2(n16342), .ZN(n21005) );
  OAI211_X1 U19759 ( .C1(n21174), .C2(n21005), .A(n16345), .B(n16344), .ZN(
        n16346) );
  OR3_X1 U19760 ( .A1(n16348), .A2(n16347), .A3(n16346), .ZN(P1_U3022) );
  NOR2_X1 U19761 ( .A1(n14304), .A2(n12518), .ZN(n16356) );
  AOI21_X1 U19762 ( .B1(n16350), .B2(n16356), .A(n16349), .ZN(n16351) );
  OAI21_X1 U19763 ( .B1(n21453), .B2(n16352), .A(n16351), .ZN(n17826) );
  INV_X1 U19764 ( .A(n17826), .ZN(n16359) );
  INV_X1 U19765 ( .A(n21733), .ZN(n16358) );
  INV_X1 U19766 ( .A(n16353), .ZN(n16354) );
  AOI22_X1 U19767 ( .A1(n21732), .A2(n16356), .B1(n16355), .B2(n16354), .ZN(
        n16357) );
  OAI21_X1 U19768 ( .B1(n16359), .B2(n16358), .A(n16357), .ZN(n16361) );
  MUX2_X1 U19769 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n16361), .S(
        n16360), .Z(P1_U3473) );
  NOR3_X1 U19770 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21575), .A3(
        n21574), .ZN(n16367) );
  OAI21_X1 U19771 ( .B1(n21632), .B2(n16393), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n16363) );
  NOR2_X1 U19772 ( .A1(n21527), .A2(n21453), .ZN(n16366) );
  INV_X1 U19773 ( .A(n16366), .ZN(n16362) );
  AOI21_X1 U19774 ( .B1(n16363), .B2(n16362), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n16364) );
  OR2_X1 U19775 ( .A1(n21393), .A2(n12902), .ZN(n16365) );
  NAND2_X1 U19776 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n16365), .ZN(n21461) );
  NAND2_X1 U19777 ( .A1(n16389), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n16370) );
  INV_X1 U19778 ( .A(n16365), .ZN(n21456) );
  AOI22_X1 U19779 ( .A1(n16366), .A2(n21586), .B1(n21190), .B2(n21456), .ZN(
        n16391) );
  INV_X1 U19780 ( .A(n16367), .ZN(n16390) );
  OAI22_X1 U19781 ( .A1(n21466), .A2(n16391), .B1(n21291), .B2(n16390), .ZN(
        n16368) );
  AOI21_X1 U19782 ( .B1(n16393), .B2(n21587), .A(n16368), .ZN(n16369) );
  OAI211_X1 U19783 ( .C1(n21590), .C2(n16396), .A(n16370), .B(n16369), .ZN(
        P1_U3145) );
  NAND2_X1 U19784 ( .A1(n16389), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n16373) );
  OAI22_X1 U19785 ( .A1(n21469), .A2(n16391), .B1(n16390), .B2(n21304), .ZN(
        n16371) );
  AOI21_X1 U19786 ( .B1(n16393), .B2(n21593), .A(n16371), .ZN(n16372) );
  OAI211_X1 U19787 ( .C1(n21596), .C2(n16396), .A(n16373), .B(n16372), .ZN(
        P1_U3146) );
  NAND2_X1 U19788 ( .A1(n16389), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n16376) );
  OAI22_X1 U19789 ( .A1(n21472), .A2(n16391), .B1(n16390), .B2(n21308), .ZN(
        n16374) );
  AOI21_X1 U19790 ( .B1(n16393), .B2(n21599), .A(n16374), .ZN(n16375) );
  OAI211_X1 U19791 ( .C1(n21602), .C2(n16396), .A(n16376), .B(n16375), .ZN(
        P1_U3147) );
  NAND2_X1 U19792 ( .A1(n16389), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n16379) );
  OAI22_X1 U19793 ( .A1(n21475), .A2(n16391), .B1(n16390), .B2(n21312), .ZN(
        n16377) );
  AOI21_X1 U19794 ( .B1(n16393), .B2(n21605), .A(n16377), .ZN(n16378) );
  OAI211_X1 U19795 ( .C1(n21608), .C2(n16396), .A(n16379), .B(n16378), .ZN(
        P1_U3148) );
  NAND2_X1 U19796 ( .A1(n16389), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n16382) );
  OAI22_X1 U19797 ( .A1(n21478), .A2(n16391), .B1(n16390), .B2(n21316), .ZN(
        n16380) );
  AOI21_X1 U19798 ( .B1(n16393), .B2(n21611), .A(n16380), .ZN(n16381) );
  OAI211_X1 U19799 ( .C1(n21614), .C2(n16396), .A(n16382), .B(n16381), .ZN(
        P1_U3149) );
  NAND2_X1 U19800 ( .A1(n16389), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n16385) );
  OAI22_X1 U19801 ( .A1(n21481), .A2(n16391), .B1(n16390), .B2(n21320), .ZN(
        n16383) );
  AOI21_X1 U19802 ( .B1(n16393), .B2(n21617), .A(n16383), .ZN(n16384) );
  OAI211_X1 U19803 ( .C1(n21620), .C2(n16396), .A(n16385), .B(n16384), .ZN(
        P1_U3150) );
  NAND2_X1 U19804 ( .A1(n16389), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n16388) );
  OAI22_X1 U19805 ( .A1(n21484), .A2(n16391), .B1(n16390), .B2(n21324), .ZN(
        n16386) );
  AOI21_X1 U19806 ( .B1(n16393), .B2(n21623), .A(n16386), .ZN(n16387) );
  OAI211_X1 U19807 ( .C1(n21626), .C2(n16396), .A(n16388), .B(n16387), .ZN(
        P1_U3151) );
  NAND2_X1 U19808 ( .A1(n16389), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n16395) );
  OAI22_X1 U19809 ( .A1(n21490), .A2(n16391), .B1(n16390), .B2(n21328), .ZN(
        n16392) );
  AOI21_X1 U19810 ( .B1(n16393), .B2(n21631), .A(n16392), .ZN(n16394) );
  OAI211_X1 U19811 ( .C1(n21637), .C2(n16396), .A(n16395), .B(n16394), .ZN(
        P1_U3152) );
  INV_X1 U19812 ( .A(n16397), .ZN(n16416) );
  INV_X1 U19813 ( .A(n16398), .ZN(n16399) );
  AOI21_X1 U19814 ( .B1(n16416), .B2(n16399), .A(n20177), .ZN(n16401) );
  OAI21_X1 U19815 ( .B1(n16401), .B2(n20107), .A(n16400), .ZN(n16408) );
  INV_X1 U19816 ( .A(n16402), .ZN(n16780) );
  AOI22_X1 U19817 ( .A1(n20150), .A2(P2_REIP_REG_28__SCAN_IN), .B1(n20126), 
        .B2(P2_EBX_REG_28__SCAN_IN), .ZN(n16404) );
  NAND2_X1 U19818 ( .A1(n20186), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16403) );
  OAI211_X1 U19819 ( .C1(n16405), .C2(n20165), .A(n16404), .B(n16403), .ZN(
        n16406) );
  AOI21_X1 U19820 ( .B1(n16780), .B2(n20185), .A(n16406), .ZN(n16407) );
  OAI211_X1 U19821 ( .C1(n20189), .C2(n16682), .A(n16408), .B(n16407), .ZN(
        P2_U2827) );
  NAND2_X1 U19822 ( .A1(n16409), .A2(n20187), .ZN(n16411) );
  AOI22_X1 U19823 ( .A1(n20150), .A2(P2_REIP_REG_27__SCAN_IN), .B1(n20126), 
        .B2(P2_EBX_REG_27__SCAN_IN), .ZN(n16410) );
  OAI211_X1 U19824 ( .C1(n20145), .C2(n16412), .A(n16411), .B(n16410), .ZN(
        n16413) );
  AOI21_X1 U19825 ( .B1(n16788), .B2(n20185), .A(n16413), .ZN(n16419) );
  AOI21_X1 U19826 ( .B1(n16414), .B2(n16415), .A(n20177), .ZN(n16417) );
  OAI21_X1 U19827 ( .B1(n20107), .B2(n16417), .A(n16416), .ZN(n16418) );
  OAI211_X1 U19828 ( .C1(n14798), .C2(n20189), .A(n16419), .B(n16418), .ZN(
        P2_U2828) );
  NAND2_X1 U19829 ( .A1(n16436), .A2(n16420), .ZN(n16421) );
  NAND2_X1 U19830 ( .A1(n10553), .A2(n16421), .ZN(n17209) );
  AOI22_X1 U19831 ( .A1(n20150), .A2(P2_REIP_REG_26__SCAN_IN), .B1(n20169), 
        .B2(P2_EBX_REG_26__SCAN_IN), .ZN(n16422) );
  OAI21_X1 U19832 ( .B1(n16423), .B2(n20145), .A(n16422), .ZN(n16428) );
  NAND2_X1 U19833 ( .A1(n16425), .A2(n16424), .ZN(n16426) );
  NAND2_X1 U19834 ( .A1(n9772), .A2(n16426), .ZN(n17208) );
  NOR2_X1 U19835 ( .A1(n17208), .A2(n20171), .ZN(n16427) );
  AOI211_X1 U19836 ( .C1(n20187), .C2(n16429), .A(n16428), .B(n16427), .ZN(
        n16433) );
  INV_X1 U19837 ( .A(n16442), .ZN(n16430) );
  AOI21_X1 U19838 ( .B1(n16430), .B2(n10330), .A(n20177), .ZN(n16431) );
  OAI21_X1 U19839 ( .B1(n16431), .B2(n20107), .A(n16414), .ZN(n16432) );
  OAI211_X1 U19840 ( .C1(n20189), .C2(n17209), .A(n16433), .B(n16432), .ZN(
        P2_U2829) );
  OR2_X1 U19841 ( .A1(n16454), .A2(n16434), .ZN(n16435) );
  NAND2_X1 U19842 ( .A1(n16436), .A2(n16435), .ZN(n17223) );
  XNOR2_X1 U19843 ( .A(n9745), .B(n16437), .ZN(n16446) );
  AOI22_X1 U19844 ( .A1(n20150), .A2(P2_REIP_REG_25__SCAN_IN), .B1(n20169), 
        .B2(P2_EBX_REG_25__SCAN_IN), .ZN(n16438) );
  OAI21_X1 U19845 ( .B1(n10354), .B2(n20145), .A(n16438), .ZN(n16445) );
  INV_X1 U19846 ( .A(n16439), .ZN(n16441) );
  INV_X1 U19847 ( .A(n16942), .ZN(n16440) );
  OAI21_X1 U19848 ( .B1(n16441), .B2(n16440), .A(n20197), .ZN(n16443) );
  AOI21_X1 U19849 ( .B1(n17819), .B2(n16443), .A(n16442), .ZN(n16444) );
  AOI211_X1 U19850 ( .C1(n20187), .C2(n16446), .A(n16445), .B(n16444), .ZN(
        n16450) );
  XOR2_X1 U19851 ( .A(n16448), .B(n16447), .Z(n17225) );
  NAND2_X1 U19852 ( .A1(n17225), .A2(n20185), .ZN(n16449) );
  OAI211_X1 U19853 ( .C1(n20189), .C2(n17223), .A(n16450), .B(n16449), .ZN(
        P2_U2830) );
  INV_X1 U19854 ( .A(n16451), .ZN(n16719) );
  INV_X1 U19855 ( .A(n16485), .ZN(n16452) );
  NAND2_X1 U19856 ( .A1(n16719), .A2(n16452), .ZN(n16483) );
  AND2_X1 U19857 ( .A1(n16483), .A2(n16453), .ZN(n16455) );
  OR2_X1 U19858 ( .A1(n16455), .A2(n16454), .ZN(n17235) );
  AND2_X1 U19859 ( .A1(n16456), .A2(n16457), .ZN(n16458) );
  OR2_X1 U19860 ( .A1(n16458), .A2(n16447), .ZN(n17234) );
  INV_X1 U19861 ( .A(n16951), .ZN(n16459) );
  AOI21_X1 U19862 ( .B1(n16477), .B2(n16459), .A(n20177), .ZN(n16460) );
  OAI21_X1 U19863 ( .B1(n16460), .B2(n20107), .A(n16439), .ZN(n16467) );
  AOI21_X1 U19864 ( .B1(n16461), .B2(P2_EBX_REG_24__SCAN_IN), .A(n20165), .ZN(
        n16465) );
  NAND2_X1 U19865 ( .A1(n20150), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n16463) );
  NAND2_X1 U19866 ( .A1(n20126), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n16462) );
  OAI211_X1 U19867 ( .C1(n20145), .C2(n11624), .A(n16463), .B(n16462), .ZN(
        n16464) );
  AOI21_X1 U19868 ( .B1(n16465), .B2(n9745), .A(n16464), .ZN(n16466) );
  OAI211_X1 U19869 ( .C1(n20171), .C2(n17234), .A(n16467), .B(n16466), .ZN(
        n16468) );
  INV_X1 U19870 ( .A(n16468), .ZN(n16469) );
  OAI21_X1 U19871 ( .B1(n17235), .B2(n20189), .A(n16469), .ZN(P2_U2831) );
  INV_X1 U19872 ( .A(n16470), .ZN(n16822) );
  NAND2_X1 U19873 ( .A1(n16822), .A2(n16471), .ZN(n16472) );
  NAND2_X1 U19874 ( .A1(n16456), .A2(n16472), .ZN(n17248) );
  INV_X1 U19875 ( .A(n16473), .ZN(n16482) );
  AOI22_X1 U19876 ( .A1(n20150), .A2(P2_REIP_REG_23__SCAN_IN), .B1(n20169), 
        .B2(P2_EBX_REG_23__SCAN_IN), .ZN(n16474) );
  OAI21_X1 U19877 ( .B1(n16475), .B2(n20145), .A(n16474), .ZN(n16481) );
  INV_X1 U19878 ( .A(n16476), .ZN(n17817) );
  OAI21_X1 U19879 ( .B1(n17817), .B2(n16962), .A(n20197), .ZN(n16479) );
  INV_X1 U19880 ( .A(n16477), .ZN(n16478) );
  AOI21_X1 U19881 ( .B1(n17819), .B2(n16479), .A(n16478), .ZN(n16480) );
  AOI211_X1 U19882 ( .C1(n20187), .C2(n16482), .A(n16481), .B(n16480), .ZN(
        n16487) );
  INV_X1 U19883 ( .A(n16483), .ZN(n16484) );
  AOI21_X1 U19884 ( .B1(n16485), .B2(n16451), .A(n16484), .ZN(n17240) );
  NAND2_X1 U19885 ( .A1(n17240), .A2(n20129), .ZN(n16486) );
  OAI211_X1 U19886 ( .C1(n20171), .C2(n17248), .A(n16487), .B(n16486), .ZN(
        P2_U2832) );
  AOI21_X1 U19887 ( .B1(n16488), .B2(n10325), .A(n20177), .ZN(n16490) );
  OAI21_X1 U19888 ( .B1(n16490), .B2(n20107), .A(n17814), .ZN(n16496) );
  AOI22_X1 U19889 ( .A1(n20150), .A2(P2_REIP_REG_21__SCAN_IN), .B1(n20126), 
        .B2(P2_EBX_REG_21__SCAN_IN), .ZN(n16492) );
  NAND2_X1 U19890 ( .A1(n20186), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16491) );
  OAI211_X1 U19891 ( .C1(n16493), .C2(n20165), .A(n16492), .B(n16491), .ZN(
        n16494) );
  INV_X1 U19892 ( .A(n16494), .ZN(n16495) );
  OAI211_X1 U19893 ( .C1(n20171), .C2(n16831), .A(n16496), .B(n16495), .ZN(
        n16497) );
  INV_X1 U19894 ( .A(n16497), .ZN(n16498) );
  OAI21_X1 U19895 ( .B1(n16725), .B2(n20189), .A(n16498), .ZN(P2_U2834) );
  AND2_X1 U19896 ( .A1(n16500), .A2(n16499), .ZN(n16501) );
  OR2_X1 U19897 ( .A1(n16501), .A2(n14863), .ZN(n17271) );
  AOI21_X1 U19898 ( .B1(n16502), .B2(n11498), .A(n14871), .ZN(n17268) );
  NAND2_X1 U19899 ( .A1(n16503), .A2(n20187), .ZN(n16505) );
  AOI22_X1 U19900 ( .A1(n20150), .A2(P2_REIP_REG_20__SCAN_IN), .B1(n20169), 
        .B2(P2_EBX_REG_20__SCAN_IN), .ZN(n16504) );
  OAI211_X1 U19901 ( .C1(n20145), .C2(n16506), .A(n16505), .B(n16504), .ZN(
        n16511) );
  INV_X1 U19902 ( .A(n16516), .ZN(n16507) );
  OAI21_X1 U19903 ( .B1(n16507), .B2(n16983), .A(n20197), .ZN(n16509) );
  INV_X1 U19904 ( .A(n16488), .ZN(n16508) );
  AOI21_X1 U19905 ( .B1(n17819), .B2(n16509), .A(n16508), .ZN(n16510) );
  AOI211_X1 U19906 ( .C1(n20185), .C2(n17268), .A(n16511), .B(n16510), .ZN(
        n16512) );
  OAI21_X1 U19907 ( .B1(n17271), .B2(n20189), .A(n16512), .ZN(P2_U2835) );
  INV_X1 U19908 ( .A(n16513), .ZN(n16514) );
  AOI21_X1 U19909 ( .B1(n16515), .B2(n16514), .A(n20177), .ZN(n16517) );
  OAI21_X1 U19910 ( .B1(n16517), .B2(n20107), .A(n16516), .ZN(n16523) );
  AOI21_X1 U19911 ( .B1(n20169), .B2(P2_EBX_REG_19__SCAN_IN), .A(n20167), .ZN(
        n16519) );
  NAND2_X1 U19912 ( .A1(n20150), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n16518) );
  OAI211_X1 U19913 ( .C1(n20145), .C2(n16520), .A(n16519), .B(n16518), .ZN(
        n16521) );
  AOI21_X1 U19914 ( .B1(n9765), .B2(n20187), .A(n16521), .ZN(n16522) );
  OAI211_X1 U19915 ( .C1(n16855), .C2(n20171), .A(n16523), .B(n16522), .ZN(
        n16524) );
  AOI21_X1 U19916 ( .B1(n16733), .B2(n20129), .A(n16524), .ZN(n16525) );
  INV_X1 U19917 ( .A(n16525), .ZN(P2_U2836) );
  OAI21_X1 U19918 ( .B1(n16528), .B2(n16527), .A(n16526), .ZN(n17276) );
  XOR2_X1 U19919 ( .A(n16993), .B(n16529), .Z(n16538) );
  AOI21_X1 U19920 ( .B1(n20169), .B2(P2_EBX_REG_18__SCAN_IN), .A(n20167), .ZN(
        n16530) );
  OAI21_X1 U19921 ( .B1(n16992), .B2(n20180), .A(n16530), .ZN(n16531) );
  AOI21_X1 U19922 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20186), .A(
        n16531), .ZN(n16532) );
  OAI21_X1 U19923 ( .B1(n16533), .B2(n20165), .A(n16532), .ZN(n16537) );
  OAI21_X1 U19924 ( .B1(n14839), .B2(n16535), .A(n16534), .ZN(n17283) );
  NOR2_X1 U19925 ( .A1(n17283), .A2(n20171), .ZN(n16536) );
  AOI211_X1 U19926 ( .C1(n20197), .C2(n16538), .A(n16537), .B(n16536), .ZN(
        n16539) );
  OAI21_X1 U19927 ( .B1(n17276), .B2(n20189), .A(n16539), .ZN(P2_U2837) );
  INV_X1 U19928 ( .A(n16540), .ZN(n17321) );
  AOI22_X1 U19929 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(n20169), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n20150), .ZN(n16541) );
  OAI211_X1 U19930 ( .C1(n20145), .C2(n10343), .A(n16541), .B(n20181), .ZN(
        n16542) );
  AOI21_X1 U19931 ( .B1(n16543), .B2(n20187), .A(n16542), .ZN(n16546) );
  OAI211_X1 U19932 ( .C1(n16544), .C2(n17041), .A(n16616), .B(n20118), .ZN(
        n16545) );
  OAI211_X1 U19933 ( .C1(n17819), .C2(n17041), .A(n16546), .B(n16545), .ZN(
        n16547) );
  AOI21_X1 U19934 ( .B1(n20185), .B2(n17321), .A(n16547), .ZN(n16548) );
  OAI21_X1 U19935 ( .B1(n20189), .B2(n17323), .A(n16548), .ZN(P2_U2842) );
  AOI21_X1 U19936 ( .B1(n20169), .B2(P2_EBX_REG_12__SCAN_IN), .A(n20167), .ZN(
        n16549) );
  OAI21_X1 U19937 ( .B1(n20867), .B2(n20180), .A(n16549), .ZN(n16552) );
  NOR2_X1 U19938 ( .A1(n16550), .A2(n20165), .ZN(n16551) );
  AOI211_X1 U19939 ( .C1(n20186), .C2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16552), .B(n16551), .ZN(n16553) );
  OAI21_X1 U19940 ( .B1(n17338), .B2(n20189), .A(n16553), .ZN(n16558) );
  INV_X1 U19941 ( .A(n16555), .ZN(n16554) );
  AOI21_X1 U19942 ( .B1(n15422), .B2(n16554), .A(n20177), .ZN(n16556) );
  NOR2_X1 U19943 ( .A1(n16649), .A2(n16555), .ZN(n16562) );
  MUX2_X1 U19944 ( .A(n16556), .B(n16562), .S(n17057), .Z(n16557) );
  AOI211_X1 U19945 ( .C1(n20185), .C2(n17335), .A(n16558), .B(n16557), .ZN(
        n16559) );
  INV_X1 U19946 ( .A(n16559), .ZN(P2_U2843) );
  INV_X1 U19947 ( .A(n17069), .ZN(n16571) );
  NAND2_X1 U19948 ( .A1(n16560), .A2(n17069), .ZN(n16561) );
  AOI22_X1 U19949 ( .A1(n16562), .A2(n16561), .B1(n20129), .B2(n17352), .ZN(
        n16570) );
  INV_X1 U19950 ( .A(n17347), .ZN(n16568) );
  AOI21_X1 U19951 ( .B1(n20169), .B2(P2_EBX_REG_11__SCAN_IN), .A(n20167), .ZN(
        n16563) );
  OAI21_X1 U19952 ( .B1(n20865), .B2(n20180), .A(n16563), .ZN(n16564) );
  AOI21_X1 U19953 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n20186), .A(
        n16564), .ZN(n16565) );
  OAI21_X1 U19954 ( .B1(n16566), .B2(n20165), .A(n16565), .ZN(n16567) );
  AOI21_X1 U19955 ( .B1(n16568), .B2(n20185), .A(n16567), .ZN(n16569) );
  OAI211_X1 U19956 ( .C1(n16571), .C2(n17819), .A(n16570), .B(n16569), .ZN(
        P2_U2844) );
  NAND2_X1 U19957 ( .A1(n16616), .A2(n20163), .ZN(n16574) );
  NOR2_X1 U19958 ( .A1(n20163), .A2(n20177), .ZN(n16572) );
  NOR2_X1 U19959 ( .A1(n20107), .A2(n16572), .ZN(n16573) );
  MUX2_X1 U19960 ( .A(n16574), .B(n16573), .S(n17116), .Z(n16582) );
  INV_X1 U19961 ( .A(n17380), .ZN(n16580) );
  AOI21_X1 U19962 ( .B1(n20169), .B2(P2_EBX_REG_8__SCAN_IN), .A(n20167), .ZN(
        n16575) );
  OAI21_X1 U19963 ( .B1(n17115), .B2(n20180), .A(n16575), .ZN(n16576) );
  AOI21_X1 U19964 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n20186), .A(
        n16576), .ZN(n16577) );
  OAI21_X1 U19965 ( .B1(n16578), .B2(n20165), .A(n16577), .ZN(n16579) );
  AOI21_X1 U19966 ( .B1(n16580), .B2(n20185), .A(n16579), .ZN(n16581) );
  OAI211_X1 U19967 ( .C1(n20189), .C2(n17386), .A(n16582), .B(n16581), .ZN(
        P2_U2847) );
  AND2_X1 U19968 ( .A1(n16584), .A2(n20197), .ZN(n16583) );
  NOR2_X1 U19969 ( .A1(n20107), .A2(n16583), .ZN(n16587) );
  INV_X1 U19970 ( .A(n16584), .ZN(n16585) );
  NAND2_X1 U19971 ( .A1(n16616), .A2(n16585), .ZN(n16586) );
  MUX2_X1 U19972 ( .A(n16587), .B(n16586), .S(n17135), .Z(n16596) );
  OAI21_X1 U19973 ( .B1(n16588), .B2(n20182), .A(n17149), .ZN(n16590) );
  NOR2_X1 U19974 ( .A1(n20180), .A2(n20856), .ZN(n16589) );
  AOI211_X1 U19975 ( .C1(n20186), .C2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16590), .B(n16589), .ZN(n16591) );
  OAI21_X1 U19976 ( .B1(n16592), .B2(n20165), .A(n16591), .ZN(n16593) );
  AOI21_X1 U19977 ( .B1(n16594), .B2(n20129), .A(n16593), .ZN(n16595) );
  OAI211_X1 U19978 ( .C1(n17408), .C2(n20171), .A(n16596), .B(n16595), .ZN(
        P2_U2849) );
  NAND2_X1 U19979 ( .A1(n16599), .A2(n16598), .ZN(n16600) );
  NAND2_X1 U19980 ( .A1(n16597), .A2(n16600), .ZN(n17443) );
  NOR2_X1 U19981 ( .A1(n16601), .A2(n20165), .ZN(n16604) );
  INV_X1 U19982 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n20851) );
  OAI22_X1 U19983 ( .A1(n20182), .A2(n16602), .B1(n20851), .B2(n20180), .ZN(
        n16603) );
  AOI211_X1 U19984 ( .C1(n20186), .C2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n16604), .B(n16603), .ZN(n16605) );
  OAI21_X1 U19985 ( .B1(n17443), .B2(n20171), .A(n16605), .ZN(n16611) );
  NAND2_X1 U19986 ( .A1(n16607), .A2(n20197), .ZN(n16606) );
  NAND2_X1 U19987 ( .A1(n17819), .A2(n16606), .ZN(n16609) );
  NOR2_X1 U19988 ( .A1(n16649), .A2(n16607), .ZN(n16608) );
  MUX2_X1 U19989 ( .A(n16609), .B(n16608), .S(n17174), .Z(n16610) );
  AOI211_X1 U19990 ( .C1(n20129), .C2(n17446), .A(n16611), .B(n16610), .ZN(
        n16612) );
  OAI21_X1 U19991 ( .B1(n20324), .B2(n20190), .A(n16612), .ZN(P2_U2852) );
  AND2_X1 U19992 ( .A1(n16614), .A2(n20197), .ZN(n16613) );
  NOR2_X1 U19993 ( .A1(n20107), .A2(n16613), .ZN(n16618) );
  INV_X1 U19994 ( .A(n16614), .ZN(n16615) );
  NAND2_X1 U19995 ( .A1(n16616), .A2(n16615), .ZN(n16617) );
  MUX2_X1 U19996 ( .A(n16618), .B(n16617), .S(n17184), .Z(n16626) );
  NAND2_X1 U19997 ( .A1(n20923), .A2(n20185), .ZN(n16622) );
  OAI22_X1 U19998 ( .A1(n16619), .A2(n20182), .B1(n20849), .B2(n20180), .ZN(
        n16620) );
  AOI21_X1 U19999 ( .B1(n20186), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n16620), .ZN(n16621) );
  OAI211_X1 U20000 ( .C1(n20165), .C2(n16623), .A(n16622), .B(n16621), .ZN(
        n16624) );
  AOI21_X1 U20001 ( .B1(n17183), .B2(n20129), .A(n16624), .ZN(n16625) );
  OAI211_X1 U20002 ( .C1(n20921), .C2(n20190), .A(n16626), .B(n16625), .ZN(
        P2_U2853) );
  NAND2_X1 U20003 ( .A1(n16627), .A2(n20197), .ZN(n16639) );
  NAND2_X1 U20004 ( .A1(n20186), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16633) );
  INV_X1 U20005 ( .A(n16628), .ZN(n16629) );
  AOI22_X1 U20006 ( .A1(n20187), .A2(n16629), .B1(n20126), .B2(
        P2_EBX_REG_1__SCAN_IN), .ZN(n16632) );
  NAND2_X1 U20007 ( .A1(n20934), .A2(n20185), .ZN(n16631) );
  NAND2_X1 U20008 ( .A1(n20150), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n16630) );
  NAND4_X1 U20009 ( .A1(n16633), .A2(n16632), .A3(n16631), .A4(n16630), .ZN(
        n16634) );
  AOI21_X1 U20010 ( .B1(n16635), .B2(n20129), .A(n16634), .ZN(n16638) );
  NAND2_X1 U20011 ( .A1(n20107), .A2(n13336), .ZN(n16637) );
  NAND2_X1 U20012 ( .A1(n20931), .A2(n16645), .ZN(n16636) );
  NAND4_X1 U20013 ( .A1(n16639), .A2(n16638), .A3(n16637), .A4(n16636), .ZN(
        P2_U2854) );
  INV_X1 U20014 ( .A(n16640), .ZN(n16648) );
  OAI21_X1 U20015 ( .B1(n20107), .B2(n20186), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16647) );
  AOI22_X1 U20016 ( .A1(n20187), .A2(n16641), .B1(n20126), .B2(
        P2_EBX_REG_0__SCAN_IN), .ZN(n16643) );
  AOI22_X1 U20017 ( .A1(n20150), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n20185), 
        .B2(n20229), .ZN(n16642) );
  OAI211_X1 U20018 ( .C1(n10780), .C2(n20189), .A(n16643), .B(n16642), .ZN(
        n16644) );
  AOI21_X1 U20019 ( .B1(n20944), .B2(n16645), .A(n16644), .ZN(n16646) );
  OAI211_X1 U20020 ( .C1(n16649), .C2(n16648), .A(n16647), .B(n16646), .ZN(
        P2_U2855) );
  AOI22_X1 U20021 ( .A1(n16662), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16664), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16652) );
  AOI22_X1 U20022 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12330), .B1(
        n16663), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16651) );
  NAND2_X1 U20023 ( .A1(n16652), .A2(n16651), .ZN(n16670) );
  AOI22_X1 U20024 ( .A1(n16658), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16656), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16655) );
  AOI22_X1 U20025 ( .A1(n12329), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16657), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16654) );
  NAND3_X1 U20026 ( .A1(n16655), .A2(n16654), .A3(n16653), .ZN(n16669) );
  AOI22_X1 U20027 ( .A1(n12329), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16656), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16661) );
  AOI22_X1 U20028 ( .A1(n16658), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16657), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16659) );
  NAND3_X1 U20029 ( .A1(n16661), .A2(n16660), .A3(n16659), .ZN(n16668) );
  AOI22_X1 U20030 ( .A1(n16662), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12330), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16666) );
  AOI22_X1 U20031 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n16664), .B1(
        n16663), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16665) );
  NAND2_X1 U20032 ( .A1(n16666), .A2(n16665), .ZN(n16667) );
  OAI22_X1 U20033 ( .A1(n16670), .A2(n16669), .B1(n16668), .B2(n16667), .ZN(
        n16671) );
  XNOR2_X1 U20034 ( .A(n16672), .B(n16671), .ZN(n16775) );
  NOR2_X1 U20035 ( .A1(n16906), .A2(n20204), .ZN(n16673) );
  AOI21_X1 U20036 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n20204), .A(n16673), .ZN(
        n16674) );
  OAI21_X1 U20037 ( .B1(n16775), .B2(n16752), .A(n16674), .ZN(P2_U2857) );
  INV_X1 U20038 ( .A(n16675), .ZN(n16676) );
  NAND3_X1 U20039 ( .A1(n9820), .A2(n16676), .A3(n16757), .ZN(n16678) );
  NAND2_X1 U20040 ( .A1(n20204), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16677) );
  OAI211_X1 U20041 ( .C1(n16916), .C2(n20204), .A(n16678), .B(n16677), .ZN(
        P2_U2858) );
  NAND2_X1 U20042 ( .A1(n12461), .A2(n16679), .ZN(n16680) );
  XOR2_X1 U20043 ( .A(n16681), .B(n16680), .Z(n16782) );
  NOR2_X1 U20044 ( .A1(n16682), .A2(n20204), .ZN(n16683) );
  AOI21_X1 U20045 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n20204), .A(n16683), .ZN(
        n16684) );
  OAI21_X1 U20046 ( .B1(n16782), .B2(n16752), .A(n16684), .ZN(P2_U2859) );
  OAI21_X1 U20047 ( .B1(n16687), .B2(n16686), .A(n16685), .ZN(n16790) );
  NAND2_X1 U20048 ( .A1(n20204), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16690) );
  NAND2_X1 U20049 ( .A1(n16688), .A2(n16760), .ZN(n16689) );
  OAI211_X1 U20050 ( .C1(n16790), .C2(n16752), .A(n16690), .B(n16689), .ZN(
        P2_U2860) );
  NOR2_X1 U20051 ( .A1(n16691), .A2(n16702), .ZN(n16701) );
  NOR2_X1 U20052 ( .A1(n16701), .A2(n16692), .ZN(n16698) );
  NOR2_X1 U20053 ( .A1(n16694), .A2(n16693), .ZN(n16695) );
  XNOR2_X1 U20054 ( .A(n16696), .B(n16695), .ZN(n16697) );
  XNOR2_X1 U20055 ( .A(n16698), .B(n16697), .ZN(n16797) );
  MUX2_X1 U20056 ( .A(n17209), .B(n16699), .S(n20204), .Z(n16700) );
  OAI21_X1 U20057 ( .B1(n16797), .B2(n16752), .A(n16700), .ZN(P2_U2861) );
  AOI21_X1 U20058 ( .B1(n16691), .B2(n16702), .A(n16701), .ZN(n16798) );
  NAND2_X1 U20059 ( .A1(n16798), .A2(n16757), .ZN(n16704) );
  NAND2_X1 U20060 ( .A1(n20204), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n16703) );
  OAI211_X1 U20061 ( .C1(n17223), .C2(n20204), .A(n16704), .B(n16703), .ZN(
        P2_U2862) );
  NOR2_X1 U20062 ( .A1(n16705), .A2(n16706), .ZN(n16810) );
  NOR2_X1 U20063 ( .A1(n16810), .A2(n16752), .ZN(n16708) );
  AOI22_X1 U20064 ( .A1(n16708), .A2(n16707), .B1(P2_EBX_REG_24__SCAN_IN), 
        .B2(n20204), .ZN(n16709) );
  OAI21_X1 U20065 ( .B1(n17235), .B2(n20204), .A(n16709), .ZN(P2_U2863) );
  INV_X1 U20066 ( .A(n16710), .ZN(n16718) );
  NAND2_X1 U20067 ( .A1(n16718), .A2(n16717), .ZN(n16716) );
  XNOR2_X1 U20068 ( .A(n16712), .B(n16711), .ZN(n16713) );
  XNOR2_X1 U20069 ( .A(n16716), .B(n16713), .ZN(n16821) );
  NAND2_X1 U20070 ( .A1(n17240), .A2(n16760), .ZN(n16715) );
  NAND2_X1 U20071 ( .A1(n20204), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n16714) );
  OAI211_X1 U20072 ( .C1(n16821), .C2(n16752), .A(n16715), .B(n16714), .ZN(
        P2_U2864) );
  OAI21_X1 U20073 ( .B1(n16718), .B2(n16717), .A(n16716), .ZN(n16830) );
  AOI21_X1 U20074 ( .B1(n16720), .B2(n14864), .A(n16719), .ZN(n17811) );
  INV_X1 U20075 ( .A(n17811), .ZN(n17259) );
  NOR2_X1 U20076 ( .A1(n17259), .A2(n20204), .ZN(n16721) );
  AOI21_X1 U20077 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n20204), .A(n16721), .ZN(
        n16722) );
  OAI21_X1 U20078 ( .B1(n16752), .B2(n16830), .A(n16722), .ZN(P2_U2865) );
  AND2_X1 U20079 ( .A1(n16723), .A2(n16728), .ZN(n16730) );
  OAI21_X1 U20080 ( .B1(n16730), .B2(n16724), .A(n16710), .ZN(n16839) );
  MUX2_X1 U20081 ( .A(n16726), .B(n16725), .S(n16760), .Z(n16727) );
  OAI21_X1 U20082 ( .B1(n16752), .B2(n16839), .A(n16727), .ZN(P2_U2866) );
  NOR2_X1 U20083 ( .A1(n16723), .A2(n16728), .ZN(n16729) );
  NOR2_X1 U20084 ( .A1(n17271), .A2(n20204), .ZN(n16731) );
  AOI21_X1 U20085 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n20204), .A(n16731), .ZN(
        n16732) );
  OAI21_X1 U20086 ( .B1(n16752), .B2(n16846), .A(n16732), .ZN(P2_U2867) );
  NAND2_X1 U20087 ( .A1(n16733), .A2(n16760), .ZN(n16736) );
  AOI21_X1 U20088 ( .B1(n16734), .B2(n16739), .A(n16723), .ZN(n16847) );
  NAND2_X1 U20089 ( .A1(n16847), .A2(n16757), .ZN(n16735) );
  OAI211_X1 U20090 ( .C1(n20207), .C2(n16737), .A(n16736), .B(n16735), .ZN(
        P2_U2868) );
  INV_X1 U20091 ( .A(n16739), .ZN(n16740) );
  AOI21_X1 U20092 ( .B1(n16741), .B2(n16738), .A(n16740), .ZN(n16856) );
  NAND2_X1 U20093 ( .A1(n16856), .A2(n16757), .ZN(n16743) );
  NAND2_X1 U20094 ( .A1(n20204), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n16742) );
  OAI211_X1 U20095 ( .C1(n17276), .C2(n20204), .A(n16743), .B(n16742), .ZN(
        P2_U2869) );
  OAI21_X1 U20096 ( .B1(n16744), .B2(n16745), .A(n16738), .ZN(n16872) );
  NOR2_X1 U20097 ( .A1(n20084), .A2(n20204), .ZN(n16746) );
  AOI21_X1 U20098 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n20204), .A(n16746), .ZN(
        n16747) );
  OAI21_X1 U20099 ( .B1(n16752), .B2(n16872), .A(n16747), .ZN(P2_U2870) );
  INV_X1 U20100 ( .A(n16744), .ZN(n16748) );
  OAI21_X1 U20101 ( .B1(n9829), .B2(n16749), .A(n16748), .ZN(n16882) );
  INV_X1 U20102 ( .A(n17012), .ZN(n20097) );
  NOR2_X1 U20103 ( .A1(n20097), .A2(n20204), .ZN(n16750) );
  AOI21_X1 U20104 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n20204), .A(n16750), .ZN(
        n16751) );
  OAI21_X1 U20105 ( .B1(n16752), .B2(n16882), .A(n16751), .ZN(P2_U2871) );
  INV_X1 U20106 ( .A(n16753), .ZN(n16754) );
  AOI21_X1 U20107 ( .B1(n16756), .B2(n16755), .A(n16754), .ZN(n20110) );
  OAI21_X1 U20108 ( .B1(n16759), .B2(n16758), .A(n16757), .ZN(n16761) );
  INV_X1 U20109 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n20104) );
  OAI22_X1 U20110 ( .A1(n16761), .A2(n9829), .B1(n16760), .B2(n20104), .ZN(
        n16762) );
  AOI21_X1 U20111 ( .B1(n20110), .B2(n20207), .A(n16762), .ZN(n16763) );
  INV_X1 U20112 ( .A(n16763), .ZN(P2_U2872) );
  INV_X1 U20113 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n16767) );
  NAND2_X1 U20114 ( .A1(n16764), .A2(n12194), .ZN(n16766) );
  AOI22_X1 U20115 ( .A1(n16873), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n20226), .ZN(n16765) );
  OAI211_X1 U20116 ( .C1(n16878), .C2(n16767), .A(n16766), .B(n16765), .ZN(
        P2_U2888) );
  INV_X1 U20117 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n16771) );
  NAND2_X1 U20118 ( .A1(n16873), .A2(BUF1_REG_30__SCAN_IN), .ZN(n16770) );
  AOI22_X1 U20119 ( .A1(n16875), .A2(n16768), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n20226), .ZN(n16769) );
  OAI211_X1 U20120 ( .C1(n16878), .C2(n16771), .A(n16770), .B(n16769), .ZN(
        n16772) );
  AOI21_X1 U20121 ( .B1(n16773), .B2(n12194), .A(n16772), .ZN(n16774) );
  OAI21_X1 U20122 ( .B1(n16775), .B2(n16883), .A(n16774), .ZN(P2_U2889) );
  INV_X1 U20123 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n16778) );
  NAND2_X1 U20124 ( .A1(n16873), .A2(BUF1_REG_28__SCAN_IN), .ZN(n16777) );
  AOI22_X1 U20125 ( .A1(n16875), .A2(n20278), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n20226), .ZN(n16776) );
  OAI211_X1 U20126 ( .C1(n16778), .C2(n16878), .A(n16777), .B(n16776), .ZN(
        n16779) );
  AOI21_X1 U20127 ( .B1(n16780), .B2(n12194), .A(n16779), .ZN(n16781) );
  OAI21_X1 U20128 ( .B1(n16782), .B2(n16883), .A(n16781), .ZN(P2_U2891) );
  INV_X1 U20129 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n16786) );
  NAND2_X1 U20130 ( .A1(n16873), .A2(BUF1_REG_27__SCAN_IN), .ZN(n16785) );
  AOI22_X1 U20131 ( .A1(n16875), .A2(n16783), .B1(P2_EAX_REG_27__SCAN_IN), 
        .B2(n20226), .ZN(n16784) );
  OAI211_X1 U20132 ( .C1(n16878), .C2(n16786), .A(n16785), .B(n16784), .ZN(
        n16787) );
  AOI21_X1 U20133 ( .B1(n16788), .B2(n12194), .A(n16787), .ZN(n16789) );
  OAI21_X1 U20134 ( .B1(n16790), .B2(n16883), .A(n16789), .ZN(P2_U2892) );
  INV_X1 U20135 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n16793) );
  AOI22_X1 U20136 ( .A1(n16875), .A2(n16791), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n20226), .ZN(n16792) );
  OAI21_X1 U20137 ( .B1(n16878), .B2(n16793), .A(n16792), .ZN(n16795) );
  NOR2_X1 U20138 ( .A1(n17208), .A2(n12497), .ZN(n16794) );
  AOI211_X1 U20139 ( .C1(n16873), .C2(BUF1_REG_26__SCAN_IN), .A(n16795), .B(
        n16794), .ZN(n16796) );
  OAI21_X1 U20140 ( .B1(n16797), .B2(n16883), .A(n16796), .ZN(P2_U2893) );
  INV_X1 U20141 ( .A(n17225), .ZN(n16804) );
  NAND2_X1 U20142 ( .A1(n16798), .A2(n20227), .ZN(n16803) );
  AOI22_X1 U20143 ( .A1(n16875), .A2(n16799), .B1(P2_EAX_REG_25__SCAN_IN), 
        .B2(n20226), .ZN(n16800) );
  OAI21_X1 U20144 ( .B1(n16878), .B2(n18018), .A(n16800), .ZN(n16801) );
  AOI21_X1 U20145 ( .B1(n16873), .B2(BUF1_REG_25__SCAN_IN), .A(n16801), .ZN(
        n16802) );
  OAI211_X1 U20146 ( .C1(n16804), .C2(n12497), .A(n16803), .B(n16802), .ZN(
        P2_U2894) );
  INV_X1 U20147 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n16807) );
  AOI22_X1 U20148 ( .A1(n16875), .A2(n16805), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n20226), .ZN(n16806) );
  OAI21_X1 U20149 ( .B1(n16878), .B2(n16807), .A(n16806), .ZN(n16809) );
  NOR2_X1 U20150 ( .A1(n17234), .A2(n12497), .ZN(n16808) );
  AOI211_X1 U20151 ( .C1(BUF1_REG_24__SCAN_IN), .C2(n16873), .A(n16809), .B(
        n16808), .ZN(n16813) );
  INV_X1 U20152 ( .A(n16810), .ZN(n16811) );
  NAND3_X1 U20153 ( .A1(n16811), .A2(n20227), .A3(n16707), .ZN(n16812) );
  NAND2_X1 U20154 ( .A1(n16813), .A2(n16812), .ZN(P2_U2895) );
  INV_X1 U20155 ( .A(n17248), .ZN(n16819) );
  INV_X1 U20156 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n16817) );
  NAND2_X1 U20157 ( .A1(n16873), .A2(BUF1_REG_23__SCAN_IN), .ZN(n16816) );
  AOI22_X1 U20158 ( .A1(n16875), .A2(n16814), .B1(P2_EAX_REG_23__SCAN_IN), 
        .B2(n20226), .ZN(n16815) );
  OAI211_X1 U20159 ( .C1(n16817), .C2(n16878), .A(n16816), .B(n16815), .ZN(
        n16818) );
  AOI21_X1 U20160 ( .B1(n16819), .B2(n12194), .A(n16818), .ZN(n16820) );
  OAI21_X1 U20161 ( .B1(n16821), .B2(n16883), .A(n16820), .ZN(P2_U2896) );
  AOI21_X1 U20162 ( .B1(n16823), .B2(n14870), .A(n16470), .ZN(n17810) );
  INV_X1 U20163 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n16827) );
  NAND2_X1 U20164 ( .A1(n16873), .A2(BUF1_REG_22__SCAN_IN), .ZN(n16826) );
  AOI22_X1 U20165 ( .A1(n16875), .A2(n16824), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n20226), .ZN(n16825) );
  OAI211_X1 U20166 ( .C1(n16827), .C2(n16878), .A(n16826), .B(n16825), .ZN(
        n16828) );
  AOI21_X1 U20167 ( .B1(n17810), .B2(n12194), .A(n16828), .ZN(n16829) );
  OAI21_X1 U20168 ( .B1(n16883), .B2(n16830), .A(n16829), .ZN(P2_U2897) );
  INV_X1 U20169 ( .A(n16831), .ZN(n16837) );
  INV_X1 U20170 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n16835) );
  NAND2_X1 U20171 ( .A1(n16873), .A2(BUF1_REG_21__SCAN_IN), .ZN(n16834) );
  AOI22_X1 U20172 ( .A1(n16875), .A2(n16832), .B1(P2_EAX_REG_21__SCAN_IN), 
        .B2(n20226), .ZN(n16833) );
  OAI211_X1 U20173 ( .C1(n16835), .C2(n16878), .A(n16834), .B(n16833), .ZN(
        n16836) );
  AOI21_X1 U20174 ( .B1(n16837), .B2(n12194), .A(n16836), .ZN(n16838) );
  OAI21_X1 U20175 ( .B1(n16883), .B2(n16839), .A(n16838), .ZN(P2_U2898) );
  INV_X1 U20176 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n16843) );
  NAND2_X1 U20177 ( .A1(n16873), .A2(BUF1_REG_20__SCAN_IN), .ZN(n16842) );
  AOI22_X1 U20178 ( .A1(n16875), .A2(n16840), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n20226), .ZN(n16841) );
  OAI211_X1 U20179 ( .C1(n16843), .C2(n16878), .A(n16842), .B(n16841), .ZN(
        n16844) );
  AOI21_X1 U20180 ( .B1(n17268), .B2(n12194), .A(n16844), .ZN(n16845) );
  OAI21_X1 U20181 ( .B1(n16883), .B2(n16846), .A(n16845), .ZN(P2_U2899) );
  NAND2_X1 U20182 ( .A1(n16847), .A2(n20227), .ZN(n16854) );
  NOR2_X1 U20183 ( .A1(n16878), .A2(n16848), .ZN(n16852) );
  OAI22_X1 U20184 ( .A1(n16850), .A2(n20302), .B1(n16897), .B2(n16849), .ZN(
        n16851) );
  AOI211_X1 U20185 ( .C1(BUF1_REG_19__SCAN_IN), .C2(n16873), .A(n16852), .B(
        n16851), .ZN(n16853) );
  OAI211_X1 U20186 ( .C1(n12497), .C2(n16855), .A(n16854), .B(n16853), .ZN(
        P2_U2900) );
  INV_X1 U20187 ( .A(n16856), .ZN(n16864) );
  INV_X1 U20188 ( .A(n17283), .ZN(n16862) );
  INV_X1 U20189 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n16860) );
  NAND2_X1 U20190 ( .A1(n16873), .A2(BUF1_REG_18__SCAN_IN), .ZN(n16859) );
  AOI22_X1 U20191 ( .A1(n16875), .A2(n16857), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n20226), .ZN(n16858) );
  OAI211_X1 U20192 ( .C1(n16860), .C2(n16878), .A(n16859), .B(n16858), .ZN(
        n16861) );
  AOI21_X1 U20193 ( .B1(n16862), .B2(n12194), .A(n16861), .ZN(n16863) );
  OAI21_X1 U20194 ( .B1(n16864), .B2(n16883), .A(n16863), .ZN(P2_U2901) );
  INV_X1 U20195 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n16868) );
  NAND2_X1 U20196 ( .A1(n16873), .A2(BUF1_REG_17__SCAN_IN), .ZN(n16867) );
  AOI22_X1 U20197 ( .A1(n16875), .A2(n16865), .B1(P2_EAX_REG_17__SCAN_IN), 
        .B2(n20226), .ZN(n16866) );
  OAI211_X1 U20198 ( .C1(n16868), .C2(n16878), .A(n16867), .B(n16866), .ZN(
        n16869) );
  AOI21_X1 U20199 ( .B1(n16870), .B2(n12194), .A(n16869), .ZN(n16871) );
  OAI21_X1 U20200 ( .B1(n16883), .B2(n16872), .A(n16871), .ZN(P2_U2902) );
  INV_X1 U20201 ( .A(n20096), .ZN(n16880) );
  NAND2_X1 U20202 ( .A1(n16873), .A2(BUF1_REG_16__SCAN_IN), .ZN(n16877) );
  AOI22_X1 U20203 ( .A1(n16875), .A2(n16874), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n20226), .ZN(n16876) );
  OAI211_X1 U20204 ( .C1(n19416), .C2(n16878), .A(n16877), .B(n16876), .ZN(
        n16879) );
  AOI21_X1 U20205 ( .B1(n16880), .B2(n12194), .A(n16879), .ZN(n16881) );
  OAI21_X1 U20206 ( .B1(n16883), .B2(n16882), .A(n16881), .ZN(P2_U2903) );
  INV_X1 U20207 ( .A(n17443), .ZN(n20917) );
  INV_X1 U20208 ( .A(n20324), .ZN(n20918) );
  XOR2_X1 U20209 ( .A(n17443), .B(n20324), .Z(n20216) );
  INV_X1 U20210 ( .A(n20921), .ZN(n16885) );
  OAI21_X1 U20211 ( .B1(n16885), .B2(n20923), .A(n16884), .ZN(n20215) );
  NAND2_X1 U20212 ( .A1(n20216), .A2(n20215), .ZN(n20214) );
  OAI21_X1 U20213 ( .B1(n20917), .B2(n20918), .A(n20214), .ZN(n16888) );
  NAND2_X1 U20214 ( .A1(n16597), .A2(n16886), .ZN(n16887) );
  NAND2_X1 U20215 ( .A1(n14777), .A2(n16887), .ZN(n20179) );
  NAND2_X1 U20216 ( .A1(n16888), .A2(n20179), .ZN(n20210) );
  INV_X1 U20217 ( .A(n16890), .ZN(n16891) );
  NAND3_X1 U20218 ( .A1(n16889), .A2(n16892), .A3(n16891), .ZN(n16893) );
  NAND2_X1 U20219 ( .A1(n16894), .A2(n16893), .ZN(n20209) );
  INV_X1 U20220 ( .A(n20209), .ZN(n16895) );
  NAND3_X1 U20221 ( .A1(n20210), .A2(n20227), .A3(n16895), .ZN(n16901) );
  INV_X1 U20222 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n16896) );
  OAI22_X1 U20223 ( .A1(n20232), .A2(n20308), .B1(n16897), .B2(n16896), .ZN(
        n16898) );
  AOI21_X1 U20224 ( .B1(n17419), .B2(n16899), .A(n16898), .ZN(n16900) );
  NAND2_X1 U20225 ( .A1(n16901), .A2(n16900), .ZN(P2_U2914) );
  OAI21_X1 U20226 ( .B1(n17187), .B2(n10327), .A(n16902), .ZN(n16903) );
  AOI21_X1 U20227 ( .B1(n16904), .B2(n17190), .A(n16903), .ZN(n16905) );
  OAI21_X1 U20228 ( .B1(n16906), .B2(n17166), .A(n16905), .ZN(n16907) );
  OAI21_X1 U20229 ( .B1(n16910), .B2(n17181), .A(n16909), .ZN(P2_U2984) );
  OAI21_X1 U20230 ( .B1(n17187), .B2(n16912), .A(n16911), .ZN(n16913) );
  AOI21_X1 U20231 ( .B1(n16914), .B2(n17190), .A(n16913), .ZN(n16915) );
  OAI21_X1 U20232 ( .B1(n16916), .B2(n17166), .A(n16915), .ZN(n16917) );
  OAI21_X1 U20233 ( .B1(n16919), .B2(n17181), .A(n16918), .ZN(P2_U2985) );
  XOR2_X1 U20234 ( .A(n16921), .B(n16920), .Z(n17214) );
  INV_X1 U20235 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17203) );
  NAND2_X1 U20236 ( .A1(n16948), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16928) );
  AOI21_X1 U20237 ( .B1(n17203), .B2(n16928), .A(n16922), .ZN(n17212) );
  NOR2_X1 U20238 ( .A1(n17149), .A2(n20891), .ZN(n17204) );
  AOI21_X1 U20239 ( .B1(n17172), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n17204), .ZN(n16923) );
  OAI21_X1 U20240 ( .B1(n16924), .B2(n17175), .A(n16923), .ZN(n16926) );
  NOR2_X1 U20241 ( .A1(n17209), .A2(n17166), .ZN(n16925) );
  AOI211_X1 U20242 ( .C1(n17212), .C2(n17196), .A(n16926), .B(n16925), .ZN(
        n16927) );
  OAI21_X1 U20243 ( .B1(n17214), .B2(n17181), .A(n16927), .ZN(P2_U2988) );
  OAI21_X1 U20244 ( .B1(n16948), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n16928), .ZN(n17228) );
  INV_X1 U20245 ( .A(n16929), .ZN(n16938) );
  INV_X1 U20246 ( .A(n16931), .ZN(n16932) );
  NAND2_X1 U20247 ( .A1(n16930), .A2(n16932), .ZN(n16947) );
  INV_X1 U20248 ( .A(n16945), .ZN(n16934) );
  OAI22_X1 U20249 ( .A1(n16947), .A2(n16933), .B1(n16934), .B2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16936) );
  OAI21_X1 U20250 ( .B1(n16934), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n16937), .ZN(n16935) );
  AOI22_X1 U20251 ( .A1(n16938), .A2(n16937), .B1(n16936), .B2(n16935), .ZN(
        n17215) );
  NAND2_X1 U20252 ( .A1(n17215), .A2(n17193), .ZN(n16944) );
  NOR2_X1 U20253 ( .A1(n17149), .A2(n20889), .ZN(n17217) );
  INV_X1 U20254 ( .A(n17217), .ZN(n16939) );
  OAI21_X1 U20255 ( .B1(n17187), .B2(n10354), .A(n16939), .ZN(n16941) );
  NOR2_X1 U20256 ( .A1(n17223), .A2(n17166), .ZN(n16940) );
  AOI211_X1 U20257 ( .C1(n17190), .C2(n16942), .A(n16941), .B(n16940), .ZN(
        n16943) );
  OAI211_X1 U20258 ( .C1(n17139), .C2(n17228), .A(n16944), .B(n16943), .ZN(
        P2_U2989) );
  XNOR2_X1 U20259 ( .A(n16945), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16946) );
  XNOR2_X1 U20260 ( .A(n16947), .B(n16946), .ZN(n17239) );
  NOR2_X1 U20261 ( .A1(n17149), .A2(n16950), .ZN(n17229) );
  NOR2_X1 U20262 ( .A1(n16951), .A2(n17175), .ZN(n16952) );
  AOI211_X1 U20263 ( .C1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n17172), .A(
        n17229), .B(n16952), .ZN(n16953) );
  OAI21_X1 U20264 ( .B1(n17235), .B2(n17166), .A(n16953), .ZN(n16954) );
  OAI21_X1 U20265 ( .B1(n17239), .B2(n17181), .A(n16955), .ZN(P2_U2990) );
  OAI21_X1 U20266 ( .B1(n16965), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16956), .ZN(n17252) );
  XOR2_X1 U20267 ( .A(n16959), .B(n16958), .Z(n17250) );
  NAND2_X1 U20268 ( .A1(n17240), .A2(n17182), .ZN(n16961) );
  NOR2_X1 U20269 ( .A1(n17149), .A2(n20886), .ZN(n17245) );
  AOI21_X1 U20270 ( .B1(n17172), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n17245), .ZN(n16960) );
  OAI211_X1 U20271 ( .C1(n17175), .C2(n16962), .A(n16961), .B(n16960), .ZN(
        n16963) );
  AOI21_X1 U20272 ( .B1(n17250), .B2(n17193), .A(n16963), .ZN(n16964) );
  OAI21_X1 U20273 ( .B1(n17139), .B2(n17252), .A(n16964), .ZN(P2_U2991) );
  OAI21_X1 U20274 ( .B1(n16966), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n10112), .ZN(n17263) );
  NAND2_X1 U20275 ( .A1(n17811), .A2(n17182), .ZN(n16970) );
  NOR2_X1 U20276 ( .A1(n17149), .A2(n16968), .ZN(n17257) );
  AOI21_X1 U20277 ( .B1(n17172), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n17257), .ZN(n16969) );
  OAI211_X1 U20278 ( .C1(n17815), .C2(n17175), .A(n16970), .B(n16969), .ZN(
        n16971) );
  AOI21_X1 U20279 ( .B1(n17261), .B2(n17193), .A(n16971), .ZN(n16972) );
  OAI21_X1 U20280 ( .B1(n17139), .B2(n17263), .A(n16972), .ZN(P2_U2992) );
  INV_X1 U20281 ( .A(n16973), .ZN(n16974) );
  NOR2_X1 U20282 ( .A1(n9825), .A2(n16976), .ZN(n16977) );
  AOI21_X1 U20283 ( .B1(n16981), .B2(n16980), .A(n16979), .ZN(n17273) );
  NOR2_X1 U20284 ( .A1(n17149), .A2(n16982), .ZN(n17267) );
  NOR2_X1 U20285 ( .A1(n16983), .A2(n17175), .ZN(n16984) );
  AOI211_X1 U20286 ( .C1(n17172), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n17267), .B(n16984), .ZN(n16985) );
  OAI21_X1 U20287 ( .B1(n17271), .B2(n17166), .A(n16985), .ZN(n16986) );
  AOI21_X1 U20288 ( .B1(n17273), .B2(n17196), .A(n16986), .ZN(n16987) );
  OAI21_X1 U20289 ( .B1(n17275), .B2(n17181), .A(n16987), .ZN(P2_U2994) );
  NOR2_X1 U20290 ( .A1(n16989), .A2(n16988), .ZN(n16990) );
  XNOR2_X1 U20291 ( .A(n14823), .B(n16990), .ZN(n17288) );
  AOI21_X1 U20292 ( .B1(n17277), .B2(n17002), .A(n16991), .ZN(n17286) );
  NOR2_X1 U20293 ( .A1(n17149), .A2(n16992), .ZN(n17280) );
  NOR2_X1 U20294 ( .A1(n16993), .A2(n17175), .ZN(n16994) );
  AOI211_X1 U20295 ( .C1(n17172), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17280), .B(n16994), .ZN(n16995) );
  OAI21_X1 U20296 ( .B1(n17276), .B2(n17166), .A(n16995), .ZN(n16996) );
  AOI21_X1 U20297 ( .B1(n17286), .B2(n17196), .A(n16996), .ZN(n16997) );
  OAI21_X1 U20298 ( .B1(n17288), .B2(n17181), .A(n16997), .ZN(P2_U2996) );
  INV_X1 U20299 ( .A(n20084), .ZN(n17001) );
  AOI21_X1 U20300 ( .B1(n17172), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16998), .ZN(n16999) );
  OAI21_X1 U20301 ( .B1(n17175), .B2(n20078), .A(n16999), .ZN(n17000) );
  AOI21_X1 U20302 ( .B1(n17001), .B2(n17182), .A(n17000), .ZN(n17005) );
  OAI211_X1 U20303 ( .C1(n17003), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n17002), .B(n17196), .ZN(n17004) );
  OAI211_X1 U20304 ( .C1(n17006), .C2(n17181), .A(n17005), .B(n17004), .ZN(
        P2_U2997) );
  XNOR2_X1 U20305 ( .A(n17021), .B(n17007), .ZN(n17015) );
  NAND2_X1 U20306 ( .A1(n17008), .A2(n17193), .ZN(n17014) );
  NAND2_X1 U20307 ( .A1(n17172), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17009) );
  OAI211_X1 U20308 ( .C1(n17175), .C2(n20095), .A(n17010), .B(n17009), .ZN(
        n17011) );
  AOI21_X1 U20309 ( .B1(n17012), .B2(n17182), .A(n17011), .ZN(n17013) );
  OAI211_X1 U20310 ( .C1(n17139), .C2(n17015), .A(n17014), .B(n17013), .ZN(
        P2_U2998) );
  NAND2_X1 U20311 ( .A1(n17017), .A2(n17016), .ZN(n17018) );
  NAND2_X1 U20312 ( .A1(n17190), .A2(n20112), .ZN(n17019) );
  OR2_X1 U20313 ( .A1(n17149), .A2(n20873), .ZN(n17289) );
  OAI211_X1 U20314 ( .C1(n17187), .C2(n17020), .A(n17019), .B(n17289), .ZN(
        n17023) );
  NOR2_X1 U20315 ( .A1(n17295), .A2(n17139), .ZN(n17022) );
  AOI211_X1 U20316 ( .C1(n17182), .C2(n20110), .A(n17023), .B(n17022), .ZN(
        n17024) );
  OAI21_X1 U20317 ( .B1(n17299), .B2(n17181), .A(n17024), .ZN(P2_U2999) );
  NAND2_X1 U20318 ( .A1(n17027), .A2(n17026), .ZN(n17028) );
  XNOR2_X1 U20319 ( .A(n17025), .B(n17028), .ZN(n17314) );
  INV_X1 U20320 ( .A(n20181), .ZN(n17089) );
  NAND2_X1 U20321 ( .A1(n17089), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n17307) );
  OAI21_X1 U20322 ( .B1(n17187), .B2(n17029), .A(n17307), .ZN(n17031) );
  NOR2_X1 U20323 ( .A1(n20127), .A2(n17166), .ZN(n17030) );
  AOI211_X1 U20324 ( .C1(n17190), .C2(n20120), .A(n17031), .B(n17030), .ZN(
        n17035) );
  NAND2_X1 U20325 ( .A1(n17056), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17036) );
  AOI21_X1 U20326 ( .B1(n17036), .B2(n17308), .A(n17033), .ZN(n17311) );
  NAND2_X1 U20327 ( .A1(n17311), .A2(n17196), .ZN(n17034) );
  OAI211_X1 U20328 ( .C1(n17314), .C2(n17181), .A(n17035), .B(n17034), .ZN(
        P2_U3000) );
  OAI21_X1 U20329 ( .B1(n17056), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n17036), .ZN(n17327) );
  NAND2_X1 U20330 ( .A1(n10440), .A2(n17039), .ZN(n17040) );
  XNOR2_X1 U20331 ( .A(n17037), .B(n17040), .ZN(n17325) );
  NOR2_X1 U20332 ( .A1(n20181), .A2(n20869), .ZN(n17320) );
  NOR2_X1 U20333 ( .A1(n17175), .A2(n17041), .ZN(n17042) );
  AOI211_X1 U20334 ( .C1(n17172), .C2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n17320), .B(n17042), .ZN(n17043) );
  OAI21_X1 U20335 ( .B1(n17323), .B2(n17166), .A(n17043), .ZN(n17044) );
  AOI21_X1 U20336 ( .B1(n17325), .B2(n17193), .A(n17044), .ZN(n17045) );
  OAI21_X1 U20337 ( .B1(n17327), .B2(n17139), .A(n17045), .ZN(P2_U3001) );
  INV_X1 U20338 ( .A(n17046), .ZN(n17049) );
  INV_X1 U20339 ( .A(n17047), .ZN(n17048) );
  AOI21_X1 U20340 ( .B1(n17064), .B2(n17065), .A(n17050), .ZN(n17055) );
  INV_X1 U20341 ( .A(n17051), .ZN(n17053) );
  NAND2_X1 U20342 ( .A1(n17053), .A2(n17052), .ZN(n17054) );
  XNOR2_X1 U20343 ( .A(n17055), .B(n17054), .ZN(n17342) );
  NOR2_X1 U20344 ( .A1(n20181), .A2(n20867), .ZN(n17328) );
  NOR2_X1 U20345 ( .A1(n17175), .A2(n17057), .ZN(n17058) );
  AOI211_X1 U20346 ( .C1(n17172), .C2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n17328), .B(n17058), .ZN(n17059) );
  OAI21_X1 U20347 ( .B1(n17338), .B2(n17166), .A(n17059), .ZN(n17060) );
  AOI21_X1 U20348 ( .B1(n17340), .B2(n17196), .A(n17060), .ZN(n17061) );
  OAI21_X1 U20349 ( .B1(n17342), .B2(n17181), .A(n17061), .ZN(P2_U3002) );
  INV_X1 U20350 ( .A(n17062), .ZN(n17063) );
  NOR2_X1 U20351 ( .A1(n17064), .A2(n17063), .ZN(n17068) );
  NAND2_X1 U20352 ( .A1(n17066), .A2(n17065), .ZN(n17067) );
  XNOR2_X1 U20353 ( .A(n17068), .B(n17067), .ZN(n17356) );
  NAND2_X1 U20354 ( .A1(n17190), .A2(n17069), .ZN(n17070) );
  NAND2_X1 U20355 ( .A1(n17089), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n17346) );
  OAI211_X1 U20356 ( .C1(n17187), .C2(n17071), .A(n17070), .B(n17346), .ZN(
        n17072) );
  AOI21_X1 U20357 ( .B1(n17352), .B2(n17182), .A(n17072), .ZN(n17076) );
  NAND2_X1 U20358 ( .A1(n17099), .A2(n17073), .ZN(n17078) );
  AOI21_X1 U20359 ( .B1(n17349), .B2(n17078), .A(n17074), .ZN(n17353) );
  NAND2_X1 U20360 ( .A1(n17353), .A2(n17196), .ZN(n17075) );
  OAI211_X1 U20361 ( .C1(n17356), .C2(n17181), .A(n17076), .B(n17075), .ZN(
        P2_U3003) );
  INV_X1 U20362 ( .A(n17099), .ZN(n17077) );
  OAI21_X1 U20363 ( .B1(n17077), .B2(n17348), .A(n17361), .ZN(n17079) );
  NAND2_X1 U20364 ( .A1(n17079), .A2(n17078), .ZN(n17369) );
  INV_X1 U20365 ( .A(n17081), .ZN(n17083) );
  OAI21_X1 U20366 ( .B1(n17125), .B2(n17083), .A(n17082), .ZN(n17098) );
  INV_X1 U20367 ( .A(n17095), .ZN(n17084) );
  OAI21_X1 U20368 ( .B1(n17098), .B2(n17084), .A(n17096), .ZN(n17088) );
  NAND2_X1 U20369 ( .A1(n17086), .A2(n17085), .ZN(n17087) );
  XNOR2_X1 U20370 ( .A(n17088), .B(n17087), .ZN(n17357) );
  NAND2_X1 U20371 ( .A1(n17357), .A2(n17193), .ZN(n17094) );
  NAND2_X1 U20372 ( .A1(n17089), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n17360) );
  OAI21_X1 U20373 ( .B1(n17187), .B2(n17090), .A(n17360), .ZN(n17092) );
  NOR2_X1 U20374 ( .A1(n20140), .A2(n17166), .ZN(n17091) );
  AOI211_X1 U20375 ( .C1(n17190), .C2(n20137), .A(n17092), .B(n17091), .ZN(
        n17093) );
  OAI211_X1 U20376 ( .C1(n17139), .C2(n17369), .A(n17094), .B(n17093), .ZN(
        P2_U3004) );
  NAND2_X1 U20377 ( .A1(n17096), .A2(n17095), .ZN(n17097) );
  XNOR2_X1 U20378 ( .A(n17098), .B(n17097), .ZN(n17379) );
  NOR2_X1 U20379 ( .A1(n20181), .A2(n20861), .ZN(n17372) );
  NOR2_X1 U20380 ( .A1(n17175), .A2(n20149), .ZN(n17100) );
  AOI211_X1 U20381 ( .C1(n17172), .C2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17372), .B(n17100), .ZN(n17101) );
  OAI21_X1 U20382 ( .B1(n20155), .B2(n17166), .A(n17101), .ZN(n17102) );
  AOI21_X1 U20383 ( .B1(n17376), .B2(n17196), .A(n17102), .ZN(n17103) );
  OAI21_X1 U20384 ( .B1(n17379), .B2(n17181), .A(n17103), .ZN(P2_U3005) );
  XNOR2_X1 U20385 ( .A(n17107), .B(n17105), .ZN(n17121) );
  AOI22_X1 U20386 ( .A1(n17121), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B1(
        n17107), .B2(n17106), .ZN(n17108) );
  XOR2_X1 U20387 ( .A(n17109), .B(n17108), .Z(n17391) );
  NAND2_X1 U20388 ( .A1(n17111), .A2(n17110), .ZN(n17114) );
  INV_X1 U20389 ( .A(n17123), .ZN(n17112) );
  AOI21_X1 U20390 ( .B1(n17125), .B2(n17122), .A(n17112), .ZN(n17113) );
  XOR2_X1 U20391 ( .A(n17114), .B(n17113), .Z(n17389) );
  NOR2_X1 U20392 ( .A1(n20181), .A2(n17115), .ZN(n17382) );
  AOI21_X1 U20393 ( .B1(n17172), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17382), .ZN(n17118) );
  NAND2_X1 U20394 ( .A1(n17190), .A2(n17116), .ZN(n17117) );
  OAI211_X1 U20395 ( .C1(n17386), .C2(n17166), .A(n17118), .B(n17117), .ZN(
        n17119) );
  AOI21_X1 U20396 ( .B1(n17389), .B2(n17193), .A(n17119), .ZN(n17120) );
  OAI21_X1 U20397 ( .B1(n17391), .B2(n17139), .A(n17120), .ZN(P2_U3006) );
  XNOR2_X1 U20398 ( .A(n17121), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17402) );
  NAND2_X1 U20399 ( .A1(n17123), .A2(n17122), .ZN(n17124) );
  XNOR2_X1 U20400 ( .A(n17125), .B(n17124), .ZN(n17400) );
  NAND2_X1 U20401 ( .A1(n20167), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n17392) );
  OAI21_X1 U20402 ( .B1(n17187), .B2(n17126), .A(n17392), .ZN(n17127) );
  AOI21_X1 U20403 ( .B1(n17190), .B2(n20161), .A(n17127), .ZN(n17128) );
  OAI21_X1 U20404 ( .B1(n20173), .B2(n17166), .A(n17128), .ZN(n17129) );
  AOI21_X1 U20405 ( .B1(n17400), .B2(n17193), .A(n17129), .ZN(n17130) );
  OAI21_X1 U20406 ( .B1(n17139), .B2(n17402), .A(n17130), .ZN(P2_U3007) );
  XNOR2_X1 U20407 ( .A(n17131), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17416) );
  XOR2_X1 U20408 ( .A(n17132), .B(n17133), .Z(n17413) );
  NOR2_X1 U20409 ( .A1(n17409), .A2(n17166), .ZN(n17137) );
  AOI22_X1 U20410 ( .A1(n17172), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n20167), .ZN(n17134) );
  OAI21_X1 U20411 ( .B1(n17175), .B2(n17135), .A(n17134), .ZN(n17136) );
  AOI211_X1 U20412 ( .C1(n17413), .C2(n17193), .A(n17137), .B(n17136), .ZN(
        n17138) );
  OAI21_X1 U20413 ( .B1(n17416), .B2(n17139), .A(n17138), .ZN(P2_U3008) );
  XNOR2_X1 U20414 ( .A(n17141), .B(n17140), .ZN(n17428) );
  INV_X1 U20415 ( .A(n17142), .ZN(n17147) );
  AOI21_X1 U20416 ( .B1(n17146), .B2(n17144), .A(n17143), .ZN(n17145) );
  AOI21_X1 U20417 ( .B1(n17147), .B2(n17146), .A(n17145), .ZN(n17426) );
  NOR2_X1 U20418 ( .A1(n17149), .A2(n17148), .ZN(n17418) );
  AOI21_X1 U20419 ( .B1(n17172), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n17418), .ZN(n17152) );
  NAND2_X1 U20420 ( .A1(n17190), .A2(n17150), .ZN(n17151) );
  OAI211_X1 U20421 ( .C1(n17153), .C2(n17166), .A(n17152), .B(n17151), .ZN(
        n17154) );
  AOI21_X1 U20422 ( .B1(n17426), .B2(n17196), .A(n17154), .ZN(n17155) );
  OAI21_X1 U20423 ( .B1(n17428), .B2(n17181), .A(n17155), .ZN(P2_U3009) );
  XNOR2_X1 U20424 ( .A(n17156), .B(n17157), .ZN(n17438) );
  XNOR2_X1 U20425 ( .A(n17158), .B(n17432), .ZN(n17159) );
  XNOR2_X1 U20426 ( .A(n17160), .B(n17159), .ZN(n17436) );
  NAND2_X1 U20427 ( .A1(n17162), .A2(n17161), .ZN(n17163) );
  NAND2_X1 U20428 ( .A1(n14609), .A2(n17163), .ZN(n20203) );
  AOI22_X1 U20429 ( .A1(n17172), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n20167), .ZN(n17165) );
  NAND2_X1 U20430 ( .A1(n17190), .A2(n20195), .ZN(n17164) );
  OAI211_X1 U20431 ( .C1(n20203), .C2(n17166), .A(n17165), .B(n17164), .ZN(
        n17167) );
  AOI21_X1 U20432 ( .B1(n17436), .B2(n17196), .A(n17167), .ZN(n17168) );
  OAI21_X1 U20433 ( .B1(n17438), .B2(n17181), .A(n17168), .ZN(P2_U3010) );
  NAND2_X1 U20434 ( .A1(n9799), .A2(n17169), .ZN(n17171) );
  XNOR2_X1 U20435 ( .A(n17171), .B(n17170), .ZN(n17450) );
  AOI22_X1 U20436 ( .A1(n17172), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_REIP_REG_3__SCAN_IN), .B2(n20167), .ZN(n17173) );
  OAI21_X1 U20437 ( .B1(n17175), .B2(n17174), .A(n17173), .ZN(n17176) );
  AOI21_X1 U20438 ( .B1(n17446), .B2(n17182), .A(n17176), .ZN(n17180) );
  NAND2_X1 U20439 ( .A1(n9918), .A2(n17178), .ZN(n17447) );
  NAND3_X1 U20440 ( .A1(n17177), .A2(n17447), .A3(n17196), .ZN(n17179) );
  OAI211_X1 U20441 ( .C1(n17450), .C2(n17181), .A(n17180), .B(n17179), .ZN(
        P2_U3011) );
  NAND2_X1 U20442 ( .A1(n17183), .A2(n17182), .ZN(n17201) );
  INV_X1 U20443 ( .A(n17184), .ZN(n17189) );
  INV_X1 U20444 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17186) );
  OAI21_X1 U20445 ( .B1(n17187), .B2(n17186), .A(n17185), .ZN(n17188) );
  AOI21_X1 U20446 ( .B1(n17190), .B2(n17189), .A(n17188), .ZN(n17200) );
  INV_X1 U20447 ( .A(n17191), .ZN(n17194) );
  NAND3_X1 U20448 ( .A1(n17194), .A2(n17193), .A3(n17192), .ZN(n17199) );
  NAND3_X1 U20449 ( .A1(n17197), .A2(n17196), .A3(n17195), .ZN(n17198) );
  NAND4_X1 U20450 ( .A1(n17201), .A2(n17200), .A3(n17199), .A4(n17198), .ZN(
        P2_U3012) );
  AOI211_X1 U20451 ( .C1(n17218), .C2(n17203), .A(n17202), .B(n17216), .ZN(
        n17205) );
  NOR2_X1 U20452 ( .A1(n17205), .A2(n17204), .ZN(n17207) );
  NAND3_X1 U20453 ( .A1(n17230), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n17220), .ZN(n17206) );
  OAI211_X1 U20454 ( .C1(n17208), .C2(n17444), .A(n17207), .B(n17206), .ZN(
        n17211) );
  NOR2_X1 U20455 ( .A1(n17209), .A2(n17429), .ZN(n17210) );
  AOI211_X1 U20456 ( .C1(n17212), .C2(n17454), .A(n17211), .B(n17210), .ZN(
        n17213) );
  OAI21_X1 U20457 ( .B1(n17214), .B2(n17458), .A(n17213), .ZN(P2_U3020) );
  NAND2_X1 U20458 ( .A1(n17215), .A2(n17412), .ZN(n17227) );
  INV_X1 U20459 ( .A(n17216), .ZN(n17219) );
  AOI21_X1 U20460 ( .B1(n17219), .B2(n17218), .A(n17217), .ZN(n17222) );
  NAND3_X1 U20461 ( .A1(n17230), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n17220), .ZN(n17221) );
  OAI211_X1 U20462 ( .C1(n17223), .C2(n17429), .A(n17222), .B(n17221), .ZN(
        n17224) );
  AOI21_X1 U20463 ( .B1(n17461), .B2(n17225), .A(n17224), .ZN(n17226) );
  OAI211_X1 U20464 ( .C1(n17228), .C2(n17415), .A(n17227), .B(n17226), .ZN(
        P2_U3021) );
  INV_X1 U20465 ( .A(n17229), .ZN(n17233) );
  OAI21_X1 U20466 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17231), .A(
        n17230), .ZN(n17232) );
  OAI211_X1 U20467 ( .C1(n17234), .C2(n17444), .A(n17233), .B(n17232), .ZN(
        n17237) );
  NOR2_X1 U20468 ( .A1(n17235), .A2(n17429), .ZN(n17236) );
  OAI21_X1 U20469 ( .B1(n17239), .B2(n17458), .A(n17238), .ZN(P2_U3022) );
  NAND2_X1 U20470 ( .A1(n17240), .A2(n17456), .ZN(n17247) );
  INV_X1 U20471 ( .A(n17241), .ZN(n17254) );
  OAI21_X1 U20472 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n17242), .ZN(n17243) );
  NOR2_X1 U20473 ( .A1(n17253), .A2(n17243), .ZN(n17244) );
  AOI211_X1 U20474 ( .C1(n17254), .C2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n17245), .B(n17244), .ZN(n17246) );
  OAI211_X1 U20475 ( .C1(n17444), .C2(n17248), .A(n17247), .B(n17246), .ZN(
        n17249) );
  AOI21_X1 U20476 ( .B1(n17250), .B2(n17412), .A(n17249), .ZN(n17251) );
  OAI21_X1 U20477 ( .B1(n17415), .B2(n17252), .A(n17251), .ZN(P2_U3023) );
  INV_X1 U20478 ( .A(n17253), .ZN(n17255) );
  MUX2_X1 U20479 ( .A(n17255), .B(n17254), .S(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17256) );
  AOI211_X1 U20480 ( .C1(n17810), .C2(n17461), .A(n17257), .B(n17256), .ZN(
        n17258) );
  OAI21_X1 U20481 ( .B1(n17259), .B2(n17429), .A(n17258), .ZN(n17260) );
  AOI21_X1 U20482 ( .B1(n17261), .B2(n17412), .A(n17260), .ZN(n17262) );
  OAI21_X1 U20483 ( .B1(n17415), .B2(n17263), .A(n17262), .ZN(P2_U3024) );
  XNOR2_X1 U20484 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17264) );
  NOR2_X1 U20485 ( .A1(n17265), .A2(n17264), .ZN(n17266) );
  AOI211_X1 U20486 ( .C1(n17281), .C2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n17267), .B(n17266), .ZN(n17270) );
  NAND2_X1 U20487 ( .A1(n17268), .A2(n17461), .ZN(n17269) );
  OAI211_X1 U20488 ( .C1(n17271), .C2(n17429), .A(n17270), .B(n17269), .ZN(
        n17272) );
  AOI21_X1 U20489 ( .B1(n17273), .B2(n17454), .A(n17272), .ZN(n17274) );
  OAI21_X1 U20490 ( .B1(n17275), .B2(n17458), .A(n17274), .ZN(P2_U3026) );
  NOR2_X1 U20491 ( .A1(n17276), .A2(n17429), .ZN(n17285) );
  AND3_X1 U20492 ( .A1(n17291), .A2(n17278), .A3(n17277), .ZN(n17279) );
  AOI211_X1 U20493 ( .C1(n17281), .C2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17280), .B(n17279), .ZN(n17282) );
  OAI21_X1 U20494 ( .B1(n17283), .B2(n17444), .A(n17282), .ZN(n17284) );
  AOI211_X1 U20495 ( .C1(n17286), .C2(n17454), .A(n17285), .B(n17284), .ZN(
        n17287) );
  OAI21_X1 U20496 ( .B1(n17288), .B2(n17458), .A(n17287), .ZN(P2_U3028) );
  INV_X1 U20497 ( .A(n17289), .ZN(n17290) );
  AOI21_X1 U20498 ( .B1(n17291), .B2(n10458), .A(n17290), .ZN(n17294) );
  NAND2_X1 U20499 ( .A1(n17292), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17293) );
  OAI211_X1 U20500 ( .C1(n20108), .C2(n17444), .A(n17294), .B(n17293), .ZN(
        n17297) );
  AOI211_X1 U20501 ( .C1(n20110), .C2(n17456), .A(n17297), .B(n17296), .ZN(
        n17298) );
  OAI21_X1 U20502 ( .B1(n17299), .B2(n17458), .A(n17298), .ZN(P2_U3031) );
  AND2_X1 U20503 ( .A1(n17301), .A2(n17300), .ZN(n17330) );
  INV_X1 U20504 ( .A(n17301), .ZN(n17305) );
  NAND2_X1 U20505 ( .A1(n10181), .A2(n17305), .ZN(n17302) );
  NAND2_X1 U20506 ( .A1(n17303), .A2(n17302), .ZN(n17334) );
  AOI21_X1 U20507 ( .B1(n17330), .B2(n17304), .A(n17334), .ZN(n17316) );
  NOR3_X1 U20508 ( .A1(n17305), .A2(n17329), .A3(n17370), .ZN(n17315) );
  NAND3_X1 U20509 ( .A1(n17315), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n17308), .ZN(n17306) );
  OAI211_X1 U20510 ( .C1(n17316), .C2(n17308), .A(n17307), .B(n17306), .ZN(
        n17310) );
  NOR2_X1 U20511 ( .A1(n20127), .A2(n17429), .ZN(n17309) );
  AOI211_X1 U20512 ( .C1(n17461), .C2(n20128), .A(n17310), .B(n17309), .ZN(
        n17313) );
  NAND2_X1 U20513 ( .A1(n17311), .A2(n17454), .ZN(n17312) );
  OAI211_X1 U20514 ( .C1(n17314), .C2(n17458), .A(n17313), .B(n17312), .ZN(
        P2_U3032) );
  INV_X1 U20515 ( .A(n17315), .ZN(n17317) );
  AOI21_X1 U20516 ( .B1(n17318), .B2(n17317), .A(n17316), .ZN(n17319) );
  AOI211_X1 U20517 ( .C1(n17461), .C2(n17321), .A(n17320), .B(n17319), .ZN(
        n17322) );
  OAI21_X1 U20518 ( .B1(n17429), .B2(n17323), .A(n17322), .ZN(n17324) );
  AOI21_X1 U20519 ( .B1(n17325), .B2(n17412), .A(n17324), .ZN(n17326) );
  OAI21_X1 U20520 ( .B1(n17327), .B2(n17415), .A(n17326), .ZN(P2_U3033) );
  INV_X1 U20521 ( .A(n17328), .ZN(n17332) );
  NAND2_X1 U20522 ( .A1(n17330), .A2(n17329), .ZN(n17331) );
  NAND2_X1 U20523 ( .A1(n17332), .A2(n17331), .ZN(n17333) );
  AOI21_X1 U20524 ( .B1(n17334), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17333), .ZN(n17337) );
  NAND2_X1 U20525 ( .A1(n17335), .A2(n17461), .ZN(n17336) );
  OAI211_X1 U20526 ( .C1(n17338), .C2(n17429), .A(n17337), .B(n17336), .ZN(
        n17339) );
  AOI21_X1 U20527 ( .B1(n17340), .B2(n17454), .A(n17339), .ZN(n17341) );
  OAI21_X1 U20528 ( .B1(n17342), .B2(n17458), .A(n17341), .ZN(P2_U3034) );
  NOR2_X1 U20529 ( .A1(n17370), .A2(n17348), .ZN(n17358) );
  NOR2_X1 U20530 ( .A1(n17361), .A2(n17349), .ZN(n17343) );
  AOI21_X1 U20531 ( .B1(n17361), .B2(n17349), .A(n17343), .ZN(n17344) );
  NAND2_X1 U20532 ( .A1(n17358), .A2(n17344), .ZN(n17345) );
  OAI211_X1 U20533 ( .C1(n17347), .C2(n17444), .A(n17346), .B(n17345), .ZN(
        n17351) );
  NOR2_X1 U20534 ( .A1(n17378), .A2(n17348), .ZN(n17363) );
  NOR3_X1 U20535 ( .A1(n17363), .A2(n17362), .A3(n17349), .ZN(n17350) );
  AOI211_X1 U20536 ( .C1(n17352), .C2(n17456), .A(n17351), .B(n17350), .ZN(
        n17355) );
  NAND2_X1 U20537 ( .A1(n17353), .A2(n17454), .ZN(n17354) );
  OAI211_X1 U20538 ( .C1(n17356), .C2(n17458), .A(n17355), .B(n17354), .ZN(
        P2_U3035) );
  NAND2_X1 U20539 ( .A1(n17357), .A2(n17412), .ZN(n17368) );
  NAND2_X1 U20540 ( .A1(n17358), .A2(n17361), .ZN(n17359) );
  OAI211_X1 U20541 ( .C1(n20139), .C2(n17444), .A(n17360), .B(n17359), .ZN(
        n17365) );
  NOR3_X1 U20542 ( .A1(n17363), .A2(n17362), .A3(n17361), .ZN(n17364) );
  AOI211_X1 U20543 ( .C1(n17366), .C2(n17456), .A(n17365), .B(n17364), .ZN(
        n17367) );
  OAI211_X1 U20544 ( .C1(n17369), .C2(n17415), .A(n17368), .B(n17367), .ZN(
        P2_U3036) );
  NOR2_X1 U20545 ( .A1(n17370), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17371) );
  NOR2_X1 U20546 ( .A1(n17372), .A2(n17371), .ZN(n17375) );
  NAND2_X1 U20547 ( .A1(n17373), .A2(n17461), .ZN(n17374) );
  OAI211_X1 U20548 ( .C1(n20155), .C2(n17429), .A(n17375), .B(n17374), .ZN(
        n17377) );
  NAND3_X1 U20549 ( .A1(n17406), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n17397), .ZN(n17396) );
  AOI21_X1 U20550 ( .B1(n17405), .B2(n10181), .A(n17404), .ZN(n17398) );
  AOI21_X1 U20551 ( .B1(n17396), .B2(n17398), .A(n17384), .ZN(n17388) );
  NOR2_X1 U20552 ( .A1(n17380), .A2(n17444), .ZN(n17381) );
  AOI211_X1 U20553 ( .C1(n17384), .C2(n17383), .A(n17382), .B(n17381), .ZN(
        n17385) );
  OAI21_X1 U20554 ( .B1(n17429), .B2(n17386), .A(n17385), .ZN(n17387) );
  AOI211_X1 U20555 ( .C1(n17389), .C2(n17412), .A(n17388), .B(n17387), .ZN(
        n17390) );
  OAI21_X1 U20556 ( .B1(n17391), .B2(n17415), .A(n17390), .ZN(P2_U3038) );
  INV_X1 U20557 ( .A(n20173), .ZN(n17394) );
  OAI21_X1 U20558 ( .B1(n20172), .B2(n17444), .A(n17392), .ZN(n17393) );
  AOI21_X1 U20559 ( .B1(n17394), .B2(n17456), .A(n17393), .ZN(n17395) );
  OAI211_X1 U20560 ( .C1(n17398), .C2(n17397), .A(n17396), .B(n17395), .ZN(
        n17399) );
  AOI21_X1 U20561 ( .B1(n17400), .B2(n17412), .A(n17399), .ZN(n17401) );
  OAI21_X1 U20562 ( .B1(n17415), .B2(n17402), .A(n17401), .ZN(P2_U3039) );
  NOR2_X1 U20563 ( .A1(n20856), .A2(n17149), .ZN(n17403) );
  AOI221_X1 U20564 ( .B1(n17406), .B2(n17405), .C1(n17404), .C2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n17403), .ZN(n17407) );
  INV_X1 U20565 ( .A(n17407), .ZN(n17411) );
  OAI22_X1 U20566 ( .A1(n17409), .A2(n17429), .B1(n17444), .B2(n17408), .ZN(
        n17410) );
  AOI211_X1 U20567 ( .C1(n17413), .C2(n17412), .A(n17411), .B(n17410), .ZN(
        n17414) );
  OAI21_X1 U20568 ( .B1(n17416), .B2(n17415), .A(n17414), .ZN(P2_U3040) );
  AOI211_X1 U20569 ( .C1(n17423), .C2(n17432), .A(n17417), .B(n17433), .ZN(
        n17425) );
  AOI21_X1 U20570 ( .B1(n17461), .B2(n17419), .A(n17418), .ZN(n17422) );
  NAND2_X1 U20571 ( .A1(n17420), .A2(n17456), .ZN(n17421) );
  OAI211_X1 U20572 ( .C1(n17431), .C2(n17423), .A(n17422), .B(n17421), .ZN(
        n17424) );
  AOI211_X1 U20573 ( .C1(n17426), .C2(n17454), .A(n17425), .B(n17424), .ZN(
        n17427) );
  OAI21_X1 U20574 ( .B1(n17428), .B2(n17458), .A(n17427), .ZN(P2_U3041) );
  OAI22_X1 U20575 ( .A1(n20203), .A2(n17429), .B1(n17444), .B2(n20179), .ZN(
        n17435) );
  NAND2_X1 U20576 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n20167), .ZN(n17430) );
  OAI221_X1 U20577 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n17433), .C1(
        n17432), .C2(n17431), .A(n17430), .ZN(n17434) );
  AOI211_X1 U20578 ( .C1(n17454), .C2(n17436), .A(n17435), .B(n17434), .ZN(
        n17437) );
  OAI21_X1 U20579 ( .B1(n17438), .B2(n17458), .A(n17437), .ZN(P2_U3042) );
  MUX2_X1 U20580 ( .A(n17440), .B(n17439), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n17441) );
  AOI21_X1 U20581 ( .B1(n20167), .B2(P2_REIP_REG_3__SCAN_IN), .A(n17441), .ZN(
        n17442) );
  OAI21_X1 U20582 ( .B1(n17444), .B2(n17443), .A(n17442), .ZN(n17445) );
  AOI21_X1 U20583 ( .B1(n17456), .B2(n17446), .A(n17445), .ZN(n17449) );
  NAND3_X1 U20584 ( .A1(n17177), .A2(n17447), .A3(n17454), .ZN(n17448) );
  OAI211_X1 U20585 ( .C1(n17450), .C2(n17458), .A(n17449), .B(n17448), .ZN(
        P2_U3043) );
  MUX2_X1 U20586 ( .A(n17452), .B(n17451), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n17464) );
  AOI22_X1 U20587 ( .A1(n17456), .A2(n17455), .B1(n17454), .B2(n17453), .ZN(
        n17463) );
  NOR2_X1 U20588 ( .A1(n17458), .A2(n17457), .ZN(n17459) );
  AOI211_X1 U20589 ( .C1(n20229), .C2(n17461), .A(n17460), .B(n17459), .ZN(
        n17462) );
  NAND3_X1 U20590 ( .A1(n17464), .A2(n17463), .A3(n17462), .ZN(P2_U3046) );
  OAI222_X1 U20591 ( .A1(n17484), .A2(n12229), .B1(n11055), .B2(n17467), .C1(
        n17476), .C2(n17465), .ZN(n17466) );
  MUX2_X1 U20592 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n17466), .S(
        n17478), .Z(P2_U3601) );
  NAND3_X1 U20593 ( .A1(n17468), .A2(P2_STATE2_REG_1__SCAN_IN), .A3(n17467), 
        .ZN(n17472) );
  AOI22_X1 U20594 ( .A1(n20931), .A2(n17470), .B1(n20911), .B2(n17469), .ZN(
        n17471) );
  NAND2_X1 U20595 ( .A1(n17472), .A2(n17471), .ZN(n17473) );
  MUX2_X1 U20596 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n17473), .S(
        n17478), .Z(P2_U3600) );
  OAI22_X1 U20597 ( .A1(n20324), .A2(n17484), .B1(n17474), .B2(n17476), .ZN(
        n17475) );
  MUX2_X1 U20598 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n17475), .S(
        n17478), .Z(P2_U3596) );
  NOR2_X1 U20599 ( .A1(n17477), .A2(n17476), .ZN(n17479) );
  MUX2_X1 U20600 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n17479), .S(
        n17478), .Z(P2_U3595) );
  OAI21_X1 U20601 ( .B1(n20476), .B2(n20529), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n17487) );
  NAND2_X1 U20602 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20920), .ZN(
        n20451) );
  INV_X1 U20603 ( .A(n20451), .ZN(n20503) );
  NAND2_X1 U20604 ( .A1(n20419), .A2(n20503), .ZN(n17486) );
  NAND2_X1 U20605 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20947), .ZN(
        n20357) );
  NOR2_X1 U20606 ( .A1(n20357), .A2(n20451), .ZN(n20495) );
  NOR2_X1 U20607 ( .A1(n20495), .A2(n20939), .ZN(n17481) );
  NAND2_X1 U20608 ( .A1(n10903), .A2(n17481), .ZN(n17492) );
  OAI211_X1 U20609 ( .C1(n20495), .C2(n17491), .A(n17492), .B(n20697), .ZN(
        n17485) );
  AOI21_X1 U20610 ( .B1(n17487), .B2(n17486), .A(n17485), .ZN(n20482) );
  INV_X1 U20611 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17498) );
  AOI22_X1 U20612 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20315), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n20314), .ZN(n20701) );
  AOI22_X1 U20613 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20315), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20314), .ZN(n20663) );
  INV_X1 U20614 ( .A(n20663), .ZN(n20756) );
  AOI22_X1 U20615 ( .A1(n20476), .A2(n20757), .B1(n20529), .B2(n20756), .ZN(
        n17497) );
  NAND3_X1 U20616 ( .A1(n20419), .A2(n20503), .A3(n17491), .ZN(n17494) );
  INV_X1 U20617 ( .A(n17492), .ZN(n17493) );
  NOR2_X2 U20618 ( .A1(n20510), .A2(n20233), .ZN(n20692) );
  NOR2_X2 U20619 ( .A1(n20317), .A2(n17495), .ZN(n20691) );
  AOI22_X1 U20620 ( .A1(n20496), .A2(n20692), .B1(n20691), .B2(n20495), .ZN(
        n17496) );
  OAI211_X1 U20621 ( .C1(n20482), .C2(n17498), .A(n17497), .B(n17496), .ZN(
        P2_U3096) );
  OAI21_X1 U20622 ( .B1(n20747), .B2(n20821), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n17500) );
  NAND2_X1 U20623 ( .A1(n17500), .A2(n20958), .ZN(n17502) );
  NAND3_X1 U20624 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n17518) );
  NOR2_X1 U20625 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n17518), .ZN(
        n20746) );
  NAND3_X1 U20626 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20938), .ZN(n20693) );
  NOR2_X1 U20627 ( .A1(n20947), .A2(n20693), .ZN(n20720) );
  NOR2_X1 U20628 ( .A1(n20746), .A2(n20720), .ZN(n17505) );
  OAI21_X1 U20629 ( .B1(n17503), .B2(n20746), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17501) );
  INV_X1 U20630 ( .A(n20748), .ZN(n17514) );
  INV_X1 U20631 ( .A(n20692), .ZN(n20754) );
  INV_X1 U20632 ( .A(n17502), .ZN(n17506) );
  AOI211_X1 U20633 ( .C1(n17503), .C2(n17491), .A(n20958), .B(n20746), .ZN(
        n17504) );
  INV_X1 U20634 ( .A(n20752), .ZN(n17512) );
  NOR2_X1 U20635 ( .A1(n20701), .A2(n17507), .ZN(n17511) );
  INV_X1 U20636 ( .A(n20691), .ZN(n20753) );
  INV_X1 U20637 ( .A(n20746), .ZN(n17508) );
  OAI22_X1 U20638 ( .A1(n20663), .A2(n17509), .B1(n20753), .B2(n17508), .ZN(
        n17510) );
  AOI211_X1 U20639 ( .C1(n17512), .C2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n17511), .B(n17510), .ZN(n17513) );
  OAI21_X1 U20640 ( .B1(n17514), .B2(n20754), .A(n17513), .ZN(P2_U3160) );
  NAND2_X1 U20641 ( .A1(n20918), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20624) );
  INV_X1 U20642 ( .A(n20624), .ZN(n20565) );
  NAND2_X1 U20643 ( .A1(n20565), .A2(n20501), .ZN(n17517) );
  NAND2_X1 U20644 ( .A1(n20814), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n17515) );
  NOR2_X1 U20645 ( .A1(n10820), .A2(n17515), .ZN(n17521) );
  INV_X1 U20646 ( .A(n20814), .ZN(n20290) );
  OAI21_X1 U20647 ( .B1(n20290), .B2(n17491), .A(n20697), .ZN(n17516) );
  INV_X1 U20648 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17527) );
  INV_X1 U20649 ( .A(n17518), .ZN(n17519) );
  AOI21_X1 U20650 ( .B1(n17491), .B2(n17519), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17520) );
  INV_X1 U20651 ( .A(n20816), .ZN(n17525) );
  NOR2_X2 U20652 ( .A1(n20225), .A2(n20510), .ZN(n20730) );
  NOR2_X2 U20653 ( .A1(n20317), .A2(n9989), .ZN(n20727) );
  INV_X1 U20654 ( .A(n20727), .ZN(n17523) );
  AOI22_X1 U20655 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20315), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20314), .ZN(n20666) );
  AOI22_X1 U20656 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20315), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n20314), .ZN(n20704) );
  INV_X1 U20657 ( .A(n20704), .ZN(n20729) );
  AOI22_X1 U20658 ( .A1(n20819), .A2(n20728), .B1(n20821), .B2(n20729), .ZN(
        n17522) );
  OAI21_X1 U20659 ( .B1(n17523), .B2(n20814), .A(n17522), .ZN(n17524) );
  AOI21_X1 U20660 ( .B1(n17525), .B2(n20730), .A(n17524), .ZN(n17526) );
  OAI21_X1 U20661 ( .B1(n20825), .B2(n17527), .A(n17526), .ZN(P2_U3169) );
  INV_X1 U20662 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n18205) );
  INV_X1 U20663 ( .A(n18533), .ZN(n17528) );
  NAND3_X1 U20664 ( .A1(n17528), .A2(n18576), .A3(P3_EBX_REG_21__SCAN_IN), 
        .ZN(n17679) );
  NAND3_X1 U20665 ( .A1(n17679), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n18586), 
        .ZN(n17544) );
  INV_X1 U20666 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17529) );
  NOR2_X1 U20667 ( .A1(n18541), .A2(n17529), .ZN(n17535) );
  AOI22_X1 U20668 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17533) );
  AOI22_X1 U20669 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17532) );
  AOI22_X1 U20670 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17531) );
  NAND2_X1 U20671 ( .A1(n11944), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n17530) );
  NAND4_X1 U20672 ( .A1(n17533), .A2(n17532), .A3(n17531), .A4(n17530), .ZN(
        n17534) );
  AOI211_X1 U20673 ( .C1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .C2(n18523), .A(
        n17535), .B(n17534), .ZN(n17542) );
  AOI22_X1 U20674 ( .A1(n17705), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17541) );
  AOI22_X1 U20675 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17540) );
  INV_X1 U20676 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17537) );
  OAI22_X1 U20677 ( .A1(n18464), .A2(n17537), .B1(n17767), .B2(n17536), .ZN(
        n17538) );
  AOI21_X1 U20678 ( .B1(n9867), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(n17538), .ZN(n17539) );
  NAND4_X1 U20679 ( .A1(n17542), .A2(n17541), .A3(n17540), .A4(n17539), .ZN(
        n18637) );
  NAND2_X1 U20680 ( .A1(n18590), .A2(n18637), .ZN(n17543) );
  OAI211_X1 U20681 ( .C1(n17679), .C2(P3_EBX_REG_22__SCAN_IN), .A(n17544), .B(
        n17543), .ZN(P3_U2681) );
  NAND2_X1 U20682 ( .A1(n18533), .A2(n18586), .ZN(n18536) );
  NOR2_X1 U20683 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17549), .ZN(n17546) );
  OAI22_X1 U20684 ( .A1(n18536), .A2(n17546), .B1(n17545), .B2(n18586), .ZN(
        P3_U2683) );
  OAI21_X1 U20685 ( .B1(n9842), .B2(P3_EBX_REG_19__SCAN_IN), .A(n18586), .ZN(
        n17548) );
  OAI22_X1 U20686 ( .A1(n17549), .A2(n17548), .B1(n17547), .B2(n18586), .ZN(
        P3_U2684) );
  NAND2_X1 U20687 ( .A1(n17639), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17552) );
  NAND2_X1 U20688 ( .A1(n17552), .A2(n19121), .ZN(n17576) );
  NAND2_X1 U20689 ( .A1(n17609), .A2(n18978), .ZN(n17553) );
  NAND2_X1 U20690 ( .A1(n17576), .A2(n17553), .ZN(n17579) );
  NOR2_X1 U20691 ( .A1(n17554), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17555) );
  NAND2_X1 U20692 ( .A1(n17651), .A2(n17555), .ZN(n17617) );
  XNOR2_X1 U20693 ( .A(n9855), .B(n10296), .ZN(n18084) );
  INV_X1 U20694 ( .A(n17556), .ZN(n17558) );
  INV_X1 U20695 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n17557) );
  NOR2_X1 U20696 ( .A1(n19110), .A2(n17557), .ZN(n17619) );
  AOI21_X1 U20697 ( .B1(n17558), .B2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n17619), .ZN(n17559) );
  OAI21_X1 U20698 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n17560), .A(
        n17559), .ZN(n17561) );
  AOI21_X1 U20699 ( .B1(n18977), .B2(n18084), .A(n17561), .ZN(n17562) );
  OAI21_X1 U20700 ( .B1(n18933), .B2(n17617), .A(n17562), .ZN(n17563) );
  AOI21_X1 U20701 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17579), .A(
        n17563), .ZN(n17564) );
  XOR2_X1 U20702 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n17565), .Z(
        n17630) );
  NAND4_X1 U20703 ( .A1(n17609), .A2(n17566), .A3(n18813), .A4(n18978), .ZN(
        n17575) );
  INV_X1 U20704 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n17567) );
  NOR2_X1 U20705 ( .A1(n19349), .A2(n17567), .ZN(n17627) );
  NOR3_X1 U20706 ( .A1(n17569), .A2(n17588), .A3(n17568), .ZN(n17570) );
  AOI211_X1 U20707 ( .C1(n17571), .C2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n17627), .B(n17570), .ZN(n17574) );
  AOI21_X1 U20708 ( .B1(n12123), .B2(n17572), .A(n9855), .ZN(n18092) );
  NAND2_X1 U20709 ( .A1(n19122), .A2(n18092), .ZN(n17573) );
  NAND3_X1 U20710 ( .A1(n17575), .A2(n17574), .A3(n17573), .ZN(n17578) );
  INV_X1 U20711 ( .A(n17639), .ZN(n17611) );
  NOR2_X1 U20712 ( .A1(n17576), .A2(n17611), .ZN(n17577) );
  AOI211_X1 U20713 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n17579), .A(
        n17578), .B(n17577), .ZN(n17580) );
  OAI21_X1 U20714 ( .B1(n17630), .B2(n19034), .A(n17580), .ZN(P3_U2801) );
  NOR2_X1 U20715 ( .A1(n17582), .A2(n17581), .ZN(n17583) );
  XNOR2_X1 U20716 ( .A(n17583), .B(n18950), .ZN(n17668) );
  OAI21_X1 U20717 ( .B1(n18933), .B2(n17584), .A(n17662), .ZN(n17594) );
  AOI21_X1 U20718 ( .B1(n17586), .B2(n18115), .A(n17585), .ZN(n18114) );
  INV_X1 U20719 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n17587) );
  NOR2_X1 U20720 ( .A1(n19349), .A2(n17587), .ZN(n17666) );
  NOR3_X1 U20721 ( .A1(n18891), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17588), .ZN(n17589) );
  AOI211_X1 U20722 ( .C1(n18977), .C2(n18114), .A(n17666), .B(n17589), .ZN(
        n17590) );
  OAI21_X1 U20723 ( .B1(n17591), .B2(n18115), .A(n17590), .ZN(n17592) );
  AOI21_X1 U20724 ( .B1(n17594), .B2(n17593), .A(n17592), .ZN(n17595) );
  OAI21_X1 U20725 ( .B1(n17668), .B2(n19034), .A(n17595), .ZN(P3_U2803) );
  INV_X1 U20726 ( .A(n18815), .ZN(n17596) );
  AOI21_X1 U20727 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17597), .A(
        n17596), .ZN(n17678) );
  NOR2_X1 U20728 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17598), .ZN(
        n17675) );
  AOI22_X1 U20729 ( .A1(n18978), .A2(n19236), .B1(n19121), .B2(n19230), .ZN(
        n18932) );
  OAI21_X1 U20730 ( .B1(n17671), .B2(n18933), .A(n18932), .ZN(n18834) );
  INV_X1 U20731 ( .A(n18834), .ZN(n17605) );
  NOR2_X1 U20732 ( .A1(n18891), .A2(n17600), .ZN(n18810) );
  INV_X1 U20733 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18156) );
  NAND2_X1 U20734 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17599), .ZN(
        n18059) );
  AND2_X1 U20735 ( .A1(n17600), .A2(n19801), .ZN(n18829) );
  AOI211_X1 U20736 ( .C1(n17601), .C2(n18059), .A(n18829), .B(n19096), .ZN(
        n18827) );
  OAI21_X1 U20737 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18868), .A(
        n18827), .ZN(n18825) );
  INV_X1 U20738 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19989) );
  NOR2_X1 U20739 ( .A1(n18156), .A2(n18066), .ZN(n18070) );
  AOI21_X1 U20740 ( .B1(n18156), .B2(n18066), .A(n18070), .ZN(n18151) );
  INV_X1 U20741 ( .A(n18151), .ZN(n17602) );
  OAI22_X1 U20742 ( .A1(n19349), .A2(n19989), .B1(n18985), .B2(n17602), .ZN(
        n17603) );
  AOI221_X1 U20743 ( .B1(n18810), .B2(n18156), .C1(n18825), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17603), .ZN(n17604) );
  OAI21_X1 U20744 ( .B1(n10160), .B2(n17605), .A(n17604), .ZN(n17606) );
  AOI21_X1 U20745 ( .B1(n18847), .B2(n17675), .A(n17606), .ZN(n17607) );
  OAI21_X1 U20746 ( .B1(n17678), .B2(n19034), .A(n17607), .ZN(P3_U2806) );
  AND2_X1 U20747 ( .A1(n19370), .A2(n17608), .ZN(n17610) );
  AOI22_X1 U20748 ( .A1(n17611), .A2(n19351), .B1(n17610), .B2(n17609), .ZN(
        n17625) );
  OAI211_X1 U20749 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n19377), .A(
        n17625), .B(n17612), .ZN(n17620) );
  NAND2_X1 U20750 ( .A1(n19280), .A2(n19875), .ZN(n17614) );
  NAND2_X1 U20751 ( .A1(n19281), .A2(n19263), .ZN(n17613) );
  NAND2_X1 U20752 ( .A1(n17614), .A2(n17613), .ZN(n19197) );
  NAND2_X1 U20753 ( .A1(n19197), .A2(n10157), .ZN(n17616) );
  INV_X1 U20754 ( .A(n19139), .ZN(n17615) );
  NAND2_X1 U20755 ( .A1(n17616), .A2(n17615), .ZN(n19167) );
  INV_X1 U20756 ( .A(n19192), .ZN(n19181) );
  NOR2_X1 U20757 ( .A1(n19181), .A2(n17617), .ZN(n17618) );
  AOI211_X1 U20758 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n17620), .A(
        n17619), .B(n17618), .ZN(n17621) );
  OAI21_X1 U20759 ( .B1(n17622), .B2(n19311), .A(n17621), .ZN(P3_U2832) );
  OAI211_X1 U20760 ( .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n19289), .A(
        n17623), .B(n19341), .ZN(n17635) );
  NAND2_X1 U20761 ( .A1(n17635), .A2(n19110), .ZN(n17624) );
  OAI211_X1 U20762 ( .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n19361), .A(
        n17625), .B(n17624), .ZN(n17628) );
  NOR3_X1 U20763 ( .A1(n19181), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n17636), .ZN(n17626) );
  AOI211_X1 U20764 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n17628), .A(
        n17627), .B(n17626), .ZN(n17629) );
  OAI21_X1 U20765 ( .B1(n17630), .B2(n19311), .A(n17629), .ZN(P3_U2833) );
  AOI22_X1 U20766 ( .A1(n17633), .A2(n19370), .B1(n19192), .B2(n17631), .ZN(
        n17649) );
  NAND2_X1 U20767 ( .A1(n19391), .A2(n17632), .ZN(n19326) );
  NOR3_X1 U20768 ( .A1(n17634), .A2(n17633), .A3(n19326), .ZN(n17641) );
  INV_X1 U20769 ( .A(n17635), .ZN(n17638) );
  OAI21_X1 U20770 ( .B1(n19236), .B2(n17636), .A(n19263), .ZN(n17637) );
  OAI211_X1 U20771 ( .C1(n17639), .C2(n19387), .A(n17638), .B(n17637), .ZN(
        n17640) );
  OAI211_X1 U20772 ( .C1(n17641), .C2(n17640), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n19110), .ZN(n17648) );
  INV_X1 U20773 ( .A(n17642), .ZN(n17643) );
  NOR3_X1 U20774 ( .A1(n17644), .A2(n17643), .A3(n19311), .ZN(n17646) );
  NOR2_X1 U20775 ( .A1(n17646), .A2(n17645), .ZN(n17647) );
  OAI211_X1 U20776 ( .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n17649), .A(
        n17648), .B(n17647), .ZN(P3_U2834) );
  INV_X1 U20777 ( .A(n19167), .ZN(n17650) );
  NOR2_X1 U20778 ( .A1(n17650), .A2(n18797), .ZN(n19151) );
  AOI21_X1 U20779 ( .B1(n19151), .B2(n17651), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17664) );
  INV_X1 U20780 ( .A(n19168), .ZN(n18839) );
  NOR2_X1 U20781 ( .A1(n19198), .A2(n18839), .ZN(n19155) );
  OAI211_X1 U20782 ( .C1(n19306), .C2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n19155), .ZN(n17669) );
  NAND2_X1 U20783 ( .A1(n19220), .A2(n19306), .ZN(n19380) );
  OAI21_X1 U20784 ( .B1(n19133), .B2(n17669), .A(n19380), .ZN(n19135) );
  INV_X1 U20785 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n19140) );
  NAND2_X1 U20786 ( .A1(n19160), .A2(n19140), .ZN(n17658) );
  INV_X1 U20787 ( .A(n17652), .ZN(n17654) );
  AOI22_X1 U20788 ( .A1(n19283), .A2(n17654), .B1(n19263), .B2(n17653), .ZN(
        n17657) );
  INV_X1 U20789 ( .A(n17655), .ZN(n17656) );
  NAND3_X1 U20790 ( .A1(n17658), .A2(n17657), .A3(n17656), .ZN(n17659) );
  AOI21_X1 U20791 ( .B1(n19875), .B2(n17660), .A(n17659), .ZN(n17661) );
  NAND2_X1 U20792 ( .A1(n19135), .A2(n17661), .ZN(n19128) );
  AOI211_X1 U20793 ( .C1(n18799), .C2(n19160), .A(n17662), .B(n19128), .ZN(
        n17663) );
  NOR3_X1 U20794 ( .A1(n17664), .A2(n19399), .A3(n17663), .ZN(n17665) );
  AOI211_X1 U20795 ( .C1(n19396), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17666), .B(n17665), .ZN(n17667) );
  OAI21_X1 U20796 ( .B1(n17668), .B2(n19311), .A(n17667), .ZN(P3_U2835) );
  NOR2_X1 U20797 ( .A1(n19875), .A2(n19263), .ZN(n19286) );
  AOI21_X1 U20798 ( .B1(n19380), .B2(n17669), .A(n19396), .ZN(n17670) );
  OAI211_X1 U20799 ( .C1(n17671), .C2(n19286), .A(n19223), .B(n17670), .ZN(
        n17674) );
  NOR2_X1 U20800 ( .A1(n17672), .A2(n17674), .ZN(n17673) );
  OAI21_X1 U20801 ( .B1(n18797), .B2(n19156), .A(n19876), .ZN(n19134) );
  AOI21_X1 U20802 ( .B1(n17673), .B2(n19134), .A(n19302), .ZN(n19150) );
  OAI211_X1 U20803 ( .C1(n17674), .C2(n19318), .A(n19150), .B(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17677) );
  AOI22_X1 U20804 ( .A1(n19192), .A2(n17675), .B1(n19302), .B2(
        P3_REIP_REG_24__SCAN_IN), .ZN(n17676) );
  OAI211_X1 U20805 ( .C1(n17678), .C2(n19311), .A(n17677), .B(n17676), .ZN(
        P3_U2838) );
  INV_X1 U20806 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n18447) );
  INV_X1 U20807 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n18140) );
  INV_X1 U20808 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n18172) );
  NAND3_X1 U20809 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(n18511), .ZN(n18501) );
  NOR2_X2 U20810 ( .A1(n18140), .A2(n18501), .ZN(n18505) );
  INV_X1 U20811 ( .A(n18492), .ZN(n17796) );
  AOI21_X1 U20812 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n18586), .A(n18496), .ZN(
        n17795) );
  INV_X1 U20813 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17681) );
  INV_X1 U20814 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17680) );
  OAI22_X1 U20815 ( .A1(n17681), .A2(n18539), .B1(n18541), .B2(n17680), .ZN(
        n17694) );
  AOI22_X1 U20816 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17705), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17686) );
  AOI22_X1 U20817 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17784), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17685) );
  AOI22_X1 U20818 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17684) );
  NAND2_X1 U20819 ( .A1(n17682), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n17683) );
  NAND4_X1 U20820 ( .A1(n17686), .A2(n17685), .A3(n17684), .A4(n17683), .ZN(
        n17693) );
  AOI22_X1 U20821 ( .A1(n17762), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17691) );
  AOI22_X1 U20822 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17690) );
  AOI22_X1 U20823 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17689) );
  INV_X1 U20824 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17687) );
  OR2_X1 U20825 ( .A1(n18545), .A2(n17687), .ZN(n17688) );
  NAND4_X1 U20826 ( .A1(n17691), .A2(n17690), .A3(n17689), .A4(n17688), .ZN(
        n17692) );
  NOR3_X1 U20827 ( .A1(n17694), .A2(n17693), .A3(n17692), .ZN(n17793) );
  INV_X1 U20828 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17696) );
  AOI22_X1 U20829 ( .A1(n17762), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17695) );
  OAI21_X1 U20830 ( .B1(n17696), .B2(n17765), .A(n17695), .ZN(n17711) );
  INV_X1 U20831 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17698) );
  INV_X1 U20832 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17697) );
  OAI22_X1 U20833 ( .A1(n18541), .A2(n17698), .B1(n18539), .B2(n17697), .ZN(
        n17710) );
  AOI22_X1 U20834 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18552), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17704) );
  AOI22_X1 U20835 ( .A1(n17699), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17784), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17703) );
  AOI22_X1 U20836 ( .A1(n17700), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17702) );
  NAND2_X1 U20837 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n17701) );
  NAND4_X1 U20838 ( .A1(n17704), .A2(n17703), .A3(n17702), .A4(n17701), .ZN(
        n17709) );
  AOI22_X1 U20839 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17705), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17707) );
  AOI22_X1 U20840 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17706) );
  NAND2_X1 U20841 ( .A1(n17707), .A2(n17706), .ZN(n17708) );
  NOR4_X1 U20842 ( .A1(n17711), .A2(n17710), .A3(n17709), .A4(n17708), .ZN(
        n18507) );
  AOI22_X1 U20843 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17718) );
  NAND2_X1 U20844 ( .A1(n17785), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n17714) );
  NAND2_X1 U20845 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n17713) );
  NAND2_X1 U20846 ( .A1(n17784), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n17712) );
  AND3_X1 U20847 ( .A1(n17714), .A2(n17713), .A3(n17712), .ZN(n17717) );
  AOI22_X1 U20848 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17716) );
  AOI22_X1 U20849 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17715) );
  NAND4_X1 U20850 ( .A1(n17718), .A2(n17717), .A3(n17716), .A4(n17715), .ZN(
        n17724) );
  AOI22_X1 U20851 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17722) );
  AOI22_X1 U20852 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17721) );
  AOI22_X1 U20853 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17720) );
  OR2_X1 U20854 ( .A1(n18545), .A2(n13550), .ZN(n17719) );
  NAND4_X1 U20855 ( .A1(n17722), .A2(n17721), .A3(n17720), .A4(n17719), .ZN(
        n17723) );
  OR2_X1 U20856 ( .A1(n17724), .A2(n17723), .ZN(n18513) );
  AOI22_X1 U20857 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n11716), .B1(
        n18524), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17732) );
  NAND2_X1 U20858 ( .A1(n17785), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n17726) );
  NAND2_X1 U20859 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n17725) );
  OAI211_X1 U20860 ( .C1(n9756), .C2(n17727), .A(n17726), .B(n17725), .ZN(
        n17728) );
  INV_X1 U20861 ( .A(n17728), .ZN(n17731) );
  AOI22_X1 U20862 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18550), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17730) );
  AOI22_X1 U20863 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17729) );
  NAND4_X1 U20864 ( .A1(n17732), .A2(n17731), .A3(n17730), .A4(n17729), .ZN(
        n17738) );
  AOI22_X1 U20865 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17736) );
  AOI22_X1 U20866 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17735) );
  AOI22_X1 U20867 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17734) );
  OR2_X1 U20868 ( .A1(n18545), .A2(n13723), .ZN(n17733) );
  NAND4_X1 U20869 ( .A1(n17736), .A2(n17735), .A3(n17734), .A4(n17733), .ZN(
        n17737) );
  OR2_X1 U20870 ( .A1(n17738), .A2(n17737), .ZN(n18514) );
  NAND2_X1 U20871 ( .A1(n18513), .A2(n18514), .ZN(n18512) );
  NOR2_X1 U20872 ( .A1(n18507), .A2(n18512), .ZN(n18506) );
  INV_X1 U20873 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17740) );
  INV_X1 U20874 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17739) );
  OAI22_X1 U20875 ( .A1(n18541), .A2(n17740), .B1(n18539), .B2(n17739), .ZN(
        n17751) );
  AOI22_X1 U20876 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17744) );
  AOI22_X1 U20877 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17743) );
  AOI22_X1 U20878 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17742) );
  INV_X1 U20879 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18540) );
  OR2_X1 U20880 ( .A1(n18545), .A2(n18540), .ZN(n17741) );
  NAND4_X1 U20881 ( .A1(n17744), .A2(n17743), .A3(n17742), .A4(n17741), .ZN(
        n17750) );
  AOI22_X1 U20882 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17748) );
  AOI22_X1 U20883 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17747) );
  AOI22_X1 U20884 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17746) );
  NAND2_X1 U20885 ( .A1(n17785), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n17745) );
  NAND4_X1 U20886 ( .A1(n17748), .A2(n17747), .A3(n17746), .A4(n17745), .ZN(
        n17749) );
  OR3_X1 U20887 ( .A1(n17751), .A2(n17750), .A3(n17749), .ZN(n18503) );
  NAND2_X1 U20888 ( .A1(n18506), .A2(n18503), .ZN(n18502) );
  INV_X1 U20889 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17753) );
  OAI22_X1 U20890 ( .A1(n9746), .A2(n17753), .B1(n9756), .B2(n17752), .ZN(
        n17754) );
  AOI21_X1 U20891 ( .B1(n13472), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n17754), .ZN(n17759) );
  AOI22_X1 U20892 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17758) );
  AOI22_X1 U20893 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17755), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17757) );
  AOI22_X1 U20894 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17756) );
  NAND4_X1 U20895 ( .A1(n17759), .A2(n17758), .A3(n17757), .A4(n17756), .ZN(
        n17773) );
  INV_X1 U20896 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17760) );
  OAI22_X1 U20897 ( .A1(n17799), .A2(n17761), .B1(n18464), .B2(n17760), .ZN(
        n17772) );
  AOI22_X1 U20898 ( .A1(n17762), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17763) );
  OAI21_X1 U20899 ( .B1(n17765), .B2(n17764), .A(n17763), .ZN(n17771) );
  INV_X1 U20900 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17768) );
  OAI22_X1 U20901 ( .A1(n17769), .A2(n17768), .B1(n17767), .B2(n17766), .ZN(
        n17770) );
  NOR4_X1 U20902 ( .A1(n17773), .A2(n17772), .A3(n17771), .A4(n17770), .ZN(
        n18498) );
  NOR2_X1 U20903 ( .A1(n18502), .A2(n18498), .ZN(n18497) );
  AOI22_X1 U20904 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17779) );
  AOI22_X1 U20905 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17778) );
  AOI22_X1 U20906 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17777) );
  INV_X1 U20907 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17775) );
  OR2_X1 U20908 ( .A1(n18545), .A2(n17775), .ZN(n17776) );
  NAND4_X1 U20909 ( .A1(n17779), .A2(n17778), .A3(n17777), .A4(n17776), .ZN(
        n17792) );
  INV_X1 U20910 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17781) );
  OAI22_X1 U20911 ( .A1(n18541), .A2(n17781), .B1(n18539), .B2(n17780), .ZN(
        n17791) );
  AOI22_X1 U20912 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17789) );
  AOI22_X1 U20913 ( .A1(n17783), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17788) );
  AOI22_X1 U20914 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17784), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17787) );
  NAND2_X1 U20915 ( .A1(n17785), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n17786) );
  NAND4_X1 U20916 ( .A1(n17789), .A2(n17788), .A3(n17787), .A4(n17786), .ZN(
        n17790) );
  OR3_X1 U20917 ( .A1(n17792), .A2(n17791), .A3(n17790), .ZN(n18494) );
  NAND2_X1 U20918 ( .A1(n18497), .A2(n18494), .ZN(n18493) );
  NOR2_X1 U20919 ( .A1(n18493), .A2(n17793), .ZN(n18490) );
  AOI21_X1 U20920 ( .B1(n17793), .B2(n18493), .A(n18490), .ZN(n17794) );
  INV_X1 U20921 ( .A(n17794), .ZN(n18609) );
  OAI22_X1 U20922 ( .A1(n17796), .A2(n17795), .B1(n18586), .B2(n18609), .ZN(
        P3_U2675) );
  INV_X1 U20923 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19874) );
  OR2_X1 U20924 ( .A1(n17797), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n17807) );
  INV_X1 U20925 ( .A(n17807), .ZN(n17798) );
  NAND2_X1 U20926 ( .A1(n17799), .A2(n17798), .ZN(n19402) );
  INV_X1 U20927 ( .A(n20015), .ZN(n17802) );
  INV_X1 U20928 ( .A(n17800), .ZN(n17801) );
  AOI21_X1 U20929 ( .B1(n19402), .B2(n17802), .A(n17801), .ZN(n17803) );
  AND2_X1 U20930 ( .A1(n19455), .A2(n17803), .ZN(n19405) );
  NOR2_X1 U20931 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20016), .ZN(
        n19454) );
  NOR3_X1 U20932 ( .A1(n19405), .A2(n19454), .A3(n19858), .ZN(n17805) );
  INV_X1 U20933 ( .A(n19408), .ZN(n19762) );
  INV_X1 U20934 ( .A(n19405), .ZN(n19413) );
  OAI22_X1 U20935 ( .A1(n19404), .A2(n20037), .B1(n12049), .B2(n20016), .ZN(
        n19407) );
  AOI21_X1 U20936 ( .B1(n19413), .B2(n19407), .A(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n17804) );
  AOI21_X1 U20937 ( .B1(n17805), .B2(n19762), .A(n17804), .ZN(P3_U2864) );
  AND2_X1 U20938 ( .A1(n17807), .A2(n17806), .ZN(n19885) );
  NAND3_X1 U20939 ( .A1(n17809), .A2(n20048), .A3(n19885), .ZN(n17808) );
  OAI21_X1 U20940 ( .B1(n17809), .B2(n19874), .A(n17808), .ZN(P3_U3284) );
  AOI22_X1 U20941 ( .A1(n17811), .A2(n20129), .B1(n20185), .B2(n17810), .ZN(
        n17824) );
  AOI22_X1 U20942 ( .A1(n20150), .A2(P2_REIP_REG_22__SCAN_IN), .B1(n20169), 
        .B2(P2_EBX_REG_22__SCAN_IN), .ZN(n17812) );
  OAI21_X1 U20943 ( .B1(n17813), .B2(n20145), .A(n17812), .ZN(n17821) );
  INV_X1 U20944 ( .A(n17814), .ZN(n17816) );
  OAI21_X1 U20945 ( .B1(n17816), .B2(n17815), .A(n20197), .ZN(n17818) );
  AOI21_X1 U20946 ( .B1(n17819), .B2(n17818), .A(n17817), .ZN(n17820) );
  AOI211_X1 U20947 ( .C1(n20187), .C2(n17822), .A(n17821), .B(n17820), .ZN(
        n17823) );
  NAND2_X1 U20948 ( .A1(n17824), .A2(n17823), .ZN(P2_U2833) );
  NAND2_X1 U20949 ( .A1(n17826), .A2(n17825), .ZN(n17830) );
  AOI21_X1 U20950 ( .B1(n17830), .B2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n21289), .ZN(n17828) );
  NOR2_X1 U20951 ( .A1(n17828), .A2(n17827), .ZN(n17829) );
  AOI21_X1 U20952 ( .B1(n17830), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n17829), .ZN(n17831) );
  AOI222_X1 U20953 ( .A1(n17832), .A2(n21392), .B1(n17832), .B2(n17831), .C1(
        n21392), .C2(n17831), .ZN(n17834) );
  AOI21_X1 U20954 ( .B1(n17834), .B2(n17833), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n17836) );
  NOR2_X1 U20955 ( .A1(n17834), .A2(n17833), .ZN(n17835) );
  OAI21_X1 U20956 ( .B1(n17836), .B2(n17835), .A(n21184), .ZN(n17845) );
  OAI21_X1 U20957 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n17837), .ZN(n17838) );
  OAI211_X1 U20958 ( .C1(n17840), .C2(n12588), .A(n17839), .B(n17838), .ZN(
        n17841) );
  NOR2_X1 U20959 ( .A1(n17842), .A2(n17841), .ZN(n17844) );
  NAND3_X1 U20960 ( .A1(n17845), .A2(n17844), .A3(n17843), .ZN(n17853) );
  NAND4_X1 U20961 ( .A1(n13119), .A2(n12924), .A3(n17847), .A4(n17846), .ZN(
        n17851) );
  OAI21_X1 U20962 ( .B1(n21759), .B2(n17849), .A(n17848), .ZN(n17850) );
  NAND2_X1 U20963 ( .A1(n17851), .A2(n17850), .ZN(n17930) );
  NOR2_X1 U20964 ( .A1(n17855), .A2(n21638), .ZN(n17933) );
  OAI211_X1 U20965 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21759), .A(n17933), 
        .B(n17852), .ZN(n17931) );
  AOI21_X1 U20966 ( .B1(n17854), .B2(n17853), .A(n17931), .ZN(n17859) );
  AOI21_X1 U20967 ( .B1(n21732), .B2(n21765), .A(n17855), .ZN(n17856) );
  INV_X1 U20968 ( .A(n17856), .ZN(n17857) );
  AOI22_X1 U20969 ( .A1(n17859), .A2(n17858), .B1(n21638), .B2(n17857), .ZN(
        P1_U3161) );
  INV_X1 U20970 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n18026) );
  NOR2_X1 U20971 ( .A1(n21139), .A2(n18026), .ZN(P1_U2905) );
  AOI21_X1 U20972 ( .B1(n20951), .B2(n14104), .A(n17860), .ZN(n17861) );
  NOR2_X1 U20973 ( .A1(n20697), .A2(n17861), .ZN(n20948) );
  INV_X1 U20974 ( .A(n20948), .ZN(n20945) );
  NOR2_X1 U20975 ( .A1(n17862), .A2(n20945), .ZN(P2_U3047) );
  AOI22_X1 U20976 ( .A1(n17870), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n17906), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n17869) );
  NAND2_X1 U20977 ( .A1(n17864), .A2(n17863), .ZN(n17865) );
  NAND2_X1 U20978 ( .A1(n17866), .A2(n17865), .ZN(n17901) );
  INV_X1 U20979 ( .A(n17867), .ZN(n21022) );
  AOI22_X1 U20980 ( .A1(n17901), .A2(n17883), .B1(n21022), .B2(n17882), .ZN(
        n17868) );
  OAI211_X1 U20981 ( .C1(n17877), .C2(n21025), .A(n17869), .B(n17868), .ZN(
        P1_U2992) );
  AOI22_X1 U20982 ( .A1(n17870), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n17906), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n17876) );
  NAND2_X1 U20983 ( .A1(n17873), .A2(n17872), .ZN(n17874) );
  XNOR2_X1 U20984 ( .A(n17871), .B(n17874), .ZN(n17908) );
  AOI22_X1 U20985 ( .A1(n17883), .A2(n17908), .B1(n21037), .B2(n17882), .ZN(
        n17875) );
  OAI211_X1 U20986 ( .C1(n17877), .C2(n21039), .A(n17876), .B(n17875), .ZN(
        P1_U2993) );
  XOR2_X1 U20987 ( .A(n17878), .B(n17879), .Z(n17916) );
  INV_X1 U20988 ( .A(n21051), .ZN(n17881) );
  AOI222_X1 U20989 ( .A1(n17916), .A2(n17883), .B1(n17882), .B2(n21106), .C1(
        n17881), .C2(n17880), .ZN(n17884) );
  NAND2_X1 U20990 ( .A1(n17906), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n17915) );
  OAI211_X1 U20991 ( .C1(n21044), .C2(n17885), .A(n17884), .B(n17915), .ZN(
        P1_U2994) );
  INV_X1 U20992 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17898) );
  NAND2_X1 U20993 ( .A1(n17887), .A2(n17917), .ZN(n17924) );
  AOI21_X1 U20994 ( .B1(n17888), .B2(n17887), .A(n17886), .ZN(n17890) );
  NOR2_X1 U20995 ( .A1(n17890), .A2(n17889), .ZN(n17918) );
  OAI211_X1 U20996 ( .C1(n17891), .C2(n17924), .A(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n17918), .ZN(n17909) );
  NAND2_X1 U20997 ( .A1(n17892), .A2(n17909), .ZN(n17903) );
  OAI22_X1 U20998 ( .A1(n21174), .A2(n17893), .B1(n21674), .B2(n17899), .ZN(
        n17895) );
  INV_X1 U20999 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17904) );
  NAND2_X1 U21000 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17910), .ZN(
        n17905) );
  AOI221_X1 U21001 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n17898), .C2(n17904), .A(
        n17905), .ZN(n17894) );
  AOI211_X1 U21002 ( .C1(n17907), .C2(n17896), .A(n17895), .B(n17894), .ZN(
        n17897) );
  OAI21_X1 U21003 ( .B1(n17898), .B2(n17903), .A(n17897), .ZN(P1_U3023) );
  INV_X1 U21004 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21673) );
  OAI22_X1 U21005 ( .A1(n21174), .A2(n21020), .B1(n21673), .B2(n17899), .ZN(
        n17900) );
  AOI21_X1 U21006 ( .B1(n17901), .B2(n17907), .A(n17900), .ZN(n17902) );
  OAI221_X1 U21007 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17905), .C1(
        n17904), .C2(n17903), .A(n17902), .ZN(P1_U3024) );
  AOI22_X1 U21008 ( .A1(n17908), .A2(n17907), .B1(n17906), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n17912) );
  OAI21_X1 U21009 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17910), .A(
        n17909), .ZN(n17911) );
  OAI211_X1 U21010 ( .C1(n21027), .C2(n21174), .A(n17912), .B(n17911), .ZN(
        P1_U3025) );
  NAND2_X1 U21011 ( .A1(n14584), .A2(n17913), .ZN(n17914) );
  AND2_X1 U21012 ( .A1(n14772), .A2(n17914), .ZN(n21105) );
  INV_X1 U21013 ( .A(n17915), .ZN(n17921) );
  INV_X1 U21014 ( .A(n17916), .ZN(n17919) );
  OAI22_X1 U21015 ( .A1(n17919), .A2(n21175), .B1(n17918), .B2(n17917), .ZN(
        n17920) );
  AOI211_X1 U21016 ( .C1(n17922), .C2(n21105), .A(n17921), .B(n17920), .ZN(
        n17923) );
  OAI21_X1 U21017 ( .B1(n17925), .B2(n17924), .A(n17923), .ZN(P1_U3026) );
  NAND4_X1 U21018 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n21641), .A4(n21759), .ZN(n17926) );
  AND2_X1 U21019 ( .A1(n17927), .A2(n17926), .ZN(n21639) );
  NAND2_X1 U21020 ( .A1(n21639), .A2(n17928), .ZN(n17929) );
  AOI22_X1 U21021 ( .A1(n13237), .A2(n17931), .B1(n17930), .B2(n17929), .ZN(
        P1_U3162) );
  OAI21_X1 U21022 ( .B1(n17933), .B2(n21530), .A(n17932), .ZN(P1_U3466) );
  NOR3_X1 U21023 ( .A1(P3_BE_N_REG_3__SCAN_IN), .A2(P3_BE_N_REG_1__SCAN_IN), 
        .A3(P3_W_R_N_REG_SCAN_IN), .ZN(n17935) );
  NOR4_X1 U21024 ( .A1(P3_BE_N_REG_0__SCAN_IN), .A2(P3_BE_N_REG_2__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17934) );
  INV_X2 U21025 ( .A(n18025), .ZN(U215) );
  NAND4_X1 U21026 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17935), .A3(n17934), .A4(
        U215), .ZN(U213) );
  INV_X1 U21027 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20234) );
  INV_X2 U21028 ( .A(U214), .ZN(n17987) );
  OAI222_X1 U21029 ( .A1(U212), .A2(n20234), .B1(n17989), .B2(n17937), .C1(
        U214), .C2(n18026), .ZN(U216) );
  AOI222_X1 U21030 ( .A1(n17979), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n17992), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n17987), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n17938) );
  INV_X1 U21031 ( .A(n17938), .ZN(U217) );
  INV_X1 U21032 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n17940) );
  AOI22_X1 U21033 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n17979), .ZN(n17939) );
  OAI21_X1 U21034 ( .B1(n17940), .B2(n17989), .A(n17939), .ZN(U218) );
  AOI222_X1 U21035 ( .A1(n17987), .A2(P1_DATAO_REG_28__SCAN_IN), .B1(n17992), 
        .B2(BUF1_REG_28__SCAN_IN), .C1(n17979), .C2(P2_DATAO_REG_28__SCAN_IN), 
        .ZN(n17941) );
  INV_X1 U21036 ( .A(n17941), .ZN(U219) );
  INV_X1 U21037 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n17943) );
  AOI22_X1 U21038 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17979), .ZN(n17942) );
  OAI21_X1 U21039 ( .B1(n17943), .B2(n17989), .A(n17942), .ZN(U220) );
  INV_X1 U21040 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n17945) );
  AOI22_X1 U21041 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17979), .ZN(n17944) );
  OAI21_X1 U21042 ( .B1(n17945), .B2(n17989), .A(n17944), .ZN(U221) );
  INV_X1 U21043 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n17947) );
  AOI22_X1 U21044 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n17979), .ZN(n17946) );
  OAI21_X1 U21045 ( .B1(n17947), .B2(n17989), .A(n17946), .ZN(U222) );
  AOI222_X1 U21046 ( .A1(n17979), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(n17992), 
        .B2(BUF1_REG_24__SCAN_IN), .C1(n17987), .C2(P1_DATAO_REG_24__SCAN_IN), 
        .ZN(n17948) );
  INV_X1 U21047 ( .A(n17948), .ZN(U223) );
  INV_X1 U21048 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n17950) );
  AOI22_X1 U21049 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17979), .ZN(n17949) );
  OAI21_X1 U21050 ( .B1(n17950), .B2(n17989), .A(n17949), .ZN(U224) );
  INV_X1 U21051 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n17952) );
  AOI22_X1 U21052 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n17979), .ZN(n17951) );
  OAI21_X1 U21053 ( .B1(n17952), .B2(n17989), .A(n17951), .ZN(U225) );
  INV_X1 U21054 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n17954) );
  AOI22_X1 U21055 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n17979), .ZN(n17953) );
  OAI21_X1 U21056 ( .B1(n17954), .B2(n17989), .A(n17953), .ZN(U226) );
  AOI22_X1 U21057 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17979), .ZN(n17955) );
  OAI21_X1 U21058 ( .B1(n17956), .B2(n17989), .A(n17955), .ZN(U227) );
  AOI22_X1 U21059 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n17979), .ZN(n17957) );
  OAI21_X1 U21060 ( .B1(n17958), .B2(n17989), .A(n17957), .ZN(U228) );
  INV_X1 U21061 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n18010) );
  OAI222_X1 U21062 ( .A1(U212), .A2(n18010), .B1(n17989), .B2(n17959), .C1(
        U214), .C2(n21119), .ZN(U229) );
  AOI222_X1 U21063 ( .A1(n17979), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n17992), 
        .B2(BUF1_REG_17__SCAN_IN), .C1(n17987), .C2(P1_DATAO_REG_17__SCAN_IN), 
        .ZN(n17960) );
  INV_X1 U21064 ( .A(n17960), .ZN(U230) );
  INV_X1 U21065 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n17962) );
  AOI22_X1 U21066 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17979), .ZN(n17961) );
  OAI21_X1 U21067 ( .B1(n17962), .B2(n17989), .A(n17961), .ZN(U231) );
  AOI22_X1 U21068 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n17979), .ZN(n17963) );
  OAI21_X1 U21069 ( .B1(n13675), .B2(n17989), .A(n17963), .ZN(U232) );
  INV_X1 U21070 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n17965) );
  AOI22_X1 U21071 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n17979), .ZN(n17964) );
  OAI21_X1 U21072 ( .B1(n17965), .B2(n17989), .A(n17964), .ZN(U233) );
  INV_X1 U21073 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n17967) );
  OAI222_X1 U21074 ( .A1(U214), .A2(n17967), .B1(n17989), .B2(n17966), .C1(
        U212), .C2(n20243), .ZN(U234) );
  INV_X1 U21075 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n17969) );
  AOI22_X1 U21076 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n17979), .ZN(n17968) );
  OAI21_X1 U21077 ( .B1(n17969), .B2(n17989), .A(n17968), .ZN(U235) );
  INV_X1 U21078 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n17971) );
  AOI22_X1 U21079 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n17979), .ZN(n17970) );
  OAI21_X1 U21080 ( .B1(n17971), .B2(n17989), .A(n17970), .ZN(U236) );
  INV_X1 U21081 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n17973) );
  AOI22_X1 U21082 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n17979), .ZN(n17972) );
  OAI21_X1 U21083 ( .B1(n17973), .B2(n17989), .A(n17972), .ZN(U237) );
  INV_X1 U21084 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n17975) );
  AOI22_X1 U21085 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n17979), .ZN(n17974) );
  OAI21_X1 U21086 ( .B1(n17975), .B2(n17989), .A(n17974), .ZN(U238) );
  INV_X1 U21087 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n17977) );
  AOI22_X1 U21088 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n17979), .ZN(n17976) );
  OAI21_X1 U21089 ( .B1(n17977), .B2(n17989), .A(n17976), .ZN(U239) );
  INV_X1 U21090 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n18000) );
  INV_X1 U21091 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n21137) );
  OAI222_X1 U21092 ( .A1(U212), .A2(n18000), .B1(n17989), .B2(n17978), .C1(
        U214), .C2(n21137), .ZN(U240) );
  AOI222_X1 U21093 ( .A1(n17979), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n17992), 
        .B2(BUF1_REG_6__SCAN_IN), .C1(n17987), .C2(P1_DATAO_REG_6__SCAN_IN), 
        .ZN(n17980) );
  INV_X1 U21094 ( .A(n17980), .ZN(U241) );
  INV_X1 U21095 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n17982) );
  AOI22_X1 U21096 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n17979), .ZN(n17981) );
  OAI21_X1 U21097 ( .B1(n17982), .B2(n17989), .A(n17981), .ZN(U242) );
  INV_X1 U21098 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n17984) );
  AOI22_X1 U21099 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n17979), .ZN(n17983) );
  OAI21_X1 U21100 ( .B1(n17984), .B2(n17989), .A(n17983), .ZN(U243) );
  AOI22_X1 U21101 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n17979), .ZN(n17985) );
  OAI21_X1 U21102 ( .B1(n17986), .B2(n17989), .A(n17985), .ZN(U244) );
  INV_X1 U21103 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n17990) );
  AOI22_X1 U21104 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n17987), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n17979), .ZN(n17988) );
  OAI21_X1 U21105 ( .B1(n17990), .B2(n17989), .A(n17988), .ZN(U245) );
  INV_X1 U21106 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n20270) );
  AOI22_X1 U21107 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n17992), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n17987), .ZN(n17991) );
  OAI21_X1 U21108 ( .B1(n20270), .B2(U212), .A(n17991), .ZN(U246) );
  INV_X1 U21109 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n17994) );
  AOI22_X1 U21110 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n17992), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n17987), .ZN(n17993) );
  OAI21_X1 U21111 ( .B1(n17994), .B2(U212), .A(n17993), .ZN(U247) );
  AOI22_X1 U21112 ( .A1(n18025), .A2(n17994), .B1(n13564), .B2(U215), .ZN(U251) );
  AOI22_X1 U21113 ( .A1(n18016), .A2(n20270), .B1(n13462), .B2(U215), .ZN(U252) );
  INV_X1 U21114 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n17995) );
  AOI22_X1 U21115 ( .A1(n18025), .A2(n17995), .B1(n19424), .B2(U215), .ZN(U253) );
  INV_X1 U21116 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n17996) );
  AOI22_X1 U21117 ( .A1(n18025), .A2(n17996), .B1(n19430), .B2(U215), .ZN(U254) );
  INV_X1 U21118 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n17997) );
  AOI22_X1 U21119 ( .A1(n18025), .A2(n17997), .B1(n19435), .B2(U215), .ZN(U255) );
  INV_X1 U21120 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n17998) );
  AOI22_X1 U21121 ( .A1(n18016), .A2(n17998), .B1(n19439), .B2(U215), .ZN(U256) );
  INV_X1 U21122 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n17999) );
  AOI22_X1 U21123 ( .A1(n18025), .A2(n17999), .B1(n13243), .B2(U215), .ZN(U257) );
  AOI22_X1 U21124 ( .A1(n18016), .A2(n18000), .B1(n19446), .B2(U215), .ZN(U258) );
  OAI22_X1 U21125 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n18025), .ZN(n18001) );
  INV_X1 U21126 ( .A(n18001), .ZN(U259) );
  INV_X1 U21127 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n18002) );
  AOI22_X1 U21128 ( .A1(n18016), .A2(n18002), .B1(n18778), .B2(U215), .ZN(U260) );
  INV_X1 U21129 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n18003) );
  AOI22_X1 U21130 ( .A1(n18025), .A2(n18003), .B1(n18780), .B2(U215), .ZN(U261) );
  INV_X1 U21131 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n18004) );
  AOI22_X1 U21132 ( .A1(n18025), .A2(n18004), .B1(n18782), .B2(U215), .ZN(U262) );
  INV_X1 U21133 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n18005) );
  AOI22_X1 U21134 ( .A1(n18016), .A2(n18005), .B1(n18784), .B2(U215), .ZN(U263) );
  AOI22_X1 U21135 ( .A1(n18025), .A2(n20243), .B1(n12209), .B2(U215), .ZN(U264) );
  OAI22_X1 U21136 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n18025), .ZN(n18006) );
  INV_X1 U21137 ( .A(n18006), .ZN(U265) );
  OAI22_X1 U21138 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n18025), .ZN(n18007) );
  INV_X1 U21139 ( .A(n18007), .ZN(U266) );
  INV_X1 U21140 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n18008) );
  AOI22_X1 U21141 ( .A1(n18016), .A2(n18008), .B1(n19416), .B2(U215), .ZN(U267) );
  OAI22_X1 U21142 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18025), .ZN(n18009) );
  INV_X1 U21143 ( .A(n18009), .ZN(U268) );
  AOI22_X1 U21144 ( .A1(n18016), .A2(n18010), .B1(n16860), .B2(U215), .ZN(U269) );
  OAI22_X1 U21145 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18025), .ZN(n18011) );
  INV_X1 U21146 ( .A(n18011), .ZN(U270) );
  OAI22_X1 U21147 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n18025), .ZN(n18012) );
  INV_X1 U21148 ( .A(n18012), .ZN(U271) );
  OAI22_X1 U21149 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n18016), .ZN(n18013) );
  INV_X1 U21150 ( .A(n18013), .ZN(U272) );
  INV_X1 U21151 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n18014) );
  AOI22_X1 U21152 ( .A1(n18025), .A2(n18014), .B1(n16827), .B2(U215), .ZN(U273) );
  OAI22_X1 U21153 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18016), .ZN(n18015) );
  INV_X1 U21154 ( .A(n18015), .ZN(U274) );
  OAI22_X1 U21155 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18016), .ZN(n18017) );
  INV_X1 U21156 ( .A(n18017), .ZN(U275) );
  INV_X1 U21157 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n18019) );
  AOI22_X1 U21158 ( .A1(n18025), .A2(n18019), .B1(n18018), .B2(U215), .ZN(U276) );
  OAI22_X1 U21159 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18025), .ZN(n18020) );
  INV_X1 U21160 ( .A(n18020), .ZN(U277) );
  OAI22_X1 U21161 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18025), .ZN(n18021) );
  INV_X1 U21162 ( .A(n18021), .ZN(U278) );
  AOI22_X1 U21163 ( .A1(n18025), .A2(n20238), .B1(n16778), .B2(U215), .ZN(U279) );
  OAI22_X1 U21164 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18025), .ZN(n18023) );
  INV_X1 U21165 ( .A(n18023), .ZN(U280) );
  AOI22_X1 U21166 ( .A1(n18025), .A2(n18024), .B1(n16771), .B2(U215), .ZN(U281) );
  AOI22_X1 U21167 ( .A1(n18025), .A2(n20234), .B1(n16767), .B2(U215), .ZN(U282) );
  INV_X1 U21168 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n18680) );
  AOI222_X1 U21169 ( .A1(n18026), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20234), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n18680), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n18027) );
  INV_X2 U21170 ( .A(n18029), .ZN(n18028) );
  INV_X1 U21171 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19962) );
  INV_X1 U21172 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20864) );
  AOI22_X1 U21173 ( .A1(n18028), .A2(n19962), .B1(n20864), .B2(n18029), .ZN(
        U347) );
  INV_X1 U21174 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20862) );
  AOI22_X1 U21175 ( .A1(n18028), .A2(n19960), .B1(n20862), .B2(n18029), .ZN(
        U348) );
  INV_X1 U21176 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19957) );
  INV_X1 U21177 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20860) );
  AOI22_X1 U21178 ( .A1(n18028), .A2(n19957), .B1(n20860), .B2(n18029), .ZN(
        U349) );
  INV_X1 U21179 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19956) );
  INV_X1 U21180 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20859) );
  AOI22_X1 U21181 ( .A1(n18028), .A2(n19956), .B1(n20859), .B2(n18029), .ZN(
        U350) );
  INV_X1 U21182 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19954) );
  INV_X1 U21183 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20857) );
  AOI22_X1 U21184 ( .A1(n18028), .A2(n19954), .B1(n20857), .B2(n18029), .ZN(
        U351) );
  INV_X1 U21185 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19951) );
  INV_X1 U21186 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20855) );
  AOI22_X1 U21187 ( .A1(n18028), .A2(n19951), .B1(n20855), .B2(n18029), .ZN(
        U352) );
  INV_X1 U21188 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19950) );
  INV_X1 U21189 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20854) );
  AOI22_X1 U21190 ( .A1(n18028), .A2(n19950), .B1(n20854), .B2(n18029), .ZN(
        U353) );
  INV_X1 U21191 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19948) );
  AOI22_X1 U21192 ( .A1(n18028), .A2(n19948), .B1(n20852), .B2(n18029), .ZN(
        U354) );
  INV_X1 U21193 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n20001) );
  INV_X1 U21194 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20901) );
  AOI22_X1 U21195 ( .A1(n18028), .A2(n20001), .B1(n20901), .B2(n18029), .ZN(
        U355) );
  INV_X1 U21196 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19998) );
  INV_X1 U21197 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20897) );
  AOI22_X1 U21198 ( .A1(n18028), .A2(n19998), .B1(n20897), .B2(n18029), .ZN(
        U356) );
  INV_X1 U21199 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19997) );
  INV_X1 U21200 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20895) );
  AOI22_X1 U21201 ( .A1(n18028), .A2(n19997), .B1(n20895), .B2(n18029), .ZN(
        U357) );
  INV_X1 U21202 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19995) );
  INV_X1 U21203 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20893) );
  AOI22_X1 U21204 ( .A1(n18028), .A2(n19995), .B1(n20893), .B2(n18029), .ZN(
        U358) );
  INV_X1 U21205 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19994) );
  INV_X1 U21206 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20892) );
  AOI22_X1 U21207 ( .A1(n18028), .A2(n19994), .B1(n20892), .B2(n18029), .ZN(
        U359) );
  INV_X1 U21208 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19992) );
  INV_X1 U21209 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20890) );
  AOI22_X1 U21210 ( .A1(n18028), .A2(n19992), .B1(n20890), .B2(n18029), .ZN(
        U360) );
  INV_X1 U21211 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19990) );
  INV_X1 U21212 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20888) );
  AOI22_X1 U21213 ( .A1(n18028), .A2(n19990), .B1(n20888), .B2(n18029), .ZN(
        U361) );
  INV_X1 U21214 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19987) );
  INV_X1 U21215 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20887) );
  AOI22_X1 U21216 ( .A1(n18028), .A2(n19987), .B1(n20887), .B2(n18029), .ZN(
        U362) );
  INV_X1 U21217 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19986) );
  INV_X1 U21218 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20885) );
  AOI22_X1 U21219 ( .A1(n18028), .A2(n19986), .B1(n20885), .B2(n18029), .ZN(
        U363) );
  INV_X1 U21220 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19983) );
  INV_X1 U21221 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20884) );
  AOI22_X1 U21222 ( .A1(n18028), .A2(n19983), .B1(n20884), .B2(n18029), .ZN(
        U364) );
  INV_X1 U21223 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19946) );
  INV_X1 U21224 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20850) );
  AOI22_X1 U21225 ( .A1(n18028), .A2(n19946), .B1(n20850), .B2(n18029), .ZN(
        U365) );
  INV_X1 U21226 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19982) );
  INV_X1 U21227 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20882) );
  AOI22_X1 U21228 ( .A1(n18028), .A2(n19982), .B1(n20882), .B2(n18029), .ZN(
        U366) );
  INV_X1 U21229 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19979) );
  INV_X1 U21230 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20881) );
  AOI22_X1 U21231 ( .A1(n18028), .A2(n19979), .B1(n20881), .B2(n18029), .ZN(
        U367) );
  INV_X1 U21232 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20879) );
  AOI22_X1 U21233 ( .A1(n18028), .A2(n19978), .B1(n20879), .B2(n18029), .ZN(
        U368) );
  INV_X1 U21234 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20878) );
  AOI22_X1 U21235 ( .A1(n18028), .A2(n19975), .B1(n20878), .B2(n18029), .ZN(
        U369) );
  INV_X1 U21236 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19974) );
  INV_X1 U21237 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20876) );
  AOI22_X1 U21238 ( .A1(n18028), .A2(n19974), .B1(n20876), .B2(n18029), .ZN(
        U370) );
  INV_X1 U21239 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19972) );
  INV_X1 U21240 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20874) );
  AOI22_X1 U21241 ( .A1(n18028), .A2(n19972), .B1(n20874), .B2(n18029), .ZN(
        U371) );
  INV_X1 U21242 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19969) );
  INV_X1 U21243 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20872) );
  AOI22_X1 U21244 ( .A1(n18028), .A2(n19969), .B1(n20872), .B2(n18029), .ZN(
        U372) );
  INV_X1 U21245 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19968) );
  INV_X1 U21246 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20870) );
  AOI22_X1 U21247 ( .A1(n18028), .A2(n19968), .B1(n20870), .B2(n18029), .ZN(
        U373) );
  INV_X1 U21248 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19966) );
  INV_X1 U21249 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20868) );
  AOI22_X1 U21250 ( .A1(n18028), .A2(n19966), .B1(n20868), .B2(n18029), .ZN(
        U374) );
  INV_X1 U21251 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19964) );
  INV_X1 U21252 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20866) );
  AOI22_X1 U21253 ( .A1(n18028), .A2(n19964), .B1(n20866), .B2(n18029), .ZN(
        U375) );
  INV_X1 U21254 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19944) );
  INV_X1 U21255 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20848) );
  AOI22_X1 U21256 ( .A1(n18028), .A2(n19944), .B1(n20848), .B2(n18029), .ZN(
        U376) );
  INV_X1 U21257 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n18031) );
  NAND3_X1 U21258 ( .A1(n19943), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n18030) );
  OR2_X1 U21259 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n19931) );
  NAND2_X1 U21260 ( .A1(n18030), .A2(n19931), .ZN(n20014) );
  OAI21_X1 U21261 ( .B1(n19930), .B2(n18031), .A(n20011), .ZN(P3_U2633) );
  NAND2_X1 U21262 ( .A1(n20047), .A2(n20016), .ZN(n18035) );
  INV_X1 U21263 ( .A(n18032), .ZN(n18040) );
  OAI21_X1 U21264 ( .B1(n18040), .B2(n18033), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n18034) );
  OAI21_X1 U21265 ( .B1(n18035), .B2(n19920), .A(n18034), .ZN(P3_U2634) );
  AOI22_X1 U21266 ( .A1(P3_D_C_N_REG_SCAN_IN), .A2(n20026), .B1(n19928), .B2(
        n19930), .ZN(n18036) );
  OAI21_X1 U21267 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n20026), .A(n18036), 
        .ZN(P3_U2635) );
  OAI21_X1 U21268 ( .B1(n19928), .B2(BS16), .A(n20014), .ZN(n20012) );
  OAI21_X1 U21269 ( .B1(n20014), .B2(n18037), .A(n20012), .ZN(P3_U2636) );
  NOR3_X1 U21270 ( .A1(n18040), .A2(n18039), .A3(n18038), .ZN(n19871) );
  NOR2_X1 U21271 ( .A1(n19871), .A2(n19914), .ZN(n20028) );
  OAI21_X1 U21272 ( .B1(n20028), .B2(n19401), .A(n18041), .ZN(P3_U2637) );
  NOR4_X1 U21273 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18045) );
  NOR4_X1 U21274 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18044) );
  NOR4_X1 U21275 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18043) );
  NOR4_X1 U21276 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18042) );
  NAND4_X1 U21277 ( .A1(n18045), .A2(n18044), .A3(n18043), .A4(n18042), .ZN(
        n18051) );
  NOR4_X1 U21278 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n18049) );
  AOI211_X1 U21279 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_21__SCAN_IN), .B(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18048) );
  NOR4_X1 U21280 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18047) );
  NOR4_X1 U21281 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n18046) );
  NAND4_X1 U21282 ( .A1(n18049), .A2(n18048), .A3(n18047), .A4(n18046), .ZN(
        n18050) );
  NOR2_X1 U21283 ( .A1(n18051), .A2(n18050), .ZN(n20025) );
  INV_X1 U21284 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20007) );
  NOR3_X1 U21285 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18053) );
  OAI21_X1 U21286 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18053), .A(n20025), .ZN(
        n18052) );
  OAI21_X1 U21287 ( .B1(n20025), .B2(n20007), .A(n18052), .ZN(P3_U2638) );
  INV_X1 U21288 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20013) );
  AOI21_X1 U21289 ( .B1(n20018), .B2(n20013), .A(n18053), .ZN(n18054) );
  INV_X1 U21290 ( .A(n20025), .ZN(n20020) );
  AOI22_X1 U21291 ( .A1(n20025), .A2(n18054), .B1(n20004), .B2(n20020), .ZN(
        P3_U2639) );
  INV_X1 U21292 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19981) );
  INV_X1 U21293 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19963) );
  INV_X1 U21294 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19952) );
  NAND2_X1 U21295 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n18431) );
  NOR2_X1 U21296 ( .A1(n19947), .A2(n18431), .ZN(n18391) );
  NAND2_X1 U21297 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n18391), .ZN(n18376) );
  NOR2_X1 U21298 ( .A1(n19952), .A2(n18376), .ZN(n18374) );
  NAND4_X1 U21299 ( .A1(n18374), .A2(P3_REIP_REG_8__SCAN_IN), .A3(
        P3_REIP_REG_7__SCAN_IN), .A4(P3_REIP_REG_6__SCAN_IN), .ZN(n18311) );
  NAND2_X1 U21300 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n18320) );
  NOR3_X1 U21301 ( .A1(n19963), .A2(n18311), .A3(n18320), .ZN(n18291) );
  NAND2_X1 U21302 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18291), .ZN(n18273) );
  NOR2_X1 U21303 ( .A1(n19967), .A2(n18273), .ZN(n18260) );
  NAND2_X1 U21304 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n18260), .ZN(n18261) );
  NAND2_X1 U21305 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n18238) );
  NOR2_X1 U21306 ( .A1(n18261), .A2(n18238), .ZN(n18224) );
  NAND2_X1 U21307 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n18224), .ZN(n18222) );
  NAND2_X1 U21308 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n18198) );
  NOR3_X1 U21309 ( .A1(n19981), .A2(n18222), .A3(n18198), .ZN(n18169) );
  NAND4_X1 U21310 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .A3(n18169), .A4(P3_REIP_REG_22__SCAN_IN), .ZN(n18072) );
  NOR2_X1 U21311 ( .A1(n18408), .A2(n18072), .ZN(n18145) );
  NAND2_X1 U21312 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n18145), .ZN(n18137) );
  NAND2_X1 U21313 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n18071) );
  NOR2_X1 U21314 ( .A1(n18137), .A2(n18071), .ZN(n18111) );
  NAND4_X1 U21315 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n18111), .ZN(n18075) );
  NOR3_X1 U21316 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n17557), .A3(n18075), 
        .ZN(n18055) );
  AOI21_X1 U21317 ( .B1(n18392), .B2(P3_EBX_REG_31__SCAN_IN), .A(n18055), .ZN(
        n18080) );
  INV_X1 U21318 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n18577) );
  NAND2_X1 U21319 ( .A1(n18419), .A2(n18577), .ZN(n18415) );
  INV_X1 U21320 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n18337) );
  NAND2_X1 U21321 ( .A1(n18338), .A2(n18337), .ZN(n18334) );
  INV_X1 U21322 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n18307) );
  NAND2_X1 U21323 ( .A1(n18312), .A2(n18307), .ZN(n18306) );
  INV_X1 U21324 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n18285) );
  NAND2_X1 U21325 ( .A1(n18233), .A2(n18227), .ZN(n18226) );
  INV_X1 U21326 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n18537) );
  INV_X1 U21327 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n18162) );
  NAND2_X1 U21328 ( .A1(n18171), .A2(n18162), .ZN(n18161) );
  INV_X1 U21329 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n18098) );
  NAND2_X1 U21330 ( .A1(n18102), .A2(n18098), .ZN(n18082) );
  NOR2_X1 U21331 ( .A1(n18436), .A2(n18082), .ZN(n18087) );
  INV_X1 U21332 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n18453) );
  INV_X1 U21333 ( .A(n18056), .ZN(n18105) );
  INV_X1 U21334 ( .A(n18057), .ZN(n18069) );
  AOI21_X1 U21335 ( .B1(n13198), .B2(n18069), .A(n18058), .ZN(n18796) );
  INV_X1 U21336 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18173) );
  NOR2_X1 U21337 ( .A1(n19125), .A2(n18848), .ZN(n18065) );
  NAND2_X1 U21338 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18065), .ZN(
        n18060) );
  INV_X1 U21339 ( .A(n18059), .ZN(n18067) );
  AOI21_X1 U21340 ( .B1(n18173), .B2(n18060), .A(n18067), .ZN(n18846) );
  INV_X2 U21341 ( .A(n18064), .ZN(n18339) );
  NOR2_X1 U21342 ( .A1(n19125), .A2(n18890), .ZN(n18881) );
  NAND2_X1 U21343 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18881), .ZN(
        n18211) );
  INV_X1 U21344 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18946) );
  NOR2_X1 U21345 ( .A1(n19125), .A2(n18922), .ZN(n18923) );
  INV_X1 U21346 ( .A(n18923), .ZN(n18246) );
  NOR2_X1 U21347 ( .A1(n18946), .A2(n18246), .ZN(n18245) );
  NAND2_X1 U21348 ( .A1(n18245), .A2(n18324), .ZN(n18253) );
  NOR2_X1 U21349 ( .A1(n18211), .A2(n18253), .ZN(n18199) );
  AND2_X1 U21350 ( .A1(n18199), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18061) );
  INV_X1 U21351 ( .A(n18881), .ZN(n18220) );
  NOR2_X1 U21352 ( .A1(n18892), .A2(n18220), .ZN(n18844) );
  INV_X1 U21353 ( .A(n18065), .ZN(n18062) );
  OAI21_X1 U21354 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18844), .A(
        n18062), .ZN(n18063) );
  INV_X1 U21355 ( .A(n18063), .ZN(n18873) );
  XNOR2_X1 U21356 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n18065), .ZN(
        n18856) );
  INV_X1 U21357 ( .A(n18856), .ZN(n18181) );
  NOR2_X1 U21358 ( .A1(n18179), .A2(n18339), .ZN(n18168) );
  NOR2_X1 U21359 ( .A1(n18846), .A2(n18168), .ZN(n18167) );
  OAI21_X1 U21360 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18067), .A(
        n18066), .ZN(n18068) );
  INV_X1 U21361 ( .A(n18068), .ZN(n18833) );
  NOR2_X1 U21362 ( .A1(n18157), .A2(n18339), .ZN(n18149) );
  NOR2_X1 U21363 ( .A1(n18151), .A2(n18149), .ZN(n18150) );
  OAI21_X1 U21364 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18070), .A(
        n18069), .ZN(n18812) );
  INV_X1 U21365 ( .A(n18812), .ZN(n18134) );
  NOR2_X1 U21366 ( .A1(n18112), .A2(n18339), .ZN(n18103) );
  NOR2_X1 U21367 ( .A1(n18105), .A2(n18103), .ZN(n18104) );
  NOR2_X1 U21368 ( .A1(n18104), .A2(n18339), .ZN(n18090) );
  NOR3_X1 U21369 ( .A1(n18084), .A2(n18083), .A3(n18247), .ZN(n18078) );
  NAND3_X1 U21370 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n18074) );
  INV_X1 U21371 ( .A(n18071), .ZN(n18073) );
  NOR2_X1 U21372 ( .A1(n18072), .A2(n18385), .ZN(n18146) );
  AND2_X1 U21373 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n18146), .ZN(n18141) );
  NOR2_X1 U21374 ( .A1(n18432), .A2(n18385), .ZN(n18438) );
  AOI21_X1 U21375 ( .B1(n18073), .B2(n18141), .A(n18438), .ZN(n18129) );
  AOI21_X1 U21376 ( .B1(n18432), .B2(n18074), .A(n18129), .ZN(n18101) );
  NOR2_X1 U21377 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n18075), .ZN(n18086) );
  INV_X1 U21378 ( .A(n18086), .ZN(n18076) );
  AOI21_X1 U21379 ( .B1(n18101), .B2(n18076), .A(n20000), .ZN(n18077) );
  OAI211_X1 U21380 ( .C1(n18081), .C2(n18435), .A(n18080), .B(n18079), .ZN(
        P3_U2640) );
  NAND2_X1 U21381 ( .A1(n18416), .A2(n18082), .ZN(n18096) );
  OAI22_X1 U21382 ( .A1(n18101), .A2(n17557), .B1(n10296), .B2(n18435), .ZN(
        n18085) );
  OAI21_X1 U21383 ( .B1(n18392), .B2(n18087), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n18088) );
  AOI211_X1 U21384 ( .C1(n18092), .C2(n18090), .A(n18091), .B(n19923), .ZN(
        n18095) );
  NAND3_X1 U21385 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n18111), .ZN(n18093) );
  OAI22_X1 U21386 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n18093), .B1(n12123), 
        .B2(n18435), .ZN(n18094) );
  AOI211_X1 U21387 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n18392), .A(n18095), .B(
        n18094), .ZN(n18100) );
  INV_X1 U21388 ( .A(n18096), .ZN(n18097) );
  OAI21_X1 U21389 ( .B1(n18102), .B2(n18098), .A(n18097), .ZN(n18099) );
  OAI211_X1 U21390 ( .C1(n18101), .C2(n17567), .A(n18100), .B(n18099), .ZN(
        P3_U2642) );
  AOI22_X1 U21391 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18129), .B1(n18392), 
        .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n18110) );
  AOI22_X1 U21392 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .B1(n17587), .B2(n13202), .ZN(n18108) );
  AOI211_X1 U21393 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n18118), .A(n18102), .B(
        n18436), .ZN(n18107) );
  AOI211_X1 U21394 ( .C1(n18105), .C2(n18103), .A(n18104), .B(n19923), .ZN(
        n18106) );
  OAI211_X1 U21395 ( .C1(n13201), .C2(n18435), .A(n18110), .B(n18109), .ZN(
        P3_U2643) );
  INV_X1 U21396 ( .A(n18111), .ZN(n18121) );
  AOI211_X1 U21397 ( .C1(n18114), .C2(n18113), .A(n18112), .B(n19923), .ZN(
        n18117) );
  OAI22_X1 U21398 ( .A1(n18115), .A2(n18435), .B1(n18437), .B2(n18447), .ZN(
        n18116) );
  AOI211_X1 U21399 ( .C1(n18129), .C2(P3_REIP_REG_27__SCAN_IN), .A(n18117), 
        .B(n18116), .ZN(n18120) );
  OAI211_X1 U21400 ( .C1(n18122), .C2(n18447), .A(n18416), .B(n18118), .ZN(
        n18119) );
  OAI211_X1 U21401 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n18121), .A(n18120), 
        .B(n18119), .ZN(P3_U2644) );
  INV_X1 U21402 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19991) );
  INV_X1 U21403 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19993) );
  OAI21_X1 U21404 ( .B1(n19991), .B2(n18137), .A(n19993), .ZN(n18128) );
  AOI211_X1 U21405 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n18123), .A(n18122), .B(
        n18436), .ZN(n18127) );
  AOI211_X1 U21406 ( .C1(n18796), .C2(n18125), .A(n18124), .B(n19923), .ZN(
        n18126) );
  AOI211_X1 U21407 ( .C1(n18129), .C2(n18128), .A(n18127), .B(n18126), .ZN(
        n18131) );
  NAND2_X1 U21408 ( .A1(n18392), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n18130) );
  OAI211_X1 U21409 ( .C1(n18435), .C2(n13198), .A(n18131), .B(n18130), .ZN(
        P3_U2645) );
  INV_X1 U21410 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18144) );
  NOR2_X1 U21411 ( .A1(n18135), .A2(n18436), .ZN(n18147) );
  AOI211_X1 U21412 ( .C1(n18134), .C2(n18133), .A(n18132), .B(n19923), .ZN(
        n18139) );
  AOI21_X1 U21413 ( .B1(n18416), .B2(n18135), .A(n18392), .ZN(n18136) );
  OAI22_X1 U21414 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n18137), .B1(n18136), 
        .B2(n18140), .ZN(n18138) );
  AOI211_X1 U21415 ( .C1(n18147), .C2(n18140), .A(n18139), .B(n18138), .ZN(
        n18143) );
  OR3_X1 U21416 ( .A1(n18438), .A2(n18141), .A3(n19991), .ZN(n18142) );
  OAI211_X1 U21417 ( .C1(n18435), .C2(n18144), .A(n18143), .B(n18142), .ZN(
        P3_U2646) );
  AOI22_X1 U21418 ( .A1(n18392), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n18145), 
        .B2(n19989), .ZN(n18155) );
  NOR2_X1 U21419 ( .A1(n18438), .A2(n18146), .ZN(n18160) );
  INV_X1 U21420 ( .A(n18147), .ZN(n18148) );
  AOI21_X1 U21421 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18161), .A(n18148), .ZN(
        n18153) );
  AOI211_X1 U21422 ( .C1(n18151), .C2(n18149), .A(n18150), .B(n19923), .ZN(
        n18152) );
  AOI211_X1 U21423 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n18160), .A(n18153), 
        .B(n18152), .ZN(n18154) );
  OAI211_X1 U21424 ( .C1(n18156), .C2(n18435), .A(n18155), .B(n18154), .ZN(
        P3_U2647) );
  AOI22_X1 U21425 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18402), .B1(
        n18392), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n18166) );
  AOI211_X1 U21426 ( .C1(n18833), .C2(n18158), .A(n18157), .B(n19923), .ZN(
        n18159) );
  AOI21_X1 U21427 ( .B1(n18160), .B2(P3_REIP_REG_23__SCAN_IN), .A(n18159), 
        .ZN(n18165) );
  OAI211_X1 U21428 ( .C1(n18171), .C2(n18162), .A(n18416), .B(n18161), .ZN(
        n18164) );
  INV_X1 U21429 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19984) );
  NOR2_X1 U21430 ( .A1(n19984), .A2(n19985), .ZN(n18170) );
  INV_X1 U21431 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19988) );
  NAND4_X1 U21432 ( .A1(n18432), .A2(n18169), .A3(n18170), .A4(n19988), .ZN(
        n18163) );
  NAND4_X1 U21433 ( .A1(n18166), .A2(n18165), .A3(n18164), .A4(n18163), .ZN(
        P3_U2648) );
  OAI21_X1 U21434 ( .B1(n18408), .B2(n18169), .A(n18441), .ZN(n18184) );
  INV_X1 U21435 ( .A(n18184), .ZN(n18197) );
  AOI211_X1 U21436 ( .C1(n18846), .C2(n18168), .A(n18167), .B(n19923), .ZN(
        n18177) );
  NAND2_X1 U21437 ( .A1(n18432), .A2(n18169), .ZN(n18188) );
  AOI211_X1 U21438 ( .C1(n19984), .C2(n19985), .A(n18170), .B(n18188), .ZN(
        n18176) );
  AOI211_X1 U21439 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n18185), .A(n18171), .B(
        n18436), .ZN(n18175) );
  OAI22_X1 U21440 ( .A1(n18173), .A2(n18435), .B1(n18437), .B2(n18172), .ZN(
        n18174) );
  NOR4_X1 U21441 ( .A1(n18177), .A2(n18176), .A3(n18175), .A4(n18174), .ZN(
        n18178) );
  OAI21_X1 U21442 ( .B1(n19985), .B2(n18197), .A(n18178), .ZN(P3_U2649) );
  AOI211_X1 U21443 ( .C1(n18181), .C2(n18180), .A(n18179), .B(n19923), .ZN(
        n18183) );
  INV_X1 U21444 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18859) );
  OAI22_X1 U21445 ( .A1(n18859), .A2(n18435), .B1(n18437), .B2(n18537), .ZN(
        n18182) );
  AOI211_X1 U21446 ( .C1(n18184), .C2(P3_REIP_REG_21__SCAN_IN), .A(n18183), 
        .B(n18182), .ZN(n18187) );
  OAI211_X1 U21447 ( .C1(n18191), .C2(n18537), .A(n18416), .B(n18185), .ZN(
        n18186) );
  OAI211_X1 U21448 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n18188), .A(n18187), 
        .B(n18186), .ZN(P3_U2650) );
  AOI22_X1 U21449 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18402), .B1(
        n18392), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n18196) );
  NOR4_X1 U21450 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n18408), .A3(n18222), 
        .A4(n18198), .ZN(n18194) );
  AOI211_X1 U21451 ( .C1(n18873), .C2(n18190), .A(n18189), .B(n19923), .ZN(
        n18193) );
  AOI211_X1 U21452 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n18204), .A(n18191), .B(
        n18436), .ZN(n18192) );
  NOR3_X1 U21453 ( .A1(n18194), .A2(n18193), .A3(n18192), .ZN(n18195) );
  OAI211_X1 U21454 ( .C1(n19981), .C2(n18197), .A(n18196), .B(n18195), .ZN(
        P3_U2651) );
  INV_X1 U21455 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18208) );
  AOI21_X1 U21456 ( .B1(n18432), .B2(n18222), .A(n18385), .ZN(n18232) );
  INV_X1 U21457 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19980) );
  NOR2_X1 U21458 ( .A1(n18408), .A2(n18222), .ZN(n18209) );
  OAI211_X1 U21459 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n18209), .B(n18198), .ZN(n18202) );
  AOI21_X1 U21460 ( .B1(n18208), .B2(n18211), .A(n18844), .ZN(n18882) );
  NOR2_X1 U21461 ( .A1(n18199), .A2(n18339), .ZN(n18213) );
  AOI21_X1 U21462 ( .B1(n18882), .B2(n18213), .A(n19923), .ZN(n18200) );
  OAI21_X1 U21463 ( .B1(n18882), .B2(n18213), .A(n18200), .ZN(n18201) );
  OAI211_X1 U21464 ( .C1(n18232), .C2(n19980), .A(n18202), .B(n18201), .ZN(
        n18203) );
  AOI211_X1 U21465 ( .C1(n18392), .C2(P3_EBX_REG_19__SCAN_IN), .A(n19302), .B(
        n18203), .ZN(n18207) );
  OAI211_X1 U21466 ( .C1(n18210), .C2(n18205), .A(n18416), .B(n18204), .ZN(
        n18206) );
  OAI211_X1 U21467 ( .C1(n18435), .C2(n18208), .A(n18207), .B(n18206), .ZN(
        P3_U2652) );
  INV_X1 U21468 ( .A(n18209), .ZN(n18219) );
  INV_X1 U21469 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19977) );
  AOI211_X1 U21470 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n18226), .A(n18210), .B(
        n18436), .ZN(n18217) );
  INV_X1 U21471 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18899) );
  INV_X1 U21472 ( .A(n19302), .ZN(n19349) );
  OAI21_X1 U21473 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18881), .A(
        n18211), .ZN(n18896) );
  INV_X1 U21474 ( .A(n18896), .ZN(n18214) );
  NOR2_X1 U21475 ( .A1(n18406), .A2(n19923), .ZN(n18389) );
  AOI221_X1 U21476 ( .B1(n18220), .B2(n18214), .C1(n18253), .C2(n18214), .A(
        n19923), .ZN(n18212) );
  OAI22_X1 U21477 ( .A1(n18214), .A2(n18213), .B1(n18389), .B2(n18212), .ZN(
        n18215) );
  OAI211_X1 U21478 ( .C1(n18899), .C2(n18435), .A(n19349), .B(n18215), .ZN(
        n18216) );
  AOI211_X1 U21479 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n18392), .A(n18217), .B(
        n18216), .ZN(n18218) );
  OAI221_X1 U21480 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n18219), .C1(n19977), 
        .C2(n18232), .A(n18218), .ZN(P3_U2653) );
  INV_X1 U21481 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19976) );
  NOR2_X1 U21482 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19125), .ZN(
        n18340) );
  AOI21_X1 U21483 ( .B1(n18908), .B2(n18340), .A(n18339), .ZN(n18221) );
  NOR2_X1 U21484 ( .A1(n18926), .A2(n18246), .ZN(n18234) );
  OAI21_X1 U21485 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18234), .A(
        n18220), .ZN(n18909) );
  XNOR2_X1 U21486 ( .A(n18221), .B(n18909), .ZN(n18225) );
  AND2_X1 U21487 ( .A1(n18222), .A2(n18432), .ZN(n18223) );
  AOI22_X1 U21488 ( .A1(n18414), .A2(n18225), .B1(n18224), .B2(n18223), .ZN(
        n18229) );
  OAI211_X1 U21489 ( .C1(n18233), .C2(n18227), .A(n18416), .B(n18226), .ZN(
        n18228) );
  OAI211_X1 U21490 ( .C1(n18435), .C2(n10295), .A(n18229), .B(n18228), .ZN(
        n18230) );
  AOI211_X1 U21491 ( .C1(n18392), .C2(P3_EBX_REG_17__SCAN_IN), .A(n19302), .B(
        n18230), .ZN(n18231) );
  OAI21_X1 U21492 ( .B1(n18232), .B2(n19976), .A(n18231), .ZN(P3_U2654) );
  INV_X1 U21493 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18244) );
  AOI211_X1 U21494 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n18255), .A(n18233), .B(
        n18436), .ZN(n18242) );
  AOI21_X1 U21495 ( .B1(n18432), .B2(n18261), .A(n18385), .ZN(n18272) );
  INV_X1 U21496 ( .A(n18234), .ZN(n18235) );
  OAI21_X1 U21497 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18245), .A(
        n18235), .ZN(n18929) );
  NAND2_X1 U21498 ( .A1(n18406), .A2(n18253), .ZN(n18237) );
  AOI21_X1 U21499 ( .B1(n18929), .B2(n18237), .A(n19923), .ZN(n18236) );
  OAI21_X1 U21500 ( .B1(n18929), .B2(n18237), .A(n18236), .ZN(n18240) );
  NOR2_X1 U21501 ( .A1(n18408), .A2(n18261), .ZN(n18248) );
  OAI211_X1 U21502 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n18248), .B(n18238), .ZN(n18239) );
  OAI211_X1 U21503 ( .C1(n18272), .C2(n19973), .A(n18240), .B(n18239), .ZN(
        n18241) );
  AOI211_X1 U21504 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n18392), .A(n18242), .B(
        n18241), .ZN(n18243) );
  OAI211_X1 U21505 ( .C1(n18244), .C2(n18435), .A(n18243), .B(n19110), .ZN(
        P3_U2655) );
  AOI21_X1 U21506 ( .B1(n18946), .B2(n18246), .A(n18245), .ZN(n18935) );
  NOR2_X1 U21507 ( .A1(n18935), .A2(n18247), .ZN(n18254) );
  OAI21_X1 U21508 ( .B1(n18946), .B2(n18435), .A(n19349), .ZN(n18252) );
  INV_X1 U21509 ( .A(n18248), .ZN(n18250) );
  INV_X1 U21510 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19971) );
  OAI211_X1 U21511 ( .C1(n18923), .C2(n18389), .A(n18935), .B(n18276), .ZN(
        n18249) );
  OAI221_X1 U21512 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n18250), .C1(n19971), 
        .C2(n18272), .A(n18249), .ZN(n18251) );
  AOI211_X1 U21513 ( .C1(n18254), .C2(n18253), .A(n18252), .B(n18251), .ZN(
        n18257) );
  OAI211_X1 U21514 ( .C1(n18259), .C2(n18258), .A(n18416), .B(n18255), .ZN(
        n18256) );
  OAI211_X1 U21515 ( .C1(n18258), .C2(n18437), .A(n18257), .B(n18256), .ZN(
        P3_U2656) );
  INV_X1 U21516 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19970) );
  AOI211_X1 U21517 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n18282), .A(n18259), .B(
        n18436), .ZN(n18265) );
  INV_X1 U21518 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n18263) );
  NAND3_X1 U21519 ( .A1(n18261), .A2(n18432), .A3(n18260), .ZN(n18262) );
  OAI211_X1 U21520 ( .C1(n18437), .C2(n18263), .A(n19349), .B(n18262), .ZN(
        n18264) );
  AOI211_X1 U21521 ( .C1(n18402), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n18265), .B(n18264), .ZN(n18271) );
  INV_X1 U21522 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18267) );
  NOR2_X1 U21523 ( .A1(n18954), .A2(n18363), .ZN(n18970) );
  NAND2_X1 U21524 ( .A1(n18968), .A2(n18970), .ZN(n18266) );
  AOI21_X1 U21525 ( .B1(n18267), .B2(n18266), .A(n18923), .ZN(n18958) );
  INV_X1 U21526 ( .A(n18971), .ZN(n18268) );
  INV_X1 U21527 ( .A(n18340), .ZN(n18423) );
  OAI21_X1 U21528 ( .B1(n18268), .B2(n18423), .A(n18406), .ZN(n18289) );
  OAI21_X1 U21529 ( .B1(n18968), .B2(n18339), .A(n18289), .ZN(n18274) );
  AOI21_X1 U21530 ( .B1(n18958), .B2(n18274), .A(n19923), .ZN(n18269) );
  OAI21_X1 U21531 ( .B1(n18958), .B2(n18274), .A(n18269), .ZN(n18270) );
  OAI211_X1 U21532 ( .C1(n18272), .C2(n19970), .A(n18271), .B(n18270), .ZN(
        P3_U2657) );
  NOR3_X1 U21533 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n18408), .A3(n18273), 
        .ZN(n18281) );
  OAI21_X1 U21534 ( .B1(n18408), .B2(n18291), .A(n18441), .ZN(n18286) );
  NOR2_X1 U21535 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18408), .ZN(n18290) );
  OAI21_X1 U21536 ( .B1(n18286), .B2(n18290), .A(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n18279) );
  NAND2_X1 U21537 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18970), .ZN(
        n18288) );
  AOI22_X1 U21538 ( .A1(n18970), .A2(n18968), .B1(n18973), .B2(n18288), .ZN(
        n18976) );
  INV_X1 U21539 ( .A(n18976), .ZN(n18275) );
  NAND3_X1 U21540 ( .A1(n18414), .A2(n18275), .A3(n18274), .ZN(n18278) );
  OAI211_X1 U21541 ( .C1(n18389), .C2(n18973), .A(n18976), .B(n18276), .ZN(
        n18277) );
  NAND4_X1 U21542 ( .A1(n19349), .A2(n18279), .A3(n18278), .A4(n18277), .ZN(
        n18280) );
  AOI211_X1 U21543 ( .C1(n18402), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n18281), .B(n18280), .ZN(n18284) );
  OAI211_X1 U21544 ( .C1(n18287), .C2(n18285), .A(n18416), .B(n18282), .ZN(
        n18283) );
  OAI211_X1 U21545 ( .C1(n18285), .C2(n18437), .A(n18284), .B(n18283), .ZN(
        P3_U2658) );
  INV_X1 U21546 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19965) );
  INV_X1 U21547 ( .A(n18286), .ZN(n18303) );
  AOI211_X1 U21548 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n18306), .A(n18287), .B(
        n18436), .ZN(n18296) );
  OAI21_X1 U21549 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18970), .A(
        n18288), .ZN(n18984) );
  XOR2_X1 U21550 ( .A(n18984), .B(n18289), .Z(n18292) );
  AOI22_X1 U21551 ( .A1(n18414), .A2(n18292), .B1(n18291), .B2(n18290), .ZN(
        n18293) );
  OAI211_X1 U21552 ( .C1(n18437), .C2(n18294), .A(n18293), .B(n19349), .ZN(
        n18295) );
  AOI211_X1 U21553 ( .C1(n18402), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n18296), .B(n18295), .ZN(n18297) );
  OAI21_X1 U21554 ( .B1(n19965), .B2(n18303), .A(n18297), .ZN(P3_U2659) );
  INV_X1 U21555 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18310) );
  INV_X1 U21556 ( .A(n18320), .ZN(n18299) );
  NAND3_X1 U21557 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .ZN(n18298) );
  NAND2_X1 U21558 ( .A1(n18432), .A2(n18374), .ZN(n18354) );
  NOR2_X1 U21559 ( .A1(n18298), .A2(n18354), .ZN(n18332) );
  AOI21_X1 U21560 ( .B1(n18299), .B2(n18332), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n18304) );
  INV_X1 U21561 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n19010) );
  NAND2_X1 U21562 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18325), .ZN(
        n18323) );
  NOR2_X1 U21563 ( .A1(n19010), .A2(n18323), .ZN(n18313) );
  AOI21_X1 U21564 ( .B1(n18313), .B2(n18324), .A(n18339), .ZN(n18301) );
  INV_X1 U21565 ( .A(n18970), .ZN(n18300) );
  OAI21_X1 U21566 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18313), .A(
        n18300), .ZN(n18998) );
  XOR2_X1 U21567 ( .A(n18301), .B(n18998), .Z(n18302) );
  OAI22_X1 U21568 ( .A1(n18304), .A2(n18303), .B1(n19923), .B2(n18302), .ZN(
        n18305) );
  AOI211_X1 U21569 ( .C1(n18392), .C2(P3_EBX_REG_11__SCAN_IN), .A(n19302), .B(
        n18305), .ZN(n18309) );
  OAI211_X1 U21570 ( .C1(n18312), .C2(n18307), .A(n18416), .B(n18306), .ZN(
        n18308) );
  OAI211_X1 U21571 ( .C1(n18435), .C2(n18310), .A(n18309), .B(n18308), .ZN(
        P3_U2660) );
  AOI21_X1 U21572 ( .B1(n18432), .B2(n18311), .A(n18385), .ZN(n18350) );
  INV_X1 U21573 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19961) );
  AOI211_X1 U21574 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n18334), .A(n18312), .B(
        n18436), .ZN(n18319) );
  AOI21_X1 U21575 ( .B1(n19010), .B2(n18323), .A(n18313), .ZN(n19013) );
  INV_X1 U21576 ( .A(n18323), .ZN(n18314) );
  AOI21_X1 U21577 ( .B1(n18314), .B2(n18324), .A(n18339), .ZN(n18328) );
  AOI21_X1 U21578 ( .B1(n19013), .B2(n18328), .A(n19923), .ZN(n18315) );
  OAI21_X1 U21579 ( .B1(n19013), .B2(n18328), .A(n18315), .ZN(n18316) );
  OAI211_X1 U21580 ( .C1(n18437), .C2(n18317), .A(n19349), .B(n18316), .ZN(
        n18318) );
  AOI211_X1 U21581 ( .C1(n18402), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n18319), .B(n18318), .ZN(n18322) );
  OAI211_X1 U21582 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n18332), .B(n18320), .ZN(n18321) );
  OAI211_X1 U21583 ( .C1(n18350), .C2(n19961), .A(n18322), .B(n18321), .ZN(
        P3_U2661) );
  INV_X1 U21584 ( .A(n18350), .ZN(n18333) );
  INV_X1 U21585 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19959) );
  OAI21_X1 U21586 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18325), .A(
        n18323), .ZN(n19029) );
  INV_X1 U21587 ( .A(n19029), .ZN(n18329) );
  AOI21_X1 U21588 ( .B1(n18325), .B2(n18324), .A(n19029), .ZN(n18326) );
  NOR2_X1 U21589 ( .A1(n18326), .A2(n19923), .ZN(n18327) );
  OAI22_X1 U21590 ( .A1(n18329), .A2(n18328), .B1(n18389), .B2(n18327), .ZN(
        n18330) );
  OAI211_X1 U21591 ( .C1(n19025), .C2(n18435), .A(n19349), .B(n18330), .ZN(
        n18331) );
  AOI221_X1 U21592 ( .B1(n18333), .B2(P3_REIP_REG_9__SCAN_IN), .C1(n18332), 
        .C2(n19959), .A(n18331), .ZN(n18336) );
  OAI211_X1 U21593 ( .C1(n18338), .C2(n18337), .A(n18416), .B(n18334), .ZN(
        n18335) );
  OAI211_X1 U21594 ( .C1(n18337), .C2(n18437), .A(n18336), .B(n18335), .ZN(
        P3_U2662) );
  INV_X1 U21595 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19958) );
  AOI22_X1 U21596 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18402), .B1(
        n18392), .B2(P3_EBX_REG_8__SCAN_IN), .ZN(n18349) );
  AOI211_X1 U21597 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n18359), .A(n18338), .B(
        n18436), .ZN(n18347) );
  NAND2_X1 U21598 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n18355) );
  NOR3_X1 U21599 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n18355), .A3(n18354), .ZN(
        n18346) );
  AOI21_X1 U21600 ( .B1(n18341), .B2(n18340), .A(n18339), .ZN(n18343) );
  OAI21_X1 U21601 ( .B1(n18344), .B2(n18343), .A(n18414), .ZN(n18342) );
  AOI21_X1 U21602 ( .B1(n18344), .B2(n18343), .A(n18342), .ZN(n18345) );
  NOR4_X1 U21603 ( .A1(n19302), .A2(n18347), .A3(n18346), .A4(n18345), .ZN(
        n18348) );
  OAI211_X1 U21604 ( .C1(n19958), .C2(n18350), .A(n18349), .B(n18348), .ZN(
        P3_U2663) );
  OAI21_X1 U21605 ( .B1(n18374), .B2(n18408), .A(n18441), .ZN(n18380) );
  OAI21_X1 U21606 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18363), .A(
        n18406), .ZN(n18362) );
  OAI21_X1 U21607 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18352), .A(
        n18351), .ZN(n19048) );
  OAI21_X1 U21608 ( .B1(n18362), .B2(n19048), .A(n18414), .ZN(n18353) );
  AOI21_X1 U21609 ( .B1(n18362), .B2(n19048), .A(n18353), .ZN(n18358) );
  INV_X1 U21610 ( .A(n18354), .ZN(n18364) );
  OAI211_X1 U21611 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(P3_REIP_REG_6__SCAN_IN), 
        .A(n18364), .B(n18355), .ZN(n18356) );
  OAI211_X1 U21612 ( .C1(n18437), .C2(n18564), .A(n19349), .B(n18356), .ZN(
        n18357) );
  AOI211_X1 U21613 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(n18380), .A(n18358), .B(
        n18357), .ZN(n18361) );
  OAI211_X1 U21614 ( .C1(n18366), .C2(n18564), .A(n18416), .B(n18359), .ZN(
        n18360) );
  OAI211_X1 U21615 ( .C1(n18435), .C2(n19036), .A(n18361), .B(n18360), .ZN(
        P3_U2664) );
  AOI22_X1 U21616 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18402), .B1(
        n18392), .B2(P3_EBX_REG_6__SCAN_IN), .ZN(n18372) );
  NOR2_X1 U21617 ( .A1(n18362), .A2(n19923), .ZN(n18365) );
  OAI21_X1 U21618 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18373), .A(
        n18363), .ZN(n19057) );
  INV_X1 U21619 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19953) );
  AOI22_X1 U21620 ( .A1(n18365), .A2(n19057), .B1(n18364), .B2(n19953), .ZN(
        n18371) );
  AOI211_X1 U21621 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n18381), .A(n18366), .B(
        n18436), .ZN(n18369) );
  AOI211_X1 U21622 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18406), .A(
        n19057), .B(n18367), .ZN(n18368) );
  AOI211_X1 U21623 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n18380), .A(n18369), .B(
        n18368), .ZN(n18370) );
  NAND4_X1 U21624 ( .A1(n18372), .A2(n18371), .A3(n18370), .A4(n19349), .ZN(
        P3_U2665) );
  OAI22_X1 U21625 ( .A1(n19068), .A2(n18435), .B1(n18437), .B2(n18382), .ZN(
        n18379) );
  AOI21_X1 U21626 ( .B1(n19068), .B2(n18388), .A(n18373), .ZN(n19070) );
  OAI21_X1 U21627 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18388), .A(
        n18406), .ZN(n18394) );
  XOR2_X1 U21628 ( .A(n19070), .B(n18394), .Z(n18377) );
  OR2_X1 U21629 ( .A1(n18408), .A2(n18374), .ZN(n18375) );
  OAI22_X1 U21630 ( .A1(n19923), .A2(n18377), .B1(n18376), .B2(n18375), .ZN(
        n18378) );
  AOI211_X1 U21631 ( .C1(P3_REIP_REG_5__SCAN_IN), .C2(n18380), .A(n18379), .B(
        n18378), .ZN(n18384) );
  OAI211_X1 U21632 ( .C1(n18387), .C2(n18382), .A(n18416), .B(n18381), .ZN(
        n18383) );
  NAND3_X1 U21633 ( .A1(n18384), .A2(n19349), .A3(n18383), .ZN(P3_U2666) );
  INV_X1 U21634 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19949) );
  INV_X1 U21635 ( .A(n18391), .ZN(n18386) );
  AOI21_X1 U21636 ( .B1(n18432), .B2(n18386), .A(n18385), .ZN(n18407) );
  AOI211_X1 U21637 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n18415), .A(n18387), .B(
        n18436), .ZN(n18401) );
  INV_X1 U21638 ( .A(n19080), .ZN(n18393) );
  NOR2_X1 U21639 ( .A1(n19125), .A2(n18393), .ZN(n18404) );
  OAI21_X1 U21640 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18404), .A(
        n18388), .ZN(n19083) );
  INV_X1 U21641 ( .A(n18389), .ZN(n18425) );
  NOR2_X1 U21642 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n18408), .ZN(n18390) );
  AOI22_X1 U21643 ( .A1(n18392), .A2(P3_EBX_REG_4__SCAN_IN), .B1(n18391), .B2(
        n18390), .ZN(n18399) );
  INV_X1 U21644 ( .A(n19083), .ZN(n18395) );
  OR2_X1 U21645 ( .A1(n18393), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19088) );
  OAI22_X1 U21646 ( .A1(n18395), .A2(n18394), .B1(n18423), .B2(n19088), .ZN(
        n18397) );
  AOI21_X1 U21647 ( .B1(n19874), .B2(n18541), .A(n18445), .ZN(n18396) );
  AOI211_X1 U21648 ( .C1(n18397), .C2(n18414), .A(n19302), .B(n18396), .ZN(
        n18398) );
  OAI211_X1 U21649 ( .C1(n19083), .C2(n18425), .A(n18399), .B(n18398), .ZN(
        n18400) );
  AOI211_X1 U21650 ( .C1(n18402), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n18401), .B(n18400), .ZN(n18403) );
  OAI21_X1 U21651 ( .B1(n19949), .B2(n18407), .A(n18403), .ZN(P3_U2667) );
  NAND2_X1 U21652 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18421) );
  AOI21_X1 U21653 ( .B1(n19095), .B2(n18421), .A(n18404), .ZN(n19099) );
  OAI21_X1 U21654 ( .B1(n18405), .B2(n18423), .A(n18406), .ZN(n18422) );
  XNOR2_X1 U21655 ( .A(n19099), .B(n18422), .ZN(n18413) );
  AOI221_X1 U21656 ( .B1(n18408), .B2(n19947), .C1(n18431), .C2(n19947), .A(
        n18407), .ZN(n18412) );
  OAI21_X1 U21657 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18409), .A(
        n18541), .ZN(n18410) );
  OAI22_X1 U21658 ( .A1(n18435), .A2(n19095), .B1(n18445), .B2(n18410), .ZN(
        n18411) );
  AOI211_X1 U21659 ( .C1(n18414), .C2(n18413), .A(n18412), .B(n18411), .ZN(
        n18418) );
  OAI211_X1 U21660 ( .C1(n18419), .C2(n18577), .A(n18416), .B(n18415), .ZN(
        n18417) );
  OAI211_X1 U21661 ( .C1(n18577), .C2(n18437), .A(n18418), .B(n18417), .ZN(
        P3_U2668) );
  AOI211_X1 U21662 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n18420), .A(n18419), .B(
        n18436), .ZN(n18430) );
  OAI21_X1 U21663 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n18421), .ZN(n18426) );
  INV_X1 U21664 ( .A(n18426), .ZN(n19114) );
  AOI211_X1 U21665 ( .C1(n19114), .C2(n18423), .A(n19923), .B(n18422), .ZN(
        n18429) );
  INV_X1 U21666 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19945) );
  OAI22_X1 U21667 ( .A1(n19945), .A2(n18441), .B1(n18424), .B2(n18445), .ZN(
        n18428) );
  OAI22_X1 U21668 ( .A1(n18437), .A2(n9877), .B1(n18426), .B2(n18425), .ZN(
        n18427) );
  NOR4_X1 U21669 ( .A1(n18430), .A2(n18429), .A3(n18428), .A4(n18427), .ZN(
        n18434) );
  OAI211_X1 U21670 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n18432), .B(n18431), .ZN(n18433) );
  OAI211_X1 U21671 ( .C1(n18435), .C2(n18405), .A(n18434), .B(n18433), .ZN(
        P3_U2669) );
  NAND2_X1 U21672 ( .A1(n18437), .A2(n18436), .ZN(n18440) );
  INV_X1 U21673 ( .A(n18438), .ZN(n18439) );
  AOI22_X1 U21674 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n18440), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n18439), .ZN(n18444) );
  NAND3_X1 U21675 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18442), .A3(
        n18441), .ZN(n18443) );
  OAI211_X1 U21676 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18445), .A(
        n18444), .B(n18443), .ZN(P3_U2671) );
  INV_X1 U21677 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n18448) );
  NAND4_X1 U21678 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n18446)
         );
  NOR4_X1 U21679 ( .A1(n18448), .A2(n18447), .A3(n18533), .A4(n18446), .ZN(
        n18449) );
  NAND4_X1 U21680 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(P3_EBX_REG_23__SCAN_IN), .A4(n18449), .ZN(n18452) );
  NOR2_X1 U21681 ( .A1(n18453), .A2(n18452), .ZN(n18488) );
  NAND2_X1 U21682 ( .A1(n18586), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n18451) );
  NAND2_X1 U21683 ( .A1(n18488), .A2(n18576), .ZN(n18450) );
  OAI22_X1 U21684 ( .A1(n18488), .A2(n18451), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n18450), .ZN(P3_U2672) );
  NAND2_X1 U21685 ( .A1(n18453), .A2(n18452), .ZN(n18454) );
  NAND2_X1 U21686 ( .A1(n18454), .A2(n18586), .ZN(n18487) );
  INV_X1 U21687 ( .A(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18455) );
  NOR2_X1 U21688 ( .A1(n18539), .A2(n18455), .ZN(n18461) );
  AOI22_X1 U21689 ( .A1(n12008), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18459) );
  AOI22_X1 U21690 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18458) );
  AOI22_X1 U21691 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18457) );
  NAND2_X1 U21692 ( .A1(n11944), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n18456) );
  NAND4_X1 U21693 ( .A1(n18459), .A2(n18458), .A3(n18457), .A4(n18456), .ZN(
        n18460) );
  AOI211_X1 U21694 ( .C1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .C2(n18524), .A(
        n18461), .B(n18460), .ZN(n18469) );
  AOI22_X1 U21695 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18468) );
  AOI22_X1 U21696 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18467) );
  OAI22_X1 U21697 ( .A1(n18464), .A2(n18463), .B1(n17767), .B2(n18462), .ZN(
        n18465) );
  AOI21_X1 U21698 ( .B1(n9867), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(n18465), .ZN(n18466) );
  NAND4_X1 U21699 ( .A1(n18469), .A2(n18468), .A3(n18467), .A4(n18466), .ZN(
        n18489) );
  NAND2_X1 U21700 ( .A1(n18490), .A2(n18489), .ZN(n18486) );
  INV_X1 U21701 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18470) );
  OAI22_X1 U21702 ( .A1(n18471), .A2(n18541), .B1(n18539), .B2(n18470), .ZN(
        n18484) );
  AOI22_X1 U21703 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18476) );
  AOI22_X1 U21704 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18475) );
  AOI22_X1 U21705 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18474) );
  NAND2_X1 U21706 ( .A1(n9867), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n18473) );
  NAND4_X1 U21707 ( .A1(n18476), .A2(n18475), .A3(n18474), .A4(n18473), .ZN(
        n18483) );
  AOI22_X1 U21708 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n17782), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18481) );
  AOI22_X1 U21709 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18480) );
  AOI22_X1 U21710 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18479) );
  NAND2_X1 U21711 ( .A1(n17762), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n18478) );
  NAND4_X1 U21712 ( .A1(n18481), .A2(n18480), .A3(n18479), .A4(n18478), .ZN(
        n18482) );
  NOR3_X1 U21713 ( .A1(n18484), .A2(n18483), .A3(n18482), .ZN(n18485) );
  XNOR2_X1 U21714 ( .A(n18486), .B(n18485), .ZN(n18601) );
  OAI22_X1 U21715 ( .A1(n18488), .A2(n18487), .B1(n18601), .B2(n18586), .ZN(
        P3_U2673) );
  XNOR2_X1 U21716 ( .A(n18490), .B(n18489), .ZN(n18605) );
  OAI221_X1 U21717 ( .B1(n18492), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n18586), 
        .C2(n18605), .A(n18491), .ZN(P3_U2674) );
  AOI21_X1 U21718 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n18586), .A(n9748), .ZN(
        n18495) );
  OAI21_X1 U21719 ( .B1(n18497), .B2(n18494), .A(n18493), .ZN(n18613) );
  OAI22_X1 U21720 ( .A1(n18496), .A2(n18495), .B1(n18586), .B2(n18613), .ZN(
        P3_U2676) );
  AOI21_X1 U21721 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18586), .A(n18505), .ZN(
        n18500) );
  AOI21_X1 U21722 ( .B1(n18498), .B2(n18502), .A(n18497), .ZN(n18499) );
  INV_X1 U21723 ( .A(n18499), .ZN(n18618) );
  OAI22_X1 U21724 ( .A1(n9748), .A2(n18500), .B1(n18586), .B2(n18618), .ZN(
        P3_U2677) );
  INV_X1 U21725 ( .A(n18501), .ZN(n18510) );
  AOI21_X1 U21726 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18586), .A(n18510), .ZN(
        n18504) );
  OAI21_X1 U21727 ( .B1(n18506), .B2(n18503), .A(n18502), .ZN(n18623) );
  OAI22_X1 U21728 ( .A1(n18505), .A2(n18504), .B1(n18586), .B2(n18623), .ZN(
        P3_U2678) );
  AOI22_X1 U21729 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n18586), .B1(
        P3_EBX_REG_23__SCAN_IN), .B2(n18511), .ZN(n18509) );
  AOI21_X1 U21730 ( .B1(n18507), .B2(n18512), .A(n18506), .ZN(n18508) );
  INV_X1 U21731 ( .A(n18508), .ZN(n18628) );
  OAI22_X1 U21732 ( .A1(n18510), .A2(n18509), .B1(n18586), .B2(n18628), .ZN(
        P3_U2679) );
  INV_X1 U21733 ( .A(n18511), .ZN(n18516) );
  OAI21_X1 U21734 ( .B1(n18514), .B2(n18513), .A(n18512), .ZN(n18633) );
  NAND3_X1 U21735 ( .A1(n18516), .A2(P3_EBX_REG_23__SCAN_IN), .A3(n18586), 
        .ZN(n18515) );
  OAI221_X1 U21736 ( .B1(n18516), .B2(P3_EBX_REG_23__SCAN_IN), .C1(n18586), 
        .C2(n18633), .A(n18515), .ZN(P3_U2680) );
  NAND2_X1 U21737 ( .A1(n18576), .A2(n18537), .ZN(n18532) );
  AOI22_X1 U21738 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n18522) );
  AOI22_X1 U21739 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18521) );
  AOI22_X1 U21740 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18520) );
  OR2_X1 U21741 ( .A1(n18545), .A2(n18518), .ZN(n18519) );
  AND4_X1 U21742 ( .A1(n18522), .A2(n18521), .A3(n18520), .A4(n18519), .ZN(
        n18531) );
  AOI22_X1 U21743 ( .A1(n18524), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18523), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18530) );
  AOI22_X1 U21744 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18528) );
  AOI22_X1 U21745 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18527) );
  AOI22_X1 U21746 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18526) );
  NAND2_X1 U21747 ( .A1(n17762), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n18525) );
  AND4_X1 U21748 ( .A1(n18528), .A2(n18527), .A3(n18526), .A4(n18525), .ZN(
        n18529) );
  AND3_X1 U21749 ( .A1(n18531), .A2(n18530), .A3(n18529), .ZN(n18645) );
  OAI22_X1 U21750 ( .A1(n18533), .A2(n18532), .B1(n18645), .B2(n18586), .ZN(
        n18534) );
  INV_X1 U21751 ( .A(n18534), .ZN(n18535) );
  OAI21_X1 U21752 ( .B1(n18537), .B2(n18536), .A(n18535), .ZN(P3_U2682) );
  NAND2_X1 U21753 ( .A1(n9824), .A2(n18576), .ZN(n18562) );
  INV_X1 U21754 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18538) );
  OAI22_X1 U21755 ( .A1(n18541), .A2(n18540), .B1(n18539), .B2(n18538), .ZN(
        n18559) );
  AOI22_X1 U21756 ( .A1(n17774), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n18542), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18549) );
  AOI22_X1 U21757 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9690), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18548) );
  AOI22_X1 U21758 ( .A1(n17705), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18543), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18547) );
  INV_X1 U21759 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18544) );
  OR2_X1 U21760 ( .A1(n18545), .A2(n18544), .ZN(n18546) );
  NAND4_X1 U21761 ( .A1(n18549), .A2(n18548), .A3(n18547), .A4(n18546), .ZN(
        n18558) );
  AOI22_X1 U21762 ( .A1(n17782), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17700), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18556) );
  AOI22_X1 U21763 ( .A1(n18550), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13472), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18555) );
  AOI22_X1 U21764 ( .A1(n18552), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18551), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18554) );
  NAND2_X1 U21765 ( .A1(n11944), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n18553) );
  NAND4_X1 U21766 ( .A1(n18556), .A2(n18555), .A3(n18554), .A4(n18553), .ZN(
        n18557) );
  OR3_X1 U21767 ( .A1(n18559), .A2(n18558), .A3(n18557), .ZN(n18652) );
  OAI21_X1 U21768 ( .B1(n9824), .B2(n10253), .A(n18586), .ZN(n18560) );
  OAI21_X1 U21769 ( .B1(n18586), .B2(n18652), .A(n18560), .ZN(n18561) );
  OAI21_X1 U21770 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n18562), .A(n18561), .ZN(
        P3_U2685) );
  NOR2_X1 U21771 ( .A1(n18563), .A2(n19448), .ZN(n18567) );
  AOI22_X1 U21772 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n18565), .B1(n18567), .B2(
        n18564), .ZN(n18566) );
  OAI21_X1 U21773 ( .B1(n19453), .B2(n18586), .A(n18566), .ZN(P3_U2696) );
  NOR3_X1 U21774 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18590), .A3(n18569), .ZN(
        n18568) );
  AOI211_X1 U21775 ( .C1(n18590), .C2(n13816), .A(n18568), .B(n18567), .ZN(
        P3_U2697) );
  INV_X1 U21776 ( .A(n18573), .ZN(n18571) );
  NOR2_X1 U21777 ( .A1(n18590), .A2(n18569), .ZN(n18570) );
  OAI21_X1 U21778 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n18571), .A(n18570), .ZN(
        n18572) );
  OAI21_X1 U21779 ( .B1(n18586), .B2(n13699), .A(n18572), .ZN(P3_U2698) );
  OAI21_X1 U21780 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18574), .A(n18573), .ZN(
        n18575) );
  AOI22_X1 U21781 ( .A1(n18590), .A2(n13594), .B1(n18575), .B2(n18586), .ZN(
        P3_U2699) );
  NAND2_X1 U21782 ( .A1(n18587), .A2(n18576), .ZN(n18592) );
  NOR3_X1 U21783 ( .A1(n9877), .A2(n18581), .A3(n18592), .ZN(n18584) );
  NOR2_X1 U21784 ( .A1(n18590), .A2(n18577), .ZN(n18579) );
  OAI22_X1 U21785 ( .A1(n18584), .A2(n18579), .B1(n18578), .B2(n18592), .ZN(
        n18580) );
  OAI21_X1 U21786 ( .B1(n18586), .B2(n19434), .A(n18580), .ZN(P3_U2700) );
  INV_X1 U21787 ( .A(n18581), .ZN(n18582) );
  OR2_X1 U21788 ( .A1(n19448), .A2(n18582), .ZN(n18583) );
  AOI21_X1 U21789 ( .B1(n18587), .B2(n18583), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n18585) );
  AOI211_X1 U21790 ( .C1(n18590), .C2(n19429), .A(n18585), .B(n18584), .ZN(
        P3_U2701) );
  OAI222_X1 U21791 ( .A1(n18592), .A2(n18588), .B1(n9878), .B2(n18587), .C1(
        n19423), .C2(n18586), .ZN(P3_U2702) );
  AOI22_X1 U21792 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18590), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n18589), .ZN(n18591) );
  OAI21_X1 U21793 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n18592), .A(n18591), .ZN(
        P3_U2703) );
  INV_X1 U21794 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18686) );
  INV_X1 U21795 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n18690) );
  INV_X1 U21796 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18697) );
  INV_X1 U21797 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18699) );
  NOR2_X1 U21798 ( .A1(n18699), .A2(n18701), .ZN(n18593) );
  NAND4_X1 U21799 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .A4(n18593), .ZN(n18634) );
  NOR2_X1 U21800 ( .A1(n18629), .A2(n19448), .ZN(n18625) );
  NAND2_X1 U21801 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18625), .ZN(n18624) );
  NAND2_X1 U21802 ( .A1(n18598), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n18597) );
  OAI22_X1 U21803 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n18636), .B1(n18677), 
        .B2(n18598), .ZN(n18595) );
  AOI22_X1 U21804 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18653), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n18595), .ZN(n18596) );
  OAI21_X1 U21805 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n18597), .A(n18596), .ZN(
        P3_U2704) );
  AOI22_X1 U21806 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18648), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n18653), .ZN(n18600) );
  OAI211_X1 U21807 ( .C1(n18598), .C2(P3_EAX_REG_30__SCAN_IN), .A(n18662), .B(
        n18597), .ZN(n18599) );
  OAI211_X1 U21808 ( .C1(n18601), .C2(n18638), .A(n18600), .B(n18599), .ZN(
        P3_U2705) );
  AOI22_X1 U21809 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18648), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18653), .ZN(n18604) );
  OAI211_X1 U21810 ( .C1(n9753), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18662), .B(
        n18602), .ZN(n18603) );
  OAI211_X1 U21811 ( .C1(n18638), .C2(n18605), .A(n18604), .B(n18603), .ZN(
        P3_U2706) );
  AOI22_X1 U21812 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18648), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n18653), .ZN(n18608) );
  AOI211_X1 U21813 ( .C1(n18686), .C2(n18610), .A(n9753), .B(n18677), .ZN(
        n18606) );
  INV_X1 U21814 ( .A(n18606), .ZN(n18607) );
  OAI211_X1 U21815 ( .C1(n18638), .C2(n18609), .A(n18608), .B(n18607), .ZN(
        P3_U2707) );
  AOI22_X1 U21816 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18648), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18653), .ZN(n18612) );
  OAI211_X1 U21817 ( .C1(n18614), .C2(P3_EAX_REG_27__SCAN_IN), .A(n18662), .B(
        n18610), .ZN(n18611) );
  OAI211_X1 U21818 ( .C1(n18638), .C2(n18613), .A(n18612), .B(n18611), .ZN(
        P3_U2708) );
  AOI22_X1 U21819 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18648), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18653), .ZN(n18617) );
  AOI211_X1 U21820 ( .C1(n18690), .C2(n18619), .A(n18614), .B(n18677), .ZN(
        n18615) );
  INV_X1 U21821 ( .A(n18615), .ZN(n18616) );
  OAI211_X1 U21822 ( .C1(n18638), .C2(n18618), .A(n18617), .B(n18616), .ZN(
        P3_U2709) );
  AOI22_X1 U21823 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18648), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18653), .ZN(n18622) );
  OAI211_X1 U21824 ( .C1(n18620), .C2(P3_EAX_REG_25__SCAN_IN), .A(n18662), .B(
        n18619), .ZN(n18621) );
  OAI211_X1 U21825 ( .C1(n18638), .C2(n18623), .A(n18622), .B(n18621), .ZN(
        P3_U2710) );
  AOI22_X1 U21826 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18648), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18653), .ZN(n18627) );
  OAI211_X1 U21827 ( .C1(n18625), .C2(P3_EAX_REG_24__SCAN_IN), .A(n18662), .B(
        n18624), .ZN(n18626) );
  OAI211_X1 U21828 ( .C1(n18638), .C2(n18628), .A(n18627), .B(n18626), .ZN(
        P3_U2711) );
  AOI22_X1 U21829 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18648), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18653), .ZN(n18632) );
  OAI211_X1 U21830 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n18630), .A(n18662), .B(
        n18629), .ZN(n18631) );
  OAI211_X1 U21831 ( .C1(n18638), .C2(n18633), .A(n18632), .B(n18631), .ZN(
        P3_U2712) );
  NOR2_X1 U21832 ( .A1(n18635), .A2(n18634), .ZN(n18643) );
  OR2_X1 U21833 ( .A1(n18677), .A2(n18647), .ZN(n18651) );
  OAI21_X1 U21834 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18636), .A(n18651), .ZN(
        n18642) );
  INV_X1 U21835 ( .A(n18637), .ZN(n18639) );
  OAI22_X1 U21836 ( .A1(n18640), .A2(n16827), .B1(n18639), .B2(n18638), .ZN(
        n18641) );
  AOI221_X1 U21837 ( .B1(n18643), .B2(n18697), .C1(n18642), .C2(
        P3_EAX_REG_22__SCAN_IN), .A(n18641), .ZN(n18644) );
  OAI21_X1 U21838 ( .B1(n13243), .B2(n18658), .A(n18644), .ZN(P3_U2713) );
  INV_X1 U21839 ( .A(n18645), .ZN(n18646) );
  AOI22_X1 U21840 ( .A1(n18653), .A2(BUF2_REG_21__SCAN_IN), .B1(n18673), .B2(
        n18646), .ZN(n18650) );
  AOI22_X1 U21841 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18648), .B1(n18647), .B2(
        n18699), .ZN(n18649) );
  OAI211_X1 U21842 ( .C1(n18699), .C2(n18651), .A(n18650), .B(n18649), .ZN(
        P3_U2714) );
  AOI22_X1 U21843 ( .A1(n18653), .A2(BUF2_REG_18__SCAN_IN), .B1(n18673), .B2(
        n18652), .ZN(n18657) );
  OAI211_X1 U21844 ( .C1(n18655), .C2(P3_EAX_REG_18__SCAN_IN), .A(n18662), .B(
        n18654), .ZN(n18656) );
  OAI211_X1 U21845 ( .C1(n18658), .C2(n19424), .A(n18657), .B(n18656), .ZN(
        P3_U2717) );
  NAND2_X1 U21846 ( .A1(n18660), .A2(n18659), .ZN(n18666) );
  NAND2_X1 U21847 ( .A1(n18662), .A2(n18661), .ZN(n18669) );
  INV_X1 U21848 ( .A(n18663), .ZN(n18664) );
  AOI22_X1 U21849 ( .A1(n18674), .A2(BUF2_REG_15__SCAN_IN), .B1(n18673), .B2(
        n18664), .ZN(n18665) );
  OAI221_X1 U21850 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n18666), .C1(n18794), 
        .C2(n18669), .A(n18665), .ZN(P3_U2720) );
  INV_X1 U21851 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n18789) );
  AOI22_X1 U21852 ( .A1(n18674), .A2(BUF2_REG_14__SCAN_IN), .B1(n18673), .B2(
        n18667), .ZN(n18668) );
  OAI221_X1 U21853 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n18670), .C1(n18789), 
        .C2(n18669), .A(n18668), .ZN(P3_U2721) );
  XNOR2_X1 U21854 ( .A(P3_EAX_REG_10__SCAN_IN), .B(n18671), .ZN(n18676) );
  AOI22_X1 U21855 ( .A1(n18674), .A2(BUF2_REG_10__SCAN_IN), .B1(n18673), .B2(
        n18672), .ZN(n18675) );
  OAI21_X1 U21856 ( .B1(n18677), .B2(n18676), .A(n18675), .ZN(P3_U2725) );
  OR2_X1 U21857 ( .A1(n18678), .A2(n18969), .ZN(n18741) );
  INV_X2 U21858 ( .A(n18741), .ZN(n20041) );
  NOR2_X1 U21859 ( .A1(n18733), .A2(n18680), .ZN(P3_U2736) );
  INV_X1 U21860 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18764) );
  AND2_X1 U21861 ( .A1(n18738), .A2(n18681), .ZN(n18703) );
  AOI22_X1 U21862 ( .A1(n20041), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18682) );
  OAI21_X1 U21863 ( .B1(n18764), .B2(n18708), .A(n18682), .ZN(P3_U2737) );
  INV_X1 U21864 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18684) );
  INV_X2 U21865 ( .A(n18733), .ZN(n18737) );
  AOI22_X1 U21866 ( .A1(n20041), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18683) );
  OAI21_X1 U21867 ( .B1(n18684), .B2(n18708), .A(n18683), .ZN(P3_U2738) );
  AOI22_X1 U21868 ( .A1(n20041), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18685) );
  OAI21_X1 U21869 ( .B1(n18686), .B2(n18708), .A(n18685), .ZN(P3_U2739) );
  INV_X1 U21870 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18688) );
  AOI22_X1 U21871 ( .A1(n20041), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18687) );
  OAI21_X1 U21872 ( .B1(n18688), .B2(n18708), .A(n18687), .ZN(P3_U2740) );
  AOI22_X1 U21873 ( .A1(n20041), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18689) );
  OAI21_X1 U21874 ( .B1(n18690), .B2(n18708), .A(n18689), .ZN(P3_U2741) );
  INV_X1 U21875 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n18692) );
  AOI22_X1 U21876 ( .A1(n20041), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18691) );
  OAI21_X1 U21877 ( .B1(n18692), .B2(n18708), .A(n18691), .ZN(P3_U2742) );
  INV_X1 U21878 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n18757) );
  AOI22_X1 U21879 ( .A1(n20041), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18693) );
  OAI21_X1 U21880 ( .B1(n18757), .B2(n18708), .A(n18693), .ZN(P3_U2743) );
  AOI22_X1 U21881 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n18703), .B1(n20041), 
        .B2(P3_UWORD_REG_7__SCAN_IN), .ZN(n18694) );
  OAI21_X1 U21882 ( .B1(n18695), .B2(n18733), .A(n18694), .ZN(P3_U2744) );
  AOI22_X1 U21883 ( .A1(n20041), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18696) );
  OAI21_X1 U21884 ( .B1(n18697), .B2(n18708), .A(n18696), .ZN(P3_U2745) );
  AOI22_X1 U21885 ( .A1(n20041), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18698) );
  OAI21_X1 U21886 ( .B1(n18699), .B2(n18708), .A(n18698), .ZN(P3_U2746) );
  AOI22_X1 U21887 ( .A1(n20041), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18700) );
  OAI21_X1 U21888 ( .B1(n18701), .B2(n18708), .A(n18700), .ZN(P3_U2747) );
  AOI222_X1 U21889 ( .A1(n18737), .A2(P3_DATAO_REG_19__SCAN_IN), .B1(n18703), 
        .B2(P3_EAX_REG_19__SCAN_IN), .C1(n20041), .C2(P3_UWORD_REG_3__SCAN_IN), 
        .ZN(n18702) );
  INV_X1 U21890 ( .A(n18702), .ZN(P3_U2748) );
  AOI22_X1 U21891 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18703), .B1(n20041), 
        .B2(P3_UWORD_REG_2__SCAN_IN), .ZN(n18704) );
  OAI21_X1 U21892 ( .B1(n18705), .B2(n18733), .A(n18704), .ZN(P3_U2749) );
  AOI22_X1 U21893 ( .A1(n20041), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18706) );
  OAI21_X1 U21894 ( .B1(n18749), .B2(n18708), .A(n18706), .ZN(P3_U2750) );
  INV_X1 U21895 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18747) );
  AOI22_X1 U21896 ( .A1(n20041), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18707) );
  OAI21_X1 U21897 ( .B1(n18747), .B2(n18708), .A(n18707), .ZN(P3_U2751) );
  AOI22_X1 U21898 ( .A1(n20041), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18709) );
  OAI21_X1 U21899 ( .B1(n18794), .B2(n18736), .A(n18709), .ZN(P3_U2752) );
  AOI22_X1 U21900 ( .A1(n20041), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18710) );
  OAI21_X1 U21901 ( .B1(n18789), .B2(n18736), .A(n18710), .ZN(P3_U2753) );
  INV_X1 U21902 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18712) );
  AOI22_X1 U21903 ( .A1(n20041), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18711) );
  OAI21_X1 U21904 ( .B1(n18712), .B2(n18736), .A(n18711), .ZN(P3_U2754) );
  INV_X1 U21905 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18714) );
  AOI22_X1 U21906 ( .A1(n20041), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18713) );
  OAI21_X1 U21907 ( .B1(n18714), .B2(n18736), .A(n18713), .ZN(P3_U2755) );
  INV_X1 U21908 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18716) );
  AOI22_X1 U21909 ( .A1(n20041), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18715) );
  OAI21_X1 U21910 ( .B1(n18716), .B2(n18736), .A(n18715), .ZN(P3_U2756) );
  INV_X1 U21911 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18718) );
  AOI22_X1 U21912 ( .A1(n20041), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18717) );
  OAI21_X1 U21913 ( .B1(n18718), .B2(n18736), .A(n18717), .ZN(P3_U2757) );
  AOI22_X1 U21914 ( .A1(n20041), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18719) );
  OAI21_X1 U21915 ( .B1(n18720), .B2(n18736), .A(n18719), .ZN(P3_U2758) );
  AOI22_X1 U21916 ( .A1(n20041), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18721) );
  OAI21_X1 U21917 ( .B1(n18776), .B2(n18736), .A(n18721), .ZN(P3_U2759) );
  INV_X1 U21918 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18723) );
  AOI22_X1 U21919 ( .A1(n20041), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18722) );
  OAI21_X1 U21920 ( .B1(n18723), .B2(n18736), .A(n18722), .ZN(P3_U2760) );
  INV_X1 U21921 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18725) );
  AOI22_X1 U21922 ( .A1(n20041), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18724) );
  OAI21_X1 U21923 ( .B1(n18725), .B2(n18736), .A(n18724), .ZN(P3_U2761) );
  AOI22_X1 U21924 ( .A1(n20041), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18726) );
  OAI21_X1 U21925 ( .B1(n18727), .B2(n18736), .A(n18726), .ZN(P3_U2762) );
  INV_X1 U21926 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18729) );
  AOI22_X1 U21927 ( .A1(n20041), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18728) );
  OAI21_X1 U21928 ( .B1(n18729), .B2(n18736), .A(n18728), .ZN(P3_U2763) );
  AOI22_X1 U21929 ( .A1(n20041), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18730) );
  OAI21_X1 U21930 ( .B1(n18731), .B2(n18736), .A(n18730), .ZN(P3_U2764) );
  AOI22_X1 U21931 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18738), .B1(n20041), .B2(
        P3_LWORD_REG_2__SCAN_IN), .ZN(n18732) );
  OAI21_X1 U21932 ( .B1(n18734), .B2(n18733), .A(n18732), .ZN(P3_U2765) );
  AOI22_X1 U21933 ( .A1(n20041), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18737), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18735) );
  OAI21_X1 U21934 ( .B1(n18768), .B2(n18736), .A(n18735), .ZN(P3_U2766) );
  AOI22_X1 U21935 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18738), .B1(n18737), .B2(
        P3_DATAO_REG_0__SCAN_IN), .ZN(n18739) );
  OAI21_X1 U21936 ( .B1(n18741), .B2(n18740), .A(n18739), .ZN(P3_U2767) );
  NOR2_X1 U21937 ( .A1(n18745), .A2(n20031), .ZN(n19905) );
  NAND2_X1 U21938 ( .A1(n18742), .A2(n19905), .ZN(n18793) );
  NAND2_X1 U21939 ( .A1(n20031), .A2(n20032), .ZN(n18743) );
  NAND2_X1 U21940 ( .A1(n18743), .A2(n18742), .ZN(n18744) );
  OR2_X2 U21941 ( .A1(n18745), .A2(n18744), .ZN(n18790) );
  AOI22_X1 U21942 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18791), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18790), .ZN(n18746) );
  OAI21_X1 U21943 ( .B1(n18747), .B2(n18793), .A(n18746), .ZN(P3_U2768) );
  AOI22_X1 U21944 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18791), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18790), .ZN(n18748) );
  OAI21_X1 U21945 ( .B1(n18749), .B2(n18793), .A(n18748), .ZN(P3_U2769) );
  AOI22_X1 U21946 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18785), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18790), .ZN(n18750) );
  OAI21_X1 U21947 ( .B1(n19424), .B2(n18787), .A(n18750), .ZN(P3_U2770) );
  AOI22_X1 U21948 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18785), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18790), .ZN(n18751) );
  OAI21_X1 U21949 ( .B1(n19430), .B2(n18787), .A(n18751), .ZN(P3_U2771) );
  AOI22_X1 U21950 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18785), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18790), .ZN(n18752) );
  OAI21_X1 U21951 ( .B1(n19435), .B2(n18787), .A(n18752), .ZN(P3_U2772) );
  AOI22_X1 U21952 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n18785), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18790), .ZN(n18753) );
  OAI21_X1 U21953 ( .B1(n19439), .B2(n18787), .A(n18753), .ZN(P3_U2773) );
  AOI22_X1 U21954 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18785), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18790), .ZN(n18754) );
  OAI21_X1 U21955 ( .B1(n13243), .B2(n18787), .A(n18754), .ZN(P3_U2774) );
  AOI22_X1 U21956 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n18785), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18790), .ZN(n18755) );
  OAI21_X1 U21957 ( .B1(n19446), .B2(n18787), .A(n18755), .ZN(P3_U2775) );
  AOI22_X1 U21958 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18791), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18790), .ZN(n18756) );
  OAI21_X1 U21959 ( .B1(n18757), .B2(n18793), .A(n18756), .ZN(P3_U2776) );
  AOI22_X1 U21960 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n18785), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18790), .ZN(n18758) );
  OAI21_X1 U21961 ( .B1(n18778), .B2(n18787), .A(n18758), .ZN(P3_U2777) );
  AOI22_X1 U21962 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n18785), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18790), .ZN(n18759) );
  OAI21_X1 U21963 ( .B1(n18780), .B2(n18787), .A(n18759), .ZN(P3_U2778) );
  AOI22_X1 U21964 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n18785), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18790), .ZN(n18760) );
  OAI21_X1 U21965 ( .B1(n18782), .B2(n18787), .A(n18760), .ZN(P3_U2779) );
  AOI22_X1 U21966 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18785), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18790), .ZN(n18761) );
  OAI21_X1 U21967 ( .B1(n18784), .B2(n18787), .A(n18761), .ZN(P3_U2780) );
  AOI22_X1 U21968 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18785), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18790), .ZN(n18762) );
  OAI21_X1 U21969 ( .B1(n12209), .B2(n18787), .A(n18762), .ZN(P3_U2781) );
  AOI22_X1 U21970 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18791), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18790), .ZN(n18763) );
  OAI21_X1 U21971 ( .B1(n18764), .B2(n18793), .A(n18763), .ZN(P3_U2782) );
  AOI22_X1 U21972 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18791), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18790), .ZN(n18765) );
  OAI21_X1 U21973 ( .B1(n18766), .B2(n18793), .A(n18765), .ZN(P3_U2783) );
  AOI22_X1 U21974 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18791), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18790), .ZN(n18767) );
  OAI21_X1 U21975 ( .B1(n18768), .B2(n18793), .A(n18767), .ZN(P3_U2784) );
  AOI22_X1 U21976 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18785), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18790), .ZN(n18769) );
  OAI21_X1 U21977 ( .B1(n19424), .B2(n18787), .A(n18769), .ZN(P3_U2785) );
  AOI22_X1 U21978 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18785), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18790), .ZN(n18770) );
  OAI21_X1 U21979 ( .B1(n19430), .B2(n18787), .A(n18770), .ZN(P3_U2786) );
  AOI22_X1 U21980 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18785), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18790), .ZN(n18771) );
  OAI21_X1 U21981 ( .B1(n19435), .B2(n18787), .A(n18771), .ZN(P3_U2787) );
  AOI22_X1 U21982 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18785), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18790), .ZN(n18772) );
  OAI21_X1 U21983 ( .B1(n19439), .B2(n18787), .A(n18772), .ZN(P3_U2788) );
  AOI22_X1 U21984 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18785), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18790), .ZN(n18773) );
  OAI21_X1 U21985 ( .B1(n13243), .B2(n18787), .A(n18773), .ZN(P3_U2789) );
  AOI22_X1 U21986 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n18785), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18790), .ZN(n18774) );
  OAI21_X1 U21987 ( .B1(n19446), .B2(n18787), .A(n18774), .ZN(P3_U2790) );
  AOI22_X1 U21988 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18791), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18790), .ZN(n18775) );
  OAI21_X1 U21989 ( .B1(n18776), .B2(n18793), .A(n18775), .ZN(P3_U2791) );
  AOI22_X1 U21990 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18785), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18790), .ZN(n18777) );
  OAI21_X1 U21991 ( .B1(n18778), .B2(n18787), .A(n18777), .ZN(P3_U2792) );
  AOI22_X1 U21992 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18785), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18790), .ZN(n18779) );
  OAI21_X1 U21993 ( .B1(n18780), .B2(n18787), .A(n18779), .ZN(P3_U2793) );
  AOI22_X1 U21994 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n18785), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18790), .ZN(n18781) );
  OAI21_X1 U21995 ( .B1(n18782), .B2(n18787), .A(n18781), .ZN(P3_U2794) );
  AOI22_X1 U21996 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18785), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18790), .ZN(n18783) );
  OAI21_X1 U21997 ( .B1(n18784), .B2(n18787), .A(n18783), .ZN(P3_U2795) );
  AOI22_X1 U21998 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18785), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18790), .ZN(n18786) );
  OAI21_X1 U21999 ( .B1(n12209), .B2(n18787), .A(n18786), .ZN(P3_U2796) );
  AOI22_X1 U22000 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18791), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18790), .ZN(n18788) );
  OAI21_X1 U22001 ( .B1(n18789), .B2(n18793), .A(n18788), .ZN(P3_U2797) );
  AOI22_X1 U22002 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18791), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18790), .ZN(n18792) );
  OAI21_X1 U22003 ( .B1(n18794), .B2(n18793), .A(n18792), .ZN(P3_U2798) );
  AOI21_X1 U22004 ( .B1(n18795), .B2(n19801), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18805) );
  AOI22_X1 U22005 ( .A1(n19302), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n18796), 
        .B2(n19122), .ZN(n18804) );
  NOR3_X1 U22006 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n19140), .A3(
        n19133), .ZN(n19127) );
  NOR2_X1 U22007 ( .A1(n18797), .A2(n18933), .ZN(n18835) );
  INV_X1 U22008 ( .A(n19129), .ZN(n18801) );
  OAI22_X1 U22009 ( .A1(n18801), .A2(n19034), .B1(n18800), .B2(n18799), .ZN(
        n18802) );
  AOI21_X1 U22010 ( .B1(n19127), .B2(n18835), .A(n18802), .ZN(n18803) );
  OAI211_X1 U22011 ( .C1(n18806), .C2(n18805), .A(n18804), .B(n18803), .ZN(
        P3_U2804) );
  NAND2_X1 U22012 ( .A1(n18807), .A2(n19141), .ZN(n18808) );
  XNOR2_X1 U22013 ( .A(n18808), .B(n19140), .ZN(n19144) );
  OAI211_X1 U22014 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n18810), .B(n18809), .ZN(n18811) );
  NAND2_X1 U22015 ( .A1(n19302), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n19146) );
  OAI211_X1 U22016 ( .C1(n18985), .C2(n18812), .A(n18811), .B(n19146), .ZN(
        n18824) );
  NAND2_X1 U22017 ( .A1(n19141), .A2(n18813), .ZN(n18814) );
  XOR2_X1 U22018 ( .A(n18814), .B(n19140), .Z(n19137) );
  INV_X1 U22019 ( .A(n19137), .ZN(n18822) );
  XNOR2_X1 U22020 ( .A(n18815), .B(n19140), .ZN(n18818) );
  NOR2_X1 U22021 ( .A1(n18816), .A2(n19140), .ZN(n18817) );
  MUX2_X1 U22022 ( .A(n18818), .B(n18817), .S(n18966), .Z(n18819) );
  INV_X1 U22023 ( .A(n18819), .ZN(n18820) );
  OAI21_X1 U22024 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18821), .A(
        n18820), .ZN(n19148) );
  OAI22_X1 U22025 ( .A1(n19004), .A2(n18822), .B1(n19034), .B2(n19148), .ZN(
        n18823) );
  AOI211_X1 U22026 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n18825), .A(
        n18824), .B(n18823), .ZN(n18826) );
  OAI21_X1 U22027 ( .B1(n19112), .B2(n19144), .A(n18826), .ZN(P3_U2805) );
  INV_X1 U22028 ( .A(n18827), .ZN(n18828) );
  AOI22_X1 U22029 ( .A1(n17599), .A2(n18829), .B1(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18828), .ZN(n18838) );
  AND2_X1 U22030 ( .A1(n18862), .A2(n18855), .ZN(n18841) );
  NAND2_X1 U22031 ( .A1(n18950), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18831) );
  OAI211_X1 U22032 ( .C1(n9813), .C2(n18841), .A(n18830), .B(n18831), .ZN(
        n18832) );
  XNOR2_X1 U22033 ( .A(n18832), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n19149) );
  AOI22_X1 U22034 ( .A1(n19015), .A2(n19149), .B1(n18833), .B2(n19122), .ZN(
        n18837) );
  OAI21_X1 U22035 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18835), .A(
        n18834), .ZN(n18836) );
  NAND2_X1 U22036 ( .A1(n19302), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n19153) );
  NAND4_X1 U22037 ( .A1(n18838), .A2(n18837), .A3(n18836), .A4(n19153), .ZN(
        P3_U2807) );
  NOR2_X1 U22038 ( .A1(n11856), .A2(n18839), .ZN(n18840) );
  OAI21_X1 U22039 ( .B1(n18841), .B2(n18840), .A(n18830), .ZN(n18842) );
  XNOR2_X1 U22040 ( .A(n18842), .B(n19164), .ZN(n19171) );
  INV_X1 U22041 ( .A(n18843), .ZN(n18874) );
  OAI21_X1 U22042 ( .B1(n18874), .B2(n19168), .A(n18932), .ZN(n18865) );
  NOR2_X1 U22043 ( .A1(n18844), .A2(n18969), .ZN(n18845) );
  AOI211_X1 U22044 ( .C1(n19404), .C2(n18848), .A(n19096), .B(n18845), .ZN(
        n18871) );
  OAI21_X1 U22045 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18868), .A(
        n18871), .ZN(n18858) );
  AOI22_X1 U22046 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18858), .B1(
        n18977), .B2(n18846), .ZN(n18852) );
  NAND2_X1 U22047 ( .A1(n19302), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n19169) );
  NAND3_X1 U22048 ( .A1(n18847), .A2(n19168), .A3(n19164), .ZN(n18851) );
  NOR2_X1 U22049 ( .A1(n18891), .A2(n18848), .ZN(n18860) );
  OAI211_X1 U22050 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n18860), .B(n18849), .ZN(n18850) );
  NAND4_X1 U22051 ( .A1(n18852), .A2(n19169), .A3(n18851), .A4(n18850), .ZN(
        n18853) );
  AOI21_X1 U22052 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18865), .A(
        n18853), .ZN(n18854) );
  OAI21_X1 U22053 ( .B1(n19034), .B2(n19171), .A(n18854), .ZN(P3_U2808) );
  NAND4_X1 U22054 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n19199), .A3(
        n19176), .A4(n18855), .ZN(n19182) );
  OAI22_X1 U22055 ( .A1(n19349), .A2(n19984), .B1(n18985), .B2(n18856), .ZN(
        n18857) );
  AOI221_X1 U22056 ( .B1(n18860), .B2(n18859), .C1(n18858), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18857), .ZN(n18867) );
  INV_X1 U22057 ( .A(n18861), .ZN(n18863) );
  NOR4_X1 U22058 ( .A1(n11856), .A2(n19203), .A3(n19157), .A4(n18950), .ZN(
        n18884) );
  AOI22_X1 U22059 ( .A1(n18863), .A2(n18862), .B1(n19176), .B2(n18884), .ZN(
        n18864) );
  XNOR2_X1 U22060 ( .A(n18864), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n19172) );
  AOI22_X1 U22061 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18865), .B1(
        n19015), .B2(n19172), .ZN(n18866) );
  OAI211_X1 U22062 ( .C1(n18933), .C2(n19182), .A(n18867), .B(n18866), .ZN(
        P3_U2809) );
  NOR2_X1 U22063 ( .A1(n19157), .A2(n19203), .ZN(n19173) );
  NAND2_X1 U22064 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19173), .ZN(
        n19159) );
  NOR2_X1 U22065 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n19159), .ZN(
        n19183) );
  INV_X1 U22066 ( .A(n19183), .ZN(n18880) );
  AOI21_X1 U22067 ( .B1(n18869), .B2(n19801), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18870) );
  OAI22_X1 U22068 ( .A1(n18871), .A2(n18870), .B1(n19349), .B2(n19981), .ZN(
        n18872) );
  AOI221_X1 U22069 ( .B1(n18977), .B2(n18873), .C1(n13199), .C2(n18873), .A(
        n18872), .ZN(n18879) );
  INV_X1 U22070 ( .A(n19159), .ZN(n19185) );
  OAI21_X1 U22071 ( .B1(n18874), .B2(n19185), .A(n18932), .ZN(n18889) );
  INV_X1 U22072 ( .A(n18901), .ZN(n18883) );
  NAND2_X1 U22073 ( .A1(n18883), .A2(n18885), .ZN(n18875) );
  OAI211_X1 U22074 ( .C1(n18884), .C2(n18885), .A(n18830), .B(n18875), .ZN(
        n18877) );
  XNOR2_X1 U22075 ( .A(n18877), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n19184) );
  AOI22_X1 U22076 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18889), .B1(
        n19015), .B2(n19184), .ZN(n18878) );
  OAI211_X1 U22077 ( .C1(n18933), .C2(n18880), .A(n18879), .B(n18878), .ZN(
        P3_U2810) );
  AOI21_X1 U22078 ( .B1(n19404), .B2(n18890), .A(n19096), .ZN(n18910) );
  OAI21_X1 U22079 ( .B1(n18881), .B2(n18969), .A(n18910), .ZN(n18898) );
  AOI22_X1 U22080 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18898), .B1(
        n18977), .B2(n18882), .ZN(n18895) );
  NOR2_X1 U22081 ( .A1(n18861), .A2(n18883), .ZN(n18904) );
  NOR2_X1 U22082 ( .A1(n18904), .A2(n18884), .ZN(n18886) );
  XNOR2_X1 U22083 ( .A(n18886), .B(n18885), .ZN(n19195) );
  NOR3_X1 U22084 ( .A1(n19203), .A2(n19157), .A3(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n19191) );
  INV_X1 U22085 ( .A(n19191), .ZN(n18887) );
  OAI22_X1 U22086 ( .A1(n19195), .A2(n19034), .B1(n18933), .B2(n18887), .ZN(
        n18888) );
  AOI21_X1 U22087 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18889), .A(
        n18888), .ZN(n18894) );
  NAND2_X1 U22088 ( .A1(n19302), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n19194) );
  NOR2_X1 U22089 ( .A1(n18891), .A2(n18890), .ZN(n18900) );
  OAI211_X1 U22090 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18900), .B(n18892), .ZN(n18893) );
  NAND4_X1 U22091 ( .A1(n18895), .A2(n18894), .A3(n19194), .A4(n18893), .ZN(
        P3_U2811) );
  NAND2_X1 U22092 ( .A1(n19199), .A2(n19203), .ZN(n19209) );
  OAI22_X1 U22093 ( .A1(n19349), .A2(n19977), .B1(n18985), .B2(n18896), .ZN(
        n18897) );
  AOI221_X1 U22094 ( .B1(n18900), .B2(n18899), .C1(n18898), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n18897), .ZN(n18907) );
  OAI21_X1 U22095 ( .B1(n18933), .B2(n19199), .A(n18932), .ZN(n18916) );
  NOR2_X1 U22096 ( .A1(n18950), .A2(n19203), .ZN(n18903) );
  NOR2_X1 U22097 ( .A1(n18903), .A2(n18901), .ZN(n18902) );
  MUX2_X1 U22098 ( .A(n18903), .B(n18902), .S(n18861), .Z(n18905) );
  OR2_X1 U22099 ( .A1(n18905), .A2(n18904), .ZN(n19206) );
  AOI22_X1 U22100 ( .A1(n18916), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n19015), .B2(n19206), .ZN(n18906) );
  OAI211_X1 U22101 ( .C1(n18933), .C2(n19209), .A(n18907), .B(n18906), .ZN(
        P3_U2812) );
  NAND2_X1 U22102 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n19210), .ZN(
        n19216) );
  AOI21_X1 U22103 ( .B1(n19801), .B2(n18908), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18911) );
  OAI22_X1 U22104 ( .A1(n18911), .A2(n18910), .B1(n19084), .B2(n18909), .ZN(
        n18912) );
  AOI21_X1 U22105 ( .B1(n19302), .B2(P3_REIP_REG_17__SCAN_IN), .A(n18912), 
        .ZN(n18918) );
  NAND2_X1 U22106 ( .A1(n11856), .A2(n19199), .ZN(n18913) );
  OAI211_X1 U22107 ( .C1(n18915), .C2(n19210), .A(n18914), .B(n18913), .ZN(
        n19213) );
  AOI22_X1 U22108 ( .A1(n18916), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n19015), .B2(n19213), .ZN(n18917) );
  OAI211_X1 U22109 ( .C1(n18933), .C2(n19216), .A(n18918), .B(n18917), .ZN(
        P3_U2813) );
  INV_X1 U22110 ( .A(n11856), .ZN(n18920) );
  OAI21_X1 U22111 ( .B1(n18920), .B2(n18950), .A(n18919), .ZN(n18921) );
  XNOR2_X1 U22112 ( .A(n18921), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n19225) );
  AOI21_X1 U22113 ( .B1(n19404), .B2(n18922), .A(n19096), .ZN(n18956) );
  OAI21_X1 U22114 ( .B1(n18923), .B2(n18969), .A(n18956), .ZN(n18936) );
  AOI22_X1 U22115 ( .A1(n19302), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18936), .ZN(n18928) );
  NAND2_X1 U22116 ( .A1(n18968), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18925) );
  NAND2_X1 U22117 ( .A1(n18971), .A2(n18924), .ZN(n18988) );
  NOR2_X1 U22118 ( .A1(n18925), .A2(n18988), .ZN(n18947) );
  OAI211_X1 U22119 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18947), .B(n18926), .ZN(n18927) );
  OAI211_X1 U22120 ( .C1(n18985), .C2(n18929), .A(n18928), .B(n18927), .ZN(
        n18930) );
  AOI21_X1 U22121 ( .B1(n19015), .B2(n19225), .A(n18930), .ZN(n18931) );
  OAI221_X1 U22122 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18933), 
        .C1(n19228), .C2(n18932), .A(n18931), .ZN(P3_U2814) );
  INV_X1 U22123 ( .A(n19281), .ZN(n18934) );
  NOR2_X1 U22124 ( .A1(n18934), .A2(n19222), .ZN(n18959) );
  NOR2_X1 U22125 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18959), .ZN(
        n19238) );
  NAND2_X1 U22126 ( .A1(n18978), .A2(n19236), .ZN(n18949) );
  AOI22_X1 U22127 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18936), .B1(
        n18977), .B2(n18935), .ZN(n18937) );
  NAND2_X1 U22128 ( .A1(n19302), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n19243) );
  NAND2_X1 U22129 ( .A1(n18937), .A2(n19243), .ZN(n18945) );
  NAND2_X1 U22130 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18939) );
  NAND2_X1 U22131 ( .A1(n19247), .A2(n19280), .ZN(n19259) );
  NOR2_X1 U22132 ( .A1(n18939), .A2(n19259), .ZN(n18960) );
  NOR2_X1 U22133 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18960), .ZN(
        n19233) );
  NAND2_X1 U22134 ( .A1(n19121), .A2(n19230), .ZN(n18943) );
  NOR2_X1 U22135 ( .A1(n18938), .A2(n18966), .ZN(n18982) );
  NOR3_X1 U22136 ( .A1(n18963), .A2(n18939), .A3(n19272), .ZN(n18940) );
  AOI21_X1 U22137 ( .B1(n11852), .B2(n18982), .A(n18940), .ZN(n18941) );
  AOI221_X1 U22138 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n11850), 
        .C1(n18950), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n18941), .ZN(
        n18942) );
  XNOR2_X1 U22139 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18942), .ZN(
        n19231) );
  OAI22_X1 U22140 ( .A1(n19233), .A2(n18943), .B1(n19034), .B2(n19231), .ZN(
        n18944) );
  AOI211_X1 U22141 ( .C1(n18947), .C2(n18946), .A(n18945), .B(n18944), .ZN(
        n18948) );
  OAI21_X1 U22142 ( .B1(n19238), .B2(n18949), .A(n18948), .ZN(P3_U2815) );
  NOR2_X1 U22143 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18952) );
  NOR2_X1 U22144 ( .A1(n18951), .A2(n18950), .ZN(n19020) );
  INV_X1 U22145 ( .A(n19247), .ZN(n19269) );
  NOR2_X1 U22146 ( .A1(n19269), .A2(n11852), .ZN(n19246) );
  AOI22_X1 U22147 ( .A1(n18982), .A2(n18952), .B1(n19020), .B2(n19246), .ZN(
        n18953) );
  XOR2_X1 U22148 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18953), .Z(
        n19257) );
  NAND3_X1 U22149 ( .A1(n19801), .A2(n19054), .A3(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19023) );
  NOR2_X1 U22150 ( .A1(n18954), .A2(n19023), .ZN(n19000) );
  AOI21_X1 U22151 ( .B1(n18968), .B2(n19000), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18955) );
  NAND2_X1 U22152 ( .A1(n19302), .A2(P3_REIP_REG_14__SCAN_IN), .ZN(n19255) );
  OAI21_X1 U22153 ( .B1(n18956), .B2(n18955), .A(n19255), .ZN(n18957) );
  AOI21_X1 U22154 ( .B1(n18958), .B2(n19122), .A(n18957), .ZN(n18962) );
  NAND2_X1 U22155 ( .A1(n19281), .A2(n19247), .ZN(n19262) );
  AOI221_X1 U22156 ( .B1(n11852), .B2(n11851), .C1(n19262), .C2(n11851), .A(
        n18959), .ZN(n19249) );
  AOI221_X1 U22157 ( .B1(n11852), .B2(n11851), .C1(n19259), .C2(n11851), .A(
        n18960), .ZN(n19250) );
  AOI22_X1 U22158 ( .A1(n18978), .A2(n19249), .B1(n19121), .B2(n19250), .ZN(
        n18961) );
  OAI211_X1 U22159 ( .C1(n19257), .C2(n19034), .A(n18962), .B(n18961), .ZN(
        P3_U2816) );
  OAI22_X1 U22160 ( .A1(n18963), .A2(n19269), .B1(n18966), .B2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18964) );
  OAI21_X1 U22161 ( .B1(n18966), .B2(n18965), .A(n18964), .ZN(n18967) );
  XNOR2_X1 U22162 ( .A(n18967), .B(n11852), .ZN(n19268) );
  AOI211_X1 U22163 ( .C1(n18987), .C2(n18973), .A(n18968), .B(n18988), .ZN(
        n18975) );
  OAI22_X1 U22164 ( .A1(n18971), .A2(n19079), .B1(n18970), .B2(n18969), .ZN(
        n18972) );
  NOR2_X1 U22165 ( .A1(n19096), .A2(n18972), .ZN(n18986) );
  OAI22_X1 U22166 ( .A1(n18986), .A2(n18973), .B1(n19349), .B2(n19967), .ZN(
        n18974) );
  AOI211_X1 U22167 ( .C1(n18977), .C2(n18976), .A(n18975), .B(n18974), .ZN(
        n18981) );
  AOI22_X1 U22168 ( .A1(n19259), .A2(n19121), .B1(n19262), .B2(n18978), .ZN(
        n18979) );
  INV_X1 U22169 ( .A(n18979), .ZN(n18991) );
  NOR2_X1 U22170 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n19269), .ZN(
        n19258) );
  AOI22_X1 U22171 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18991), .B1(
        n19258), .B2(n19031), .ZN(n18980) );
  OAI211_X1 U22172 ( .C1(n19034), .C2(n19268), .A(n18981), .B(n18980), .ZN(
        P3_U2817) );
  INV_X1 U22173 ( .A(n19272), .ZN(n19288) );
  AOI21_X1 U22174 ( .B1(n19020), .B2(n19288), .A(n18982), .ZN(n18983) );
  XNOR2_X1 U22175 ( .A(n18983), .B(n11850), .ZN(n19278) );
  NOR2_X1 U22176 ( .A1(n18985), .A2(n18984), .ZN(n18990) );
  NAND2_X1 U22177 ( .A1(n19302), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n19276) );
  OAI221_X1 U22178 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18988), .C1(
        n18987), .C2(n18986), .A(n19276), .ZN(n18989) );
  AOI211_X1 U22179 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18991), .A(
        n18990), .B(n18989), .ZN(n18993) );
  NAND3_X1 U22180 ( .A1(n19288), .A2(n11850), .A3(n19031), .ZN(n18992) );
  OAI211_X1 U22181 ( .C1(n19278), .C2(n19034), .A(n18993), .B(n18992), .ZN(
        P3_U2818) );
  NOR2_X1 U22182 ( .A1(n18994), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n19021) );
  NOR2_X1 U22183 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19019) );
  AOI22_X1 U22184 ( .A1(n19021), .A2(n19019), .B1(n19020), .B2(n19287), .ZN(
        n18995) );
  XOR2_X1 U22185 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18995), .Z(
        n19293) );
  INV_X1 U22186 ( .A(n19287), .ZN(n18996) );
  NOR2_X1 U22187 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18996), .ZN(
        n19279) );
  NOR2_X1 U22188 ( .A1(n19110), .A2(n19963), .ZN(n19002) );
  INV_X1 U22189 ( .A(n19023), .ZN(n19037) );
  NAND2_X1 U22190 ( .A1(n18997), .A2(n19037), .ZN(n19027) );
  NOR2_X1 U22191 ( .A1(n19010), .A2(n19027), .ZN(n19009) );
  AOI21_X1 U22192 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19008), .A(
        n19009), .ZN(n18999) );
  OAI22_X1 U22193 ( .A1(n19000), .A2(n18999), .B1(n19084), .B2(n18998), .ZN(
        n19001) );
  AOI211_X1 U22194 ( .C1(n19279), .C2(n19031), .A(n19002), .B(n19001), .ZN(
        n19006) );
  INV_X1 U22195 ( .A(n19031), .ZN(n19003) );
  NOR2_X1 U22196 ( .A1(n19287), .A2(n19003), .ZN(n19007) );
  OAI22_X1 U22197 ( .A1(n19281), .A2(n19004), .B1(n19112), .B2(n19280), .ZN(
        n19032) );
  OAI21_X1 U22198 ( .B1(n19007), .B2(n19032), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n19005) );
  OAI211_X1 U22199 ( .C1(n19293), .C2(n19034), .A(n19006), .B(n19005), .ZN(
        P3_U2819) );
  INV_X1 U22200 ( .A(n19007), .ZN(n19018) );
  INV_X1 U22201 ( .A(n19008), .ZN(n19126) );
  AOI211_X1 U22202 ( .C1(n19027), .C2(n19010), .A(n19126), .B(n19009), .ZN(
        n19012) );
  NOR2_X1 U22203 ( .A1(n19349), .A2(n19961), .ZN(n19011) );
  AOI211_X1 U22204 ( .C1(n19013), .C2(n19122), .A(n19012), .B(n19011), .ZN(
        n19017) );
  AOI22_X1 U22205 ( .A1(n19021), .A2(n11849), .B1(n19020), .B2(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n19014) );
  XNOR2_X1 U22206 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n19014), .ZN(
        n19296) );
  AOI22_X1 U22207 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n19032), .B1(
        n19015), .B2(n19296), .ZN(n19016) );
  OAI211_X1 U22208 ( .C1(n19019), .C2(n19018), .A(n19017), .B(n19016), .ZN(
        P3_U2820) );
  NOR2_X1 U22209 ( .A1(n19021), .A2(n19020), .ZN(n19022) );
  XNOR2_X1 U22210 ( .A(n19022), .B(n11849), .ZN(n19312) );
  OAI22_X1 U22211 ( .A1(n19126), .A2(n19025), .B1(n19024), .B2(n19023), .ZN(
        n19026) );
  AOI22_X1 U22212 ( .A1(n19302), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n19027), 
        .B2(n19026), .ZN(n19028) );
  OAI21_X1 U22213 ( .B1(n19084), .B2(n19029), .A(n19028), .ZN(n19030) );
  AOI221_X1 U22214 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19032), .C1(
        n11849), .C2(n19031), .A(n19030), .ZN(n19033) );
  OAI21_X1 U22215 ( .B1(n19312), .B2(n19034), .A(n19033), .ZN(P3_U2821) );
  INV_X1 U22216 ( .A(n19035), .ZN(n19038) );
  INV_X1 U22217 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19955) );
  NOR2_X1 U22218 ( .A1(n19349), .A2(n19955), .ZN(n19333) );
  AOI221_X1 U22219 ( .B1(n19038), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n19037), .C2(n19036), .A(n19333), .ZN(n19047) );
  AOI21_X1 U22220 ( .B1(n19041), .B2(n19040), .A(n19039), .ZN(n19042) );
  XNOR2_X1 U22221 ( .A(n19042), .B(n19317), .ZN(n19335) );
  OAI21_X1 U22222 ( .B1(n19044), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n19043), .ZN(n19045) );
  INV_X1 U22223 ( .A(n19045), .ZN(n19334) );
  AOI22_X1 U22224 ( .A1(n19335), .A2(n19121), .B1(n19119), .B2(n19334), .ZN(
        n19046) );
  OAI211_X1 U22225 ( .C1(n19084), .C2(n19048), .A(n19047), .B(n19046), .ZN(
        P3_U2823) );
  NAND2_X1 U22226 ( .A1(n19801), .A2(n19054), .ZN(n19061) );
  OR2_X1 U22227 ( .A1(n19050), .A2(n19049), .ZN(n19051) );
  NAND2_X1 U22228 ( .A1(n19052), .A2(n19051), .ZN(n19344) );
  INV_X1 U22229 ( .A(n19344), .ZN(n19053) );
  AOI22_X1 U22230 ( .A1(n19053), .A2(n19119), .B1(n19302), .B2(
        P3_REIP_REG_6__SCAN_IN), .ZN(n19060) );
  AOI21_X1 U22231 ( .B1(n19054), .B2(n19801), .A(n19126), .ZN(n19072) );
  OAI21_X1 U22232 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n19056), .A(
        n19055), .ZN(n19342) );
  OAI22_X1 U22233 ( .A1(n19084), .A2(n19057), .B1(n19112), .B2(n19342), .ZN(
        n19058) );
  AOI21_X1 U22234 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19072), .A(
        n19058), .ZN(n19059) );
  OAI211_X1 U22235 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19061), .A(
        n19060), .B(n19059), .ZN(P3_U2824) );
  OAI21_X1 U22236 ( .B1(n19064), .B2(n19063), .A(n19062), .ZN(n19350) );
  OR2_X1 U22237 ( .A1(n19065), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n19066) );
  AND2_X1 U22238 ( .A1(n19067), .A2(n19066), .ZN(n19353) );
  AOI22_X1 U22239 ( .A1(n19119), .A2(n19353), .B1(n19302), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n19074) );
  OAI21_X1 U22240 ( .B1(n19096), .B2(n19069), .A(n19068), .ZN(n19071) );
  AOI22_X1 U22241 ( .A1(n19072), .A2(n19071), .B1(n19070), .B2(n19122), .ZN(
        n19073) );
  OAI211_X1 U22242 ( .C1(n19112), .C2(n19350), .A(n19074), .B(n19073), .ZN(
        P3_U2825) );
  OAI21_X1 U22243 ( .B1(n19077), .B2(n19076), .A(n19075), .ZN(n19078) );
  INV_X1 U22244 ( .A(n19078), .ZN(n19359) );
  NOR2_X1 U22245 ( .A1(n19110), .A2(n19949), .ZN(n19358) );
  AOI21_X1 U22246 ( .B1(n19119), .B2(n19359), .A(n19358), .ZN(n19087) );
  OAI21_X1 U22247 ( .B1(n19080), .B2(n19079), .A(n19116), .ZN(n19098) );
  OAI21_X1 U22248 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19082), .A(
        n19081), .ZN(n19367) );
  OAI22_X1 U22249 ( .A1(n19084), .A2(n19083), .B1(n19112), .B2(n19367), .ZN(
        n19085) );
  AOI21_X1 U22250 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19098), .A(
        n19085), .ZN(n19086) );
  OAI211_X1 U22251 ( .C1(n19636), .C2(n19088), .A(n19087), .B(n19086), .ZN(
        P3_U2826) );
  OAI21_X1 U22252 ( .B1(n19091), .B2(n19090), .A(n19089), .ZN(n19376) );
  OAI21_X1 U22253 ( .B1(n19093), .B2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n19092), .ZN(n19094) );
  INV_X1 U22254 ( .A(n19094), .ZN(n19369) );
  AND2_X1 U22255 ( .A1(n19302), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n19368) );
  AOI21_X1 U22256 ( .B1(n19119), .B2(n19369), .A(n19368), .ZN(n19101) );
  OAI21_X1 U22257 ( .B1(n19096), .B2(n18405), .A(n19095), .ZN(n19097) );
  AOI22_X1 U22258 ( .A1(n19099), .A2(n19122), .B1(n19098), .B2(n19097), .ZN(
        n19100) );
  OAI211_X1 U22259 ( .C1(n19112), .C2(n19376), .A(n19101), .B(n19100), .ZN(
        P3_U2827) );
  OR2_X1 U22260 ( .A1(n19103), .A2(n19102), .ZN(n19104) );
  NAND2_X1 U22261 ( .A1(n19105), .A2(n19104), .ZN(n19386) );
  OR2_X1 U22262 ( .A1(n19107), .A2(n19106), .ZN(n19108) );
  AND2_X1 U22263 ( .A1(n19109), .A2(n19108), .ZN(n19390) );
  NOR2_X1 U22264 ( .A1(n19110), .A2(n19945), .ZN(n19395) );
  AOI21_X1 U22265 ( .B1(n19119), .B2(n19390), .A(n19395), .ZN(n19111) );
  OAI21_X1 U22266 ( .B1(n19112), .B2(n19386), .A(n19111), .ZN(n19113) );
  AOI21_X1 U22267 ( .B1(n19122), .B2(n19114), .A(n19113), .ZN(n19115) );
  OAI221_X1 U22268 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19636), .C1(
        n18405), .C2(n19116), .A(n19115), .ZN(P3_U2828) );
  INV_X1 U22269 ( .A(n19117), .ZN(n19118) );
  AOI22_X1 U22270 ( .A1(n19119), .A2(n19118), .B1(n19302), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n19124) );
  AOI22_X1 U22271 ( .A1(n19122), .A2(n19125), .B1(n19121), .B2(n19120), .ZN(
        n19123) );
  OAI211_X1 U22272 ( .C1(n19126), .C2(n19125), .A(n19124), .B(n19123), .ZN(
        P3_U2829) );
  AOI22_X1 U22273 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n19128), .B1(
        n19151), .B2(n19127), .ZN(n19132) );
  AOI22_X1 U22274 ( .A1(n19129), .A2(n19297), .B1(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n19396), .ZN(n19131) );
  NAND2_X1 U22275 ( .A1(n19302), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n19130) );
  OAI211_X1 U22276 ( .C1(n19399), .C2(n19132), .A(n19131), .B(n19130), .ZN(
        P3_U2836) );
  INV_X1 U22277 ( .A(n19133), .ZN(n19136) );
  OAI211_X1 U22278 ( .C1(n19136), .C2(n19382), .A(n19135), .B(n19134), .ZN(
        n19138) );
  AOI22_X1 U22279 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n19138), .B1(
        n19263), .B2(n19137), .ZN(n19143) );
  NAND3_X1 U22280 ( .A1(n19141), .A2(n19140), .A3(n19139), .ZN(n19142) );
  OAI211_X1 U22281 ( .C1(n19144), .C2(n19387), .A(n19143), .B(n19142), .ZN(
        n19145) );
  AOI22_X1 U22282 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n19396), .B1(
        n19341), .B2(n19145), .ZN(n19147) );
  OAI211_X1 U22283 ( .C1(n19148), .C2(n19311), .A(n19147), .B(n19146), .ZN(
        P3_U2837) );
  INV_X1 U22284 ( .A(n19149), .ZN(n19154) );
  OAI221_X1 U22285 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n19151), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n19360), .A(n19150), .ZN(
        n19152) );
  OAI211_X1 U22286 ( .C1(n19154), .C2(n19311), .A(n19153), .B(n19152), .ZN(
        P3_U2839) );
  OAI221_X1 U22287 ( .B1(n19306), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C1(
        n19306), .C2(n19155), .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n19163) );
  OAI21_X1 U22288 ( .B1(n19157), .B2(n19156), .A(n19876), .ZN(n19158) );
  INV_X1 U22289 ( .A(n19158), .ZN(n19201) );
  AOI221_X1 U22290 ( .B1(n19198), .B2(n19160), .C1(n19159), .C2(n19160), .A(
        n19201), .ZN(n19161) );
  OAI211_X1 U22291 ( .C1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n19382), .A(
        n19223), .B(n19161), .ZN(n19174) );
  OAI22_X1 U22292 ( .A1(n19220), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n19168), .B2(n19286), .ZN(n19178) );
  OAI22_X1 U22293 ( .A1(n19289), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n19176), .B2(n19382), .ZN(n19162) );
  NOR4_X1 U22294 ( .A1(n19163), .A2(n19174), .A3(n19178), .A4(n19162), .ZN(
        n19165) );
  OAI22_X1 U22295 ( .A1(n19399), .A2(n19165), .B1(n19164), .B2(n19360), .ZN(
        n19166) );
  OAI221_X1 U22296 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n19168), 
        .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n19167), .A(n19166), .ZN(
        n19170) );
  OAI211_X1 U22297 ( .C1(n19171), .C2(n19311), .A(n19170), .B(n19169), .ZN(
        P3_U2840) );
  AOI22_X1 U22298 ( .A1(n19302), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n19297), 
        .B2(n19172), .ZN(n19180) );
  AOI21_X1 U22299 ( .B1(n19217), .B2(n19173), .A(n19306), .ZN(n19175) );
  OAI21_X1 U22300 ( .B1(n19176), .B2(n19187), .A(n19186), .ZN(n19177) );
  OAI211_X1 U22301 ( .C1(n19178), .C2(n19177), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n19110), .ZN(n19179) );
  OAI211_X1 U22302 ( .C1(n19182), .C2(n19181), .A(n19180), .B(n19179), .ZN(
        P3_U2841) );
  AOI22_X1 U22303 ( .A1(n19297), .A2(n19184), .B1(n19192), .B2(n19183), .ZN(
        n19190) );
  NOR3_X1 U22304 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19187), .A3(
        n20047), .ZN(n19188) );
  OAI21_X1 U22305 ( .B1(n19193), .B2(n19188), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n19189) );
  OAI211_X1 U22306 ( .C1(n19981), .C2(n19349), .A(n19190), .B(n19189), .ZN(
        P3_U2842) );
  OAI22_X1 U22307 ( .A1(n19382), .A2(n19313), .B1(n19378), .B2(n19314), .ZN(
        n19319) );
  INV_X1 U22308 ( .A(n19319), .ZN(n19371) );
  NOR2_X1 U22309 ( .A1(n19371), .A2(n19196), .ZN(n19234) );
  NAND2_X1 U22310 ( .A1(n10157), .A2(n19301), .ZN(n19229) );
  NOR2_X1 U22311 ( .A1(n19306), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n19385) );
  OR3_X1 U22312 ( .A1(n19198), .A2(n19228), .A3(n19385), .ZN(n19202) );
  OAI211_X1 U22313 ( .C1(n19199), .C2(n19286), .A(n19223), .B(n19341), .ZN(
        n19200) );
  AOI211_X1 U22314 ( .C1(n19380), .C2(n19202), .A(n19201), .B(n19200), .ZN(
        n19211) );
  NAND2_X1 U22315 ( .A1(n19210), .A2(n19380), .ZN(n19204) );
  AOI211_X1 U22316 ( .C1(n19211), .C2(n19204), .A(n19302), .B(n19203), .ZN(
        n19205) );
  AOI21_X1 U22317 ( .B1(n19297), .B2(n19206), .A(n19205), .ZN(n19208) );
  NAND2_X1 U22318 ( .A1(n19302), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n19207) );
  OAI211_X1 U22319 ( .C1(n19209), .C2(n19229), .A(n19208), .B(n19207), .ZN(
        P3_U2844) );
  NOR3_X1 U22320 ( .A1(n19211), .A2(n19302), .A3(n19210), .ZN(n19212) );
  AOI21_X1 U22321 ( .B1(n19297), .B2(n19213), .A(n19212), .ZN(n19215) );
  NAND2_X1 U22322 ( .A1(n19302), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n19214) );
  OAI211_X1 U22323 ( .C1(n19216), .C2(n19229), .A(n19215), .B(n19214), .ZN(
        P3_U2845) );
  INV_X1 U22324 ( .A(n19318), .ZN(n19316) );
  INV_X1 U22325 ( .A(n19289), .ZN(n19294) );
  AOI21_X1 U22326 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n19306), .A(
        n19217), .ZN(n19221) );
  OAI22_X1 U22327 ( .A1(n19220), .A2(n19219), .B1(n19218), .B2(n19382), .ZN(
        n19303) );
  AOI211_X1 U22328 ( .C1(n19294), .C2(n19222), .A(n19221), .B(n19303), .ZN(
        n19240) );
  OAI211_X1 U22329 ( .C1(n19316), .C2(n19240), .A(n19223), .B(n19341), .ZN(
        n19224) );
  NAND2_X1 U22330 ( .A1(n19349), .A2(n19224), .ZN(n19227) );
  AOI22_X1 U22331 ( .A1(n19302), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n19297), 
        .B2(n19225), .ZN(n19226) );
  OAI221_X1 U22332 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n19229), 
        .C1(n19228), .C2(n19227), .A(n19226), .ZN(P3_U2846) );
  NAND2_X1 U22333 ( .A1(n19875), .A2(n19230), .ZN(n19232) );
  OAI22_X1 U22334 ( .A1(n19233), .A2(n19232), .B1(n19326), .B2(n19231), .ZN(
        n19242) );
  NAND3_X1 U22335 ( .A1(n19247), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n19234), .ZN(n19253) );
  INV_X1 U22336 ( .A(n19253), .ZN(n19235) );
  AOI21_X1 U22337 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n19235), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n19239) );
  NAND2_X1 U22338 ( .A1(n19263), .A2(n19236), .ZN(n19237) );
  OAI22_X1 U22339 ( .A1(n19240), .A2(n19239), .B1(n19238), .B2(n19237), .ZN(
        n19241) );
  OAI21_X1 U22340 ( .B1(n19242), .B2(n19241), .A(n19341), .ZN(n19244) );
  OAI211_X1 U22341 ( .C1(n19360), .C2(n19245), .A(n19244), .B(n19243), .ZN(
        P3_U2847) );
  INV_X1 U22342 ( .A(n19246), .ZN(n19248) );
  INV_X1 U22343 ( .A(n19282), .ZN(n19305) );
  AOI21_X1 U22344 ( .B1(n19247), .B2(n19305), .A(n19306), .ZN(n19265) );
  AOI211_X1 U22345 ( .C1(n19318), .C2(n19248), .A(n19265), .B(n19303), .ZN(
        n19252) );
  AOI22_X1 U22346 ( .A1(n19875), .A2(n19250), .B1(n19263), .B2(n19249), .ZN(
        n19251) );
  OAI221_X1 U22347 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n19253), 
        .C1(n11851), .C2(n19252), .A(n19251), .ZN(n19254) );
  AOI22_X1 U22348 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n19396), .B1(
        n19341), .B2(n19254), .ZN(n19256) );
  OAI211_X1 U22349 ( .C1(n19257), .C2(n19311), .A(n19256), .B(n19255), .ZN(
        P3_U2848) );
  AOI22_X1 U22350 ( .A1(n19302), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n19301), 
        .B2(n19258), .ZN(n19267) );
  AOI22_X1 U22351 ( .A1(n19294), .A2(n19272), .B1(n19259), .B2(n19875), .ZN(
        n19260) );
  INV_X1 U22352 ( .A(n19260), .ZN(n19261) );
  AOI211_X1 U22353 ( .C1(n19263), .C2(n19262), .A(n19303), .B(n19261), .ZN(
        n19271) );
  OAI211_X1 U22354 ( .C1(n19289), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n19271), .B(n19341), .ZN(n19264) );
  OAI211_X1 U22355 ( .C1(n19265), .C2(n19264), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n19110), .ZN(n19266) );
  OAI211_X1 U22356 ( .C1(n19268), .C2(n19311), .A(n19267), .B(n19266), .ZN(
        P3_U2849) );
  OAI22_X1 U22357 ( .A1(n19283), .A2(n11850), .B1(n19269), .B2(n19282), .ZN(
        n19270) );
  AOI21_X1 U22358 ( .B1(n19271), .B2(n19270), .A(n19399), .ZN(n19275) );
  OAI21_X1 U22359 ( .B1(n19273), .B2(n19272), .A(n11850), .ZN(n19274) );
  AOI22_X1 U22360 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n19396), .B1(
        n19275), .B2(n19274), .ZN(n19277) );
  OAI211_X1 U22361 ( .C1(n19278), .C2(n19311), .A(n19277), .B(n19276), .ZN(
        P3_U2850) );
  AOI22_X1 U22362 ( .A1(n19302), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n19301), 
        .B2(n19279), .ZN(n19292) );
  NOR2_X1 U22363 ( .A1(n19399), .A2(n19303), .ZN(n19285) );
  OAI22_X1 U22364 ( .A1(n19281), .A2(n19322), .B1(n19387), .B2(n19280), .ZN(
        n19308) );
  AOI221_X1 U22365 ( .B1(n11849), .B2(n19283), .C1(n19282), .C2(n19283), .A(
        n19308), .ZN(n19284) );
  OAI211_X1 U22366 ( .C1(n19287), .C2(n19286), .A(n19285), .B(n19284), .ZN(
        n19295) );
  OAI22_X1 U22367 ( .A1(n19289), .A2(n19288), .B1(n19306), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19290) );
  OAI211_X1 U22368 ( .C1(n19295), .C2(n19290), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n19110), .ZN(n19291) );
  OAI211_X1 U22369 ( .C1(n19293), .C2(n19311), .A(n19292), .B(n19291), .ZN(
        P3_U2851) );
  NAND2_X1 U22370 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n19301), .ZN(
        n19300) );
  OAI221_X1 U22371 ( .B1(n19295), .B2(n19294), .C1(n19295), .C2(n11849), .A(
        n19110), .ZN(n19299) );
  AOI22_X1 U22372 ( .A1(n19302), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n19297), 
        .B2(n19296), .ZN(n19298) );
  OAI221_X1 U22373 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n19300), 
        .C1(n11847), .C2(n19299), .A(n19298), .ZN(P3_U2852) );
  AOI22_X1 U22374 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n19302), .B1(n19301), 
        .B2(n11849), .ZN(n19310) );
  INV_X1 U22375 ( .A(n19303), .ZN(n19304) );
  OAI211_X1 U22376 ( .C1(n19306), .C2(n19305), .A(n19304), .B(n19341), .ZN(
        n19307) );
  OAI211_X1 U22377 ( .C1(n19308), .C2(n19307), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n19110), .ZN(n19309) );
  OAI211_X1 U22378 ( .C1(n19312), .C2(n19311), .A(n19310), .B(n19309), .ZN(
        P3_U2853) );
  INV_X1 U22379 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n19346) );
  AND2_X1 U22380 ( .A1(n19876), .A2(n19313), .ZN(n19389) );
  AOI211_X1 U22381 ( .C1(n19380), .C2(n19314), .A(n19389), .B(n19385), .ZN(
        n19372) );
  OAI21_X1 U22382 ( .B1(n19316), .B2(n19315), .A(n19372), .ZN(n19340) );
  AOI211_X1 U22383 ( .C1(n19318), .C2(n19346), .A(n19317), .B(n19340), .ZN(
        n19339) );
  OAI21_X1 U22384 ( .B1(n19339), .B2(n19361), .A(n19360), .ZN(n19329) );
  NAND3_X1 U22385 ( .A1(n19320), .A2(n10305), .A3(n19319), .ZN(n19321) );
  OAI21_X1 U22386 ( .B1(n14570), .B2(n19322), .A(n19321), .ZN(n19323) );
  AOI21_X1 U22387 ( .B1(n19324), .B2(n19875), .A(n19323), .ZN(n19325) );
  OAI21_X1 U22388 ( .B1(n19327), .B2(n19326), .A(n19325), .ZN(n19328) );
  AOI22_X1 U22389 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n19329), .B1(
        n19341), .B2(n19328), .ZN(n19330) );
  OAI21_X1 U22390 ( .B1(n19349), .B2(n19958), .A(n19330), .ZN(P3_U2854) );
  NOR2_X1 U22391 ( .A1(n19371), .A2(n19331), .ZN(n19332) );
  OAI21_X1 U22392 ( .B1(n19332), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n19341), .ZN(n19338) );
  AOI21_X1 U22393 ( .B1(n19396), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n19333), .ZN(n19337) );
  AOI22_X1 U22394 ( .A1(n19335), .A2(n19351), .B1(n19370), .B2(n19334), .ZN(
        n19336) );
  OAI211_X1 U22395 ( .C1(n19339), .C2(n19338), .A(n19337), .B(n19336), .ZN(
        P3_U2855) );
  AOI21_X1 U22396 ( .B1(n19341), .B2(n19340), .A(n19396), .ZN(n19355) );
  OAI222_X1 U22397 ( .A1(n19344), .A2(n19343), .B1(n19355), .B2(n19346), .C1(
        n19377), .C2(n19342), .ZN(n19345) );
  INV_X1 U22398 ( .A(n19345), .ZN(n19348) );
  NOR3_X1 U22399 ( .A1(n19399), .A2(n19371), .A3(n9976), .ZN(n19363) );
  NAND4_X1 U22400 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n19363), .A4(n19346), .ZN(
        n19347) );
  OAI211_X1 U22401 ( .C1(n19953), .C2(n19349), .A(n19348), .B(n19347), .ZN(
        P3_U2856) );
  NAND2_X1 U22402 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n19363), .ZN(
        n19357) );
  INV_X1 U22403 ( .A(n19350), .ZN(n19352) );
  AOI222_X1 U22404 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n19302), .B1(n19370), 
        .B2(n19353), .C1(n19352), .C2(n19351), .ZN(n19354) );
  OAI221_X1 U22405 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n19357), .C1(
        n19356), .C2(n19355), .A(n19354), .ZN(P3_U2857) );
  AOI21_X1 U22406 ( .B1(n19359), .B2(n19370), .A(n19358), .ZN(n19366) );
  OAI221_X1 U22407 ( .B1(n19361), .B2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C1(
        n19361), .C2(n19372), .A(n19360), .ZN(n19364) );
  AOI22_X1 U22408 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n19364), .B1(
        n19363), .B2(n19362), .ZN(n19365) );
  OAI211_X1 U22409 ( .C1(n19377), .C2(n19367), .A(n19366), .B(n19365), .ZN(
        P3_U2858) );
  AOI21_X1 U22410 ( .B1(n19370), .B2(n19369), .A(n19368), .ZN(n19375) );
  AOI221_X1 U22411 ( .B1(n19372), .B2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C1(
        n19371), .C2(n9976), .A(n19399), .ZN(n19373) );
  AOI21_X1 U22412 ( .B1(n19396), .B2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n19373), .ZN(n19374) );
  OAI211_X1 U22413 ( .C1(n19377), .C2(n19376), .A(n19375), .B(n19374), .ZN(
        P3_U2859) );
  OR3_X1 U22414 ( .A1(n19379), .A2(n19378), .A3(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19394) );
  INV_X1 U22415 ( .A(n19380), .ZN(n19383) );
  NAND2_X1 U22416 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19381) );
  OAI22_X1 U22417 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19383), .B1(
        n19382), .B2(n19381), .ZN(n19384) );
  OAI21_X1 U22418 ( .B1(n19385), .B2(n19384), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19393) );
  NOR2_X1 U22419 ( .A1(n19387), .A2(n19386), .ZN(n19388) );
  AOI211_X1 U22420 ( .C1(n19391), .C2(n19390), .A(n19389), .B(n19388), .ZN(
        n19392) );
  AND3_X1 U22421 ( .A1(n19394), .A2(n19393), .A3(n19392), .ZN(n19398) );
  AOI21_X1 U22422 ( .B1(n19396), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n19395), .ZN(n19397) );
  OAI21_X1 U22423 ( .B1(n19399), .B2(n19398), .A(n19397), .ZN(P3_U2860) );
  AOI21_X1 U22424 ( .B1(n19402), .B2(n19401), .A(n19400), .ZN(n19912) );
  OAI21_X1 U22425 ( .B1(n19912), .B2(n19454), .A(n19413), .ZN(n19403) );
  OAI221_X1 U22426 ( .B1(n12049), .B2(n20037), .C1(n12049), .C2(n19413), .A(
        n19403), .ZN(P3_U2863) );
  OAI21_X1 U22427 ( .B1(n19404), .B2(n20037), .A(n20016), .ZN(n19406) );
  AOI211_X1 U22428 ( .C1(n19406), .C2(n19858), .A(n19405), .B(n19454), .ZN(
        n19410) );
  OAI221_X1 U22429 ( .B1(n19408), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n19408), .C2(n19407), .A(n19413), .ZN(n19411) );
  AOI22_X1 U22430 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19410), .B1(
        n19411), .B2(n19409), .ZN(P3_U2865) );
  NOR2_X1 U22431 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19409), .ZN(
        n19588) );
  INV_X1 U22432 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19889) );
  NOR2_X1 U22433 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19889), .ZN(
        n19688) );
  NOR2_X1 U22434 ( .A1(n19588), .A2(n19688), .ZN(n19412) );
  OAI22_X1 U22435 ( .A1(n19412), .A2(n19411), .B1(n19889), .B2(n19410), .ZN(
        P3_U2866) );
  NOR2_X1 U22436 ( .A1(n19890), .A2(n19413), .ZN(P3_U2867) );
  NAND2_X1 U22437 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19860) );
  NAND2_X1 U22438 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19735) );
  NOR2_X2 U22439 ( .A1(n19860), .A2(n19735), .ZN(n19821) );
  NAND2_X1 U22440 ( .A1(n19858), .A2(n12049), .ZN(n19864) );
  NOR2_X1 U22441 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19456) );
  INV_X1 U22442 ( .A(n19456), .ZN(n19497) );
  NOR2_X1 U22443 ( .A1(n19864), .A2(n19497), .ZN(n19517) );
  NOR2_X1 U22444 ( .A1(n19821), .A2(n19505), .ZN(n19477) );
  OAI21_X1 U22445 ( .B1(n12049), .B2(n20016), .A(n19765), .ZN(n19564) );
  NOR2_X1 U22446 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n12049), .ZN(
        n19457) );
  INV_X1 U22447 ( .A(n19457), .ZN(n19637) );
  NOR2_X2 U22448 ( .A1(n19637), .A2(n19735), .ZN(n19847) );
  INV_X1 U22449 ( .A(n19735), .ZN(n19737) );
  NAND2_X1 U22450 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19737), .ZN(
        n19795) );
  NOR2_X2 U22451 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19795), .ZN(
        n19773) );
  NOR2_X1 U22452 ( .A1(n19847), .A2(n19773), .ZN(n19761) );
  OAI22_X1 U22453 ( .A1(n19477), .A2(n19564), .B1(n19761), .B2(n19636), .ZN(
        n19452) );
  NAND2_X1 U22454 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19801), .ZN(n19805) );
  INV_X1 U22455 ( .A(n19805), .ZN(n19760) );
  NOR2_X2 U22456 ( .A1(n19455), .A2(n13564), .ZN(n19796) );
  NOR2_X1 U22457 ( .A1(n19918), .A2(n19477), .ZN(n19447) );
  AOI22_X1 U22458 ( .A1(n19760), .A2(n19847), .B1(n19796), .B2(n19447), .ZN(
        n19418) );
  NOR2_X1 U22459 ( .A1(n19415), .A2(n19414), .ZN(n19449) );
  INV_X1 U22460 ( .A(n19449), .ZN(n19425) );
  NOR2_X2 U22461 ( .A1(n10081), .A2(n19425), .ZN(n19802) );
  NOR2_X1 U22462 ( .A1(n19636), .A2(n19416), .ZN(n19797) );
  AOI22_X1 U22463 ( .A1(n19802), .A2(n19505), .B1(n19797), .B2(n19773), .ZN(
        n19417) );
  OAI211_X1 U22464 ( .C1(n19419), .C2(n19452), .A(n19418), .B(n19417), .ZN(
        P3_U2868) );
  NOR2_X2 U22465 ( .A1(n19455), .A2(n13462), .ZN(n19806) );
  NAND2_X1 U22466 ( .A1(n19801), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19812) );
  INV_X1 U22467 ( .A(n19812), .ZN(n19769) );
  AOI22_X1 U22468 ( .A1(n19806), .A2(n19447), .B1(n19769), .B2(n19773), .ZN(
        n19422) );
  NAND2_X1 U22469 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19801), .ZN(n19772) );
  INV_X1 U22470 ( .A(n19772), .ZN(n19807) );
  NOR2_X2 U22471 ( .A1(n19420), .A2(n19425), .ZN(n19808) );
  AOI22_X1 U22472 ( .A1(n19807), .A2(n19847), .B1(n19808), .B2(n19505), .ZN(
        n19421) );
  OAI211_X1 U22473 ( .C1(n19423), .C2(n19452), .A(n19422), .B(n19421), .ZN(
        P3_U2869) );
  NAND2_X1 U22474 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19801), .ZN(n19778) );
  INV_X1 U22475 ( .A(n19778), .ZN(n19814) );
  NOR2_X2 U22476 ( .A1(n19455), .A2(n19424), .ZN(n19813) );
  AOI22_X1 U22477 ( .A1(n19814), .A2(n19847), .B1(n19813), .B2(n19447), .ZN(
        n19428) );
  OR2_X1 U22478 ( .A1(n19426), .A2(n19425), .ZN(n19818) );
  INV_X1 U22479 ( .A(n19818), .ZN(n19774) );
  NOR2_X2 U22480 ( .A1(n19636), .A2(n16860), .ZN(n19815) );
  AOI22_X1 U22481 ( .A1(n19774), .A2(n19505), .B1(n19815), .B2(n19773), .ZN(
        n19427) );
  OAI211_X1 U22482 ( .C1(n19429), .C2(n19452), .A(n19428), .B(n19427), .ZN(
        P3_U2870) );
  NAND2_X1 U22483 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19801), .ZN(n19826) );
  INV_X1 U22484 ( .A(n19826), .ZN(n19779) );
  NOR2_X2 U22485 ( .A1(n19455), .A2(n19430), .ZN(n19820) );
  AOI22_X1 U22486 ( .A1(n19779), .A2(n19847), .B1(n19820), .B2(n19447), .ZN(
        n19433) );
  AND2_X1 U22487 ( .A1(n19431), .A2(n19449), .ZN(n19822) );
  AND2_X1 U22488 ( .A1(n19801), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19819) );
  AOI22_X1 U22489 ( .A1(n19822), .A2(n19505), .B1(n19819), .B2(n19773), .ZN(
        n19432) );
  OAI211_X1 U22490 ( .C1(n19434), .C2(n19452), .A(n19433), .B(n19432), .ZN(
        P3_U2871) );
  AND2_X1 U22491 ( .A1(n19801), .A2(BUF2_REG_20__SCAN_IN), .ZN(n19829) );
  NOR2_X2 U22492 ( .A1(n19455), .A2(n19435), .ZN(n19827) );
  AOI22_X1 U22493 ( .A1(n19829), .A2(n19773), .B1(n19827), .B2(n19447), .ZN(
        n19438) );
  NAND2_X1 U22494 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19801), .ZN(n19723) );
  INV_X1 U22495 ( .A(n19723), .ZN(n19828) );
  AND2_X1 U22496 ( .A1(n19436), .A2(n19449), .ZN(n19720) );
  AOI22_X1 U22497 ( .A1(n19828), .A2(n19847), .B1(n19720), .B2(n19517), .ZN(
        n19437) );
  OAI211_X1 U22498 ( .C1(n13594), .C2(n19452), .A(n19438), .B(n19437), .ZN(
        P3_U2872) );
  NOR2_X2 U22499 ( .A1(n19455), .A2(n19439), .ZN(n19833) );
  AOI22_X1 U22500 ( .A1(n19835), .A2(n19773), .B1(n19833), .B2(n19447), .ZN(
        n19442) );
  NAND2_X1 U22501 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19801), .ZN(n19753) );
  INV_X1 U22502 ( .A(n19753), .ZN(n19834) );
  AND2_X1 U22503 ( .A1(n19440), .A2(n19449), .ZN(n19749) );
  AOI22_X1 U22504 ( .A1(n19834), .A2(n19847), .B1(n19749), .B2(n19517), .ZN(
        n19441) );
  OAI211_X1 U22505 ( .C1(n13699), .C2(n19452), .A(n19442), .B(n19441), .ZN(
        P3_U2873) );
  NOR2_X2 U22506 ( .A1(n19636), .A2(n16827), .ZN(n19840) );
  NOR2_X2 U22507 ( .A1(n19455), .A2(n13243), .ZN(n19839) );
  AOI22_X1 U22508 ( .A1(n19840), .A2(n19773), .B1(n19839), .B2(n19447), .ZN(
        n19445) );
  AND2_X1 U22509 ( .A1(n19449), .A2(n19443), .ZN(n19657) );
  NOR2_X2 U22510 ( .A1(n16771), .A2(n19636), .ZN(n19841) );
  AOI22_X1 U22511 ( .A1(n19657), .A2(n19505), .B1(n19841), .B2(n19847), .ZN(
        n19444) );
  OAI211_X1 U22512 ( .C1(n13816), .C2(n19452), .A(n19445), .B(n19444), .ZN(
        P3_U2874) );
  AND2_X1 U22513 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19801), .ZN(n19848) );
  NOR2_X2 U22514 ( .A1(n19446), .A2(n19455), .ZN(n19846) );
  AOI22_X1 U22515 ( .A1(n19848), .A2(n19773), .B1(n19846), .B2(n19447), .ZN(
        n19451) );
  AND2_X1 U22516 ( .A1(n19449), .A2(n19448), .ZN(n19472) );
  NOR2_X2 U22517 ( .A1(n19636), .A2(n16767), .ZN(n19850) );
  AOI22_X1 U22518 ( .A1(n19472), .A2(n19505), .B1(n19850), .B2(n19847), .ZN(
        n19450) );
  OAI211_X1 U22519 ( .C1(n19453), .C2(n19452), .A(n19451), .B(n19450), .ZN(
        P3_U2875) );
  INV_X1 U22520 ( .A(n19773), .ZN(n19794) );
  NAND2_X1 U22521 ( .A1(n19858), .A2(n19907), .ZN(n19734) );
  NOR2_X1 U22522 ( .A1(n19497), .A2(n19734), .ZN(n19473) );
  AOI22_X1 U22523 ( .A1(n19797), .A2(n19821), .B1(n19796), .B2(n19473), .ZN(
        n19459) );
  INV_X1 U22524 ( .A(n19795), .ZN(n19799) );
  NOR2_X1 U22525 ( .A1(n19455), .A2(n19454), .ZN(n19798) );
  INV_X1 U22526 ( .A(n19798), .ZN(n19634) );
  NOR2_X1 U22527 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19634), .ZN(
        n19736) );
  AOI22_X1 U22528 ( .A1(n19801), .A2(n19799), .B1(n19456), .B2(n19736), .ZN(
        n19474) );
  NAND2_X1 U22529 ( .A1(n19457), .A2(n19456), .ZN(n19535) );
  INV_X1 U22530 ( .A(n19535), .ZN(n19539) );
  AOI22_X1 U22531 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19474), .B1(
        n19539), .B2(n19802), .ZN(n19458) );
  OAI211_X1 U22532 ( .C1(n19805), .C2(n19794), .A(n19459), .B(n19458), .ZN(
        P3_U2876) );
  AOI22_X1 U22533 ( .A1(n19806), .A2(n19473), .B1(n19769), .B2(n19821), .ZN(
        n19461) );
  AOI22_X1 U22534 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19474), .B1(
        n19539), .B2(n19808), .ZN(n19460) );
  OAI211_X1 U22535 ( .C1(n19772), .C2(n19794), .A(n19461), .B(n19460), .ZN(
        P3_U2877) );
  AOI22_X1 U22536 ( .A1(n19814), .A2(n19773), .B1(n19813), .B2(n19473), .ZN(
        n19463) );
  AOI22_X1 U22537 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19474), .B1(
        n19815), .B2(n19821), .ZN(n19462) );
  OAI211_X1 U22538 ( .C1(n19535), .C2(n19818), .A(n19463), .B(n19462), .ZN(
        P3_U2878) );
  INV_X1 U22539 ( .A(n19822), .ZN(n19782) );
  AOI22_X1 U22540 ( .A1(n19779), .A2(n19773), .B1(n19820), .B2(n19473), .ZN(
        n19465) );
  AOI22_X1 U22541 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19474), .B1(
        n19819), .B2(n19821), .ZN(n19464) );
  OAI211_X1 U22542 ( .C1(n19535), .C2(n19782), .A(n19465), .B(n19464), .ZN(
        P3_U2879) );
  INV_X1 U22543 ( .A(n19720), .ZN(n19832) );
  AOI22_X1 U22544 ( .A1(n19828), .A2(n19773), .B1(n19827), .B2(n19473), .ZN(
        n19467) );
  AOI22_X1 U22545 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19474), .B1(
        n19829), .B2(n19821), .ZN(n19466) );
  OAI211_X1 U22546 ( .C1(n19535), .C2(n19832), .A(n19467), .B(n19466), .ZN(
        P3_U2880) );
  AOI22_X1 U22547 ( .A1(n19835), .A2(n19821), .B1(n19833), .B2(n19473), .ZN(
        n19469) );
  AOI22_X1 U22548 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19474), .B1(
        n19539), .B2(n19749), .ZN(n19468) );
  OAI211_X1 U22549 ( .C1(n19753), .C2(n19794), .A(n19469), .B(n19468), .ZN(
        P3_U2881) );
  AOI22_X1 U22550 ( .A1(n19839), .A2(n19473), .B1(n19841), .B2(n19773), .ZN(
        n19471) );
  AOI22_X1 U22551 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19474), .B1(
        n19840), .B2(n19821), .ZN(n19470) );
  OAI211_X1 U22552 ( .C1(n19535), .C2(n19844), .A(n19471), .B(n19470), .ZN(
        P3_U2882) );
  INV_X1 U22553 ( .A(n19472), .ZN(n19855) );
  AOI22_X1 U22554 ( .A1(n19846), .A2(n19473), .B1(n19850), .B2(n19773), .ZN(
        n19476) );
  AOI22_X1 U22555 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19474), .B1(
        n19848), .B2(n19821), .ZN(n19475) );
  OAI211_X1 U22556 ( .C1(n19535), .C2(n19855), .A(n19476), .B(n19475), .ZN(
        P3_U2883) );
  INV_X1 U22557 ( .A(n19821), .ZN(n19854) );
  NOR2_X1 U22558 ( .A1(n19858), .A2(n19497), .ZN(n19543) );
  NAND2_X1 U22559 ( .A1(n12049), .A2(n19543), .ZN(n19556) );
  NOR2_X1 U22560 ( .A1(n19539), .A2(n19560), .ZN(n19521) );
  NOR2_X1 U22561 ( .A1(n19918), .A2(n19521), .ZN(n19493) );
  AOI22_X1 U22562 ( .A1(n19797), .A2(n19505), .B1(n19796), .B2(n19493), .ZN(
        n19480) );
  OAI21_X1 U22563 ( .B1(n19477), .B2(n19762), .A(n19521), .ZN(n19478) );
  OAI211_X1 U22564 ( .C1(n19560), .C2(n20016), .A(n19765), .B(n19478), .ZN(
        n19494) );
  AOI22_X1 U22565 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19494), .B1(
        n19560), .B2(n19802), .ZN(n19479) );
  OAI211_X1 U22566 ( .C1(n19805), .C2(n19854), .A(n19480), .B(n19479), .ZN(
        P3_U2884) );
  AOI22_X1 U22567 ( .A1(n19806), .A2(n19493), .B1(n19769), .B2(n19505), .ZN(
        n19482) );
  AOI22_X1 U22568 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19494), .B1(
        n19560), .B2(n19808), .ZN(n19481) );
  OAI211_X1 U22569 ( .C1(n19772), .C2(n19854), .A(n19482), .B(n19481), .ZN(
        P3_U2885) );
  AOI22_X1 U22570 ( .A1(n19814), .A2(n19821), .B1(n19813), .B2(n19493), .ZN(
        n19484) );
  AOI22_X1 U22571 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19494), .B1(
        n19815), .B2(n19505), .ZN(n19483) );
  OAI211_X1 U22572 ( .C1(n19556), .C2(n19818), .A(n19484), .B(n19483), .ZN(
        P3_U2886) );
  AOI22_X1 U22573 ( .A1(n19779), .A2(n19821), .B1(n19820), .B2(n19493), .ZN(
        n19486) );
  AOI22_X1 U22574 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19494), .B1(
        n19819), .B2(n19517), .ZN(n19485) );
  OAI211_X1 U22575 ( .C1(n19556), .C2(n19782), .A(n19486), .B(n19485), .ZN(
        P3_U2887) );
  AOI22_X1 U22576 ( .A1(n19828), .A2(n19821), .B1(n19827), .B2(n19493), .ZN(
        n19488) );
  AOI22_X1 U22577 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19494), .B1(
        n19829), .B2(n19505), .ZN(n19487) );
  OAI211_X1 U22578 ( .C1(n19556), .C2(n19832), .A(n19488), .B(n19487), .ZN(
        P3_U2888) );
  INV_X1 U22579 ( .A(n19749), .ZN(n19838) );
  AOI22_X1 U22580 ( .A1(n19834), .A2(n19821), .B1(n19833), .B2(n19493), .ZN(
        n19490) );
  AOI22_X1 U22581 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19494), .B1(
        n19835), .B2(n19505), .ZN(n19489) );
  OAI211_X1 U22582 ( .C1(n19556), .C2(n19838), .A(n19490), .B(n19489), .ZN(
        P3_U2889) );
  AOI22_X1 U22583 ( .A1(n19840), .A2(n19505), .B1(n19839), .B2(n19493), .ZN(
        n19492) );
  AOI22_X1 U22584 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19494), .B1(
        n19841), .B2(n19821), .ZN(n19491) );
  OAI211_X1 U22585 ( .C1(n19556), .C2(n19844), .A(n19492), .B(n19491), .ZN(
        P3_U2890) );
  AOI22_X1 U22586 ( .A1(n19848), .A2(n19505), .B1(n19846), .B2(n19493), .ZN(
        n19496) );
  AOI22_X1 U22587 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19494), .B1(
        n19850), .B2(n19821), .ZN(n19495) );
  OAI211_X1 U22588 ( .C1(n19556), .C2(n19855), .A(n19496), .B(n19495), .ZN(
        P3_U2891) );
  AOI211_X1 U22589 ( .C1(n19858), .C2(n19762), .A(n19497), .B(n19634), .ZN(
        n19515) );
  AND2_X1 U22590 ( .A1(n19907), .A2(n19543), .ZN(n19516) );
  AOI22_X1 U22591 ( .A1(n19760), .A2(n19505), .B1(n19796), .B2(n19516), .ZN(
        n19499) );
  NOR2_X2 U22592 ( .A1(n19860), .A2(n19497), .ZN(n19583) );
  AOI22_X1 U22593 ( .A1(n19539), .A2(n19797), .B1(n19583), .B2(n19802), .ZN(
        n19498) );
  OAI211_X1 U22594 ( .C1(n19515), .C2(n19500), .A(n19499), .B(n19498), .ZN(
        P3_U2892) );
  AOI22_X1 U22595 ( .A1(n19539), .A2(n19769), .B1(n19806), .B2(n19516), .ZN(
        n19502) );
  AOI22_X1 U22596 ( .A1(n19583), .A2(n19808), .B1(n19807), .B2(n19517), .ZN(
        n19501) );
  OAI211_X1 U22597 ( .C1(n19515), .C2(n17698), .A(n19502), .B(n19501), .ZN(
        P3_U2893) );
  AOI22_X1 U22598 ( .A1(n19539), .A2(n19815), .B1(n19813), .B2(n19516), .ZN(
        n19504) );
  INV_X1 U22599 ( .A(n19515), .ZN(n19518) );
  AOI22_X1 U22600 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19518), .B1(
        n19814), .B2(n19517), .ZN(n19503) );
  OAI211_X1 U22601 ( .C1(n19579), .C2(n19818), .A(n19504), .B(n19503), .ZN(
        P3_U2894) );
  AOI22_X1 U22602 ( .A1(n19779), .A2(n19505), .B1(n19820), .B2(n19516), .ZN(
        n19507) );
  AOI22_X1 U22603 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19518), .B1(
        n19539), .B2(n19819), .ZN(n19506) );
  OAI211_X1 U22604 ( .C1(n19579), .C2(n19782), .A(n19507), .B(n19506), .ZN(
        P3_U2895) );
  AOI22_X1 U22605 ( .A1(n19539), .A2(n19829), .B1(n19827), .B2(n19516), .ZN(
        n19509) );
  AOI22_X1 U22606 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19518), .B1(
        n19828), .B2(n19517), .ZN(n19508) );
  OAI211_X1 U22607 ( .C1(n19579), .C2(n19832), .A(n19509), .B(n19508), .ZN(
        P3_U2896) );
  AOI22_X1 U22608 ( .A1(n19539), .A2(n19835), .B1(n19833), .B2(n19516), .ZN(
        n19511) );
  AOI22_X1 U22609 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19518), .B1(
        n19834), .B2(n19517), .ZN(n19510) );
  OAI211_X1 U22610 ( .C1(n19579), .C2(n19838), .A(n19511), .B(n19510), .ZN(
        P3_U2897) );
  AOI22_X1 U22611 ( .A1(n19539), .A2(n19840), .B1(n19839), .B2(n19516), .ZN(
        n19513) );
  AOI22_X1 U22612 ( .A1(n19583), .A2(n19657), .B1(n19841), .B2(n19517), .ZN(
        n19512) );
  OAI211_X1 U22613 ( .C1(n19515), .C2(n19514), .A(n19513), .B(n19512), .ZN(
        P3_U2898) );
  AOI22_X1 U22614 ( .A1(n19539), .A2(n19848), .B1(n19846), .B2(n19516), .ZN(
        n19520) );
  AOI22_X1 U22615 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19518), .B1(
        n19850), .B2(n19517), .ZN(n19519) );
  OAI211_X1 U22616 ( .C1(n19579), .C2(n19855), .A(n19520), .B(n19519), .ZN(
        P3_U2899) );
  INV_X1 U22617 ( .A(n19588), .ZN(n19589) );
  INV_X1 U22618 ( .A(n9683), .ZN(n19600) );
  AOI21_X1 U22619 ( .B1(n19600), .B2(n19579), .A(n19918), .ZN(n19538) );
  AOI22_X1 U22620 ( .A1(n19560), .A2(n19797), .B1(n19796), .B2(n19538), .ZN(
        n19524) );
  AOI221_X1 U22621 ( .B1(n19521), .B2(n19579), .C1(n19762), .C2(n19579), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19522) );
  OAI21_X1 U22622 ( .B1(n9683), .B2(n19522), .A(n19765), .ZN(n19540) );
  AOI22_X1 U22623 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19540), .B1(
        n9683), .B2(n19802), .ZN(n19523) );
  OAI211_X1 U22624 ( .C1(n19805), .C2(n19535), .A(n19524), .B(n19523), .ZN(
        P3_U2900) );
  AOI22_X1 U22625 ( .A1(n19560), .A2(n19769), .B1(n19538), .B2(n19806), .ZN(
        n19526) );
  AOI22_X1 U22626 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19540), .B1(
        n9683), .B2(n19808), .ZN(n19525) );
  OAI211_X1 U22627 ( .C1(n19535), .C2(n19772), .A(n19526), .B(n19525), .ZN(
        P3_U2901) );
  AOI22_X1 U22628 ( .A1(n19560), .A2(n19815), .B1(n19538), .B2(n19813), .ZN(
        n19528) );
  AOI22_X1 U22629 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19540), .B1(
        n9683), .B2(n19774), .ZN(n19527) );
  OAI211_X1 U22630 ( .C1(n19535), .C2(n19778), .A(n19528), .B(n19527), .ZN(
        P3_U2902) );
  AOI22_X1 U22631 ( .A1(n19560), .A2(n19819), .B1(n19538), .B2(n19820), .ZN(
        n19530) );
  AOI22_X1 U22632 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19540), .B1(
        n9683), .B2(n19822), .ZN(n19529) );
  OAI211_X1 U22633 ( .C1(n19535), .C2(n19826), .A(n19530), .B(n19529), .ZN(
        P3_U2903) );
  AOI22_X1 U22634 ( .A1(n19560), .A2(n19829), .B1(n19538), .B2(n19827), .ZN(
        n19532) );
  AOI22_X1 U22635 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19540), .B1(
        n9683), .B2(n19720), .ZN(n19531) );
  OAI211_X1 U22636 ( .C1(n19535), .C2(n19723), .A(n19532), .B(n19531), .ZN(
        P3_U2904) );
  AOI22_X1 U22637 ( .A1(n19560), .A2(n19835), .B1(n19538), .B2(n19833), .ZN(
        n19534) );
  AOI22_X1 U22638 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19540), .B1(
        n9683), .B2(n19749), .ZN(n19533) );
  OAI211_X1 U22639 ( .C1(n19535), .C2(n19753), .A(n19534), .B(n19533), .ZN(
        P3_U2905) );
  AOI22_X1 U22640 ( .A1(n19539), .A2(n19841), .B1(n19538), .B2(n19839), .ZN(
        n19537) );
  AOI22_X1 U22641 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19540), .B1(
        n19560), .B2(n19840), .ZN(n19536) );
  OAI211_X1 U22642 ( .C1(n19600), .C2(n19844), .A(n19537), .B(n19536), .ZN(
        P3_U2906) );
  AOI22_X1 U22643 ( .A1(n19539), .A2(n19850), .B1(n19538), .B2(n19846), .ZN(
        n19542) );
  AOI22_X1 U22644 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19540), .B1(
        n19560), .B2(n19848), .ZN(n19541) );
  OAI211_X1 U22645 ( .C1(n19600), .C2(n19855), .A(n19542), .B(n19541), .ZN(
        P3_U2907) );
  INV_X1 U22646 ( .A(n19797), .ZN(n19768) );
  NOR2_X1 U22647 ( .A1(n19589), .A2(n19734), .ZN(n19559) );
  AOI22_X1 U22648 ( .A1(n19760), .A2(n19560), .B1(n19796), .B2(n19559), .ZN(
        n19545) );
  AOI22_X1 U22649 ( .A1(n19801), .A2(n19543), .B1(n19588), .B2(n19736), .ZN(
        n19561) );
  NOR2_X2 U22650 ( .A1(n19637), .A2(n19589), .ZN(n19628) );
  AOI22_X1 U22651 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19561), .B1(
        n19802), .B2(n19628), .ZN(n19544) );
  OAI211_X1 U22652 ( .C1(n19579), .C2(n19768), .A(n19545), .B(n19544), .ZN(
        P3_U2908) );
  AOI22_X1 U22653 ( .A1(n19560), .A2(n19807), .B1(n19806), .B2(n19559), .ZN(
        n19547) );
  AOI22_X1 U22654 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19561), .B1(
        n19808), .B2(n19628), .ZN(n19546) );
  OAI211_X1 U22655 ( .C1(n19579), .C2(n19812), .A(n19547), .B(n19546), .ZN(
        P3_U2909) );
  AOI22_X1 U22656 ( .A1(n19583), .A2(n19815), .B1(n19813), .B2(n19559), .ZN(
        n19549) );
  AOI22_X1 U22657 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19561), .B1(
        n19774), .B2(n19628), .ZN(n19548) );
  OAI211_X1 U22658 ( .C1(n19556), .C2(n19778), .A(n19549), .B(n19548), .ZN(
        P3_U2910) );
  AOI22_X1 U22659 ( .A1(n19583), .A2(n19819), .B1(n19820), .B2(n19559), .ZN(
        n19551) );
  AOI22_X1 U22660 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19561), .B1(
        n19822), .B2(n19628), .ZN(n19550) );
  OAI211_X1 U22661 ( .C1(n19556), .C2(n19826), .A(n19551), .B(n19550), .ZN(
        P3_U2911) );
  INV_X1 U22662 ( .A(n19628), .ZN(n19625) );
  AOI22_X1 U22663 ( .A1(n19560), .A2(n19828), .B1(n19827), .B2(n19559), .ZN(
        n19553) );
  AOI22_X1 U22664 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19561), .B1(
        n19583), .B2(n19829), .ZN(n19552) );
  OAI211_X1 U22665 ( .C1(n19832), .C2(n19625), .A(n19553), .B(n19552), .ZN(
        P3_U2912) );
  AOI22_X1 U22666 ( .A1(n19583), .A2(n19835), .B1(n19833), .B2(n19559), .ZN(
        n19555) );
  AOI22_X1 U22667 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19561), .B1(
        n19749), .B2(n19628), .ZN(n19554) );
  OAI211_X1 U22668 ( .C1(n19556), .C2(n19753), .A(n19555), .B(n19554), .ZN(
        P3_U2913) );
  AOI22_X1 U22669 ( .A1(n19583), .A2(n19840), .B1(n19839), .B2(n19559), .ZN(
        n19558) );
  AOI22_X1 U22670 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19561), .B1(
        n19560), .B2(n19841), .ZN(n19557) );
  OAI211_X1 U22671 ( .C1(n19844), .C2(n19625), .A(n19558), .B(n19557), .ZN(
        P3_U2914) );
  AOI22_X1 U22672 ( .A1(n19560), .A2(n19850), .B1(n19846), .B2(n19559), .ZN(
        n19563) );
  AOI22_X1 U22673 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19561), .B1(
        n19583), .B2(n19848), .ZN(n19562) );
  OAI211_X1 U22674 ( .C1(n19855), .C2(n19625), .A(n19563), .B(n19562), .ZN(
        P3_U2915) );
  NAND2_X1 U22675 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19588), .ZN(
        n19635) );
  NOR2_X1 U22676 ( .A1(n19628), .A2(n19656), .ZN(n19610) );
  NOR2_X1 U22677 ( .A1(n19918), .A2(n19610), .ZN(n19582) );
  AOI22_X1 U22678 ( .A1(n19760), .A2(n19583), .B1(n19796), .B2(n19582), .ZN(
        n19568) );
  NOR2_X1 U22679 ( .A1(n9683), .A2(n19583), .ZN(n19565) );
  AOI221_X1 U22680 ( .B1(n19610), .B2(n19762), .C1(n19610), .C2(n19565), .A(
        n19564), .ZN(n19566) );
  INV_X1 U22681 ( .A(n19566), .ZN(n19584) );
  AOI22_X1 U22682 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19584), .B1(
        n19802), .B2(n19656), .ZN(n19567) );
  OAI211_X1 U22683 ( .C1(n19600), .C2(n19768), .A(n19568), .B(n19567), .ZN(
        P3_U2916) );
  AOI22_X1 U22684 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19584), .B1(
        n19806), .B2(n19582), .ZN(n19570) );
  AOI22_X1 U22685 ( .A1(n9683), .A2(n19769), .B1(n19808), .B2(n19656), .ZN(
        n19569) );
  OAI211_X1 U22686 ( .C1(n19579), .C2(n19772), .A(n19570), .B(n19569), .ZN(
        P3_U2917) );
  AOI22_X1 U22687 ( .A1(n9683), .A2(n19815), .B1(n19813), .B2(n19582), .ZN(
        n19572) );
  AOI22_X1 U22688 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19584), .B1(
        n19774), .B2(n19656), .ZN(n19571) );
  OAI211_X1 U22689 ( .C1(n19579), .C2(n19778), .A(n19572), .B(n19571), .ZN(
        P3_U2918) );
  INV_X1 U22690 ( .A(n19656), .ZN(n19614) );
  AOI22_X1 U22691 ( .A1(n19583), .A2(n19779), .B1(n19820), .B2(n19582), .ZN(
        n19574) );
  AOI22_X1 U22692 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19584), .B1(
        n9683), .B2(n19819), .ZN(n19573) );
  OAI211_X1 U22693 ( .C1(n19782), .C2(n19614), .A(n19574), .B(n19573), .ZN(
        P3_U2919) );
  AOI22_X1 U22694 ( .A1(n19583), .A2(n19828), .B1(n19827), .B2(n19582), .ZN(
        n19576) );
  AOI22_X1 U22695 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19584), .B1(
        n9683), .B2(n19829), .ZN(n19575) );
  OAI211_X1 U22696 ( .C1(n19832), .C2(n19614), .A(n19576), .B(n19575), .ZN(
        P3_U2920) );
  AOI22_X1 U22697 ( .A1(n9683), .A2(n19835), .B1(n19833), .B2(n19582), .ZN(
        n19578) );
  AOI22_X1 U22698 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19584), .B1(
        n19749), .B2(n19656), .ZN(n19577) );
  OAI211_X1 U22699 ( .C1(n19579), .C2(n19753), .A(n19578), .B(n19577), .ZN(
        P3_U2921) );
  AOI22_X1 U22700 ( .A1(n9683), .A2(n19840), .B1(n19839), .B2(n19582), .ZN(
        n19581) );
  AOI22_X1 U22701 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19584), .B1(
        n19583), .B2(n19841), .ZN(n19580) );
  OAI211_X1 U22702 ( .C1(n19844), .C2(n19614), .A(n19581), .B(n19580), .ZN(
        P3_U2922) );
  AOI22_X1 U22703 ( .A1(n19583), .A2(n19850), .B1(n19846), .B2(n19582), .ZN(
        n19586) );
  AOI22_X1 U22704 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19584), .B1(
        n9683), .B2(n19848), .ZN(n19585) );
  OAI211_X1 U22705 ( .C1(n19855), .C2(n19614), .A(n19586), .B(n19585), .ZN(
        P3_U2923) );
  NOR2_X1 U22706 ( .A1(n19918), .A2(n19635), .ZN(n19605) );
  AOI22_X1 U22707 ( .A1(n19760), .A2(n9683), .B1(n19796), .B2(n19605), .ZN(
        n19591) );
  AOI21_X1 U22708 ( .B1(n19858), .B2(n19762), .A(n19634), .ZN(n19587) );
  NAND2_X1 U22709 ( .A1(n19588), .A2(n19587), .ZN(n19607) );
  NOR2_X2 U22710 ( .A1(n19860), .A2(n19589), .ZN(n19683) );
  AOI22_X1 U22711 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19607), .B1(
        n19802), .B2(n19683), .ZN(n19590) );
  OAI211_X1 U22712 ( .C1(n19768), .C2(n19625), .A(n19591), .B(n19590), .ZN(
        P3_U2924) );
  AOI22_X1 U22713 ( .A1(n19806), .A2(n19605), .B1(n19769), .B2(n19628), .ZN(
        n19593) );
  AOI22_X1 U22714 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19607), .B1(
        n19808), .B2(n19683), .ZN(n19592) );
  OAI211_X1 U22715 ( .C1(n19600), .C2(n19772), .A(n19593), .B(n19592), .ZN(
        P3_U2925) );
  INV_X1 U22716 ( .A(n19683), .ZN(n19678) );
  AOI22_X1 U22717 ( .A1(n9683), .A2(n19814), .B1(n19813), .B2(n19605), .ZN(
        n19595) );
  AOI22_X1 U22718 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19607), .B1(
        n19815), .B2(n19628), .ZN(n19594) );
  OAI211_X1 U22719 ( .C1(n19818), .C2(n19678), .A(n19595), .B(n19594), .ZN(
        P3_U2926) );
  AOI22_X1 U22720 ( .A1(n9683), .A2(n19779), .B1(n19820), .B2(n19605), .ZN(
        n19597) );
  AOI22_X1 U22721 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19607), .B1(
        n19819), .B2(n19628), .ZN(n19596) );
  OAI211_X1 U22722 ( .C1(n19782), .C2(n19678), .A(n19597), .B(n19596), .ZN(
        P3_U2927) );
  AOI22_X1 U22723 ( .A1(n19829), .A2(n19628), .B1(n19827), .B2(n19605), .ZN(
        n19599) );
  AOI22_X1 U22724 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19607), .B1(
        n19720), .B2(n19683), .ZN(n19598) );
  OAI211_X1 U22725 ( .C1(n19600), .C2(n19723), .A(n19599), .B(n19598), .ZN(
        P3_U2928) );
  AOI22_X1 U22726 ( .A1(n9683), .A2(n19834), .B1(n19833), .B2(n19605), .ZN(
        n19602) );
  AOI22_X1 U22727 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19607), .B1(
        n19835), .B2(n19628), .ZN(n19601) );
  OAI211_X1 U22728 ( .C1(n19838), .C2(n19678), .A(n19602), .B(n19601), .ZN(
        P3_U2929) );
  AOI22_X1 U22729 ( .A1(n9683), .A2(n19841), .B1(n19839), .B2(n19605), .ZN(
        n19604) );
  AOI22_X1 U22730 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19607), .B1(
        n19840), .B2(n19628), .ZN(n19603) );
  OAI211_X1 U22731 ( .C1(n19844), .C2(n19678), .A(n19604), .B(n19603), .ZN(
        P3_U2930) );
  AOI22_X1 U22732 ( .A1(n9683), .A2(n19850), .B1(n19846), .B2(n19605), .ZN(
        n19609) );
  AOI22_X1 U22733 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19607), .B1(
        n19848), .B2(n19628), .ZN(n19608) );
  OAI211_X1 U22734 ( .C1(n19855), .C2(n19678), .A(n19609), .B(n19608), .ZN(
        P3_U2931) );
  NOR2_X2 U22735 ( .A1(n19864), .A2(n19689), .ZN(n19706) );
  NOR2_X1 U22736 ( .A1(n19683), .A2(n19706), .ZN(n19666) );
  NOR2_X1 U22737 ( .A1(n19918), .A2(n19666), .ZN(n19629) );
  AOI22_X1 U22738 ( .A1(n19760), .A2(n19628), .B1(n19796), .B2(n19629), .ZN(
        n19613) );
  OAI21_X1 U22739 ( .B1(n19610), .B2(n19762), .A(n19666), .ZN(n19611) );
  OAI211_X1 U22740 ( .C1(n19706), .C2(n20016), .A(n19765), .B(n19611), .ZN(
        n19630) );
  AOI22_X1 U22741 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19630), .B1(
        n19802), .B2(n19706), .ZN(n19612) );
  OAI211_X1 U22742 ( .C1(n19768), .C2(n19614), .A(n19613), .B(n19612), .ZN(
        P3_U2932) );
  AOI22_X1 U22743 ( .A1(n19806), .A2(n19629), .B1(n19769), .B2(n19656), .ZN(
        n19616) );
  AOI22_X1 U22744 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19630), .B1(
        n19808), .B2(n19706), .ZN(n19615) );
  OAI211_X1 U22745 ( .C1(n19772), .C2(n19625), .A(n19616), .B(n19615), .ZN(
        P3_U2933) );
  AOI22_X1 U22746 ( .A1(n19815), .A2(n19656), .B1(n19813), .B2(n19629), .ZN(
        n19618) );
  AOI22_X1 U22747 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19630), .B1(
        n19774), .B2(n19706), .ZN(n19617) );
  OAI211_X1 U22748 ( .C1(n19778), .C2(n19625), .A(n19618), .B(n19617), .ZN(
        P3_U2934) );
  AOI22_X1 U22749 ( .A1(n19820), .A2(n19629), .B1(n19819), .B2(n19656), .ZN(
        n19620) );
  AOI22_X1 U22750 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19630), .B1(
        n19822), .B2(n19706), .ZN(n19619) );
  OAI211_X1 U22751 ( .C1(n19826), .C2(n19625), .A(n19620), .B(n19619), .ZN(
        P3_U2935) );
  AOI22_X1 U22752 ( .A1(n19829), .A2(n19656), .B1(n19827), .B2(n19629), .ZN(
        n19622) );
  AOI22_X1 U22753 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19630), .B1(
        n19720), .B2(n19706), .ZN(n19621) );
  OAI211_X1 U22754 ( .C1(n19723), .C2(n19625), .A(n19622), .B(n19621), .ZN(
        P3_U2936) );
  AOI22_X1 U22755 ( .A1(n19835), .A2(n19656), .B1(n19833), .B2(n19629), .ZN(
        n19624) );
  AOI22_X1 U22756 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19630), .B1(
        n19749), .B2(n19706), .ZN(n19623) );
  OAI211_X1 U22757 ( .C1(n19753), .C2(n19625), .A(n19624), .B(n19623), .ZN(
        P3_U2937) );
  INV_X1 U22758 ( .A(n19706), .ZN(n19702) );
  AOI22_X1 U22759 ( .A1(n19839), .A2(n19629), .B1(n19841), .B2(n19628), .ZN(
        n19627) );
  AOI22_X1 U22760 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19630), .B1(
        n19840), .B2(n19656), .ZN(n19626) );
  OAI211_X1 U22761 ( .C1(n19844), .C2(n19702), .A(n19627), .B(n19626), .ZN(
        P3_U2938) );
  AOI22_X1 U22762 ( .A1(n19846), .A2(n19629), .B1(n19850), .B2(n19628), .ZN(
        n19632) );
  AOI22_X1 U22763 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19630), .B1(
        n19848), .B2(n19656), .ZN(n19631) );
  OAI211_X1 U22764 ( .C1(n19855), .C2(n19702), .A(n19632), .B(n19631), .ZN(
        P3_U2939) );
  NAND2_X1 U22765 ( .A1(n19688), .A2(n19858), .ZN(n19633) );
  OAI22_X1 U22766 ( .A1(n19636), .A2(n19635), .B1(n19634), .B2(n19633), .ZN(
        n19662) );
  NOR2_X1 U22767 ( .A1(n19689), .A2(n19734), .ZN(n19661) );
  AOI22_X1 U22768 ( .A1(n19760), .A2(n19656), .B1(n19796), .B2(n19661), .ZN(
        n19639) );
  NOR2_X2 U22769 ( .A1(n19637), .A2(n19689), .ZN(n19730) );
  AOI22_X1 U22770 ( .A1(n19802), .A2(n19730), .B1(n19797), .B2(n19683), .ZN(
        n19638) );
  OAI211_X1 U22771 ( .C1(n19640), .C2(n19662), .A(n19639), .B(n19638), .ZN(
        P3_U2940) );
  AOI22_X1 U22772 ( .A1(n19807), .A2(n19656), .B1(n19806), .B2(n19661), .ZN(
        n19642) );
  AOI22_X1 U22773 ( .A1(n19808), .A2(n19730), .B1(n19769), .B2(n19683), .ZN(
        n19641) );
  OAI211_X1 U22774 ( .C1(n19643), .C2(n19662), .A(n19642), .B(n19641), .ZN(
        P3_U2941) );
  AOI22_X1 U22775 ( .A1(n19815), .A2(n19683), .B1(n19813), .B2(n19661), .ZN(
        n19645) );
  AOI22_X1 U22776 ( .A1(n19814), .A2(n19656), .B1(n19774), .B2(n19730), .ZN(
        n19644) );
  OAI211_X1 U22777 ( .C1(n19646), .C2(n19662), .A(n19645), .B(n19644), .ZN(
        P3_U2942) );
  AOI22_X1 U22778 ( .A1(n19779), .A2(n19656), .B1(n19820), .B2(n19661), .ZN(
        n19648) );
  AOI22_X1 U22779 ( .A1(n19822), .A2(n19730), .B1(n19819), .B2(n19683), .ZN(
        n19647) );
  OAI211_X1 U22780 ( .C1(n19649), .C2(n19662), .A(n19648), .B(n19647), .ZN(
        P3_U2943) );
  AOI22_X1 U22781 ( .A1(n19828), .A2(n19656), .B1(n19827), .B2(n19661), .ZN(
        n19651) );
  AOI22_X1 U22782 ( .A1(n19720), .A2(n19730), .B1(n19829), .B2(n19683), .ZN(
        n19650) );
  OAI211_X1 U22783 ( .C1(n19652), .C2(n19662), .A(n19651), .B(n19650), .ZN(
        P3_U2944) );
  AOI22_X1 U22784 ( .A1(n19835), .A2(n19683), .B1(n19833), .B2(n19661), .ZN(
        n19654) );
  AOI22_X1 U22785 ( .A1(n19834), .A2(n19656), .B1(n19749), .B2(n19730), .ZN(
        n19653) );
  OAI211_X1 U22786 ( .C1(n19655), .C2(n19662), .A(n19654), .B(n19653), .ZN(
        P3_U2945) );
  INV_X1 U22787 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n19660) );
  AOI22_X1 U22788 ( .A1(n19839), .A2(n19661), .B1(n19841), .B2(n19656), .ZN(
        n19659) );
  AOI22_X1 U22789 ( .A1(n19840), .A2(n19683), .B1(n19657), .B2(n19730), .ZN(
        n19658) );
  OAI211_X1 U22790 ( .C1(n19660), .C2(n19662), .A(n19659), .B(n19658), .ZN(
        P3_U2946) );
  INV_X1 U22791 ( .A(n19730), .ZN(n19726) );
  AOI22_X1 U22792 ( .A1(n19846), .A2(n19661), .B1(n19850), .B2(n19656), .ZN(
        n19665) );
  INV_X1 U22793 ( .A(n19662), .ZN(n19663) );
  AOI22_X1 U22794 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19663), .B1(
        n19848), .B2(n19683), .ZN(n19664) );
  OAI211_X1 U22795 ( .C1(n19855), .C2(n19726), .A(n19665), .B(n19664), .ZN(
        P3_U2947) );
  NOR2_X1 U22796 ( .A1(n19858), .A2(n19689), .ZN(n19738) );
  NAND2_X1 U22797 ( .A1(n12049), .A2(n19738), .ZN(n19752) );
  NOR2_X1 U22798 ( .A1(n19730), .A2(n19756), .ZN(n19710) );
  OAI21_X1 U22799 ( .B1(n19666), .B2(n19762), .A(n19710), .ZN(n19667) );
  OAI211_X1 U22800 ( .C1(n19756), .C2(n20016), .A(n19765), .B(n19667), .ZN(
        n19685) );
  NOR2_X1 U22801 ( .A1(n19918), .A2(n19710), .ZN(n19684) );
  AOI22_X1 U22802 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19685), .B1(
        n19796), .B2(n19684), .ZN(n19669) );
  AOI22_X1 U22803 ( .A1(n19802), .A2(n19756), .B1(n19797), .B2(n19706), .ZN(
        n19668) );
  OAI211_X1 U22804 ( .C1(n19805), .C2(n19678), .A(n19669), .B(n19668), .ZN(
        P3_U2948) );
  AOI22_X1 U22805 ( .A1(n19806), .A2(n19684), .B1(n19769), .B2(n19706), .ZN(
        n19671) );
  AOI22_X1 U22806 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19685), .B1(
        n19808), .B2(n19756), .ZN(n19670) );
  OAI211_X1 U22807 ( .C1(n19772), .C2(n19678), .A(n19671), .B(n19670), .ZN(
        P3_U2949) );
  AOI22_X1 U22808 ( .A1(n19814), .A2(n19683), .B1(n19813), .B2(n19684), .ZN(
        n19673) );
  AOI22_X1 U22809 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19685), .B1(
        n19815), .B2(n19706), .ZN(n19672) );
  OAI211_X1 U22810 ( .C1(n19818), .C2(n19752), .A(n19673), .B(n19672), .ZN(
        P3_U2950) );
  AOI22_X1 U22811 ( .A1(n19779), .A2(n19683), .B1(n19820), .B2(n19684), .ZN(
        n19675) );
  AOI22_X1 U22812 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19685), .B1(
        n19819), .B2(n19706), .ZN(n19674) );
  OAI211_X1 U22813 ( .C1(n19782), .C2(n19752), .A(n19675), .B(n19674), .ZN(
        P3_U2951) );
  AOI22_X1 U22814 ( .A1(n19829), .A2(n19706), .B1(n19827), .B2(n19684), .ZN(
        n19677) );
  AOI22_X1 U22815 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19685), .B1(
        n19720), .B2(n19756), .ZN(n19676) );
  OAI211_X1 U22816 ( .C1(n19723), .C2(n19678), .A(n19677), .B(n19676), .ZN(
        P3_U2952) );
  AOI22_X1 U22817 ( .A1(n19834), .A2(n19683), .B1(n19833), .B2(n19684), .ZN(
        n19680) );
  AOI22_X1 U22818 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19685), .B1(
        n19835), .B2(n19706), .ZN(n19679) );
  OAI211_X1 U22819 ( .C1(n19838), .C2(n19752), .A(n19680), .B(n19679), .ZN(
        P3_U2953) );
  AOI22_X1 U22820 ( .A1(n19839), .A2(n19684), .B1(n19841), .B2(n19683), .ZN(
        n19682) );
  AOI22_X1 U22821 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19685), .B1(
        n19840), .B2(n19706), .ZN(n19681) );
  OAI211_X1 U22822 ( .C1(n19844), .C2(n19752), .A(n19682), .B(n19681), .ZN(
        P3_U2954) );
  AOI22_X1 U22823 ( .A1(n19846), .A2(n19684), .B1(n19850), .B2(n19683), .ZN(
        n19687) );
  AOI22_X1 U22824 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19685), .B1(
        n19848), .B2(n19706), .ZN(n19686) );
  OAI211_X1 U22825 ( .C1(n19855), .C2(n19752), .A(n19687), .B(n19686), .ZN(
        P3_U2955) );
  AND2_X1 U22826 ( .A1(n19907), .A2(n19738), .ZN(n19705) );
  AOI22_X1 U22827 ( .A1(n19760), .A2(n19706), .B1(n19796), .B2(n19705), .ZN(
        n19691) );
  OAI211_X1 U22828 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n19801), .A(
        n19798), .B(n19688), .ZN(n19707) );
  NOR2_X2 U22829 ( .A1(n19860), .A2(n19689), .ZN(n19790) );
  AOI22_X1 U22830 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19707), .B1(
        n19802), .B2(n19790), .ZN(n19690) );
  OAI211_X1 U22831 ( .C1(n19768), .C2(n19726), .A(n19691), .B(n19690), .ZN(
        P3_U2956) );
  AOI22_X1 U22832 ( .A1(n19806), .A2(n19705), .B1(n19769), .B2(n19730), .ZN(
        n19693) );
  AOI22_X1 U22833 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19707), .B1(
        n19808), .B2(n19790), .ZN(n19692) );
  OAI211_X1 U22834 ( .C1(n19772), .C2(n19702), .A(n19693), .B(n19692), .ZN(
        P3_U2957) );
  AOI22_X1 U22835 ( .A1(n19815), .A2(n19730), .B1(n19813), .B2(n19705), .ZN(
        n19695) );
  AOI22_X1 U22836 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19707), .B1(
        n19774), .B2(n19790), .ZN(n19694) );
  OAI211_X1 U22837 ( .C1(n19778), .C2(n19702), .A(n19695), .B(n19694), .ZN(
        P3_U2958) );
  AOI22_X1 U22838 ( .A1(n19820), .A2(n19705), .B1(n19819), .B2(n19730), .ZN(
        n19697) );
  AOI22_X1 U22839 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19707), .B1(
        n19822), .B2(n19790), .ZN(n19696) );
  OAI211_X1 U22840 ( .C1(n19826), .C2(n19702), .A(n19697), .B(n19696), .ZN(
        P3_U2959) );
  AOI22_X1 U22841 ( .A1(n19829), .A2(n19730), .B1(n19827), .B2(n19705), .ZN(
        n19699) );
  AOI22_X1 U22842 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19707), .B1(
        n19720), .B2(n19790), .ZN(n19698) );
  OAI211_X1 U22843 ( .C1(n19723), .C2(n19702), .A(n19699), .B(n19698), .ZN(
        P3_U2960) );
  AOI22_X1 U22844 ( .A1(n19835), .A2(n19730), .B1(n19833), .B2(n19705), .ZN(
        n19701) );
  AOI22_X1 U22845 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19707), .B1(
        n19749), .B2(n19790), .ZN(n19700) );
  OAI211_X1 U22846 ( .C1(n19753), .C2(n19702), .A(n19701), .B(n19700), .ZN(
        P3_U2961) );
  INV_X1 U22847 ( .A(n19790), .ZN(n19777) );
  AOI22_X1 U22848 ( .A1(n19839), .A2(n19705), .B1(n19841), .B2(n19706), .ZN(
        n19704) );
  AOI22_X1 U22849 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19707), .B1(
        n19840), .B2(n19730), .ZN(n19703) );
  OAI211_X1 U22850 ( .C1(n19844), .C2(n19777), .A(n19704), .B(n19703), .ZN(
        P3_U2962) );
  AOI22_X1 U22851 ( .A1(n19848), .A2(n19730), .B1(n19846), .B2(n19705), .ZN(
        n19709) );
  AOI22_X1 U22852 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19707), .B1(
        n19850), .B2(n19706), .ZN(n19708) );
  OAI211_X1 U22853 ( .C1(n19855), .C2(n19777), .A(n19709), .B(n19708), .ZN(
        P3_U2963) );
  NOR2_X1 U22854 ( .A1(n19790), .A2(n9684), .ZN(n19763) );
  NOR2_X1 U22855 ( .A1(n19918), .A2(n19763), .ZN(n19729) );
  AOI22_X1 U22856 ( .A1(n19797), .A2(n19756), .B1(n19796), .B2(n19729), .ZN(
        n19713) );
  OAI21_X1 U22857 ( .B1(n19710), .B2(n19762), .A(n19763), .ZN(n19711) );
  OAI211_X1 U22858 ( .C1(n9684), .C2(n20016), .A(n19765), .B(n19711), .ZN(
        n19731) );
  AOI22_X1 U22859 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19731), .B1(
        n19802), .B2(n9684), .ZN(n19712) );
  OAI211_X1 U22860 ( .C1(n19805), .C2(n19726), .A(n19713), .B(n19712), .ZN(
        P3_U2964) );
  AOI22_X1 U22861 ( .A1(n19806), .A2(n19729), .B1(n19769), .B2(n19756), .ZN(
        n19715) );
  AOI22_X1 U22862 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19731), .B1(
        n19808), .B2(n9684), .ZN(n19714) );
  OAI211_X1 U22863 ( .C1(n19772), .C2(n19726), .A(n19715), .B(n19714), .ZN(
        P3_U2965) );
  AOI22_X1 U22864 ( .A1(n19815), .A2(n19756), .B1(n19813), .B2(n19729), .ZN(
        n19717) );
  AOI22_X1 U22865 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19731), .B1(
        n19774), .B2(n9684), .ZN(n19716) );
  OAI211_X1 U22866 ( .C1(n19778), .C2(n19726), .A(n19717), .B(n19716), .ZN(
        P3_U2966) );
  AOI22_X1 U22867 ( .A1(n19820), .A2(n19729), .B1(n19819), .B2(n19756), .ZN(
        n19719) );
  AOI22_X1 U22868 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19731), .B1(
        n19822), .B2(n9684), .ZN(n19718) );
  OAI211_X1 U22869 ( .C1(n19826), .C2(n19726), .A(n19719), .B(n19718), .ZN(
        P3_U2967) );
  AOI22_X1 U22870 ( .A1(n19829), .A2(n19756), .B1(n19827), .B2(n19729), .ZN(
        n19722) );
  AOI22_X1 U22871 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19731), .B1(
        n19720), .B2(n9684), .ZN(n19721) );
  OAI211_X1 U22872 ( .C1(n19723), .C2(n19726), .A(n19722), .B(n19721), .ZN(
        P3_U2968) );
  AOI22_X1 U22873 ( .A1(n19835), .A2(n19756), .B1(n19833), .B2(n19729), .ZN(
        n19725) );
  AOI22_X1 U22874 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19731), .B1(
        n19749), .B2(n9684), .ZN(n19724) );
  OAI211_X1 U22875 ( .C1(n19753), .C2(n19726), .A(n19725), .B(n19724), .ZN(
        P3_U2969) );
  INV_X1 U22876 ( .A(n9684), .ZN(n19825) );
  AOI22_X1 U22877 ( .A1(n19840), .A2(n19756), .B1(n19839), .B2(n19729), .ZN(
        n19728) );
  AOI22_X1 U22878 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19731), .B1(
        n19841), .B2(n19730), .ZN(n19727) );
  OAI211_X1 U22879 ( .C1(n19844), .C2(n19825), .A(n19728), .B(n19727), .ZN(
        P3_U2970) );
  AOI22_X1 U22880 ( .A1(n19848), .A2(n19756), .B1(n19846), .B2(n19729), .ZN(
        n19733) );
  AOI22_X1 U22881 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19731), .B1(
        n19850), .B2(n19730), .ZN(n19732) );
  OAI211_X1 U22882 ( .C1(n19855), .C2(n19825), .A(n19733), .B(n19732), .ZN(
        P3_U2971) );
  NOR2_X1 U22883 ( .A1(n19735), .A2(n19734), .ZN(n19800) );
  AOI22_X1 U22884 ( .A1(n19760), .A2(n19756), .B1(n19796), .B2(n19800), .ZN(
        n19740) );
  AOI22_X1 U22885 ( .A1(n19801), .A2(n19738), .B1(n19737), .B2(n19736), .ZN(
        n19757) );
  AOI22_X1 U22886 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19757), .B1(
        n19802), .B2(n19847), .ZN(n19739) );
  OAI211_X1 U22887 ( .C1(n19768), .C2(n19777), .A(n19740), .B(n19739), .ZN(
        P3_U2972) );
  AOI22_X1 U22888 ( .A1(n19807), .A2(n19756), .B1(n19806), .B2(n19800), .ZN(
        n19742) );
  AOI22_X1 U22889 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19757), .B1(
        n19808), .B2(n19847), .ZN(n19741) );
  OAI211_X1 U22890 ( .C1(n19812), .C2(n19777), .A(n19742), .B(n19741), .ZN(
        P3_U2973) );
  INV_X1 U22891 ( .A(n19847), .ZN(n19811) );
  AOI22_X1 U22892 ( .A1(n19814), .A2(n19756), .B1(n19813), .B2(n19800), .ZN(
        n19744) );
  AOI22_X1 U22893 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19757), .B1(
        n19815), .B2(n19790), .ZN(n19743) );
  OAI211_X1 U22894 ( .C1(n19818), .C2(n19811), .A(n19744), .B(n19743), .ZN(
        P3_U2974) );
  AOI22_X1 U22895 ( .A1(n19820), .A2(n19800), .B1(n19819), .B2(n19790), .ZN(
        n19746) );
  AOI22_X1 U22896 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19757), .B1(
        n19822), .B2(n19847), .ZN(n19745) );
  OAI211_X1 U22897 ( .C1(n19826), .C2(n19752), .A(n19746), .B(n19745), .ZN(
        P3_U2975) );
  AOI22_X1 U22898 ( .A1(n19828), .A2(n19756), .B1(n19827), .B2(n19800), .ZN(
        n19748) );
  AOI22_X1 U22899 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19757), .B1(
        n19829), .B2(n19790), .ZN(n19747) );
  OAI211_X1 U22900 ( .C1(n19832), .C2(n19811), .A(n19748), .B(n19747), .ZN(
        P3_U2976) );
  AOI22_X1 U22901 ( .A1(n19835), .A2(n19790), .B1(n19833), .B2(n19800), .ZN(
        n19751) );
  AOI22_X1 U22902 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19757), .B1(
        n19749), .B2(n19847), .ZN(n19750) );
  OAI211_X1 U22903 ( .C1(n19753), .C2(n19752), .A(n19751), .B(n19750), .ZN(
        P3_U2977) );
  AOI22_X1 U22904 ( .A1(n19839), .A2(n19800), .B1(n19841), .B2(n19756), .ZN(
        n19755) );
  AOI22_X1 U22905 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19757), .B1(
        n19840), .B2(n19790), .ZN(n19754) );
  OAI211_X1 U22906 ( .C1(n19844), .C2(n19811), .A(n19755), .B(n19754), .ZN(
        P3_U2978) );
  AOI22_X1 U22907 ( .A1(n19846), .A2(n19800), .B1(n19850), .B2(n19756), .ZN(
        n19759) );
  AOI22_X1 U22908 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19757), .B1(
        n19848), .B2(n19790), .ZN(n19758) );
  OAI211_X1 U22909 ( .C1(n19855), .C2(n19811), .A(n19759), .B(n19758), .ZN(
        P3_U2979) );
  NOR2_X1 U22910 ( .A1(n19918), .A2(n19761), .ZN(n19789) );
  AOI22_X1 U22911 ( .A1(n19760), .A2(n19790), .B1(n19796), .B2(n19789), .ZN(
        n19767) );
  OAI21_X1 U22912 ( .B1(n19763), .B2(n19762), .A(n19761), .ZN(n19764) );
  OAI211_X1 U22913 ( .C1(n19773), .C2(n20016), .A(n19765), .B(n19764), .ZN(
        n19791) );
  AOI22_X1 U22914 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19791), .B1(
        n19802), .B2(n19773), .ZN(n19766) );
  OAI211_X1 U22915 ( .C1(n19768), .C2(n19825), .A(n19767), .B(n19766), .ZN(
        P3_U2980) );
  AOI22_X1 U22916 ( .A1(n19806), .A2(n19789), .B1(n19769), .B2(n9684), .ZN(
        n19771) );
  AOI22_X1 U22917 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19791), .B1(
        n19808), .B2(n19773), .ZN(n19770) );
  OAI211_X1 U22918 ( .C1(n19772), .C2(n19777), .A(n19771), .B(n19770), .ZN(
        P3_U2981) );
  AOI22_X1 U22919 ( .A1(n19815), .A2(n9684), .B1(n19813), .B2(n19789), .ZN(
        n19776) );
  AOI22_X1 U22920 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19791), .B1(
        n19774), .B2(n19773), .ZN(n19775) );
  OAI211_X1 U22921 ( .C1(n19778), .C2(n19777), .A(n19776), .B(n19775), .ZN(
        P3_U2982) );
  AOI22_X1 U22922 ( .A1(n19779), .A2(n19790), .B1(n19820), .B2(n19789), .ZN(
        n19781) );
  AOI22_X1 U22923 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19791), .B1(
        n19819), .B2(n9684), .ZN(n19780) );
  OAI211_X1 U22924 ( .C1(n19782), .C2(n19794), .A(n19781), .B(n19780), .ZN(
        P3_U2983) );
  AOI22_X1 U22925 ( .A1(n19828), .A2(n19790), .B1(n19827), .B2(n19789), .ZN(
        n19784) );
  AOI22_X1 U22926 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19791), .B1(
        n19829), .B2(n9684), .ZN(n19783) );
  OAI211_X1 U22927 ( .C1(n19832), .C2(n19794), .A(n19784), .B(n19783), .ZN(
        P3_U2984) );
  AOI22_X1 U22928 ( .A1(n19834), .A2(n19790), .B1(n19833), .B2(n19789), .ZN(
        n19786) );
  AOI22_X1 U22929 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19791), .B1(
        n19835), .B2(n9684), .ZN(n19785) );
  OAI211_X1 U22930 ( .C1(n19838), .C2(n19794), .A(n19786), .B(n19785), .ZN(
        P3_U2985) );
  AOI22_X1 U22931 ( .A1(n19839), .A2(n19789), .B1(n19841), .B2(n19790), .ZN(
        n19788) );
  AOI22_X1 U22932 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19791), .B1(
        n19840), .B2(n9684), .ZN(n19787) );
  OAI211_X1 U22933 ( .C1(n19844), .C2(n19794), .A(n19788), .B(n19787), .ZN(
        P3_U2986) );
  AOI22_X1 U22934 ( .A1(n19848), .A2(n9684), .B1(n19846), .B2(n19789), .ZN(
        n19793) );
  AOI22_X1 U22935 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19791), .B1(
        n19850), .B2(n19790), .ZN(n19792) );
  OAI211_X1 U22936 ( .C1(n19855), .C2(n19794), .A(n19793), .B(n19792), .ZN(
        P3_U2987) );
  NOR2_X1 U22937 ( .A1(n19918), .A2(n19795), .ZN(n19845) );
  AOI22_X1 U22938 ( .A1(n19797), .A2(n19847), .B1(n19796), .B2(n19845), .ZN(
        n19804) );
  AOI22_X1 U22939 ( .A1(n19801), .A2(n19800), .B1(n19799), .B2(n19798), .ZN(
        n19851) );
  AOI22_X1 U22940 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19851), .B1(
        n19802), .B2(n19821), .ZN(n19803) );
  OAI211_X1 U22941 ( .C1(n19805), .C2(n19825), .A(n19804), .B(n19803), .ZN(
        P3_U2988) );
  AOI22_X1 U22942 ( .A1(n19807), .A2(n9684), .B1(n19806), .B2(n19845), .ZN(
        n19810) );
  AOI22_X1 U22943 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19851), .B1(
        n19808), .B2(n19821), .ZN(n19809) );
  OAI211_X1 U22944 ( .C1(n19812), .C2(n19811), .A(n19810), .B(n19809), .ZN(
        P3_U2989) );
  AOI22_X1 U22945 ( .A1(n19814), .A2(n9684), .B1(n19813), .B2(n19845), .ZN(
        n19817) );
  AOI22_X1 U22946 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19851), .B1(
        n19815), .B2(n19847), .ZN(n19816) );
  OAI211_X1 U22947 ( .C1(n19818), .C2(n19854), .A(n19817), .B(n19816), .ZN(
        P3_U2990) );
  AOI22_X1 U22948 ( .A1(n19820), .A2(n19845), .B1(n19819), .B2(n19847), .ZN(
        n19824) );
  AOI22_X1 U22949 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19851), .B1(
        n19822), .B2(n19821), .ZN(n19823) );
  OAI211_X1 U22950 ( .C1(n19826), .C2(n19825), .A(n19824), .B(n19823), .ZN(
        P3_U2991) );
  AOI22_X1 U22951 ( .A1(n19828), .A2(n9684), .B1(n19827), .B2(n19845), .ZN(
        n19831) );
  AOI22_X1 U22952 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19851), .B1(
        n19829), .B2(n19847), .ZN(n19830) );
  OAI211_X1 U22953 ( .C1(n19832), .C2(n19854), .A(n19831), .B(n19830), .ZN(
        P3_U2992) );
  AOI22_X1 U22954 ( .A1(n19834), .A2(n9684), .B1(n19833), .B2(n19845), .ZN(
        n19837) );
  AOI22_X1 U22955 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19851), .B1(
        n19835), .B2(n19847), .ZN(n19836) );
  OAI211_X1 U22956 ( .C1(n19838), .C2(n19854), .A(n19837), .B(n19836), .ZN(
        P3_U2993) );
  AOI22_X1 U22957 ( .A1(n19840), .A2(n19847), .B1(n19839), .B2(n19845), .ZN(
        n19843) );
  AOI22_X1 U22958 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19851), .B1(
        n19841), .B2(n9684), .ZN(n19842) );
  OAI211_X1 U22959 ( .C1(n19844), .C2(n19854), .A(n19843), .B(n19842), .ZN(
        P3_U2994) );
  AOI22_X1 U22960 ( .A1(n19848), .A2(n19847), .B1(n19846), .B2(n19845), .ZN(
        n19853) );
  AOI22_X1 U22961 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n9684), .ZN(n19852) );
  OAI211_X1 U22962 ( .C1(n19855), .C2(n19854), .A(n19853), .B(n19852), .ZN(
        P3_U2995) );
  NAND2_X1 U22963 ( .A1(n19897), .A2(n19856), .ZN(n19857) );
  OAI21_X1 U22964 ( .B1(n19897), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n19857), .ZN(n19892) );
  INV_X1 U22965 ( .A(n19861), .ZN(n19863) );
  OAI21_X1 U22966 ( .B1(n19861), .B2(n19860), .A(n19859), .ZN(n19862) );
  OAI21_X1 U22967 ( .B1(n19863), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n19862), .ZN(n19866) );
  INV_X1 U22968 ( .A(n19864), .ZN(n19865) );
  AOI21_X1 U22969 ( .B1(n19897), .B2(n19866), .A(n19865), .ZN(n19867) );
  OAI21_X1 U22970 ( .B1(n19892), .B2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n19867), .ZN(n19869) );
  AOI21_X1 U22971 ( .B1(n19892), .B2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19868) );
  NAND2_X1 U22972 ( .A1(n19869), .A2(n19868), .ZN(n19900) );
  INV_X1 U22973 ( .A(n19870), .ZN(n19873) );
  OAI21_X1 U22974 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n19871), .ZN(n19872) );
  OAI211_X1 U22975 ( .C1(n19874), .C2(n19897), .A(n19873), .B(n19872), .ZN(
        n19887) );
  NOR2_X1 U22976 ( .A1(n19876), .A2(n19875), .ZN(n19877) );
  OAI22_X1 U22977 ( .A1(n19880), .A2(n19879), .B1(n19878), .B2(n19877), .ZN(
        n19881) );
  INV_X1 U22978 ( .A(n19881), .ZN(n19882) );
  OAI21_X1 U22979 ( .B1(n19884), .B2(n19883), .A(n19882), .ZN(n20029) );
  OR2_X1 U22980 ( .A1(n20029), .A2(n19885), .ZN(n19886) );
  NOR2_X1 U22981 ( .A1(n19887), .A2(n19886), .ZN(n19888) );
  OAI21_X1 U22982 ( .B1(n19900), .B2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19888), .ZN(n19902) );
  NAND2_X1 U22983 ( .A1(n19890), .A2(n19889), .ZN(n19891) );
  AND2_X1 U22984 ( .A1(n19892), .A2(n19891), .ZN(n19899) );
  NOR2_X1 U22985 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19893), .ZN(
        n19896) );
  NAND2_X1 U22986 ( .A1(n19897), .A2(n19894), .ZN(n19895) );
  AOI22_X1 U22987 ( .A1(n19897), .A2(n19896), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19895), .ZN(n19898) );
  AOI21_X1 U22988 ( .B1(n19900), .B2(n19899), .A(n19898), .ZN(n19901) );
  INV_X1 U22989 ( .A(n19904), .ZN(n19915) );
  INV_X1 U22990 ( .A(n19903), .ZN(n19906) );
  AOI211_X1 U22991 ( .C1(n19906), .C2(n19905), .A(n19914), .B(n19904), .ZN(
        n19919) );
  NOR2_X1 U22992 ( .A1(n19919), .A2(n20035), .ZN(n20017) );
  NAND2_X1 U22993 ( .A1(n20032), .A2(n20047), .ZN(n19916) );
  OAI211_X1 U22994 ( .C1(P3_STATE2_REG_1__SCAN_IN), .C2(n19907), .A(n20017), 
        .B(n19916), .ZN(n19911) );
  INV_X1 U22995 ( .A(n20034), .ZN(n19908) );
  AOI22_X1 U22996 ( .A1(n19909), .A2(n19908), .B1(n20032), .B2(n20041), .ZN(
        n19910) );
  OAI22_X1 U22997 ( .A1(n19912), .A2(n19911), .B1(P3_STATE2_REG_0__SCAN_IN), 
        .B2(n19910), .ZN(n19913) );
  OAI21_X1 U22998 ( .B1(n19915), .B2(n19914), .A(n19913), .ZN(P3_U2996) );
  NAND2_X1 U22999 ( .A1(n20032), .A2(n20041), .ZN(n19922) );
  INV_X1 U23000 ( .A(n19916), .ZN(n19917) );
  NAND3_X1 U23001 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(n19917), .ZN(n19924) );
  OR4_X1 U23002 ( .A1(n19920), .A2(n19919), .A3(n19918), .A4(n19917), .ZN(
        n19921) );
  NAND4_X1 U23003 ( .A1(n19923), .A2(n19922), .A3(n19924), .A4(n19921), .ZN(
        P3_U2997) );
  AND4_X1 U23004 ( .A1(n20034), .A2(n19925), .A3(n20015), .A4(n19924), .ZN(
        P3_U2998) );
  AND2_X1 U23005 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n20011), .ZN(
        P3_U2999) );
  AND2_X1 U23006 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n20011), .ZN(
        P3_U3000) );
  AND2_X1 U23007 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n20011), .ZN(
        P3_U3001) );
  AND2_X1 U23008 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n20011), .ZN(
        P3_U3002) );
  AND2_X1 U23009 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n20011), .ZN(
        P3_U3003) );
  AND2_X1 U23010 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n20011), .ZN(
        P3_U3004) );
  AND2_X1 U23011 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n20011), .ZN(
        P3_U3005) );
  AND2_X1 U23012 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n20011), .ZN(
        P3_U3006) );
  AND2_X1 U23013 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n20011), .ZN(
        P3_U3007) );
  AND2_X1 U23014 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n20011), .ZN(
        P3_U3008) );
  NOR2_X1 U23015 ( .A1(n19926), .A2(n20014), .ZN(P3_U3009) );
  AND2_X1 U23016 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n20011), .ZN(
        P3_U3010) );
  AND2_X1 U23017 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n20011), .ZN(
        P3_U3011) );
  AND2_X1 U23018 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n20011), .ZN(
        P3_U3012) );
  AND2_X1 U23019 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n20011), .ZN(
        P3_U3013) );
  AND2_X1 U23020 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n20011), .ZN(
        P3_U3014) );
  AND2_X1 U23021 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n20011), .ZN(
        P3_U3015) );
  AND2_X1 U23022 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n20011), .ZN(
        P3_U3016) );
  AND2_X1 U23023 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n20011), .ZN(
        P3_U3017) );
  AND2_X1 U23024 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n20011), .ZN(
        P3_U3018) );
  AND2_X1 U23025 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n20011), .ZN(
        P3_U3019) );
  NOR2_X1 U23026 ( .A1(n19927), .A2(n20014), .ZN(P3_U3020) );
  AND2_X1 U23027 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n20011), .ZN(P3_U3021) );
  AND2_X1 U23028 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n20011), .ZN(P3_U3022) );
  AND2_X1 U23029 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n20011), .ZN(P3_U3023) );
  AND2_X1 U23030 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n20011), .ZN(P3_U3024) );
  AND2_X1 U23031 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n20011), .ZN(P3_U3025) );
  AND2_X1 U23032 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n20011), .ZN(P3_U3026) );
  AND2_X1 U23033 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n20011), .ZN(P3_U3027) );
  AND2_X1 U23034 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n20011), .ZN(P3_U3028) );
  OAI21_X1 U23035 ( .B1(n21647), .B2(n19928), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19929) );
  INV_X1 U23036 ( .A(n19929), .ZN(n19933) );
  AOI21_X1 U23037 ( .B1(n20032), .B2(P3_STATE_REG_1__SCAN_IN), .A(n19930), 
        .ZN(n19939) );
  INV_X1 U23038 ( .A(NA), .ZN(n21653) );
  OAI21_X1 U23039 ( .B1(n21653), .B2(n19931), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n19938) );
  INV_X1 U23040 ( .A(n19938), .ZN(n19932) );
  OAI22_X1 U23041 ( .A1(n19996), .A2(n19933), .B1(n19939), .B2(n19932), .ZN(
        P3_U3029) );
  OAI22_X1 U23042 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(n21647), .B2(n19943), .ZN(n19936)
         );
  OAI21_X1 U23043 ( .B1(P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n19940) );
  NAND2_X1 U23044 ( .A1(n20032), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19935) );
  OAI211_X1 U23045 ( .C1(n19936), .C2(n19940), .A(n19934), .B(n19935), .ZN(
        P3_U3030) );
  INV_X1 U23046 ( .A(n19935), .ZN(n19937) );
  AOI21_X1 U23047 ( .B1(n19937), .B2(n21653), .A(n19936), .ZN(n19941) );
  OAI22_X1 U23048 ( .A1(n19941), .A2(n19940), .B1(n19939), .B2(n19938), .ZN(
        P3_U3031) );
  OAI222_X1 U23049 ( .A1(n20018), .A2(n20002), .B1(n19944), .B2(n19996), .C1(
        n19945), .C2(n19999), .ZN(P3_U3032) );
  OAI222_X1 U23050 ( .A1(n19999), .A2(n19947), .B1(n19946), .B2(n19996), .C1(
        n19945), .C2(n20002), .ZN(P3_U3033) );
  OAI222_X1 U23051 ( .A1(n19999), .A2(n19949), .B1(n19948), .B2(n19996), .C1(
        n19947), .C2(n20002), .ZN(P3_U3034) );
  OAI222_X1 U23052 ( .A1(n19999), .A2(n19952), .B1(n19950), .B2(n19996), .C1(
        n19949), .C2(n20002), .ZN(P3_U3035) );
  OAI222_X1 U23053 ( .A1(n19952), .A2(n20002), .B1(n19951), .B2(n19996), .C1(
        n19953), .C2(n19999), .ZN(P3_U3036) );
  OAI222_X1 U23054 ( .A1(n19999), .A2(n19955), .B1(n19954), .B2(n19996), .C1(
        n19953), .C2(n20002), .ZN(P3_U3037) );
  OAI222_X1 U23055 ( .A1(n19999), .A2(n19958), .B1(n19956), .B2(n19996), .C1(
        n19955), .C2(n20002), .ZN(P3_U3038) );
  OAI222_X1 U23056 ( .A1(n19958), .A2(n20002), .B1(n19957), .B2(n19996), .C1(
        n19959), .C2(n19999), .ZN(P3_U3039) );
  OAI222_X1 U23057 ( .A1(n19999), .A2(n19961), .B1(n19960), .B2(n19996), .C1(
        n19959), .C2(n20002), .ZN(P3_U3040) );
  OAI222_X1 U23058 ( .A1(n19999), .A2(n19963), .B1(n19962), .B2(n19996), .C1(
        n19961), .C2(n20002), .ZN(P3_U3041) );
  OAI222_X1 U23059 ( .A1(n19999), .A2(n19965), .B1(n19964), .B2(n19996), .C1(
        n19963), .C2(n20002), .ZN(P3_U3042) );
  OAI222_X1 U23060 ( .A1(n19999), .A2(n19967), .B1(n19966), .B2(n19996), .C1(
        n19965), .C2(n20002), .ZN(P3_U3043) );
  OAI222_X1 U23061 ( .A1(n19999), .A2(n19970), .B1(n19968), .B2(n19996), .C1(
        n19967), .C2(n20002), .ZN(P3_U3044) );
  OAI222_X1 U23062 ( .A1(n19970), .A2(n20002), .B1(n19969), .B2(n19996), .C1(
        n19971), .C2(n19999), .ZN(P3_U3045) );
  OAI222_X1 U23063 ( .A1(n19999), .A2(n19973), .B1(n19972), .B2(n19996), .C1(
        n19971), .C2(n20002), .ZN(P3_U3046) );
  OAI222_X1 U23064 ( .A1(n19999), .A2(n19976), .B1(n19974), .B2(n19996), .C1(
        n19973), .C2(n20002), .ZN(P3_U3047) );
  OAI222_X1 U23065 ( .A1(n19976), .A2(n20002), .B1(n19975), .B2(n19996), .C1(
        n19977), .C2(n19999), .ZN(P3_U3048) );
  OAI222_X1 U23066 ( .A1(n19999), .A2(n19980), .B1(n19978), .B2(n19996), .C1(
        n19977), .C2(n20002), .ZN(P3_U3049) );
  OAI222_X1 U23067 ( .A1(n19980), .A2(n20002), .B1(n19979), .B2(n19996), .C1(
        n19981), .C2(n19999), .ZN(P3_U3050) );
  OAI222_X1 U23068 ( .A1(n19999), .A2(n19984), .B1(n19982), .B2(n19996), .C1(
        n19981), .C2(n20002), .ZN(P3_U3051) );
  OAI222_X1 U23069 ( .A1(n19984), .A2(n20002), .B1(n19983), .B2(n19996), .C1(
        n19985), .C2(n19999), .ZN(P3_U3052) );
  OAI222_X1 U23070 ( .A1(n19999), .A2(n19988), .B1(n19986), .B2(n19996), .C1(
        n19985), .C2(n20002), .ZN(P3_U3053) );
  OAI222_X1 U23071 ( .A1(n19988), .A2(n20002), .B1(n19987), .B2(n19996), .C1(
        n19989), .C2(n19999), .ZN(P3_U3054) );
  OAI222_X1 U23072 ( .A1(n19999), .A2(n19991), .B1(n19990), .B2(n19996), .C1(
        n19989), .C2(n20002), .ZN(P3_U3055) );
  OAI222_X1 U23073 ( .A1(n19999), .A2(n19993), .B1(n19992), .B2(n19996), .C1(
        n19991), .C2(n20002), .ZN(P3_U3056) );
  OAI222_X1 U23074 ( .A1(n19999), .A2(n17587), .B1(n19994), .B2(n19996), .C1(
        n19993), .C2(n20002), .ZN(P3_U3057) );
  OAI222_X1 U23075 ( .A1(n19999), .A2(n13202), .B1(n19995), .B2(n19996), .C1(
        n17587), .C2(n20002), .ZN(P3_U3058) );
  OAI222_X1 U23076 ( .A1(n13202), .A2(n20002), .B1(n19997), .B2(n19996), .C1(
        n17567), .C2(n19999), .ZN(P3_U3059) );
  OAI222_X1 U23077 ( .A1(n19999), .A2(n17557), .B1(n19998), .B2(n19996), .C1(
        n17567), .C2(n20002), .ZN(P3_U3060) );
  OAI222_X1 U23078 ( .A1(n20002), .A2(n17557), .B1(n20001), .B2(n19996), .C1(
        n20000), .C2(n19999), .ZN(P3_U3061) );
  AOI22_X1 U23079 ( .A1(n19996), .A2(n20004), .B1(n20003), .B2(n20026), .ZN(
        P3_U3274) );
  INV_X1 U23080 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n20005) );
  AOI22_X1 U23081 ( .A1(n19996), .A2(n20021), .B1(n20005), .B2(n20026), .ZN(
        P3_U3275) );
  AOI22_X1 U23082 ( .A1(n19996), .A2(n20007), .B1(n20006), .B2(n20026), .ZN(
        P3_U3276) );
  INV_X1 U23083 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20024) );
  INV_X1 U23084 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n20008) );
  AOI22_X1 U23085 ( .A1(n19996), .A2(n20024), .B1(n20008), .B2(n20026), .ZN(
        P3_U3277) );
  INV_X1 U23086 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20010) );
  INV_X1 U23087 ( .A(n20012), .ZN(n20009) );
  AOI21_X1 U23088 ( .B1(n20011), .B2(n20010), .A(n20009), .ZN(P3_U3280) );
  OAI21_X1 U23089 ( .B1(n20014), .B2(n20013), .A(n20012), .ZN(P3_U3281) );
  OAI21_X1 U23090 ( .B1(n20017), .B2(n20016), .A(n20015), .ZN(P3_U3282) );
  AOI21_X1 U23091 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20019) );
  AOI22_X1 U23092 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n20019), .B2(n20018), .ZN(n20022) );
  AOI22_X1 U23093 ( .A1(n20025), .A2(n20022), .B1(n20021), .B2(n20020), .ZN(
        P3_U3292) );
  OAI21_X1 U23094 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n20025), .ZN(n20023) );
  OAI21_X1 U23095 ( .B1(n20025), .B2(n20024), .A(n20023), .ZN(P3_U3293) );
  INV_X1 U23096 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n20027) );
  AOI22_X1 U23097 ( .A1(n19996), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n20027), 
        .B2(n20026), .ZN(P3_U3294) );
  MUX2_X1 U23098 ( .A(P3_MORE_REG_SCAN_IN), .B(n20029), .S(n20028), .Z(
        P3_U3295) );
  OAI21_X1 U23099 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n20031), .A(n20030), 
        .ZN(n20033) );
  AOI211_X1 U23100 ( .C1(n20046), .C2(n20033), .A(n20032), .B(n20047), .ZN(
        n20036) );
  OAI21_X1 U23101 ( .B1(n20036), .B2(n20035), .A(n20034), .ZN(n20043) );
  INV_X1 U23102 ( .A(n20051), .ZN(n20044) );
  OAI21_X1 U23103 ( .B1(n20038), .B2(n20037), .A(n20044), .ZN(n20039) );
  AOI21_X1 U23104 ( .B1(n20041), .B2(n20040), .A(n20039), .ZN(n20042) );
  MUX2_X1 U23105 ( .A(n20043), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n20042), 
        .Z(P3_U3296) );
  MUX2_X1 U23106 ( .A(P3_M_IO_N_REG_SCAN_IN), .B(P3_MEMORYFETCH_REG_SCAN_IN), 
        .S(n19996), .Z(P3_U3297) );
  AOI21_X1 U23107 ( .B1(n20048), .B2(n20047), .A(P3_READREQUEST_REG_SCAN_IN), 
        .ZN(n20045) );
  AOI22_X1 U23108 ( .A1(n20051), .A2(n20046), .B1(n20045), .B2(n20044), .ZN(
        P3_U3298) );
  AOI21_X1 U23109 ( .B1(n20048), .B2(n20047), .A(P3_MEMORYFETCH_REG_SCAN_IN), 
        .ZN(n20050) );
  OAI21_X1 U23110 ( .B1(n20051), .B2(n20050), .A(n20049), .ZN(P3_U3299) );
  INV_X1 U23111 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20829) );
  INV_X1 U23112 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n20052) );
  INV_X1 U23113 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20846) );
  NAND2_X1 U23114 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20846), .ZN(n20836) );
  AOI22_X1 U23115 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20836), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n20829), .ZN(n20909) );
  OAI21_X1 U23116 ( .B1(n20829), .B2(n20052), .A(n20828), .ZN(P2_U2815) );
  INV_X1 U23117 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n20054) );
  OAI22_X1 U23118 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20055), .B1(n20054), 
        .B2(n20053), .ZN(P2_U2816) );
  INV_X1 U23119 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20839) );
  INV_X2 U23120 ( .A(n20976), .ZN(n20979) );
  OR2_X1 U23121 ( .A1(n20838), .A2(n20979), .ZN(n20832) );
  AOI21_X1 U23122 ( .B1(n20829), .B2(n20832), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n20056) );
  AOI21_X1 U23123 ( .B1(n20979), .B2(P2_CODEFETCH_REG_SCAN_IN), .A(n20056), 
        .ZN(P2_U2817) );
  OAI21_X1 U23124 ( .B1(n20838), .B2(BS16), .A(n20909), .ZN(n20907) );
  OAI21_X1 U23125 ( .B1(n20909), .B2(n20910), .A(n20907), .ZN(P2_U2818) );
  NOR4_X1 U23126 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20067) );
  NOR4_X1 U23127 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20066) );
  NOR4_X1 U23128 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(P2_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20057) );
  NAND2_X1 U23129 ( .A1(n20058), .A2(n20057), .ZN(n20064) );
  NOR4_X1 U23130 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20062) );
  NOR4_X1 U23131 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20061) );
  NOR4_X1 U23132 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20060) );
  NOR4_X1 U23133 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20059) );
  NAND4_X1 U23134 ( .A1(n20062), .A2(n20061), .A3(n20060), .A4(n20059), .ZN(
        n20063) );
  AOI211_X1 U23135 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20064), .B(n20063), .ZN(n20065) );
  NAND3_X1 U23136 ( .A1(n20067), .A2(n20066), .A3(n20065), .ZN(n20068) );
  NOR2_X1 U23137 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n20068), .ZN(n20070) );
  INV_X1 U23138 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20905) );
  AOI22_X1 U23139 ( .A1(n20070), .A2(n20071), .B1(n20068), .B2(n20905), .ZN(
        P2_U2820) );
  INV_X1 U23140 ( .A(n20068), .ZN(n20076) );
  NOR2_X1 U23141 ( .A1(n20076), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20069)
         );
  OR4_X1 U23142 ( .A1(n20068), .A2(P2_REIP_REG_0__SCAN_IN), .A3(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A4(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20075) );
  OAI21_X1 U23143 ( .B1(n20070), .B2(n20069), .A(n20075), .ZN(P2_U2821) );
  INV_X1 U23144 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20908) );
  NAND2_X1 U23145 ( .A1(n20070), .A2(n20908), .ZN(n20074) );
  OAI21_X1 U23146 ( .B1(n20847), .B2(n20071), .A(n20076), .ZN(n20072) );
  OAI21_X1 U23147 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n20076), .A(n20072), 
        .ZN(n20073) );
  OAI221_X1 U23148 ( .B1(n20074), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n20074), .C2(P2_REIP_REG_0__SCAN_IN), .A(n20073), .ZN(P2_U2822) );
  INV_X1 U23149 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20903) );
  OAI211_X1 U23150 ( .C1(n20076), .C2(n20903), .A(n20075), .B(n20074), .ZN(
        P2_U2823) );
  AOI21_X1 U23151 ( .B1(n20093), .B2(n20095), .A(n20147), .ZN(n20077) );
  XOR2_X1 U23152 ( .A(n20078), .B(n20077), .Z(n20088) );
  AOI21_X1 U23153 ( .B1(n20169), .B2(P2_EBX_REG_17__SCAN_IN), .A(n20167), .ZN(
        n20079) );
  OAI21_X1 U23154 ( .B1(n20877), .B2(n20180), .A(n20079), .ZN(n20082) );
  NOR2_X1 U23155 ( .A1(n20080), .A2(n20165), .ZN(n20081) );
  AOI211_X1 U23156 ( .C1(n20186), .C2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n20082), .B(n20081), .ZN(n20087) );
  OAI22_X1 U23157 ( .A1(n20084), .A2(n20189), .B1(n20083), .B2(n20171), .ZN(
        n20085) );
  INV_X1 U23158 ( .A(n20085), .ZN(n20086) );
  OAI211_X1 U23159 ( .C1(n20177), .C2(n20088), .A(n20087), .B(n20086), .ZN(
        P2_U2838) );
  INV_X1 U23160 ( .A(n20089), .ZN(n20092) );
  AOI21_X1 U23161 ( .B1(n20169), .B2(P2_EBX_REG_16__SCAN_IN), .A(n20167), .ZN(
        n20090) );
  OAI21_X1 U23162 ( .B1(n20875), .B2(n20180), .A(n20090), .ZN(n20091) );
  AOI21_X1 U23163 ( .B1(n20092), .B2(n20187), .A(n20091), .ZN(n20101) );
  INV_X1 U23164 ( .A(n20093), .ZN(n20094) );
  NAND2_X1 U23165 ( .A1(n10322), .A2(n20094), .ZN(n20111) );
  XOR2_X1 U23166 ( .A(n20111), .B(n20095), .Z(n20099) );
  OAI22_X1 U23167 ( .A1(n20097), .A2(n20189), .B1(n20096), .B2(n20171), .ZN(
        n20098) );
  AOI21_X1 U23168 ( .B1(n20099), .B2(n20197), .A(n20098), .ZN(n20100) );
  OAI211_X1 U23169 ( .C1(n20102), .C2(n20145), .A(n20101), .B(n20100), .ZN(
        P2_U2839) );
  NAND2_X1 U23170 ( .A1(n20150), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n20103) );
  OAI211_X1 U23171 ( .C1(n20182), .C2(n20104), .A(n20181), .B(n20103), .ZN(
        n20105) );
  AOI21_X1 U23172 ( .B1(n20106), .B2(n20187), .A(n20105), .ZN(n20117) );
  AOI22_X1 U23173 ( .A1(n20107), .A2(n20112), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n20186), .ZN(n20116) );
  INV_X1 U23174 ( .A(n20108), .ZN(n20109) );
  AOI22_X1 U23175 ( .A1(n20110), .A2(n20129), .B1(n20109), .B2(n20185), .ZN(
        n20115) );
  AOI211_X1 U23176 ( .C1(n20112), .C2(n20121), .A(n20177), .B(n20111), .ZN(
        n20113) );
  INV_X1 U23177 ( .A(n20113), .ZN(n20114) );
  NAND4_X1 U23178 ( .A1(n20117), .A2(n20116), .A3(n20115), .A4(n20114), .ZN(
        P2_U2840) );
  NAND2_X1 U23179 ( .A1(n20118), .A2(n20120), .ZN(n20119) );
  MUX2_X1 U23180 ( .A(n20120), .B(n20119), .S(n10322), .Z(n20122) );
  NAND2_X1 U23181 ( .A1(n20122), .A2(n20121), .ZN(n20133) );
  AOI22_X1 U23182 ( .A1(n20123), .A2(n20187), .B1(n20186), .B2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n20124) );
  OAI21_X1 U23183 ( .B1(n20871), .B2(n20180), .A(n20124), .ZN(n20125) );
  AOI211_X1 U23184 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n20126), .A(n20167), .B(
        n20125), .ZN(n20132) );
  INV_X1 U23185 ( .A(n20127), .ZN(n20130) );
  AOI22_X1 U23186 ( .A1(n20130), .A2(n20129), .B1(n20128), .B2(n20185), .ZN(
        n20131) );
  OAI211_X1 U23187 ( .C1(n20177), .C2(n20133), .A(n20132), .B(n20131), .ZN(
        P2_U2841) );
  OAI22_X1 U23188 ( .A1(n20134), .A2(n20165), .B1(n20863), .B2(n20180), .ZN(
        n20135) );
  AOI211_X1 U23189 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n20169), .A(n20167), .B(
        n20135), .ZN(n20144) );
  NAND2_X1 U23190 ( .A1(n10322), .A2(n20136), .ZN(n20138) );
  XNOR2_X1 U23191 ( .A(n20138), .B(n20137), .ZN(n20142) );
  OAI22_X1 U23192 ( .A1(n20140), .A2(n20189), .B1(n20139), .B2(n20171), .ZN(
        n20141) );
  AOI21_X1 U23193 ( .B1(n20142), .B2(n20197), .A(n20141), .ZN(n20143) );
  OAI211_X1 U23194 ( .C1(n17090), .C2(n20145), .A(n20144), .B(n20143), .ZN(
        P2_U2845) );
  NOR2_X1 U23195 ( .A1(n20147), .A2(n20146), .ZN(n20148) );
  XOR2_X1 U23196 ( .A(n20149), .B(n20148), .Z(n20159) );
  AOI22_X1 U23197 ( .A1(n20151), .A2(n20187), .B1(n20150), .B2(
        P2_REIP_REG_9__SCAN_IN), .ZN(n20152) );
  OAI211_X1 U23198 ( .C1(n20153), .C2(n20182), .A(n20152), .B(n17149), .ZN(
        n20157) );
  OAI22_X1 U23199 ( .A1(n20155), .A2(n20189), .B1(n20154), .B2(n20171), .ZN(
        n20156) );
  AOI211_X1 U23200 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n20186), .A(
        n20157), .B(n20156), .ZN(n20158) );
  OAI21_X1 U23201 ( .B1(n20159), .B2(n20177), .A(n20158), .ZN(P2_U2846) );
  NAND2_X1 U23202 ( .A1(n10322), .A2(n20160), .ZN(n20162) );
  MUX2_X1 U23203 ( .A(n10322), .B(n20162), .S(n20161), .Z(n20164) );
  NAND2_X1 U23204 ( .A1(n20164), .A2(n20163), .ZN(n20178) );
  OAI22_X1 U23205 ( .A1(n20166), .A2(n20165), .B1(n20858), .B2(n20180), .ZN(
        n20168) );
  AOI211_X1 U23206 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n20169), .A(n20168), .B(
        n20167), .ZN(n20170) );
  INV_X1 U23207 ( .A(n20170), .ZN(n20175) );
  OAI22_X1 U23208 ( .A1(n20173), .A2(n20189), .B1(n20172), .B2(n20171), .ZN(
        n20174) );
  AOI211_X1 U23209 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n20186), .A(
        n20175), .B(n20174), .ZN(n20176) );
  OAI21_X1 U23210 ( .B1(n20178), .B2(n20177), .A(n20176), .ZN(P2_U2848) );
  INV_X1 U23211 ( .A(n20179), .ZN(n20208) );
  INV_X1 U23212 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n20853) );
  NOR2_X1 U23213 ( .A1(n20180), .A2(n20853), .ZN(n20184) );
  OAI21_X1 U23214 ( .B1(n20182), .B2(n11105), .A(n20181), .ZN(n20183) );
  AOI211_X1 U23215 ( .C1(n20208), .C2(n20185), .A(n20184), .B(n20183), .ZN(
        n20202) );
  AOI22_X1 U23216 ( .A1(n20188), .A2(n20187), .B1(n20186), .B2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20201) );
  OAI22_X1 U23217 ( .A1(n20209), .A2(n20190), .B1(n20189), .B2(n20203), .ZN(
        n20191) );
  INV_X1 U23218 ( .A(n20191), .ZN(n20200) );
  NAND2_X1 U23219 ( .A1(n20192), .A2(n20195), .ZN(n20194) );
  MUX2_X1 U23220 ( .A(n20195), .B(n20194), .S(n10322), .Z(n20198) );
  NAND3_X1 U23221 ( .A1(n20198), .A2(n20197), .A3(n20196), .ZN(n20199) );
  NAND4_X1 U23222 ( .A1(n20202), .A2(n20201), .A3(n20200), .A4(n20199), .ZN(
        P2_U2851) );
  OAI22_X1 U23223 ( .A1(n20209), .A2(n16752), .B1(n20204), .B2(n20203), .ZN(
        n20205) );
  INV_X1 U23224 ( .A(n20205), .ZN(n20206) );
  OAI21_X1 U23225 ( .B1(n20207), .B2(n11105), .A(n20206), .ZN(P2_U2883) );
  AOI22_X1 U23226 ( .A1(n20208), .A2(n12194), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n20226), .ZN(n20213) );
  XNOR2_X1 U23227 ( .A(n20210), .B(n20209), .ZN(n20211) );
  NAND2_X1 U23228 ( .A1(n20211), .A2(n20227), .ZN(n20212) );
  OAI211_X1 U23229 ( .C1(n20305), .C2(n20232), .A(n20213), .B(n20212), .ZN(
        P2_U2915) );
  AOI22_X1 U23230 ( .A1(n12194), .A2(n20917), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n20226), .ZN(n20219) );
  OAI21_X1 U23231 ( .B1(n20216), .B2(n20215), .A(n20214), .ZN(n20217) );
  NAND2_X1 U23232 ( .A1(n20217), .A2(n20227), .ZN(n20218) );
  OAI211_X1 U23233 ( .C1(n20302), .C2(n20232), .A(n20219), .B(n20218), .ZN(
        P2_U2916) );
  AOI22_X1 U23234 ( .A1(n12194), .A2(n20934), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n20226), .ZN(n20224) );
  OAI21_X1 U23235 ( .B1(n20221), .B2(n20228), .A(n20220), .ZN(n20222) );
  NAND2_X1 U23236 ( .A1(n20222), .A2(n20227), .ZN(n20223) );
  OAI211_X1 U23237 ( .C1(n20225), .C2(n20232), .A(n20224), .B(n20223), .ZN(
        P2_U2918) );
  AOI22_X1 U23238 ( .A1(n12194), .A2(n20229), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n20226), .ZN(n20231) );
  OAI211_X1 U23239 ( .C1(n20944), .C2(n20229), .A(n20228), .B(n20227), .ZN(
        n20230) );
  OAI211_X1 U23240 ( .C1(n20233), .C2(n20232), .A(n20231), .B(n20230), .ZN(
        P2_U2919) );
  NOR2_X1 U23241 ( .A1(n20271), .A2(n20234), .ZN(P2_U2920) );
  INV_X1 U23242 ( .A(n20235), .ZN(n20236) );
  AOI22_X1 U23243 ( .A1(n20236), .A2(P2_EAX_REG_28__SCAN_IN), .B1(
        P2_UWORD_REG_12__SCAN_IN), .B2(n20273), .ZN(n20237) );
  OAI21_X1 U23244 ( .B1(n20238), .B2(n20271), .A(n20237), .ZN(P2_U2923) );
  AOI22_X1 U23245 ( .A1(n20273), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n20240), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n20239) );
  OAI21_X1 U23246 ( .B1(n20276), .B2(n13235), .A(n20239), .ZN(P2_U2936) );
  AOI22_X1 U23247 ( .A1(n20273), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n20240), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n20241) );
  OAI21_X1 U23248 ( .B1(n20276), .B2(n20242), .A(n20241), .ZN(P2_U2937) );
  INV_X1 U23249 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n20245) );
  OAI222_X1 U23250 ( .A1(n20245), .A2(n20962), .B1(n20244), .B2(n20276), .C1(
        n20243), .C2(n20271), .ZN(P2_U2938) );
  INV_X1 U23251 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n20247) );
  AOI22_X1 U23252 ( .A1(n20273), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n20272), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n20246) );
  OAI21_X1 U23253 ( .B1(n20276), .B2(n20247), .A(n20246), .ZN(P2_U2939) );
  AOI22_X1 U23254 ( .A1(n20273), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n20272), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n20248) );
  OAI21_X1 U23255 ( .B1(n20276), .B2(n20249), .A(n20248), .ZN(P2_U2940) );
  AOI22_X1 U23256 ( .A1(n20273), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n20272), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n20250) );
  OAI21_X1 U23257 ( .B1(n20276), .B2(n20251), .A(n20250), .ZN(P2_U2941) );
  AOI22_X1 U23258 ( .A1(n20273), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n20272), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n20252) );
  OAI21_X1 U23259 ( .B1(n20276), .B2(n20253), .A(n20252), .ZN(P2_U2942) );
  AOI22_X1 U23260 ( .A1(n20273), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n20272), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n20254) );
  OAI21_X1 U23261 ( .B1(n20276), .B2(n20255), .A(n20254), .ZN(P2_U2943) );
  AOI22_X1 U23262 ( .A1(n20273), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n20272), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n20256) );
  OAI21_X1 U23263 ( .B1(n20276), .B2(n20257), .A(n20256), .ZN(P2_U2944) );
  AOI22_X1 U23264 ( .A1(n20273), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n20272), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n20258) );
  OAI21_X1 U23265 ( .B1(n20276), .B2(n20259), .A(n20258), .ZN(P2_U2945) );
  AOI22_X1 U23266 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n20260), .B1(n20272), .B2(
        P2_DATAO_REG_5__SCAN_IN), .ZN(n20261) );
  OAI21_X1 U23267 ( .B1(n13997), .B2(n20962), .A(n20261), .ZN(P2_U2946) );
  INV_X1 U23268 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n20263) );
  AOI22_X1 U23269 ( .A1(n20273), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n20272), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n20262) );
  OAI21_X1 U23270 ( .B1(n20276), .B2(n20263), .A(n20262), .ZN(P2_U2947) );
  INV_X1 U23271 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n20265) );
  AOI22_X1 U23272 ( .A1(n20273), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n20272), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n20264) );
  OAI21_X1 U23273 ( .B1(n20276), .B2(n20265), .A(n20264), .ZN(P2_U2948) );
  INV_X1 U23274 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n20267) );
  AOI22_X1 U23275 ( .A1(n20273), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n20272), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n20266) );
  OAI21_X1 U23276 ( .B1(n20276), .B2(n20267), .A(n20266), .ZN(P2_U2949) );
  INV_X1 U23277 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n20269) );
  OAI222_X1 U23278 ( .A1(n20271), .A2(n20270), .B1(n20269), .B2(n20276), .C1(
        n20268), .C2(n20962), .ZN(P2_U2950) );
  INV_X1 U23279 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n20275) );
  AOI22_X1 U23280 ( .A1(n20273), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n20272), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n20274) );
  OAI21_X1 U23281 ( .B1(n20276), .B2(n20275), .A(n20274), .ZN(P2_U2951) );
  AOI22_X1 U23282 ( .A1(P2_UWORD_REG_12__SCAN_IN), .A2(n20277), .B1(n20281), 
        .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n20280) );
  NAND2_X1 U23283 ( .A1(n20279), .A2(n20278), .ZN(n20283) );
  NAND2_X1 U23284 ( .A1(n20280), .A2(n20283), .ZN(P2_U2964) );
  AOI22_X1 U23285 ( .A1(P2_LWORD_REG_12__SCAN_IN), .A2(n20282), .B1(n20281), 
        .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n20284) );
  NAND2_X1 U23286 ( .A1(n20284), .A2(n20283), .ZN(P2_U2979) );
  NAND2_X1 U23287 ( .A1(n20920), .A2(n20927), .ZN(n20388) );
  OR2_X1 U23288 ( .A1(n20388), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20330) );
  NOR2_X1 U23289 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20330), .ZN(
        n20318) );
  AOI22_X1 U23290 ( .A1(n20757), .A2(n20819), .B1(n20691), .B2(n20318), .ZN(
        n20295) );
  AOI21_X1 U23291 ( .B1(n20285), .B2(n20355), .A(n20910), .ZN(n20286) );
  NOR2_X1 U23292 ( .A1(n20286), .A2(n20563), .ZN(n20289) );
  OAI21_X1 U23293 ( .B1(n20291), .B2(n20939), .A(n17491), .ZN(n20287) );
  AOI21_X1 U23294 ( .B1(n20289), .B2(n20814), .A(n20287), .ZN(n20288) );
  OAI21_X1 U23295 ( .B1(n20288), .B2(n20318), .A(n20697), .ZN(n20321) );
  OAI21_X1 U23296 ( .B1(n20290), .B2(n20318), .A(n20289), .ZN(n20293) );
  OAI21_X1 U23297 ( .B1(n20291), .B2(n20318), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20292) );
  AOI22_X1 U23298 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20321), .B1(
        n20692), .B2(n20320), .ZN(n20294) );
  OAI211_X1 U23299 ( .C1(n20663), .C2(n20355), .A(n20295), .B(n20294), .ZN(
        P2_U3048) );
  AOI22_X1 U23300 ( .A1(n20729), .A2(n20819), .B1(n20727), .B2(n20318), .ZN(
        n20297) );
  AOI22_X1 U23301 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20321), .B1(
        n20730), .B2(n20320), .ZN(n20296) );
  OAI211_X1 U23302 ( .C1(n20666), .C2(n20355), .A(n20297), .B(n20296), .ZN(
        P2_U3049) );
  AOI22_X1 U23303 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20315), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20314), .ZN(n20669) );
  AOI22_X1 U23304 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n20314), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n20315), .ZN(n20707) );
  NOR2_X2 U23305 ( .A1(n20317), .A2(n20298), .ZN(n20762) );
  AOI22_X1 U23306 ( .A1(n20767), .A2(n20819), .B1(n20762), .B2(n20318), .ZN(
        n20301) );
  NOR2_X2 U23307 ( .A1(n20510), .A2(n20299), .ZN(n20761) );
  AOI22_X1 U23308 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20321), .B1(
        n20761), .B2(n20320), .ZN(n20300) );
  OAI211_X1 U23309 ( .C1(n20669), .C2(n20355), .A(n20301), .B(n20300), .ZN(
        P2_U3050) );
  AOI22_X1 U23310 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20315), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20314), .ZN(n20672) );
  AOI22_X1 U23311 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20315), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n20314), .ZN(n20710) );
  AOI22_X1 U23312 ( .A1(n20776), .A2(n20819), .B1(n20772), .B2(n20318), .ZN(
        n20304) );
  NOR2_X2 U23313 ( .A1(n20302), .A2(n20510), .ZN(n20771) );
  AOI22_X1 U23314 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20321), .B1(
        n20771), .B2(n20320), .ZN(n20303) );
  OAI211_X1 U23315 ( .C1(n20672), .C2(n20355), .A(n20304), .B(n20303), .ZN(
        P2_U3051) );
  AOI22_X1 U23316 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20315), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20314), .ZN(n20675) );
  AOI22_X1 U23317 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n20314), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n20315), .ZN(n20713) );
  NOR2_X2 U23318 ( .A1(n20317), .A2(n9921), .ZN(n20782) );
  AOI22_X1 U23319 ( .A1(n20787), .A2(n20819), .B1(n20782), .B2(n20318), .ZN(
        n20307) );
  NOR2_X2 U23320 ( .A1(n20510), .A2(n20305), .ZN(n20781) );
  AOI22_X1 U23321 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20321), .B1(
        n20781), .B2(n20320), .ZN(n20306) );
  OAI211_X1 U23322 ( .C1(n20675), .C2(n20355), .A(n20307), .B(n20306), .ZN(
        P2_U3052) );
  AOI22_X1 U23323 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20315), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n20314), .ZN(n20678) );
  AOI22_X1 U23324 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n20314), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n20315), .ZN(n20716) );
  INV_X1 U23325 ( .A(n20716), .ZN(n20796) );
  NOR2_X2 U23326 ( .A1(n20317), .A2(n11473), .ZN(n20792) );
  AOI22_X1 U23327 ( .A1(n20796), .A2(n20819), .B1(n20792), .B2(n20318), .ZN(
        n20310) );
  NOR2_X2 U23328 ( .A1(n20308), .A2(n20510), .ZN(n20791) );
  AOI22_X1 U23329 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20321), .B1(
        n20791), .B2(n20320), .ZN(n20309) );
  OAI211_X1 U23330 ( .C1(n20678), .C2(n20355), .A(n20310), .B(n20309), .ZN(
        P2_U3053) );
  AOI22_X1 U23331 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20315), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n20314), .ZN(n20681) );
  AOI22_X1 U23332 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n20314), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n20315), .ZN(n20719) );
  INV_X1 U23333 ( .A(n20719), .ZN(n20806) );
  NOR2_X2 U23334 ( .A1(n20317), .A2(n13913), .ZN(n20802) );
  AOI22_X1 U23335 ( .A1(n20806), .A2(n20819), .B1(n20802), .B2(n20318), .ZN(
        n20313) );
  NOR2_X2 U23336 ( .A1(n20510), .A2(n20311), .ZN(n20801) );
  AOI22_X1 U23337 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20321), .B1(
        n20801), .B2(n20320), .ZN(n20312) );
  OAI211_X1 U23338 ( .C1(n20681), .C2(n20355), .A(n20313), .B(n20312), .ZN(
        P2_U3054) );
  AOI22_X1 U23339 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20315), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n20314), .ZN(n20688) );
  AOI22_X1 U23340 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20315), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n20314), .ZN(n20726) );
  INV_X1 U23341 ( .A(n20726), .ZN(n20820) );
  NOR2_X2 U23342 ( .A1(n20317), .A2(n20316), .ZN(n20812) );
  AOI22_X1 U23343 ( .A1(n20820), .A2(n20819), .B1(n20812), .B2(n20318), .ZN(
        n20323) );
  NOR2_X2 U23344 ( .A1(n20319), .A2(n20510), .ZN(n20811) );
  AOI22_X1 U23345 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20321), .B1(
        n20811), .B2(n20320), .ZN(n20322) );
  OAI211_X1 U23346 ( .C1(n20688), .C2(n20355), .A(n20323), .B(n20322), .ZN(
        P2_U3055) );
  NAND2_X1 U23347 ( .A1(n20324), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20507) );
  OAI21_X1 U23348 ( .B1(n20507), .B2(n20562), .A(n20330), .ZN(n20328) );
  OAI21_X1 U23349 ( .B1(n10909), .B2(n20939), .A(n17491), .ZN(n20326) );
  NAND2_X1 U23350 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20938), .ZN(
        n20450) );
  NOR2_X1 U23351 ( .A1(n20450), .A2(n20388), .ZN(n20350) );
  INV_X1 U23352 ( .A(n20350), .ZN(n20325) );
  AOI21_X1 U23353 ( .B1(n20326), .B2(n20325), .A(n20510), .ZN(n20327) );
  OAI21_X1 U23354 ( .B1(n10909), .B2(n20350), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20329) );
  OAI21_X1 U23355 ( .B1(n20330), .B2(n20563), .A(n20329), .ZN(n20351) );
  AOI22_X1 U23356 ( .A1(n20351), .A2(n20692), .B1(n20691), .B2(n20350), .ZN(
        n20332) );
  AOI22_X1 U23357 ( .A1(n20346), .A2(n20757), .B1(n20383), .B2(n20756), .ZN(
        n20331) );
  OAI211_X1 U23358 ( .C1(n20339), .C2(n20333), .A(n20332), .B(n20331), .ZN(
        P2_U3056) );
  AOI22_X1 U23359 ( .A1(n20351), .A2(n20730), .B1(n20727), .B2(n20350), .ZN(
        n20335) );
  AOI22_X1 U23360 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20352), .B1(
        n20383), .B2(n20728), .ZN(n20334) );
  OAI211_X1 U23361 ( .C1(n20704), .C2(n20355), .A(n20335), .B(n20334), .ZN(
        P2_U3057) );
  AOI22_X1 U23362 ( .A1(n20351), .A2(n20761), .B1(n20762), .B2(n20350), .ZN(
        n20337) );
  AOI22_X1 U23363 ( .A1(n20346), .A2(n20767), .B1(n20383), .B2(n20766), .ZN(
        n20336) );
  OAI211_X1 U23364 ( .C1(n20339), .C2(n20338), .A(n20337), .B(n20336), .ZN(
        P2_U3058) );
  AOI22_X1 U23365 ( .A1(n20351), .A2(n20771), .B1(n20772), .B2(n20350), .ZN(
        n20341) );
  AOI22_X1 U23366 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20352), .B1(
        n20383), .B2(n20777), .ZN(n20340) );
  OAI211_X1 U23367 ( .C1(n20710), .C2(n20355), .A(n20341), .B(n20340), .ZN(
        P2_U3059) );
  AOI22_X1 U23368 ( .A1(n20351), .A2(n20781), .B1(n20782), .B2(n20350), .ZN(
        n20343) );
  INV_X1 U23369 ( .A(n20675), .ZN(n20786) );
  AOI22_X1 U23370 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20352), .B1(
        n20383), .B2(n20786), .ZN(n20342) );
  OAI211_X1 U23371 ( .C1(n20713), .C2(n20355), .A(n20343), .B(n20342), .ZN(
        P2_U3060) );
  AOI22_X1 U23372 ( .A1(n20351), .A2(n20791), .B1(n20792), .B2(n20350), .ZN(
        n20345) );
  AOI22_X1 U23373 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20352), .B1(
        n20383), .B2(n20797), .ZN(n20344) );
  OAI211_X1 U23374 ( .C1(n20716), .C2(n20355), .A(n20345), .B(n20344), .ZN(
        P2_U3061) );
  INV_X1 U23375 ( .A(n20383), .ZN(n20349) );
  AOI22_X1 U23376 ( .A1(n20351), .A2(n20801), .B1(n20802), .B2(n20350), .ZN(
        n20348) );
  AOI22_X1 U23377 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20352), .B1(
        n20346), .B2(n20806), .ZN(n20347) );
  OAI211_X1 U23378 ( .C1(n20681), .C2(n20349), .A(n20348), .B(n20347), .ZN(
        P2_U3062) );
  AOI22_X1 U23379 ( .A1(n20351), .A2(n20811), .B1(n20812), .B2(n20350), .ZN(
        n20354) );
  AOI22_X1 U23380 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20352), .B1(
        n20383), .B2(n20818), .ZN(n20353) );
  OAI211_X1 U23381 ( .C1(n20726), .C2(n20355), .A(n20354), .B(n20353), .ZN(
        P2_U3063) );
  INV_X1 U23382 ( .A(n20424), .ZN(n20356) );
  NOR2_X1 U23383 ( .A1(n20357), .A2(n20388), .ZN(n20381) );
  OAI21_X1 U23384 ( .B1(n20361), .B2(n20381), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20360) );
  INV_X1 U23385 ( .A(n20388), .ZN(n20358) );
  NAND2_X1 U23386 ( .A1(n20359), .A2(n20358), .ZN(n20363) );
  NAND2_X1 U23387 ( .A1(n20360), .A2(n20363), .ZN(n20382) );
  AOI22_X1 U23388 ( .A1(n20382), .A2(n20692), .B1(n20691), .B2(n20381), .ZN(
        n20368) );
  INV_X1 U23389 ( .A(n20361), .ZN(n20362) );
  AOI21_X1 U23390 ( .B1(n20362), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20366) );
  OAI21_X1 U23391 ( .B1(n20405), .B2(n20383), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20364) );
  NAND3_X1 U23392 ( .A1(n20364), .A2(n20958), .A3(n20363), .ZN(n20365) );
  OAI211_X1 U23393 ( .C1(n20381), .C2(n20366), .A(n20365), .B(n20697), .ZN(
        n20384) );
  AOI22_X1 U23394 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20384), .B1(
        n20383), .B2(n20757), .ZN(n20367) );
  OAI211_X1 U23395 ( .C1(n20663), .C2(n20417), .A(n20368), .B(n20367), .ZN(
        P2_U3064) );
  AOI22_X1 U23396 ( .A1(n20382), .A2(n20730), .B1(n20727), .B2(n20381), .ZN(
        n20370) );
  AOI22_X1 U23397 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20384), .B1(
        n20383), .B2(n20729), .ZN(n20369) );
  OAI211_X1 U23398 ( .C1(n20666), .C2(n20417), .A(n20370), .B(n20369), .ZN(
        P2_U3065) );
  AOI22_X1 U23399 ( .A1(n20382), .A2(n20761), .B1(n20762), .B2(n20381), .ZN(
        n20372) );
  AOI22_X1 U23400 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20384), .B1(
        n20383), .B2(n20767), .ZN(n20371) );
  OAI211_X1 U23401 ( .C1(n20669), .C2(n20417), .A(n20372), .B(n20371), .ZN(
        P2_U3066) );
  AOI22_X1 U23402 ( .A1(n20382), .A2(n20771), .B1(n20772), .B2(n20381), .ZN(
        n20374) );
  AOI22_X1 U23403 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20384), .B1(
        n20383), .B2(n20776), .ZN(n20373) );
  OAI211_X1 U23404 ( .C1(n20672), .C2(n20417), .A(n20374), .B(n20373), .ZN(
        P2_U3067) );
  AOI22_X1 U23405 ( .A1(n20382), .A2(n20781), .B1(n20782), .B2(n20381), .ZN(
        n20376) );
  AOI22_X1 U23406 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20384), .B1(
        n20383), .B2(n20787), .ZN(n20375) );
  OAI211_X1 U23407 ( .C1(n20675), .C2(n20417), .A(n20376), .B(n20375), .ZN(
        P2_U3068) );
  AOI22_X1 U23408 ( .A1(n20382), .A2(n20791), .B1(n20792), .B2(n20381), .ZN(
        n20378) );
  AOI22_X1 U23409 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20384), .B1(
        n20383), .B2(n20796), .ZN(n20377) );
  OAI211_X1 U23410 ( .C1(n20678), .C2(n20417), .A(n20378), .B(n20377), .ZN(
        P2_U3069) );
  AOI22_X1 U23411 ( .A1(n20382), .A2(n20801), .B1(n20802), .B2(n20381), .ZN(
        n20380) );
  AOI22_X1 U23412 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20384), .B1(
        n20383), .B2(n20806), .ZN(n20379) );
  OAI211_X1 U23413 ( .C1(n20681), .C2(n20417), .A(n20380), .B(n20379), .ZN(
        P2_U3070) );
  AOI22_X1 U23414 ( .A1(n20382), .A2(n20811), .B1(n20812), .B2(n20381), .ZN(
        n20386) );
  AOI22_X1 U23415 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20384), .B1(
        n20383), .B2(n20820), .ZN(n20385) );
  OAI211_X1 U23416 ( .C1(n20688), .C2(n20417), .A(n20386), .B(n20385), .ZN(
        P2_U3071) );
  NOR2_X1 U23417 ( .A1(n20387), .A2(n20388), .ZN(n20412) );
  AOI22_X1 U23418 ( .A1(n20756), .A2(n20446), .B1(n20691), .B2(n20412), .ZN(
        n20398) );
  OAI21_X1 U23419 ( .B1(n20507), .B2(n20629), .A(n20958), .ZN(n20396) );
  NOR2_X1 U23420 ( .A1(n20938), .A2(n20388), .ZN(n20392) );
  INV_X1 U23421 ( .A(n20393), .ZN(n20390) );
  INV_X1 U23422 ( .A(n20412), .ZN(n20389) );
  OAI211_X1 U23423 ( .C1(n20390), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20563), 
        .B(n20389), .ZN(n20391) );
  OAI211_X1 U23424 ( .C1(n20396), .C2(n20392), .A(n20697), .B(n20391), .ZN(
        n20414) );
  INV_X1 U23425 ( .A(n20392), .ZN(n20395) );
  OAI21_X1 U23426 ( .B1(n20393), .B2(n20412), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20394) );
  AOI22_X1 U23427 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20414), .B1(
        n20692), .B2(n20413), .ZN(n20397) );
  OAI211_X1 U23428 ( .C1(n20701), .C2(n20417), .A(n20398), .B(n20397), .ZN(
        P2_U3072) );
  AOI22_X1 U23429 ( .A1(n20728), .A2(n20446), .B1(n20727), .B2(n20412), .ZN(
        n20400) );
  AOI22_X1 U23430 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20414), .B1(
        n20730), .B2(n20413), .ZN(n20399) );
  OAI211_X1 U23431 ( .C1(n20704), .C2(n20417), .A(n20400), .B(n20399), .ZN(
        P2_U3073) );
  AOI22_X1 U23432 ( .A1(n20767), .A2(n20405), .B1(n20412), .B2(n20762), .ZN(
        n20402) );
  AOI22_X1 U23433 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20414), .B1(
        n20761), .B2(n20413), .ZN(n20401) );
  OAI211_X1 U23434 ( .C1(n20669), .C2(n20443), .A(n20402), .B(n20401), .ZN(
        P2_U3074) );
  AOI22_X1 U23435 ( .A1(n20777), .A2(n20446), .B1(n20412), .B2(n20772), .ZN(
        n20404) );
  AOI22_X1 U23436 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20414), .B1(
        n20771), .B2(n20413), .ZN(n20403) );
  OAI211_X1 U23437 ( .C1(n20710), .C2(n20417), .A(n20404), .B(n20403), .ZN(
        P2_U3075) );
  AOI22_X1 U23438 ( .A1(n20787), .A2(n20405), .B1(n20412), .B2(n20782), .ZN(
        n20407) );
  AOI22_X1 U23439 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20414), .B1(
        n20781), .B2(n20413), .ZN(n20406) );
  OAI211_X1 U23440 ( .C1(n20675), .C2(n20443), .A(n20407), .B(n20406), .ZN(
        P2_U3076) );
  AOI22_X1 U23441 ( .A1(n20797), .A2(n20446), .B1(n20412), .B2(n20792), .ZN(
        n20409) );
  AOI22_X1 U23442 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20414), .B1(
        n20791), .B2(n20413), .ZN(n20408) );
  OAI211_X1 U23443 ( .C1(n20716), .C2(n20417), .A(n20409), .B(n20408), .ZN(
        P2_U3077) );
  AOI22_X1 U23444 ( .A1(n20807), .A2(n20446), .B1(n20412), .B2(n20802), .ZN(
        n20411) );
  AOI22_X1 U23445 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20414), .B1(
        n20801), .B2(n20413), .ZN(n20410) );
  OAI211_X1 U23446 ( .C1(n20719), .C2(n20417), .A(n20411), .B(n20410), .ZN(
        P2_U3078) );
  AOI22_X1 U23447 ( .A1(n20818), .A2(n20446), .B1(n20412), .B2(n20812), .ZN(
        n20416) );
  AOI22_X1 U23448 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20414), .B1(
        n20811), .B2(n20413), .ZN(n20415) );
  OAI211_X1 U23449 ( .C1(n20726), .C2(n20417), .A(n20416), .B(n20415), .ZN(
        P2_U3079) );
  INV_X1 U23450 ( .A(n20418), .ZN(n20421) );
  INV_X1 U23451 ( .A(n20419), .ZN(n20420) );
  NAND2_X1 U23452 ( .A1(n20421), .A2(n20420), .ZN(n20658) );
  NOR2_X1 U23453 ( .A1(n20658), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20428) );
  INV_X1 U23454 ( .A(n20428), .ZN(n20423) );
  NOR3_X2 U23455 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n20451), .ZN(n20444) );
  OAI21_X1 U23456 ( .B1(n10945), .B2(n20444), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20422) );
  AOI22_X1 U23457 ( .A1(n20445), .A2(n20692), .B1(n20691), .B2(n20444), .ZN(
        n20430) );
  AOI21_X1 U23458 ( .B1(n20443), .B2(n20481), .A(n20910), .ZN(n20427) );
  INV_X1 U23459 ( .A(n20444), .ZN(n20425) );
  OAI211_X1 U23460 ( .C1(n10900), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20563), 
        .B(n20425), .ZN(n20426) );
  OAI211_X1 U23461 ( .C1(n20428), .C2(n20427), .A(n20426), .B(n20697), .ZN(
        n20447) );
  AOI22_X1 U23462 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20447), .B1(
        n20470), .B2(n20756), .ZN(n20429) );
  OAI211_X1 U23463 ( .C1(n20701), .C2(n20443), .A(n20430), .B(n20429), .ZN(
        P2_U3080) );
  AOI22_X1 U23464 ( .A1(n20445), .A2(n20730), .B1(n20727), .B2(n20444), .ZN(
        n20432) );
  AOI22_X1 U23465 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20447), .B1(
        n20470), .B2(n20728), .ZN(n20431) );
  OAI211_X1 U23466 ( .C1(n20704), .C2(n20443), .A(n20432), .B(n20431), .ZN(
        P2_U3081) );
  AOI22_X1 U23467 ( .A1(n20445), .A2(n20761), .B1(n20762), .B2(n20444), .ZN(
        n20434) );
  AOI22_X1 U23468 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20447), .B1(
        n20470), .B2(n20766), .ZN(n20433) );
  OAI211_X1 U23469 ( .C1(n20707), .C2(n20443), .A(n20434), .B(n20433), .ZN(
        P2_U3082) );
  AOI22_X1 U23470 ( .A1(n20445), .A2(n20771), .B1(n20772), .B2(n20444), .ZN(
        n20436) );
  AOI22_X1 U23471 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20447), .B1(
        n20446), .B2(n20776), .ZN(n20435) );
  OAI211_X1 U23472 ( .C1(n20672), .C2(n20481), .A(n20436), .B(n20435), .ZN(
        P2_U3083) );
  AOI22_X1 U23473 ( .A1(n20445), .A2(n20781), .B1(n20782), .B2(n20444), .ZN(
        n20438) );
  AOI22_X1 U23474 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20447), .B1(
        n20446), .B2(n20787), .ZN(n20437) );
  OAI211_X1 U23475 ( .C1(n20675), .C2(n20481), .A(n20438), .B(n20437), .ZN(
        P2_U3084) );
  AOI22_X1 U23476 ( .A1(n20445), .A2(n20791), .B1(n20792), .B2(n20444), .ZN(
        n20440) );
  AOI22_X1 U23477 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20447), .B1(
        n20470), .B2(n20797), .ZN(n20439) );
  OAI211_X1 U23478 ( .C1(n20716), .C2(n20443), .A(n20440), .B(n20439), .ZN(
        P2_U3085) );
  AOI22_X1 U23479 ( .A1(n20445), .A2(n20801), .B1(n20802), .B2(n20444), .ZN(
        n20442) );
  AOI22_X1 U23480 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20447), .B1(
        n20470), .B2(n20807), .ZN(n20441) );
  OAI211_X1 U23481 ( .C1(n20719), .C2(n20443), .A(n20442), .B(n20441), .ZN(
        P2_U3086) );
  AOI22_X1 U23482 ( .A1(n20445), .A2(n20811), .B1(n20812), .B2(n20444), .ZN(
        n20449) );
  AOI22_X1 U23483 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20447), .B1(
        n20446), .B2(n20820), .ZN(n20448) );
  OAI211_X1 U23484 ( .C1(n20688), .C2(n20481), .A(n20449), .B(n20448), .ZN(
        P2_U3087) );
  NOR2_X1 U23485 ( .A1(n20450), .A2(n20451), .ZN(n20475) );
  AOI22_X1 U23486 ( .A1(n20756), .A2(n20476), .B1(n20691), .B2(n20475), .ZN(
        n20461) );
  OAI21_X1 U23487 ( .B1(n20507), .B2(n20695), .A(n20958), .ZN(n20459) );
  NOR2_X1 U23488 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20451), .ZN(
        n20455) );
  INV_X1 U23489 ( .A(n20456), .ZN(n20453) );
  INV_X1 U23490 ( .A(n20475), .ZN(n20452) );
  OAI211_X1 U23491 ( .C1(n20453), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20563), 
        .B(n20452), .ZN(n20454) );
  OAI211_X1 U23492 ( .C1(n20459), .C2(n20455), .A(n20697), .B(n20454), .ZN(
        n20478) );
  INV_X1 U23493 ( .A(n20455), .ZN(n20458) );
  OAI21_X1 U23494 ( .B1(n20456), .B2(n20475), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20457) );
  AOI22_X1 U23495 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20478), .B1(
        n20692), .B2(n20477), .ZN(n20460) );
  OAI211_X1 U23496 ( .C1(n20701), .C2(n20481), .A(n20461), .B(n20460), .ZN(
        P2_U3088) );
  AOI22_X1 U23497 ( .A1(n20728), .A2(n20476), .B1(n20727), .B2(n20475), .ZN(
        n20463) );
  AOI22_X1 U23498 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20478), .B1(
        n20730), .B2(n20477), .ZN(n20462) );
  OAI211_X1 U23499 ( .C1(n20704), .C2(n20481), .A(n20463), .B(n20462), .ZN(
        P2_U3089) );
  AOI22_X1 U23500 ( .A1(n20767), .A2(n20470), .B1(n20762), .B2(n20475), .ZN(
        n20465) );
  AOI22_X1 U23501 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20478), .B1(
        n20761), .B2(n20477), .ZN(n20464) );
  OAI211_X1 U23502 ( .C1(n20669), .C2(n17480), .A(n20465), .B(n20464), .ZN(
        P2_U3090) );
  AOI22_X1 U23503 ( .A1(n20776), .A2(n20470), .B1(n20772), .B2(n20475), .ZN(
        n20467) );
  AOI22_X1 U23504 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20478), .B1(
        n20771), .B2(n20477), .ZN(n20466) );
  OAI211_X1 U23505 ( .C1(n20672), .C2(n17480), .A(n20467), .B(n20466), .ZN(
        P2_U3091) );
  AOI22_X1 U23506 ( .A1(n20786), .A2(n20476), .B1(n20475), .B2(n20782), .ZN(
        n20469) );
  AOI22_X1 U23507 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20478), .B1(
        n20781), .B2(n20477), .ZN(n20468) );
  OAI211_X1 U23508 ( .C1(n20713), .C2(n20481), .A(n20469), .B(n20468), .ZN(
        P2_U3092) );
  AOI22_X1 U23509 ( .A1(n20796), .A2(n20470), .B1(n20792), .B2(n20475), .ZN(
        n20472) );
  AOI22_X1 U23510 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20478), .B1(
        n20791), .B2(n20477), .ZN(n20471) );
  OAI211_X1 U23511 ( .C1(n20678), .C2(n17480), .A(n20472), .B(n20471), .ZN(
        P2_U3093) );
  AOI22_X1 U23512 ( .A1(n20807), .A2(n20476), .B1(n20475), .B2(n20802), .ZN(
        n20474) );
  AOI22_X1 U23513 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20478), .B1(
        n20801), .B2(n20477), .ZN(n20473) );
  OAI211_X1 U23514 ( .C1(n20719), .C2(n20481), .A(n20474), .B(n20473), .ZN(
        P2_U3094) );
  AOI22_X1 U23515 ( .A1(n20818), .A2(n20476), .B1(n20475), .B2(n20812), .ZN(
        n20480) );
  AOI22_X1 U23516 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20478), .B1(
        n20811), .B2(n20477), .ZN(n20479) );
  OAI211_X1 U23517 ( .C1(n20726), .C2(n20481), .A(n20480), .B(n20479), .ZN(
        P2_U3095) );
  AOI22_X1 U23518 ( .A1(n20496), .A2(n20730), .B1(n20495), .B2(n20727), .ZN(
        n20484) );
  AOI22_X1 U23519 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20497), .B1(
        n20529), .B2(n20728), .ZN(n20483) );
  OAI211_X1 U23520 ( .C1(n20704), .C2(n17480), .A(n20484), .B(n20483), .ZN(
        P2_U3097) );
  AOI22_X1 U23521 ( .A1(n20496), .A2(n20761), .B1(n20495), .B2(n20762), .ZN(
        n20486) );
  AOI22_X1 U23522 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20497), .B1(
        n20529), .B2(n20766), .ZN(n20485) );
  OAI211_X1 U23523 ( .C1(n20707), .C2(n17480), .A(n20486), .B(n20485), .ZN(
        P2_U3098) );
  AOI22_X1 U23524 ( .A1(n20496), .A2(n20771), .B1(n20495), .B2(n20772), .ZN(
        n20488) );
  AOI22_X1 U23525 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20497), .B1(
        n20529), .B2(n20777), .ZN(n20487) );
  OAI211_X1 U23526 ( .C1(n20710), .C2(n17480), .A(n20488), .B(n20487), .ZN(
        P2_U3099) );
  AOI22_X1 U23527 ( .A1(n20496), .A2(n20781), .B1(n20495), .B2(n20782), .ZN(
        n20490) );
  AOI22_X1 U23528 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20497), .B1(
        n20529), .B2(n20786), .ZN(n20489) );
  OAI211_X1 U23529 ( .C1(n20713), .C2(n17480), .A(n20490), .B(n20489), .ZN(
        P2_U3100) );
  AOI22_X1 U23530 ( .A1(n20496), .A2(n20791), .B1(n20495), .B2(n20792), .ZN(
        n20492) );
  AOI22_X1 U23531 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20497), .B1(
        n20529), .B2(n20797), .ZN(n20491) );
  OAI211_X1 U23532 ( .C1(n20716), .C2(n17480), .A(n20492), .B(n20491), .ZN(
        P2_U3101) );
  AOI22_X1 U23533 ( .A1(n20496), .A2(n20801), .B1(n20495), .B2(n20802), .ZN(
        n20494) );
  AOI22_X1 U23534 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20497), .B1(
        n20529), .B2(n20807), .ZN(n20493) );
  OAI211_X1 U23535 ( .C1(n20719), .C2(n17480), .A(n20494), .B(n20493), .ZN(
        P2_U3102) );
  AOI22_X1 U23536 ( .A1(n20496), .A2(n20811), .B1(n20495), .B2(n20812), .ZN(
        n20499) );
  AOI22_X1 U23537 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20497), .B1(
        n20529), .B2(n20818), .ZN(n20498) );
  OAI211_X1 U23538 ( .C1(n20726), .C2(n17480), .A(n20499), .B(n20498), .ZN(
        P2_U3103) );
  INV_X1 U23539 ( .A(n20500), .ZN(n20502) );
  NAND2_X1 U23540 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20503), .ZN(
        n20508) );
  OR2_X1 U23541 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20508), .ZN(n20505) );
  AND2_X1 U23542 ( .A1(n20504), .A2(n20503), .ZN(n20536) );
  NOR3_X1 U23543 ( .A1(n10912), .A2(n20536), .A3(n20939), .ZN(n20509) );
  AOI21_X1 U23544 ( .B1(n20939), .B2(n20505), .A(n20509), .ZN(n20528) );
  AOI22_X1 U23545 ( .A1(n20528), .A2(n20692), .B1(n20691), .B2(n20536), .ZN(
        n20515) );
  NOR2_X1 U23546 ( .A1(n20507), .A2(n20506), .ZN(n20916) );
  INV_X1 U23547 ( .A(n20508), .ZN(n20513) );
  INV_X1 U23548 ( .A(n20536), .ZN(n20511) );
  AOI211_X1 U23549 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20511), .A(n20510), 
        .B(n20509), .ZN(n20512) );
  AOI22_X1 U23550 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20530), .B1(
        n20529), .B2(n20757), .ZN(n20514) );
  OAI211_X1 U23551 ( .C1(n20663), .C2(n20555), .A(n20515), .B(n20514), .ZN(
        P2_U3104) );
  AOI22_X1 U23552 ( .A1(n20528), .A2(n20730), .B1(n20536), .B2(n20727), .ZN(
        n20517) );
  AOI22_X1 U23553 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20530), .B1(
        n20529), .B2(n20729), .ZN(n20516) );
  OAI211_X1 U23554 ( .C1(n20666), .C2(n20555), .A(n20517), .B(n20516), .ZN(
        P2_U3105) );
  AOI22_X1 U23555 ( .A1(n20528), .A2(n20761), .B1(n20536), .B2(n20762), .ZN(
        n20519) );
  AOI22_X1 U23556 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20530), .B1(
        n20529), .B2(n20767), .ZN(n20518) );
  OAI211_X1 U23557 ( .C1(n20669), .C2(n20555), .A(n20519), .B(n20518), .ZN(
        P2_U3106) );
  AOI22_X1 U23558 ( .A1(n20528), .A2(n20771), .B1(n20536), .B2(n20772), .ZN(
        n20521) );
  AOI22_X1 U23559 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20530), .B1(
        n20529), .B2(n20776), .ZN(n20520) );
  OAI211_X1 U23560 ( .C1(n20672), .C2(n20555), .A(n20521), .B(n20520), .ZN(
        P2_U3107) );
  AOI22_X1 U23561 ( .A1(n20528), .A2(n20781), .B1(n20536), .B2(n20782), .ZN(
        n20523) );
  AOI22_X1 U23562 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20530), .B1(
        n20529), .B2(n20787), .ZN(n20522) );
  OAI211_X1 U23563 ( .C1(n20675), .C2(n20555), .A(n20523), .B(n20522), .ZN(
        P2_U3108) );
  AOI22_X1 U23564 ( .A1(n20528), .A2(n20791), .B1(n20536), .B2(n20792), .ZN(
        n20525) );
  AOI22_X1 U23565 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20530), .B1(
        n20529), .B2(n20796), .ZN(n20524) );
  OAI211_X1 U23566 ( .C1(n20678), .C2(n20555), .A(n20525), .B(n20524), .ZN(
        P2_U3109) );
  AOI22_X1 U23567 ( .A1(n20528), .A2(n20801), .B1(n20536), .B2(n20802), .ZN(
        n20527) );
  AOI22_X1 U23568 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20530), .B1(
        n20529), .B2(n20806), .ZN(n20526) );
  OAI211_X1 U23569 ( .C1(n20681), .C2(n20555), .A(n20527), .B(n20526), .ZN(
        P2_U3110) );
  AOI22_X1 U23570 ( .A1(n20528), .A2(n20811), .B1(n20536), .B2(n20812), .ZN(
        n20532) );
  AOI22_X1 U23571 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20530), .B1(
        n20529), .B2(n20820), .ZN(n20531) );
  OAI211_X1 U23572 ( .C1(n20688), .C2(n20555), .A(n20532), .B(n20531), .ZN(
        P2_U3111) );
  INV_X1 U23573 ( .A(n20650), .ZN(n20533) );
  INV_X1 U23574 ( .A(n20562), .ZN(n20564) );
  NAND3_X1 U23575 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20927), .A3(
        n20938), .ZN(n20570) );
  NOR2_X1 U23576 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20570), .ZN(
        n20556) );
  AOI22_X1 U23577 ( .A1(n20757), .A2(n20557), .B1(n20691), .B2(n20556), .ZN(
        n20542) );
  INV_X1 U23578 ( .A(n20537), .ZN(n20534) );
  OAI21_X1 U23579 ( .B1(n20535), .B2(n20556), .A(n20697), .ZN(n20559) );
  NOR2_X1 U23580 ( .A1(n20536), .A2(n20556), .ZN(n20539) );
  OAI21_X1 U23581 ( .B1(n20537), .B2(n20556), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20538) );
  AOI22_X1 U23582 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20559), .B1(
        n20692), .B2(n20558), .ZN(n20541) );
  OAI211_X1 U23583 ( .C1(n20663), .C2(n20592), .A(n20542), .B(n20541), .ZN(
        P2_U3112) );
  AOI22_X1 U23584 ( .A1(n20728), .A2(n20584), .B1(n20727), .B2(n20556), .ZN(
        n20544) );
  AOI22_X1 U23585 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20559), .B1(
        n20558), .B2(n20730), .ZN(n20543) );
  OAI211_X1 U23586 ( .C1(n20704), .C2(n20555), .A(n20544), .B(n20543), .ZN(
        P2_U3113) );
  AOI22_X1 U23587 ( .A1(n20767), .A2(n20557), .B1(n20762), .B2(n20556), .ZN(
        n20546) );
  AOI22_X1 U23588 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20559), .B1(
        n20558), .B2(n20761), .ZN(n20545) );
  OAI211_X1 U23589 ( .C1(n20669), .C2(n20592), .A(n20546), .B(n20545), .ZN(
        P2_U3114) );
  AOI22_X1 U23590 ( .A1(n20777), .A2(n20584), .B1(n20772), .B2(n20556), .ZN(
        n20548) );
  AOI22_X1 U23591 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20559), .B1(
        n20558), .B2(n20771), .ZN(n20547) );
  OAI211_X1 U23592 ( .C1(n20710), .C2(n20555), .A(n20548), .B(n20547), .ZN(
        P2_U3115) );
  AOI22_X1 U23593 ( .A1(n20787), .A2(n20557), .B1(n20782), .B2(n20556), .ZN(
        n20550) );
  AOI22_X1 U23594 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20559), .B1(
        n20558), .B2(n20781), .ZN(n20549) );
  OAI211_X1 U23595 ( .C1(n20675), .C2(n20592), .A(n20550), .B(n20549), .ZN(
        P2_U3116) );
  AOI22_X1 U23596 ( .A1(n20797), .A2(n20584), .B1(n20792), .B2(n20556), .ZN(
        n20552) );
  AOI22_X1 U23597 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20559), .B1(
        n20558), .B2(n20791), .ZN(n20551) );
  OAI211_X1 U23598 ( .C1(n20716), .C2(n20555), .A(n20552), .B(n20551), .ZN(
        P2_U3117) );
  AOI22_X1 U23599 ( .A1(n20807), .A2(n20584), .B1(n20802), .B2(n20556), .ZN(
        n20554) );
  AOI22_X1 U23600 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20559), .B1(
        n20558), .B2(n20801), .ZN(n20553) );
  OAI211_X1 U23601 ( .C1(n20719), .C2(n20555), .A(n20554), .B(n20553), .ZN(
        P2_U3118) );
  AOI22_X1 U23602 ( .A1(n20820), .A2(n20557), .B1(n20812), .B2(n20556), .ZN(
        n20561) );
  AOI22_X1 U23603 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20559), .B1(
        n20558), .B2(n20811), .ZN(n20560) );
  OAI211_X1 U23604 ( .C1(n20688), .C2(n20592), .A(n20561), .B(n20560), .ZN(
        P2_U3119) );
  NOR2_X1 U23605 ( .A1(n20947), .A2(n20570), .ZN(n20587) );
  AOI22_X1 U23606 ( .A1(n20757), .A2(n20584), .B1(n20691), .B2(n20587), .ZN(
        n20573) );
  INV_X1 U23607 ( .A(n20587), .ZN(n20598) );
  NAND2_X1 U23608 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20598), .ZN(n20567) );
  NOR2_X1 U23609 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n17491), .ZN(
        n20941) );
  AOI21_X1 U23610 ( .B1(n20565), .B2(n20564), .A(n20563), .ZN(n20568) );
  OAI22_X1 U23611 ( .A1(n20941), .A2(n20570), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20568), .ZN(n20566) );
  OAI211_X1 U23612 ( .C1(n10910), .C2(n20567), .A(n20566), .B(n20697), .ZN(
        n20589) );
  INV_X1 U23613 ( .A(n20568), .ZN(n20571) );
  OAI21_X1 U23614 ( .B1(n10910), .B2(n20587), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20569) );
  AOI22_X1 U23615 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20589), .B1(
        n20692), .B2(n20588), .ZN(n20572) );
  OAI211_X1 U23616 ( .C1(n20663), .C2(n20621), .A(n20573), .B(n20572), .ZN(
        P2_U3120) );
  AOI22_X1 U23617 ( .A1(n20728), .A2(n10555), .B1(n20727), .B2(n20587), .ZN(
        n20575) );
  AOI22_X1 U23618 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20589), .B1(
        n20730), .B2(n20588), .ZN(n20574) );
  OAI211_X1 U23619 ( .C1(n20704), .C2(n20592), .A(n20575), .B(n20574), .ZN(
        P2_U3121) );
  AOI22_X1 U23620 ( .A1(n20766), .A2(n10555), .B1(n20587), .B2(n20762), .ZN(
        n20577) );
  AOI22_X1 U23621 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20589), .B1(
        n20761), .B2(n20588), .ZN(n20576) );
  OAI211_X1 U23622 ( .C1(n20707), .C2(n20592), .A(n20577), .B(n20576), .ZN(
        P2_U3122) );
  AOI22_X1 U23623 ( .A1(n20776), .A2(n20584), .B1(n20587), .B2(n20772), .ZN(
        n20579) );
  AOI22_X1 U23624 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20589), .B1(
        n20771), .B2(n20588), .ZN(n20578) );
  OAI211_X1 U23625 ( .C1(n20672), .C2(n20621), .A(n20579), .B(n20578), .ZN(
        P2_U3123) );
  AOI22_X1 U23626 ( .A1(n20787), .A2(n20584), .B1(n20587), .B2(n20782), .ZN(
        n20581) );
  AOI22_X1 U23627 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20589), .B1(
        n20781), .B2(n20588), .ZN(n20580) );
  OAI211_X1 U23628 ( .C1(n20675), .C2(n20621), .A(n20581), .B(n20580), .ZN(
        P2_U3124) );
  AOI22_X1 U23629 ( .A1(n20796), .A2(n20584), .B1(n20587), .B2(n20792), .ZN(
        n20583) );
  AOI22_X1 U23630 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20589), .B1(
        n20791), .B2(n20588), .ZN(n20582) );
  OAI211_X1 U23631 ( .C1(n20678), .C2(n20621), .A(n20583), .B(n20582), .ZN(
        P2_U3125) );
  AOI22_X1 U23632 ( .A1(n20806), .A2(n20584), .B1(n20587), .B2(n20802), .ZN(
        n20586) );
  AOI22_X1 U23633 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20589), .B1(
        n20801), .B2(n20588), .ZN(n20585) );
  OAI211_X1 U23634 ( .C1(n20681), .C2(n20621), .A(n20586), .B(n20585), .ZN(
        P2_U3126) );
  AOI22_X1 U23635 ( .A1(n20818), .A2(n10555), .B1(n20587), .B2(n20812), .ZN(
        n20591) );
  AOI22_X1 U23636 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20589), .B1(
        n20811), .B2(n20588), .ZN(n20590) );
  OAI211_X1 U23637 ( .C1(n20726), .C2(n20592), .A(n20591), .B(n20590), .ZN(
        P2_U3127) );
  NAND3_X1 U23638 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20927), .ZN(n20625) );
  NOR2_X1 U23639 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20625), .ZN(
        n20616) );
  AOI22_X1 U23640 ( .A1(n20757), .A2(n10555), .B1(n20691), .B2(n20616), .ZN(
        n20603) );
  OAI21_X1 U23641 ( .B1(n10564), .B2(n10555), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20593) );
  NAND2_X1 U23642 ( .A1(n20593), .A2(n20958), .ZN(n20601) );
  INV_X1 U23643 ( .A(n20601), .ZN(n20595) );
  OAI21_X1 U23644 ( .B1(n10917), .B2(n20939), .A(n17491), .ZN(n20594) );
  AOI21_X1 U23645 ( .B1(n20595), .B2(n20598), .A(n20594), .ZN(n20596) );
  OAI21_X1 U23646 ( .B1(n20616), .B2(n20596), .A(n20697), .ZN(n20618) );
  INV_X1 U23647 ( .A(n20616), .ZN(n20597) );
  AND2_X1 U23648 ( .A1(n20598), .A2(n20597), .ZN(n20600) );
  OAI21_X1 U23649 ( .B1(n10917), .B2(n20616), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20599) );
  AOI22_X1 U23650 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20618), .B1(
        n20692), .B2(n20617), .ZN(n20602) );
  OAI211_X1 U23651 ( .C1(n20663), .C2(n20649), .A(n20603), .B(n20602), .ZN(
        P2_U3128) );
  AOI22_X1 U23652 ( .A1(n20729), .A2(n10555), .B1(n20727), .B2(n20616), .ZN(
        n20605) );
  AOI22_X1 U23653 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20618), .B1(
        n20730), .B2(n20617), .ZN(n20604) );
  OAI211_X1 U23654 ( .C1(n20666), .C2(n20649), .A(n20605), .B(n20604), .ZN(
        P2_U3129) );
  AOI22_X1 U23655 ( .A1(n20766), .A2(n10564), .B1(n20762), .B2(n20616), .ZN(
        n20607) );
  AOI22_X1 U23656 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20618), .B1(
        n20761), .B2(n20617), .ZN(n20606) );
  OAI211_X1 U23657 ( .C1(n20707), .C2(n20621), .A(n20607), .B(n20606), .ZN(
        P2_U3130) );
  AOI22_X1 U23658 ( .A1(n20777), .A2(n10564), .B1(n20616), .B2(n20772), .ZN(
        n20609) );
  AOI22_X1 U23659 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20618), .B1(
        n20771), .B2(n20617), .ZN(n20608) );
  OAI211_X1 U23660 ( .C1(n20710), .C2(n20621), .A(n20609), .B(n20608), .ZN(
        P2_U3131) );
  AOI22_X1 U23661 ( .A1(n20786), .A2(n10564), .B1(n20616), .B2(n20782), .ZN(
        n20611) );
  AOI22_X1 U23662 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20618), .B1(
        n20781), .B2(n20617), .ZN(n20610) );
  OAI211_X1 U23663 ( .C1(n20713), .C2(n20621), .A(n20611), .B(n20610), .ZN(
        P2_U3132) );
  AOI22_X1 U23664 ( .A1(n20797), .A2(n10564), .B1(n20616), .B2(n20792), .ZN(
        n20613) );
  AOI22_X1 U23665 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20618), .B1(
        n20791), .B2(n20617), .ZN(n20612) );
  OAI211_X1 U23666 ( .C1(n20716), .C2(n20621), .A(n20613), .B(n20612), .ZN(
        P2_U3133) );
  AOI22_X1 U23667 ( .A1(n20807), .A2(n10564), .B1(n20616), .B2(n20802), .ZN(
        n20615) );
  AOI22_X1 U23668 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20618), .B1(
        n20801), .B2(n20617), .ZN(n20614) );
  OAI211_X1 U23669 ( .C1(n20719), .C2(n20621), .A(n20615), .B(n20614), .ZN(
        P2_U3134) );
  AOI22_X1 U23670 ( .A1(n20818), .A2(n10564), .B1(n20812), .B2(n20616), .ZN(
        n20620) );
  AOI22_X1 U23671 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20618), .B1(
        n20811), .B2(n20617), .ZN(n20619) );
  OAI211_X1 U23672 ( .C1(n20726), .C2(n20621), .A(n20620), .B(n20619), .ZN(
        P2_U3135) );
  NOR2_X1 U23673 ( .A1(n20947), .A2(n20625), .ZN(n20644) );
  OAI21_X1 U23674 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20625), .A(n20939), 
        .ZN(n20623) );
  AOI22_X1 U23675 ( .A1(n20645), .A2(n20692), .B1(n20691), .B2(n20644), .ZN(
        n20631) );
  OR2_X1 U23676 ( .A1(n20624), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20694) );
  OAI22_X1 U23677 ( .A1(n20629), .A2(n20694), .B1(n20941), .B2(n20625), .ZN(
        n20627) );
  NAND3_X1 U23678 ( .A1(n20627), .A2(n20697), .A3(n20626), .ZN(n20646) );
  AOI22_X1 U23679 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20646), .B1(
        n20684), .B2(n20756), .ZN(n20630) );
  OAI211_X1 U23680 ( .C1(n20701), .C2(n20649), .A(n20631), .B(n20630), .ZN(
        P2_U3136) );
  AOI22_X1 U23681 ( .A1(n20645), .A2(n20730), .B1(n20727), .B2(n20644), .ZN(
        n20633) );
  AOI22_X1 U23682 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20646), .B1(
        n20684), .B2(n20728), .ZN(n20632) );
  OAI211_X1 U23683 ( .C1(n20704), .C2(n20649), .A(n20633), .B(n20632), .ZN(
        P2_U3137) );
  AOI22_X1 U23684 ( .A1(n20645), .A2(n20761), .B1(n20762), .B2(n20644), .ZN(
        n20635) );
  AOI22_X1 U23685 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20646), .B1(
        n20684), .B2(n20766), .ZN(n20634) );
  OAI211_X1 U23686 ( .C1(n20707), .C2(n20649), .A(n20635), .B(n20634), .ZN(
        P2_U3138) );
  AOI22_X1 U23687 ( .A1(n20645), .A2(n20771), .B1(n20772), .B2(n20644), .ZN(
        n20637) );
  AOI22_X1 U23688 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20646), .B1(
        n20684), .B2(n20777), .ZN(n20636) );
  OAI211_X1 U23689 ( .C1(n20710), .C2(n20649), .A(n20637), .B(n20636), .ZN(
        P2_U3139) );
  AOI22_X1 U23690 ( .A1(n20645), .A2(n20781), .B1(n20782), .B2(n20644), .ZN(
        n20639) );
  AOI22_X1 U23691 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20646), .B1(
        n20684), .B2(n20786), .ZN(n20638) );
  OAI211_X1 U23692 ( .C1(n20713), .C2(n20649), .A(n20639), .B(n20638), .ZN(
        P2_U3140) );
  AOI22_X1 U23693 ( .A1(n20645), .A2(n20791), .B1(n20792), .B2(n20644), .ZN(
        n20641) );
  AOI22_X1 U23694 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20646), .B1(
        n20684), .B2(n20797), .ZN(n20640) );
  OAI211_X1 U23695 ( .C1(n20716), .C2(n20649), .A(n20641), .B(n20640), .ZN(
        P2_U3141) );
  AOI22_X1 U23696 ( .A1(n20645), .A2(n20801), .B1(n20802), .B2(n20644), .ZN(
        n20643) );
  AOI22_X1 U23697 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20646), .B1(
        n20684), .B2(n20807), .ZN(n20642) );
  OAI211_X1 U23698 ( .C1(n20719), .C2(n20649), .A(n20643), .B(n20642), .ZN(
        P2_U3142) );
  AOI22_X1 U23699 ( .A1(n20645), .A2(n20811), .B1(n20812), .B2(n20644), .ZN(
        n20648) );
  AOI22_X1 U23700 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20646), .B1(
        n20684), .B2(n20818), .ZN(n20647) );
  OAI211_X1 U23701 ( .C1(n20726), .C2(n20649), .A(n20648), .B(n20647), .ZN(
        P2_U3143) );
  INV_X1 U23702 ( .A(n20651), .ZN(n20654) );
  NOR2_X1 U23703 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20693), .ZN(
        n20682) );
  OAI21_X1 U23704 ( .B1(n20652), .B2(n20682), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20653) );
  AOI22_X1 U23705 ( .A1(n20683), .A2(n20692), .B1(n20691), .B2(n20682), .ZN(
        n20662) );
  AOI21_X1 U23706 ( .B1(n20655), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20660) );
  OAI21_X1 U23707 ( .B1(n20656), .B2(n20684), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20657) );
  OAI21_X1 U23708 ( .B1(n20658), .B2(n20920), .A(n20657), .ZN(n20659) );
  OAI211_X1 U23709 ( .C1(n20682), .C2(n20660), .A(n20659), .B(n20697), .ZN(
        n20685) );
  AOI22_X1 U23710 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20685), .B1(
        n20684), .B2(n20757), .ZN(n20661) );
  OAI211_X1 U23711 ( .C1(n20663), .C2(n20725), .A(n20662), .B(n20661), .ZN(
        P2_U3144) );
  AOI22_X1 U23712 ( .A1(n20683), .A2(n20730), .B1(n20727), .B2(n20682), .ZN(
        n20665) );
  AOI22_X1 U23713 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20685), .B1(
        n20684), .B2(n20729), .ZN(n20664) );
  OAI211_X1 U23714 ( .C1(n20666), .C2(n20725), .A(n20665), .B(n20664), .ZN(
        P2_U3145) );
  AOI22_X1 U23715 ( .A1(n20683), .A2(n20761), .B1(n20762), .B2(n20682), .ZN(
        n20668) );
  AOI22_X1 U23716 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20685), .B1(
        n20684), .B2(n20767), .ZN(n20667) );
  OAI211_X1 U23717 ( .C1(n20669), .C2(n20725), .A(n20668), .B(n20667), .ZN(
        P2_U3146) );
  AOI22_X1 U23718 ( .A1(n20683), .A2(n20771), .B1(n20772), .B2(n20682), .ZN(
        n20671) );
  AOI22_X1 U23719 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20685), .B1(
        n20684), .B2(n20776), .ZN(n20670) );
  OAI211_X1 U23720 ( .C1(n20672), .C2(n20725), .A(n20671), .B(n20670), .ZN(
        P2_U3147) );
  AOI22_X1 U23721 ( .A1(n20683), .A2(n20781), .B1(n20782), .B2(n20682), .ZN(
        n20674) );
  AOI22_X1 U23722 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20685), .B1(
        n20684), .B2(n20787), .ZN(n20673) );
  OAI211_X1 U23723 ( .C1(n20675), .C2(n20725), .A(n20674), .B(n20673), .ZN(
        P2_U3148) );
  AOI22_X1 U23724 ( .A1(n20683), .A2(n20791), .B1(n20792), .B2(n20682), .ZN(
        n20677) );
  AOI22_X1 U23725 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20685), .B1(
        n20684), .B2(n20796), .ZN(n20676) );
  OAI211_X1 U23726 ( .C1(n20678), .C2(n20725), .A(n20677), .B(n20676), .ZN(
        P2_U3149) );
  AOI22_X1 U23727 ( .A1(n20683), .A2(n20801), .B1(n20802), .B2(n20682), .ZN(
        n20680) );
  AOI22_X1 U23728 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20685), .B1(
        n20684), .B2(n20806), .ZN(n20679) );
  OAI211_X1 U23729 ( .C1(n20681), .C2(n20725), .A(n20680), .B(n20679), .ZN(
        P2_U3150) );
  AOI22_X1 U23730 ( .A1(n20683), .A2(n20811), .B1(n20812), .B2(n20682), .ZN(
        n20687) );
  AOI22_X1 U23731 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20685), .B1(
        n20684), .B2(n20820), .ZN(n20686) );
  OAI211_X1 U23732 ( .C1(n20688), .C2(n20725), .A(n20687), .B(n20686), .ZN(
        P2_U3151) );
  OAI21_X1 U23733 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20693), .A(n20939), 
        .ZN(n20690) );
  AOI22_X1 U23734 ( .A1(n20721), .A2(n20692), .B1(n20691), .B2(n20720), .ZN(
        n20700) );
  OAI22_X1 U23735 ( .A1(n20695), .A2(n20694), .B1(n20941), .B2(n20693), .ZN(
        n20698) );
  NAND3_X1 U23736 ( .A1(n20698), .A2(n20697), .A3(n20696), .ZN(n20722) );
  AOI22_X1 U23737 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20722), .B1(
        n20747), .B2(n20756), .ZN(n20699) );
  OAI211_X1 U23738 ( .C1(n20701), .C2(n20725), .A(n20700), .B(n20699), .ZN(
        P2_U3152) );
  AOI22_X1 U23739 ( .A1(n20721), .A2(n20730), .B1(n20727), .B2(n20720), .ZN(
        n20703) );
  AOI22_X1 U23740 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20722), .B1(
        n20747), .B2(n20728), .ZN(n20702) );
  OAI211_X1 U23741 ( .C1(n20704), .C2(n20725), .A(n20703), .B(n20702), .ZN(
        P2_U3153) );
  AOI22_X1 U23742 ( .A1(n20721), .A2(n20761), .B1(n20762), .B2(n20720), .ZN(
        n20706) );
  AOI22_X1 U23743 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20722), .B1(
        n20747), .B2(n20766), .ZN(n20705) );
  OAI211_X1 U23744 ( .C1(n20707), .C2(n20725), .A(n20706), .B(n20705), .ZN(
        P2_U3154) );
  AOI22_X1 U23745 ( .A1(n20721), .A2(n20771), .B1(n20772), .B2(n20720), .ZN(
        n20709) );
  AOI22_X1 U23746 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20722), .B1(
        n20747), .B2(n20777), .ZN(n20708) );
  OAI211_X1 U23747 ( .C1(n20710), .C2(n20725), .A(n20709), .B(n20708), .ZN(
        P2_U3155) );
  AOI22_X1 U23748 ( .A1(n20721), .A2(n20781), .B1(n20782), .B2(n20720), .ZN(
        n20712) );
  AOI22_X1 U23749 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20722), .B1(
        n20747), .B2(n20786), .ZN(n20711) );
  OAI211_X1 U23750 ( .C1(n20713), .C2(n20725), .A(n20712), .B(n20711), .ZN(
        P2_U3156) );
  AOI22_X1 U23751 ( .A1(n20721), .A2(n20791), .B1(n20792), .B2(n20720), .ZN(
        n20715) );
  AOI22_X1 U23752 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20722), .B1(
        n20747), .B2(n20797), .ZN(n20714) );
  OAI211_X1 U23753 ( .C1(n20716), .C2(n20725), .A(n20715), .B(n20714), .ZN(
        P2_U3157) );
  AOI22_X1 U23754 ( .A1(n20721), .A2(n20801), .B1(n20802), .B2(n20720), .ZN(
        n20718) );
  AOI22_X1 U23755 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20722), .B1(
        n20747), .B2(n20807), .ZN(n20717) );
  OAI211_X1 U23756 ( .C1(n20719), .C2(n20725), .A(n20718), .B(n20717), .ZN(
        P2_U3158) );
  AOI22_X1 U23757 ( .A1(n20721), .A2(n20811), .B1(n20812), .B2(n20720), .ZN(
        n20724) );
  AOI22_X1 U23758 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20722), .B1(
        n20747), .B2(n20818), .ZN(n20723) );
  OAI211_X1 U23759 ( .C1(n20726), .C2(n20725), .A(n20724), .B(n20723), .ZN(
        P2_U3159) );
  AOI22_X1 U23760 ( .A1(n20728), .A2(n20821), .B1(n20746), .B2(n20727), .ZN(
        n20732) );
  AOI22_X1 U23761 ( .A1(n20730), .A2(n20748), .B1(n20747), .B2(n20729), .ZN(
        n20731) );
  OAI211_X1 U23762 ( .C1(n20752), .C2(n10823), .A(n20732), .B(n20731), .ZN(
        P2_U3161) );
  INV_X1 U23763 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n20735) );
  AOI22_X1 U23764 ( .A1(n20766), .A2(n20821), .B1(n20746), .B2(n20762), .ZN(
        n20734) );
  AOI22_X1 U23765 ( .A1(n20761), .A2(n20748), .B1(n20747), .B2(n20767), .ZN(
        n20733) );
  OAI211_X1 U23766 ( .C1(n20752), .C2(n20735), .A(n20734), .B(n20733), .ZN(
        P2_U3162) );
  AOI22_X1 U23767 ( .A1(n20776), .A2(n20747), .B1(n20746), .B2(n20772), .ZN(
        n20737) );
  AOI22_X1 U23768 ( .A1(n20771), .A2(n20748), .B1(n20821), .B2(n20777), .ZN(
        n20736) );
  OAI211_X1 U23769 ( .C1(n20752), .C2(n10790), .A(n20737), .B(n20736), .ZN(
        P2_U3163) );
  INV_X1 U23770 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n20740) );
  AOI22_X1 U23771 ( .A1(n20786), .A2(n20821), .B1(n20746), .B2(n20782), .ZN(
        n20739) );
  AOI22_X1 U23772 ( .A1(n20781), .A2(n20748), .B1(n20747), .B2(n20787), .ZN(
        n20738) );
  OAI211_X1 U23773 ( .C1(n20752), .C2(n20740), .A(n20739), .B(n20738), .ZN(
        P2_U3164) );
  AOI22_X1 U23774 ( .A1(n20796), .A2(n20747), .B1(n20746), .B2(n20792), .ZN(
        n20742) );
  AOI22_X1 U23775 ( .A1(n20791), .A2(n20748), .B1(n20821), .B2(n20797), .ZN(
        n20741) );
  OAI211_X1 U23776 ( .C1(n20752), .C2(n10901), .A(n20742), .B(n20741), .ZN(
        P2_U3165) );
  AOI22_X1 U23777 ( .A1(n20806), .A2(n20747), .B1(n20746), .B2(n20802), .ZN(
        n20744) );
  AOI22_X1 U23778 ( .A1(n20801), .A2(n20748), .B1(n20821), .B2(n20807), .ZN(
        n20743) );
  OAI211_X1 U23779 ( .C1(n20752), .C2(n20745), .A(n20744), .B(n20743), .ZN(
        P2_U3166) );
  INV_X1 U23780 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n20751) );
  AOI22_X1 U23781 ( .A1(n20820), .A2(n20747), .B1(n20746), .B2(n20812), .ZN(
        n20750) );
  AOI22_X1 U23782 ( .A1(n20811), .A2(n20748), .B1(n20821), .B2(n20818), .ZN(
        n20749) );
  OAI211_X1 U23783 ( .C1(n20752), .C2(n20751), .A(n20750), .B(n20749), .ZN(
        P2_U3167) );
  OAI22_X1 U23784 ( .A1(n20816), .A2(n20754), .B1(n20814), .B2(n20753), .ZN(
        n20755) );
  INV_X1 U23785 ( .A(n20755), .ZN(n20759) );
  AOI22_X1 U23786 ( .A1(n20821), .A2(n20757), .B1(n20819), .B2(n20756), .ZN(
        n20758) );
  OAI211_X1 U23787 ( .C1(n20825), .C2(n20760), .A(n20759), .B(n20758), .ZN(
        P2_U3168) );
  INV_X1 U23788 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n20770) );
  INV_X1 U23789 ( .A(n20761), .ZN(n20764) );
  INV_X1 U23790 ( .A(n20762), .ZN(n20763) );
  OAI22_X1 U23791 ( .A1(n20816), .A2(n20764), .B1(n20814), .B2(n20763), .ZN(
        n20765) );
  INV_X1 U23792 ( .A(n20765), .ZN(n20769) );
  AOI22_X1 U23793 ( .A1(n20821), .A2(n20767), .B1(n20819), .B2(n20766), .ZN(
        n20768) );
  OAI211_X1 U23794 ( .C1(n20825), .C2(n20770), .A(n20769), .B(n20768), .ZN(
        P2_U3170) );
  INV_X1 U23795 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n20780) );
  INV_X1 U23796 ( .A(n20771), .ZN(n20774) );
  INV_X1 U23797 ( .A(n20772), .ZN(n20773) );
  OAI22_X1 U23798 ( .A1(n20816), .A2(n20774), .B1(n20814), .B2(n20773), .ZN(
        n20775) );
  INV_X1 U23799 ( .A(n20775), .ZN(n20779) );
  AOI22_X1 U23800 ( .A1(n20819), .A2(n20777), .B1(n20821), .B2(n20776), .ZN(
        n20778) );
  OAI211_X1 U23801 ( .C1(n20825), .C2(n20780), .A(n20779), .B(n20778), .ZN(
        P2_U3171) );
  INV_X1 U23802 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n20790) );
  INV_X1 U23803 ( .A(n20781), .ZN(n20784) );
  INV_X1 U23804 ( .A(n20782), .ZN(n20783) );
  OAI22_X1 U23805 ( .A1(n20816), .A2(n20784), .B1(n20814), .B2(n20783), .ZN(
        n20785) );
  INV_X1 U23806 ( .A(n20785), .ZN(n20789) );
  AOI22_X1 U23807 ( .A1(n20821), .A2(n20787), .B1(n20819), .B2(n20786), .ZN(
        n20788) );
  OAI211_X1 U23808 ( .C1(n20825), .C2(n20790), .A(n20789), .B(n20788), .ZN(
        P2_U3172) );
  INV_X1 U23809 ( .A(n20791), .ZN(n20794) );
  INV_X1 U23810 ( .A(n20792), .ZN(n20793) );
  OAI22_X1 U23811 ( .A1(n20816), .A2(n20794), .B1(n20814), .B2(n20793), .ZN(
        n20795) );
  INV_X1 U23812 ( .A(n20795), .ZN(n20799) );
  AOI22_X1 U23813 ( .A1(n20819), .A2(n20797), .B1(n20821), .B2(n20796), .ZN(
        n20798) );
  OAI211_X1 U23814 ( .C1(n20825), .C2(n20800), .A(n20799), .B(n20798), .ZN(
        P2_U3173) );
  INV_X1 U23815 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n20810) );
  INV_X1 U23816 ( .A(n20801), .ZN(n20804) );
  INV_X1 U23817 ( .A(n20802), .ZN(n20803) );
  OAI22_X1 U23818 ( .A1(n20816), .A2(n20804), .B1(n20814), .B2(n20803), .ZN(
        n20805) );
  INV_X1 U23819 ( .A(n20805), .ZN(n20809) );
  AOI22_X1 U23820 ( .A1(n20819), .A2(n20807), .B1(n20821), .B2(n20806), .ZN(
        n20808) );
  OAI211_X1 U23821 ( .C1(n20825), .C2(n20810), .A(n20809), .B(n20808), .ZN(
        P2_U3174) );
  INV_X1 U23822 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n20824) );
  INV_X1 U23823 ( .A(n20811), .ZN(n20815) );
  INV_X1 U23824 ( .A(n20812), .ZN(n20813) );
  OAI22_X1 U23825 ( .A1(n20816), .A2(n20815), .B1(n20814), .B2(n20813), .ZN(
        n20817) );
  INV_X1 U23826 ( .A(n20817), .ZN(n20823) );
  AOI22_X1 U23827 ( .A1(n20821), .A2(n20820), .B1(n20819), .B2(n20818), .ZN(
        n20822) );
  OAI211_X1 U23828 ( .C1(n20825), .C2(n20824), .A(n20823), .B(n20822), .ZN(
        P2_U3175) );
  AND2_X1 U23829 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20828), .ZN(
        P2_U3179) );
  AND2_X1 U23830 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20828), .ZN(
        P2_U3180) );
  AND2_X1 U23831 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20828), .ZN(
        P2_U3181) );
  AND2_X1 U23832 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20828), .ZN(
        P2_U3182) );
  AND2_X1 U23833 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20828), .ZN(
        P2_U3183) );
  AND2_X1 U23834 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20828), .ZN(
        P2_U3184) );
  AND2_X1 U23835 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20828), .ZN(
        P2_U3185) );
  AND2_X1 U23836 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20828), .ZN(
        P2_U3186) );
  AND2_X1 U23837 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20828), .ZN(
        P2_U3187) );
  AND2_X1 U23838 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20828), .ZN(
        P2_U3188) );
  AND2_X1 U23839 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20828), .ZN(
        P2_U3189) );
  AND2_X1 U23840 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20828), .ZN(
        P2_U3190) );
  AND2_X1 U23841 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20828), .ZN(
        P2_U3191) );
  AND2_X1 U23842 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20828), .ZN(
        P2_U3192) );
  AND2_X1 U23843 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20828), .ZN(
        P2_U3193) );
  AND2_X1 U23844 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20828), .ZN(
        P2_U3194) );
  AND2_X1 U23845 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20828), .ZN(
        P2_U3195) );
  AND2_X1 U23846 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20828), .ZN(
        P2_U3196) );
  NOR2_X1 U23847 ( .A1(n20826), .A2(n20909), .ZN(P2_U3197) );
  AND2_X1 U23848 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20828), .ZN(
        P2_U3198) );
  AND2_X1 U23849 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20828), .ZN(
        P2_U3199) );
  NOR2_X1 U23850 ( .A1(n20827), .A2(n20909), .ZN(P2_U3200) );
  AND2_X1 U23851 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20828), .ZN(P2_U3201) );
  AND2_X1 U23852 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20828), .ZN(P2_U3202) );
  AND2_X1 U23853 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20828), .ZN(P2_U3203) );
  AND2_X1 U23854 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20828), .ZN(P2_U3204) );
  AND2_X1 U23855 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20828), .ZN(P2_U3205) );
  AND2_X1 U23856 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20828), .ZN(P2_U3206) );
  AND2_X1 U23857 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20828), .ZN(P2_U3207) );
  AND2_X1 U23858 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20828), .ZN(P2_U3208) );
  INV_X1 U23859 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20974) );
  NOR2_X1 U23860 ( .A1(n20966), .A2(n20839), .ZN(n20837) );
  OR3_X1 U23861 ( .A1(n20974), .A2(n20829), .A3(n20837), .ZN(n20830) );
  NOR3_X1 U23862 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .A3(n21653), .ZN(n20843) );
  AOI21_X1 U23863 ( .B1(n20846), .B2(n20830), .A(n20843), .ZN(n20831) );
  OAI221_X1 U23864 ( .B1(n20832), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .C1(
        n20832), .C2(n21647), .A(n20831), .ZN(P2_U3209) );
  AOI21_X1 U23865 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21647), .A(n20846), 
        .ZN(n20840) );
  NOR3_X1 U23866 ( .A1(n20840), .A2(n20974), .A3(n20829), .ZN(n20833) );
  NOR2_X1 U23867 ( .A1(n20833), .A2(n20837), .ZN(n20835) );
  OAI211_X1 U23868 ( .C1(n21647), .C2(n20836), .A(n20835), .B(n20834), .ZN(
        P2_U3210) );
  AOI22_X1 U23869 ( .A1(n20838), .A2(n20974), .B1(n20837), .B2(n21653), .ZN(
        n20845) );
  OAI21_X1 U23870 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n20844) );
  NOR2_X1 U23871 ( .A1(n20846), .A2(n20839), .ZN(n20841) );
  AOI21_X1 U23872 ( .B1(n20841), .B2(n20963), .A(n20840), .ZN(n20842) );
  OAI22_X1 U23873 ( .A1(n20845), .A2(n20844), .B1(n20843), .B2(n20842), .ZN(
        P2_U3211) );
  OAI222_X1 U23874 ( .A1(n20898), .A2(n20849), .B1(n20848), .B2(n20979), .C1(
        n20847), .C2(n20899), .ZN(P2_U3212) );
  OAI222_X1 U23875 ( .A1(n20898), .A2(n20851), .B1(n20850), .B2(n20979), .C1(
        n20849), .C2(n20899), .ZN(P2_U3213) );
  OAI222_X1 U23876 ( .A1(n20898), .A2(n20853), .B1(n20852), .B2(n20979), .C1(
        n20851), .C2(n20899), .ZN(P2_U3214) );
  OAI222_X1 U23877 ( .A1(n20898), .A2(n17148), .B1(n20854), .B2(n20979), .C1(
        n20853), .C2(n20899), .ZN(P2_U3215) );
  OAI222_X1 U23878 ( .A1(n20898), .A2(n20856), .B1(n20855), .B2(n20979), .C1(
        n17148), .C2(n20899), .ZN(P2_U3216) );
  OAI222_X1 U23879 ( .A1(n20898), .A2(n20858), .B1(n20857), .B2(n20979), .C1(
        n20856), .C2(n20899), .ZN(P2_U3217) );
  OAI222_X1 U23880 ( .A1(n20898), .A2(n17115), .B1(n20859), .B2(n20979), .C1(
        n20858), .C2(n20899), .ZN(P2_U3218) );
  OAI222_X1 U23881 ( .A1(n20898), .A2(n20861), .B1(n20860), .B2(n20979), .C1(
        n17115), .C2(n20899), .ZN(P2_U3219) );
  OAI222_X1 U23882 ( .A1(n20898), .A2(n20863), .B1(n20862), .B2(n20979), .C1(
        n20861), .C2(n20899), .ZN(P2_U3220) );
  OAI222_X1 U23883 ( .A1(n20898), .A2(n20865), .B1(n20864), .B2(n20979), .C1(
        n20863), .C2(n20899), .ZN(P2_U3221) );
  OAI222_X1 U23884 ( .A1(n20898), .A2(n20867), .B1(n20866), .B2(n20979), .C1(
        n20865), .C2(n20899), .ZN(P2_U3222) );
  OAI222_X1 U23885 ( .A1(n20898), .A2(n20869), .B1(n20868), .B2(n20979), .C1(
        n20867), .C2(n20899), .ZN(P2_U3223) );
  OAI222_X1 U23886 ( .A1(n20898), .A2(n20871), .B1(n20870), .B2(n20979), .C1(
        n20869), .C2(n20899), .ZN(P2_U3224) );
  OAI222_X1 U23887 ( .A1(n20898), .A2(n20873), .B1(n20872), .B2(n20979), .C1(
        n20871), .C2(n20899), .ZN(P2_U3225) );
  OAI222_X1 U23888 ( .A1(n20898), .A2(n20875), .B1(n20874), .B2(n20979), .C1(
        n20873), .C2(n20899), .ZN(P2_U3226) );
  OAI222_X1 U23889 ( .A1(n20898), .A2(n20877), .B1(n20876), .B2(n20979), .C1(
        n20875), .C2(n20899), .ZN(P2_U3227) );
  OAI222_X1 U23890 ( .A1(n20898), .A2(n16992), .B1(n20878), .B2(n20979), .C1(
        n20877), .C2(n20899), .ZN(P2_U3228) );
  OAI222_X1 U23891 ( .A1(n20898), .A2(n20880), .B1(n20879), .B2(n20979), .C1(
        n16992), .C2(n20899), .ZN(P2_U3229) );
  OAI222_X1 U23892 ( .A1(n20898), .A2(n16982), .B1(n20881), .B2(n20979), .C1(
        n20880), .C2(n20899), .ZN(P2_U3230) );
  OAI222_X1 U23893 ( .A1(n20898), .A2(n20883), .B1(n20882), .B2(n20979), .C1(
        n16982), .C2(n20899), .ZN(P2_U3231) );
  OAI222_X1 U23894 ( .A1(n20898), .A2(n16968), .B1(n20884), .B2(n20979), .C1(
        n20883), .C2(n20899), .ZN(P2_U3232) );
  OAI222_X1 U23895 ( .A1(n20898), .A2(n20886), .B1(n20885), .B2(n20979), .C1(
        n16968), .C2(n20899), .ZN(P2_U3233) );
  OAI222_X1 U23896 ( .A1(n20898), .A2(n16950), .B1(n20887), .B2(n20979), .C1(
        n20886), .C2(n20899), .ZN(P2_U3234) );
  OAI222_X1 U23897 ( .A1(n20898), .A2(n20889), .B1(n20888), .B2(n20979), .C1(
        n16950), .C2(n20899), .ZN(P2_U3235) );
  OAI222_X1 U23898 ( .A1(n20898), .A2(n20891), .B1(n20890), .B2(n20979), .C1(
        n20889), .C2(n20899), .ZN(P2_U3236) );
  INV_X1 U23899 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20894) );
  OAI222_X1 U23900 ( .A1(n20898), .A2(n20894), .B1(n20892), .B2(n20979), .C1(
        n20891), .C2(n20899), .ZN(P2_U3237) );
  OAI222_X1 U23901 ( .A1(n20899), .A2(n20894), .B1(n20893), .B2(n20979), .C1(
        n14894), .C2(n20898), .ZN(P2_U3238) );
  OAI222_X1 U23902 ( .A1(n20898), .A2(n20896), .B1(n20895), .B2(n20979), .C1(
        n14894), .C2(n20899), .ZN(P2_U3239) );
  INV_X1 U23903 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20900) );
  OAI222_X1 U23904 ( .A1(n20898), .A2(n20900), .B1(n20897), .B2(n20979), .C1(
        n20896), .C2(n20899), .ZN(P2_U3240) );
  OAI222_X1 U23905 ( .A1(n20898), .A2(n11561), .B1(n20901), .B2(n20979), .C1(
        n20900), .C2(n20899), .ZN(P2_U3241) );
  INV_X1 U23906 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20902) );
  AOI22_X1 U23907 ( .A1(n20979), .A2(n20903), .B1(n20902), .B2(n20976), .ZN(
        P2_U3585) );
  MUX2_X1 U23908 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20979), .Z(P2_U3586) );
  MUX2_X1 U23909 ( .A(P2_BE_N_REG_1__SCAN_IN), .B(P2_BYTEENABLE_REG_1__SCAN_IN), .S(n20979), .Z(P2_U3587) );
  INV_X1 U23910 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20904) );
  AOI22_X1 U23911 ( .A1(n20979), .A2(n20905), .B1(n20904), .B2(n20976), .ZN(
        P2_U3588) );
  OAI21_X1 U23912 ( .B1(n20909), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20907), 
        .ZN(n20906) );
  INV_X1 U23913 ( .A(n20906), .ZN(P2_U3591) );
  OAI21_X1 U23914 ( .B1(n20909), .B2(n20908), .A(n20907), .ZN(P2_U3592) );
  INV_X1 U23915 ( .A(n20943), .ZN(n20915) );
  NOR3_X1 U23916 ( .A1(n20912), .A2(n20911), .A3(n20910), .ZN(n20914) );
  AND2_X1 U23917 ( .A1(n20958), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20928) );
  NAND2_X1 U23918 ( .A1(n20913), .A2(n20928), .ZN(n20922) );
  OAI21_X1 U23919 ( .B1(n20915), .B2(n20914), .A(n20922), .ZN(n20925) );
  AOI222_X1 U23920 ( .A1(n20925), .A2(n20918), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20917), .C1(n20958), .C2(n20916), .ZN(n20919) );
  AOI22_X1 U23921 ( .A1(n20948), .A2(n20920), .B1(n20919), .B2(n20945), .ZN(
        P2_U3602) );
  NAND2_X1 U23922 ( .A1(n20922), .A2(n20921), .ZN(n20924) );
  AOI22_X1 U23923 ( .A1(n20925), .A2(n20924), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20923), .ZN(n20926) );
  AOI22_X1 U23924 ( .A1(n20948), .A2(n20927), .B1(n20926), .B2(n20945), .ZN(
        P2_U3603) );
  INV_X1 U23925 ( .A(n20928), .ZN(n20933) );
  INV_X1 U23926 ( .A(n20929), .ZN(n20930) );
  NAND2_X1 U23927 ( .A1(n20943), .A2(n20930), .ZN(n20932) );
  MUX2_X1 U23928 ( .A(n20933), .B(n20932), .S(n20931), .Z(n20936) );
  NAND2_X1 U23929 ( .A1(n20934), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20935) );
  AND2_X1 U23930 ( .A1(n20936), .A2(n20935), .ZN(n20937) );
  AOI22_X1 U23931 ( .A1(n20948), .A2(n20938), .B1(n20937), .B2(n20945), .ZN(
        P2_U3604) );
  NOR2_X1 U23932 ( .A1(n20940), .A2(n20939), .ZN(n20942) );
  AOI211_X1 U23933 ( .C1(n20944), .C2(n20943), .A(n20942), .B(n20941), .ZN(
        n20946) );
  AOI22_X1 U23934 ( .A1(n20948), .A2(n20947), .B1(n20946), .B2(n20945), .ZN(
        P2_U3605) );
  INV_X1 U23935 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20949) );
  AOI22_X1 U23936 ( .A1(n20979), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20949), 
        .B2(n20976), .ZN(P2_U3608) );
  OAI22_X1 U23937 ( .A1(n20953), .A2(n20952), .B1(n20951), .B2(n20950), .ZN(
        n20954) );
  OR2_X1 U23938 ( .A1(n20955), .A2(n20954), .ZN(n20957) );
  MUX2_X1 U23939 ( .A(P2_MORE_REG_SCAN_IN), .B(n20957), .S(n20956), .Z(
        P2_U3609) );
  AOI21_X1 U23940 ( .B1(n20959), .B2(n17491), .A(n20958), .ZN(n20960) );
  OAI211_X1 U23941 ( .C1(n20963), .C2(n20962), .A(n20961), .B(n20960), .ZN(
        n20975) );
  AOI211_X1 U23942 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n20965), .A(n11573), 
        .B(n20964), .ZN(n20972) );
  OAI211_X1 U23943 ( .C1(n20968), .C2(n20967), .A(P2_STATE2_REG_2__SCAN_IN), 
        .B(n20966), .ZN(n20970) );
  AND2_X1 U23944 ( .A1(n20970), .A2(n20969), .ZN(n20971) );
  OAI21_X1 U23945 ( .B1(n20972), .B2(n20971), .A(n20975), .ZN(n20973) );
  OAI21_X1 U23946 ( .B1(n20975), .B2(n20974), .A(n20973), .ZN(P2_U3610) );
  INV_X1 U23947 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n20977) );
  AOI22_X1 U23948 ( .A1(n20979), .A2(n20978), .B1(n20977), .B2(n20976), .ZN(
        P2_U3611) );
  AOI21_X1 U23949 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n12627), .A(n21657), 
        .ZN(n20987) );
  INV_X1 U23950 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20980) );
  AOI21_X1 U23951 ( .B1(n20987), .B2(n20980), .A(n21770), .ZN(P1_U2802) );
  INV_X1 U23952 ( .A(n20981), .ZN(n20983) );
  OAI21_X1 U23953 ( .B1(n20983), .B2(n20982), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20984) );
  OAI21_X1 U23954 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20985), .A(n20984), 
        .ZN(P1_U2803) );
  NOR2_X1 U23955 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20988) );
  OAI21_X1 U23956 ( .B1(n20988), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21755), .ZN(
        n20986) );
  OAI21_X1 U23957 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21755), .A(n20986), 
        .ZN(P1_U2804) );
  NOR2_X1 U23958 ( .A1(n21770), .A2(n20987), .ZN(n21730) );
  OAI21_X1 U23959 ( .B1(BS16), .B2(n20988), .A(n21730), .ZN(n21728) );
  OAI21_X1 U23960 ( .B1(n21730), .B2(n21426), .A(n21728), .ZN(P1_U2805) );
  OAI21_X1 U23961 ( .B1(n20991), .B2(n20990), .A(n20989), .ZN(P1_U2806) );
  NOR4_X1 U23962 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20995) );
  NOR4_X1 U23963 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20994) );
  NOR4_X1 U23964 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20993) );
  NOR4_X1 U23965 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20992) );
  NAND4_X1 U23966 ( .A1(n20995), .A2(n20994), .A3(n20993), .A4(n20992), .ZN(
        n21001) );
  NOR4_X1 U23967 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20999) );
  AOI211_X1 U23968 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_14__SCAN_IN), .B(
        P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n20998) );
  NOR4_X1 U23969 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_11__SCAN_IN), .A3(P1_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20997) );
  NOR4_X1 U23970 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20996) );
  NAND4_X1 U23971 ( .A1(n20999), .A2(n20998), .A3(n20997), .A4(n20996), .ZN(
        n21000) );
  NOR2_X1 U23972 ( .A1(n21001), .A2(n21000), .ZN(n21754) );
  INV_X1 U23973 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21723) );
  NOR3_X1 U23974 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n21003) );
  OAI21_X1 U23975 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n21003), .A(n21754), .ZN(
        n21002) );
  OAI21_X1 U23976 ( .B1(n21754), .B2(n21723), .A(n21002), .ZN(P1_U2807) );
  INV_X1 U23977 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21729) );
  AOI21_X1 U23978 ( .B1(n21660), .B2(n21729), .A(n21003), .ZN(n21004) );
  INV_X1 U23979 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21720) );
  INV_X1 U23980 ( .A(n21754), .ZN(n21751) );
  AOI22_X1 U23981 ( .A1(n21754), .A2(n21004), .B1(n21720), .B2(n21751), .ZN(
        P1_U2808) );
  INV_X1 U23982 ( .A(n21005), .ZN(n21101) );
  AOI22_X1 U23983 ( .A1(n21101), .A2(n21041), .B1(n21040), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n21006) );
  OAI211_X1 U23984 ( .C1(n21068), .C2(n21007), .A(n21006), .B(n21042), .ZN(
        n21008) );
  AOI221_X1 U23985 ( .B1(n21010), .B2(n21677), .C1(n21009), .C2(
        P1_REIP_REG_9__SCAN_IN), .A(n21008), .ZN(n21015) );
  INV_X1 U23986 ( .A(n21011), .ZN(n21102) );
  AOI22_X1 U23987 ( .A1(n21102), .A2(n21036), .B1(n9698), .B2(n21012), .ZN(
        n21014) );
  NAND2_X1 U23988 ( .A1(n21015), .A2(n21014), .ZN(P1_U2831) );
  NAND3_X1 U23989 ( .A1(n21081), .A2(n21029), .A3(n21673), .ZN(n21016) );
  OAI211_X1 U23990 ( .C1(n21068), .C2(n21017), .A(n21016), .B(n21042), .ZN(
        n21018) );
  AOI21_X1 U23991 ( .B1(n21040), .B2(P1_EBX_REG_7__SCAN_IN), .A(n21018), .ZN(
        n21019) );
  OAI21_X1 U23992 ( .B1(n21086), .B2(n21020), .A(n21019), .ZN(n21021) );
  AOI21_X1 U23993 ( .B1(n21022), .B2(n21036), .A(n21021), .ZN(n21024) );
  OAI21_X1 U23994 ( .B1(n21029), .B2(n21087), .A(n21074), .ZN(n21026) );
  NAND2_X1 U23995 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n21026), .ZN(n21023) );
  OAI211_X1 U23996 ( .C1(n21094), .C2(n21025), .A(n21024), .B(n21023), .ZN(
        P1_U2833) );
  AOI22_X1 U23997 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n21082), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n21026), .ZN(n21034) );
  INV_X1 U23998 ( .A(n21027), .ZN(n21032) );
  OAI21_X1 U23999 ( .B1(n21089), .B2(n13013), .A(n21042), .ZN(n21031) );
  NOR3_X1 U24000 ( .A1(n21087), .A2(n21029), .A3(n21028), .ZN(n21030) );
  AOI211_X1 U24001 ( .C1(n21041), .C2(n21032), .A(n21031), .B(n21030), .ZN(
        n21033) );
  NAND2_X1 U24002 ( .A1(n21034), .A2(n21033), .ZN(n21035) );
  AOI21_X1 U24003 ( .B1(n21037), .B2(n21036), .A(n21035), .ZN(n21038) );
  OAI21_X1 U24004 ( .B1(n21039), .B2(n9697), .A(n21038), .ZN(P1_U2834) );
  NOR2_X1 U24005 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n21087), .ZN(n21046) );
  AOI22_X1 U24006 ( .A1(n21041), .A2(n21105), .B1(n21040), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n21043) );
  OAI211_X1 U24007 ( .C1(n21068), .C2(n21044), .A(n21043), .B(n21042), .ZN(
        n21045) );
  AOI21_X1 U24008 ( .B1(n21046), .B2(n21047), .A(n21045), .ZN(n21050) );
  OR2_X1 U24009 ( .A1(n21087), .A2(n21047), .ZN(n21048) );
  NAND2_X1 U24010 ( .A1(n21048), .A2(n21074), .ZN(n21061) );
  AOI22_X1 U24011 ( .A1(n21106), .A2(n21096), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n21061), .ZN(n21049) );
  OAI211_X1 U24012 ( .C1(n21051), .C2(n9697), .A(n21050), .B(n21049), .ZN(
        P1_U2835) );
  NOR3_X1 U24013 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n21087), .A3(n21052), .ZN(
        n21059) );
  INV_X1 U24014 ( .A(n21053), .ZN(n21055) );
  OAI22_X1 U24015 ( .A1(n21055), .A2(n21054), .B1(n14549), .B2(n21068), .ZN(
        n21058) );
  OAI22_X1 U24016 ( .A1(n21086), .A2(n21056), .B1(n21089), .B2(n13003), .ZN(
        n21057) );
  NOR4_X1 U24017 ( .A1(n21060), .A2(n21059), .A3(n21058), .A4(n21057), .ZN(
        n21064) );
  AOI22_X1 U24018 ( .A1(n21062), .A2(n21096), .B1(P1_REIP_REG_4__SCAN_IN), 
        .B2(n21061), .ZN(n21063) );
  OAI211_X1 U24019 ( .C1(n21065), .C2(n21094), .A(n21064), .B(n21063), .ZN(
        P1_U2836) );
  INV_X1 U24020 ( .A(n21066), .ZN(n21079) );
  AND2_X1 U24021 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n21075) );
  NAND2_X1 U24022 ( .A1(n21075), .A2(n21665), .ZN(n21067) );
  OAI22_X1 U24023 ( .A1(n21086), .A2(n21109), .B1(n21087), .B2(n21067), .ZN(
        n21072) );
  INV_X1 U24024 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n21115) );
  OAI22_X1 U24025 ( .A1(n21089), .A2(n21115), .B1(n21069), .B2(n21068), .ZN(
        n21071) );
  AND2_X1 U24026 ( .A1(n21739), .A2(n21083), .ZN(n21070) );
  NOR3_X1 U24027 ( .A1(n21072), .A2(n21071), .A3(n21070), .ZN(n21078) );
  INV_X1 U24028 ( .A(n21073), .ZN(n21113) );
  OAI21_X1 U24029 ( .B1(n21087), .B2(n21075), .A(n21074), .ZN(n21076) );
  AOI22_X1 U24030 ( .A1(n21113), .A2(n21096), .B1(P1_REIP_REG_3__SCAN_IN), 
        .B2(n21076), .ZN(n21077) );
  OAI211_X1 U24031 ( .C1(n21079), .C2(n9697), .A(n21078), .B(n21077), .ZN(
        P1_U2837) );
  AOI21_X1 U24032 ( .B1(n21081), .B2(n21660), .A(n21080), .ZN(n21100) );
  INV_X1 U24033 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21663) );
  AOI22_X1 U24034 ( .A1(n21083), .A2(n21192), .B1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n21082), .ZN(n21084) );
  OAI21_X1 U24035 ( .B1(n21086), .B2(n21085), .A(n21084), .ZN(n21092) );
  OR3_X1 U24036 ( .A1(n21087), .A2(P1_REIP_REG_2__SCAN_IN), .A3(n21660), .ZN(
        n21088) );
  OAI21_X1 U24037 ( .B1(n21090), .B2(n21089), .A(n21088), .ZN(n21091) );
  NOR2_X1 U24038 ( .A1(n21092), .A2(n21091), .ZN(n21099) );
  NOR2_X1 U24039 ( .A1(n9697), .A2(n21093), .ZN(n21095) );
  AOI21_X1 U24040 ( .B1(n21097), .B2(n21096), .A(n21095), .ZN(n21098) );
  OAI211_X1 U24041 ( .C1(n21100), .C2(n21663), .A(n21099), .B(n21098), .ZN(
        P1_U2838) );
  AOI22_X1 U24042 ( .A1(n21102), .A2(n21112), .B1(n21111), .B2(n21101), .ZN(
        n21103) );
  OAI21_X1 U24043 ( .B1(n21116), .B2(n21104), .A(n21103), .ZN(P1_U2863) );
  AOI22_X1 U24044 ( .A1(n21106), .A2(n21112), .B1(n21111), .B2(n21105), .ZN(
        n21107) );
  OAI21_X1 U24045 ( .B1(n21116), .B2(n21108), .A(n21107), .ZN(P1_U2867) );
  INV_X1 U24046 ( .A(n21109), .ZN(n21110) );
  AOI22_X1 U24047 ( .A1(n21113), .A2(n21112), .B1(n21111), .B2(n21110), .ZN(
        n21114) );
  OAI21_X1 U24048 ( .B1(n21116), .B2(n21115), .A(n21114), .ZN(P1_U2869) );
  INV_X1 U24049 ( .A(n21117), .ZN(n21120) );
  AOI22_X1 U24050 ( .A1(n21120), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n21760), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n21118) );
  OAI21_X1 U24051 ( .B1(n21119), .B2(n21139), .A(n21118), .ZN(P1_U2918) );
  AOI22_X1 U24052 ( .A1(n21120), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n21760), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n21121) );
  OAI21_X1 U24053 ( .B1(n21122), .B2(n21139), .A(n21121), .ZN(P1_U2919) );
  AOI22_X1 U24054 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n21123) );
  OAI21_X1 U24055 ( .B1(n21124), .B2(n21151), .A(n21123), .ZN(P1_U2921) );
  AOI22_X1 U24056 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n21125) );
  OAI21_X1 U24057 ( .B1(n21126), .B2(n21151), .A(n21125), .ZN(P1_U2922) );
  INV_X1 U24058 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n21128) );
  AOI22_X1 U24059 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n21127) );
  OAI21_X1 U24060 ( .B1(n21128), .B2(n21151), .A(n21127), .ZN(P1_U2923) );
  INV_X1 U24061 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n21130) );
  AOI22_X1 U24062 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n21129) );
  OAI21_X1 U24063 ( .B1(n21130), .B2(n21151), .A(n21129), .ZN(P1_U2924) );
  AOI22_X1 U24064 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n21131) );
  OAI21_X1 U24065 ( .B1(n15886), .B2(n21151), .A(n21131), .ZN(P1_U2925) );
  AOI22_X1 U24066 ( .A1(P1_EAX_REG_10__SCAN_IN), .A2(n21132), .B1(n13826), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n21133) );
  OAI21_X1 U24067 ( .B1(n21134), .B2(n21142), .A(n21133), .ZN(P1_U2926) );
  AOI22_X1 U24068 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n21135) );
  OAI21_X1 U24069 ( .B1(n14956), .B2(n21151), .A(n21135), .ZN(P1_U2927) );
  AOI22_X1 U24070 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n21136) );
  OAI21_X1 U24071 ( .B1(n14927), .B2(n21151), .A(n21136), .ZN(P1_U2928) );
  OAI222_X1 U24072 ( .A1(n21142), .A2(n21138), .B1(n21151), .B2(n14757), .C1(
        n21139), .C2(n21137), .ZN(P1_U2929) );
  INV_X1 U24073 ( .A(P1_LWORD_REG_6__SCAN_IN), .ZN(n21141) );
  OAI222_X1 U24074 ( .A1(n21142), .A2(n21141), .B1(n21151), .B2(n14749), .C1(
        n21140), .C2(n21139), .ZN(P1_U2930) );
  AOI22_X1 U24075 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n21143) );
  OAI21_X1 U24076 ( .B1(n14652), .B2(n21151), .A(n21143), .ZN(P1_U2931) );
  AOI22_X1 U24077 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n21144) );
  OAI21_X1 U24078 ( .B1(n21145), .B2(n21151), .A(n21144), .ZN(P1_U2932) );
  AOI22_X1 U24079 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n21146) );
  OAI21_X1 U24080 ( .B1(n21147), .B2(n21151), .A(n21146), .ZN(P1_U2933) );
  AOI22_X1 U24081 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n21148) );
  OAI21_X1 U24082 ( .B1(n13880), .B2(n21151), .A(n21148), .ZN(P1_U2934) );
  AOI22_X1 U24083 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n21149) );
  OAI21_X1 U24084 ( .B1(n13681), .B2(n21151), .A(n21149), .ZN(P1_U2935) );
  AOI22_X1 U24085 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n21760), .B1(n13826), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n21150) );
  OAI21_X1 U24086 ( .B1(n21152), .B2(n21151), .A(n21150), .ZN(P1_U2936) );
  AOI22_X1 U24087 ( .A1(n21170), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n21169), .ZN(n21154) );
  NAND2_X1 U24088 ( .A1(n21161), .A2(n21153), .ZN(n21163) );
  NAND2_X1 U24089 ( .A1(n21154), .A2(n21163), .ZN(P1_U2947) );
  AOI22_X1 U24090 ( .A1(n21155), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n21169), .ZN(n21157) );
  NAND2_X1 U24091 ( .A1(n21161), .A2(n21156), .ZN(n21165) );
  NAND2_X1 U24092 ( .A1(n21157), .A2(n21165), .ZN(P1_U2948) );
  AOI22_X1 U24093 ( .A1(n21170), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n21169), .ZN(n21159) );
  NAND2_X1 U24094 ( .A1(n21161), .A2(n21158), .ZN(n21167) );
  NAND2_X1 U24095 ( .A1(n21159), .A2(n21167), .ZN(P1_U2949) );
  AOI22_X1 U24096 ( .A1(n21170), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n21169), .ZN(n21162) );
  NAND2_X1 U24097 ( .A1(n21161), .A2(n21160), .ZN(n21171) );
  NAND2_X1 U24098 ( .A1(n21162), .A2(n21171), .ZN(P1_U2950) );
  AOI22_X1 U24099 ( .A1(n21170), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n21169), .ZN(n21164) );
  NAND2_X1 U24100 ( .A1(n21164), .A2(n21163), .ZN(P1_U2962) );
  AOI22_X1 U24101 ( .A1(n21170), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n21169), .ZN(n21166) );
  NAND2_X1 U24102 ( .A1(n21166), .A2(n21165), .ZN(P1_U2963) );
  AOI22_X1 U24103 ( .A1(n21170), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n21169), .ZN(n21168) );
  NAND2_X1 U24104 ( .A1(n21168), .A2(n21167), .ZN(P1_U2964) );
  AOI22_X1 U24105 ( .A1(n21170), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n21169), .ZN(n21172) );
  NAND2_X1 U24106 ( .A1(n21172), .A2(n21171), .ZN(P1_U2965) );
  OAI22_X1 U24107 ( .A1(n21176), .A2(n21175), .B1(n21174), .B2(n21173), .ZN(
        n21177) );
  INV_X1 U24108 ( .A(n21177), .ZN(n21183) );
  OAI22_X1 U24109 ( .A1(n21180), .A2(n21179), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21178), .ZN(n21181) );
  NAND3_X1 U24110 ( .A1(n21183), .A2(n21182), .A3(n21181), .ZN(P1_U3031) );
  NOR2_X1 U24111 ( .A1(n21184), .A2(n21747), .ZN(P1_U3032) );
  NOR2_X1 U24112 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21290) );
  INV_X1 U24113 ( .A(n21290), .ZN(n21187) );
  NOR2_X1 U24114 ( .A1(n21187), .A2(n21522), .ZN(n21195) );
  INV_X1 U24115 ( .A(n21195), .ZN(n21220) );
  OAI22_X1 U24116 ( .A1(n21636), .A2(n21538), .B1(n21220), .B2(n21291), .ZN(
        n21188) );
  INV_X1 U24117 ( .A(n21188), .ZN(n21201) );
  NAND3_X1 U24118 ( .A1(n21251), .A2(n21586), .A3(n21636), .ZN(n21191) );
  NAND2_X1 U24119 ( .A1(n21191), .A2(n21742), .ZN(n21196) );
  OR2_X1 U24120 ( .A1(n21739), .A2(n21192), .ZN(n21254) );
  OR2_X1 U24121 ( .A1(n21254), .A2(n21526), .ZN(n21198) );
  INV_X1 U24122 ( .A(n21394), .ZN(n21193) );
  NAND2_X1 U24123 ( .A1(n21193), .A2(n21393), .ZN(n21197) );
  AOI22_X1 U24124 ( .A1(n21196), .A2(n21198), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21197), .ZN(n21194) );
  INV_X1 U24125 ( .A(n21196), .ZN(n21199) );
  AOI22_X1 U24126 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n21223), .B1(
        n21577), .B2(n21222), .ZN(n21200) );
  OAI211_X1 U24127 ( .C1(n21590), .C2(n21251), .A(n21201), .B(n21200), .ZN(
        P1_U3033) );
  OAI22_X1 U24128 ( .A1(n21636), .A2(n21542), .B1(n21220), .B2(n21304), .ZN(
        n21202) );
  INV_X1 U24129 ( .A(n21202), .ZN(n21204) );
  AOI22_X1 U24130 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n21223), .B1(
        n21591), .B2(n21222), .ZN(n21203) );
  OAI211_X1 U24131 ( .C1(n21596), .C2(n21251), .A(n21204), .B(n21203), .ZN(
        P1_U3034) );
  OAI22_X1 U24132 ( .A1(n21636), .A2(n21546), .B1(n21220), .B2(n21308), .ZN(
        n21205) );
  INV_X1 U24133 ( .A(n21205), .ZN(n21207) );
  AOI22_X1 U24134 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n21223), .B1(
        n21597), .B2(n21222), .ZN(n21206) );
  OAI211_X1 U24135 ( .C1(n21602), .C2(n21251), .A(n21207), .B(n21206), .ZN(
        P1_U3035) );
  OAI22_X1 U24136 ( .A1(n21636), .A2(n21550), .B1(n21220), .B2(n21312), .ZN(
        n21208) );
  INV_X1 U24137 ( .A(n21208), .ZN(n21210) );
  AOI22_X1 U24138 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n21223), .B1(
        n21603), .B2(n21222), .ZN(n21209) );
  OAI211_X1 U24139 ( .C1(n21608), .C2(n21251), .A(n21210), .B(n21209), .ZN(
        P1_U3036) );
  OAI22_X1 U24140 ( .A1(n21636), .A2(n21554), .B1(n21220), .B2(n21316), .ZN(
        n21211) );
  INV_X1 U24141 ( .A(n21211), .ZN(n21213) );
  AOI22_X1 U24142 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n21223), .B1(
        n21609), .B2(n21222), .ZN(n21212) );
  OAI211_X1 U24143 ( .C1(n21614), .C2(n21251), .A(n21213), .B(n21212), .ZN(
        P1_U3037) );
  OAI22_X1 U24144 ( .A1(n21636), .A2(n21558), .B1(n21220), .B2(n21320), .ZN(
        n21214) );
  INV_X1 U24145 ( .A(n21214), .ZN(n21216) );
  AOI22_X1 U24146 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n21223), .B1(
        n21615), .B2(n21222), .ZN(n21215) );
  OAI211_X1 U24147 ( .C1(n21620), .C2(n21251), .A(n21216), .B(n21215), .ZN(
        P1_U3038) );
  OAI22_X1 U24148 ( .A1(n21636), .A2(n21562), .B1(n21220), .B2(n21324), .ZN(
        n21217) );
  INV_X1 U24149 ( .A(n21217), .ZN(n21219) );
  AOI22_X1 U24150 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n21223), .B1(
        n21621), .B2(n21222), .ZN(n21218) );
  OAI211_X1 U24151 ( .C1(n21626), .C2(n21251), .A(n21219), .B(n21218), .ZN(
        P1_U3039) );
  OAI22_X1 U24152 ( .A1(n21636), .A2(n21570), .B1(n21220), .B2(n21328), .ZN(
        n21221) );
  INV_X1 U24153 ( .A(n21221), .ZN(n21225) );
  AOI22_X1 U24154 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n21223), .B1(
        n21627), .B2(n21222), .ZN(n21224) );
  OAI211_X1 U24155 ( .C1(n21637), .C2(n21251), .A(n21225), .B(n21224), .ZN(
        P1_U3040) );
  INV_X1 U24156 ( .A(n21254), .ZN(n21296) );
  NAND2_X1 U24157 ( .A1(n21290), .A2(n21575), .ZN(n21226) );
  NOR2_X1 U24158 ( .A1(n21422), .A2(n21226), .ZN(n21245) );
  AOI21_X1 U24159 ( .B1(n21296), .B2(n21423), .A(n21245), .ZN(n21227) );
  OAI22_X1 U24160 ( .A1(n21227), .A2(n21584), .B1(n21226), .B2(n21641), .ZN(
        n21246) );
  AOI22_X1 U24161 ( .A1(n21246), .A2(n21577), .B1(n21578), .B2(n21245), .ZN(
        n21231) );
  INV_X1 U24162 ( .A(n21226), .ZN(n21229) );
  OAI21_X1 U24163 ( .B1(n21293), .B2(n21426), .A(n21227), .ZN(n21228) );
  OAI221_X1 U24164 ( .B1(n21586), .B2(n21229), .C1(n21584), .C2(n21228), .A(
        n21582), .ZN(n21248) );
  INV_X1 U24165 ( .A(n21283), .ZN(n21247) );
  AOI22_X1 U24166 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n21248), .B1(
        n21247), .B2(n21523), .ZN(n21230) );
  OAI211_X1 U24167 ( .C1(n21538), .C2(n21251), .A(n21231), .B(n21230), .ZN(
        P1_U3041) );
  AOI22_X1 U24168 ( .A1(n21246), .A2(n21591), .B1(n21592), .B2(n21245), .ZN(
        n21233) );
  INV_X1 U24169 ( .A(n21251), .ZN(n21240) );
  AOI22_X1 U24170 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n21248), .B1(
        n21240), .B2(n21593), .ZN(n21232) );
  OAI211_X1 U24171 ( .C1(n21596), .C2(n21283), .A(n21233), .B(n21232), .ZN(
        P1_U3042) );
  AOI22_X1 U24172 ( .A1(n21246), .A2(n21597), .B1(n21598), .B2(n21245), .ZN(
        n21235) );
  AOI22_X1 U24173 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n21248), .B1(
        n21240), .B2(n21599), .ZN(n21234) );
  OAI211_X1 U24174 ( .C1(n21602), .C2(n21283), .A(n21235), .B(n21234), .ZN(
        P1_U3043) );
  AOI22_X1 U24175 ( .A1(n21246), .A2(n21603), .B1(n21604), .B2(n21245), .ZN(
        n21237) );
  AOI22_X1 U24176 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n21248), .B1(
        n21247), .B2(n21547), .ZN(n21236) );
  OAI211_X1 U24177 ( .C1(n21550), .C2(n21251), .A(n21237), .B(n21236), .ZN(
        P1_U3044) );
  AOI22_X1 U24178 ( .A1(n21246), .A2(n21609), .B1(n21610), .B2(n21245), .ZN(
        n21239) );
  AOI22_X1 U24179 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n21248), .B1(
        n21240), .B2(n21611), .ZN(n21238) );
  OAI211_X1 U24180 ( .C1(n21614), .C2(n21283), .A(n21239), .B(n21238), .ZN(
        P1_U3045) );
  AOI22_X1 U24181 ( .A1(n21246), .A2(n21615), .B1(n21616), .B2(n21245), .ZN(
        n21242) );
  AOI22_X1 U24182 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n21248), .B1(
        n21240), .B2(n21617), .ZN(n21241) );
  OAI211_X1 U24183 ( .C1(n21620), .C2(n21283), .A(n21242), .B(n21241), .ZN(
        P1_U3046) );
  AOI22_X1 U24184 ( .A1(n21246), .A2(n21621), .B1(n21622), .B2(n21245), .ZN(
        n21244) );
  AOI22_X1 U24185 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n21248), .B1(
        n21247), .B2(n21559), .ZN(n21243) );
  OAI211_X1 U24186 ( .C1(n21562), .C2(n21251), .A(n21244), .B(n21243), .ZN(
        P1_U3047) );
  AOI22_X1 U24187 ( .A1(n21246), .A2(n21627), .B1(n21630), .B2(n21245), .ZN(
        n21250) );
  AOI22_X1 U24188 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n21248), .B1(
        n21247), .B2(n21563), .ZN(n21249) );
  OAI211_X1 U24189 ( .C1(n21570), .C2(n21251), .A(n21250), .B(n21249), .ZN(
        P1_U3048) );
  NAND2_X1 U24190 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21290), .ZN(
        n21299) );
  OR2_X1 U24191 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21299), .ZN(
        n21282) );
  OAI22_X1 U24192 ( .A1(n21335), .A2(n21590), .B1(n21282), .B2(n21291), .ZN(
        n21252) );
  INV_X1 U24193 ( .A(n21252), .ZN(n21263) );
  NAND3_X1 U24194 ( .A1(n21335), .A2(n21283), .A3(n21586), .ZN(n21253) );
  NAND2_X1 U24195 ( .A1(n21253), .A2(n21742), .ZN(n21257) );
  OR2_X1 U24196 ( .A1(n21254), .A2(n21453), .ZN(n21260) );
  AOI22_X1 U24197 ( .A1(n21257), .A2(n21260), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21282), .ZN(n21256) );
  NAND3_X1 U24198 ( .A1(n21463), .A2(n21256), .A3(n21255), .ZN(n21286) );
  INV_X1 U24199 ( .A(n21257), .ZN(n21261) );
  INV_X1 U24200 ( .A(n21258), .ZN(n21259) );
  AOI22_X1 U24201 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n21286), .B1(
        n21577), .B2(n21285), .ZN(n21262) );
  OAI211_X1 U24202 ( .C1(n21538), .C2(n21283), .A(n21263), .B(n21262), .ZN(
        P1_U3049) );
  OAI22_X1 U24203 ( .A1(n21283), .A2(n21542), .B1(n21282), .B2(n21304), .ZN(
        n21264) );
  INV_X1 U24204 ( .A(n21264), .ZN(n21266) );
  AOI22_X1 U24205 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n21286), .B1(
        n21591), .B2(n21285), .ZN(n21265) );
  OAI211_X1 U24206 ( .C1(n21596), .C2(n21335), .A(n21266), .B(n21265), .ZN(
        P1_U3050) );
  OAI22_X1 U24207 ( .A1(n21283), .A2(n21546), .B1(n21282), .B2(n21308), .ZN(
        n21267) );
  INV_X1 U24208 ( .A(n21267), .ZN(n21269) );
  AOI22_X1 U24209 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n21286), .B1(
        n21597), .B2(n21285), .ZN(n21268) );
  OAI211_X1 U24210 ( .C1(n21602), .C2(n21335), .A(n21269), .B(n21268), .ZN(
        P1_U3051) );
  OAI22_X1 U24211 ( .A1(n21335), .A2(n21608), .B1(n21282), .B2(n21312), .ZN(
        n21270) );
  INV_X1 U24212 ( .A(n21270), .ZN(n21272) );
  AOI22_X1 U24213 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n21286), .B1(
        n21603), .B2(n21285), .ZN(n21271) );
  OAI211_X1 U24214 ( .C1(n21550), .C2(n21283), .A(n21272), .B(n21271), .ZN(
        P1_U3052) );
  OAI22_X1 U24215 ( .A1(n21283), .A2(n21554), .B1(n21282), .B2(n21316), .ZN(
        n21273) );
  INV_X1 U24216 ( .A(n21273), .ZN(n21275) );
  AOI22_X1 U24217 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n21286), .B1(
        n21609), .B2(n21285), .ZN(n21274) );
  OAI211_X1 U24218 ( .C1(n21614), .C2(n21335), .A(n21275), .B(n21274), .ZN(
        P1_U3053) );
  OAI22_X1 U24219 ( .A1(n21283), .A2(n21558), .B1(n21282), .B2(n21320), .ZN(
        n21276) );
  INV_X1 U24220 ( .A(n21276), .ZN(n21278) );
  AOI22_X1 U24221 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n21286), .B1(
        n21615), .B2(n21285), .ZN(n21277) );
  OAI211_X1 U24222 ( .C1(n21620), .C2(n21335), .A(n21278), .B(n21277), .ZN(
        P1_U3054) );
  OAI22_X1 U24223 ( .A1(n21283), .A2(n21562), .B1(n21282), .B2(n21324), .ZN(
        n21279) );
  INV_X1 U24224 ( .A(n21279), .ZN(n21281) );
  AOI22_X1 U24225 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n21286), .B1(
        n21621), .B2(n21285), .ZN(n21280) );
  OAI211_X1 U24226 ( .C1(n21626), .C2(n21335), .A(n21281), .B(n21280), .ZN(
        P1_U3055) );
  OAI22_X1 U24227 ( .A1(n21283), .A2(n21570), .B1(n21282), .B2(n21328), .ZN(
        n21284) );
  INV_X1 U24228 ( .A(n21284), .ZN(n21288) );
  AOI22_X1 U24229 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n21286), .B1(
        n21627), .B2(n21285), .ZN(n21287) );
  OAI211_X1 U24230 ( .C1(n21637), .C2(n21335), .A(n21288), .B(n21287), .ZN(
        P1_U3056) );
  NAND2_X1 U24231 ( .A1(n21290), .A2(n21289), .ZN(n21329) );
  OAI22_X1 U24232 ( .A1(n21335), .A2(n21538), .B1(n21329), .B2(n21291), .ZN(
        n21292) );
  INV_X1 U24233 ( .A(n21292), .ZN(n21303) );
  OR2_X1 U24234 ( .A1(n21293), .A2(n21580), .ZN(n21294) );
  INV_X1 U24235 ( .A(n21329), .ZN(n21295) );
  AOI21_X1 U24236 ( .B1(n21296), .B2(n21572), .A(n21295), .ZN(n21301) );
  AOI22_X1 U24237 ( .A1(n21298), .A2(n21301), .B1(n21584), .B2(n21299), .ZN(
        n21297) );
  NAND2_X1 U24238 ( .A1(n21582), .A2(n21297), .ZN(n21332) );
  INV_X1 U24239 ( .A(n21298), .ZN(n21300) );
  AOI22_X1 U24240 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n21332), .B1(
        n21577), .B2(n21331), .ZN(n21302) );
  OAI211_X1 U24241 ( .C1(n21590), .C2(n21349), .A(n21303), .B(n21302), .ZN(
        P1_U3057) );
  OAI22_X1 U24242 ( .A1(n21335), .A2(n21542), .B1(n21329), .B2(n21304), .ZN(
        n21305) );
  INV_X1 U24243 ( .A(n21305), .ZN(n21307) );
  AOI22_X1 U24244 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n21332), .B1(
        n21591), .B2(n21331), .ZN(n21306) );
  OAI211_X1 U24245 ( .C1(n21596), .C2(n21349), .A(n21307), .B(n21306), .ZN(
        P1_U3058) );
  OAI22_X1 U24246 ( .A1(n21335), .A2(n21546), .B1(n21329), .B2(n21308), .ZN(
        n21309) );
  INV_X1 U24247 ( .A(n21309), .ZN(n21311) );
  AOI22_X1 U24248 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n21332), .B1(
        n21597), .B2(n21331), .ZN(n21310) );
  OAI211_X1 U24249 ( .C1(n21602), .C2(n21349), .A(n21311), .B(n21310), .ZN(
        P1_U3059) );
  OAI22_X1 U24250 ( .A1(n21335), .A2(n21550), .B1(n21329), .B2(n21312), .ZN(
        n21313) );
  INV_X1 U24251 ( .A(n21313), .ZN(n21315) );
  AOI22_X1 U24252 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n21332), .B1(
        n21603), .B2(n21331), .ZN(n21314) );
  OAI211_X1 U24253 ( .C1(n21608), .C2(n21349), .A(n21315), .B(n21314), .ZN(
        P1_U3060) );
  OAI22_X1 U24254 ( .A1(n21335), .A2(n21554), .B1(n21329), .B2(n21316), .ZN(
        n21317) );
  INV_X1 U24255 ( .A(n21317), .ZN(n21319) );
  AOI22_X1 U24256 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n21332), .B1(
        n21609), .B2(n21331), .ZN(n21318) );
  OAI211_X1 U24257 ( .C1(n21614), .C2(n21349), .A(n21319), .B(n21318), .ZN(
        P1_U3061) );
  OAI22_X1 U24258 ( .A1(n21335), .A2(n21558), .B1(n21329), .B2(n21320), .ZN(
        n21321) );
  INV_X1 U24259 ( .A(n21321), .ZN(n21323) );
  AOI22_X1 U24260 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n21332), .B1(
        n21615), .B2(n21331), .ZN(n21322) );
  OAI211_X1 U24261 ( .C1(n21620), .C2(n21349), .A(n21323), .B(n21322), .ZN(
        P1_U3062) );
  OAI22_X1 U24262 ( .A1(n21349), .A2(n21626), .B1(n21329), .B2(n21324), .ZN(
        n21325) );
  INV_X1 U24263 ( .A(n21325), .ZN(n21327) );
  AOI22_X1 U24264 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n21332), .B1(
        n21621), .B2(n21331), .ZN(n21326) );
  OAI211_X1 U24265 ( .C1(n21562), .C2(n21335), .A(n21327), .B(n21326), .ZN(
        P1_U3063) );
  OAI22_X1 U24266 ( .A1(n21349), .A2(n21637), .B1(n21329), .B2(n21328), .ZN(
        n21330) );
  INV_X1 U24267 ( .A(n21330), .ZN(n21334) );
  AOI22_X1 U24268 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n21332), .B1(
        n21627), .B2(n21331), .ZN(n21333) );
  OAI211_X1 U24269 ( .C1(n21570), .C2(n21335), .A(n21334), .B(n21333), .ZN(
        P1_U3064) );
  INV_X1 U24270 ( .A(n21393), .ZN(n21336) );
  OAI33_X1 U24271 ( .A1(n21338), .A2(n21526), .A3(n21584), .B1(n21394), .B2(
        n21336), .B3(n21533), .ZN(n21356) );
  AOI22_X1 U24272 ( .A1(n9873), .A2(n21577), .B1(n21578), .B2(n10557), .ZN(
        n21341) );
  INV_X1 U24273 ( .A(n21388), .ZN(n21346) );
  OAI21_X1 U24274 ( .B1(n21357), .B2(n21346), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21337) );
  OAI21_X1 U24275 ( .B1(n21526), .B2(n21338), .A(n21337), .ZN(n21339) );
  AOI22_X1 U24276 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n21358), .B1(
        n21346), .B2(n21523), .ZN(n21340) );
  OAI211_X1 U24277 ( .C1(n21538), .C2(n21349), .A(n21341), .B(n21340), .ZN(
        P1_U3065) );
  AOI22_X1 U24278 ( .A1(n9873), .A2(n21591), .B1(n21592), .B2(n10557), .ZN(
        n21343) );
  AOI22_X1 U24279 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n21358), .B1(
        n21357), .B2(n21593), .ZN(n21342) );
  OAI211_X1 U24280 ( .C1(n21596), .C2(n21388), .A(n21343), .B(n21342), .ZN(
        P1_U3066) );
  AOI22_X1 U24281 ( .A1(n9873), .A2(n21597), .B1(n21598), .B2(n10557), .ZN(
        n21345) );
  AOI22_X1 U24282 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n21358), .B1(
        n21357), .B2(n21599), .ZN(n21344) );
  OAI211_X1 U24283 ( .C1(n21602), .C2(n21388), .A(n21345), .B(n21344), .ZN(
        P1_U3067) );
  AOI22_X1 U24284 ( .A1(n9873), .A2(n21603), .B1(n21604), .B2(n10557), .ZN(
        n21348) );
  AOI22_X1 U24285 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n21358), .B1(
        n21346), .B2(n21547), .ZN(n21347) );
  OAI211_X1 U24286 ( .C1(n21550), .C2(n21349), .A(n21348), .B(n21347), .ZN(
        P1_U3068) );
  AOI22_X1 U24287 ( .A1(n9873), .A2(n21609), .B1(n21610), .B2(n10557), .ZN(
        n21351) );
  AOI22_X1 U24288 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n21358), .B1(
        n21357), .B2(n21611), .ZN(n21350) );
  OAI211_X1 U24289 ( .C1(n21614), .C2(n21388), .A(n21351), .B(n21350), .ZN(
        P1_U3069) );
  AOI22_X1 U24290 ( .A1(n9873), .A2(n21615), .B1(n21616), .B2(n10557), .ZN(
        n21353) );
  AOI22_X1 U24291 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n21358), .B1(
        n21357), .B2(n21617), .ZN(n21352) );
  OAI211_X1 U24292 ( .C1(n21620), .C2(n21388), .A(n21353), .B(n21352), .ZN(
        P1_U3070) );
  AOI22_X1 U24293 ( .A1(n9873), .A2(n21621), .B1(n21622), .B2(n10557), .ZN(
        n21355) );
  AOI22_X1 U24294 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n21358), .B1(
        n21357), .B2(n21623), .ZN(n21354) );
  OAI211_X1 U24295 ( .C1(n21626), .C2(n21388), .A(n21355), .B(n21354), .ZN(
        P1_U3071) );
  AOI22_X1 U24296 ( .A1(n9873), .A2(n21627), .B1(n21630), .B2(n10557), .ZN(
        n21360) );
  AOI22_X1 U24297 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n21358), .B1(
        n21357), .B2(n21631), .ZN(n21359) );
  OAI211_X1 U24298 ( .C1(n21637), .C2(n21388), .A(n21360), .B(n21359), .ZN(
        P1_U3072) );
  NOR2_X1 U24299 ( .A1(n21361), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21367) );
  INV_X1 U24300 ( .A(n21367), .ZN(n21363) );
  NOR2_X1 U24301 ( .A1(n21422), .A2(n21363), .ZN(n21383) );
  AOI21_X1 U24302 ( .B1(n21362), .B2(n21423), .A(n21383), .ZN(n21364) );
  OAI22_X1 U24303 ( .A1(n21364), .A2(n21584), .B1(n21363), .B2(n21641), .ZN(
        n21382) );
  AOI22_X1 U24304 ( .A1(n21578), .A2(n21383), .B1(n21382), .B2(n21577), .ZN(
        n21369) );
  OAI21_X1 U24305 ( .B1(n21365), .B2(n21426), .A(n21364), .ZN(n21366) );
  OAI221_X1 U24306 ( .B1(n21586), .B2(n21367), .C1(n21584), .C2(n21366), .A(
        n21582), .ZN(n21385) );
  AOI22_X1 U24307 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n21385), .B1(
        n21384), .B2(n21523), .ZN(n21368) );
  OAI211_X1 U24308 ( .C1(n21538), .C2(n21388), .A(n21369), .B(n21368), .ZN(
        P1_U3073) );
  AOI22_X1 U24309 ( .A1(n21592), .A2(n21383), .B1(n21382), .B2(n21591), .ZN(
        n21371) );
  AOI22_X1 U24310 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n21385), .B1(
        n21384), .B2(n21539), .ZN(n21370) );
  OAI211_X1 U24311 ( .C1(n21542), .C2(n21388), .A(n21371), .B(n21370), .ZN(
        P1_U3074) );
  AOI22_X1 U24312 ( .A1(n21598), .A2(n21383), .B1(n21382), .B2(n21597), .ZN(
        n21373) );
  AOI22_X1 U24313 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n21385), .B1(
        n21384), .B2(n21543), .ZN(n21372) );
  OAI211_X1 U24314 ( .C1(n21546), .C2(n21388), .A(n21373), .B(n21372), .ZN(
        P1_U3075) );
  AOI22_X1 U24315 ( .A1(n21604), .A2(n21383), .B1(n21382), .B2(n21603), .ZN(
        n21375) );
  AOI22_X1 U24316 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n21385), .B1(
        n21384), .B2(n21547), .ZN(n21374) );
  OAI211_X1 U24317 ( .C1(n21550), .C2(n21388), .A(n21375), .B(n21374), .ZN(
        P1_U3076) );
  AOI22_X1 U24318 ( .A1(n21610), .A2(n21383), .B1(n21382), .B2(n21609), .ZN(
        n21377) );
  AOI22_X1 U24319 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n21385), .B1(
        n21384), .B2(n21551), .ZN(n21376) );
  OAI211_X1 U24320 ( .C1(n21554), .C2(n21388), .A(n21377), .B(n21376), .ZN(
        P1_U3077) );
  AOI22_X1 U24321 ( .A1(n21616), .A2(n21383), .B1(n21382), .B2(n21615), .ZN(
        n21379) );
  AOI22_X1 U24322 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n21385), .B1(
        n21384), .B2(n21555), .ZN(n21378) );
  OAI211_X1 U24323 ( .C1(n21558), .C2(n21388), .A(n21379), .B(n21378), .ZN(
        P1_U3078) );
  AOI22_X1 U24324 ( .A1(n21622), .A2(n21383), .B1(n21382), .B2(n21621), .ZN(
        n21381) );
  AOI22_X1 U24325 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n21385), .B1(
        n21384), .B2(n21559), .ZN(n21380) );
  OAI211_X1 U24326 ( .C1(n21562), .C2(n21388), .A(n21381), .B(n21380), .ZN(
        P1_U3079) );
  AOI22_X1 U24327 ( .A1(n21630), .A2(n21383), .B1(n21382), .B2(n21627), .ZN(
        n21387) );
  AOI22_X1 U24328 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n21385), .B1(
        n21384), .B2(n21563), .ZN(n21386) );
  OAI211_X1 U24329 ( .C1(n21570), .C2(n21388), .A(n21387), .B(n21386), .ZN(
        P1_U3080) );
  INV_X1 U24330 ( .A(n21389), .ZN(n21390) );
  NAND2_X1 U24331 ( .A1(n21739), .A2(n21391), .ZN(n21454) );
  NAND2_X1 U24332 ( .A1(n21392), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21495) );
  OR2_X1 U24333 ( .A1(n21522), .A2(n21495), .ZN(n21398) );
  OAI21_X1 U24334 ( .B1(n21454), .B2(n21526), .A(n21398), .ZN(n21400) );
  INV_X1 U24335 ( .A(n21400), .ZN(n21396) );
  NAND2_X1 U24336 ( .A1(n21394), .A2(n21393), .ZN(n21532) );
  OAI22_X1 U24337 ( .A1(n21396), .A2(n21584), .B1(n21395), .B2(n21532), .ZN(
        n21417) );
  INV_X1 U24338 ( .A(n21398), .ZN(n21416) );
  AOI22_X1 U24339 ( .A1(n21417), .A2(n21577), .B1(n21578), .B2(n21416), .ZN(
        n21403) );
  AOI21_X1 U24340 ( .B1(n21449), .B2(n21397), .A(n21426), .ZN(n21401) );
  NAND2_X1 U24341 ( .A1(n21398), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21399) );
  AOI22_X1 U24342 ( .A1(n21419), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n21418), .B2(n21587), .ZN(n21402) );
  OAI211_X1 U24343 ( .C1(n21590), .C2(n21449), .A(n21403), .B(n21402), .ZN(
        P1_U3097) );
  AOI22_X1 U24344 ( .A1(n21417), .A2(n21591), .B1(n21592), .B2(n21416), .ZN(
        n21405) );
  AOI22_X1 U24345 ( .A1(n21419), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n21418), .B2(n21593), .ZN(n21404) );
  OAI211_X1 U24346 ( .C1(n21596), .C2(n21449), .A(n21405), .B(n21404), .ZN(
        P1_U3098) );
  AOI22_X1 U24347 ( .A1(n21417), .A2(n21597), .B1(n21598), .B2(n21416), .ZN(
        n21407) );
  AOI22_X1 U24348 ( .A1(n21419), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n21418), .B2(n21599), .ZN(n21406) );
  OAI211_X1 U24349 ( .C1(n21602), .C2(n21449), .A(n21407), .B(n21406), .ZN(
        P1_U3099) );
  AOI22_X1 U24350 ( .A1(n21417), .A2(n21603), .B1(n21604), .B2(n21416), .ZN(
        n21409) );
  AOI22_X1 U24351 ( .A1(n21419), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n21418), .B2(n21605), .ZN(n21408) );
  OAI211_X1 U24352 ( .C1(n21608), .C2(n21449), .A(n21409), .B(n21408), .ZN(
        P1_U3100) );
  AOI22_X1 U24353 ( .A1(n21417), .A2(n21609), .B1(n21610), .B2(n21416), .ZN(
        n21411) );
  AOI22_X1 U24354 ( .A1(n21419), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n21418), .B2(n21611), .ZN(n21410) );
  OAI211_X1 U24355 ( .C1(n21614), .C2(n21449), .A(n21411), .B(n21410), .ZN(
        P1_U3101) );
  AOI22_X1 U24356 ( .A1(n21417), .A2(n21615), .B1(n21616), .B2(n21416), .ZN(
        n21413) );
  AOI22_X1 U24357 ( .A1(n21419), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n21418), .B2(n21617), .ZN(n21412) );
  OAI211_X1 U24358 ( .C1(n21620), .C2(n21449), .A(n21413), .B(n21412), .ZN(
        P1_U3102) );
  AOI22_X1 U24359 ( .A1(n21417), .A2(n21621), .B1(n21622), .B2(n21416), .ZN(
        n21415) );
  AOI22_X1 U24360 ( .A1(n21419), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n21418), .B2(n21623), .ZN(n21414) );
  OAI211_X1 U24361 ( .C1(n21626), .C2(n21449), .A(n21415), .B(n21414), .ZN(
        P1_U3103) );
  AOI22_X1 U24362 ( .A1(n21417), .A2(n21627), .B1(n21630), .B2(n21416), .ZN(
        n21421) );
  AOI22_X1 U24363 ( .A1(n21419), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n21418), .B2(n21631), .ZN(n21420) );
  OAI211_X1 U24364 ( .C1(n21637), .C2(n21449), .A(n21421), .B(n21420), .ZN(
        P1_U3104) );
  INV_X1 U24365 ( .A(n21454), .ZN(n21496) );
  NOR2_X1 U24366 ( .A1(n21495), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21428) );
  INV_X1 U24367 ( .A(n21428), .ZN(n21424) );
  NOR2_X1 U24368 ( .A1(n21422), .A2(n21424), .ZN(n21444) );
  AOI21_X1 U24369 ( .B1(n21496), .B2(n21423), .A(n21444), .ZN(n21425) );
  OAI22_X1 U24370 ( .A1(n21425), .A2(n21584), .B1(n21424), .B2(n21641), .ZN(
        n21445) );
  AOI22_X1 U24371 ( .A1(n21445), .A2(n21577), .B1(n21578), .B2(n21444), .ZN(
        n21431) );
  OAI21_X1 U24372 ( .B1(n21499), .B2(n21426), .A(n21425), .ZN(n21427) );
  AOI22_X1 U24373 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n21446), .B1(
        n21486), .B2(n21523), .ZN(n21430) );
  OAI211_X1 U24374 ( .C1(n21538), .C2(n21449), .A(n21431), .B(n21430), .ZN(
        P1_U3105) );
  AOI22_X1 U24375 ( .A1(n21445), .A2(n21591), .B1(n21592), .B2(n21444), .ZN(
        n21433) );
  AOI22_X1 U24376 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n21446), .B1(
        n21486), .B2(n21539), .ZN(n21432) );
  OAI211_X1 U24377 ( .C1(n21542), .C2(n21449), .A(n21433), .B(n21432), .ZN(
        P1_U3106) );
  AOI22_X1 U24378 ( .A1(n21445), .A2(n21597), .B1(n21598), .B2(n21444), .ZN(
        n21435) );
  AOI22_X1 U24379 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n21446), .B1(
        n21486), .B2(n21543), .ZN(n21434) );
  OAI211_X1 U24380 ( .C1(n21546), .C2(n21449), .A(n21435), .B(n21434), .ZN(
        P1_U3107) );
  AOI22_X1 U24381 ( .A1(n21445), .A2(n21603), .B1(n21604), .B2(n21444), .ZN(
        n21437) );
  AOI22_X1 U24382 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n21446), .B1(
        n21486), .B2(n21547), .ZN(n21436) );
  OAI211_X1 U24383 ( .C1(n21550), .C2(n21449), .A(n21437), .B(n21436), .ZN(
        P1_U3108) );
  AOI22_X1 U24384 ( .A1(n21445), .A2(n21609), .B1(n21610), .B2(n21444), .ZN(
        n21439) );
  AOI22_X1 U24385 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n21446), .B1(
        n21486), .B2(n21551), .ZN(n21438) );
  OAI211_X1 U24386 ( .C1(n21554), .C2(n21449), .A(n21439), .B(n21438), .ZN(
        P1_U3109) );
  AOI22_X1 U24387 ( .A1(n21445), .A2(n21615), .B1(n21616), .B2(n21444), .ZN(
        n21441) );
  AOI22_X1 U24388 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n21446), .B1(
        n21486), .B2(n21555), .ZN(n21440) );
  OAI211_X1 U24389 ( .C1(n21558), .C2(n21449), .A(n21441), .B(n21440), .ZN(
        P1_U3110) );
  AOI22_X1 U24390 ( .A1(n21445), .A2(n21621), .B1(n21622), .B2(n21444), .ZN(
        n21443) );
  AOI22_X1 U24391 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n21446), .B1(
        n21486), .B2(n21559), .ZN(n21442) );
  OAI211_X1 U24392 ( .C1(n21562), .C2(n21449), .A(n21443), .B(n21442), .ZN(
        P1_U3111) );
  AOI22_X1 U24393 ( .A1(n21445), .A2(n21627), .B1(n21630), .B2(n21444), .ZN(
        n21448) );
  AOI22_X1 U24394 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n21446), .B1(
        n21486), .B2(n21563), .ZN(n21447) );
  OAI211_X1 U24395 ( .C1(n21570), .C2(n21449), .A(n21448), .B(n21447), .ZN(
        P1_U3112) );
  INV_X1 U24396 ( .A(n21486), .ZN(n21450) );
  NAND2_X1 U24397 ( .A1(n21450), .A2(n21586), .ZN(n21452) );
  NOR2_X1 U24398 ( .A1(n21454), .A2(n21453), .ZN(n21457) );
  NOR2_X1 U24399 ( .A1(n21575), .A2(n21495), .ZN(n21501) );
  INV_X1 U24400 ( .A(n21501), .ZN(n21497) );
  NOR2_X1 U24401 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21497), .ZN(
        n21485) );
  AOI22_X1 U24402 ( .A1(n21486), .A2(n21587), .B1(n21485), .B2(n21578), .ZN(
        n21465) );
  INV_X1 U24403 ( .A(n21457), .ZN(n21459) );
  INV_X1 U24404 ( .A(n21485), .ZN(n21458) );
  AOI22_X1 U24405 ( .A1(n21460), .A2(n21459), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21458), .ZN(n21462) );
  NAND3_X1 U24406 ( .A1(n21463), .A2(n21462), .A3(n21461), .ZN(n21487) );
  AOI22_X1 U24407 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n21487), .B1(
        n21518), .B2(n21523), .ZN(n21464) );
  OAI211_X1 U24408 ( .C1(n21491), .C2(n21466), .A(n21465), .B(n21464), .ZN(
        P1_U3113) );
  AOI22_X1 U24409 ( .A1(n21486), .A2(n21593), .B1(n21485), .B2(n21592), .ZN(
        n21468) );
  AOI22_X1 U24410 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n21487), .B1(
        n21518), .B2(n21539), .ZN(n21467) );
  OAI211_X1 U24411 ( .C1(n21491), .C2(n21469), .A(n21468), .B(n21467), .ZN(
        P1_U3114) );
  AOI22_X1 U24412 ( .A1(n21486), .A2(n21599), .B1(n21485), .B2(n21598), .ZN(
        n21471) );
  AOI22_X1 U24413 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n21487), .B1(
        n21518), .B2(n21543), .ZN(n21470) );
  OAI211_X1 U24414 ( .C1(n21491), .C2(n21472), .A(n21471), .B(n21470), .ZN(
        P1_U3115) );
  AOI22_X1 U24415 ( .A1(n21518), .A2(n21547), .B1(n21485), .B2(n21604), .ZN(
        n21474) );
  AOI22_X1 U24416 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n21487), .B1(
        n21486), .B2(n21605), .ZN(n21473) );
  OAI211_X1 U24417 ( .C1(n21491), .C2(n21475), .A(n21474), .B(n21473), .ZN(
        P1_U3116) );
  AOI22_X1 U24418 ( .A1(n21518), .A2(n21551), .B1(n21485), .B2(n21610), .ZN(
        n21477) );
  AOI22_X1 U24419 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n21487), .B1(
        n21486), .B2(n21611), .ZN(n21476) );
  OAI211_X1 U24420 ( .C1(n21491), .C2(n21478), .A(n21477), .B(n21476), .ZN(
        P1_U3117) );
  AOI22_X1 U24421 ( .A1(n21486), .A2(n21617), .B1(n21485), .B2(n21616), .ZN(
        n21480) );
  AOI22_X1 U24422 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n21487), .B1(
        n21518), .B2(n21555), .ZN(n21479) );
  OAI211_X1 U24423 ( .C1(n21491), .C2(n21481), .A(n21480), .B(n21479), .ZN(
        P1_U3118) );
  AOI22_X1 U24424 ( .A1(n21486), .A2(n21623), .B1(n21485), .B2(n21622), .ZN(
        n21483) );
  AOI22_X1 U24425 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n21487), .B1(
        n21518), .B2(n21559), .ZN(n21482) );
  OAI211_X1 U24426 ( .C1(n21491), .C2(n21484), .A(n21483), .B(n21482), .ZN(
        P1_U3119) );
  AOI22_X1 U24427 ( .A1(n21486), .A2(n21631), .B1(n21485), .B2(n21630), .ZN(
        n21489) );
  AOI22_X1 U24428 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n21487), .B1(
        n21518), .B2(n21563), .ZN(n21488) );
  OAI211_X1 U24429 ( .C1(n21491), .C2(n21490), .A(n21489), .B(n21488), .ZN(
        P1_U3120) );
  INV_X1 U24430 ( .A(n21492), .ZN(n21493) );
  NOR2_X1 U24431 ( .A1(n21571), .A2(n21495), .ZN(n21516) );
  AOI21_X1 U24432 ( .B1(n21496), .B2(n21572), .A(n21516), .ZN(n21498) );
  OAI22_X1 U24433 ( .A1(n21498), .A2(n21584), .B1(n21497), .B2(n21641), .ZN(
        n21517) );
  AOI22_X1 U24434 ( .A1(n21517), .A2(n21577), .B1(n21578), .B2(n21516), .ZN(
        n21503) );
  OAI21_X1 U24435 ( .B1(n21499), .B2(n21580), .A(n21498), .ZN(n21500) );
  AOI22_X1 U24436 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n21519), .B1(
        n21518), .B2(n21587), .ZN(n21502) );
  OAI211_X1 U24437 ( .C1(n21590), .C2(n21569), .A(n21503), .B(n21502), .ZN(
        P1_U3121) );
  AOI22_X1 U24438 ( .A1(n21517), .A2(n21591), .B1(n21592), .B2(n21516), .ZN(
        n21505) );
  AOI22_X1 U24439 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n21519), .B1(
        n21518), .B2(n21593), .ZN(n21504) );
  OAI211_X1 U24440 ( .C1(n21596), .C2(n21569), .A(n21505), .B(n21504), .ZN(
        P1_U3122) );
  AOI22_X1 U24441 ( .A1(n21517), .A2(n21597), .B1(n21598), .B2(n21516), .ZN(
        n21507) );
  AOI22_X1 U24442 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n21519), .B1(
        n21518), .B2(n21599), .ZN(n21506) );
  OAI211_X1 U24443 ( .C1(n21602), .C2(n21569), .A(n21507), .B(n21506), .ZN(
        P1_U3123) );
  AOI22_X1 U24444 ( .A1(n21517), .A2(n21603), .B1(n21604), .B2(n21516), .ZN(
        n21509) );
  AOI22_X1 U24445 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n21519), .B1(
        n21518), .B2(n21605), .ZN(n21508) );
  OAI211_X1 U24446 ( .C1(n21608), .C2(n21569), .A(n21509), .B(n21508), .ZN(
        P1_U3124) );
  AOI22_X1 U24447 ( .A1(n21517), .A2(n21609), .B1(n21610), .B2(n21516), .ZN(
        n21511) );
  AOI22_X1 U24448 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n21519), .B1(
        n21518), .B2(n21611), .ZN(n21510) );
  OAI211_X1 U24449 ( .C1(n21614), .C2(n21569), .A(n21511), .B(n21510), .ZN(
        P1_U3125) );
  AOI22_X1 U24450 ( .A1(n21517), .A2(n21615), .B1(n21616), .B2(n21516), .ZN(
        n21513) );
  AOI22_X1 U24451 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n21519), .B1(
        n21518), .B2(n21617), .ZN(n21512) );
  OAI211_X1 U24452 ( .C1(n21620), .C2(n21569), .A(n21513), .B(n21512), .ZN(
        P1_U3126) );
  AOI22_X1 U24453 ( .A1(n21517), .A2(n21621), .B1(n21622), .B2(n21516), .ZN(
        n21515) );
  AOI22_X1 U24454 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n21519), .B1(
        n21518), .B2(n21623), .ZN(n21514) );
  OAI211_X1 U24455 ( .C1(n21626), .C2(n21569), .A(n21515), .B(n21514), .ZN(
        P1_U3127) );
  AOI22_X1 U24456 ( .A1(n21517), .A2(n21627), .B1(n21630), .B2(n21516), .ZN(
        n21521) );
  AOI22_X1 U24457 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n21519), .B1(
        n21518), .B2(n21631), .ZN(n21520) );
  OAI211_X1 U24458 ( .C1(n21637), .C2(n21569), .A(n21521), .B(n21520), .ZN(
        P1_U3128) );
  AOI22_X1 U24459 ( .A1(n21564), .A2(n21523), .B1(n10556), .B2(n21578), .ZN(
        n21537) );
  NAND3_X1 U24460 ( .A1(n21569), .A2(n21586), .A3(n21524), .ZN(n21525) );
  NAND2_X1 U24461 ( .A1(n21525), .A2(n21742), .ZN(n21531) );
  OR2_X1 U24462 ( .A1(n21527), .A2(n21526), .ZN(n21534) );
  AOI22_X1 U24463 ( .A1(n21531), .A2(n21534), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21532), .ZN(n21528) );
  INV_X1 U24464 ( .A(n21531), .ZN(n21535) );
  AOI22_X1 U24465 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n21566), .B1(
        n21577), .B2(n21565), .ZN(n21536) );
  OAI211_X1 U24466 ( .C1(n21538), .C2(n21569), .A(n21537), .B(n21536), .ZN(
        P1_U3129) );
  AOI22_X1 U24467 ( .A1(n21564), .A2(n21539), .B1(n10556), .B2(n21592), .ZN(
        n21541) );
  AOI22_X1 U24468 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n21566), .B1(
        n21591), .B2(n21565), .ZN(n21540) );
  OAI211_X1 U24469 ( .C1(n21542), .C2(n21569), .A(n21541), .B(n21540), .ZN(
        P1_U3130) );
  AOI22_X1 U24470 ( .A1(n21564), .A2(n21543), .B1(n10556), .B2(n21598), .ZN(
        n21545) );
  AOI22_X1 U24471 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n21566), .B1(
        n21597), .B2(n21565), .ZN(n21544) );
  OAI211_X1 U24472 ( .C1(n21546), .C2(n21569), .A(n21545), .B(n21544), .ZN(
        P1_U3131) );
  AOI22_X1 U24473 ( .A1(n21564), .A2(n21547), .B1(n10556), .B2(n21604), .ZN(
        n21549) );
  AOI22_X1 U24474 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n21566), .B1(
        n21603), .B2(n21565), .ZN(n21548) );
  OAI211_X1 U24475 ( .C1(n21550), .C2(n21569), .A(n21549), .B(n21548), .ZN(
        P1_U3132) );
  AOI22_X1 U24476 ( .A1(n21564), .A2(n21551), .B1(n10556), .B2(n21610), .ZN(
        n21553) );
  AOI22_X1 U24477 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n21566), .B1(
        n21609), .B2(n21565), .ZN(n21552) );
  OAI211_X1 U24478 ( .C1(n21554), .C2(n21569), .A(n21553), .B(n21552), .ZN(
        P1_U3133) );
  AOI22_X1 U24479 ( .A1(n21564), .A2(n21555), .B1(n10556), .B2(n21616), .ZN(
        n21557) );
  AOI22_X1 U24480 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n21566), .B1(
        n21615), .B2(n21565), .ZN(n21556) );
  OAI211_X1 U24481 ( .C1(n21558), .C2(n21569), .A(n21557), .B(n21556), .ZN(
        P1_U3134) );
  AOI22_X1 U24482 ( .A1(n21564), .A2(n21559), .B1(n10556), .B2(n21622), .ZN(
        n21561) );
  AOI22_X1 U24483 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n21566), .B1(
        n21621), .B2(n21565), .ZN(n21560) );
  OAI211_X1 U24484 ( .C1(n21562), .C2(n21569), .A(n21561), .B(n21560), .ZN(
        P1_U3135) );
  AOI22_X1 U24485 ( .A1(n21564), .A2(n21563), .B1(n10556), .B2(n21630), .ZN(
        n21568) );
  AOI22_X1 U24486 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n21566), .B1(
        n21627), .B2(n21565), .ZN(n21567) );
  OAI211_X1 U24487 ( .C1(n21570), .C2(n21569), .A(n21568), .B(n21567), .ZN(
        P1_U3136) );
  NOR2_X1 U24488 ( .A1(n21571), .A2(n21574), .ZN(n21629) );
  AOI21_X1 U24489 ( .B1(n21573), .B2(n21572), .A(n21629), .ZN(n21579) );
  NOR2_X1 U24490 ( .A1(n21575), .A2(n21574), .ZN(n21585) );
  INV_X1 U24491 ( .A(n21585), .ZN(n21576) );
  OAI22_X1 U24492 ( .A1(n21579), .A2(n21584), .B1(n21576), .B2(n21641), .ZN(
        n21628) );
  AOI22_X1 U24493 ( .A1(n21578), .A2(n21629), .B1(n21628), .B2(n21577), .ZN(
        n21589) );
  OAI21_X1 U24494 ( .B1(n21581), .B2(n21580), .A(n21579), .ZN(n21583) );
  OAI221_X1 U24495 ( .B1(n21586), .B2(n21585), .C1(n21584), .C2(n21583), .A(
        n21582), .ZN(n21633) );
  AOI22_X1 U24496 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21633), .B1(
        n21632), .B2(n21587), .ZN(n21588) );
  OAI211_X1 U24497 ( .C1(n21590), .C2(n21636), .A(n21589), .B(n21588), .ZN(
        P1_U3153) );
  AOI22_X1 U24498 ( .A1(n21592), .A2(n21629), .B1(n21628), .B2(n21591), .ZN(
        n21595) );
  AOI22_X1 U24499 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21633), .B1(
        n21632), .B2(n21593), .ZN(n21594) );
  OAI211_X1 U24500 ( .C1(n21596), .C2(n21636), .A(n21595), .B(n21594), .ZN(
        P1_U3154) );
  AOI22_X1 U24501 ( .A1(n21598), .A2(n21629), .B1(n21628), .B2(n21597), .ZN(
        n21601) );
  AOI22_X1 U24502 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21633), .B1(
        n21632), .B2(n21599), .ZN(n21600) );
  OAI211_X1 U24503 ( .C1(n21602), .C2(n21636), .A(n21601), .B(n21600), .ZN(
        P1_U3155) );
  AOI22_X1 U24504 ( .A1(n21604), .A2(n21629), .B1(n21628), .B2(n21603), .ZN(
        n21607) );
  AOI22_X1 U24505 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21633), .B1(
        n21632), .B2(n21605), .ZN(n21606) );
  OAI211_X1 U24506 ( .C1(n21608), .C2(n21636), .A(n21607), .B(n21606), .ZN(
        P1_U3156) );
  AOI22_X1 U24507 ( .A1(n21610), .A2(n21629), .B1(n21628), .B2(n21609), .ZN(
        n21613) );
  AOI22_X1 U24508 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21633), .B1(
        n21632), .B2(n21611), .ZN(n21612) );
  OAI211_X1 U24509 ( .C1(n21614), .C2(n21636), .A(n21613), .B(n21612), .ZN(
        P1_U3157) );
  AOI22_X1 U24510 ( .A1(n21616), .A2(n21629), .B1(n21628), .B2(n21615), .ZN(
        n21619) );
  AOI22_X1 U24511 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21633), .B1(
        n21632), .B2(n21617), .ZN(n21618) );
  OAI211_X1 U24512 ( .C1(n21620), .C2(n21636), .A(n21619), .B(n21618), .ZN(
        P1_U3158) );
  AOI22_X1 U24513 ( .A1(n21622), .A2(n21629), .B1(n21628), .B2(n21621), .ZN(
        n21625) );
  AOI22_X1 U24514 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21633), .B1(
        n21632), .B2(n21623), .ZN(n21624) );
  OAI211_X1 U24515 ( .C1(n21626), .C2(n21636), .A(n21625), .B(n21624), .ZN(
        P1_U3159) );
  AOI22_X1 U24516 ( .A1(n21630), .A2(n21629), .B1(n21628), .B2(n21627), .ZN(
        n21635) );
  AOI22_X1 U24517 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21633), .B1(
        n21632), .B2(n21631), .ZN(n21634) );
  OAI211_X1 U24518 ( .C1(n21637), .C2(n21636), .A(n21635), .B(n21634), .ZN(
        P1_U3160) );
  NOR2_X1 U24519 ( .A1(n21638), .A2(n13237), .ZN(n21640) );
  OAI21_X1 U24520 ( .B1(n21641), .B2(n21640), .A(n21639), .ZN(P1_U3163) );
  AND2_X1 U24521 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21726), .ZN(
        P1_U3164) );
  AND2_X1 U24522 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21726), .ZN(
        P1_U3165) );
  AND2_X1 U24523 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21726), .ZN(
        P1_U3166) );
  AND2_X1 U24524 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21726), .ZN(
        P1_U3167) );
  AND2_X1 U24525 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21726), .ZN(
        P1_U3168) );
  AND2_X1 U24526 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21726), .ZN(
        P1_U3169) );
  AND2_X1 U24527 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21726), .ZN(
        P1_U3170) );
  AND2_X1 U24528 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21726), .ZN(
        P1_U3171) );
  AND2_X1 U24529 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21726), .ZN(
        P1_U3172) );
  AND2_X1 U24530 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21726), .ZN(
        P1_U3173) );
  AND2_X1 U24531 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21726), .ZN(
        P1_U3174) );
  AND2_X1 U24532 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21726), .ZN(
        P1_U3175) );
  AND2_X1 U24533 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21726), .ZN(
        P1_U3176) );
  AND2_X1 U24534 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21726), .ZN(
        P1_U3177) );
  AND2_X1 U24535 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21726), .ZN(
        P1_U3178) );
  AND2_X1 U24536 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21726), .ZN(
        P1_U3179) );
  AND2_X1 U24537 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21726), .ZN(
        P1_U3180) );
  NOR2_X1 U24538 ( .A1(n21730), .A2(n21642), .ZN(P1_U3181) );
  NOR2_X1 U24539 ( .A1(n21730), .A2(n21643), .ZN(P1_U3182) );
  AND2_X1 U24540 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21726), .ZN(
        P1_U3183) );
  AND2_X1 U24541 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21726), .ZN(
        P1_U3184) );
  AND2_X1 U24542 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21726), .ZN(
        P1_U3185) );
  AND2_X1 U24543 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21726), .ZN(P1_U3186) );
  AND2_X1 U24544 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21726), .ZN(P1_U3187) );
  AND2_X1 U24545 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21726), .ZN(P1_U3188) );
  AND2_X1 U24546 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21726), .ZN(P1_U3189) );
  AND2_X1 U24547 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21726), .ZN(P1_U3190) );
  AND2_X1 U24548 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21726), .ZN(P1_U3191) );
  AND2_X1 U24549 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21726), .ZN(P1_U3192) );
  AND2_X1 U24550 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21726), .ZN(P1_U3193) );
  AND2_X1 U24551 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21644), .ZN(n21659) );
  INV_X1 U24552 ( .A(n21645), .ZN(n21648) );
  NAND2_X1 U24553 ( .A1(n21657), .A2(NA), .ZN(n21646) );
  OAI211_X1 U24554 ( .C1(n21648), .C2(n21647), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .B(n21646), .ZN(n21649) );
  INV_X1 U24555 ( .A(n21649), .ZN(n21650) );
  OAI22_X1 U24556 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21659), .B1(n21770), 
        .B2(n21650), .ZN(P1_U3194) );
  NAND2_X1 U24557 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21651) );
  OAI21_X1 U24558 ( .B1(NA), .B2(n21651), .A(n12627), .ZN(n21652) );
  OAI21_X1 U24559 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21653), .A(n21652), 
        .ZN(n21658) );
  INV_X1 U24560 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21655) );
  OAI211_X1 U24561 ( .C1(NA), .C2(n21759), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n12627), .ZN(n21654) );
  OAI211_X1 U24562 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21655), .A(HOLD), .B(
        n21654), .ZN(n21656) );
  OAI22_X1 U24563 ( .A1(n21659), .A2(n21658), .B1(n21657), .B2(n21656), .ZN(
        P1_U3196) );
  NAND2_X1 U24564 ( .A1(n21770), .A2(n12627), .ZN(n21714) );
  NAND2_X1 U24565 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21770), .ZN(n21718) );
  OAI222_X1 U24566 ( .A1(n21714), .A2(n21663), .B1(n21661), .B2(n21770), .C1(
        n21660), .C2(n21718), .ZN(P1_U3197) );
  INV_X1 U24567 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n21662) );
  OAI222_X1 U24568 ( .A1(n21718), .A2(n21663), .B1(n21662), .B2(n21770), .C1(
        n21665), .C2(n21714), .ZN(P1_U3198) );
  INV_X1 U24569 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21664) );
  OAI222_X1 U24570 ( .A1(n21718), .A2(n21665), .B1(n21664), .B2(n21770), .C1(
        n21667), .C2(n21714), .ZN(P1_U3199) );
  INV_X1 U24571 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21670) );
  OAI222_X1 U24572 ( .A1(n21718), .A2(n21667), .B1(n21666), .B2(n21770), .C1(
        n21670), .C2(n21714), .ZN(P1_U3200) );
  INV_X1 U24573 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n21669) );
  OAI222_X1 U24574 ( .A1(n21718), .A2(n21670), .B1(n21669), .B2(n21770), .C1(
        n21668), .C2(n21714), .ZN(P1_U3201) );
  INV_X1 U24575 ( .A(n21718), .ZN(n21709) );
  INV_X1 U24576 ( .A(n21714), .ZN(n21711) );
  AOI222_X1 U24577 ( .A1(n21709), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n21755), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n21711), .ZN(n21671) );
  INV_X1 U24578 ( .A(n21671), .ZN(P1_U3202) );
  OAI222_X1 U24579 ( .A1(n21718), .A2(n21673), .B1(n21672), .B2(n21770), .C1(
        n21674), .C2(n21714), .ZN(P1_U3203) );
  INV_X1 U24580 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n21675) );
  OAI222_X1 U24581 ( .A1(n21714), .A2(n21677), .B1(n21675), .B2(n21770), .C1(
        n21674), .C2(n21718), .ZN(P1_U3204) );
  AOI22_X1 U24582 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n21755), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n21711), .ZN(n21676) );
  OAI21_X1 U24583 ( .B1(n21677), .B2(n21718), .A(n21676), .ZN(P1_U3205) );
  AOI22_X1 U24584 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n21755), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n21709), .ZN(n21678) );
  OAI21_X1 U24585 ( .B1(n21680), .B2(n21714), .A(n21678), .ZN(P1_U3206) );
  AOI22_X1 U24586 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n21755), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n21711), .ZN(n21679) );
  OAI21_X1 U24587 ( .B1(n21680), .B2(n21718), .A(n21679), .ZN(P1_U3207) );
  AOI22_X1 U24588 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n21755), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n21709), .ZN(n21681) );
  OAI21_X1 U24589 ( .B1(n21684), .B2(n21714), .A(n21681), .ZN(P1_U3208) );
  INV_X1 U24590 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n21683) );
  OAI222_X1 U24591 ( .A1(n21718), .A2(n21684), .B1(n21683), .B2(n21770), .C1(
        n21682), .C2(n21714), .ZN(P1_U3209) );
  AOI222_X1 U24592 ( .A1(n21711), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n21755), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n21709), .ZN(n21685) );
  INV_X1 U24593 ( .A(n21685), .ZN(P1_U3210) );
  AOI222_X1 U24594 ( .A1(n21709), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n21755), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n21711), .ZN(n21686) );
  INV_X1 U24595 ( .A(n21686), .ZN(P1_U3211) );
  INV_X1 U24596 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n21687) );
  OAI222_X1 U24597 ( .A1(n21718), .A2(n21688), .B1(n21687), .B2(n21770), .C1(
        n21690), .C2(n21714), .ZN(P1_U3212) );
  AOI22_X1 U24598 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n21755), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n21711), .ZN(n21689) );
  OAI21_X1 U24599 ( .B1(n21690), .B2(n21718), .A(n21689), .ZN(P1_U3213) );
  AOI22_X1 U24600 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n21755), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n21709), .ZN(n21691) );
  OAI21_X1 U24601 ( .B1(n21693), .B2(n21714), .A(n21691), .ZN(P1_U3214) );
  AOI22_X1 U24602 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n21755), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n21711), .ZN(n21692) );
  OAI21_X1 U24603 ( .B1(n21693), .B2(n21718), .A(n21692), .ZN(P1_U3215) );
  INV_X1 U24604 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21695) );
  OAI222_X1 U24605 ( .A1(n21718), .A2(n21695), .B1(n21694), .B2(n21770), .C1(
        n21697), .C2(n21714), .ZN(P1_U3216) );
  INV_X1 U24606 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n21696) );
  OAI222_X1 U24607 ( .A1(n21718), .A2(n21697), .B1(n21696), .B2(n21770), .C1(
        n21699), .C2(n21714), .ZN(P1_U3217) );
  AOI22_X1 U24608 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n21755), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21711), .ZN(n21698) );
  OAI21_X1 U24609 ( .B1(n21699), .B2(n21718), .A(n21698), .ZN(P1_U3218) );
  AOI22_X1 U24610 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n21755), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21709), .ZN(n21700) );
  OAI21_X1 U24611 ( .B1(n21702), .B2(n21714), .A(n21700), .ZN(P1_U3219) );
  INV_X1 U24612 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n21701) );
  OAI222_X1 U24613 ( .A1(n21718), .A2(n21702), .B1(n21701), .B2(n21770), .C1(
        n21704), .C2(n21714), .ZN(P1_U3220) );
  INV_X1 U24614 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n21703) );
  OAI222_X1 U24615 ( .A1(n21718), .A2(n21704), .B1(n21703), .B2(n21716), .C1(
        n21706), .C2(n21714), .ZN(P1_U3221) );
  INV_X1 U24616 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n21705) );
  OAI222_X1 U24617 ( .A1(n21718), .A2(n21706), .B1(n21705), .B2(n21716), .C1(
        n21708), .C2(n21714), .ZN(P1_U3222) );
  AOI22_X1 U24618 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n21711), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21755), .ZN(n21707) );
  OAI21_X1 U24619 ( .B1(n21708), .B2(n21718), .A(n21707), .ZN(P1_U3223) );
  AOI22_X1 U24620 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n21709), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21755), .ZN(n21710) );
  OAI21_X1 U24621 ( .B1(n21713), .B2(n21714), .A(n21710), .ZN(P1_U3224) );
  AOI22_X1 U24622 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n21711), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21755), .ZN(n21712) );
  OAI21_X1 U24623 ( .B1(n21713), .B2(n21718), .A(n21712), .ZN(P1_U3225) );
  OAI222_X1 U24624 ( .A1(n21718), .A2(n15449), .B1(n21717), .B2(n21716), .C1(
        n21715), .C2(n21714), .ZN(P1_U3226) );
  INV_X1 U24625 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n21719) );
  AOI22_X1 U24626 ( .A1(n21770), .A2(n21720), .B1(n21719), .B2(n21755), .ZN(
        P1_U3458) );
  INV_X1 U24627 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21749) );
  AOI22_X1 U24628 ( .A1(n21770), .A2(n21749), .B1(n21721), .B2(n21755), .ZN(
        P1_U3459) );
  INV_X1 U24629 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n21722) );
  AOI22_X1 U24630 ( .A1(n21770), .A2(n21723), .B1(n21722), .B2(n21755), .ZN(
        P1_U3460) );
  INV_X1 U24631 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21752) );
  INV_X1 U24632 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n21724) );
  AOI22_X1 U24633 ( .A1(n21770), .A2(n21752), .B1(n21724), .B2(n21755), .ZN(
        P1_U3461) );
  INV_X1 U24634 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21727) );
  INV_X1 U24635 ( .A(n21728), .ZN(n21725) );
  AOI21_X1 U24636 ( .B1(n21727), .B2(n21726), .A(n21725), .ZN(P1_U3464) );
  OAI21_X1 U24637 ( .B1(n21730), .B2(n21729), .A(n21728), .ZN(P1_U3465) );
  AOI22_X1 U24638 ( .A1(n21734), .A2(n21733), .B1(n21732), .B2(n21731), .ZN(
        n21735) );
  INV_X1 U24639 ( .A(n21735), .ZN(n21738) );
  MUX2_X1 U24640 ( .A(n21738), .B(n21737), .S(n21736), .Z(P1_U3469) );
  INV_X1 U24641 ( .A(n21739), .ZN(n21741) );
  OAI22_X1 U24642 ( .A1(n21743), .A2(n21742), .B1(n21741), .B2(n21740), .ZN(
        n21744) );
  OAI21_X1 U24643 ( .B1(n21745), .B2(n21744), .A(n21747), .ZN(n21746) );
  OAI21_X1 U24644 ( .B1(n21747), .B2(n12902), .A(n21746), .ZN(P1_U3475) );
  AOI211_X1 U24645 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_REIP_REG_1__SCAN_IN), .B(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21748) );
  AOI21_X1 U24646 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n21748), .ZN(n21750) );
  AOI22_X1 U24647 ( .A1(n21754), .A2(n21750), .B1(n21749), .B2(n21751), .ZN(
        P1_U3481) );
  NOR2_X1 U24648 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n21753) );
  AOI22_X1 U24649 ( .A1(n21754), .A2(n21753), .B1(n21752), .B2(n21751), .ZN(
        P1_U3482) );
  AOI22_X1 U24650 ( .A1(n21770), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21756), 
        .B2(n21755), .ZN(P1_U3483) );
  AOI211_X1 U24651 ( .C1(n21760), .C2(n21759), .A(n21758), .B(n21757), .ZN(
        n21769) );
  INV_X1 U24652 ( .A(n21761), .ZN(n21764) );
  INV_X1 U24653 ( .A(n21762), .ZN(n21763) );
  OAI211_X1 U24654 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21764), .A(n21763), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21766) );
  AOI21_X1 U24655 ( .B1(n21766), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n21765), 
        .ZN(n21768) );
  NAND2_X1 U24656 ( .A1(n21769), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21767) );
  OAI21_X1 U24657 ( .B1(n21769), .B2(n21768), .A(n21767), .ZN(P1_U3485) );
  MUX2_X1 U24658 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n21770), .Z(P1_U3486) );
  AND2_X2 U11507 ( .A1(n13404), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11682) );
  NAND2_X2 U11914 ( .A1(n11865), .A2(n17662), .ZN(n17644) );
  NAND2_X2 U11243 ( .A1(n18798), .A2(n18799), .ZN(n10152) );
  XNOR2_X1 U11442 ( .A(n13458), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13448) );
  AND2_X2 U11512 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10249) );
  AND2_X1 U11213 ( .A1(n14304), .A2(n10275), .ZN(n12605) );
  AND2_X2 U13380 ( .A1(n10697), .A2(n14353), .ZN(n12340) );
  AND2_X2 U11503 ( .A1(n12324), .A2(n14353), .ZN(n10849) );
  XNOR2_X1 U13000 ( .A(n11572), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15422) );
  AND2_X2 U13729 ( .A1(n12317), .A2(n14353), .ZN(n10625) );
  AND2_X2 U13714 ( .A1(n12316), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10619) );
  NAND2_X2 U12964 ( .A1(n11575), .A2(n11574), .ZN(n10322) );
  AND4_X1 U11158 ( .A1(n12524), .A2(n12523), .A3(n12522), .A4(n12521), .ZN(
        n12525) );
  NOR2_X1 U11159 ( .A1(n11602), .A2(n10345), .ZN(n11157) );
  CLKBUF_X1 U11180 ( .A(n10574), .Z(n14337) );
  INV_X2 U11183 ( .A(n11725), .ZN(n18464) );
  CLKBUF_X1 U11192 ( .A(n13345), .Z(n17755) );
  NOR2_X1 U11219 ( .A1(n11632), .A2(n16412), .ZN(n11631) );
  NOR2_X1 U11273 ( .A1(n11580), .A2(n11579), .ZN(n11578) );
  CLKBUF_X1 U11355 ( .A(n11092), .Z(n11120) );
  NOR2_X1 U11460 ( .A1(n11614), .A2(n17813), .ZN(n11618) );
  AND2_X1 U11467 ( .A1(n10249), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n18409) );
  AOI211_X1 U11494 ( .C1(P1_EBX_REG_18__SCAN_IN), .C2(n21040), .A(n15634), .B(
        n15633), .ZN(n15635) );
  CLKBUF_X2 U11505 ( .A(n13113), .Z(n13610) );
  CLKBUF_X1 U11511 ( .A(n14438), .Z(n21186) );
  AND4_X1 U11515 ( .A1(n10714), .A2(n10720), .A3(n10715), .A4(n10716), .ZN(
        n11184) );
  AND3_X1 U11532 ( .A1(n11715), .A2(n11714), .A3(n11712), .ZN(n10107) );
  NAND2_X1 U11601 ( .A1(n18914), .A2(n18950), .ZN(n18830) );
  CLKBUF_X1 U11609 ( .A(n15419), .Z(n15873) );
  OAI21_X1 U11645 ( .B1(n16442), .B2(n20147), .A(n16924), .ZN(n16414) );
  INV_X1 U11661 ( .A(n10726), .ZN(n12494) );
  XNOR2_X1 U11694 ( .A(n10940), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17140) );
  CLKBUF_X1 U12251 ( .A(n21716), .Z(n21770) );
  INV_X1 U12402 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13404) );
endmodule

